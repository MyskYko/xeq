//
// Conformal-LEC Version 20.10-d131 (29-Jun-2020)
//
module top(RIc0d9478_65,RIc0d7678_1,RIc0d76f0_2,RIc0d7768_3,RIc0d94f0_66,RIc0d77e0_4,RIc0d7858_5,RIc0d9568_67,RIc0d95e0_68,
        RIc0d78d0_6,RIc0d7948_7,RIc0d9658_69,RIc0d96d0_70,RIc0d79c0_8,RIc0d7a38_9,RIc0d9748_71,RIc0d97c0_72,RIc0d7ab0_10,RIc0d7b28_11,
        RIc0d9838_73,RIc0d98b0_74,RIc0d7ba0_12,RIc0d7c18_13,RIc0d9928_75,RIc0d99a0_76,RIc0d7c90_14,RIc0d7d08_15,RIc0d9a18_77,RIc0d9a90_78,
        RIc0d7d80_16,RIc0d7df8_17,RIc0d9b08_79,RIc0d9b80_80,RIc0d7e70_18,RIc0d7ee8_19,RIc0d9bf8_81,RIc0d7f60_20,RIc0d7fd8_21,RIc0d9c70_82,
        RIc0d9ce8_83,RIc0d9d60_84,RIc0d8050_22,RIc0d80c8_23,RIc0d9dd8_85,RIc0d9e50_86,RIc0d8140_24,RIc0d81b8_25,RIc0d9ec8_87,RIc0d9f40_88,
        RIc0d8230_26,RIc0d82a8_27,RIc0d9fb8_89,RIc0da030_90,RIc0d8320_28,RIc0d8398_29,RIc0da0a8_91,RIc0da120_92,RIc0d8410_30,RIc0d8488_31,
        RIc0da198_93,RIc0da210_94,RIc0d8500_32,RIc0d8578_33,RIc0da288_95,RIc0da300_96,RIc0d85f0_34,RIc0d8668_35,RIc0da378_97,RIc0da3f0_98,
        RIc0d86e0_36,RIc0d8758_37,RIc0da468_99,RIc0d87d0_38,RIc0d8848_39,RIc0da4e0_100,RIc0da558_101,RIc0da5d0_102,RIc0d88c0_40,RIc0d8938_41,
        RIc0da648_103,RIc0da6c0_104,RIc0d89b0_42,RIc0d8a28_43,RIc0da738_105,RIc0da7b0_106,RIc0d8aa0_44,RIc0d8b18_45,RIc0da828_107,RIc0da8a0_108,
        RIc0d8b90_46,RIc0d8c08_47,RIc0da918_109,RIc0da990_110,RIc0d8c80_48,RIc0d8cf8_49,RIc0daa08_111,RIc0daa80_112,RIc0d8d70_50,RIc0d8de8_51,
        RIc0daaf8_113,RIc0dab70_114,RIc0d8e60_52,RIc0d8ed8_53,RIc0dabe8_115,RIc0dac60_116,RIc0d8f50_54,RIc0d8fc8_55,RIc0dacd8_117,RIc0d9040_56,
        RIc0d90b8_57,RIc0dad50_118,RIc0dadc8_119,RIc0dae40_120,RIc0d9130_58,RIc0d91a8_59,RIc0daeb8_121,RIc0daf30_122,RIc0d9220_60,RIc0d9298_61,
        RIc0dafa8_123,RIc0db020_124,RIc0d9310_62,RIc0d9388_63,RIc0db098_125,RIc0db110_126,RIc0db188_127,RIc0d9400_64,RIc0db200_128,R_81_84446b8,
        R_82_8444760,R_83_8444808,R_84_84448b0,R_85_8444958,R_86_8444a00,R_87_9bec6f8,R_88_9bec7a0,R_89_9bec848,R_8a_9bec8f0,R_8b_9bec998,
        R_8c_9beca40,R_8d_9becae8,R_8e_9becb90,R_8f_9becc38,R_90_9becce0,R_91_9becd88,R_92_9bece30,R_93_9beced8,R_94_9becf80,R_95_9bed028,
        R_96_9bed0d0,R_97_9bed178,R_98_9bed220,R_99_9bed2c8,R_9a_9bed370,R_9b_9bed418,R_9c_9bed4c0,R_9d_9bed568,R_9e_9bed610,R_9f_9bed6b8,
        R_a0_9bed760,R_a1_9bed808,R_a2_9bed8b0,R_a3_9bed958,R_a4_9beda00,R_a5_9bedaa8,R_a6_9bedb50,R_a7_9bedbf8,R_a8_9bedca0,R_a9_9bedd48,
        R_aa_9beddf0,R_ab_9bede98,R_ac_9bedf40,R_ad_9bedfe8,R_ae_9bee090,R_af_9bee138,R_b0_9bee1e0,R_b1_9bee288,R_b2_9bee330,R_b3_9bee3d8,
        R_b4_9bee480,R_b5_9bee528,R_b6_9bee5d0,R_b7_9bee678,R_b8_9bee720,R_b9_9bee7c8,R_ba_9bee870,R_bb_9bee918,R_bc_9bee9c0,R_bd_9beea68,
        R_be_9beeb10,R_bf_9beebb8,R_c0_9beec60,R_c1_9beed08,R_c2_9beedb0,R_c3_9beee58,R_c4_9beef00,R_c5_9beefa8,R_c6_9bef050,R_c7_9bef0f8,
        R_c8_9bef1a0,R_c9_9bef248,R_ca_9bef2f0,R_cb_9bef398,R_cc_9bef440,R_cd_9bef4e8,R_ce_9bef590,R_cf_9bef638,R_d0_9bef6e0,R_d1_9bef788,
        R_d2_9bef830,R_d3_9bef8d8,R_d4_9bef980,R_d5_9befa28,R_d6_9befad0,R_d7_9befb78,R_d8_9befc20,R_d9_9befcc8,R_da_9befd70,R_db_9befe18,
        R_dc_9befec0,R_dd_9beff68,R_de_9bf0010,R_df_9bf00b8,R_e0_9bf0160,R_e1_9bf0208,R_e2_9bf02b0,R_e3_9bf0358,R_e4_9bf0400,R_e5_9bf04a8,
        R_e6_9bf0550,R_e7_9bf05f8,R_e8_9bf06a0,R_e9_9bf0748,R_ea_9bf07f0,R_eb_9bf0898,R_ec_9bf0940,R_ed_9bf09e8,R_ee_9bf0a90,R_ef_9bf0b38,
        R_f0_9bf0be0,R_f1_9bf0c88,R_f2_9bf0d30,R_f3_9bf0dd8);
input RIc0d9478_65,RIc0d7678_1,RIc0d76f0_2,RIc0d7768_3,RIc0d94f0_66,RIc0d77e0_4,RIc0d7858_5,RIc0d9568_67,RIc0d95e0_68,
        RIc0d78d0_6,RIc0d7948_7,RIc0d9658_69,RIc0d96d0_70,RIc0d79c0_8,RIc0d7a38_9,RIc0d9748_71,RIc0d97c0_72,RIc0d7ab0_10,RIc0d7b28_11,
        RIc0d9838_73,RIc0d98b0_74,RIc0d7ba0_12,RIc0d7c18_13,RIc0d9928_75,RIc0d99a0_76,RIc0d7c90_14,RIc0d7d08_15,RIc0d9a18_77,RIc0d9a90_78,
        RIc0d7d80_16,RIc0d7df8_17,RIc0d9b08_79,RIc0d9b80_80,RIc0d7e70_18,RIc0d7ee8_19,RIc0d9bf8_81,RIc0d7f60_20,RIc0d7fd8_21,RIc0d9c70_82,
        RIc0d9ce8_83,RIc0d9d60_84,RIc0d8050_22,RIc0d80c8_23,RIc0d9dd8_85,RIc0d9e50_86,RIc0d8140_24,RIc0d81b8_25,RIc0d9ec8_87,RIc0d9f40_88,
        RIc0d8230_26,RIc0d82a8_27,RIc0d9fb8_89,RIc0da030_90,RIc0d8320_28,RIc0d8398_29,RIc0da0a8_91,RIc0da120_92,RIc0d8410_30,RIc0d8488_31,
        RIc0da198_93,RIc0da210_94,RIc0d8500_32,RIc0d8578_33,RIc0da288_95,RIc0da300_96,RIc0d85f0_34,RIc0d8668_35,RIc0da378_97,RIc0da3f0_98,
        RIc0d86e0_36,RIc0d8758_37,RIc0da468_99,RIc0d87d0_38,RIc0d8848_39,RIc0da4e0_100,RIc0da558_101,RIc0da5d0_102,RIc0d88c0_40,RIc0d8938_41,
        RIc0da648_103,RIc0da6c0_104,RIc0d89b0_42,RIc0d8a28_43,RIc0da738_105,RIc0da7b0_106,RIc0d8aa0_44,RIc0d8b18_45,RIc0da828_107,RIc0da8a0_108,
        RIc0d8b90_46,RIc0d8c08_47,RIc0da918_109,RIc0da990_110,RIc0d8c80_48,RIc0d8cf8_49,RIc0daa08_111,RIc0daa80_112,RIc0d8d70_50,RIc0d8de8_51,
        RIc0daaf8_113,RIc0dab70_114,RIc0d8e60_52,RIc0d8ed8_53,RIc0dabe8_115,RIc0dac60_116,RIc0d8f50_54,RIc0d8fc8_55,RIc0dacd8_117,RIc0d9040_56,
        RIc0d90b8_57,RIc0dad50_118,RIc0dadc8_119,RIc0dae40_120,RIc0d9130_58,RIc0d91a8_59,RIc0daeb8_121,RIc0daf30_122,RIc0d9220_60,RIc0d9298_61,
        RIc0dafa8_123,RIc0db020_124,RIc0d9310_62,RIc0d9388_63,RIc0db098_125,RIc0db110_126,RIc0db188_127,RIc0d9400_64,RIc0db200_128;
output R_81_84446b8,R_82_8444760,R_83_8444808,R_84_84448b0,R_85_8444958,R_86_8444a00,R_87_9bec6f8,R_88_9bec7a0,R_89_9bec848,
        R_8a_9bec8f0,R_8b_9bec998,R_8c_9beca40,R_8d_9becae8,R_8e_9becb90,R_8f_9becc38,R_90_9becce0,R_91_9becd88,R_92_9bece30,R_93_9beced8,
        R_94_9becf80,R_95_9bed028,R_96_9bed0d0,R_97_9bed178,R_98_9bed220,R_99_9bed2c8,R_9a_9bed370,R_9b_9bed418,R_9c_9bed4c0,R_9d_9bed568,
        R_9e_9bed610,R_9f_9bed6b8,R_a0_9bed760,R_a1_9bed808,R_a2_9bed8b0,R_a3_9bed958,R_a4_9beda00,R_a5_9bedaa8,R_a6_9bedb50,R_a7_9bedbf8,
        R_a8_9bedca0,R_a9_9bedd48,R_aa_9beddf0,R_ab_9bede98,R_ac_9bedf40,R_ad_9bedfe8,R_ae_9bee090,R_af_9bee138,R_b0_9bee1e0,R_b1_9bee288,
        R_b2_9bee330,R_b3_9bee3d8,R_b4_9bee480,R_b5_9bee528,R_b6_9bee5d0,R_b7_9bee678,R_b8_9bee720,R_b9_9bee7c8,R_ba_9bee870,R_bb_9bee918,
        R_bc_9bee9c0,R_bd_9beea68,R_be_9beeb10,R_bf_9beebb8,R_c0_9beec60,R_c1_9beed08,R_c2_9beedb0,R_c3_9beee58,R_c4_9beef00,R_c5_9beefa8,
        R_c6_9bef050,R_c7_9bef0f8,R_c8_9bef1a0,R_c9_9bef248,R_ca_9bef2f0,R_cb_9bef398,R_cc_9bef440,R_cd_9bef4e8,R_ce_9bef590,R_cf_9bef638,
        R_d0_9bef6e0,R_d1_9bef788,R_d2_9bef830,R_d3_9bef8d8,R_d4_9bef980,R_d5_9befa28,R_d6_9befad0,R_d7_9befb78,R_d8_9befc20,R_d9_9befcc8,
        R_da_9befd70,R_db_9befe18,R_dc_9befec0,R_dd_9beff68,R_de_9bf0010,R_df_9bf00b8,R_e0_9bf0160,R_e1_9bf0208,R_e2_9bf02b0,R_e3_9bf0358,
        R_e4_9bf0400,R_e5_9bf04a8,R_e6_9bf0550,R_e7_9bf05f8,R_e8_9bf06a0,R_e9_9bf0748,R_ea_9bf07f0,R_eb_9bf0898,R_ec_9bf0940,R_ed_9bf09e8,
        R_ee_9bf0a90,R_ef_9bf0b38,R_f0_9bf0be0,R_f1_9bf0c88,R_f2_9bf0d30,R_f3_9bf0dd8;

wire \244 , \245 , \246 , \247 , \248 , \249 , \250 , \251 , \252 ,
         \253 , \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 , \262 ,
         \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 , \272 ,
         \273 , \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 , \282 ,
         \283 , \284 , \285 , \286 , \287 , \288 , \289 , \290 , \291 , \292 ,
         \293 , \294 , \295 , \296 , \297 , \298 , \299 , \300 , \301 , \302 ,
         \303 , \304 , \305 , \306 , \307 , \308 , \309 , \310 , \311 , \312 ,
         \313 , \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321 , \322 ,
         \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331 , \332 ,
         \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 , \342 ,
         \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 , \351 , \352 ,
         \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 , \362 ,
         \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 ,
         \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 ,
         \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 ,
         \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 ,
         \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 ,
         \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 ,
         \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 ,
         \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 ,
         \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 ,
         \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 ,
         \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 ,
         \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 ,
         \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 ,
         \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 ,
         \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 ,
         \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 ,
         \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 ,
         \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 ,
         \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 ,
         \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 ,
         \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 ,
         \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 ,
         \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 ,
         \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 ,
         \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612_N$1 ,
         \613_N$2 , \614_N$3 , \615_N$4 , \616_N$5 , \617_N$6 , \618_N$7 , \619_N$8 , \620_N$9 , \621_N$10 , \622_N$11 ,
         \623_N$12 , \624_N$13 , \625_N$14 , \626_N$15 , \627_N$16 , \628_N$17 , \629_N$18 , \630_N$19 , \631_N$20 , \632_N$21 ,
         \633_N$22 , \634_N$23 , \635_N$24 , \636_N$25 , \637_N$26 , \638_N$27 , \639_N$28 , \640_N$29 , \641_N$30 , \642_N$31 ,
         \643_N$32 , \644_N$33 , \645_N$34 , \646_N$35 , \647_N$36 , \648_N$37 , \649_N$38 , \650_N$39 , \651_N$40 , \652_N$41 ,
         \653_N$42 , \654_N$43 , \655_N$44 , \656_N$45 , \657_N$46 , \658_N$47 , \659_N$48 , \660_N$49 , \661_N$50 , \662_N$51 ,
         \663_N$52 , \664_N$53 , \665_N$54 , \666_N$55 , \667_N$56 , \668_N$57 , \669_N$58 , \670_N$59 , \671_N$60 , \672_N$61 ,
         \673_N$62 , \674_N$63 , \675_N$64 , \676_N$65 , \677_N$66 , \678_N$67 , \679_N$68 , \680_N$69 , \681_N$70 , \682_N$71 ,
         \683_N$72 , \684_N$73 , \685_N$74 , \686_N$75 , \687_N$76 , \688_N$77 , \689_N$78 , \690_N$79 , \691_N$80 , \692_N$81 ,
         \693_N$82 , \694_N$83 , \695_N$84 , \696_N$85 , \697_N$86 , \698_N$87 , \699_N$88 , \700_N$89 , \701_N$90 , \702_N$91 ,
         \703_N$92 , \704_N$93 , \705_N$94 , \706_N$95 , \707_N$96 , \708_N$97 , \709_N$98 , \710_N$99 , \711_N$100 , \712_N$101 ,
         \713_N$102 , \714_N$103 , \715_N$104 , \716_N$105 , \717_N$106 , \718_N$107 , \719_N$108 , \720_N$109 , \721_N$110 , \722_N$111 ,
         \723_N$112 , \724_N$113 , \725_N$114 , \726_N$116 , \727_N$117 , \728_N$118 , \729_N$119 , \730_N$120 , \731_N$121 , \732_N$122 ,
         \733_N$123 , \734_N$124 , \735_N$125 , \736_N$126 , \737_N$127 , \738_N$128 , \739_N$129 , \740_N$130 , \741_N$131 , \742_N$132 ,
         \743_N$133 , \744_N$134 , \745_N$135 , \746_N$136 , \747_N$137 , \748_N$138 , \749_N$139 , \750_N$140 , \751_N$141 , \752_N$142 ,
         \753_N$143 , \754_N$144 , \755_N$145 , \756_N$146 , \757_N$147 , \758_N$148 , \759_N$149 , \760_N$150 , \761_N$151 , \762_N$152 ,
         \763_N$153 , \764_N$154 , \765_N$155 , \766_N$156 , \767_N$157 , \768_N$158 , \769_N$159 , \770_N$160 , \771_N$161 , \772_N$162 ,
         \773_N$163 , \774_N$164 , \775_N$165 , \776_N$166 , \777_N$167 , \778_N$168 , \779_N$169 , \780_N$170 , \781_N$171 , \782_N$172 ,
         \783_N$173 , \784_N$174 , \785_N$175 , \786_N$176 , \787_N$177 , \788_N$178 , \789_N$179 , \790_N$180 , \791_N$181 , \792_N$182 ,
         \793_N$183 , \794_N$184 , \795_N$185 , \796_N$186 , \797_N$187 , \798_N$188 , \799_N$189 , \800_N$190 , \801_N$191 , \802_N$192 ,
         \803_N$193 , \804_N$194 , \805_N$195 , \806_N$196 , \807_N$197 , \808_N$198 , \809_N$199 , \810_N$200 , \811_N$201 , \812_N$202 ,
         \813_N$203 , \814_N$204 , \815_N$205 , \816_N$206 , \817_N$207 , \818_N$208 , \819_N$209 , \820_N$210 , \821_N$211 , \822_N$212 ,
         \823_N$213 , \824_N$214 , \825_N$215 , \826_N$216 , \827_N$217 , \828_N$218 , \829_N$219 , \830_N$220 , \831_N$221 , \832_N$222 ,
         \833_N$223 , \834_N$224 , \835_N$225 , \836_N$226 , \837_N$227 , \838_N$228 , \839_N$229 , \840_N$230 , \841_N$231 , \842_N$232 ,
         \843_N$233 , \844_N$234 , \845_N$235 , \846_N$236 , \847_N$237 , \848_N$238 , \849_N$239 , \850_N$240 , \851_N$241 , \852_N$242 ,
         \853_N$243 , \854_N$244 , \855_N$245 , \856_N$246 , \857_N$247 , \858_N$248 , \859_N$249 , \860_N$250 , \861_N$251 , \862_N$252 ,
         \863_N$253 , \864_N$254 , \865_N$255 , \866_N$256 , \867_N$257 , \868_N$258 , \869_N$259 , \870_N$260 , \871_N$261 , \872_N$262 ,
         \873_N$263 , \874_N$264 , \875_N$265 , \876_N$266 , \877_N$267 , \878_N$268 , \879_N$269 , \880_N$270 , \881_N$271 , \882_N$272 ,
         \883_N$273 , \884_N$274 , \885_N$275 , \886_N$276 , \887_N$277 , \888_N$278 , \889_N$279 , \890_N$280 , \891_N$281 , \892_N$282 ,
         \893_N$283 , \894_N$284 , \895_N$285 , \896_N$286 , \897_N$287 , \898_N$288 , \899_N$289 , \900_N$290 , \901_N$291 , \902_N$292 ,
         \903_N$293 , \904_N$294 , \905_N$295 , \906_N$296 , \907_N$297 , \908_N$298 , \909_N$299 , \910_N$300 , \911_N$301 , \912_N$302 ,
         \913_N$303 , \914_N$304 , \915_N$305 , \916_N$306 , \917_N$307 , \918_N$308 , \919_N$309 , \920_N$310 , \921_N$311 , \922_N$312 ,
         \923_N$313 , \924_N$314 , \925_N$315 , \926_N$316 , \927_N$317 , \928_N$318 , \929_N$319 , \930_N$320 , \931_N$321 , \932_N$322 ,
         \933_N$323 , \934_N$324 , \935_N$325 , \936_N$326 , \937_N$327 , \938_N$328 , \939_N$329 , \940_N$330 , \941_N$331 , \942_N$332 ,
         \943_N$333 , \944_N$334 , \945_N$335 , \946_N$336 , \947_N$337 , \948_N$338 , \949_N$339 , \950_N$340 , \951_N$341 , \952_N$342 ,
         \953_N$343 , \954_N$344 , \955_N$345 , \956_N$346 , \957_N$347 , \958_N$348 , \959_N$349 , \960_N$350 , \961_N$351 , \962_N$352 ,
         \963_N$353 , \964_N$354 , \965_N$355 , \966_N$356 , \967_N$357 , \968_N$358 , \969_N$359 , \970_N$360 , \971_N$361 , \972_N$362 ,
         \973_N$363 , \974_N$364 , \975_N$365 , \976_N$366 , \977_N$367 , \978_N$368 , \979_N$369 , \980_ZERO , \981 , \982_N$115 ,
         \983_ONE , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 ,
         \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 ,
         \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 ,
         \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 ,
         \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 ,
         \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 ,
         \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 ,
         \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 ,
         \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 ,
         \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 ,
         \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 ,
         \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 ,
         \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 ,
         \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 ,
         \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 ,
         \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
         \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 ,
         \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 ,
         \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 ,
         \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 ,
         \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 ,
         \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 ,
         \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 ,
         \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 ,
         \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 ,
         \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 ,
         \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 ,
         \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 ,
         \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 ,
         \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 ,
         \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 ,
         \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 ,
         \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 ,
         \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 ,
         \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
         \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 ,
         \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 ,
         \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 ,
         \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 ,
         \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 ,
         \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 ,
         \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 ,
         \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 ,
         \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 ,
         \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 ,
         \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 ,
         \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 ,
         \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 ,
         \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 ,
         \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 ,
         \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 ,
         \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 ,
         \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 ,
         \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 ,
         \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 ,
         \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 ,
         \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 ,
         \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 ,
         \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 ,
         \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 ,
         \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 ,
         \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 ,
         \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 ,
         \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 ,
         \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 ,
         \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 ,
         \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 ,
         \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 ,
         \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 ,
         \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 ,
         \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 ,
         \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 ,
         \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 ,
         \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 ,
         \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 ,
         \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 ,
         \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 ,
         \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 ,
         \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 ,
         \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 ,
         \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 ,
         \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 ,
         \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 ,
         \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 ,
         \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 ,
         \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 ,
         \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 ,
         \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 ,
         \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 ,
         \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 ,
         \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 ,
         \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 ,
         \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 ,
         \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 ,
         \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 ,
         \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 ,
         \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 ,
         \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 ,
         \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 ,
         \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 ,
         \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 ,
         \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 ,
         \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 ,
         \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 ,
         \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 ,
         \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 ,
         \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 ,
         \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 ,
         \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 ,
         \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 ,
         \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 ,
         \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 ,
         \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 ,
         \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 ,
         \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 ,
         \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 ,
         \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 ,
         \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 ,
         \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 ,
         \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 ,
         \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 ,
         \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 ,
         \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 ,
         \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 ,
         \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 ,
         \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 ,
         \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 ,
         \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 ,
         \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 ,
         \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 ,
         \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 ,
         \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 ,
         \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 ,
         \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 ,
         \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 ,
         \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 ,
         \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 ,
         \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 ,
         \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 ,
         \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 ,
         \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 ,
         \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 ,
         \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 ,
         \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 ,
         \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 ,
         \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 ,
         \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 ,
         \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 ,
         \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 ,
         \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 ,
         \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 ,
         \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 ,
         \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 ,
         \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 ,
         \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 ,
         \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 ,
         \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 ,
         \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 ,
         \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 ,
         \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 ,
         \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 ,
         \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 ,
         \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 ,
         \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 ,
         \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 ,
         \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 ,
         \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 ,
         \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 ,
         \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 ,
         \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 ,
         \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 ,
         \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 ,
         \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 ,
         \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 ,
         \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 ,
         \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 ,
         \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 ,
         \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 ,
         \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 ,
         \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 ,
         \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 ,
         \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 ,
         \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 ,
         \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 ,
         \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 ,
         \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 ,
         \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 ,
         \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 ,
         \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 ,
         \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 ,
         \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 ,
         \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 ,
         \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 ,
         \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 ,
         \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 ,
         \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 ,
         \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 ,
         \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 ,
         \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 ,
         \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 ,
         \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 ,
         \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 ,
         \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 ,
         \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 ,
         \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 ,
         \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 ,
         \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 ,
         \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 ,
         \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 ,
         \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 ,
         \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 ,
         \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 ,
         \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 ,
         \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 ,
         \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 ,
         \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 ,
         \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 ,
         \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 ,
         \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 ,
         \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 ,
         \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 ,
         \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 ,
         \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 ,
         \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 ,
         \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 ,
         \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 ,
         \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 ,
         \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 ,
         \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 ,
         \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 ,
         \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 ,
         \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 ,
         \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 ,
         \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 ,
         \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 ,
         \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 ,
         \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 ,
         \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 ,
         \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 ,
         \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 ,
         \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 ,
         \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 ,
         \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 ,
         \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 ,
         \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 ,
         \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 ,
         \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 ,
         \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 ,
         \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 ,
         \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 ,
         \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 ,
         \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 ,
         \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 ,
         \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 ,
         \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 ,
         \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 ,
         \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 ,
         \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 ,
         \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 ,
         \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 ,
         \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 ,
         \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 ,
         \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 ,
         \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 ,
         \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 ,
         \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 ,
         \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 ,
         \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 ,
         \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 ,
         \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 ,
         \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 ,
         \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 ,
         \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 ,
         \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 ,
         \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 ,
         \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 ,
         \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 ,
         \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 ,
         \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 ,
         \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 ,
         \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 ,
         \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 ,
         \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 ,
         \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 ,
         \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 ,
         \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 ,
         \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 ,
         \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 ,
         \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 ,
         \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 ,
         \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 ,
         \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 ,
         \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 ,
         \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 ,
         \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 ,
         \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 ,
         \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 ,
         \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 ,
         \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 ,
         \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 ,
         \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 ,
         \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 ,
         \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 ,
         \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 ,
         \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 ,
         \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 ,
         \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 ,
         \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 ,
         \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 ,
         \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 ,
         \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 ,
         \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 ,
         \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 ,
         \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 ,
         \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 ,
         \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 ,
         \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 ,
         \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 ,
         \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 ,
         \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 ,
         \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 ,
         \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 ,
         \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 ,
         \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 ,
         \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 ,
         \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 ,
         \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 ,
         \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 ,
         \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 ,
         \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 ,
         \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 ,
         \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 ,
         \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 ,
         \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 ,
         \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 ,
         \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 ,
         \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 ,
         \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 ,
         \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 ,
         \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 ,
         \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 ,
         \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 ,
         \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 ,
         \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 ,
         \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 ,
         \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 ,
         \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 ,
         \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 ,
         \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 ,
         \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 ,
         \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 ,
         \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 ,
         \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 ,
         \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 ,
         \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 ,
         \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 ,
         \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 ,
         \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 ,
         \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 ,
         \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 ,
         \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 ,
         \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 ,
         \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 ,
         \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 ,
         \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 ,
         \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 ,
         \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 ,
         \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 ,
         \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 ,
         \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 ,
         \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 ,
         \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 ,
         \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 ,
         \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 ,
         \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 ,
         \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 ,
         \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 ,
         \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 ,
         \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 ,
         \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 ,
         \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 ,
         \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 ,
         \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 ,
         \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 ,
         \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 ,
         \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 ,
         \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 ,
         \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 ,
         \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 ,
         \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 ,
         \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 ,
         \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 ,
         \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 ,
         \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 ,
         \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 ,
         \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 ,
         \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 ,
         \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 ,
         \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 ,
         \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 ,
         \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 ,
         \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 ,
         \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 ,
         \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 ,
         \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 ,
         \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 ,
         \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 ,
         \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 ,
         \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 ,
         \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 ,
         \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 ,
         \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 ,
         \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 ,
         \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 ,
         \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 ,
         \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 ,
         \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 ,
         \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 ,
         \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 ,
         \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 ,
         \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 ,
         \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 ,
         \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 ,
         \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 ,
         \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 ,
         \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 ,
         \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 ,
         \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 ,
         \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 ,
         \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 ,
         \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 ,
         \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 ,
         \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 ,
         \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 ,
         \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 ,
         \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 ,
         \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 ,
         \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 ,
         \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 ,
         \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 ,
         \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 ,
         \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 ,
         \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 ,
         \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 ,
         \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 ,
         \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 ,
         \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 ,
         \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 ,
         \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 ,
         \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 ,
         \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 ,
         \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 ,
         \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 ,
         \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 ,
         \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 ,
         \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 ,
         \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 ,
         \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 ,
         \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 ,
         \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 ,
         \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 ,
         \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 ,
         \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 ,
         \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 ,
         \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 ,
         \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 ,
         \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 ,
         \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 ,
         \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 ,
         \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 ,
         \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 ,
         \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 ,
         \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 ,
         \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 ,
         \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 ,
         \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 ,
         \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 ,
         \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 ,
         \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 ,
         \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 ,
         \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 ,
         \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 ,
         \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 ,
         \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 ,
         \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 ,
         \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 ,
         \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 ,
         \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 ,
         \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 ,
         \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 ,
         \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 ,
         \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 ,
         \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 ,
         \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 ,
         \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 ,
         \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 ,
         \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 ,
         \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 ,
         \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 ,
         \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 ,
         \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 ,
         \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 ,
         \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 ,
         \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 ,
         \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 ,
         \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 ,
         \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 ,
         \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 ,
         \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 ,
         \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 ,
         \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 ,
         \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 ,
         \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 ,
         \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 ,
         \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 ,
         \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 ,
         \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 ,
         \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 ,
         \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 ,
         \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 ,
         \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 ,
         \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 ,
         \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 ,
         \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 ,
         \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 ,
         \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 ,
         \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 ,
         \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 ,
         \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 ,
         \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 ,
         \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 ,
         \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 ,
         \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 ,
         \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 ,
         \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 ,
         \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 ,
         \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 ,
         \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 ,
         \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 ,
         \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 ,
         \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 ,
         \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 ,
         \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 ,
         \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 ,
         \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 ,
         \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 ,
         \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 ,
         \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 ,
         \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 ,
         \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 ,
         \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 ,
         \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 ,
         \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 ,
         \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 ,
         \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 ,
         \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 ,
         \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 ,
         \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 ,
         \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 ,
         \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 ,
         \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 ,
         \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 ,
         \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 ,
         \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 ,
         \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 ,
         \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 ,
         \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 ,
         \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 ,
         \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 ,
         \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 ,
         \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 ,
         \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 ,
         \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 ,
         \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 ,
         \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 ,
         \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 ,
         \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 ,
         \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 ,
         \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 ,
         \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 ,
         \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 ,
         \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 ,
         \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 ,
         \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 ,
         \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 ,
         \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 ,
         \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 ,
         \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 ,
         \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 ,
         \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 ,
         \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 ,
         \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 ,
         \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 ,
         \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 ,
         \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 ,
         \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 ,
         \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 ,
         \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 ,
         \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 ,
         \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 ,
         \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 ,
         \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 ,
         \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 ,
         \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 ,
         \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 ,
         \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 ,
         \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 ,
         \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 ,
         \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 ,
         \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 ,
         \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 ,
         \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 ,
         \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 ,
         \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 ,
         \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 ,
         \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 ,
         \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 ,
         \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 ,
         \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 ,
         \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 ,
         \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 ,
         \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 ,
         \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 ,
         \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 ,
         \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 ,
         \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 ,
         \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 ,
         \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 ,
         \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 ,
         \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 ,
         \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 ,
         \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 ,
         \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 ,
         \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 ,
         \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 ,
         \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 ,
         \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 ,
         \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 ,
         \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 ,
         \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 ,
         \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 ,
         \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 ,
         \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 ,
         \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 ,
         \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 ,
         \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 ,
         \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 ,
         \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 ,
         \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 ,
         \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 ,
         \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 ,
         \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 ,
         \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 ,
         \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 ,
         \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 ,
         \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 ,
         \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 ,
         \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 ,
         \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 ,
         \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 ,
         \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 ,
         \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 ,
         \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 ,
         \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 ,
         \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 ,
         \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 ,
         \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 ,
         \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 ,
         \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 ,
         \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 ,
         \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 ,
         \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 ,
         \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 ,
         \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 ,
         \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 ,
         \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 ,
         \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 ,
         \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 ,
         \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 ,
         \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 ,
         \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 ,
         \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 ,
         \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 ,
         \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 ,
         \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 ,
         \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 ,
         \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 ,
         \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 ,
         \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 ,
         \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 ,
         \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 ,
         \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 ,
         \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 ,
         \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 ,
         \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 ,
         \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 ,
         \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 ,
         \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 ,
         \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 ,
         \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 ,
         \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 ,
         \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 ,
         \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 ,
         \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 ,
         \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 ,
         \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 ,
         \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 ,
         \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 ,
         \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 ,
         \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 ,
         \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 ,
         \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 ,
         \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 ,
         \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 ,
         \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 ,
         \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 ,
         \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 ,
         \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 ,
         \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 ,
         \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 ,
         \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 ,
         \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 ,
         \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 ,
         \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 ,
         \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 ,
         \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 ,
         \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 ,
         \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 ,
         \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 ,
         \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 ,
         \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 ,
         \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 ,
         \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 ,
         \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 ,
         \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 ,
         \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 ,
         \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 ,
         \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 ,
         \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 ,
         \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 ,
         \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 ,
         \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 ,
         \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 ,
         \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 ,
         \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 ,
         \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 ,
         \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 ,
         \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 ,
         \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 ,
         \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 ,
         \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 ,
         \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 ,
         \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 ,
         \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 ,
         \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 ,
         \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 ,
         \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 ,
         \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 ,
         \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 ,
         \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 ,
         \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 ,
         \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 ,
         \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 ,
         \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 ,
         \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 ,
         \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 ,
         \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 ,
         \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 ,
         \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 ,
         \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 ,
         \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 ,
         \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 ,
         \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 ,
         \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 ,
         \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 ,
         \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 ,
         \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 ,
         \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 ,
         \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 ,
         \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 ,
         \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 ,
         \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 ,
         \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 ,
         \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 ,
         \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 ,
         \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 ,
         \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 ,
         \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 ,
         \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 ,
         \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 ,
         \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 ,
         \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 ,
         \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 ,
         \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 ,
         \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 ,
         \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 ,
         \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 ,
         \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 ,
         \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 ,
         \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 ,
         \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 ,
         \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 ,
         \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 ,
         \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 ,
         \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 ,
         \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 ,
         \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 ,
         \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 ,
         \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 ,
         \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 ,
         \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 ,
         \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 ,
         \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 ,
         \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 ,
         \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 ,
         \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 ,
         \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 ,
         \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 ,
         \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 ,
         \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 ,
         \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 ,
         \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 ,
         \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 ,
         \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 ,
         \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 ,
         \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 ,
         \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 ,
         \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 ,
         \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 ,
         \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 ,
         \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 ,
         \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 ,
         \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 ,
         \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 ,
         \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 ,
         \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 ,
         \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 ,
         \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 ,
         \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 ,
         \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 ,
         \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 ,
         \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 ,
         \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 ,
         \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 ,
         \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 ,
         \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 ,
         \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 ,
         \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 ,
         \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 ,
         \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 ,
         \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 ,
         \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 ,
         \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 ,
         \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 ,
         \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 ,
         \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 ,
         \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 ,
         \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 ,
         \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 ,
         \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 ,
         \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 ,
         \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 ,
         \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 ,
         \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 ,
         \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 ,
         \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 ,
         \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 ,
         \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 ,
         \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 ,
         \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 ,
         \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 ,
         \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 ,
         \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 ,
         \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 ,
         \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 ,
         \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 ,
         \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 ,
         \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 ,
         \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 ,
         \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 ,
         \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 ,
         \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 ,
         \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 ,
         \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 ,
         \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 ,
         \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 ,
         \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 ,
         \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 ,
         \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 ,
         \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 ,
         \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 ,
         \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 ,
         \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 ,
         \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 ,
         \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 ,
         \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 ,
         \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 ,
         \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 ,
         \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 ,
         \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 ,
         \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 ,
         \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 ,
         \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 ,
         \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 ,
         \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 ,
         \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 ,
         \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 ,
         \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 ,
         \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 ,
         \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 ,
         \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 ,
         \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 ,
         \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 ,
         \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 ,
         \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 ,
         \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 ,
         \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 ,
         \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 ,
         \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 ,
         \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 ,
         \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 ,
         \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 ,
         \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 ,
         \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 ,
         \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 ,
         \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 ,
         \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 ,
         \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 ,
         \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 ,
         \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 ,
         \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 ,
         \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 ,
         \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 ,
         \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 ,
         \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 ,
         \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 ,
         \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 ,
         \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 ,
         \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 ,
         \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 ,
         \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 ,
         \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 ,
         \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 ,
         \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 ,
         \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 ,
         \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 ,
         \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 ,
         \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 ,
         \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 ,
         \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 ,
         \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 ,
         \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 ,
         \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 ,
         \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 ,
         \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 ,
         \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 ,
         \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 ,
         \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 ,
         \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 ,
         \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 ,
         \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 ,
         \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 ,
         \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 ,
         \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 ,
         \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 ,
         \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 ,
         \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 ,
         \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 ,
         \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 ,
         \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 ,
         \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 ,
         \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 ,
         \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 ,
         \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 ,
         \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 ,
         \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 ,
         \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 ,
         \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 ,
         \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 ,
         \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 ,
         \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 ,
         \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 ,
         \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 ,
         \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 ,
         \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 ,
         \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 ,
         \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 ,
         \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 ,
         \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 ,
         \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 ,
         \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 ,
         \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 ,
         \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 ,
         \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 ,
         \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 ,
         \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 ,
         \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 ,
         \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 ,
         \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 ,
         \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 ,
         \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 ,
         \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 ,
         \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 ,
         \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 ,
         \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 ,
         \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 ,
         \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 ,
         \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 ,
         \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 ,
         \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 ,
         \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 ,
         \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 ,
         \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 ,
         \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 ,
         \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 ,
         \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 ,
         \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 ,
         \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 ,
         \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 ,
         \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 ,
         \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 ,
         \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 ,
         \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 ,
         \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 ,
         \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 ,
         \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 ,
         \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 ,
         \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 ,
         \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 ,
         \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 ,
         \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 ,
         \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 ,
         \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 ,
         \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 ,
         \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 ,
         \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 ,
         \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 ,
         \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 ,
         \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 ,
         \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 ,
         \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 ,
         \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 ,
         \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 ,
         \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 ,
         \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 ,
         \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 ,
         \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 ,
         \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 ,
         \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 ,
         \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 ,
         \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 ,
         \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 ,
         \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 ,
         \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 ,
         \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 ,
         \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 ,
         \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 ,
         \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 ,
         \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 ,
         \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 ,
         \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 ,
         \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 ,
         \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 ,
         \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 ,
         \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 ,
         \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 ,
         \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 ,
         \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 ,
         \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 ,
         \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 ,
         \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 ,
         \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 ,
         \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 ,
         \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 ,
         \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 ,
         \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 ,
         \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 ,
         \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 ,
         \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 ,
         \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 ,
         \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 ,
         \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 ,
         \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 ,
         \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 ,
         \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 ,
         \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 ,
         \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 ,
         \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 ,
         \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 ,
         \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 ,
         \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 ,
         \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 ,
         \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 ,
         \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 ,
         \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 ,
         \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 ,
         \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 ,
         \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 ,
         \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 ,
         \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 ,
         \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 ,
         \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 ,
         \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 ,
         \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 ,
         \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 ,
         \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 ,
         \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 ,
         \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 ,
         \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 ,
         \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 ,
         \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 ,
         \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 ,
         \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 ,
         \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 ,
         \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 ,
         \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 ,
         \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 ,
         \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 ,
         \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 ,
         \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 ,
         \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 ,
         \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 ,
         \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 ,
         \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 ,
         \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 ,
         \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 ,
         \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 ,
         \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 ,
         \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 ,
         \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 ,
         \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 ,
         \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 ,
         \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 ,
         \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 ,
         \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 ,
         \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 ,
         \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 ,
         \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 ,
         \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 ,
         \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 ,
         \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 ,
         \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 ,
         \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 ,
         \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 ,
         \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 ,
         \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 ,
         \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 ,
         \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 ,
         \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 ,
         \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 ,
         \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 ,
         \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 ,
         \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 ,
         \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 ,
         \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 ,
         \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 ,
         \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 ,
         \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 ,
         \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 ,
         \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 ,
         \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 ,
         \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 ,
         \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 ,
         \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 ,
         \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 ,
         \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 ,
         \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 ,
         \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 ,
         \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 ,
         \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 ,
         \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 ,
         \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 ,
         \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 ,
         \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 ,
         \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 ,
         \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 ,
         \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 ,
         \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 ,
         \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 ,
         \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 ,
         \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 ,
         \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 ,
         \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 ,
         \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 ,
         \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 ,
         \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 ,
         \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 ,
         \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 ,
         \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 ,
         \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 ,
         \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 ,
         \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 ,
         \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 ,
         \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 ,
         \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 ,
         \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 ,
         \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 ,
         \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 ,
         \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 ,
         \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 ,
         \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 ,
         \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 ,
         \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 ,
         \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 ,
         \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 ,
         \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 ,
         \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 ,
         \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 ,
         \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 ,
         \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 ,
         \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 ,
         \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 ,
         \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 ,
         \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 ,
         \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 ,
         \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 ,
         \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 ,
         \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 ,
         \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 ,
         \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 ,
         \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 ,
         \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 ,
         \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 ,
         \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 ,
         \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 ,
         \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 ,
         \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 ,
         \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 ,
         \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 ,
         \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 ,
         \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 ,
         \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 ,
         \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 ,
         \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 ,
         \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 ,
         \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 ,
         \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 ,
         \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 ,
         \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 ,
         \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 ,
         \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 ,
         \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 ,
         \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 ,
         \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 ,
         \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 ,
         \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 ,
         \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 ,
         \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 ,
         \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 ,
         \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 ,
         \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 ,
         \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 ,
         \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 ,
         \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 ,
         \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 ,
         \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 ,
         \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 ,
         \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 ,
         \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 ,
         \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 ,
         \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 ,
         \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 ,
         \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 ,
         \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 ,
         \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 ,
         \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 ,
         \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 ,
         \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 ,
         \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 ,
         \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 ,
         \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 ,
         \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 ,
         \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 ,
         \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 ,
         \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 ,
         \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 ,
         \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 ,
         \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 ,
         \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 ,
         \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 ,
         \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 ,
         \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 ,
         \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 ,
         \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 ,
         \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 ,
         \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 ,
         \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 ,
         \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 ,
         \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 ,
         \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 ,
         \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 ,
         \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 ,
         \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 ,
         \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 ,
         \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 ,
         \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 ,
         \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 ,
         \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 ,
         \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 ,
         \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 ,
         \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 ,
         \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 ,
         \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 ,
         \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 ,
         \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 ,
         \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 ,
         \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 ,
         \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 ,
         \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 ,
         \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 ,
         \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 ,
         \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 ,
         \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 ,
         \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 ,
         \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 ,
         \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 ,
         \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 ,
         \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 ,
         \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 ,
         \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 ,
         \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 ,
         \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 ,
         \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 ,
         \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 ,
         \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 ,
         \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 ,
         \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 ,
         \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 ,
         \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 ,
         \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 ,
         \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 ,
         \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 ,
         \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 ,
         \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 ,
         \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 ,
         \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 ,
         \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 ,
         \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 ,
         \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 ,
         \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 ,
         \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 ,
         \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 ,
         \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 ,
         \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 ,
         \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 ,
         \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 ,
         \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 ,
         \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 ,
         \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 ,
         \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 ,
         \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 ,
         \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 ,
         \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 ,
         \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 ,
         \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 ,
         \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 ,
         \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 ,
         \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 ,
         \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 ,
         \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 ,
         \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 ,
         \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 ,
         \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 ,
         \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 ,
         \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 ,
         \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 ,
         \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 ,
         \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 ,
         \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 ,
         \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 ,
         \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 ,
         \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 ,
         \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 ,
         \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 ,
         \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 ,
         \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 ,
         \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 ,
         \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 ,
         \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 ,
         \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 ,
         \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 ,
         \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 ,
         \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 ,
         \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 ,
         \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 ,
         \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 ,
         \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 ,
         \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 ,
         \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 ,
         \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 ,
         \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 ,
         \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 ,
         \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 ,
         \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 ,
         \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 ,
         \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 ,
         \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 ,
         \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 ,
         \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 ,
         \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 ,
         \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 ,
         \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 ,
         \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 ,
         \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 ,
         \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 ,
         \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 ,
         \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 ,
         \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 ,
         \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 ,
         \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 ,
         \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 ,
         \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 ,
         \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 ,
         \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 ,
         \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 ,
         \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 ,
         \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 ,
         \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 ,
         \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 ,
         \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 ,
         \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 ,
         \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 ,
         \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 ,
         \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 ,
         \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 ,
         \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 ,
         \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 ,
         \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 ,
         \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 ,
         \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 ,
         \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 ,
         \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 ,
         \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 ,
         \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 ,
         \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 ,
         \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 ,
         \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 ,
         \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 ,
         \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 ,
         \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 ,
         \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 ,
         \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 ,
         \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 ,
         \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 ,
         \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 ,
         \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 ,
         \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 ,
         \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 ,
         \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 ,
         \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 ,
         \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 ,
         \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 ,
         \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 ,
         \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 ,
         \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 ,
         \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 ,
         \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 ,
         \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 ,
         \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 ,
         \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 ,
         \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 ,
         \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 ,
         \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 ,
         \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 ,
         \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 ,
         \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 ,
         \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 ,
         \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 ,
         \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 ,
         \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 ,
         \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 ,
         \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 ,
         \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 ,
         \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 ,
         \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 ,
         \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 ,
         \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 ,
         \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 ,
         \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 ,
         \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 ,
         \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 ,
         \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 ,
         \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 ,
         \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 ,
         \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 ,
         \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 ,
         \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 ,
         \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 ,
         \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 ,
         \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 ,
         \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 ,
         \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 ,
         \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 ,
         \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 ,
         \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 ,
         \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 ,
         \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 ,
         \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 ,
         \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 ,
         \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 ,
         \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 ,
         \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 ,
         \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 ,
         \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 ,
         \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 ,
         \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 ,
         \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 ,
         \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 ,
         \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 ,
         \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 ,
         \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 ,
         \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 ,
         \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 ,
         \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 ,
         \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 ,
         \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 ,
         \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 ,
         \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 ,
         \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 ,
         \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 ,
         \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 ,
         \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 ,
         \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 ,
         \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 ,
         \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 ,
         \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 ,
         \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 ,
         \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 ,
         \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 ,
         \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 ,
         \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 ,
         \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 ,
         \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 ,
         \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 ,
         \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 ,
         \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 ,
         \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 ,
         \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 ,
         \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 ,
         \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 ,
         \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 ,
         \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 ,
         \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 ,
         \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 ,
         \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 ,
         \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 ,
         \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 ,
         \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 ,
         \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 ,
         \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 ,
         \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 ,
         \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 ,
         \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 ,
         \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 ,
         \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 ,
         \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 ,
         \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 ,
         \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 ,
         \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 ,
         \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 ,
         \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 ,
         \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 ,
         \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 ,
         \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 ,
         \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 ,
         \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 ,
         \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 ,
         \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 ,
         \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 ,
         \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 ,
         \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 ,
         \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 ,
         \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 ,
         \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 ,
         \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 ,
         \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 ,
         \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 ,
         \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 ,
         \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 ,
         \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 ,
         \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 ,
         \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 ,
         \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 ,
         \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 ,
         \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 ,
         \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 ,
         \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 ,
         \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 ,
         \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 ,
         \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 ,
         \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 ,
         \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 ,
         \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 ,
         \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 ,
         \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 ,
         \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 ,
         \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 ,
         \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 ,
         \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 ,
         \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 ,
         \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 ,
         \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 ,
         \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 ,
         \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 ,
         \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 ,
         \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 ,
         \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 ,
         \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 ,
         \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 ,
         \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 ,
         \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 ,
         \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 ,
         \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 ,
         \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 ,
         \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 ,
         \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 ,
         \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 ,
         \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 ,
         \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 ,
         \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 ,
         \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 ,
         \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 ,
         \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 ,
         \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 ,
         \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 ,
         \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 ,
         \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 ,
         \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 ,
         \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 ,
         \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 ,
         \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 ,
         \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 ,
         \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 ,
         \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 ,
         \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 ,
         \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 ,
         \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 ,
         \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 ,
         \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 ,
         \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 ,
         \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 ,
         \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 ,
         \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 ,
         \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 ,
         \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 ,
         \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 ,
         \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 ,
         \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 ,
         \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 ,
         \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 ,
         \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 ,
         \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 ,
         \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 ,
         \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 ,
         \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 ,
         \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 ,
         \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 ,
         \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 ,
         \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 ,
         \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 ,
         \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 ,
         \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 ,
         \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 ,
         \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 ,
         \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 ,
         \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 ,
         \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 ,
         \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 ,
         \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 ,
         \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 ,
         \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 ,
         \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 ,
         \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 ,
         \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 ,
         \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 ,
         \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 ,
         \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 ,
         \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 ,
         \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 ,
         \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 ,
         \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 ,
         \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 ,
         \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 ,
         \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 ,
         \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 ,
         \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 ,
         \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 ,
         \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 ,
         \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 ,
         \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 ,
         \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 ,
         \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 ,
         \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 ,
         \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 ,
         \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 ,
         \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 ,
         \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 ,
         \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 ,
         \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 ,
         \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 ,
         \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 ,
         \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 ,
         \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 ,
         \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 ,
         \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 ,
         \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 ,
         \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 ,
         \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 ,
         \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 ,
         \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 ,
         \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 ,
         \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 ,
         \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 ,
         \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 ,
         \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 ,
         \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 ,
         \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 ,
         \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 ,
         \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 ,
         \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 ,
         \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 ,
         \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 ,
         \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 ,
         \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 ,
         \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 ,
         \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 ,
         \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 ,
         \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 ,
         \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 ,
         \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 ,
         \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 ,
         \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 ,
         \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 ,
         \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 ,
         \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 ,
         \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 ,
         \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 ,
         \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 ,
         \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 ,
         \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 ,
         \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 ,
         \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 ,
         \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 ,
         \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 ,
         \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 ,
         \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 ,
         \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 ,
         \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 ,
         \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 ,
         \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 ,
         \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 ,
         \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 ,
         \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 ,
         \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 ,
         \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 ,
         \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 ,
         \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 ,
         \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 ,
         \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 ,
         \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 ,
         \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 ,
         \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 ,
         \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 ,
         \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 ,
         \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 ,
         \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 ,
         \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 ,
         \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 ,
         \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 ,
         \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 ,
         \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 ,
         \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 ,
         \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 ,
         \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 ,
         \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 ,
         \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 ,
         \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 ,
         \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 ,
         \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 ,
         \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 ,
         \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 ,
         \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 ,
         \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 ,
         \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 ,
         \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 ,
         \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 ,
         \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 ,
         \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 ,
         \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 ,
         \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 ,
         \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 ,
         \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 ,
         \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 ,
         \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 ,
         \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 ,
         \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 ,
         \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 ,
         \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 ,
         \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 ,
         \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 ,
         \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 ,
         \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 ,
         \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 ,
         \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 ,
         \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 ,
         \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 ,
         \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 ,
         \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 ,
         \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 ,
         \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 ,
         \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 ,
         \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 ,
         \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 ,
         \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 ,
         \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 ,
         \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 ,
         \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 ,
         \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 ,
         \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 ,
         \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 ,
         \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 ,
         \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 ,
         \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 ,
         \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 ,
         \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 ,
         \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 ,
         \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 ,
         \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 ,
         \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 ,
         \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 ,
         \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 ,
         \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 ,
         \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 ,
         \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 ,
         \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 ,
         \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 ,
         \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 ,
         \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 ,
         \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 ,
         \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 ,
         \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 ,
         \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 ,
         \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 ,
         \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 ,
         \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 ,
         \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 ,
         \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 ,
         \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 ,
         \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 ,
         \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 ,
         \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 ,
         \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 ,
         \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 ,
         \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 ,
         \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 ,
         \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 ,
         \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 ,
         \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 ,
         \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 ,
         \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 ,
         \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 ,
         \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 ,
         \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 ,
         \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 ,
         \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 ,
         \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 ,
         \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 ,
         \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 ,
         \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 ,
         \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 ,
         \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 ,
         \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 ,
         \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 ,
         \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 ,
         \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 ,
         \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 ,
         \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 ,
         \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 ,
         \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 ,
         \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 ,
         \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 ,
         \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 ,
         \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 ,
         \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 ,
         \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 ,
         \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 ,
         \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 ,
         \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 ,
         \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 ,
         \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 ,
         \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 ,
         \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 ,
         \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 ,
         \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 ,
         \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 ,
         \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 ,
         \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 ,
         \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 ,
         \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 ,
         \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 ,
         \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 ,
         \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 ,
         \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 ,
         \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 ,
         \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 ,
         \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 ,
         \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 ,
         \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 ,
         \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 ,
         \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 ,
         \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 ,
         \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 ,
         \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 ,
         \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 ,
         \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 ,
         \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 ,
         \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 ,
         \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 ,
         \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 ,
         \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 ,
         \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 ,
         \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 ,
         \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 ,
         \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 ,
         \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 ,
         \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 ,
         \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 ,
         \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 ,
         \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 ,
         \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 ,
         \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 ,
         \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 ,
         \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 ,
         \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 ,
         \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 ,
         \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 ,
         \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 ,
         \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 ,
         \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 ,
         \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 ,
         \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 ,
         \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 ,
         \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 ,
         \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 ,
         \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 ,
         \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 ,
         \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 ,
         \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 ,
         \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 ,
         \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 ,
         \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 ,
         \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 ,
         \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 ,
         \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 ,
         \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 ,
         \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 ,
         \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 ,
         \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 ,
         \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 ,
         \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 ,
         \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 ,
         \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 ,
         \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 ,
         \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 ,
         \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 ,
         \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 ,
         \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 ,
         \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 ,
         \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 ,
         \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 ,
         \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 ,
         \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 ,
         \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 ,
         \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 ,
         \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 ,
         \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 ,
         \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 ,
         \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 ,
         \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 ,
         \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 ,
         \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 ,
         \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 ,
         \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 ,
         \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 ,
         \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 ,
         \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 ,
         \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 ,
         \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 ,
         \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 ,
         \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 ,
         \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 ,
         \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 ,
         \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 ,
         \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 ,
         \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 ,
         \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 ,
         \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 ,
         \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 ,
         \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 ,
         \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 ,
         \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 ,
         \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 ,
         \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 ,
         \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 ,
         \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 ,
         \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 ,
         \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 ,
         \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 ,
         \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 ,
         \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 ,
         \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 ,
         \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 ,
         \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 ,
         \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 ,
         \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 ,
         \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 ,
         \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 ,
         \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 ,
         \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 ,
         \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 ,
         \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 ,
         \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 ,
         \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 ,
         \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 ,
         \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 ,
         \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 ,
         \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 ,
         \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 ,
         \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 ,
         \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 ,
         \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 ,
         \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 ,
         \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 ,
         \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 ,
         \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 ,
         \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 ,
         \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 ,
         \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 ,
         \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 ,
         \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 ,
         \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 ,
         \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 ,
         \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 ,
         \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 ,
         \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 ,
         \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 ,
         \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 ,
         \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 ,
         \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 ,
         \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 ,
         \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 ,
         \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 ,
         \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 ,
         \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 ,
         \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 ,
         \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 ,
         \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 ,
         \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 ,
         \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 ,
         \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 ,
         \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 ,
         \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 ,
         \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 ,
         \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 ,
         \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 ,
         \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 ,
         \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 ,
         \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 ,
         \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 ,
         \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 ,
         \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 ,
         \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 ,
         \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 ,
         \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 ,
         \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 ,
         \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 ,
         \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 ,
         \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 ,
         \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 ,
         \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 ,
         \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 ,
         \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 ,
         \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 ,
         \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 ,
         \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 ,
         \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 ,
         \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 ,
         \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 ,
         \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 ,
         \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 ,
         \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 ,
         \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 ,
         \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 ,
         \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 ,
         \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 ,
         \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 ,
         \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 ,
         \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 ,
         \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 ,
         \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 ,
         \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 ,
         \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 ,
         \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 ,
         \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 ,
         \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 ,
         \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 ,
         \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 ,
         \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 ,
         \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 ,
         \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 ,
         \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 ,
         \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 ,
         \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 ,
         \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 ,
         \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 ,
         \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 ,
         \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 ,
         \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 ,
         \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 ,
         \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 ,
         \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 ,
         \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 ,
         \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 ,
         \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 ,
         \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 ,
         \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 ,
         \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 ,
         \22253 , \22254 , \22255 , \22256 , \22257_nG5617 , \22258 , \22259 , \22260 , \22261_nG561a , \22262 ,
         \22263 , \22264_nG561d , \22265 , \22266 , \22267_nG5620 , \22268 , \22269 , \22270_nG5623 , \22271 , \22272 ,
         \22273_nG5626 , \22274 , \22275 , \22276_nG5629 , \22277 , \22278 , \22279_nG562c , \22280 , \22281 , \22282_nG562f ,
         \22283 , \22284 , \22285_nG5632 , \22286 , \22287 , \22288_nG5635 , \22289 , \22290 , \22291_nG5638 , \22292 ,
         \22293 , \22294_nG563b , \22295 , \22296 , \22297_nG563e , \22298 , \22299 , \22300_nG5641 , \22301 , \22302 ,
         \22303_nG5644 , \22304 , \22305 , \22306_nG5647 , \22307 , \22308 , \22309_nG564a , \22310 , \22311 , \22312_nG564d ,
         \22313 , \22314 , \22315_nG5650 , \22316 , \22317 , \22318_nG5653 , \22319 , \22320 , \22321_nG5656 , \22322 ,
         \22323 , \22324_nG5659 , \22325 , \22326 , \22327_nG565c , \22328 , \22329 , \22330_nG565f , \22331 , \22332 ,
         \22333_nG5662 , \22334 , \22335 , \22336_nG5665 , \22337 , \22338 , \22339_nG5668 , \22340 , \22341 , \22342_nG566b ,
         \22343 , \22344 , \22345_nG566e , \22346 , \22347 , \22348_nG5671 , \22349 , \22350 , \22351_nG5674 , \22352 ,
         \22353 , \22354_nG5677 , \22355 , \22356 , \22357_nG567a , \22358 , \22359 , \22360_nG567d , \22361 , \22362 ,
         \22363_nG5680 , \22364 , \22365 , \22366_nG5683 , \22367 , \22368 , \22369_nG5686 , \22370 , \22371 , \22372_nG5689 ,
         \22373 , \22374 , \22375_nG568c , \22376 , \22377 , \22378_nG568f , \22379 , \22380 , \22381_nG5692 , \22382 ,
         \22383 , \22384_nG5695 , \22385 , \22386 , \22387_nG5698 , \22388 , \22389 , \22390_nG569b , \22391 , \22392 ,
         \22393_nG569e , \22394 , \22395 , \22396_nG56a1 , \22397 , \22398 , \22399_nG56a4 , \22400 , \22401 , \22402_nG56a7 ,
         \22403 , \22404 , \22405_nG56aa , \22406 , \22407 , \22408_nG56ad , \22409 , \22410 , \22411_nG56b0 , \22412 ,
         \22413 , \22414_nG56b3 , \22415 , \22416 , \22417_nG56b6 , \22418 , \22419 , \22420_nG56b9 , \22421 , \22422 ,
         \22423_nG56bc , \22424 , \22425 , \22426_nG56bf , \22427 , \22428 , \22429_nG56c2 , \22430 , \22431 , \22432_nG56c5 ,
         \22433 , \22434 , \22435_nG56c8 , \22436 , \22437 , \22438_nG56cb , \22439 , \22440 , \22441_nG56ce , \22442 ,
         \22443 , \22444_nG56d1 , \22445 , \22446 , \22447_nG56d4 , \22448 , \22449 , \22450_nG56d7 , \22451 , \22452 ,
         \22453_nG56da , \22454 , \22455 , \22456_nG56dd , \22457 , \22458 , \22459_nG56e0 , \22460 , \22461 , \22462_nG56e3 ,
         \22463 , \22464 , \22465_nG56e6 , \22466 , \22467 , \22468_nG56e9 , \22469 , \22470 , \22471_nG56ec , \22472 ,
         \22473 , \22474_nG56ef , \22475 , \22476 , \22477_nG56f2 , \22478 , \22479 , \22480_nG56f5 , \22481 , \22482 ,
         \22483_nG56f8 , \22484 , \22485 , \22486_nG56fb , \22487 , \22488 , \22489_nG56fe , \22490 , \22491 , \22492_nG5701 ,
         \22493 , \22494 , \22495_nG5704 , \22496 , \22497 , \22498_nG5707 , \22499 , \22500 , \22501_nG570a , \22502 ,
         \22503 , \22504_nG570d , \22505 , \22506 , \22507_nG5710 , \22508 , \22509 , \22510_nG5713 , \22511 , \22512 ,
         \22513_nG5716 , \22514 , \22515 , \22516_nG5719 , \22517 , \22518 , \22519_nG571c , \22520 , \22521 , \22522_nG571f ,
         \22523 , \22524 , \22525_nG5722 , \22526 , \22527 , \22528_nG5725 , \22529 , \22530 , \22531_nG5728 , \22532 ,
         \22533 , \22534_nG572b , \22535 , \22536 , \22537_nG572e , \22538 , \22539 , \22540_nG5731 , \22541 , \22542 ,
         \22543_nG5734 , \22544 , \22545 , \22546_nG5737 , \22547 , \22548 , \22549_nG573a , \22550 , \22551 , \22552_nG573d ,
         \22553 , \22554 , \22555_nG5740 , \22556 , \22557 , \22558_nG5743 , \22559 , \22560 , \22561_nG5746 , \22562 ,
         \22563 , \22564_nG5749 , \22565 , \22566 , \22567_nG574c , \22568 , \22569 , \22570_nG574f , \22571 , \22572 ,
         \22573_nG5752 , \22574 , \22575 , \22576_nG5755 , \22577 , \22578 , \22579_nG5758 , \22580 , \22581 , \22582_nG575b ,
         \22583 , \22584 , \22585_nG575e , \22586 , \22587 , \22588_nG5761 , \22589 , \22590 , \22591_nG5764 , \22592 ,
         \22593 , \22594_nG5767 , \22595 , \22596 , \22597_nG576a , \22598 , \22599 , \22600_nG576d , \22601 , \22602 ,
         \22603_nG5770 , \22604 , \22605 , \22606_nG5773 , \22607 , \22608 , \22609_nG5776 , \22610 , \22611 , \22612_nG5779 ,
         \22613 , \22614 , \22615_nG577c , \22616 , \22617 , \22618_nG577f , \22619 , \22620 , \22621_nG5782 , \22622 ,
         \22623 , \22624_nG5785 , \22625 , \22626 , \22627_nG5788 , \22628 , \22629 , \22630_nG578b , \22631 , \22632 ,
         \22633_nG578e , \22634 , \22635 , \22636_nG5791 , \22637 , \22638 , \22639_nG5794 , \22640 , \22641_nG2fd , \22642_nG5796 ,
         \22643_nG5797 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 ,
         \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 ,
         \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 ,
         \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 ,
         \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 ,
         \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 ,
         \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 ,
         \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 ,
         \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 ,
         \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 ,
         \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 ,
         \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 ,
         \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 ,
         \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 ,
         \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 ,
         \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 ,
         \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 ,
         \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 ,
         \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 ,
         \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 ,
         \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 ,
         \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 ,
         \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 ,
         \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 ,
         \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 ,
         \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899_nG5898 , \22900 , \22901 , \22902 ,
         \22903_nG589b , \22904 , \22905 , \22906 , \22907_nG589e , \22908 , \22909 , \22910 , \22911_nG58a1 , \22912 ,
         \22913 , \22914 , \22915_nG58a4 , \22916 , \22917 , \22918 , \22919_nG58a7 , \22920 , \22921 , \22922 ,
         \22923_nG58aa , \22924 , \22925 , \22926 , \22927_nG58ad , \22928 , \22929 , \22930 , \22931_nG58b0 , \22932 ,
         \22933 , \22934 , \22935_nG58b3 , \22936 , \22937 , \22938 , \22939_nG58b6 , \22940 , \22941 , \22942 ,
         \22943_nG58b9 , \22944 , \22945 , \22946 , \22947_nG58bc , \22948 , \22949 , \22950 , \22951_nG58bf , \22952 ,
         \22953 , \22954 , \22955_nG58c2 , \22956 , \22957 , \22958 , \22959_nG58c5 , \22960 , \22961 , \22962 ,
         \22963_nG58c8 , \22964 , \22965 , \22966 , \22967_nG58cb , \22968 , \22969 , \22970 , \22971_nG58ce , \22972 ,
         \22973 , \22974 , \22975_nG58d1 , \22976 , \22977 , \22978 , \22979_nG58d4 , \22980 , \22981 , \22982 ,
         \22983_nG58d7 , \22984 , \22985 , \22986 , \22987_nG58da , \22988 , \22989 , \22990 , \22991_nG58dd , \22992 ,
         \22993 , \22994 , \22995_nG58e0 , \22996 , \22997 , \22998 , \22999_nG58e3 , \23000 , \23001 , \23002 ,
         \23003_nG58e6 , \23004 , \23005 , \23006 , \23007_nG58e9 , \23008 , \23009 , \23010 , \23011_nG58ec , \23012 ,
         \23013 , \23014 , \23015_nG58ef , \23016 , \23017 , \23018 , \23019_nG58f2 , \23020 , \23021 , \23022 ,
         \23023_nG58f5 , \23024 , \23025 , \23026 , \23027_nG58f8 , \23028 , \23029 , \23030 , \23031_nG58fb , \23032 ,
         \23033 , \23034 , \23035_nG58fe , \23036 , \23037 , \23038 , \23039_nG5901 , \23040 , \23041 , \23042 ,
         \23043_nG5904 , \23044 , \23045 , \23046 , \23047_nG5907 , \23048 , \23049 , \23050 , \23051_nG590a , \23052 ,
         \23053 , \23054 , \23055_nG590d , \23056 , \23057 , \23058 , \23059_nG5910 , \23060 , \23061 , \23062 ,
         \23063_nG5913 , \23064 , \23065 , \23066 , \23067_nG5916 , \23068 , \23069 , \23070 , \23071_nG5919 , \23072 ,
         \23073 , \23074 , \23075_nG591c , \23076 , \23077 , \23078 , \23079_nG591f , \23080 , \23081 , \23082 ,
         \23083_nG5922 , \23084 , \23085 , \23086 , \23087_nG5925 , \23088 , \23089 , \23090 , \23091_nG5928 , \23092 ,
         \23093 , \23094 , \23095_nG592b , \23096 , \23097 , \23098 , \23099_nG592e , \23100 , \23101 , \23102 ,
         \23103_nG5931 , \23104 , \23105 , \23106 , \23107_nG5934 , \23108 , \23109 , \23110 , \23111_nG5937 , \23112 ,
         \23113 , \23114 , \23115_nG593a , \23116 , \23117 , \23118 , \23119_nG593d , \23120 , \23121 , \23122 ,
         \23123_nG5940 , \23124 , \23125 , \23126 , \23127_nG5943 , \23128 , \23129 , \23130 , \23131_nG5946 , \23132 ,
         \23133 , \23134 , \23135_nG5949 , \23136 , \23137 , \23138 , \23139_nG594c , \23140 , \23141 , \23142 ,
         \23143_nG594f , \23144 , \23145 , \23146 , \23147_nG5952 , \23148 , \23149 , \23150 , \23151_nG5955 , \23152 ,
         \23153 , \23154 , \23155_nG5958 , \23156 , \23157 , \23158 , \23159_nG595b , \23160 , \23161 , \23162 ,
         \23163_nG595e , \23164 , \23165 , \23166 , \23167_nG5961 , \23168 , \23169 , \23170 , \23171_nG5964 , \23172 ,
         \23173 , \23174 , \23175_nG5967 , \23176 , \23177 , \23178 , \23179_nG596a , \23180 , \23181 , \23182 ,
         \23183_nG596d , \23184 , \23185 , \23186 , \23187_nG5970 , \23188 , \23189 , \23190 , \23191_nG5973 , \23192 ,
         \23193 , \23194 , \23195_nG5976 , \23196 , \23197 , \23198 , \23199_nG5979 , \23200 , \23201 , \23202 ,
         \23203_nG597c , \23204 , \23205 , \23206 , \23207_nG597f , \23208 , \23209 , \23210 , \23211_nG5982 , \23212 ,
         \23213 , \23214 , \23215_nG5985 , \23216 , \23217 , \23218 , \23219_nG5988 , \23220 , \23221 , \23222 ,
         \23223_nG598b , \23224 , \23225 , \23226 , \23227_nG598e , \23228 , \23229 , \23230 , \23231_nG5991 , \23232 ,
         \23233 , \23234 , \23235_nG5994 , \23236 , \23237 , \23238 , \23239_nG5997 , \23240 , \23241 , \23242 ,
         \23243_nG599a , \23244 , \23245 , \23246 , \23247_nG599d , \23248 , \23249 , \23250 , \23251_nG59a0 , \23252 ,
         \23253 , \23254 , \23255_nG59a3 , \23256 , \23257 , \23258 , \23259_nG59a6 , \23260 , \23261 , \23262 ,
         \23263_nG59a9 , \23264 , \23265 , \23266 , \23267_nG59ac , \23268 , \23269 , \23270 , \23271_nG59af , \23272 ,
         \23273 , \23274 , \23275_nG59b2 , \23276 , \23277 , \23278 , \23279_nG59b5 , \23280 , \23281 , \23282 ,
         \23283_nG59b8 , \23284 , \23285 , \23286 , \23287_nG59bb , \23288 , \23289 , \23290 , \23291_nG59be , \23292 ,
         \23293 , \23294 , \23295_nG59c1 , \23296 , \23297 , \23298 , \23299_nG59c4 , \23300 , \23301 , \23302 ,
         \23303_nG59c7 , \23304 , \23305 , \23306 , \23307_nG59ca , \23308 , \23309 , \23310 , \23311_nG59cd , \23312 ,
         \23313 , \23314 , \23315_nG59d0 , \23316 , \23317 , \23318 , \23319_nG59d3 , \23320 , \23321 , \23322 ,
         \23323_nG59d6 , \23324 , \23325 , \23326 , \23327_nG59d9 , \23328 , \23329 , \23330 , \23331_nG59dc , \23332 ,
         \23333 , \23334 , \23335_nG59df , \23336 , \23337 , \23338 , \23339_nG59e2 , \23340 , \23341 , \23342 ,
         \23343_nG59e5 , \23344 , \23345 , \23346 , \23347_nG59e8 , \23348 , \23349 , \23350 , \23351_nG59eb , \23352 ,
         \23353 , \23354 , \23355_nG59ee , \23356 ;
buf \U$labaj2367 ( R_81_84446b8, \22900 );
buf \U$labaj2368 ( R_82_8444760, \22904 );
buf \U$labaj2369 ( R_83_8444808, \22908 );
buf \U$labaj2370 ( R_84_84448b0, \22912 );
buf \U$labaj2371 ( R_85_8444958, \22916 );
buf \U$labaj2372 ( R_86_8444a00, \22920 );
buf \U$labaj2373 ( R_87_9bec6f8, \22924 );
buf \U$labaj2374 ( R_88_9bec7a0, \22928 );
buf \U$labaj2375 ( R_89_9bec848, \22932 );
buf \U$labaj2376 ( R_8a_9bec8f0, \22936 );
buf \U$labaj2377 ( R_8b_9bec998, \22940 );
buf \U$labaj2378 ( R_8c_9beca40, \22944 );
buf \U$labaj2379 ( R_8d_9becae8, \22948 );
buf \U$labaj2380 ( R_8e_9becb90, \22952 );
buf \U$labaj2381 ( R_8f_9becc38, \22956 );
buf \U$labaj2382 ( R_90_9becce0, \22960 );
buf \U$labaj2383 ( R_91_9becd88, \22964 );
buf \U$labaj2384 ( R_92_9bece30, \22968 );
buf \U$labaj2385 ( R_93_9beced8, \22972 );
buf \U$labaj2386 ( R_94_9becf80, \22976 );
buf \U$labaj2387 ( R_95_9bed028, \22980 );
buf \U$labaj2388 ( R_96_9bed0d0, \22984 );
buf \U$labaj2389 ( R_97_9bed178, \22988 );
buf \U$labaj2390 ( R_98_9bed220, \22992 );
buf \U$labaj2391 ( R_99_9bed2c8, \22996 );
buf \U$labaj2392 ( R_9a_9bed370, \23000 );
buf \U$labaj2393 ( R_9b_9bed418, \23004 );
buf \U$labaj2394 ( R_9c_9bed4c0, \23008 );
buf \U$labaj2395 ( R_9d_9bed568, \23012 );
buf \U$labaj2396 ( R_9e_9bed610, \23016 );
buf \U$labaj2397 ( R_9f_9bed6b8, \23020 );
buf \U$labaj2398 ( R_a0_9bed760, \23024 );
buf \U$labaj2399 ( R_a1_9bed808, \23028 );
buf \U$labaj2400 ( R_a2_9bed8b0, \23032 );
buf \U$labaj2401 ( R_a3_9bed958, \23036 );
buf \U$labaj2402 ( R_a4_9beda00, \23040 );
buf \U$labaj2403 ( R_a5_9bedaa8, \23044 );
buf \U$labaj2404 ( R_a6_9bedb50, \23048 );
buf \U$labaj2405 ( R_a7_9bedbf8, \23052 );
buf \U$labaj2406 ( R_a8_9bedca0, \23056 );
buf \U$labaj2407 ( R_a9_9bedd48, \23060 );
buf \U$labaj2408 ( R_aa_9beddf0, \23064 );
buf \U$labaj2409 ( R_ab_9bede98, \23068 );
buf \U$labaj2410 ( R_ac_9bedf40, \23072 );
buf \U$labaj2411 ( R_ad_9bedfe8, \23076 );
buf \U$labaj2412 ( R_ae_9bee090, \23080 );
buf \U$labaj2413 ( R_af_9bee138, \23084 );
buf \U$labaj2414 ( R_b0_9bee1e0, \23088 );
buf \U$labaj2415 ( R_b1_9bee288, \23092 );
buf \U$labaj2416 ( R_b2_9bee330, \23096 );
buf \U$labaj2417 ( R_b3_9bee3d8, \23100 );
buf \U$labaj2418 ( R_b4_9bee480, \23104 );
buf \U$labaj2419 ( R_b5_9bee528, \23108 );
buf \U$labaj2420 ( R_b6_9bee5d0, \23112 );
buf \U$labaj2421 ( R_b7_9bee678, \23116 );
buf \U$labaj2422 ( R_b8_9bee720, \23120 );
buf \U$labaj2423 ( R_b9_9bee7c8, \23124 );
buf \U$labaj2424 ( R_ba_9bee870, \23128 );
buf \U$labaj2425 ( R_bb_9bee918, \23132 );
buf \U$labaj2426 ( R_bc_9bee9c0, \23136 );
buf \U$labaj2427 ( R_bd_9beea68, \23140 );
buf \U$labaj2428 ( R_be_9beeb10, \23144 );
buf \U$labaj2429 ( R_bf_9beebb8, \23148 );
buf \U$labaj2430 ( R_c0_9beec60, \23152 );
buf \U$labaj2431 ( R_c1_9beed08, \23156 );
buf \U$labaj2432 ( R_c2_9beedb0, \23160 );
buf \U$labaj2433 ( R_c3_9beee58, \23164 );
buf \U$labaj2434 ( R_c4_9beef00, \23168 );
buf \U$labaj2435 ( R_c5_9beefa8, \23172 );
buf \U$labaj2436 ( R_c6_9bef050, \23176 );
buf \U$labaj2437 ( R_c7_9bef0f8, \23180 );
buf \U$labaj2438 ( R_c8_9bef1a0, \23184 );
buf \U$labaj2439 ( R_c9_9bef248, \23188 );
buf \U$labaj2440 ( R_ca_9bef2f0, \23192 );
buf \U$labaj2441 ( R_cb_9bef398, \23196 );
buf \U$labaj2442 ( R_cc_9bef440, \23200 );
buf \U$labaj2443 ( R_cd_9bef4e8, \23204 );
buf \U$labaj2444 ( R_ce_9bef590, \23208 );
buf \U$labaj2445 ( R_cf_9bef638, \23212 );
buf \U$labaj2446 ( R_d0_9bef6e0, \23216 );
buf \U$labaj2447 ( R_d1_9bef788, \23220 );
buf \U$labaj2448 ( R_d2_9bef830, \23224 );
buf \U$labaj2449 ( R_d3_9bef8d8, \23228 );
buf \U$labaj2450 ( R_d4_9bef980, \23232 );
buf \U$labaj2451 ( R_d5_9befa28, \23236 );
buf \U$labaj2452 ( R_d6_9befad0, \23240 );
buf \U$labaj2453 ( R_d7_9befb78, \23244 );
buf \U$labaj2454 ( R_d8_9befc20, \23248 );
buf \U$labaj2455 ( R_d9_9befcc8, \23252 );
buf \U$labaj2456 ( R_da_9befd70, \23256 );
buf \U$labaj2457 ( R_db_9befe18, \23260 );
buf \U$labaj2458 ( R_dc_9befec0, \23264 );
buf \U$labaj2459 ( R_dd_9beff68, \23268 );
buf \U$labaj2460 ( R_de_9bf0010, \23272 );
buf \U$labaj2461 ( R_df_9bf00b8, \23276 );
buf \U$labaj2462 ( R_e0_9bf0160, \23280 );
buf \U$labaj2463 ( R_e1_9bf0208, \23284 );
buf \U$labaj2464 ( R_e2_9bf02b0, \23288 );
buf \U$labaj2465 ( R_e3_9bf0358, \23292 );
buf \U$labaj2466 ( R_e4_9bf0400, \23296 );
buf \U$labaj2467 ( R_e5_9bf04a8, \23300 );
buf \U$labaj2468 ( R_e6_9bf0550, \23304 );
buf \U$labaj2469 ( R_e7_9bf05f8, \23308 );
buf \U$labaj2470 ( R_e8_9bf06a0, \23312 );
buf \U$labaj2471 ( R_e9_9bf0748, \23316 );
buf \U$labaj2472 ( R_ea_9bf07f0, \23320 );
buf \U$labaj2473 ( R_eb_9bf0898, \23324 );
buf \U$labaj2474 ( R_ec_9bf0940, \23328 );
buf \U$labaj2475 ( R_ed_9bf09e8, \23332 );
buf \U$labaj2476 ( R_ee_9bf0a90, \23336 );
buf \U$labaj2477 ( R_ef_9bf0b38, \23340 );
buf \U$labaj2478 ( R_f0_9bf0be0, \23344 );
buf \U$labaj2479 ( R_f1_9bf0c88, \23348 );
buf \U$labaj2480 ( R_f2_9bf0d30, \23352 );
buf \U$labaj2481 ( R_f3_9bf0dd8, \23356 );
buf \U$1 ( \984 , RIc0d9478_65);
buf \U$2 ( \985 , RIc0d7678_1);
buf \U$3 ( \986 , RIc0d76f0_2);
xor \U$4 ( \987 , \985 , \986 );
buf \U$5 ( \988 , RIc0d7768_3);
xor \U$6 ( \989 , \986 , \988 );
not \U$7 ( \990 , \989 );
and \U$8 ( \991 , \987 , \990 );
and \U$9 ( \992 , \984 , \991 );
not \U$10 ( \993 , \992 );
and \U$11 ( \994 , \986 , \988 );
not \U$12 ( \995 , \994 );
and \U$13 ( \996 , \985 , \995 );
xnor \U$14 ( \997 , \993 , \996 );
buf \U$15 ( \998 , RIc0d94f0_66);
and \U$16 ( \999 , \998 , \985 );
or \U$17 ( \1000 , \997 , \999 );
not \U$18 ( \1001 , \996 );
xor \U$19 ( \1002 , \1000 , \1001 );
and \U$20 ( \1003 , \984 , \985 );
xor \U$21 ( \1004 , \1002 , \1003 );
buf \U$22 ( \1005 , RIc0d77e0_4);
buf \U$23 ( \1006 , RIc0d7858_5);
and \U$24 ( \1007 , \1005 , \1006 );
not \U$25 ( \1008 , \1007 );
and \U$26 ( \1009 , \988 , \1008 );
not \U$27 ( \1010 , \1009 );
and \U$28 ( \1011 , \998 , \991 );
and \U$29 ( \1012 , \984 , \989 );
nor \U$30 ( \1013 , \1011 , \1012 );
xnor \U$31 ( \1014 , \1013 , \996 );
and \U$32 ( \1015 , \1010 , \1014 );
buf \U$33 ( \1016 , RIc0d9568_67);
and \U$34 ( \1017 , \1016 , \985 );
and \U$35 ( \1018 , \1014 , \1017 );
and \U$36 ( \1019 , \1010 , \1017 );
or \U$37 ( \1020 , \1015 , \1018 , \1019 );
xnor \U$38 ( \1021 , \997 , \999 );
and \U$39 ( \1022 , \1020 , \1021 );
xor \U$40 ( \1023 , \1004 , \1022 );
xor \U$41 ( \1024 , \1020 , \1021 );
xor \U$42 ( \1025 , \988 , \1005 );
xor \U$43 ( \1026 , \1005 , \1006 );
not \U$44 ( \1027 , \1026 );
and \U$45 ( \1028 , \1025 , \1027 );
and \U$46 ( \1029 , \984 , \1028 );
not \U$47 ( \1030 , \1029 );
xnor \U$48 ( \1031 , \1030 , \1009 );
and \U$49 ( \1032 , \1016 , \991 );
and \U$50 ( \1033 , \998 , \989 );
nor \U$51 ( \1034 , \1032 , \1033 );
xnor \U$52 ( \1035 , \1034 , \996 );
and \U$53 ( \1036 , \1031 , \1035 );
buf \U$54 ( \1037 , RIc0d95e0_68);
and \U$55 ( \1038 , \1037 , \985 );
and \U$56 ( \1039 , \1035 , \1038 );
and \U$57 ( \1040 , \1031 , \1038 );
or \U$58 ( \1041 , \1036 , \1039 , \1040 );
buf \U$59 ( \1042 , RIc0d78d0_6);
buf \U$60 ( \1043 , RIc0d7948_7);
and \U$61 ( \1044 , \1042 , \1043 );
not \U$62 ( \1045 , \1044 );
and \U$63 ( \1046 , \1006 , \1045 );
not \U$64 ( \1047 , \1046 );
and \U$65 ( \1048 , \998 , \1028 );
and \U$66 ( \1049 , \984 , \1026 );
nor \U$67 ( \1050 , \1048 , \1049 );
xnor \U$68 ( \1051 , \1050 , \1009 );
and \U$69 ( \1052 , \1047 , \1051 );
and \U$70 ( \1053 , \1037 , \991 );
and \U$71 ( \1054 , \1016 , \989 );
nor \U$72 ( \1055 , \1053 , \1054 );
xnor \U$73 ( \1056 , \1055 , \996 );
and \U$74 ( \1057 , \1051 , \1056 );
and \U$75 ( \1058 , \1047 , \1056 );
or \U$76 ( \1059 , \1052 , \1057 , \1058 );
xor \U$77 ( \1060 , \1031 , \1035 );
xor \U$78 ( \1061 , \1060 , \1038 );
or \U$79 ( \1062 , \1059 , \1061 );
and \U$80 ( \1063 , \1041 , \1062 );
xor \U$81 ( \1064 , \1010 , \1014 );
xor \U$82 ( \1065 , \1064 , \1017 );
and \U$83 ( \1066 , \1062 , \1065 );
and \U$84 ( \1067 , \1041 , \1065 );
or \U$85 ( \1068 , \1063 , \1066 , \1067 );
and \U$86 ( \1069 , \1024 , \1068 );
xor \U$87 ( \1070 , \1024 , \1068 );
xor \U$88 ( \1071 , \1041 , \1062 );
xor \U$89 ( \1072 , \1071 , \1065 );
xor \U$90 ( \1073 , \1006 , \1042 );
xor \U$91 ( \1074 , \1042 , \1043 );
not \U$92 ( \1075 , \1074 );
and \U$93 ( \1076 , \1073 , \1075 );
and \U$94 ( \1077 , \984 , \1076 );
not \U$95 ( \1078 , \1077 );
xnor \U$96 ( \1079 , \1078 , \1046 );
and \U$97 ( \1080 , \1016 , \1028 );
and \U$98 ( \1081 , \998 , \1026 );
nor \U$99 ( \1082 , \1080 , \1081 );
xnor \U$100 ( \1083 , \1082 , \1009 );
and \U$101 ( \1084 , \1079 , \1083 );
buf \U$102 ( \1085 , RIc0d9658_69);
and \U$103 ( \1086 , \1085 , \991 );
and \U$104 ( \1087 , \1037 , \989 );
nor \U$105 ( \1088 , \1086 , \1087 );
xnor \U$106 ( \1089 , \1088 , \996 );
and \U$107 ( \1090 , \1083 , \1089 );
and \U$108 ( \1091 , \1079 , \1089 );
or \U$109 ( \1092 , \1084 , \1090 , \1091 );
buf \U$110 ( \1093 , RIc0d96d0_70);
and \U$111 ( \1094 , \1093 , \985 );
buf \U$112 ( \1095 , \1094 );
and \U$113 ( \1096 , \1092 , \1095 );
and \U$114 ( \1097 , \1085 , \985 );
and \U$115 ( \1098 , \1095 , \1097 );
and \U$116 ( \1099 , \1092 , \1097 );
or \U$117 ( \1100 , \1096 , \1098 , \1099 );
buf \U$118 ( \1101 , RIc0d79c0_8);
buf \U$119 ( \1102 , RIc0d7a38_9);
and \U$120 ( \1103 , \1101 , \1102 );
not \U$121 ( \1104 , \1103 );
and \U$122 ( \1105 , \1043 , \1104 );
not \U$123 ( \1106 , \1105 );
and \U$124 ( \1107 , \998 , \1076 );
and \U$125 ( \1108 , \984 , \1074 );
nor \U$126 ( \1109 , \1107 , \1108 );
xnor \U$127 ( \1110 , \1109 , \1046 );
and \U$128 ( \1111 , \1106 , \1110 );
and \U$129 ( \1112 , \1037 , \1028 );
and \U$130 ( \1113 , \1016 , \1026 );
nor \U$131 ( \1114 , \1112 , \1113 );
xnor \U$132 ( \1115 , \1114 , \1009 );
and \U$133 ( \1116 , \1110 , \1115 );
and \U$134 ( \1117 , \1106 , \1115 );
or \U$135 ( \1118 , \1111 , \1116 , \1117 );
xor \U$136 ( \1119 , \1079 , \1083 );
xor \U$137 ( \1120 , \1119 , \1089 );
and \U$138 ( \1121 , \1118 , \1120 );
not \U$139 ( \1122 , \1094 );
and \U$140 ( \1123 , \1120 , \1122 );
and \U$141 ( \1124 , \1118 , \1122 );
or \U$142 ( \1125 , \1121 , \1123 , \1124 );
xor \U$143 ( \1126 , \1047 , \1051 );
xor \U$144 ( \1127 , \1126 , \1056 );
and \U$145 ( \1128 , \1125 , \1127 );
xor \U$146 ( \1129 , \1092 , \1095 );
xor \U$147 ( \1130 , \1129 , \1097 );
and \U$148 ( \1131 , \1127 , \1130 );
and \U$149 ( \1132 , \1125 , \1130 );
or \U$150 ( \1133 , \1128 , \1131 , \1132 );
and \U$151 ( \1134 , \1100 , \1133 );
xnor \U$152 ( \1135 , \1059 , \1061 );
and \U$153 ( \1136 , \1133 , \1135 );
and \U$154 ( \1137 , \1100 , \1135 );
or \U$155 ( \1138 , \1134 , \1136 , \1137 );
and \U$156 ( \1139 , \1072 , \1138 );
xor \U$157 ( \1140 , \1072 , \1138 );
xor \U$158 ( \1141 , \1100 , \1133 );
xor \U$159 ( \1142 , \1141 , \1135 );
xor \U$160 ( \1143 , \1043 , \1101 );
xor \U$161 ( \1144 , \1101 , \1102 );
not \U$162 ( \1145 , \1144 );
and \U$163 ( \1146 , \1143 , \1145 );
and \U$164 ( \1147 , \984 , \1146 );
not \U$165 ( \1148 , \1147 );
xnor \U$166 ( \1149 , \1148 , \1105 );
and \U$167 ( \1150 , \1016 , \1076 );
and \U$168 ( \1151 , \998 , \1074 );
nor \U$169 ( \1152 , \1150 , \1151 );
xnor \U$170 ( \1153 , \1152 , \1046 );
and \U$171 ( \1154 , \1149 , \1153 );
and \U$172 ( \1155 , \1085 , \1028 );
and \U$173 ( \1156 , \1037 , \1026 );
nor \U$174 ( \1157 , \1155 , \1156 );
xnor \U$175 ( \1158 , \1157 , \1009 );
and \U$176 ( \1159 , \1153 , \1158 );
and \U$177 ( \1160 , \1149 , \1158 );
or \U$178 ( \1161 , \1154 , \1159 , \1160 );
buf \U$179 ( \1162 , RIc0d9748_71);
and \U$180 ( \1163 , \1162 , \991 );
and \U$181 ( \1164 , \1093 , \989 );
nor \U$182 ( \1165 , \1163 , \1164 );
xnor \U$183 ( \1166 , \1165 , \996 );
buf \U$184 ( \1167 , RIc0d97c0_72);
and \U$185 ( \1168 , \1167 , \985 );
or \U$186 ( \1169 , \1166 , \1168 );
and \U$187 ( \1170 , \1161 , \1169 );
and \U$188 ( \1171 , \1093 , \991 );
and \U$189 ( \1172 , \1085 , \989 );
nor \U$190 ( \1173 , \1171 , \1172 );
xnor \U$191 ( \1174 , \1173 , \996 );
and \U$192 ( \1175 , \1169 , \1174 );
and \U$193 ( \1176 , \1161 , \1174 );
or \U$194 ( \1177 , \1170 , \1175 , \1176 );
and \U$195 ( \1178 , \1162 , \985 );
xor \U$196 ( \1179 , \1106 , \1110 );
xor \U$197 ( \1180 , \1179 , \1115 );
and \U$198 ( \1181 , \1178 , \1180 );
and \U$199 ( \1182 , \1177 , \1181 );
xor \U$200 ( \1183 , \1118 , \1120 );
xor \U$201 ( \1184 , \1183 , \1122 );
and \U$202 ( \1185 , \1181 , \1184 );
and \U$203 ( \1186 , \1177 , \1184 );
or \U$204 ( \1187 , \1182 , \1185 , \1186 );
xor \U$205 ( \1188 , \1125 , \1127 );
xor \U$206 ( \1189 , \1188 , \1130 );
and \U$207 ( \1190 , \1187 , \1189 );
and \U$208 ( \1191 , \1142 , \1190 );
xor \U$209 ( \1192 , \1142 , \1190 );
xor \U$210 ( \1193 , \1187 , \1189 );
buf \U$211 ( \1194 , RIc0d7ab0_10);
buf \U$212 ( \1195 , RIc0d7b28_11);
and \U$213 ( \1196 , \1194 , \1195 );
not \U$214 ( \1197 , \1196 );
and \U$215 ( \1198 , \1102 , \1197 );
not \U$216 ( \1199 , \1198 );
and \U$217 ( \1200 , \998 , \1146 );
and \U$218 ( \1201 , \984 , \1144 );
nor \U$219 ( \1202 , \1200 , \1201 );
xnor \U$220 ( \1203 , \1202 , \1105 );
and \U$221 ( \1204 , \1199 , \1203 );
and \U$222 ( \1205 , \1037 , \1076 );
and \U$223 ( \1206 , \1016 , \1074 );
nor \U$224 ( \1207 , \1205 , \1206 );
xnor \U$225 ( \1208 , \1207 , \1046 );
and \U$226 ( \1209 , \1203 , \1208 );
and \U$227 ( \1210 , \1199 , \1208 );
or \U$228 ( \1211 , \1204 , \1209 , \1210 );
and \U$229 ( \1212 , \1093 , \1028 );
and \U$230 ( \1213 , \1085 , \1026 );
nor \U$231 ( \1214 , \1212 , \1213 );
xnor \U$232 ( \1215 , \1214 , \1009 );
and \U$233 ( \1216 , \1167 , \991 );
and \U$234 ( \1217 , \1162 , \989 );
nor \U$235 ( \1218 , \1216 , \1217 );
xnor \U$236 ( \1219 , \1218 , \996 );
and \U$237 ( \1220 , \1215 , \1219 );
buf \U$238 ( \1221 , RIc0d9838_73);
and \U$239 ( \1222 , \1221 , \985 );
and \U$240 ( \1223 , \1219 , \1222 );
and \U$241 ( \1224 , \1215 , \1222 );
or \U$242 ( \1225 , \1220 , \1223 , \1224 );
and \U$243 ( \1226 , \1211 , \1225 );
xnor \U$244 ( \1227 , \1166 , \1168 );
and \U$245 ( \1228 , \1225 , \1227 );
and \U$246 ( \1229 , \1211 , \1227 );
or \U$247 ( \1230 , \1226 , \1228 , \1229 );
xor \U$248 ( \1231 , \1161 , \1169 );
xor \U$249 ( \1232 , \1231 , \1174 );
and \U$250 ( \1233 , \1230 , \1232 );
xor \U$251 ( \1234 , \1178 , \1180 );
and \U$252 ( \1235 , \1232 , \1234 );
and \U$253 ( \1236 , \1230 , \1234 );
or \U$254 ( \1237 , \1233 , \1235 , \1236 );
xor \U$255 ( \1238 , \1177 , \1181 );
xor \U$256 ( \1239 , \1238 , \1184 );
and \U$257 ( \1240 , \1237 , \1239 );
and \U$258 ( \1241 , \1193 , \1240 );
xor \U$259 ( \1242 , \1193 , \1240 );
xor \U$260 ( \1243 , \1237 , \1239 );
xor \U$261 ( \1244 , \1102 , \1194 );
xor \U$262 ( \1245 , \1194 , \1195 );
not \U$263 ( \1246 , \1245 );
and \U$264 ( \1247 , \1244 , \1246 );
and \U$265 ( \1248 , \984 , \1247 );
not \U$266 ( \1249 , \1248 );
xnor \U$267 ( \1250 , \1249 , \1198 );
and \U$268 ( \1251 , \1016 , \1146 );
and \U$269 ( \1252 , \998 , \1144 );
nor \U$270 ( \1253 , \1251 , \1252 );
xnor \U$271 ( \1254 , \1253 , \1105 );
and \U$272 ( \1255 , \1250 , \1254 );
and \U$273 ( \1256 , \1085 , \1076 );
and \U$274 ( \1257 , \1037 , \1074 );
nor \U$275 ( \1258 , \1256 , \1257 );
xnor \U$276 ( \1259 , \1258 , \1046 );
and \U$277 ( \1260 , \1254 , \1259 );
and \U$278 ( \1261 , \1250 , \1259 );
or \U$279 ( \1262 , \1255 , \1260 , \1261 );
and \U$280 ( \1263 , \1162 , \1028 );
and \U$281 ( \1264 , \1093 , \1026 );
nor \U$282 ( \1265 , \1263 , \1264 );
xnor \U$283 ( \1266 , \1265 , \1009 );
and \U$284 ( \1267 , \1221 , \991 );
and \U$285 ( \1268 , \1167 , \989 );
nor \U$286 ( \1269 , \1267 , \1268 );
xnor \U$287 ( \1270 , \1269 , \996 );
and \U$288 ( \1271 , \1266 , \1270 );
buf \U$289 ( \1272 , RIc0d98b0_74);
and \U$290 ( \1273 , \1272 , \985 );
and \U$291 ( \1274 , \1270 , \1273 );
and \U$292 ( \1275 , \1266 , \1273 );
or \U$293 ( \1276 , \1271 , \1274 , \1275 );
and \U$294 ( \1277 , \1262 , \1276 );
xor \U$295 ( \1278 , \1215 , \1219 );
xor \U$296 ( \1279 , \1278 , \1222 );
and \U$297 ( \1280 , \1276 , \1279 );
and \U$298 ( \1281 , \1262 , \1279 );
or \U$299 ( \1282 , \1277 , \1280 , \1281 );
xor \U$300 ( \1283 , \1149 , \1153 );
xor \U$301 ( \1284 , \1283 , \1158 );
and \U$302 ( \1285 , \1282 , \1284 );
xor \U$303 ( \1286 , \1211 , \1225 );
xor \U$304 ( \1287 , \1286 , \1227 );
and \U$305 ( \1288 , \1284 , \1287 );
and \U$306 ( \1289 , \1282 , \1287 );
or \U$307 ( \1290 , \1285 , \1288 , \1289 );
xor \U$308 ( \1291 , \1230 , \1232 );
xor \U$309 ( \1292 , \1291 , \1234 );
and \U$310 ( \1293 , \1290 , \1292 );
and \U$311 ( \1294 , \1243 , \1293 );
xor \U$312 ( \1295 , \1243 , \1293 );
xor \U$313 ( \1296 , \1290 , \1292 );
and \U$314 ( \1297 , \1093 , \1076 );
and \U$315 ( \1298 , \1085 , \1074 );
nor \U$316 ( \1299 , \1297 , \1298 );
xnor \U$317 ( \1300 , \1299 , \1046 );
and \U$318 ( \1301 , \1167 , \1028 );
and \U$319 ( \1302 , \1162 , \1026 );
nor \U$320 ( \1303 , \1301 , \1302 );
xnor \U$321 ( \1304 , \1303 , \1009 );
and \U$322 ( \1305 , \1300 , \1304 );
and \U$323 ( \1306 , \1272 , \991 );
and \U$324 ( \1307 , \1221 , \989 );
nor \U$325 ( \1308 , \1306 , \1307 );
xnor \U$326 ( \1309 , \1308 , \996 );
and \U$327 ( \1310 , \1304 , \1309 );
and \U$328 ( \1311 , \1300 , \1309 );
or \U$329 ( \1312 , \1305 , \1310 , \1311 );
buf \U$330 ( \1313 , RIc0d7ba0_12);
buf \U$331 ( \1314 , RIc0d7c18_13);
and \U$332 ( \1315 , \1313 , \1314 );
not \U$333 ( \1316 , \1315 );
and \U$334 ( \1317 , \1195 , \1316 );
not \U$335 ( \1318 , \1317 );
and \U$336 ( \1319 , \998 , \1247 );
and \U$337 ( \1320 , \984 , \1245 );
nor \U$338 ( \1321 , \1319 , \1320 );
xnor \U$339 ( \1322 , \1321 , \1198 );
and \U$340 ( \1323 , \1318 , \1322 );
and \U$341 ( \1324 , \1037 , \1146 );
and \U$342 ( \1325 , \1016 , \1144 );
nor \U$343 ( \1326 , \1324 , \1325 );
xnor \U$344 ( \1327 , \1326 , \1105 );
and \U$345 ( \1328 , \1322 , \1327 );
and \U$346 ( \1329 , \1318 , \1327 );
or \U$347 ( \1330 , \1323 , \1328 , \1329 );
or \U$348 ( \1331 , \1312 , \1330 );
xor \U$349 ( \1332 , \1199 , \1203 );
xor \U$350 ( \1333 , \1332 , \1208 );
and \U$351 ( \1334 , \1331 , \1333 );
xor \U$352 ( \1335 , \1262 , \1276 );
xor \U$353 ( \1336 , \1335 , \1279 );
and \U$354 ( \1337 , \1333 , \1336 );
and \U$355 ( \1338 , \1331 , \1336 );
or \U$356 ( \1339 , \1334 , \1337 , \1338 );
and \U$357 ( \1340 , \1162 , \1076 );
and \U$358 ( \1341 , \1093 , \1074 );
nor \U$359 ( \1342 , \1340 , \1341 );
xnor \U$360 ( \1343 , \1342 , \1046 );
and \U$361 ( \1344 , \1221 , \1028 );
and \U$362 ( \1345 , \1167 , \1026 );
nor \U$363 ( \1346 , \1344 , \1345 );
xnor \U$364 ( \1347 , \1346 , \1009 );
and \U$365 ( \1348 , \1343 , \1347 );
buf \U$366 ( \1349 , RIc0d9928_75);
and \U$367 ( \1350 , \1349 , \991 );
and \U$368 ( \1351 , \1272 , \989 );
nor \U$369 ( \1352 , \1350 , \1351 );
xnor \U$370 ( \1353 , \1352 , \996 );
and \U$371 ( \1354 , \1347 , \1353 );
and \U$372 ( \1355 , \1343 , \1353 );
or \U$373 ( \1356 , \1348 , \1354 , \1355 );
xor \U$374 ( \1357 , \1195 , \1313 );
xor \U$375 ( \1358 , \1313 , \1314 );
not \U$376 ( \1359 , \1358 );
and \U$377 ( \1360 , \1357 , \1359 );
and \U$378 ( \1361 , \984 , \1360 );
not \U$379 ( \1362 , \1361 );
xnor \U$380 ( \1363 , \1362 , \1317 );
and \U$381 ( \1364 , \1016 , \1247 );
and \U$382 ( \1365 , \998 , \1245 );
nor \U$383 ( \1366 , \1364 , \1365 );
xnor \U$384 ( \1367 , \1366 , \1198 );
and \U$385 ( \1368 , \1363 , \1367 );
and \U$386 ( \1369 , \1085 , \1146 );
and \U$387 ( \1370 , \1037 , \1144 );
nor \U$388 ( \1371 , \1369 , \1370 );
xnor \U$389 ( \1372 , \1371 , \1105 );
and \U$390 ( \1373 , \1367 , \1372 );
and \U$391 ( \1374 , \1363 , \1372 );
or \U$392 ( \1375 , \1368 , \1373 , \1374 );
and \U$393 ( \1376 , \1356 , \1375 );
buf \U$394 ( \1377 , RIc0d99a0_76);
and \U$395 ( \1378 , \1377 , \985 );
buf \U$396 ( \1379 , \1378 );
and \U$397 ( \1380 , \1375 , \1379 );
and \U$398 ( \1381 , \1356 , \1379 );
or \U$399 ( \1382 , \1376 , \1380 , \1381 );
and \U$400 ( \1383 , \1349 , \985 );
xor \U$401 ( \1384 , \1300 , \1304 );
xor \U$402 ( \1385 , \1384 , \1309 );
and \U$403 ( \1386 , \1383 , \1385 );
xor \U$404 ( \1387 , \1318 , \1322 );
xor \U$405 ( \1388 , \1387 , \1327 );
and \U$406 ( \1389 , \1385 , \1388 );
and \U$407 ( \1390 , \1383 , \1388 );
or \U$408 ( \1391 , \1386 , \1389 , \1390 );
and \U$409 ( \1392 , \1382 , \1391 );
xor \U$410 ( \1393 , \1266 , \1270 );
xor \U$411 ( \1394 , \1393 , \1273 );
and \U$412 ( \1395 , \1391 , \1394 );
and \U$413 ( \1396 , \1382 , \1394 );
or \U$414 ( \1397 , \1392 , \1395 , \1396 );
xor \U$415 ( \1398 , \1250 , \1254 );
xor \U$416 ( \1399 , \1398 , \1259 );
xnor \U$417 ( \1400 , \1312 , \1330 );
and \U$418 ( \1401 , \1399 , \1400 );
and \U$419 ( \1402 , \1397 , \1401 );
xor \U$420 ( \1403 , \1331 , \1333 );
xor \U$421 ( \1404 , \1403 , \1336 );
and \U$422 ( \1405 , \1401 , \1404 );
and \U$423 ( \1406 , \1397 , \1404 );
or \U$424 ( \1407 , \1402 , \1405 , \1406 );
and \U$425 ( \1408 , \1339 , \1407 );
xor \U$426 ( \1409 , \1282 , \1284 );
xor \U$427 ( \1410 , \1409 , \1287 );
and \U$428 ( \1411 , \1407 , \1410 );
and \U$429 ( \1412 , \1339 , \1410 );
or \U$430 ( \1413 , \1408 , \1411 , \1412 );
and \U$431 ( \1414 , \1296 , \1413 );
xor \U$432 ( \1415 , \1296 , \1413 );
xor \U$433 ( \1416 , \1339 , \1407 );
xor \U$434 ( \1417 , \1416 , \1410 );
buf \U$435 ( \1418 , RIc0d7c90_14);
buf \U$436 ( \1419 , RIc0d7d08_15);
and \U$437 ( \1420 , \1418 , \1419 );
not \U$438 ( \1421 , \1420 );
and \U$439 ( \1422 , \1314 , \1421 );
not \U$440 ( \1423 , \1422 );
and \U$441 ( \1424 , \998 , \1360 );
and \U$442 ( \1425 , \984 , \1358 );
nor \U$443 ( \1426 , \1424 , \1425 );
xnor \U$444 ( \1427 , \1426 , \1317 );
and \U$445 ( \1428 , \1423 , \1427 );
and \U$446 ( \1429 , \1037 , \1247 );
and \U$447 ( \1430 , \1016 , \1245 );
nor \U$448 ( \1431 , \1429 , \1430 );
xnor \U$449 ( \1432 , \1431 , \1198 );
and \U$450 ( \1433 , \1427 , \1432 );
and \U$451 ( \1434 , \1423 , \1432 );
or \U$452 ( \1435 , \1428 , \1433 , \1434 );
and \U$453 ( \1436 , \1093 , \1146 );
and \U$454 ( \1437 , \1085 , \1144 );
nor \U$455 ( \1438 , \1436 , \1437 );
xnor \U$456 ( \1439 , \1438 , \1105 );
and \U$457 ( \1440 , \1167 , \1076 );
and \U$458 ( \1441 , \1162 , \1074 );
nor \U$459 ( \1442 , \1440 , \1441 );
xnor \U$460 ( \1443 , \1442 , \1046 );
and \U$461 ( \1444 , \1439 , \1443 );
and \U$462 ( \1445 , \1272 , \1028 );
and \U$463 ( \1446 , \1221 , \1026 );
nor \U$464 ( \1447 , \1445 , \1446 );
xnor \U$465 ( \1448 , \1447 , \1009 );
and \U$466 ( \1449 , \1443 , \1448 );
and \U$467 ( \1450 , \1439 , \1448 );
or \U$468 ( \1451 , \1444 , \1449 , \1450 );
and \U$469 ( \1452 , \1435 , \1451 );
and \U$470 ( \1453 , \1377 , \991 );
and \U$471 ( \1454 , \1349 , \989 );
nor \U$472 ( \1455 , \1453 , \1454 );
xnor \U$473 ( \1456 , \1455 , \996 );
buf \U$474 ( \1457 , RIc0d9a18_77);
and \U$475 ( \1458 , \1457 , \985 );
and \U$476 ( \1459 , \1456 , \1458 );
and \U$477 ( \1460 , \1451 , \1459 );
and \U$478 ( \1461 , \1435 , \1459 );
or \U$479 ( \1462 , \1452 , \1460 , \1461 );
xor \U$480 ( \1463 , \1343 , \1347 );
xor \U$481 ( \1464 , \1463 , \1353 );
xor \U$482 ( \1465 , \1363 , \1367 );
xor \U$483 ( \1466 , \1465 , \1372 );
and \U$484 ( \1467 , \1464 , \1466 );
not \U$485 ( \1468 , \1378 );
and \U$486 ( \1469 , \1466 , \1468 );
and \U$487 ( \1470 , \1464 , \1468 );
or \U$488 ( \1471 , \1467 , \1469 , \1470 );
and \U$489 ( \1472 , \1462 , \1471 );
xor \U$490 ( \1473 , \1383 , \1385 );
xor \U$491 ( \1474 , \1473 , \1388 );
and \U$492 ( \1475 , \1471 , \1474 );
and \U$493 ( \1476 , \1462 , \1474 );
or \U$494 ( \1477 , \1472 , \1475 , \1476 );
xor \U$495 ( \1478 , \1382 , \1391 );
xor \U$496 ( \1479 , \1478 , \1394 );
and \U$497 ( \1480 , \1477 , \1479 );
xor \U$498 ( \1481 , \1399 , \1400 );
and \U$499 ( \1482 , \1479 , \1481 );
and \U$500 ( \1483 , \1477 , \1481 );
or \U$501 ( \1484 , \1480 , \1482 , \1483 );
xor \U$502 ( \1485 , \1397 , \1401 );
xor \U$503 ( \1486 , \1485 , \1404 );
and \U$504 ( \1487 , \1484 , \1486 );
and \U$505 ( \1488 , \1417 , \1487 );
xor \U$506 ( \1489 , \1417 , \1487 );
xor \U$507 ( \1490 , \1484 , \1486 );
xor \U$508 ( \1491 , \1314 , \1418 );
xor \U$509 ( \1492 , \1418 , \1419 );
not \U$510 ( \1493 , \1492 );
and \U$511 ( \1494 , \1491 , \1493 );
and \U$512 ( \1495 , \984 , \1494 );
not \U$513 ( \1496 , \1495 );
xnor \U$514 ( \1497 , \1496 , \1422 );
and \U$515 ( \1498 , \1016 , \1360 );
and \U$516 ( \1499 , \998 , \1358 );
nor \U$517 ( \1500 , \1498 , \1499 );
xnor \U$518 ( \1501 , \1500 , \1317 );
and \U$519 ( \1502 , \1497 , \1501 );
and \U$520 ( \1503 , \1085 , \1247 );
and \U$521 ( \1504 , \1037 , \1245 );
nor \U$522 ( \1505 , \1503 , \1504 );
xnor \U$523 ( \1506 , \1505 , \1198 );
and \U$524 ( \1507 , \1501 , \1506 );
and \U$525 ( \1508 , \1497 , \1506 );
or \U$526 ( \1509 , \1502 , \1507 , \1508 );
and \U$527 ( \1510 , \1162 , \1146 );
and \U$528 ( \1511 , \1093 , \1144 );
nor \U$529 ( \1512 , \1510 , \1511 );
xnor \U$530 ( \1513 , \1512 , \1105 );
and \U$531 ( \1514 , \1221 , \1076 );
and \U$532 ( \1515 , \1167 , \1074 );
nor \U$533 ( \1516 , \1514 , \1515 );
xnor \U$534 ( \1517 , \1516 , \1046 );
and \U$535 ( \1518 , \1513 , \1517 );
and \U$536 ( \1519 , \1349 , \1028 );
and \U$537 ( \1520 , \1272 , \1026 );
nor \U$538 ( \1521 , \1519 , \1520 );
xnor \U$539 ( \1522 , \1521 , \1009 );
and \U$540 ( \1523 , \1517 , \1522 );
and \U$541 ( \1524 , \1513 , \1522 );
or \U$542 ( \1525 , \1518 , \1523 , \1524 );
and \U$543 ( \1526 , \1509 , \1525 );
and \U$544 ( \1527 , \1457 , \991 );
and \U$545 ( \1528 , \1377 , \989 );
nor \U$546 ( \1529 , \1527 , \1528 );
xnor \U$547 ( \1530 , \1529 , \996 );
buf \U$548 ( \1531 , RIc0d9a90_78);
and \U$549 ( \1532 , \1531 , \985 );
or \U$550 ( \1533 , \1530 , \1532 );
and \U$551 ( \1534 , \1525 , \1533 );
and \U$552 ( \1535 , \1509 , \1533 );
or \U$553 ( \1536 , \1526 , \1534 , \1535 );
xor \U$554 ( \1537 , \1423 , \1427 );
xor \U$555 ( \1538 , \1537 , \1432 );
xor \U$556 ( \1539 , \1439 , \1443 );
xor \U$557 ( \1540 , \1539 , \1448 );
and \U$558 ( \1541 , \1538 , \1540 );
xor \U$559 ( \1542 , \1456 , \1458 );
and \U$560 ( \1543 , \1540 , \1542 );
and \U$561 ( \1544 , \1538 , \1542 );
or \U$562 ( \1545 , \1541 , \1543 , \1544 );
and \U$563 ( \1546 , \1536 , \1545 );
xor \U$564 ( \1547 , \1464 , \1466 );
xor \U$565 ( \1548 , \1547 , \1468 );
and \U$566 ( \1549 , \1545 , \1548 );
and \U$567 ( \1550 , \1536 , \1548 );
or \U$568 ( \1551 , \1546 , \1549 , \1550 );
xor \U$569 ( \1552 , \1356 , \1375 );
xor \U$570 ( \1553 , \1552 , \1379 );
and \U$571 ( \1554 , \1551 , \1553 );
xor \U$572 ( \1555 , \1462 , \1471 );
xor \U$573 ( \1556 , \1555 , \1474 );
and \U$574 ( \1557 , \1553 , \1556 );
and \U$575 ( \1558 , \1551 , \1556 );
or \U$576 ( \1559 , \1554 , \1557 , \1558 );
xor \U$577 ( \1560 , \1477 , \1479 );
xor \U$578 ( \1561 , \1560 , \1481 );
and \U$579 ( \1562 , \1559 , \1561 );
and \U$580 ( \1563 , \1490 , \1562 );
xor \U$581 ( \1564 , \1490 , \1562 );
xor \U$582 ( \1565 , \1559 , \1561 );
buf \U$583 ( \1566 , RIc0d7d80_16);
buf \U$584 ( \1567 , RIc0d7df8_17);
and \U$585 ( \1568 , \1566 , \1567 );
not \U$586 ( \1569 , \1568 );
and \U$587 ( \1570 , \1419 , \1569 );
not \U$588 ( \1571 , \1570 );
and \U$589 ( \1572 , \998 , \1494 );
and \U$590 ( \1573 , \984 , \1492 );
nor \U$591 ( \1574 , \1572 , \1573 );
xnor \U$592 ( \1575 , \1574 , \1422 );
and \U$593 ( \1576 , \1571 , \1575 );
and \U$594 ( \1577 , \1037 , \1360 );
and \U$595 ( \1578 , \1016 , \1358 );
nor \U$596 ( \1579 , \1577 , \1578 );
xnor \U$597 ( \1580 , \1579 , \1317 );
and \U$598 ( \1581 , \1575 , \1580 );
and \U$599 ( \1582 , \1571 , \1580 );
or \U$600 ( \1583 , \1576 , \1581 , \1582 );
and \U$601 ( \1584 , \1377 , \1028 );
and \U$602 ( \1585 , \1349 , \1026 );
nor \U$603 ( \1586 , \1584 , \1585 );
xnor \U$604 ( \1587 , \1586 , \1009 );
and \U$605 ( \1588 , \1531 , \991 );
and \U$606 ( \1589 , \1457 , \989 );
nor \U$607 ( \1590 , \1588 , \1589 );
xnor \U$608 ( \1591 , \1590 , \996 );
and \U$609 ( \1592 , \1587 , \1591 );
buf \U$610 ( \1593 , RIc0d9b08_79);
and \U$611 ( \1594 , \1593 , \985 );
and \U$612 ( \1595 , \1591 , \1594 );
and \U$613 ( \1596 , \1587 , \1594 );
or \U$614 ( \1597 , \1592 , \1595 , \1596 );
and \U$615 ( \1598 , \1583 , \1597 );
and \U$616 ( \1599 , \1093 , \1247 );
and \U$617 ( \1600 , \1085 , \1245 );
nor \U$618 ( \1601 , \1599 , \1600 );
xnor \U$619 ( \1602 , \1601 , \1198 );
and \U$620 ( \1603 , \1167 , \1146 );
and \U$621 ( \1604 , \1162 , \1144 );
nor \U$622 ( \1605 , \1603 , \1604 );
xnor \U$623 ( \1606 , \1605 , \1105 );
and \U$624 ( \1607 , \1602 , \1606 );
and \U$625 ( \1608 , \1272 , \1076 );
and \U$626 ( \1609 , \1221 , \1074 );
nor \U$627 ( \1610 , \1608 , \1609 );
xnor \U$628 ( \1611 , \1610 , \1046 );
and \U$629 ( \1612 , \1606 , \1611 );
and \U$630 ( \1613 , \1602 , \1611 );
or \U$631 ( \1614 , \1607 , \1612 , \1613 );
and \U$632 ( \1615 , \1597 , \1614 );
and \U$633 ( \1616 , \1583 , \1614 );
or \U$634 ( \1617 , \1598 , \1615 , \1616 );
xor \U$635 ( \1618 , \1497 , \1501 );
xor \U$636 ( \1619 , \1618 , \1506 );
xor \U$637 ( \1620 , \1513 , \1517 );
xor \U$638 ( \1621 , \1620 , \1522 );
and \U$639 ( \1622 , \1619 , \1621 );
xnor \U$640 ( \1623 , \1530 , \1532 );
and \U$641 ( \1624 , \1621 , \1623 );
and \U$642 ( \1625 , \1619 , \1623 );
or \U$643 ( \1626 , \1622 , \1624 , \1625 );
and \U$644 ( \1627 , \1617 , \1626 );
xor \U$645 ( \1628 , \1538 , \1540 );
xor \U$646 ( \1629 , \1628 , \1542 );
and \U$647 ( \1630 , \1626 , \1629 );
and \U$648 ( \1631 , \1617 , \1629 );
or \U$649 ( \1632 , \1627 , \1630 , \1631 );
xor \U$650 ( \1633 , \1435 , \1451 );
xor \U$651 ( \1634 , \1633 , \1459 );
and \U$652 ( \1635 , \1632 , \1634 );
xor \U$653 ( \1636 , \1536 , \1545 );
xor \U$654 ( \1637 , \1636 , \1548 );
and \U$655 ( \1638 , \1634 , \1637 );
and \U$656 ( \1639 , \1632 , \1637 );
or \U$657 ( \1640 , \1635 , \1638 , \1639 );
xor \U$658 ( \1641 , \1551 , \1553 );
xor \U$659 ( \1642 , \1641 , \1556 );
and \U$660 ( \1643 , \1640 , \1642 );
and \U$661 ( \1644 , \1565 , \1643 );
xor \U$662 ( \1645 , \1565 , \1643 );
xor \U$663 ( \1646 , \1640 , \1642 );
and \U$664 ( \1647 , \1457 , \1028 );
and \U$665 ( \1648 , \1377 , \1026 );
nor \U$666 ( \1649 , \1647 , \1648 );
xnor \U$667 ( \1650 , \1649 , \1009 );
and \U$668 ( \1651 , \1593 , \991 );
and \U$669 ( \1652 , \1531 , \989 );
nor \U$670 ( \1653 , \1651 , \1652 );
xnor \U$671 ( \1654 , \1653 , \996 );
and \U$672 ( \1655 , \1650 , \1654 );
buf \U$673 ( \1656 , RIc0d9b80_80);
and \U$674 ( \1657 , \1656 , \985 );
and \U$675 ( \1658 , \1654 , \1657 );
and \U$676 ( \1659 , \1650 , \1657 );
or \U$677 ( \1660 , \1655 , \1658 , \1659 );
xor \U$678 ( \1661 , \1419 , \1566 );
xor \U$679 ( \1662 , \1566 , \1567 );
not \U$680 ( \1663 , \1662 );
and \U$681 ( \1664 , \1661 , \1663 );
and \U$682 ( \1665 , \984 , \1664 );
not \U$683 ( \1666 , \1665 );
xnor \U$684 ( \1667 , \1666 , \1570 );
and \U$685 ( \1668 , \1016 , \1494 );
and \U$686 ( \1669 , \998 , \1492 );
nor \U$687 ( \1670 , \1668 , \1669 );
xnor \U$688 ( \1671 , \1670 , \1422 );
and \U$689 ( \1672 , \1667 , \1671 );
and \U$690 ( \1673 , \1085 , \1360 );
and \U$691 ( \1674 , \1037 , \1358 );
nor \U$692 ( \1675 , \1673 , \1674 );
xnor \U$693 ( \1676 , \1675 , \1317 );
and \U$694 ( \1677 , \1671 , \1676 );
and \U$695 ( \1678 , \1667 , \1676 );
or \U$696 ( \1679 , \1672 , \1677 , \1678 );
and \U$697 ( \1680 , \1660 , \1679 );
and \U$698 ( \1681 , \1162 , \1247 );
and \U$699 ( \1682 , \1093 , \1245 );
nor \U$700 ( \1683 , \1681 , \1682 );
xnor \U$701 ( \1684 , \1683 , \1198 );
and \U$702 ( \1685 , \1221 , \1146 );
and \U$703 ( \1686 , \1167 , \1144 );
nor \U$704 ( \1687 , \1685 , \1686 );
xnor \U$705 ( \1688 , \1687 , \1105 );
and \U$706 ( \1689 , \1684 , \1688 );
and \U$707 ( \1690 , \1349 , \1076 );
and \U$708 ( \1691 , \1272 , \1074 );
nor \U$709 ( \1692 , \1690 , \1691 );
xnor \U$710 ( \1693 , \1692 , \1046 );
and \U$711 ( \1694 , \1688 , \1693 );
and \U$712 ( \1695 , \1684 , \1693 );
or \U$713 ( \1696 , \1689 , \1694 , \1695 );
and \U$714 ( \1697 , \1679 , \1696 );
and \U$715 ( \1698 , \1660 , \1696 );
or \U$716 ( \1699 , \1680 , \1697 , \1698 );
xor \U$717 ( \1700 , \1571 , \1575 );
xor \U$718 ( \1701 , \1700 , \1580 );
xor \U$719 ( \1702 , \1587 , \1591 );
xor \U$720 ( \1703 , \1702 , \1594 );
and \U$721 ( \1704 , \1701 , \1703 );
xor \U$722 ( \1705 , \1602 , \1606 );
xor \U$723 ( \1706 , \1705 , \1611 );
and \U$724 ( \1707 , \1703 , \1706 );
and \U$725 ( \1708 , \1701 , \1706 );
or \U$726 ( \1709 , \1704 , \1707 , \1708 );
and \U$727 ( \1710 , \1699 , \1709 );
xor \U$728 ( \1711 , \1619 , \1621 );
xor \U$729 ( \1712 , \1711 , \1623 );
and \U$730 ( \1713 , \1709 , \1712 );
and \U$731 ( \1714 , \1699 , \1712 );
or \U$732 ( \1715 , \1710 , \1713 , \1714 );
xor \U$733 ( \1716 , \1509 , \1525 );
xor \U$734 ( \1717 , \1716 , \1533 );
and \U$735 ( \1718 , \1715 , \1717 );
xor \U$736 ( \1719 , \1617 , \1626 );
xor \U$737 ( \1720 , \1719 , \1629 );
and \U$738 ( \1721 , \1717 , \1720 );
and \U$739 ( \1722 , \1715 , \1720 );
or \U$740 ( \1723 , \1718 , \1721 , \1722 );
xor \U$741 ( \1724 , \1632 , \1634 );
xor \U$742 ( \1725 , \1724 , \1637 );
and \U$743 ( \1726 , \1723 , \1725 );
and \U$744 ( \1727 , \1646 , \1726 );
xor \U$745 ( \1728 , \1646 , \1726 );
xor \U$746 ( \1729 , \1723 , \1725 );
and \U$747 ( \1730 , \1093 , \1360 );
and \U$748 ( \1731 , \1085 , \1358 );
nor \U$749 ( \1732 , \1730 , \1731 );
xnor \U$750 ( \1733 , \1732 , \1317 );
and \U$751 ( \1734 , \1167 , \1247 );
and \U$752 ( \1735 , \1162 , \1245 );
nor \U$753 ( \1736 , \1734 , \1735 );
xnor \U$754 ( \1737 , \1736 , \1198 );
and \U$755 ( \1738 , \1733 , \1737 );
and \U$756 ( \1739 , \1272 , \1146 );
and \U$757 ( \1740 , \1221 , \1144 );
nor \U$758 ( \1741 , \1739 , \1740 );
xnor \U$759 ( \1742 , \1741 , \1105 );
and \U$760 ( \1743 , \1737 , \1742 );
and \U$761 ( \1744 , \1733 , \1742 );
or \U$762 ( \1745 , \1738 , \1743 , \1744 );
buf \U$763 ( \1746 , RIc0d7e70_18);
buf \U$764 ( \1747 , RIc0d7ee8_19);
and \U$765 ( \1748 , \1746 , \1747 );
not \U$766 ( \1749 , \1748 );
and \U$767 ( \1750 , \1567 , \1749 );
not \U$768 ( \1751 , \1750 );
and \U$769 ( \1752 , \998 , \1664 );
and \U$770 ( \1753 , \984 , \1662 );
nor \U$771 ( \1754 , \1752 , \1753 );
xnor \U$772 ( \1755 , \1754 , \1570 );
and \U$773 ( \1756 , \1751 , \1755 );
and \U$774 ( \1757 , \1037 , \1494 );
and \U$775 ( \1758 , \1016 , \1492 );
nor \U$776 ( \1759 , \1757 , \1758 );
xnor \U$777 ( \1760 , \1759 , \1422 );
and \U$778 ( \1761 , \1755 , \1760 );
and \U$779 ( \1762 , \1751 , \1760 );
or \U$780 ( \1763 , \1756 , \1761 , \1762 );
and \U$781 ( \1764 , \1745 , \1763 );
and \U$782 ( \1765 , \1377 , \1076 );
and \U$783 ( \1766 , \1349 , \1074 );
nor \U$784 ( \1767 , \1765 , \1766 );
xnor \U$785 ( \1768 , \1767 , \1046 );
and \U$786 ( \1769 , \1531 , \1028 );
and \U$787 ( \1770 , \1457 , \1026 );
nor \U$788 ( \1771 , \1769 , \1770 );
xnor \U$789 ( \1772 , \1771 , \1009 );
and \U$790 ( \1773 , \1768 , \1772 );
and \U$791 ( \1774 , \1656 , \991 );
and \U$792 ( \1775 , \1593 , \989 );
nor \U$793 ( \1776 , \1774 , \1775 );
xnor \U$794 ( \1777 , \1776 , \996 );
and \U$795 ( \1778 , \1772 , \1777 );
and \U$796 ( \1779 , \1768 , \1777 );
or \U$797 ( \1780 , \1773 , \1778 , \1779 );
and \U$798 ( \1781 , \1763 , \1780 );
and \U$799 ( \1782 , \1745 , \1780 );
or \U$800 ( \1783 , \1764 , \1781 , \1782 );
xor \U$801 ( \1784 , \1650 , \1654 );
xor \U$802 ( \1785 , \1784 , \1657 );
xor \U$803 ( \1786 , \1684 , \1688 );
xor \U$804 ( \1787 , \1786 , \1693 );
or \U$805 ( \1788 , \1785 , \1787 );
and \U$806 ( \1789 , \1783 , \1788 );
xor \U$807 ( \1790 , \1701 , \1703 );
xor \U$808 ( \1791 , \1790 , \1706 );
and \U$809 ( \1792 , \1788 , \1791 );
and \U$810 ( \1793 , \1783 , \1791 );
or \U$811 ( \1794 , \1789 , \1792 , \1793 );
xor \U$812 ( \1795 , \1583 , \1597 );
xor \U$813 ( \1796 , \1795 , \1614 );
and \U$814 ( \1797 , \1794 , \1796 );
xor \U$815 ( \1798 , \1699 , \1709 );
xor \U$816 ( \1799 , \1798 , \1712 );
and \U$817 ( \1800 , \1796 , \1799 );
and \U$818 ( \1801 , \1794 , \1799 );
or \U$819 ( \1802 , \1797 , \1800 , \1801 );
xor \U$820 ( \1803 , \1715 , \1717 );
xor \U$821 ( \1804 , \1803 , \1720 );
and \U$822 ( \1805 , \1802 , \1804 );
and \U$823 ( \1806 , \1729 , \1805 );
xor \U$824 ( \1807 , \1729 , \1805 );
xor \U$825 ( \1808 , \1802 , \1804 );
and \U$826 ( \1809 , \1162 , \1360 );
and \U$827 ( \1810 , \1093 , \1358 );
nor \U$828 ( \1811 , \1809 , \1810 );
xnor \U$829 ( \1812 , \1811 , \1317 );
and \U$830 ( \1813 , \1221 , \1247 );
and \U$831 ( \1814 , \1167 , \1245 );
nor \U$832 ( \1815 , \1813 , \1814 );
xnor \U$833 ( \1816 , \1815 , \1198 );
and \U$834 ( \1817 , \1812 , \1816 );
and \U$835 ( \1818 , \1349 , \1146 );
and \U$836 ( \1819 , \1272 , \1144 );
nor \U$837 ( \1820 , \1818 , \1819 );
xnor \U$838 ( \1821 , \1820 , \1105 );
and \U$839 ( \1822 , \1816 , \1821 );
and \U$840 ( \1823 , \1812 , \1821 );
or \U$841 ( \1824 , \1817 , \1822 , \1823 );
xor \U$842 ( \1825 , \1567 , \1746 );
xor \U$843 ( \1826 , \1746 , \1747 );
not \U$844 ( \1827 , \1826 );
and \U$845 ( \1828 , \1825 , \1827 );
and \U$846 ( \1829 , \984 , \1828 );
not \U$847 ( \1830 , \1829 );
xnor \U$848 ( \1831 , \1830 , \1750 );
and \U$849 ( \1832 , \1016 , \1664 );
and \U$850 ( \1833 , \998 , \1662 );
nor \U$851 ( \1834 , \1832 , \1833 );
xnor \U$852 ( \1835 , \1834 , \1570 );
and \U$853 ( \1836 , \1831 , \1835 );
and \U$854 ( \1837 , \1085 , \1494 );
and \U$855 ( \1838 , \1037 , \1492 );
nor \U$856 ( \1839 , \1837 , \1838 );
xnor \U$857 ( \1840 , \1839 , \1422 );
and \U$858 ( \1841 , \1835 , \1840 );
and \U$859 ( \1842 , \1831 , \1840 );
or \U$860 ( \1843 , \1836 , \1841 , \1842 );
and \U$861 ( \1844 , \1824 , \1843 );
and \U$862 ( \1845 , \1457 , \1076 );
and \U$863 ( \1846 , \1377 , \1074 );
nor \U$864 ( \1847 , \1845 , \1846 );
xnor \U$865 ( \1848 , \1847 , \1046 );
and \U$866 ( \1849 , \1593 , \1028 );
and \U$867 ( \1850 , \1531 , \1026 );
nor \U$868 ( \1851 , \1849 , \1850 );
xnor \U$869 ( \1852 , \1851 , \1009 );
and \U$870 ( \1853 , \1848 , \1852 );
buf \U$871 ( \1854 , RIc0d9bf8_81);
and \U$872 ( \1855 , \1854 , \991 );
and \U$873 ( \1856 , \1656 , \989 );
nor \U$874 ( \1857 , \1855 , \1856 );
xnor \U$875 ( \1858 , \1857 , \996 );
and \U$876 ( \1859 , \1852 , \1858 );
and \U$877 ( \1860 , \1848 , \1858 );
or \U$878 ( \1861 , \1853 , \1859 , \1860 );
and \U$879 ( \1862 , \1843 , \1861 );
and \U$880 ( \1863 , \1824 , \1861 );
or \U$881 ( \1864 , \1844 , \1862 , \1863 );
and \U$882 ( \1865 , \1854 , \985 );
xor \U$883 ( \1866 , \1733 , \1737 );
xor \U$884 ( \1867 , \1866 , \1742 );
and \U$885 ( \1868 , \1865 , \1867 );
xor \U$886 ( \1869 , \1768 , \1772 );
xor \U$887 ( \1870 , \1869 , \1777 );
and \U$888 ( \1871 , \1867 , \1870 );
and \U$889 ( \1872 , \1865 , \1870 );
or \U$890 ( \1873 , \1868 , \1871 , \1872 );
and \U$891 ( \1874 , \1864 , \1873 );
xor \U$892 ( \1875 , \1667 , \1671 );
xor \U$893 ( \1876 , \1875 , \1676 );
and \U$894 ( \1877 , \1873 , \1876 );
and \U$895 ( \1878 , \1864 , \1876 );
or \U$896 ( \1879 , \1874 , \1877 , \1878 );
xor \U$897 ( \1880 , \1660 , \1679 );
xor \U$898 ( \1881 , \1880 , \1696 );
and \U$899 ( \1882 , \1879 , \1881 );
xor \U$900 ( \1883 , \1783 , \1788 );
xor \U$901 ( \1884 , \1883 , \1791 );
and \U$902 ( \1885 , \1881 , \1884 );
and \U$903 ( \1886 , \1879 , \1884 );
or \U$904 ( \1887 , \1882 , \1885 , \1886 );
buf \U$905 ( \1888 , RIc0d7f60_20);
buf \U$906 ( \1889 , RIc0d7fd8_21);
and \U$907 ( \1890 , \1888 , \1889 );
not \U$908 ( \1891 , \1890 );
and \U$909 ( \1892 , \1747 , \1891 );
not \U$910 ( \1893 , \1892 );
and \U$911 ( \1894 , \998 , \1828 );
and \U$912 ( \1895 , \984 , \1826 );
nor \U$913 ( \1896 , \1894 , \1895 );
xnor \U$914 ( \1897 , \1896 , \1750 );
and \U$915 ( \1898 , \1893 , \1897 );
and \U$916 ( \1899 , \1037 , \1664 );
and \U$917 ( \1900 , \1016 , \1662 );
nor \U$918 ( \1901 , \1899 , \1900 );
xnor \U$919 ( \1902 , \1901 , \1570 );
and \U$920 ( \1903 , \1897 , \1902 );
and \U$921 ( \1904 , \1893 , \1902 );
or \U$922 ( \1905 , \1898 , \1903 , \1904 );
and \U$923 ( \1906 , \1093 , \1494 );
and \U$924 ( \1907 , \1085 , \1492 );
nor \U$925 ( \1908 , \1906 , \1907 );
xnor \U$926 ( \1909 , \1908 , \1422 );
and \U$927 ( \1910 , \1167 , \1360 );
and \U$928 ( \1911 , \1162 , \1358 );
nor \U$929 ( \1912 , \1910 , \1911 );
xnor \U$930 ( \1913 , \1912 , \1317 );
and \U$931 ( \1914 , \1909 , \1913 );
and \U$932 ( \1915 , \1272 , \1247 );
and \U$933 ( \1916 , \1221 , \1245 );
nor \U$934 ( \1917 , \1915 , \1916 );
xnor \U$935 ( \1918 , \1917 , \1198 );
and \U$936 ( \1919 , \1913 , \1918 );
and \U$937 ( \1920 , \1909 , \1918 );
or \U$938 ( \1921 , \1914 , \1919 , \1920 );
and \U$939 ( \1922 , \1905 , \1921 );
and \U$940 ( \1923 , \1377 , \1146 );
and \U$941 ( \1924 , \1349 , \1144 );
nor \U$942 ( \1925 , \1923 , \1924 );
xnor \U$943 ( \1926 , \1925 , \1105 );
and \U$944 ( \1927 , \1531 , \1076 );
and \U$945 ( \1928 , \1457 , \1074 );
nor \U$946 ( \1929 , \1927 , \1928 );
xnor \U$947 ( \1930 , \1929 , \1046 );
and \U$948 ( \1931 , \1926 , \1930 );
and \U$949 ( \1932 , \1656 , \1028 );
and \U$950 ( \1933 , \1593 , \1026 );
nor \U$951 ( \1934 , \1932 , \1933 );
xnor \U$952 ( \1935 , \1934 , \1009 );
and \U$953 ( \1936 , \1930 , \1935 );
and \U$954 ( \1937 , \1926 , \1935 );
or \U$955 ( \1938 , \1931 , \1936 , \1937 );
and \U$956 ( \1939 , \1921 , \1938 );
and \U$957 ( \1940 , \1905 , \1938 );
or \U$958 ( \1941 , \1922 , \1939 , \1940 );
buf \U$959 ( \1942 , RIc0d9c70_82);
and \U$960 ( \1943 , \1942 , \985 );
xor \U$961 ( \1944 , \1848 , \1852 );
xor \U$962 ( \1945 , \1944 , \1858 );
or \U$963 ( \1946 , \1943 , \1945 );
and \U$964 ( \1947 , \1941 , \1946 );
xor \U$965 ( \1948 , \1812 , \1816 );
xor \U$966 ( \1949 , \1948 , \1821 );
xor \U$967 ( \1950 , \1831 , \1835 );
xor \U$968 ( \1951 , \1950 , \1840 );
and \U$969 ( \1952 , \1949 , \1951 );
and \U$970 ( \1953 , \1946 , \1952 );
and \U$971 ( \1954 , \1941 , \1952 );
or \U$972 ( \1955 , \1947 , \1953 , \1954 );
xor \U$973 ( \1956 , \1751 , \1755 );
xor \U$974 ( \1957 , \1956 , \1760 );
xor \U$975 ( \1958 , \1824 , \1843 );
xor \U$976 ( \1959 , \1958 , \1861 );
and \U$977 ( \1960 , \1957 , \1959 );
xor \U$978 ( \1961 , \1865 , \1867 );
xor \U$979 ( \1962 , \1961 , \1870 );
and \U$980 ( \1963 , \1959 , \1962 );
and \U$981 ( \1964 , \1957 , \1962 );
or \U$982 ( \1965 , \1960 , \1963 , \1964 );
and \U$983 ( \1966 , \1955 , \1965 );
xnor \U$984 ( \1967 , \1785 , \1787 );
and \U$985 ( \1968 , \1965 , \1967 );
and \U$986 ( \1969 , \1955 , \1967 );
or \U$987 ( \1970 , \1966 , \1968 , \1969 );
xor \U$988 ( \1971 , \1745 , \1763 );
xor \U$989 ( \1972 , \1971 , \1780 );
xor \U$990 ( \1973 , \1864 , \1873 );
xor \U$991 ( \1974 , \1973 , \1876 );
and \U$992 ( \1975 , \1972 , \1974 );
and \U$993 ( \1976 , \1970 , \1975 );
xor \U$994 ( \1977 , \1879 , \1881 );
xor \U$995 ( \1978 , \1977 , \1884 );
and \U$996 ( \1979 , \1975 , \1978 );
and \U$997 ( \1980 , \1970 , \1978 );
or \U$998 ( \1981 , \1976 , \1979 , \1980 );
and \U$999 ( \1982 , \1887 , \1981 );
xor \U$1000 ( \1983 , \1794 , \1796 );
xor \U$1001 ( \1984 , \1983 , \1799 );
and \U$1002 ( \1985 , \1981 , \1984 );
and \U$1003 ( \1986 , \1887 , \1984 );
or \U$1004 ( \1987 , \1982 , \1985 , \1986 );
and \U$1005 ( \1988 , \1808 , \1987 );
xor \U$1006 ( \1989 , \1808 , \1987 );
xor \U$1007 ( \1990 , \1887 , \1981 );
xor \U$1008 ( \1991 , \1990 , \1984 );
and \U$1009 ( \1992 , \1457 , \1146 );
and \U$1010 ( \1993 , \1377 , \1144 );
nor \U$1011 ( \1994 , \1992 , \1993 );
xnor \U$1012 ( \1995 , \1994 , \1105 );
and \U$1013 ( \1996 , \1593 , \1076 );
and \U$1014 ( \1997 , \1531 , \1074 );
nor \U$1015 ( \1998 , \1996 , \1997 );
xnor \U$1016 ( \1999 , \1998 , \1046 );
and \U$1017 ( \2000 , \1995 , \1999 );
and \U$1018 ( \2001 , \1854 , \1028 );
and \U$1019 ( \2002 , \1656 , \1026 );
nor \U$1020 ( \2003 , \2001 , \2002 );
xnor \U$1021 ( \2004 , \2003 , \1009 );
and \U$1022 ( \2005 , \1999 , \2004 );
and \U$1023 ( \2006 , \1995 , \2004 );
or \U$1024 ( \2007 , \2000 , \2005 , \2006 );
and \U$1025 ( \2008 , \1162 , \1494 );
and \U$1026 ( \2009 , \1093 , \1492 );
nor \U$1027 ( \2010 , \2008 , \2009 );
xnor \U$1028 ( \2011 , \2010 , \1422 );
and \U$1029 ( \2012 , \1221 , \1360 );
and \U$1030 ( \2013 , \1167 , \1358 );
nor \U$1031 ( \2014 , \2012 , \2013 );
xnor \U$1032 ( \2015 , \2014 , \1317 );
and \U$1033 ( \2016 , \2011 , \2015 );
and \U$1034 ( \2017 , \1349 , \1247 );
and \U$1035 ( \2018 , \1272 , \1245 );
nor \U$1036 ( \2019 , \2017 , \2018 );
xnor \U$1037 ( \2020 , \2019 , \1198 );
and \U$1038 ( \2021 , \2015 , \2020 );
and \U$1039 ( \2022 , \2011 , \2020 );
or \U$1040 ( \2023 , \2016 , \2021 , \2022 );
and \U$1041 ( \2024 , \2007 , \2023 );
xor \U$1042 ( \2025 , \1747 , \1888 );
xor \U$1043 ( \2026 , \1888 , \1889 );
not \U$1044 ( \2027 , \2026 );
and \U$1045 ( \2028 , \2025 , \2027 );
and \U$1046 ( \2029 , \984 , \2028 );
not \U$1047 ( \2030 , \2029 );
xnor \U$1048 ( \2031 , \2030 , \1892 );
and \U$1049 ( \2032 , \1016 , \1828 );
and \U$1050 ( \2033 , \998 , \1826 );
nor \U$1051 ( \2034 , \2032 , \2033 );
xnor \U$1052 ( \2035 , \2034 , \1750 );
and \U$1053 ( \2036 , \2031 , \2035 );
and \U$1054 ( \2037 , \1085 , \1664 );
and \U$1055 ( \2038 , \1037 , \1662 );
nor \U$1056 ( \2039 , \2037 , \2038 );
xnor \U$1057 ( \2040 , \2039 , \1570 );
and \U$1058 ( \2041 , \2035 , \2040 );
and \U$1059 ( \2042 , \2031 , \2040 );
or \U$1060 ( \2043 , \2036 , \2041 , \2042 );
and \U$1061 ( \2044 , \2023 , \2043 );
and \U$1062 ( \2045 , \2007 , \2043 );
or \U$1063 ( \2046 , \2024 , \2044 , \2045 );
buf \U$1064 ( \2047 , RIc0d9ce8_83);
and \U$1065 ( \2048 , \2047 , \991 );
and \U$1066 ( \2049 , \1942 , \989 );
nor \U$1067 ( \2050 , \2048 , \2049 );
xnor \U$1068 ( \2051 , \2050 , \996 );
buf \U$1069 ( \2052 , RIc0d9d60_84);
and \U$1070 ( \2053 , \2052 , \985 );
or \U$1071 ( \2054 , \2051 , \2053 );
and \U$1072 ( \2055 , \1942 , \991 );
and \U$1073 ( \2056 , \1854 , \989 );
nor \U$1074 ( \2057 , \2055 , \2056 );
xnor \U$1075 ( \2058 , \2057 , \996 );
and \U$1076 ( \2059 , \2054 , \2058 );
and \U$1077 ( \2060 , \2047 , \985 );
and \U$1078 ( \2061 , \2058 , \2060 );
and \U$1079 ( \2062 , \2054 , \2060 );
or \U$1080 ( \2063 , \2059 , \2061 , \2062 );
and \U$1081 ( \2064 , \2046 , \2063 );
xor \U$1082 ( \2065 , \1893 , \1897 );
xor \U$1083 ( \2066 , \2065 , \1902 );
xor \U$1084 ( \2067 , \1909 , \1913 );
xor \U$1085 ( \2068 , \2067 , \1918 );
and \U$1086 ( \2069 , \2066 , \2068 );
xor \U$1087 ( \2070 , \1926 , \1930 );
xor \U$1088 ( \2071 , \2070 , \1935 );
and \U$1089 ( \2072 , \2068 , \2071 );
and \U$1090 ( \2073 , \2066 , \2071 );
or \U$1091 ( \2074 , \2069 , \2072 , \2073 );
and \U$1092 ( \2075 , \2063 , \2074 );
and \U$1093 ( \2076 , \2046 , \2074 );
or \U$1094 ( \2077 , \2064 , \2075 , \2076 );
xor \U$1095 ( \2078 , \1905 , \1921 );
xor \U$1096 ( \2079 , \2078 , \1938 );
xnor \U$1097 ( \2080 , \1943 , \1945 );
and \U$1098 ( \2081 , \2079 , \2080 );
xor \U$1099 ( \2082 , \1949 , \1951 );
and \U$1100 ( \2083 , \2080 , \2082 );
and \U$1101 ( \2084 , \2079 , \2082 );
or \U$1102 ( \2085 , \2081 , \2083 , \2084 );
and \U$1103 ( \2086 , \2077 , \2085 );
xor \U$1104 ( \2087 , \1957 , \1959 );
xor \U$1105 ( \2088 , \2087 , \1962 );
and \U$1106 ( \2089 , \2085 , \2088 );
and \U$1107 ( \2090 , \2077 , \2088 );
or \U$1108 ( \2091 , \2086 , \2089 , \2090 );
xor \U$1109 ( \2092 , \1955 , \1965 );
xor \U$1110 ( \2093 , \2092 , \1967 );
and \U$1111 ( \2094 , \2091 , \2093 );
xor \U$1112 ( \2095 , \1972 , \1974 );
and \U$1113 ( \2096 , \2093 , \2095 );
and \U$1114 ( \2097 , \2091 , \2095 );
or \U$1115 ( \2098 , \2094 , \2096 , \2097 );
xor \U$1116 ( \2099 , \1970 , \1975 );
xor \U$1117 ( \2100 , \2099 , \1978 );
and \U$1118 ( \2101 , \2098 , \2100 );
and \U$1119 ( \2102 , \1991 , \2101 );
xor \U$1120 ( \2103 , \1991 , \2101 );
xor \U$1121 ( \2104 , \2098 , \2100 );
buf \U$1122 ( \2105 , RIc0d8050_22);
buf \U$1123 ( \2106 , RIc0d80c8_23);
and \U$1124 ( \2107 , \2105 , \2106 );
not \U$1125 ( \2108 , \2107 );
and \U$1126 ( \2109 , \1889 , \2108 );
not \U$1127 ( \2110 , \2109 );
and \U$1128 ( \2111 , \998 , \2028 );
and \U$1129 ( \2112 , \984 , \2026 );
nor \U$1130 ( \2113 , \2111 , \2112 );
xnor \U$1131 ( \2114 , \2113 , \1892 );
and \U$1132 ( \2115 , \2110 , \2114 );
and \U$1133 ( \2116 , \1037 , \1828 );
and \U$1134 ( \2117 , \1016 , \1826 );
nor \U$1135 ( \2118 , \2116 , \2117 );
xnor \U$1136 ( \2119 , \2118 , \1750 );
and \U$1137 ( \2120 , \2114 , \2119 );
and \U$1138 ( \2121 , \2110 , \2119 );
or \U$1139 ( \2122 , \2115 , \2120 , \2121 );
and \U$1140 ( \2123 , \1377 , \1247 );
and \U$1141 ( \2124 , \1349 , \1245 );
nor \U$1142 ( \2125 , \2123 , \2124 );
xnor \U$1143 ( \2126 , \2125 , \1198 );
and \U$1144 ( \2127 , \1531 , \1146 );
and \U$1145 ( \2128 , \1457 , \1144 );
nor \U$1146 ( \2129 , \2127 , \2128 );
xnor \U$1147 ( \2130 , \2129 , \1105 );
and \U$1148 ( \2131 , \2126 , \2130 );
and \U$1149 ( \2132 , \1656 , \1076 );
and \U$1150 ( \2133 , \1593 , \1074 );
nor \U$1151 ( \2134 , \2132 , \2133 );
xnor \U$1152 ( \2135 , \2134 , \1046 );
and \U$1153 ( \2136 , \2130 , \2135 );
and \U$1154 ( \2137 , \2126 , \2135 );
or \U$1155 ( \2138 , \2131 , \2136 , \2137 );
and \U$1156 ( \2139 , \2122 , \2138 );
and \U$1157 ( \2140 , \1093 , \1664 );
and \U$1158 ( \2141 , \1085 , \1662 );
nor \U$1159 ( \2142 , \2140 , \2141 );
xnor \U$1160 ( \2143 , \2142 , \1570 );
and \U$1161 ( \2144 , \1167 , \1494 );
and \U$1162 ( \2145 , \1162 , \1492 );
nor \U$1163 ( \2146 , \2144 , \2145 );
xnor \U$1164 ( \2147 , \2146 , \1422 );
and \U$1165 ( \2148 , \2143 , \2147 );
and \U$1166 ( \2149 , \1272 , \1360 );
and \U$1167 ( \2150 , \1221 , \1358 );
nor \U$1168 ( \2151 , \2149 , \2150 );
xnor \U$1169 ( \2152 , \2151 , \1317 );
and \U$1170 ( \2153 , \2147 , \2152 );
and \U$1171 ( \2154 , \2143 , \2152 );
or \U$1172 ( \2155 , \2148 , \2153 , \2154 );
and \U$1173 ( \2156 , \2138 , \2155 );
and \U$1174 ( \2157 , \2122 , \2155 );
or \U$1175 ( \2158 , \2139 , \2156 , \2157 );
and \U$1176 ( \2159 , \1942 , \1028 );
and \U$1177 ( \2160 , \1854 , \1026 );
nor \U$1178 ( \2161 , \2159 , \2160 );
xnor \U$1179 ( \2162 , \2161 , \1009 );
and \U$1180 ( \2163 , \2052 , \991 );
and \U$1181 ( \2164 , \2047 , \989 );
nor \U$1182 ( \2165 , \2163 , \2164 );
xnor \U$1183 ( \2166 , \2165 , \996 );
and \U$1184 ( \2167 , \2162 , \2166 );
buf \U$1185 ( \2168 , RIc0d9dd8_85);
and \U$1186 ( \2169 , \2168 , \985 );
and \U$1187 ( \2170 , \2166 , \2169 );
and \U$1188 ( \2171 , \2162 , \2169 );
or \U$1189 ( \2172 , \2167 , \2170 , \2171 );
xor \U$1190 ( \2173 , \1995 , \1999 );
xor \U$1191 ( \2174 , \2173 , \2004 );
and \U$1192 ( \2175 , \2172 , \2174 );
xnor \U$1193 ( \2176 , \2051 , \2053 );
and \U$1194 ( \2177 , \2174 , \2176 );
and \U$1195 ( \2178 , \2172 , \2176 );
or \U$1196 ( \2179 , \2175 , \2177 , \2178 );
and \U$1197 ( \2180 , \2158 , \2179 );
xor \U$1198 ( \2181 , \2011 , \2015 );
xor \U$1199 ( \2182 , \2181 , \2020 );
xor \U$1200 ( \2183 , \2031 , \2035 );
xor \U$1201 ( \2184 , \2183 , \2040 );
and \U$1202 ( \2185 , \2182 , \2184 );
and \U$1203 ( \2186 , \2179 , \2185 );
and \U$1204 ( \2187 , \2158 , \2185 );
or \U$1205 ( \2188 , \2180 , \2186 , \2187 );
xor \U$1206 ( \2189 , \2007 , \2023 );
xor \U$1207 ( \2190 , \2189 , \2043 );
xor \U$1208 ( \2191 , \2054 , \2058 );
xor \U$1209 ( \2192 , \2191 , \2060 );
and \U$1210 ( \2193 , \2190 , \2192 );
xor \U$1211 ( \2194 , \2066 , \2068 );
xor \U$1212 ( \2195 , \2194 , \2071 );
and \U$1213 ( \2196 , \2192 , \2195 );
and \U$1214 ( \2197 , \2190 , \2195 );
or \U$1215 ( \2198 , \2193 , \2196 , \2197 );
and \U$1216 ( \2199 , \2188 , \2198 );
xor \U$1217 ( \2200 , \2079 , \2080 );
xor \U$1218 ( \2201 , \2200 , \2082 );
and \U$1219 ( \2202 , \2198 , \2201 );
and \U$1220 ( \2203 , \2188 , \2201 );
or \U$1221 ( \2204 , \2199 , \2202 , \2203 );
xor \U$1222 ( \2205 , \1941 , \1946 );
xor \U$1223 ( \2206 , \2205 , \1952 );
and \U$1224 ( \2207 , \2204 , \2206 );
xor \U$1225 ( \2208 , \2077 , \2085 );
xor \U$1226 ( \2209 , \2208 , \2088 );
and \U$1227 ( \2210 , \2206 , \2209 );
and \U$1228 ( \2211 , \2204 , \2209 );
or \U$1229 ( \2212 , \2207 , \2210 , \2211 );
xor \U$1230 ( \2213 , \2091 , \2093 );
xor \U$1231 ( \2214 , \2213 , \2095 );
and \U$1232 ( \2215 , \2212 , \2214 );
and \U$1233 ( \2216 , \2104 , \2215 );
xor \U$1234 ( \2217 , \2104 , \2215 );
xor \U$1235 ( \2218 , \2212 , \2214 );
xor \U$1236 ( \2219 , \1889 , \2105 );
xor \U$1237 ( \2220 , \2105 , \2106 );
not \U$1238 ( \2221 , \2220 );
and \U$1239 ( \2222 , \2219 , \2221 );
and \U$1240 ( \2223 , \984 , \2222 );
not \U$1241 ( \2224 , \2223 );
xnor \U$1242 ( \2225 , \2224 , \2109 );
and \U$1243 ( \2226 , \1016 , \2028 );
and \U$1244 ( \2227 , \998 , \2026 );
nor \U$1245 ( \2228 , \2226 , \2227 );
xnor \U$1246 ( \2229 , \2228 , \1892 );
and \U$1247 ( \2230 , \2225 , \2229 );
and \U$1248 ( \2231 , \1085 , \1828 );
and \U$1249 ( \2232 , \1037 , \1826 );
nor \U$1250 ( \2233 , \2231 , \2232 );
xnor \U$1251 ( \2234 , \2233 , \1750 );
and \U$1252 ( \2235 , \2229 , \2234 );
and \U$1253 ( \2236 , \2225 , \2234 );
or \U$1254 ( \2237 , \2230 , \2235 , \2236 );
and \U$1255 ( \2238 , \1457 , \1247 );
and \U$1256 ( \2239 , \1377 , \1245 );
nor \U$1257 ( \2240 , \2238 , \2239 );
xnor \U$1258 ( \2241 , \2240 , \1198 );
and \U$1259 ( \2242 , \1593 , \1146 );
and \U$1260 ( \2243 , \1531 , \1144 );
nor \U$1261 ( \2244 , \2242 , \2243 );
xnor \U$1262 ( \2245 , \2244 , \1105 );
and \U$1263 ( \2246 , \2241 , \2245 );
and \U$1264 ( \2247 , \1854 , \1076 );
and \U$1265 ( \2248 , \1656 , \1074 );
nor \U$1266 ( \2249 , \2247 , \2248 );
xnor \U$1267 ( \2250 , \2249 , \1046 );
and \U$1268 ( \2251 , \2245 , \2250 );
and \U$1269 ( \2252 , \2241 , \2250 );
or \U$1270 ( \2253 , \2246 , \2251 , \2252 );
and \U$1271 ( \2254 , \2237 , \2253 );
and \U$1272 ( \2255 , \1162 , \1664 );
and \U$1273 ( \2256 , \1093 , \1662 );
nor \U$1274 ( \2257 , \2255 , \2256 );
xnor \U$1275 ( \2258 , \2257 , \1570 );
and \U$1276 ( \2259 , \1221 , \1494 );
and \U$1277 ( \2260 , \1167 , \1492 );
nor \U$1278 ( \2261 , \2259 , \2260 );
xnor \U$1279 ( \2262 , \2261 , \1422 );
and \U$1280 ( \2263 , \2258 , \2262 );
and \U$1281 ( \2264 , \1349 , \1360 );
and \U$1282 ( \2265 , \1272 , \1358 );
nor \U$1283 ( \2266 , \2264 , \2265 );
xnor \U$1284 ( \2267 , \2266 , \1317 );
and \U$1285 ( \2268 , \2262 , \2267 );
and \U$1286 ( \2269 , \2258 , \2267 );
or \U$1287 ( \2270 , \2263 , \2268 , \2269 );
and \U$1288 ( \2271 , \2253 , \2270 );
and \U$1289 ( \2272 , \2237 , \2270 );
or \U$1290 ( \2273 , \2254 , \2271 , \2272 );
and \U$1291 ( \2274 , \2047 , \1028 );
and \U$1292 ( \2275 , \1942 , \1026 );
nor \U$1293 ( \2276 , \2274 , \2275 );
xnor \U$1294 ( \2277 , \2276 , \1009 );
and \U$1295 ( \2278 , \2168 , \991 );
and \U$1296 ( \2279 , \2052 , \989 );
nor \U$1297 ( \2280 , \2278 , \2279 );
xnor \U$1298 ( \2281 , \2280 , \996 );
and \U$1299 ( \2282 , \2277 , \2281 );
buf \U$1300 ( \2283 , RIc0d9e50_86);
and \U$1301 ( \2284 , \2283 , \985 );
and \U$1302 ( \2285 , \2281 , \2284 );
and \U$1303 ( \2286 , \2277 , \2284 );
or \U$1304 ( \2287 , \2282 , \2285 , \2286 );
xor \U$1305 ( \2288 , \2162 , \2166 );
xor \U$1306 ( \2289 , \2288 , \2169 );
and \U$1307 ( \2290 , \2287 , \2289 );
xor \U$1308 ( \2291 , \2126 , \2130 );
xor \U$1309 ( \2292 , \2291 , \2135 );
and \U$1310 ( \2293 , \2289 , \2292 );
and \U$1311 ( \2294 , \2287 , \2292 );
or \U$1312 ( \2295 , \2290 , \2293 , \2294 );
and \U$1313 ( \2296 , \2273 , \2295 );
xor \U$1314 ( \2297 , \2110 , \2114 );
xor \U$1315 ( \2298 , \2297 , \2119 );
xor \U$1316 ( \2299 , \2143 , \2147 );
xor \U$1317 ( \2300 , \2299 , \2152 );
and \U$1318 ( \2301 , \2298 , \2300 );
and \U$1319 ( \2302 , \2295 , \2301 );
and \U$1320 ( \2303 , \2273 , \2301 );
or \U$1321 ( \2304 , \2296 , \2302 , \2303 );
xor \U$1322 ( \2305 , \2122 , \2138 );
xor \U$1323 ( \2306 , \2305 , \2155 );
xor \U$1324 ( \2307 , \2172 , \2174 );
xor \U$1325 ( \2308 , \2307 , \2176 );
and \U$1326 ( \2309 , \2306 , \2308 );
xor \U$1327 ( \2310 , \2182 , \2184 );
and \U$1328 ( \2311 , \2308 , \2310 );
and \U$1329 ( \2312 , \2306 , \2310 );
or \U$1330 ( \2313 , \2309 , \2311 , \2312 );
and \U$1331 ( \2314 , \2304 , \2313 );
xor \U$1332 ( \2315 , \2190 , \2192 );
xor \U$1333 ( \2316 , \2315 , \2195 );
and \U$1334 ( \2317 , \2313 , \2316 );
and \U$1335 ( \2318 , \2304 , \2316 );
or \U$1336 ( \2319 , \2314 , \2317 , \2318 );
xor \U$1337 ( \2320 , \2046 , \2063 );
xor \U$1338 ( \2321 , \2320 , \2074 );
and \U$1339 ( \2322 , \2319 , \2321 );
xor \U$1340 ( \2323 , \2188 , \2198 );
xor \U$1341 ( \2324 , \2323 , \2201 );
and \U$1342 ( \2325 , \2321 , \2324 );
and \U$1343 ( \2326 , \2319 , \2324 );
or \U$1344 ( \2327 , \2322 , \2325 , \2326 );
xor \U$1345 ( \2328 , \2204 , \2206 );
xor \U$1346 ( \2329 , \2328 , \2209 );
and \U$1347 ( \2330 , \2327 , \2329 );
and \U$1348 ( \2331 , \2218 , \2330 );
xor \U$1349 ( \2332 , \2218 , \2330 );
xor \U$1350 ( \2333 , \2327 , \2329 );
buf \U$1351 ( \2334 , RIc0d8140_24);
buf \U$1352 ( \2335 , RIc0d81b8_25);
and \U$1353 ( \2336 , \2334 , \2335 );
not \U$1354 ( \2337 , \2336 );
and \U$1355 ( \2338 , \2106 , \2337 );
not \U$1356 ( \2339 , \2338 );
and \U$1357 ( \2340 , \998 , \2222 );
and \U$1358 ( \2341 , \984 , \2220 );
nor \U$1359 ( \2342 , \2340 , \2341 );
xnor \U$1360 ( \2343 , \2342 , \2109 );
and \U$1361 ( \2344 , \2339 , \2343 );
and \U$1362 ( \2345 , \1037 , \2028 );
and \U$1363 ( \2346 , \1016 , \2026 );
nor \U$1364 ( \2347 , \2345 , \2346 );
xnor \U$1365 ( \2348 , \2347 , \1892 );
and \U$1366 ( \2349 , \2343 , \2348 );
and \U$1367 ( \2350 , \2339 , \2348 );
or \U$1368 ( \2351 , \2344 , \2349 , \2350 );
and \U$1369 ( \2352 , \1093 , \1828 );
and \U$1370 ( \2353 , \1085 , \1826 );
nor \U$1371 ( \2354 , \2352 , \2353 );
xnor \U$1372 ( \2355 , \2354 , \1750 );
and \U$1373 ( \2356 , \1167 , \1664 );
and \U$1374 ( \2357 , \1162 , \1662 );
nor \U$1375 ( \2358 , \2356 , \2357 );
xnor \U$1376 ( \2359 , \2358 , \1570 );
and \U$1377 ( \2360 , \2355 , \2359 );
and \U$1378 ( \2361 , \1272 , \1494 );
and \U$1379 ( \2362 , \1221 , \1492 );
nor \U$1380 ( \2363 , \2361 , \2362 );
xnor \U$1381 ( \2364 , \2363 , \1422 );
and \U$1382 ( \2365 , \2359 , \2364 );
and \U$1383 ( \2366 , \2355 , \2364 );
or \U$1384 ( \2367 , \2360 , \2365 , \2366 );
and \U$1385 ( \2368 , \2351 , \2367 );
and \U$1386 ( \2369 , \1377 , \1360 );
and \U$1387 ( \2370 , \1349 , \1358 );
nor \U$1388 ( \2371 , \2369 , \2370 );
xnor \U$1389 ( \2372 , \2371 , \1317 );
and \U$1390 ( \2373 , \1531 , \1247 );
and \U$1391 ( \2374 , \1457 , \1245 );
nor \U$1392 ( \2375 , \2373 , \2374 );
xnor \U$1393 ( \2376 , \2375 , \1198 );
and \U$1394 ( \2377 , \2372 , \2376 );
and \U$1395 ( \2378 , \1656 , \1146 );
and \U$1396 ( \2379 , \1593 , \1144 );
nor \U$1397 ( \2380 , \2378 , \2379 );
xnor \U$1398 ( \2381 , \2380 , \1105 );
and \U$1399 ( \2382 , \2376 , \2381 );
and \U$1400 ( \2383 , \2372 , \2381 );
or \U$1401 ( \2384 , \2377 , \2382 , \2383 );
and \U$1402 ( \2385 , \2367 , \2384 );
and \U$1403 ( \2386 , \2351 , \2384 );
or \U$1404 ( \2387 , \2368 , \2385 , \2386 );
xor \U$1405 ( \2388 , \2225 , \2229 );
xor \U$1406 ( \2389 , \2388 , \2234 );
xor \U$1407 ( \2390 , \2241 , \2245 );
xor \U$1408 ( \2391 , \2390 , \2250 );
and \U$1409 ( \2392 , \2389 , \2391 );
xor \U$1410 ( \2393 , \2258 , \2262 );
xor \U$1411 ( \2394 , \2393 , \2267 );
and \U$1412 ( \2395 , \2391 , \2394 );
and \U$1413 ( \2396 , \2389 , \2394 );
or \U$1414 ( \2397 , \2392 , \2395 , \2396 );
and \U$1415 ( \2398 , \2387 , \2397 );
and \U$1416 ( \2399 , \1942 , \1076 );
and \U$1417 ( \2400 , \1854 , \1074 );
nor \U$1418 ( \2401 , \2399 , \2400 );
xnor \U$1419 ( \2402 , \2401 , \1046 );
and \U$1420 ( \2403 , \2052 , \1028 );
and \U$1421 ( \2404 , \2047 , \1026 );
nor \U$1422 ( \2405 , \2403 , \2404 );
xnor \U$1423 ( \2406 , \2405 , \1009 );
and \U$1424 ( \2407 , \2402 , \2406 );
and \U$1425 ( \2408 , \2283 , \991 );
and \U$1426 ( \2409 , \2168 , \989 );
nor \U$1427 ( \2410 , \2408 , \2409 );
xnor \U$1428 ( \2411 , \2410 , \996 );
and \U$1429 ( \2412 , \2406 , \2411 );
and \U$1430 ( \2413 , \2402 , \2411 );
or \U$1431 ( \2414 , \2407 , \2412 , \2413 );
xor \U$1432 ( \2415 , \2277 , \2281 );
xor \U$1433 ( \2416 , \2415 , \2284 );
or \U$1434 ( \2417 , \2414 , \2416 );
and \U$1435 ( \2418 , \2397 , \2417 );
and \U$1436 ( \2419 , \2387 , \2417 );
or \U$1437 ( \2420 , \2398 , \2418 , \2419 );
xor \U$1438 ( \2421 , \2237 , \2253 );
xor \U$1439 ( \2422 , \2421 , \2270 );
xor \U$1440 ( \2423 , \2287 , \2289 );
xor \U$1441 ( \2424 , \2423 , \2292 );
and \U$1442 ( \2425 , \2422 , \2424 );
xor \U$1443 ( \2426 , \2298 , \2300 );
and \U$1444 ( \2427 , \2424 , \2426 );
and \U$1445 ( \2428 , \2422 , \2426 );
or \U$1446 ( \2429 , \2425 , \2427 , \2428 );
and \U$1447 ( \2430 , \2420 , \2429 );
xor \U$1448 ( \2431 , \2306 , \2308 );
xor \U$1449 ( \2432 , \2431 , \2310 );
and \U$1450 ( \2433 , \2429 , \2432 );
and \U$1451 ( \2434 , \2420 , \2432 );
or \U$1452 ( \2435 , \2430 , \2433 , \2434 );
xor \U$1453 ( \2436 , \2158 , \2179 );
xor \U$1454 ( \2437 , \2436 , \2185 );
and \U$1455 ( \2438 , \2435 , \2437 );
xor \U$1456 ( \2439 , \2304 , \2313 );
xor \U$1457 ( \2440 , \2439 , \2316 );
and \U$1458 ( \2441 , \2437 , \2440 );
and \U$1459 ( \2442 , \2435 , \2440 );
or \U$1460 ( \2443 , \2438 , \2441 , \2442 );
xor \U$1461 ( \2444 , \2319 , \2321 );
xor \U$1462 ( \2445 , \2444 , \2324 );
and \U$1463 ( \2446 , \2443 , \2445 );
and \U$1464 ( \2447 , \2333 , \2446 );
xor \U$1465 ( \2448 , \2333 , \2446 );
xor \U$1466 ( \2449 , \2443 , \2445 );
and \U$1467 ( \2450 , \2047 , \1076 );
and \U$1468 ( \2451 , \1942 , \1074 );
nor \U$1469 ( \2452 , \2450 , \2451 );
xnor \U$1470 ( \2453 , \2452 , \1046 );
and \U$1471 ( \2454 , \2168 , \1028 );
and \U$1472 ( \2455 , \2052 , \1026 );
nor \U$1473 ( \2456 , \2454 , \2455 );
xnor \U$1474 ( \2457 , \2456 , \1009 );
and \U$1475 ( \2458 , \2453 , \2457 );
buf \U$1476 ( \2459 , RIc0d9ec8_87);
and \U$1477 ( \2460 , \2459 , \991 );
and \U$1478 ( \2461 , \2283 , \989 );
nor \U$1479 ( \2462 , \2460 , \2461 );
xnor \U$1480 ( \2463 , \2462 , \996 );
and \U$1481 ( \2464 , \2457 , \2463 );
and \U$1482 ( \2465 , \2453 , \2463 );
or \U$1483 ( \2466 , \2458 , \2464 , \2465 );
buf \U$1484 ( \2467 , RIc0d9f40_88);
and \U$1485 ( \2468 , \2467 , \985 );
buf \U$1486 ( \2469 , \2468 );
and \U$1487 ( \2470 , \2466 , \2469 );
and \U$1488 ( \2471 , \2459 , \985 );
and \U$1489 ( \2472 , \2469 , \2471 );
and \U$1490 ( \2473 , \2466 , \2471 );
or \U$1491 ( \2474 , \2470 , \2472 , \2473 );
and \U$1492 ( \2475 , \1162 , \1828 );
and \U$1493 ( \2476 , \1093 , \1826 );
nor \U$1494 ( \2477 , \2475 , \2476 );
xnor \U$1495 ( \2478 , \2477 , \1750 );
and \U$1496 ( \2479 , \1221 , \1664 );
and \U$1497 ( \2480 , \1167 , \1662 );
nor \U$1498 ( \2481 , \2479 , \2480 );
xnor \U$1499 ( \2482 , \2481 , \1570 );
and \U$1500 ( \2483 , \2478 , \2482 );
and \U$1501 ( \2484 , \1349 , \1494 );
and \U$1502 ( \2485 , \1272 , \1492 );
nor \U$1503 ( \2486 , \2484 , \2485 );
xnor \U$1504 ( \2487 , \2486 , \1422 );
and \U$1505 ( \2488 , \2482 , \2487 );
and \U$1506 ( \2489 , \2478 , \2487 );
or \U$1507 ( \2490 , \2483 , \2488 , \2489 );
xor \U$1508 ( \2491 , \2106 , \2334 );
xor \U$1509 ( \2492 , \2334 , \2335 );
not \U$1510 ( \2493 , \2492 );
and \U$1511 ( \2494 , \2491 , \2493 );
and \U$1512 ( \2495 , \984 , \2494 );
not \U$1513 ( \2496 , \2495 );
xnor \U$1514 ( \2497 , \2496 , \2338 );
and \U$1515 ( \2498 , \1016 , \2222 );
and \U$1516 ( \2499 , \998 , \2220 );
nor \U$1517 ( \2500 , \2498 , \2499 );
xnor \U$1518 ( \2501 , \2500 , \2109 );
and \U$1519 ( \2502 , \2497 , \2501 );
and \U$1520 ( \2503 , \1085 , \2028 );
and \U$1521 ( \2504 , \1037 , \2026 );
nor \U$1522 ( \2505 , \2503 , \2504 );
xnor \U$1523 ( \2506 , \2505 , \1892 );
and \U$1524 ( \2507 , \2501 , \2506 );
and \U$1525 ( \2508 , \2497 , \2506 );
or \U$1526 ( \2509 , \2502 , \2507 , \2508 );
and \U$1527 ( \2510 , \2490 , \2509 );
and \U$1528 ( \2511 , \1457 , \1360 );
and \U$1529 ( \2512 , \1377 , \1358 );
nor \U$1530 ( \2513 , \2511 , \2512 );
xnor \U$1531 ( \2514 , \2513 , \1317 );
and \U$1532 ( \2515 , \1593 , \1247 );
and \U$1533 ( \2516 , \1531 , \1245 );
nor \U$1534 ( \2517 , \2515 , \2516 );
xnor \U$1535 ( \2518 , \2517 , \1198 );
and \U$1536 ( \2519 , \2514 , \2518 );
and \U$1537 ( \2520 , \1854 , \1146 );
and \U$1538 ( \2521 , \1656 , \1144 );
nor \U$1539 ( \2522 , \2520 , \2521 );
xnor \U$1540 ( \2523 , \2522 , \1105 );
and \U$1541 ( \2524 , \2518 , \2523 );
and \U$1542 ( \2525 , \2514 , \2523 );
or \U$1543 ( \2526 , \2519 , \2524 , \2525 );
and \U$1544 ( \2527 , \2509 , \2526 );
and \U$1545 ( \2528 , \2490 , \2526 );
or \U$1546 ( \2529 , \2510 , \2527 , \2528 );
and \U$1547 ( \2530 , \2474 , \2529 );
xor \U$1548 ( \2531 , \2355 , \2359 );
xor \U$1549 ( \2532 , \2531 , \2364 );
xor \U$1550 ( \2533 , \2402 , \2406 );
xor \U$1551 ( \2534 , \2533 , \2411 );
and \U$1552 ( \2535 , \2532 , \2534 );
xor \U$1553 ( \2536 , \2372 , \2376 );
xor \U$1554 ( \2537 , \2536 , \2381 );
and \U$1555 ( \2538 , \2534 , \2537 );
and \U$1556 ( \2539 , \2532 , \2537 );
or \U$1557 ( \2540 , \2535 , \2538 , \2539 );
and \U$1558 ( \2541 , \2529 , \2540 );
and \U$1559 ( \2542 , \2474 , \2540 );
or \U$1560 ( \2543 , \2530 , \2541 , \2542 );
xor \U$1561 ( \2544 , \2351 , \2367 );
xor \U$1562 ( \2545 , \2544 , \2384 );
xor \U$1563 ( \2546 , \2389 , \2391 );
xor \U$1564 ( \2547 , \2546 , \2394 );
and \U$1565 ( \2548 , \2545 , \2547 );
xnor \U$1566 ( \2549 , \2414 , \2416 );
and \U$1567 ( \2550 , \2547 , \2549 );
and \U$1568 ( \2551 , \2545 , \2549 );
or \U$1569 ( \2552 , \2548 , \2550 , \2551 );
and \U$1570 ( \2553 , \2543 , \2552 );
xor \U$1571 ( \2554 , \2422 , \2424 );
xor \U$1572 ( \2555 , \2554 , \2426 );
and \U$1573 ( \2556 , \2552 , \2555 );
and \U$1574 ( \2557 , \2543 , \2555 );
or \U$1575 ( \2558 , \2553 , \2556 , \2557 );
xor \U$1576 ( \2559 , \2273 , \2295 );
xor \U$1577 ( \2560 , \2559 , \2301 );
and \U$1578 ( \2561 , \2558 , \2560 );
xor \U$1579 ( \2562 , \2420 , \2429 );
xor \U$1580 ( \2563 , \2562 , \2432 );
and \U$1581 ( \2564 , \2560 , \2563 );
and \U$1582 ( \2565 , \2558 , \2563 );
or \U$1583 ( \2566 , \2561 , \2564 , \2565 );
xor \U$1584 ( \2567 , \2435 , \2437 );
xor \U$1585 ( \2568 , \2567 , \2440 );
and \U$1586 ( \2569 , \2566 , \2568 );
and \U$1587 ( \2570 , \2449 , \2569 );
xor \U$1588 ( \2571 , \2449 , \2569 );
xor \U$1589 ( \2572 , \2566 , \2568 );
and \U$1590 ( \2573 , \1377 , \1494 );
and \U$1591 ( \2574 , \1349 , \1492 );
nor \U$1592 ( \2575 , \2573 , \2574 );
xnor \U$1593 ( \2576 , \2575 , \1422 );
and \U$1594 ( \2577 , \1531 , \1360 );
and \U$1595 ( \2578 , \1457 , \1358 );
nor \U$1596 ( \2579 , \2577 , \2578 );
xnor \U$1597 ( \2580 , \2579 , \1317 );
and \U$1598 ( \2581 , \2576 , \2580 );
and \U$1599 ( \2582 , \1656 , \1247 );
and \U$1600 ( \2583 , \1593 , \1245 );
nor \U$1601 ( \2584 , \2582 , \2583 );
xnor \U$1602 ( \2585 , \2584 , \1198 );
and \U$1603 ( \2586 , \2580 , \2585 );
and \U$1604 ( \2587 , \2576 , \2585 );
or \U$1605 ( \2588 , \2581 , \2586 , \2587 );
and \U$1606 ( \2589 , \1093 , \2028 );
and \U$1607 ( \2590 , \1085 , \2026 );
nor \U$1608 ( \2591 , \2589 , \2590 );
xnor \U$1609 ( \2592 , \2591 , \1892 );
and \U$1610 ( \2593 , \1167 , \1828 );
and \U$1611 ( \2594 , \1162 , \1826 );
nor \U$1612 ( \2595 , \2593 , \2594 );
xnor \U$1613 ( \2596 , \2595 , \1750 );
and \U$1614 ( \2597 , \2592 , \2596 );
and \U$1615 ( \2598 , \1272 , \1664 );
and \U$1616 ( \2599 , \1221 , \1662 );
nor \U$1617 ( \2600 , \2598 , \2599 );
xnor \U$1618 ( \2601 , \2600 , \1570 );
and \U$1619 ( \2602 , \2596 , \2601 );
and \U$1620 ( \2603 , \2592 , \2601 );
or \U$1621 ( \2604 , \2597 , \2602 , \2603 );
and \U$1622 ( \2605 , \2588 , \2604 );
buf \U$1623 ( \2606 , RIc0d8230_26);
buf \U$1624 ( \2607 , RIc0d82a8_27);
and \U$1625 ( \2608 , \2606 , \2607 );
not \U$1626 ( \2609 , \2608 );
and \U$1627 ( \2610 , \2335 , \2609 );
not \U$1628 ( \2611 , \2610 );
and \U$1629 ( \2612 , \998 , \2494 );
and \U$1630 ( \2613 , \984 , \2492 );
nor \U$1631 ( \2614 , \2612 , \2613 );
xnor \U$1632 ( \2615 , \2614 , \2338 );
and \U$1633 ( \2616 , \2611 , \2615 );
and \U$1634 ( \2617 , \1037 , \2222 );
and \U$1635 ( \2618 , \1016 , \2220 );
nor \U$1636 ( \2619 , \2617 , \2618 );
xnor \U$1637 ( \2620 , \2619 , \2109 );
and \U$1638 ( \2621 , \2615 , \2620 );
and \U$1639 ( \2622 , \2611 , \2620 );
or \U$1640 ( \2623 , \2616 , \2621 , \2622 );
and \U$1641 ( \2624 , \2604 , \2623 );
and \U$1642 ( \2625 , \2588 , \2623 );
or \U$1643 ( \2626 , \2605 , \2624 , \2625 );
xor \U$1644 ( \2627 , \2478 , \2482 );
xor \U$1645 ( \2628 , \2627 , \2487 );
xor \U$1646 ( \2629 , \2497 , \2501 );
xor \U$1647 ( \2630 , \2629 , \2506 );
and \U$1648 ( \2631 , \2628 , \2630 );
xor \U$1649 ( \2632 , \2514 , \2518 );
xor \U$1650 ( \2633 , \2632 , \2523 );
and \U$1651 ( \2634 , \2630 , \2633 );
and \U$1652 ( \2635 , \2628 , \2633 );
or \U$1653 ( \2636 , \2631 , \2634 , \2635 );
and \U$1654 ( \2637 , \2626 , \2636 );
and \U$1655 ( \2638 , \1942 , \1146 );
and \U$1656 ( \2639 , \1854 , \1144 );
nor \U$1657 ( \2640 , \2638 , \2639 );
xnor \U$1658 ( \2641 , \2640 , \1105 );
and \U$1659 ( \2642 , \2052 , \1076 );
and \U$1660 ( \2643 , \2047 , \1074 );
nor \U$1661 ( \2644 , \2642 , \2643 );
xnor \U$1662 ( \2645 , \2644 , \1046 );
and \U$1663 ( \2646 , \2641 , \2645 );
and \U$1664 ( \2647 , \2283 , \1028 );
and \U$1665 ( \2648 , \2168 , \1026 );
nor \U$1666 ( \2649 , \2647 , \2648 );
xnor \U$1667 ( \2650 , \2649 , \1009 );
and \U$1668 ( \2651 , \2645 , \2650 );
and \U$1669 ( \2652 , \2641 , \2650 );
or \U$1670 ( \2653 , \2646 , \2651 , \2652 );
xor \U$1671 ( \2654 , \2453 , \2457 );
xor \U$1672 ( \2655 , \2654 , \2463 );
and \U$1673 ( \2656 , \2653 , \2655 );
not \U$1674 ( \2657 , \2468 );
and \U$1675 ( \2658 , \2655 , \2657 );
and \U$1676 ( \2659 , \2653 , \2657 );
or \U$1677 ( \2660 , \2656 , \2658 , \2659 );
and \U$1678 ( \2661 , \2636 , \2660 );
and \U$1679 ( \2662 , \2626 , \2660 );
or \U$1680 ( \2663 , \2637 , \2661 , \2662 );
xor \U$1681 ( \2664 , \2339 , \2343 );
xor \U$1682 ( \2665 , \2664 , \2348 );
xor \U$1683 ( \2666 , \2466 , \2469 );
xor \U$1684 ( \2667 , \2666 , \2471 );
and \U$1685 ( \2668 , \2665 , \2667 );
xor \U$1686 ( \2669 , \2532 , \2534 );
xor \U$1687 ( \2670 , \2669 , \2537 );
and \U$1688 ( \2671 , \2667 , \2670 );
and \U$1689 ( \2672 , \2665 , \2670 );
or \U$1690 ( \2673 , \2668 , \2671 , \2672 );
and \U$1691 ( \2674 , \2663 , \2673 );
xor \U$1692 ( \2675 , \2545 , \2547 );
xor \U$1693 ( \2676 , \2675 , \2549 );
and \U$1694 ( \2677 , \2673 , \2676 );
and \U$1695 ( \2678 , \2663 , \2676 );
or \U$1696 ( \2679 , \2674 , \2677 , \2678 );
xor \U$1697 ( \2680 , \2387 , \2397 );
xor \U$1698 ( \2681 , \2680 , \2417 );
and \U$1699 ( \2682 , \2679 , \2681 );
xor \U$1700 ( \2683 , \2543 , \2552 );
xor \U$1701 ( \2684 , \2683 , \2555 );
and \U$1702 ( \2685 , \2681 , \2684 );
and \U$1703 ( \2686 , \2679 , \2684 );
or \U$1704 ( \2687 , \2682 , \2685 , \2686 );
xor \U$1705 ( \2688 , \2558 , \2560 );
xor \U$1706 ( \2689 , \2688 , \2563 );
and \U$1707 ( \2690 , \2687 , \2689 );
and \U$1708 ( \2691 , \2572 , \2690 );
xor \U$1709 ( \2692 , \2572 , \2690 );
xor \U$1710 ( \2693 , \2687 , \2689 );
and \U$1711 ( \2694 , \2047 , \1146 );
and \U$1712 ( \2695 , \1942 , \1144 );
nor \U$1713 ( \2696 , \2694 , \2695 );
xnor \U$1714 ( \2697 , \2696 , \1105 );
and \U$1715 ( \2698 , \2168 , \1076 );
and \U$1716 ( \2699 , \2052 , \1074 );
nor \U$1717 ( \2700 , \2698 , \2699 );
xnor \U$1718 ( \2701 , \2700 , \1046 );
and \U$1719 ( \2702 , \2697 , \2701 );
and \U$1720 ( \2703 , \2459 , \1028 );
and \U$1721 ( \2704 , \2283 , \1026 );
nor \U$1722 ( \2705 , \2703 , \2704 );
xnor \U$1723 ( \2706 , \2705 , \1009 );
and \U$1724 ( \2707 , \2701 , \2706 );
and \U$1725 ( \2708 , \2697 , \2706 );
or \U$1726 ( \2709 , \2702 , \2707 , \2708 );
buf \U$1727 ( \2710 , RIc0d9fb8_89);
and \U$1728 ( \2711 , \2710 , \991 );
and \U$1729 ( \2712 , \2467 , \989 );
nor \U$1730 ( \2713 , \2711 , \2712 );
xnor \U$1731 ( \2714 , \2713 , \996 );
buf \U$1732 ( \2715 , RIc0da030_90);
and \U$1733 ( \2716 , \2715 , \985 );
or \U$1734 ( \2717 , \2714 , \2716 );
and \U$1735 ( \2718 , \2709 , \2717 );
and \U$1736 ( \2719 , \2467 , \991 );
and \U$1737 ( \2720 , \2459 , \989 );
nor \U$1738 ( \2721 , \2719 , \2720 );
xnor \U$1739 ( \2722 , \2721 , \996 );
and \U$1740 ( \2723 , \2717 , \2722 );
and \U$1741 ( \2724 , \2709 , \2722 );
or \U$1742 ( \2725 , \2718 , \2723 , \2724 );
and \U$1743 ( \2726 , \1457 , \1494 );
and \U$1744 ( \2727 , \1377 , \1492 );
nor \U$1745 ( \2728 , \2726 , \2727 );
xnor \U$1746 ( \2729 , \2728 , \1422 );
and \U$1747 ( \2730 , \1593 , \1360 );
and \U$1748 ( \2731 , \1531 , \1358 );
nor \U$1749 ( \2732 , \2730 , \2731 );
xnor \U$1750 ( \2733 , \2732 , \1317 );
and \U$1751 ( \2734 , \2729 , \2733 );
and \U$1752 ( \2735 , \1854 , \1247 );
and \U$1753 ( \2736 , \1656 , \1245 );
nor \U$1754 ( \2737 , \2735 , \2736 );
xnor \U$1755 ( \2738 , \2737 , \1198 );
and \U$1756 ( \2739 , \2733 , \2738 );
and \U$1757 ( \2740 , \2729 , \2738 );
or \U$1758 ( \2741 , \2734 , \2739 , \2740 );
and \U$1759 ( \2742 , \1162 , \2028 );
and \U$1760 ( \2743 , \1093 , \2026 );
nor \U$1761 ( \2744 , \2742 , \2743 );
xnor \U$1762 ( \2745 , \2744 , \1892 );
and \U$1763 ( \2746 , \1221 , \1828 );
and \U$1764 ( \2747 , \1167 , \1826 );
nor \U$1765 ( \2748 , \2746 , \2747 );
xnor \U$1766 ( \2749 , \2748 , \1750 );
and \U$1767 ( \2750 , \2745 , \2749 );
and \U$1768 ( \2751 , \1349 , \1664 );
and \U$1769 ( \2752 , \1272 , \1662 );
nor \U$1770 ( \2753 , \2751 , \2752 );
xnor \U$1771 ( \2754 , \2753 , \1570 );
and \U$1772 ( \2755 , \2749 , \2754 );
and \U$1773 ( \2756 , \2745 , \2754 );
or \U$1774 ( \2757 , \2750 , \2755 , \2756 );
and \U$1775 ( \2758 , \2741 , \2757 );
xor \U$1776 ( \2759 , \2335 , \2606 );
xor \U$1777 ( \2760 , \2606 , \2607 );
not \U$1778 ( \2761 , \2760 );
and \U$1779 ( \2762 , \2759 , \2761 );
and \U$1780 ( \2763 , \984 , \2762 );
not \U$1781 ( \2764 , \2763 );
xnor \U$1782 ( \2765 , \2764 , \2610 );
and \U$1783 ( \2766 , \1016 , \2494 );
and \U$1784 ( \2767 , \998 , \2492 );
nor \U$1785 ( \2768 , \2766 , \2767 );
xnor \U$1786 ( \2769 , \2768 , \2338 );
and \U$1787 ( \2770 , \2765 , \2769 );
and \U$1788 ( \2771 , \1085 , \2222 );
and \U$1789 ( \2772 , \1037 , \2220 );
nor \U$1790 ( \2773 , \2771 , \2772 );
xnor \U$1791 ( \2774 , \2773 , \2109 );
and \U$1792 ( \2775 , \2769 , \2774 );
and \U$1793 ( \2776 , \2765 , \2774 );
or \U$1794 ( \2777 , \2770 , \2775 , \2776 );
and \U$1795 ( \2778 , \2757 , \2777 );
and \U$1796 ( \2779 , \2741 , \2777 );
or \U$1797 ( \2780 , \2758 , \2778 , \2779 );
and \U$1798 ( \2781 , \2725 , \2780 );
and \U$1799 ( \2782 , \2710 , \985 );
xor \U$1800 ( \2783 , \2576 , \2580 );
xor \U$1801 ( \2784 , \2783 , \2585 );
and \U$1802 ( \2785 , \2782 , \2784 );
xor \U$1803 ( \2786 , \2641 , \2645 );
xor \U$1804 ( \2787 , \2786 , \2650 );
and \U$1805 ( \2788 , \2784 , \2787 );
and \U$1806 ( \2789 , \2782 , \2787 );
or \U$1807 ( \2790 , \2785 , \2788 , \2789 );
and \U$1808 ( \2791 , \2780 , \2790 );
and \U$1809 ( \2792 , \2725 , \2790 );
or \U$1810 ( \2793 , \2781 , \2791 , \2792 );
xor \U$1811 ( \2794 , \2588 , \2604 );
xor \U$1812 ( \2795 , \2794 , \2623 );
xor \U$1813 ( \2796 , \2628 , \2630 );
xor \U$1814 ( \2797 , \2796 , \2633 );
and \U$1815 ( \2798 , \2795 , \2797 );
xor \U$1816 ( \2799 , \2653 , \2655 );
xor \U$1817 ( \2800 , \2799 , \2657 );
and \U$1818 ( \2801 , \2797 , \2800 );
and \U$1819 ( \2802 , \2795 , \2800 );
or \U$1820 ( \2803 , \2798 , \2801 , \2802 );
and \U$1821 ( \2804 , \2793 , \2803 );
xor \U$1822 ( \2805 , \2490 , \2509 );
xor \U$1823 ( \2806 , \2805 , \2526 );
and \U$1824 ( \2807 , \2803 , \2806 );
and \U$1825 ( \2808 , \2793 , \2806 );
or \U$1826 ( \2809 , \2804 , \2807 , \2808 );
xor \U$1827 ( \2810 , \2626 , \2636 );
xor \U$1828 ( \2811 , \2810 , \2660 );
xor \U$1829 ( \2812 , \2665 , \2667 );
xor \U$1830 ( \2813 , \2812 , \2670 );
and \U$1831 ( \2814 , \2811 , \2813 );
and \U$1832 ( \2815 , \2809 , \2814 );
xor \U$1833 ( \2816 , \2474 , \2529 );
xor \U$1834 ( \2817 , \2816 , \2540 );
and \U$1835 ( \2818 , \2814 , \2817 );
and \U$1836 ( \2819 , \2809 , \2817 );
or \U$1837 ( \2820 , \2815 , \2818 , \2819 );
xor \U$1838 ( \2821 , \2679 , \2681 );
xor \U$1839 ( \2822 , \2821 , \2684 );
and \U$1840 ( \2823 , \2820 , \2822 );
and \U$1841 ( \2824 , \2693 , \2823 );
xor \U$1842 ( \2825 , \2693 , \2823 );
xor \U$1843 ( \2826 , \2820 , \2822 );
buf \U$1844 ( \2827 , RIc0d8320_28);
buf \U$1845 ( \2828 , RIc0d8398_29);
and \U$1846 ( \2829 , \2827 , \2828 );
not \U$1847 ( \2830 , \2829 );
and \U$1848 ( \2831 , \2607 , \2830 );
not \U$1849 ( \2832 , \2831 );
and \U$1850 ( \2833 , \998 , \2762 );
and \U$1851 ( \2834 , \984 , \2760 );
nor \U$1852 ( \2835 , \2833 , \2834 );
xnor \U$1853 ( \2836 , \2835 , \2610 );
and \U$1854 ( \2837 , \2832 , \2836 );
and \U$1855 ( \2838 , \1037 , \2494 );
and \U$1856 ( \2839 , \1016 , \2492 );
nor \U$1857 ( \2840 , \2838 , \2839 );
xnor \U$1858 ( \2841 , \2840 , \2338 );
and \U$1859 ( \2842 , \2836 , \2841 );
and \U$1860 ( \2843 , \2832 , \2841 );
or \U$1861 ( \2844 , \2837 , \2842 , \2843 );
and \U$1862 ( \2845 , \1093 , \2222 );
and \U$1863 ( \2846 , \1085 , \2220 );
nor \U$1864 ( \2847 , \2845 , \2846 );
xnor \U$1865 ( \2848 , \2847 , \2109 );
and \U$1866 ( \2849 , \1167 , \2028 );
and \U$1867 ( \2850 , \1162 , \2026 );
nor \U$1868 ( \2851 , \2849 , \2850 );
xnor \U$1869 ( \2852 , \2851 , \1892 );
and \U$1870 ( \2853 , \2848 , \2852 );
and \U$1871 ( \2854 , \1272 , \1828 );
and \U$1872 ( \2855 , \1221 , \1826 );
nor \U$1873 ( \2856 , \2854 , \2855 );
xnor \U$1874 ( \2857 , \2856 , \1750 );
and \U$1875 ( \2858 , \2852 , \2857 );
and \U$1876 ( \2859 , \2848 , \2857 );
or \U$1877 ( \2860 , \2853 , \2858 , \2859 );
and \U$1878 ( \2861 , \2844 , \2860 );
and \U$1879 ( \2862 , \1377 , \1664 );
and \U$1880 ( \2863 , \1349 , \1662 );
nor \U$1881 ( \2864 , \2862 , \2863 );
xnor \U$1882 ( \2865 , \2864 , \1570 );
and \U$1883 ( \2866 , \1531 , \1494 );
and \U$1884 ( \2867 , \1457 , \1492 );
nor \U$1885 ( \2868 , \2866 , \2867 );
xnor \U$1886 ( \2869 , \2868 , \1422 );
and \U$1887 ( \2870 , \2865 , \2869 );
and \U$1888 ( \2871 , \1656 , \1360 );
and \U$1889 ( \2872 , \1593 , \1358 );
nor \U$1890 ( \2873 , \2871 , \2872 );
xnor \U$1891 ( \2874 , \2873 , \1317 );
and \U$1892 ( \2875 , \2869 , \2874 );
and \U$1893 ( \2876 , \2865 , \2874 );
or \U$1894 ( \2877 , \2870 , \2875 , \2876 );
and \U$1895 ( \2878 , \2860 , \2877 );
and \U$1896 ( \2879 , \2844 , \2877 );
or \U$1897 ( \2880 , \2861 , \2878 , \2879 );
xor \U$1898 ( \2881 , \2729 , \2733 );
xor \U$1899 ( \2882 , \2881 , \2738 );
xor \U$1900 ( \2883 , \2745 , \2749 );
xor \U$1901 ( \2884 , \2883 , \2754 );
and \U$1902 ( \2885 , \2882 , \2884 );
xor \U$1903 ( \2886 , \2697 , \2701 );
xor \U$1904 ( \2887 , \2886 , \2706 );
and \U$1905 ( \2888 , \2884 , \2887 );
and \U$1906 ( \2889 , \2882 , \2887 );
or \U$1907 ( \2890 , \2885 , \2888 , \2889 );
and \U$1908 ( \2891 , \2880 , \2890 );
and \U$1909 ( \2892 , \2467 , \1028 );
and \U$1910 ( \2893 , \2459 , \1026 );
nor \U$1911 ( \2894 , \2892 , \2893 );
xnor \U$1912 ( \2895 , \2894 , \1009 );
and \U$1913 ( \2896 , \2715 , \991 );
and \U$1914 ( \2897 , \2710 , \989 );
nor \U$1915 ( \2898 , \2896 , \2897 );
xnor \U$1916 ( \2899 , \2898 , \996 );
and \U$1917 ( \2900 , \2895 , \2899 );
buf \U$1918 ( \2901 , RIc0da0a8_91);
and \U$1919 ( \2902 , \2901 , \985 );
and \U$1920 ( \2903 , \2899 , \2902 );
and \U$1921 ( \2904 , \2895 , \2902 );
or \U$1922 ( \2905 , \2900 , \2903 , \2904 );
and \U$1923 ( \2906 , \1942 , \1247 );
and \U$1924 ( \2907 , \1854 , \1245 );
nor \U$1925 ( \2908 , \2906 , \2907 );
xnor \U$1926 ( \2909 , \2908 , \1198 );
and \U$1927 ( \2910 , \2052 , \1146 );
and \U$1928 ( \2911 , \2047 , \1144 );
nor \U$1929 ( \2912 , \2910 , \2911 );
xnor \U$1930 ( \2913 , \2912 , \1105 );
and \U$1931 ( \2914 , \2909 , \2913 );
and \U$1932 ( \2915 , \2283 , \1076 );
and \U$1933 ( \2916 , \2168 , \1074 );
nor \U$1934 ( \2917 , \2915 , \2916 );
xnor \U$1935 ( \2918 , \2917 , \1046 );
and \U$1936 ( \2919 , \2913 , \2918 );
and \U$1937 ( \2920 , \2909 , \2918 );
or \U$1938 ( \2921 , \2914 , \2919 , \2920 );
and \U$1939 ( \2922 , \2905 , \2921 );
xnor \U$1940 ( \2923 , \2714 , \2716 );
and \U$1941 ( \2924 , \2921 , \2923 );
and \U$1942 ( \2925 , \2905 , \2923 );
or \U$1943 ( \2926 , \2922 , \2924 , \2925 );
and \U$1944 ( \2927 , \2890 , \2926 );
and \U$1945 ( \2928 , \2880 , \2926 );
or \U$1946 ( \2929 , \2891 , \2927 , \2928 );
xor \U$1947 ( \2930 , \2592 , \2596 );
xor \U$1948 ( \2931 , \2930 , \2601 );
xor \U$1949 ( \2932 , \2611 , \2615 );
xor \U$1950 ( \2933 , \2932 , \2620 );
and \U$1951 ( \2934 , \2931 , \2933 );
xor \U$1952 ( \2935 , \2782 , \2784 );
xor \U$1953 ( \2936 , \2935 , \2787 );
and \U$1954 ( \2937 , \2933 , \2936 );
and \U$1955 ( \2938 , \2931 , \2936 );
or \U$1956 ( \2939 , \2934 , \2937 , \2938 );
and \U$1957 ( \2940 , \2929 , \2939 );
xor \U$1958 ( \2941 , \2795 , \2797 );
xor \U$1959 ( \2942 , \2941 , \2800 );
and \U$1960 ( \2943 , \2939 , \2942 );
and \U$1961 ( \2944 , \2929 , \2942 );
or \U$1962 ( \2945 , \2940 , \2943 , \2944 );
xor \U$1963 ( \2946 , \2793 , \2803 );
xor \U$1964 ( \2947 , \2946 , \2806 );
and \U$1965 ( \2948 , \2945 , \2947 );
xor \U$1966 ( \2949 , \2811 , \2813 );
and \U$1967 ( \2950 , \2947 , \2949 );
and \U$1968 ( \2951 , \2945 , \2949 );
or \U$1969 ( \2952 , \2948 , \2950 , \2951 );
xor \U$1970 ( \2953 , \2809 , \2814 );
xor \U$1971 ( \2954 , \2953 , \2817 );
and \U$1972 ( \2955 , \2952 , \2954 );
xor \U$1973 ( \2956 , \2663 , \2673 );
xor \U$1974 ( \2957 , \2956 , \2676 );
and \U$1975 ( \2958 , \2954 , \2957 );
and \U$1976 ( \2959 , \2952 , \2957 );
or \U$1977 ( \2960 , \2955 , \2958 , \2959 );
and \U$1978 ( \2961 , \2826 , \2960 );
xor \U$1979 ( \2962 , \2826 , \2960 );
xor \U$1980 ( \2963 , \2952 , \2954 );
xor \U$1981 ( \2964 , \2963 , \2957 );
xor \U$1982 ( \2965 , \2607 , \2827 );
xor \U$1983 ( \2966 , \2827 , \2828 );
not \U$1984 ( \2967 , \2966 );
and \U$1985 ( \2968 , \2965 , \2967 );
and \U$1986 ( \2969 , \984 , \2968 );
not \U$1987 ( \2970 , \2969 );
xnor \U$1988 ( \2971 , \2970 , \2831 );
and \U$1989 ( \2972 , \1016 , \2762 );
and \U$1990 ( \2973 , \998 , \2760 );
nor \U$1991 ( \2974 , \2972 , \2973 );
xnor \U$1992 ( \2975 , \2974 , \2610 );
and \U$1993 ( \2976 , \2971 , \2975 );
and \U$1994 ( \2977 , \1085 , \2494 );
and \U$1995 ( \2978 , \1037 , \2492 );
nor \U$1996 ( \2979 , \2977 , \2978 );
xnor \U$1997 ( \2980 , \2979 , \2338 );
and \U$1998 ( \2981 , \2975 , \2980 );
and \U$1999 ( \2982 , \2971 , \2980 );
or \U$2000 ( \2983 , \2976 , \2981 , \2982 );
and \U$2001 ( \2984 , \1162 , \2222 );
and \U$2002 ( \2985 , \1093 , \2220 );
nor \U$2003 ( \2986 , \2984 , \2985 );
xnor \U$2004 ( \2987 , \2986 , \2109 );
and \U$2005 ( \2988 , \1221 , \2028 );
and \U$2006 ( \2989 , \1167 , \2026 );
nor \U$2007 ( \2990 , \2988 , \2989 );
xnor \U$2008 ( \2991 , \2990 , \1892 );
and \U$2009 ( \2992 , \2987 , \2991 );
and \U$2010 ( \2993 , \1349 , \1828 );
and \U$2011 ( \2994 , \1272 , \1826 );
nor \U$2012 ( \2995 , \2993 , \2994 );
xnor \U$2013 ( \2996 , \2995 , \1750 );
and \U$2014 ( \2997 , \2991 , \2996 );
and \U$2015 ( \2998 , \2987 , \2996 );
or \U$2016 ( \2999 , \2992 , \2997 , \2998 );
and \U$2017 ( \3000 , \2983 , \2999 );
and \U$2018 ( \3001 , \1457 , \1664 );
and \U$2019 ( \3002 , \1377 , \1662 );
nor \U$2020 ( \3003 , \3001 , \3002 );
xnor \U$2021 ( \3004 , \3003 , \1570 );
and \U$2022 ( \3005 , \1593 , \1494 );
and \U$2023 ( \3006 , \1531 , \1492 );
nor \U$2024 ( \3007 , \3005 , \3006 );
xnor \U$2025 ( \3008 , \3007 , \1422 );
and \U$2026 ( \3009 , \3004 , \3008 );
and \U$2027 ( \3010 , \1854 , \1360 );
and \U$2028 ( \3011 , \1656 , \1358 );
nor \U$2029 ( \3012 , \3010 , \3011 );
xnor \U$2030 ( \3013 , \3012 , \1317 );
and \U$2031 ( \3014 , \3008 , \3013 );
and \U$2032 ( \3015 , \3004 , \3013 );
or \U$2033 ( \3016 , \3009 , \3014 , \3015 );
and \U$2034 ( \3017 , \2999 , \3016 );
and \U$2035 ( \3018 , \2983 , \3016 );
or \U$2036 ( \3019 , \3000 , \3017 , \3018 );
and \U$2037 ( \3020 , \2047 , \1247 );
and \U$2038 ( \3021 , \1942 , \1245 );
nor \U$2039 ( \3022 , \3020 , \3021 );
xnor \U$2040 ( \3023 , \3022 , \1198 );
and \U$2041 ( \3024 , \2168 , \1146 );
and \U$2042 ( \3025 , \2052 , \1144 );
nor \U$2043 ( \3026 , \3024 , \3025 );
xnor \U$2044 ( \3027 , \3026 , \1105 );
and \U$2045 ( \3028 , \3023 , \3027 );
and \U$2046 ( \3029 , \2459 , \1076 );
and \U$2047 ( \3030 , \2283 , \1074 );
nor \U$2048 ( \3031 , \3029 , \3030 );
xnor \U$2049 ( \3032 , \3031 , \1046 );
and \U$2050 ( \3033 , \3027 , \3032 );
and \U$2051 ( \3034 , \3023 , \3032 );
or \U$2052 ( \3035 , \3028 , \3033 , \3034 );
and \U$2053 ( \3036 , \2710 , \1028 );
and \U$2054 ( \3037 , \2467 , \1026 );
nor \U$2055 ( \3038 , \3036 , \3037 );
xnor \U$2056 ( \3039 , \3038 , \1009 );
and \U$2057 ( \3040 , \2901 , \991 );
and \U$2058 ( \3041 , \2715 , \989 );
nor \U$2059 ( \3042 , \3040 , \3041 );
xnor \U$2060 ( \3043 , \3042 , \996 );
and \U$2061 ( \3044 , \3039 , \3043 );
buf \U$2062 ( \3045 , RIc0da120_92);
and \U$2063 ( \3046 , \3045 , \985 );
and \U$2064 ( \3047 , \3043 , \3046 );
and \U$2065 ( \3048 , \3039 , \3046 );
or \U$2066 ( \3049 , \3044 , \3047 , \3048 );
and \U$2067 ( \3050 , \3035 , \3049 );
xor \U$2068 ( \3051 , \2895 , \2899 );
xor \U$2069 ( \3052 , \3051 , \2902 );
and \U$2070 ( \3053 , \3049 , \3052 );
and \U$2071 ( \3054 , \3035 , \3052 );
or \U$2072 ( \3055 , \3050 , \3053 , \3054 );
and \U$2073 ( \3056 , \3019 , \3055 );
xor \U$2074 ( \3057 , \2848 , \2852 );
xor \U$2075 ( \3058 , \3057 , \2857 );
xor \U$2076 ( \3059 , \2909 , \2913 );
xor \U$2077 ( \3060 , \3059 , \2918 );
and \U$2078 ( \3061 , \3058 , \3060 );
xor \U$2079 ( \3062 , \2865 , \2869 );
xor \U$2080 ( \3063 , \3062 , \2874 );
and \U$2081 ( \3064 , \3060 , \3063 );
and \U$2082 ( \3065 , \3058 , \3063 );
or \U$2083 ( \3066 , \3061 , \3064 , \3065 );
and \U$2084 ( \3067 , \3055 , \3066 );
and \U$2085 ( \3068 , \3019 , \3066 );
or \U$2086 ( \3069 , \3056 , \3067 , \3068 );
xor \U$2087 ( \3070 , \2765 , \2769 );
xor \U$2088 ( \3071 , \3070 , \2774 );
xor \U$2089 ( \3072 , \2882 , \2884 );
xor \U$2090 ( \3073 , \3072 , \2887 );
and \U$2091 ( \3074 , \3071 , \3073 );
xor \U$2092 ( \3075 , \2905 , \2921 );
xor \U$2093 ( \3076 , \3075 , \2923 );
and \U$2094 ( \3077 , \3073 , \3076 );
and \U$2095 ( \3078 , \3071 , \3076 );
or \U$2096 ( \3079 , \3074 , \3077 , \3078 );
and \U$2097 ( \3080 , \3069 , \3079 );
xor \U$2098 ( \3081 , \2709 , \2717 );
xor \U$2099 ( \3082 , \3081 , \2722 );
and \U$2100 ( \3083 , \3079 , \3082 );
and \U$2101 ( \3084 , \3069 , \3082 );
or \U$2102 ( \3085 , \3080 , \3083 , \3084 );
xor \U$2103 ( \3086 , \2741 , \2757 );
xor \U$2104 ( \3087 , \3086 , \2777 );
xor \U$2105 ( \3088 , \2880 , \2890 );
xor \U$2106 ( \3089 , \3088 , \2926 );
and \U$2107 ( \3090 , \3087 , \3089 );
xor \U$2108 ( \3091 , \2931 , \2933 );
xor \U$2109 ( \3092 , \3091 , \2936 );
and \U$2110 ( \3093 , \3089 , \3092 );
and \U$2111 ( \3094 , \3087 , \3092 );
or \U$2112 ( \3095 , \3090 , \3093 , \3094 );
and \U$2113 ( \3096 , \3085 , \3095 );
xor \U$2114 ( \3097 , \2725 , \2780 );
xor \U$2115 ( \3098 , \3097 , \2790 );
and \U$2116 ( \3099 , \3095 , \3098 );
and \U$2117 ( \3100 , \3085 , \3098 );
or \U$2118 ( \3101 , \3096 , \3099 , \3100 );
and \U$2119 ( \3102 , \1093 , \2494 );
and \U$2120 ( \3103 , \1085 , \2492 );
nor \U$2121 ( \3104 , \3102 , \3103 );
xnor \U$2122 ( \3105 , \3104 , \2338 );
and \U$2123 ( \3106 , \1167 , \2222 );
and \U$2124 ( \3107 , \1162 , \2220 );
nor \U$2125 ( \3108 , \3106 , \3107 );
xnor \U$2126 ( \3109 , \3108 , \2109 );
and \U$2127 ( \3110 , \3105 , \3109 );
and \U$2128 ( \3111 , \1272 , \2028 );
and \U$2129 ( \3112 , \1221 , \2026 );
nor \U$2130 ( \3113 , \3111 , \3112 );
xnor \U$2131 ( \3114 , \3113 , \1892 );
and \U$2132 ( \3115 , \3109 , \3114 );
and \U$2133 ( \3116 , \3105 , \3114 );
or \U$2134 ( \3117 , \3110 , \3115 , \3116 );
buf \U$2135 ( \3118 , RIc0d8410_30);
buf \U$2136 ( \3119 , RIc0d8488_31);
and \U$2137 ( \3120 , \3118 , \3119 );
not \U$2138 ( \3121 , \3120 );
and \U$2139 ( \3122 , \2828 , \3121 );
not \U$2140 ( \3123 , \3122 );
and \U$2141 ( \3124 , \998 , \2968 );
and \U$2142 ( \3125 , \984 , \2966 );
nor \U$2143 ( \3126 , \3124 , \3125 );
xnor \U$2144 ( \3127 , \3126 , \2831 );
and \U$2145 ( \3128 , \3123 , \3127 );
and \U$2146 ( \3129 , \1037 , \2762 );
and \U$2147 ( \3130 , \1016 , \2760 );
nor \U$2148 ( \3131 , \3129 , \3130 );
xnor \U$2149 ( \3132 , \3131 , \2610 );
and \U$2150 ( \3133 , \3127 , \3132 );
and \U$2151 ( \3134 , \3123 , \3132 );
or \U$2152 ( \3135 , \3128 , \3133 , \3134 );
and \U$2153 ( \3136 , \3117 , \3135 );
and \U$2154 ( \3137 , \1377 , \1828 );
and \U$2155 ( \3138 , \1349 , \1826 );
nor \U$2156 ( \3139 , \3137 , \3138 );
xnor \U$2157 ( \3140 , \3139 , \1750 );
and \U$2158 ( \3141 , \1531 , \1664 );
and \U$2159 ( \3142 , \1457 , \1662 );
nor \U$2160 ( \3143 , \3141 , \3142 );
xnor \U$2161 ( \3144 , \3143 , \1570 );
and \U$2162 ( \3145 , \3140 , \3144 );
and \U$2163 ( \3146 , \1656 , \1494 );
and \U$2164 ( \3147 , \1593 , \1492 );
nor \U$2165 ( \3148 , \3146 , \3147 );
xnor \U$2166 ( \3149 , \3148 , \1422 );
and \U$2167 ( \3150 , \3144 , \3149 );
and \U$2168 ( \3151 , \3140 , \3149 );
or \U$2169 ( \3152 , \3145 , \3150 , \3151 );
and \U$2170 ( \3153 , \3135 , \3152 );
and \U$2171 ( \3154 , \3117 , \3152 );
or \U$2172 ( \3155 , \3136 , \3153 , \3154 );
xor \U$2173 ( \3156 , \3023 , \3027 );
xor \U$2174 ( \3157 , \3156 , \3032 );
xor \U$2175 ( \3158 , \3039 , \3043 );
xor \U$2176 ( \3159 , \3158 , \3046 );
and \U$2177 ( \3160 , \3157 , \3159 );
xor \U$2178 ( \3161 , \3004 , \3008 );
xor \U$2179 ( \3162 , \3161 , \3013 );
and \U$2180 ( \3163 , \3159 , \3162 );
and \U$2181 ( \3164 , \3157 , \3162 );
or \U$2182 ( \3165 , \3160 , \3163 , \3164 );
and \U$2183 ( \3166 , \3155 , \3165 );
and \U$2184 ( \3167 , \2467 , \1076 );
and \U$2185 ( \3168 , \2459 , \1074 );
nor \U$2186 ( \3169 , \3167 , \3168 );
xnor \U$2187 ( \3170 , \3169 , \1046 );
and \U$2188 ( \3171 , \2715 , \1028 );
and \U$2189 ( \3172 , \2710 , \1026 );
nor \U$2190 ( \3173 , \3171 , \3172 );
xnor \U$2191 ( \3174 , \3173 , \1009 );
and \U$2192 ( \3175 , \3170 , \3174 );
and \U$2193 ( \3176 , \3045 , \991 );
and \U$2194 ( \3177 , \2901 , \989 );
nor \U$2195 ( \3178 , \3176 , \3177 );
xnor \U$2196 ( \3179 , \3178 , \996 );
and \U$2197 ( \3180 , \3174 , \3179 );
and \U$2198 ( \3181 , \3170 , \3179 );
or \U$2199 ( \3182 , \3175 , \3180 , \3181 );
and \U$2200 ( \3183 , \1942 , \1360 );
and \U$2201 ( \3184 , \1854 , \1358 );
nor \U$2202 ( \3185 , \3183 , \3184 );
xnor \U$2203 ( \3186 , \3185 , \1317 );
and \U$2204 ( \3187 , \2052 , \1247 );
and \U$2205 ( \3188 , \2047 , \1245 );
nor \U$2206 ( \3189 , \3187 , \3188 );
xnor \U$2207 ( \3190 , \3189 , \1198 );
and \U$2208 ( \3191 , \3186 , \3190 );
and \U$2209 ( \3192 , \2283 , \1146 );
and \U$2210 ( \3193 , \2168 , \1144 );
nor \U$2211 ( \3194 , \3192 , \3193 );
xnor \U$2212 ( \3195 , \3194 , \1105 );
and \U$2213 ( \3196 , \3190 , \3195 );
and \U$2214 ( \3197 , \3186 , \3195 );
or \U$2215 ( \3198 , \3191 , \3196 , \3197 );
or \U$2216 ( \3199 , \3182 , \3198 );
and \U$2217 ( \3200 , \3165 , \3199 );
and \U$2218 ( \3201 , \3155 , \3199 );
or \U$2219 ( \3202 , \3166 , \3200 , \3201 );
xor \U$2220 ( \3203 , \2832 , \2836 );
xor \U$2221 ( \3204 , \3203 , \2841 );
xor \U$2222 ( \3205 , \3035 , \3049 );
xor \U$2223 ( \3206 , \3205 , \3052 );
and \U$2224 ( \3207 , \3204 , \3206 );
xor \U$2225 ( \3208 , \3058 , \3060 );
xor \U$2226 ( \3209 , \3208 , \3063 );
and \U$2227 ( \3210 , \3206 , \3209 );
and \U$2228 ( \3211 , \3204 , \3209 );
or \U$2229 ( \3212 , \3207 , \3210 , \3211 );
and \U$2230 ( \3213 , \3202 , \3212 );
xor \U$2231 ( \3214 , \2844 , \2860 );
xor \U$2232 ( \3215 , \3214 , \2877 );
and \U$2233 ( \3216 , \3212 , \3215 );
and \U$2234 ( \3217 , \3202 , \3215 );
or \U$2235 ( \3218 , \3213 , \3216 , \3217 );
xor \U$2236 ( \3219 , \3069 , \3079 );
xor \U$2237 ( \3220 , \3219 , \3082 );
and \U$2238 ( \3221 , \3218 , \3220 );
xor \U$2239 ( \3222 , \3087 , \3089 );
xor \U$2240 ( \3223 , \3222 , \3092 );
and \U$2241 ( \3224 , \3220 , \3223 );
and \U$2242 ( \3225 , \3218 , \3223 );
or \U$2243 ( \3226 , \3221 , \3224 , \3225 );
xor \U$2244 ( \3227 , \3085 , \3095 );
xor \U$2245 ( \3228 , \3227 , \3098 );
and \U$2246 ( \3229 , \3226 , \3228 );
xor \U$2247 ( \3230 , \2929 , \2939 );
xor \U$2248 ( \3231 , \3230 , \2942 );
and \U$2249 ( \3232 , \3228 , \3231 );
and \U$2250 ( \3233 , \3226 , \3231 );
or \U$2251 ( \3234 , \3229 , \3232 , \3233 );
and \U$2252 ( \3235 , \3101 , \3234 );
xor \U$2253 ( \3236 , \2945 , \2947 );
xor \U$2254 ( \3237 , \3236 , \2949 );
and \U$2255 ( \3238 , \3234 , \3237 );
and \U$2256 ( \3239 , \3101 , \3237 );
or \U$2257 ( \3240 , \3235 , \3238 , \3239 );
and \U$2258 ( \3241 , \2964 , \3240 );
xor \U$2259 ( \3242 , \2964 , \3240 );
xor \U$2260 ( \3243 , \3101 , \3234 );
xor \U$2261 ( \3244 , \3243 , \3237 );
and \U$2262 ( \3245 , \1162 , \2494 );
and \U$2263 ( \3246 , \1093 , \2492 );
nor \U$2264 ( \3247 , \3245 , \3246 );
xnor \U$2265 ( \3248 , \3247 , \2338 );
and \U$2266 ( \3249 , \1221 , \2222 );
and \U$2267 ( \3250 , \1167 , \2220 );
nor \U$2268 ( \3251 , \3249 , \3250 );
xnor \U$2269 ( \3252 , \3251 , \2109 );
and \U$2270 ( \3253 , \3248 , \3252 );
and \U$2271 ( \3254 , \1349 , \2028 );
and \U$2272 ( \3255 , \1272 , \2026 );
nor \U$2273 ( \3256 , \3254 , \3255 );
xnor \U$2274 ( \3257 , \3256 , \1892 );
and \U$2275 ( \3258 , \3252 , \3257 );
and \U$2276 ( \3259 , \3248 , \3257 );
or \U$2277 ( \3260 , \3253 , \3258 , \3259 );
xor \U$2278 ( \3261 , \2828 , \3118 );
xor \U$2279 ( \3262 , \3118 , \3119 );
not \U$2280 ( \3263 , \3262 );
and \U$2281 ( \3264 , \3261 , \3263 );
and \U$2282 ( \3265 , \984 , \3264 );
not \U$2283 ( \3266 , \3265 );
xnor \U$2284 ( \3267 , \3266 , \3122 );
and \U$2285 ( \3268 , \1016 , \2968 );
and \U$2286 ( \3269 , \998 , \2966 );
nor \U$2287 ( \3270 , \3268 , \3269 );
xnor \U$2288 ( \3271 , \3270 , \2831 );
and \U$2289 ( \3272 , \3267 , \3271 );
and \U$2290 ( \3273 , \1085 , \2762 );
and \U$2291 ( \3274 , \1037 , \2760 );
nor \U$2292 ( \3275 , \3273 , \3274 );
xnor \U$2293 ( \3276 , \3275 , \2610 );
and \U$2294 ( \3277 , \3271 , \3276 );
and \U$2295 ( \3278 , \3267 , \3276 );
or \U$2296 ( \3279 , \3272 , \3277 , \3278 );
and \U$2297 ( \3280 , \3260 , \3279 );
and \U$2298 ( \3281 , \1457 , \1828 );
and \U$2299 ( \3282 , \1377 , \1826 );
nor \U$2300 ( \3283 , \3281 , \3282 );
xnor \U$2301 ( \3284 , \3283 , \1750 );
and \U$2302 ( \3285 , \1593 , \1664 );
and \U$2303 ( \3286 , \1531 , \1662 );
nor \U$2304 ( \3287 , \3285 , \3286 );
xnor \U$2305 ( \3288 , \3287 , \1570 );
and \U$2306 ( \3289 , \3284 , \3288 );
and \U$2307 ( \3290 , \1854 , \1494 );
and \U$2308 ( \3291 , \1656 , \1492 );
nor \U$2309 ( \3292 , \3290 , \3291 );
xnor \U$2310 ( \3293 , \3292 , \1422 );
and \U$2311 ( \3294 , \3288 , \3293 );
and \U$2312 ( \3295 , \3284 , \3293 );
or \U$2313 ( \3296 , \3289 , \3294 , \3295 );
and \U$2314 ( \3297 , \3279 , \3296 );
and \U$2315 ( \3298 , \3260 , \3296 );
or \U$2316 ( \3299 , \3280 , \3297 , \3298 );
and \U$2317 ( \3300 , \2710 , \1076 );
and \U$2318 ( \3301 , \2467 , \1074 );
nor \U$2319 ( \3302 , \3300 , \3301 );
xnor \U$2320 ( \3303 , \3302 , \1046 );
and \U$2321 ( \3304 , \2901 , \1028 );
and \U$2322 ( \3305 , \2715 , \1026 );
nor \U$2323 ( \3306 , \3304 , \3305 );
xnor \U$2324 ( \3307 , \3306 , \1009 );
and \U$2325 ( \3308 , \3303 , \3307 );
buf \U$2326 ( \3309 , RIc0da198_93);
and \U$2327 ( \3310 , \3309 , \991 );
and \U$2328 ( \3311 , \3045 , \989 );
nor \U$2329 ( \3312 , \3310 , \3311 );
xnor \U$2330 ( \3313 , \3312 , \996 );
and \U$2331 ( \3314 , \3307 , \3313 );
and \U$2332 ( \3315 , \3303 , \3313 );
or \U$2333 ( \3316 , \3308 , \3314 , \3315 );
and \U$2334 ( \3317 , \2047 , \1360 );
and \U$2335 ( \3318 , \1942 , \1358 );
nor \U$2336 ( \3319 , \3317 , \3318 );
xnor \U$2337 ( \3320 , \3319 , \1317 );
and \U$2338 ( \3321 , \2168 , \1247 );
and \U$2339 ( \3322 , \2052 , \1245 );
nor \U$2340 ( \3323 , \3321 , \3322 );
xnor \U$2341 ( \3324 , \3323 , \1198 );
and \U$2342 ( \3325 , \3320 , \3324 );
and \U$2343 ( \3326 , \2459 , \1146 );
and \U$2344 ( \3327 , \2283 , \1144 );
nor \U$2345 ( \3328 , \3326 , \3327 );
xnor \U$2346 ( \3329 , \3328 , \1105 );
and \U$2347 ( \3330 , \3324 , \3329 );
and \U$2348 ( \3331 , \3320 , \3329 );
or \U$2349 ( \3332 , \3325 , \3330 , \3331 );
and \U$2350 ( \3333 , \3316 , \3332 );
buf \U$2351 ( \3334 , RIc0da210_94);
and \U$2352 ( \3335 , \3334 , \985 );
buf \U$2353 ( \3336 , \3335 );
and \U$2354 ( \3337 , \3332 , \3336 );
and \U$2355 ( \3338 , \3316 , \3336 );
or \U$2356 ( \3339 , \3333 , \3337 , \3338 );
and \U$2357 ( \3340 , \3299 , \3339 );
and \U$2358 ( \3341 , \3309 , \985 );
xor \U$2359 ( \3342 , \3170 , \3174 );
xor \U$2360 ( \3343 , \3342 , \3179 );
and \U$2361 ( \3344 , \3341 , \3343 );
xor \U$2362 ( \3345 , \3186 , \3190 );
xor \U$2363 ( \3346 , \3345 , \3195 );
and \U$2364 ( \3347 , \3343 , \3346 );
and \U$2365 ( \3348 , \3341 , \3346 );
or \U$2366 ( \3349 , \3344 , \3347 , \3348 );
and \U$2367 ( \3350 , \3339 , \3349 );
and \U$2368 ( \3351 , \3299 , \3349 );
or \U$2369 ( \3352 , \3340 , \3350 , \3351 );
xor \U$2370 ( \3353 , \3105 , \3109 );
xor \U$2371 ( \3354 , \3353 , \3114 );
xor \U$2372 ( \3355 , \3123 , \3127 );
xor \U$2373 ( \3356 , \3355 , \3132 );
and \U$2374 ( \3357 , \3354 , \3356 );
xor \U$2375 ( \3358 , \3140 , \3144 );
xor \U$2376 ( \3359 , \3358 , \3149 );
and \U$2377 ( \3360 , \3356 , \3359 );
and \U$2378 ( \3361 , \3354 , \3359 );
or \U$2379 ( \3362 , \3357 , \3360 , \3361 );
xor \U$2380 ( \3363 , \2971 , \2975 );
xor \U$2381 ( \3364 , \3363 , \2980 );
and \U$2382 ( \3365 , \3362 , \3364 );
xor \U$2383 ( \3366 , \2987 , \2991 );
xor \U$2384 ( \3367 , \3366 , \2996 );
and \U$2385 ( \3368 , \3364 , \3367 );
and \U$2386 ( \3369 , \3362 , \3367 );
or \U$2387 ( \3370 , \3365 , \3368 , \3369 );
and \U$2388 ( \3371 , \3352 , \3370 );
xor \U$2389 ( \3372 , \3117 , \3135 );
xor \U$2390 ( \3373 , \3372 , \3152 );
xor \U$2391 ( \3374 , \3157 , \3159 );
xor \U$2392 ( \3375 , \3374 , \3162 );
and \U$2393 ( \3376 , \3373 , \3375 );
xnor \U$2394 ( \3377 , \3182 , \3198 );
and \U$2395 ( \3378 , \3375 , \3377 );
and \U$2396 ( \3379 , \3373 , \3377 );
or \U$2397 ( \3380 , \3376 , \3378 , \3379 );
and \U$2398 ( \3381 , \3370 , \3380 );
and \U$2399 ( \3382 , \3352 , \3380 );
or \U$2400 ( \3383 , \3371 , \3381 , \3382 );
xor \U$2401 ( \3384 , \2983 , \2999 );
xor \U$2402 ( \3385 , \3384 , \3016 );
xor \U$2403 ( \3386 , \3155 , \3165 );
xor \U$2404 ( \3387 , \3386 , \3199 );
and \U$2405 ( \3388 , \3385 , \3387 );
xor \U$2406 ( \3389 , \3204 , \3206 );
xor \U$2407 ( \3390 , \3389 , \3209 );
and \U$2408 ( \3391 , \3387 , \3390 );
and \U$2409 ( \3392 , \3385 , \3390 );
or \U$2410 ( \3393 , \3388 , \3391 , \3392 );
and \U$2411 ( \3394 , \3383 , \3393 );
xor \U$2412 ( \3395 , \3071 , \3073 );
xor \U$2413 ( \3396 , \3395 , \3076 );
and \U$2414 ( \3397 , \3393 , \3396 );
and \U$2415 ( \3398 , \3383 , \3396 );
or \U$2416 ( \3399 , \3394 , \3397 , \3398 );
xor \U$2417 ( \3400 , \3019 , \3055 );
xor \U$2418 ( \3401 , \3400 , \3066 );
xor \U$2419 ( \3402 , \3202 , \3212 );
xor \U$2420 ( \3403 , \3402 , \3215 );
and \U$2421 ( \3404 , \3401 , \3403 );
and \U$2422 ( \3405 , \3399 , \3404 );
xor \U$2423 ( \3406 , \3218 , \3220 );
xor \U$2424 ( \3407 , \3406 , \3223 );
and \U$2425 ( \3408 , \3404 , \3407 );
and \U$2426 ( \3409 , \3399 , \3407 );
or \U$2427 ( \3410 , \3405 , \3408 , \3409 );
xor \U$2428 ( \3411 , \3226 , \3228 );
xor \U$2429 ( \3412 , \3411 , \3231 );
and \U$2430 ( \3413 , \3410 , \3412 );
and \U$2431 ( \3414 , \3244 , \3413 );
xor \U$2432 ( \3415 , \3244 , \3413 );
xor \U$2433 ( \3416 , \3410 , \3412 );
and \U$2434 ( \3417 , \1377 , \2028 );
and \U$2435 ( \3418 , \1349 , \2026 );
nor \U$2436 ( \3419 , \3417 , \3418 );
xnor \U$2437 ( \3420 , \3419 , \1892 );
and \U$2438 ( \3421 , \1531 , \1828 );
and \U$2439 ( \3422 , \1457 , \1826 );
nor \U$2440 ( \3423 , \3421 , \3422 );
xnor \U$2441 ( \3424 , \3423 , \1750 );
and \U$2442 ( \3425 , \3420 , \3424 );
and \U$2443 ( \3426 , \1656 , \1664 );
and \U$2444 ( \3427 , \1593 , \1662 );
nor \U$2445 ( \3428 , \3426 , \3427 );
xnor \U$2446 ( \3429 , \3428 , \1570 );
and \U$2447 ( \3430 , \3424 , \3429 );
and \U$2448 ( \3431 , \3420 , \3429 );
or \U$2449 ( \3432 , \3425 , \3430 , \3431 );
buf \U$2450 ( \3433 , RIc0d8500_32);
buf \U$2451 ( \3434 , RIc0d8578_33);
and \U$2452 ( \3435 , \3433 , \3434 );
not \U$2453 ( \3436 , \3435 );
and \U$2454 ( \3437 , \3119 , \3436 );
not \U$2455 ( \3438 , \3437 );
and \U$2456 ( \3439 , \998 , \3264 );
and \U$2457 ( \3440 , \984 , \3262 );
nor \U$2458 ( \3441 , \3439 , \3440 );
xnor \U$2459 ( \3442 , \3441 , \3122 );
and \U$2460 ( \3443 , \3438 , \3442 );
and \U$2461 ( \3444 , \1037 , \2968 );
and \U$2462 ( \3445 , \1016 , \2966 );
nor \U$2463 ( \3446 , \3444 , \3445 );
xnor \U$2464 ( \3447 , \3446 , \2831 );
and \U$2465 ( \3448 , \3442 , \3447 );
and \U$2466 ( \3449 , \3438 , \3447 );
or \U$2467 ( \3450 , \3443 , \3448 , \3449 );
and \U$2468 ( \3451 , \3432 , \3450 );
and \U$2469 ( \3452 , \1093 , \2762 );
and \U$2470 ( \3453 , \1085 , \2760 );
nor \U$2471 ( \3454 , \3452 , \3453 );
xnor \U$2472 ( \3455 , \3454 , \2610 );
and \U$2473 ( \3456 , \1167 , \2494 );
and \U$2474 ( \3457 , \1162 , \2492 );
nor \U$2475 ( \3458 , \3456 , \3457 );
xnor \U$2476 ( \3459 , \3458 , \2338 );
and \U$2477 ( \3460 , \3455 , \3459 );
and \U$2478 ( \3461 , \1272 , \2222 );
and \U$2479 ( \3462 , \1221 , \2220 );
nor \U$2480 ( \3463 , \3461 , \3462 );
xnor \U$2481 ( \3464 , \3463 , \2109 );
and \U$2482 ( \3465 , \3459 , \3464 );
and \U$2483 ( \3466 , \3455 , \3464 );
or \U$2484 ( \3467 , \3460 , \3465 , \3466 );
and \U$2485 ( \3468 , \3450 , \3467 );
and \U$2486 ( \3469 , \3432 , \3467 );
or \U$2487 ( \3470 , \3451 , \3468 , \3469 );
and \U$2488 ( \3471 , \2467 , \1146 );
and \U$2489 ( \3472 , \2459 , \1144 );
nor \U$2490 ( \3473 , \3471 , \3472 );
xnor \U$2491 ( \3474 , \3473 , \1105 );
and \U$2492 ( \3475 , \2715 , \1076 );
and \U$2493 ( \3476 , \2710 , \1074 );
nor \U$2494 ( \3477 , \3475 , \3476 );
xnor \U$2495 ( \3478 , \3477 , \1046 );
and \U$2496 ( \3479 , \3474 , \3478 );
and \U$2497 ( \3480 , \3045 , \1028 );
and \U$2498 ( \3481 , \2901 , \1026 );
nor \U$2499 ( \3482 , \3480 , \3481 );
xnor \U$2500 ( \3483 , \3482 , \1009 );
and \U$2501 ( \3484 , \3478 , \3483 );
and \U$2502 ( \3485 , \3474 , \3483 );
or \U$2503 ( \3486 , \3479 , \3484 , \3485 );
and \U$2504 ( \3487 , \1942 , \1494 );
and \U$2505 ( \3488 , \1854 , \1492 );
nor \U$2506 ( \3489 , \3487 , \3488 );
xnor \U$2507 ( \3490 , \3489 , \1422 );
and \U$2508 ( \3491 , \2052 , \1360 );
and \U$2509 ( \3492 , \2047 , \1358 );
nor \U$2510 ( \3493 , \3491 , \3492 );
xnor \U$2511 ( \3494 , \3493 , \1317 );
and \U$2512 ( \3495 , \3490 , \3494 );
and \U$2513 ( \3496 , \2283 , \1247 );
and \U$2514 ( \3497 , \2168 , \1245 );
nor \U$2515 ( \3498 , \3496 , \3497 );
xnor \U$2516 ( \3499 , \3498 , \1198 );
and \U$2517 ( \3500 , \3494 , \3499 );
and \U$2518 ( \3501 , \3490 , \3499 );
or \U$2519 ( \3502 , \3495 , \3500 , \3501 );
and \U$2520 ( \3503 , \3486 , \3502 );
and \U$2521 ( \3504 , \3334 , \991 );
and \U$2522 ( \3505 , \3309 , \989 );
nor \U$2523 ( \3506 , \3504 , \3505 );
xnor \U$2524 ( \3507 , \3506 , \996 );
buf \U$2525 ( \3508 , RIc0da288_95);
and \U$2526 ( \3509 , \3508 , \985 );
and \U$2527 ( \3510 , \3507 , \3509 );
and \U$2528 ( \3511 , \3502 , \3510 );
and \U$2529 ( \3512 , \3486 , \3510 );
or \U$2530 ( \3513 , \3503 , \3511 , \3512 );
and \U$2531 ( \3514 , \3470 , \3513 );
xor \U$2532 ( \3515 , \3303 , \3307 );
xor \U$2533 ( \3516 , \3515 , \3313 );
xor \U$2534 ( \3517 , \3320 , \3324 );
xor \U$2535 ( \3518 , \3517 , \3329 );
and \U$2536 ( \3519 , \3516 , \3518 );
not \U$2537 ( \3520 , \3335 );
and \U$2538 ( \3521 , \3518 , \3520 );
and \U$2539 ( \3522 , \3516 , \3520 );
or \U$2540 ( \3523 , \3519 , \3521 , \3522 );
and \U$2541 ( \3524 , \3513 , \3523 );
and \U$2542 ( \3525 , \3470 , \3523 );
or \U$2543 ( \3526 , \3514 , \3524 , \3525 );
xor \U$2544 ( \3527 , \3248 , \3252 );
xor \U$2545 ( \3528 , \3527 , \3257 );
xor \U$2546 ( \3529 , \3267 , \3271 );
xor \U$2547 ( \3530 , \3529 , \3276 );
and \U$2548 ( \3531 , \3528 , \3530 );
xor \U$2549 ( \3532 , \3284 , \3288 );
xor \U$2550 ( \3533 , \3532 , \3293 );
and \U$2551 ( \3534 , \3530 , \3533 );
and \U$2552 ( \3535 , \3528 , \3533 );
or \U$2553 ( \3536 , \3531 , \3534 , \3535 );
xor \U$2554 ( \3537 , \3354 , \3356 );
xor \U$2555 ( \3538 , \3537 , \3359 );
and \U$2556 ( \3539 , \3536 , \3538 );
xor \U$2557 ( \3540 , \3341 , \3343 );
xor \U$2558 ( \3541 , \3540 , \3346 );
and \U$2559 ( \3542 , \3538 , \3541 );
and \U$2560 ( \3543 , \3536 , \3541 );
or \U$2561 ( \3544 , \3539 , \3542 , \3543 );
and \U$2562 ( \3545 , \3526 , \3544 );
xor \U$2563 ( \3546 , \3260 , \3279 );
xor \U$2564 ( \3547 , \3546 , \3296 );
xor \U$2565 ( \3548 , \3316 , \3332 );
xor \U$2566 ( \3549 , \3548 , \3336 );
and \U$2567 ( \3550 , \3547 , \3549 );
and \U$2568 ( \3551 , \3544 , \3550 );
and \U$2569 ( \3552 , \3526 , \3550 );
or \U$2570 ( \3553 , \3545 , \3551 , \3552 );
xor \U$2571 ( \3554 , \3299 , \3339 );
xor \U$2572 ( \3555 , \3554 , \3349 );
xor \U$2573 ( \3556 , \3362 , \3364 );
xor \U$2574 ( \3557 , \3556 , \3367 );
and \U$2575 ( \3558 , \3555 , \3557 );
xor \U$2576 ( \3559 , \3373 , \3375 );
xor \U$2577 ( \3560 , \3559 , \3377 );
and \U$2578 ( \3561 , \3557 , \3560 );
and \U$2579 ( \3562 , \3555 , \3560 );
or \U$2580 ( \3563 , \3558 , \3561 , \3562 );
and \U$2581 ( \3564 , \3553 , \3563 );
xor \U$2582 ( \3565 , \3385 , \3387 );
xor \U$2583 ( \3566 , \3565 , \3390 );
and \U$2584 ( \3567 , \3563 , \3566 );
and \U$2585 ( \3568 , \3553 , \3566 );
or \U$2586 ( \3569 , \3564 , \3567 , \3568 );
xor \U$2587 ( \3570 , \3383 , \3393 );
xor \U$2588 ( \3571 , \3570 , \3396 );
and \U$2589 ( \3572 , \3569 , \3571 );
xor \U$2590 ( \3573 , \3401 , \3403 );
and \U$2591 ( \3574 , \3571 , \3573 );
and \U$2592 ( \3575 , \3569 , \3573 );
or \U$2593 ( \3576 , \3572 , \3574 , \3575 );
xor \U$2594 ( \3577 , \3399 , \3404 );
xor \U$2595 ( \3578 , \3577 , \3407 );
and \U$2596 ( \3579 , \3576 , \3578 );
and \U$2597 ( \3580 , \3416 , \3579 );
xor \U$2598 ( \3581 , \3416 , \3579 );
xor \U$2599 ( \3582 , \3576 , \3578 );
xor \U$2600 ( \3583 , \3119 , \3433 );
xor \U$2601 ( \3584 , \3433 , \3434 );
not \U$2602 ( \3585 , \3584 );
and \U$2603 ( \3586 , \3583 , \3585 );
and \U$2604 ( \3587 , \984 , \3586 );
not \U$2605 ( \3588 , \3587 );
xnor \U$2606 ( \3589 , \3588 , \3437 );
and \U$2607 ( \3590 , \1016 , \3264 );
and \U$2608 ( \3591 , \998 , \3262 );
nor \U$2609 ( \3592 , \3590 , \3591 );
xnor \U$2610 ( \3593 , \3592 , \3122 );
and \U$2611 ( \3594 , \3589 , \3593 );
and \U$2612 ( \3595 , \1085 , \2968 );
and \U$2613 ( \3596 , \1037 , \2966 );
nor \U$2614 ( \3597 , \3595 , \3596 );
xnor \U$2615 ( \3598 , \3597 , \2831 );
and \U$2616 ( \3599 , \3593 , \3598 );
and \U$2617 ( \3600 , \3589 , \3598 );
or \U$2618 ( \3601 , \3594 , \3599 , \3600 );
and \U$2619 ( \3602 , \1457 , \2028 );
and \U$2620 ( \3603 , \1377 , \2026 );
nor \U$2621 ( \3604 , \3602 , \3603 );
xnor \U$2622 ( \3605 , \3604 , \1892 );
and \U$2623 ( \3606 , \1593 , \1828 );
and \U$2624 ( \3607 , \1531 , \1826 );
nor \U$2625 ( \3608 , \3606 , \3607 );
xnor \U$2626 ( \3609 , \3608 , \1750 );
and \U$2627 ( \3610 , \3605 , \3609 );
and \U$2628 ( \3611 , \1854 , \1664 );
and \U$2629 ( \3612 , \1656 , \1662 );
nor \U$2630 ( \3613 , \3611 , \3612 );
xnor \U$2631 ( \3614 , \3613 , \1570 );
and \U$2632 ( \3615 , \3609 , \3614 );
and \U$2633 ( \3616 , \3605 , \3614 );
or \U$2634 ( \3617 , \3610 , \3615 , \3616 );
and \U$2635 ( \3618 , \3601 , \3617 );
and \U$2636 ( \3619 , \1162 , \2762 );
and \U$2637 ( \3620 , \1093 , \2760 );
nor \U$2638 ( \3621 , \3619 , \3620 );
xnor \U$2639 ( \3622 , \3621 , \2610 );
and \U$2640 ( \3623 , \1221 , \2494 );
and \U$2641 ( \3624 , \1167 , \2492 );
nor \U$2642 ( \3625 , \3623 , \3624 );
xnor \U$2643 ( \3626 , \3625 , \2338 );
and \U$2644 ( \3627 , \3622 , \3626 );
and \U$2645 ( \3628 , \1349 , \2222 );
and \U$2646 ( \3629 , \1272 , \2220 );
nor \U$2647 ( \3630 , \3628 , \3629 );
xnor \U$2648 ( \3631 , \3630 , \2109 );
and \U$2649 ( \3632 , \3626 , \3631 );
and \U$2650 ( \3633 , \3622 , \3631 );
or \U$2651 ( \3634 , \3627 , \3632 , \3633 );
and \U$2652 ( \3635 , \3617 , \3634 );
and \U$2653 ( \3636 , \3601 , \3634 );
or \U$2654 ( \3637 , \3618 , \3635 , \3636 );
and \U$2655 ( \3638 , \2710 , \1146 );
and \U$2656 ( \3639 , \2467 , \1144 );
nor \U$2657 ( \3640 , \3638 , \3639 );
xnor \U$2658 ( \3641 , \3640 , \1105 );
and \U$2659 ( \3642 , \2901 , \1076 );
and \U$2660 ( \3643 , \2715 , \1074 );
nor \U$2661 ( \3644 , \3642 , \3643 );
xnor \U$2662 ( \3645 , \3644 , \1046 );
and \U$2663 ( \3646 , \3641 , \3645 );
and \U$2664 ( \3647 , \3309 , \1028 );
and \U$2665 ( \3648 , \3045 , \1026 );
nor \U$2666 ( \3649 , \3647 , \3648 );
xnor \U$2667 ( \3650 , \3649 , \1009 );
and \U$2668 ( \3651 , \3645 , \3650 );
and \U$2669 ( \3652 , \3641 , \3650 );
or \U$2670 ( \3653 , \3646 , \3651 , \3652 );
and \U$2671 ( \3654 , \2047 , \1494 );
and \U$2672 ( \3655 , \1942 , \1492 );
nor \U$2673 ( \3656 , \3654 , \3655 );
xnor \U$2674 ( \3657 , \3656 , \1422 );
and \U$2675 ( \3658 , \2168 , \1360 );
and \U$2676 ( \3659 , \2052 , \1358 );
nor \U$2677 ( \3660 , \3658 , \3659 );
xnor \U$2678 ( \3661 , \3660 , \1317 );
and \U$2679 ( \3662 , \3657 , \3661 );
and \U$2680 ( \3663 , \2459 , \1247 );
and \U$2681 ( \3664 , \2283 , \1245 );
nor \U$2682 ( \3665 , \3663 , \3664 );
xnor \U$2683 ( \3666 , \3665 , \1198 );
and \U$2684 ( \3667 , \3661 , \3666 );
and \U$2685 ( \3668 , \3657 , \3666 );
or \U$2686 ( \3669 , \3662 , \3667 , \3668 );
and \U$2687 ( \3670 , \3653 , \3669 );
and \U$2688 ( \3671 , \3508 , \991 );
and \U$2689 ( \3672 , \3334 , \989 );
nor \U$2690 ( \3673 , \3671 , \3672 );
xnor \U$2691 ( \3674 , \3673 , \996 );
buf \U$2692 ( \3675 , RIc0da300_96);
and \U$2693 ( \3676 , \3675 , \985 );
or \U$2694 ( \3677 , \3674 , \3676 );
and \U$2695 ( \3678 , \3669 , \3677 );
and \U$2696 ( \3679 , \3653 , \3677 );
or \U$2697 ( \3680 , \3670 , \3678 , \3679 );
and \U$2698 ( \3681 , \3637 , \3680 );
xor \U$2699 ( \3682 , \3474 , \3478 );
xor \U$2700 ( \3683 , \3682 , \3483 );
xor \U$2701 ( \3684 , \3490 , \3494 );
xor \U$2702 ( \3685 , \3684 , \3499 );
and \U$2703 ( \3686 , \3683 , \3685 );
xor \U$2704 ( \3687 , \3507 , \3509 );
and \U$2705 ( \3688 , \3685 , \3687 );
and \U$2706 ( \3689 , \3683 , \3687 );
or \U$2707 ( \3690 , \3686 , \3688 , \3689 );
and \U$2708 ( \3691 , \3680 , \3690 );
and \U$2709 ( \3692 , \3637 , \3690 );
or \U$2710 ( \3693 , \3681 , \3691 , \3692 );
xor \U$2711 ( \3694 , \3420 , \3424 );
xor \U$2712 ( \3695 , \3694 , \3429 );
xor \U$2713 ( \3696 , \3438 , \3442 );
xor \U$2714 ( \3697 , \3696 , \3447 );
and \U$2715 ( \3698 , \3695 , \3697 );
xor \U$2716 ( \3699 , \3455 , \3459 );
xor \U$2717 ( \3700 , \3699 , \3464 );
and \U$2718 ( \3701 , \3697 , \3700 );
and \U$2719 ( \3702 , \3695 , \3700 );
or \U$2720 ( \3703 , \3698 , \3701 , \3702 );
xor \U$2721 ( \3704 , \3528 , \3530 );
xor \U$2722 ( \3705 , \3704 , \3533 );
and \U$2723 ( \3706 , \3703 , \3705 );
xor \U$2724 ( \3707 , \3516 , \3518 );
xor \U$2725 ( \3708 , \3707 , \3520 );
and \U$2726 ( \3709 , \3705 , \3708 );
and \U$2727 ( \3710 , \3703 , \3708 );
or \U$2728 ( \3711 , \3706 , \3709 , \3710 );
and \U$2729 ( \3712 , \3693 , \3711 );
xor \U$2730 ( \3713 , \3432 , \3450 );
xor \U$2731 ( \3714 , \3713 , \3467 );
xor \U$2732 ( \3715 , \3486 , \3502 );
xor \U$2733 ( \3716 , \3715 , \3510 );
and \U$2734 ( \3717 , \3714 , \3716 );
and \U$2735 ( \3718 , \3711 , \3717 );
and \U$2736 ( \3719 , \3693 , \3717 );
or \U$2737 ( \3720 , \3712 , \3718 , \3719 );
xor \U$2738 ( \3721 , \3470 , \3513 );
xor \U$2739 ( \3722 , \3721 , \3523 );
xor \U$2740 ( \3723 , \3536 , \3538 );
xor \U$2741 ( \3724 , \3723 , \3541 );
and \U$2742 ( \3725 , \3722 , \3724 );
xor \U$2743 ( \3726 , \3547 , \3549 );
and \U$2744 ( \3727 , \3724 , \3726 );
and \U$2745 ( \3728 , \3722 , \3726 );
or \U$2746 ( \3729 , \3725 , \3727 , \3728 );
and \U$2747 ( \3730 , \3720 , \3729 );
xor \U$2748 ( \3731 , \3555 , \3557 );
xor \U$2749 ( \3732 , \3731 , \3560 );
and \U$2750 ( \3733 , \3729 , \3732 );
and \U$2751 ( \3734 , \3720 , \3732 );
or \U$2752 ( \3735 , \3730 , \3733 , \3734 );
xor \U$2753 ( \3736 , \3352 , \3370 );
xor \U$2754 ( \3737 , \3736 , \3380 );
and \U$2755 ( \3738 , \3735 , \3737 );
xor \U$2756 ( \3739 , \3553 , \3563 );
xor \U$2757 ( \3740 , \3739 , \3566 );
and \U$2758 ( \3741 , \3737 , \3740 );
and \U$2759 ( \3742 , \3735 , \3740 );
or \U$2760 ( \3743 , \3738 , \3741 , \3742 );
xor \U$2761 ( \3744 , \3569 , \3571 );
xor \U$2762 ( \3745 , \3744 , \3573 );
and \U$2763 ( \3746 , \3743 , \3745 );
and \U$2764 ( \3747 , \3582 , \3746 );
xor \U$2765 ( \3748 , \3582 , \3746 );
xor \U$2766 ( \3749 , \3743 , \3745 );
and \U$2767 ( \3750 , \1093 , \2968 );
and \U$2768 ( \3751 , \1085 , \2966 );
nor \U$2769 ( \3752 , \3750 , \3751 );
xnor \U$2770 ( \3753 , \3752 , \2831 );
and \U$2771 ( \3754 , \1167 , \2762 );
and \U$2772 ( \3755 , \1162 , \2760 );
nor \U$2773 ( \3756 , \3754 , \3755 );
xnor \U$2774 ( \3757 , \3756 , \2610 );
and \U$2775 ( \3758 , \3753 , \3757 );
and \U$2776 ( \3759 , \1272 , \2494 );
and \U$2777 ( \3760 , \1221 , \2492 );
nor \U$2778 ( \3761 , \3759 , \3760 );
xnor \U$2779 ( \3762 , \3761 , \2338 );
and \U$2780 ( \3763 , \3757 , \3762 );
and \U$2781 ( \3764 , \3753 , \3762 );
or \U$2782 ( \3765 , \3758 , \3763 , \3764 );
and \U$2783 ( \3766 , \1377 , \2222 );
and \U$2784 ( \3767 , \1349 , \2220 );
nor \U$2785 ( \3768 , \3766 , \3767 );
xnor \U$2786 ( \3769 , \3768 , \2109 );
and \U$2787 ( \3770 , \1531 , \2028 );
and \U$2788 ( \3771 , \1457 , \2026 );
nor \U$2789 ( \3772 , \3770 , \3771 );
xnor \U$2790 ( \3773 , \3772 , \1892 );
and \U$2791 ( \3774 , \3769 , \3773 );
and \U$2792 ( \3775 , \1656 , \1828 );
and \U$2793 ( \3776 , \1593 , \1826 );
nor \U$2794 ( \3777 , \3775 , \3776 );
xnor \U$2795 ( \3778 , \3777 , \1750 );
and \U$2796 ( \3779 , \3773 , \3778 );
and \U$2797 ( \3780 , \3769 , \3778 );
or \U$2798 ( \3781 , \3774 , \3779 , \3780 );
and \U$2799 ( \3782 , \3765 , \3781 );
buf \U$2800 ( \3783 , RIc0d85f0_34);
buf \U$2801 ( \3784 , RIc0d8668_35);
and \U$2802 ( \3785 , \3783 , \3784 );
not \U$2803 ( \3786 , \3785 );
and \U$2804 ( \3787 , \3434 , \3786 );
not \U$2805 ( \3788 , \3787 );
and \U$2806 ( \3789 , \998 , \3586 );
and \U$2807 ( \3790 , \984 , \3584 );
nor \U$2808 ( \3791 , \3789 , \3790 );
xnor \U$2809 ( \3792 , \3791 , \3437 );
and \U$2810 ( \3793 , \3788 , \3792 );
and \U$2811 ( \3794 , \1037 , \3264 );
and \U$2812 ( \3795 , \1016 , \3262 );
nor \U$2813 ( \3796 , \3794 , \3795 );
xnor \U$2814 ( \3797 , \3796 , \3122 );
and \U$2815 ( \3798 , \3792 , \3797 );
and \U$2816 ( \3799 , \3788 , \3797 );
or \U$2817 ( \3800 , \3793 , \3798 , \3799 );
and \U$2818 ( \3801 , \3781 , \3800 );
and \U$2819 ( \3802 , \3765 , \3800 );
or \U$2820 ( \3803 , \3782 , \3801 , \3802 );
and \U$2821 ( \3804 , \3334 , \1028 );
and \U$2822 ( \3805 , \3309 , \1026 );
nor \U$2823 ( \3806 , \3804 , \3805 );
xnor \U$2824 ( \3807 , \3806 , \1009 );
and \U$2825 ( \3808 , \3675 , \991 );
and \U$2826 ( \3809 , \3508 , \989 );
nor \U$2827 ( \3810 , \3808 , \3809 );
xnor \U$2828 ( \3811 , \3810 , \996 );
and \U$2829 ( \3812 , \3807 , \3811 );
buf \U$2830 ( \3813 , RIc0da378_97);
and \U$2831 ( \3814 , \3813 , \985 );
and \U$2832 ( \3815 , \3811 , \3814 );
and \U$2833 ( \3816 , \3807 , \3814 );
or \U$2834 ( \3817 , \3812 , \3815 , \3816 );
and \U$2835 ( \3818 , \2467 , \1247 );
and \U$2836 ( \3819 , \2459 , \1245 );
nor \U$2837 ( \3820 , \3818 , \3819 );
xnor \U$2838 ( \3821 , \3820 , \1198 );
and \U$2839 ( \3822 , \2715 , \1146 );
and \U$2840 ( \3823 , \2710 , \1144 );
nor \U$2841 ( \3824 , \3822 , \3823 );
xnor \U$2842 ( \3825 , \3824 , \1105 );
and \U$2843 ( \3826 , \3821 , \3825 );
and \U$2844 ( \3827 , \3045 , \1076 );
and \U$2845 ( \3828 , \2901 , \1074 );
nor \U$2846 ( \3829 , \3827 , \3828 );
xnor \U$2847 ( \3830 , \3829 , \1046 );
and \U$2848 ( \3831 , \3825 , \3830 );
and \U$2849 ( \3832 , \3821 , \3830 );
or \U$2850 ( \3833 , \3826 , \3831 , \3832 );
and \U$2851 ( \3834 , \3817 , \3833 );
and \U$2852 ( \3835 , \1942 , \1664 );
and \U$2853 ( \3836 , \1854 , \1662 );
nor \U$2854 ( \3837 , \3835 , \3836 );
xnor \U$2855 ( \3838 , \3837 , \1570 );
and \U$2856 ( \3839 , \2052 , \1494 );
and \U$2857 ( \3840 , \2047 , \1492 );
nor \U$2858 ( \3841 , \3839 , \3840 );
xnor \U$2859 ( \3842 , \3841 , \1422 );
and \U$2860 ( \3843 , \3838 , \3842 );
and \U$2861 ( \3844 , \2283 , \1360 );
and \U$2862 ( \3845 , \2168 , \1358 );
nor \U$2863 ( \3846 , \3844 , \3845 );
xnor \U$2864 ( \3847 , \3846 , \1317 );
and \U$2865 ( \3848 , \3842 , \3847 );
and \U$2866 ( \3849 , \3838 , \3847 );
or \U$2867 ( \3850 , \3843 , \3848 , \3849 );
and \U$2868 ( \3851 , \3833 , \3850 );
and \U$2869 ( \3852 , \3817 , \3850 );
or \U$2870 ( \3853 , \3834 , \3851 , \3852 );
and \U$2871 ( \3854 , \3803 , \3853 );
xor \U$2872 ( \3855 , \3641 , \3645 );
xor \U$2873 ( \3856 , \3855 , \3650 );
xor \U$2874 ( \3857 , \3657 , \3661 );
xor \U$2875 ( \3858 , \3857 , \3666 );
and \U$2876 ( \3859 , \3856 , \3858 );
xnor \U$2877 ( \3860 , \3674 , \3676 );
and \U$2878 ( \3861 , \3858 , \3860 );
and \U$2879 ( \3862 , \3856 , \3860 );
or \U$2880 ( \3863 , \3859 , \3861 , \3862 );
and \U$2881 ( \3864 , \3853 , \3863 );
and \U$2882 ( \3865 , \3803 , \3863 );
or \U$2883 ( \3866 , \3854 , \3864 , \3865 );
xor \U$2884 ( \3867 , \3589 , \3593 );
xor \U$2885 ( \3868 , \3867 , \3598 );
xor \U$2886 ( \3869 , \3605 , \3609 );
xor \U$2887 ( \3870 , \3869 , \3614 );
and \U$2888 ( \3871 , \3868 , \3870 );
xor \U$2889 ( \3872 , \3622 , \3626 );
xor \U$2890 ( \3873 , \3872 , \3631 );
and \U$2891 ( \3874 , \3870 , \3873 );
and \U$2892 ( \3875 , \3868 , \3873 );
or \U$2893 ( \3876 , \3871 , \3874 , \3875 );
xor \U$2894 ( \3877 , \3695 , \3697 );
xor \U$2895 ( \3878 , \3877 , \3700 );
and \U$2896 ( \3879 , \3876 , \3878 );
xor \U$2897 ( \3880 , \3683 , \3685 );
xor \U$2898 ( \3881 , \3880 , \3687 );
and \U$2899 ( \3882 , \3878 , \3881 );
and \U$2900 ( \3883 , \3876 , \3881 );
or \U$2901 ( \3884 , \3879 , \3882 , \3883 );
and \U$2902 ( \3885 , \3866 , \3884 );
xor \U$2903 ( \3886 , \3601 , \3617 );
xor \U$2904 ( \3887 , \3886 , \3634 );
xor \U$2905 ( \3888 , \3653 , \3669 );
xor \U$2906 ( \3889 , \3888 , \3677 );
and \U$2907 ( \3890 , \3887 , \3889 );
and \U$2908 ( \3891 , \3884 , \3890 );
and \U$2909 ( \3892 , \3866 , \3890 );
or \U$2910 ( \3893 , \3885 , \3891 , \3892 );
xor \U$2911 ( \3894 , \3637 , \3680 );
xor \U$2912 ( \3895 , \3894 , \3690 );
xor \U$2913 ( \3896 , \3703 , \3705 );
xor \U$2914 ( \3897 , \3896 , \3708 );
and \U$2915 ( \3898 , \3895 , \3897 );
xor \U$2916 ( \3899 , \3714 , \3716 );
and \U$2917 ( \3900 , \3897 , \3899 );
and \U$2918 ( \3901 , \3895 , \3899 );
or \U$2919 ( \3902 , \3898 , \3900 , \3901 );
and \U$2920 ( \3903 , \3893 , \3902 );
xor \U$2921 ( \3904 , \3722 , \3724 );
xor \U$2922 ( \3905 , \3904 , \3726 );
and \U$2923 ( \3906 , \3902 , \3905 );
and \U$2924 ( \3907 , \3893 , \3905 );
or \U$2925 ( \3908 , \3903 , \3906 , \3907 );
xor \U$2926 ( \3909 , \3526 , \3544 );
xor \U$2927 ( \3910 , \3909 , \3550 );
and \U$2928 ( \3911 , \3908 , \3910 );
xor \U$2929 ( \3912 , \3720 , \3729 );
xor \U$2930 ( \3913 , \3912 , \3732 );
and \U$2931 ( \3914 , \3910 , \3913 );
and \U$2932 ( \3915 , \3908 , \3913 );
or \U$2933 ( \3916 , \3911 , \3914 , \3915 );
xor \U$2934 ( \3917 , \3735 , \3737 );
xor \U$2935 ( \3918 , \3917 , \3740 );
and \U$2936 ( \3919 , \3916 , \3918 );
and \U$2937 ( \3920 , \3749 , \3919 );
xor \U$2938 ( \3921 , \3749 , \3919 );
xor \U$2939 ( \3922 , \3916 , \3918 );
and \U$2940 ( \3923 , \3508 , \1028 );
and \U$2941 ( \3924 , \3334 , \1026 );
nor \U$2942 ( \3925 , \3923 , \3924 );
xnor \U$2943 ( \3926 , \3925 , \1009 );
and \U$2944 ( \3927 , \3813 , \991 );
and \U$2945 ( \3928 , \3675 , \989 );
nor \U$2946 ( \3929 , \3927 , \3928 );
xnor \U$2947 ( \3930 , \3929 , \996 );
and \U$2948 ( \3931 , \3926 , \3930 );
buf \U$2949 ( \3932 , RIc0da3f0_98);
and \U$2950 ( \3933 , \3932 , \985 );
and \U$2951 ( \3934 , \3930 , \3933 );
and \U$2952 ( \3935 , \3926 , \3933 );
or \U$2953 ( \3936 , \3931 , \3934 , \3935 );
and \U$2954 ( \3937 , \2710 , \1247 );
and \U$2955 ( \3938 , \2467 , \1245 );
nor \U$2956 ( \3939 , \3937 , \3938 );
xnor \U$2957 ( \3940 , \3939 , \1198 );
and \U$2958 ( \3941 , \2901 , \1146 );
and \U$2959 ( \3942 , \2715 , \1144 );
nor \U$2960 ( \3943 , \3941 , \3942 );
xnor \U$2961 ( \3944 , \3943 , \1105 );
and \U$2962 ( \3945 , \3940 , \3944 );
and \U$2963 ( \3946 , \3309 , \1076 );
and \U$2964 ( \3947 , \3045 , \1074 );
nor \U$2965 ( \3948 , \3946 , \3947 );
xnor \U$2966 ( \3949 , \3948 , \1046 );
and \U$2967 ( \3950 , \3944 , \3949 );
and \U$2968 ( \3951 , \3940 , \3949 );
or \U$2969 ( \3952 , \3945 , \3950 , \3951 );
and \U$2970 ( \3953 , \3936 , \3952 );
and \U$2971 ( \3954 , \2047 , \1664 );
and \U$2972 ( \3955 , \1942 , \1662 );
nor \U$2973 ( \3956 , \3954 , \3955 );
xnor \U$2974 ( \3957 , \3956 , \1570 );
and \U$2975 ( \3958 , \2168 , \1494 );
and \U$2976 ( \3959 , \2052 , \1492 );
nor \U$2977 ( \3960 , \3958 , \3959 );
xnor \U$2978 ( \3961 , \3960 , \1422 );
and \U$2979 ( \3962 , \3957 , \3961 );
and \U$2980 ( \3963 , \2459 , \1360 );
and \U$2981 ( \3964 , \2283 , \1358 );
nor \U$2982 ( \3965 , \3963 , \3964 );
xnor \U$2983 ( \3966 , \3965 , \1317 );
and \U$2984 ( \3967 , \3961 , \3966 );
and \U$2985 ( \3968 , \3957 , \3966 );
or \U$2986 ( \3969 , \3962 , \3967 , \3968 );
and \U$2987 ( \3970 , \3952 , \3969 );
and \U$2988 ( \3971 , \3936 , \3969 );
or \U$2989 ( \3972 , \3953 , \3970 , \3971 );
and \U$2990 ( \3973 , \1162 , \2968 );
and \U$2991 ( \3974 , \1093 , \2966 );
nor \U$2992 ( \3975 , \3973 , \3974 );
xnor \U$2993 ( \3976 , \3975 , \2831 );
and \U$2994 ( \3977 , \1221 , \2762 );
and \U$2995 ( \3978 , \1167 , \2760 );
nor \U$2996 ( \3979 , \3977 , \3978 );
xnor \U$2997 ( \3980 , \3979 , \2610 );
and \U$2998 ( \3981 , \3976 , \3980 );
and \U$2999 ( \3982 , \1349 , \2494 );
and \U$3000 ( \3983 , \1272 , \2492 );
nor \U$3001 ( \3984 , \3982 , \3983 );
xnor \U$3002 ( \3985 , \3984 , \2338 );
and \U$3003 ( \3986 , \3980 , \3985 );
and \U$3004 ( \3987 , \3976 , \3985 );
or \U$3005 ( \3988 , \3981 , \3986 , \3987 );
xor \U$3006 ( \3989 , \3434 , \3783 );
xor \U$3007 ( \3990 , \3783 , \3784 );
not \U$3008 ( \3991 , \3990 );
and \U$3009 ( \3992 , \3989 , \3991 );
and \U$3010 ( \3993 , \984 , \3992 );
not \U$3011 ( \3994 , \3993 );
xnor \U$3012 ( \3995 , \3994 , \3787 );
and \U$3013 ( \3996 , \1016 , \3586 );
and \U$3014 ( \3997 , \998 , \3584 );
nor \U$3015 ( \3998 , \3996 , \3997 );
xnor \U$3016 ( \3999 , \3998 , \3437 );
and \U$3017 ( \4000 , \3995 , \3999 );
and \U$3018 ( \4001 , \1085 , \3264 );
and \U$3019 ( \4002 , \1037 , \3262 );
nor \U$3020 ( \4003 , \4001 , \4002 );
xnor \U$3021 ( \4004 , \4003 , \3122 );
and \U$3022 ( \4005 , \3999 , \4004 );
and \U$3023 ( \4006 , \3995 , \4004 );
or \U$3024 ( \4007 , \4000 , \4005 , \4006 );
and \U$3025 ( \4008 , \3988 , \4007 );
and \U$3026 ( \4009 , \1457 , \2222 );
and \U$3027 ( \4010 , \1377 , \2220 );
nor \U$3028 ( \4011 , \4009 , \4010 );
xnor \U$3029 ( \4012 , \4011 , \2109 );
and \U$3030 ( \4013 , \1593 , \2028 );
and \U$3031 ( \4014 , \1531 , \2026 );
nor \U$3032 ( \4015 , \4013 , \4014 );
xnor \U$3033 ( \4016 , \4015 , \1892 );
and \U$3034 ( \4017 , \4012 , \4016 );
and \U$3035 ( \4018 , \1854 , \1828 );
and \U$3036 ( \4019 , \1656 , \1826 );
nor \U$3037 ( \4020 , \4018 , \4019 );
xnor \U$3038 ( \4021 , \4020 , \1750 );
and \U$3039 ( \4022 , \4016 , \4021 );
and \U$3040 ( \4023 , \4012 , \4021 );
or \U$3041 ( \4024 , \4017 , \4022 , \4023 );
and \U$3042 ( \4025 , \4007 , \4024 );
and \U$3043 ( \4026 , \3988 , \4024 );
or \U$3044 ( \4027 , \4008 , \4025 , \4026 );
and \U$3045 ( \4028 , \3972 , \4027 );
xor \U$3046 ( \4029 , \3807 , \3811 );
xor \U$3047 ( \4030 , \4029 , \3814 );
xor \U$3048 ( \4031 , \3821 , \3825 );
xor \U$3049 ( \4032 , \4031 , \3830 );
and \U$3050 ( \4033 , \4030 , \4032 );
xor \U$3051 ( \4034 , \3838 , \3842 );
xor \U$3052 ( \4035 , \4034 , \3847 );
and \U$3053 ( \4036 , \4032 , \4035 );
and \U$3054 ( \4037 , \4030 , \4035 );
or \U$3055 ( \4038 , \4033 , \4036 , \4037 );
and \U$3056 ( \4039 , \4027 , \4038 );
and \U$3057 ( \4040 , \3972 , \4038 );
or \U$3058 ( \4041 , \4028 , \4039 , \4040 );
xor \U$3059 ( \4042 , \3753 , \3757 );
xor \U$3060 ( \4043 , \4042 , \3762 );
xor \U$3061 ( \4044 , \3769 , \3773 );
xor \U$3062 ( \4045 , \4044 , \3778 );
and \U$3063 ( \4046 , \4043 , \4045 );
xor \U$3064 ( \4047 , \3788 , \3792 );
xor \U$3065 ( \4048 , \4047 , \3797 );
and \U$3066 ( \4049 , \4045 , \4048 );
and \U$3067 ( \4050 , \4043 , \4048 );
or \U$3068 ( \4051 , \4046 , \4049 , \4050 );
xor \U$3069 ( \4052 , \3868 , \3870 );
xor \U$3070 ( \4053 , \4052 , \3873 );
and \U$3071 ( \4054 , \4051 , \4053 );
xor \U$3072 ( \4055 , \3856 , \3858 );
xor \U$3073 ( \4056 , \4055 , \3860 );
and \U$3074 ( \4057 , \4053 , \4056 );
and \U$3075 ( \4058 , \4051 , \4056 );
or \U$3076 ( \4059 , \4054 , \4057 , \4058 );
and \U$3077 ( \4060 , \4041 , \4059 );
xor \U$3078 ( \4061 , \3765 , \3781 );
xor \U$3079 ( \4062 , \4061 , \3800 );
xor \U$3080 ( \4063 , \3817 , \3833 );
xor \U$3081 ( \4064 , \4063 , \3850 );
and \U$3082 ( \4065 , \4062 , \4064 );
and \U$3083 ( \4066 , \4059 , \4065 );
and \U$3084 ( \4067 , \4041 , \4065 );
or \U$3085 ( \4068 , \4060 , \4066 , \4067 );
xor \U$3086 ( \4069 , \3803 , \3853 );
xor \U$3087 ( \4070 , \4069 , \3863 );
xor \U$3088 ( \4071 , \3876 , \3878 );
xor \U$3089 ( \4072 , \4071 , \3881 );
and \U$3090 ( \4073 , \4070 , \4072 );
xor \U$3091 ( \4074 , \3887 , \3889 );
and \U$3092 ( \4075 , \4072 , \4074 );
and \U$3093 ( \4076 , \4070 , \4074 );
or \U$3094 ( \4077 , \4073 , \4075 , \4076 );
and \U$3095 ( \4078 , \4068 , \4077 );
xor \U$3096 ( \4079 , \3895 , \3897 );
xor \U$3097 ( \4080 , \4079 , \3899 );
and \U$3098 ( \4081 , \4077 , \4080 );
and \U$3099 ( \4082 , \4068 , \4080 );
or \U$3100 ( \4083 , \4078 , \4081 , \4082 );
xor \U$3101 ( \4084 , \3693 , \3711 );
xor \U$3102 ( \4085 , \4084 , \3717 );
and \U$3103 ( \4086 , \4083 , \4085 );
xor \U$3104 ( \4087 , \3893 , \3902 );
xor \U$3105 ( \4088 , \4087 , \3905 );
and \U$3106 ( \4089 , \4085 , \4088 );
and \U$3107 ( \4090 , \4083 , \4088 );
or \U$3108 ( \4091 , \4086 , \4089 , \4090 );
xor \U$3109 ( \4092 , \3908 , \3910 );
xor \U$3110 ( \4093 , \4092 , \3913 );
and \U$3111 ( \4094 , \4091 , \4093 );
and \U$3112 ( \4095 , \3922 , \4094 );
xor \U$3113 ( \4096 , \3922 , \4094 );
xor \U$3114 ( \4097 , \4091 , \4093 );
and \U$3115 ( \4098 , \1377 , \2494 );
and \U$3116 ( \4099 , \1349 , \2492 );
nor \U$3117 ( \4100 , \4098 , \4099 );
xnor \U$3118 ( \4101 , \4100 , \2338 );
and \U$3119 ( \4102 , \1531 , \2222 );
and \U$3120 ( \4103 , \1457 , \2220 );
nor \U$3121 ( \4104 , \4102 , \4103 );
xnor \U$3122 ( \4105 , \4104 , \2109 );
and \U$3123 ( \4106 , \4101 , \4105 );
and \U$3124 ( \4107 , \1656 , \2028 );
and \U$3125 ( \4108 , \1593 , \2026 );
nor \U$3126 ( \4109 , \4107 , \4108 );
xnor \U$3127 ( \4110 , \4109 , \1892 );
and \U$3128 ( \4111 , \4105 , \4110 );
and \U$3129 ( \4112 , \4101 , \4110 );
or \U$3130 ( \4113 , \4106 , \4111 , \4112 );
buf \U$3131 ( \4114 , RIc0d86e0_36);
buf \U$3132 ( \4115 , RIc0d8758_37);
and \U$3133 ( \4116 , \4114 , \4115 );
not \U$3134 ( \4117 , \4116 );
and \U$3135 ( \4118 , \3784 , \4117 );
not \U$3136 ( \4119 , \4118 );
and \U$3137 ( \4120 , \998 , \3992 );
and \U$3138 ( \4121 , \984 , \3990 );
nor \U$3139 ( \4122 , \4120 , \4121 );
xnor \U$3140 ( \4123 , \4122 , \3787 );
and \U$3141 ( \4124 , \4119 , \4123 );
and \U$3142 ( \4125 , \1037 , \3586 );
and \U$3143 ( \4126 , \1016 , \3584 );
nor \U$3144 ( \4127 , \4125 , \4126 );
xnor \U$3145 ( \4128 , \4127 , \3437 );
and \U$3146 ( \4129 , \4123 , \4128 );
and \U$3147 ( \4130 , \4119 , \4128 );
or \U$3148 ( \4131 , \4124 , \4129 , \4130 );
and \U$3149 ( \4132 , \4113 , \4131 );
and \U$3150 ( \4133 , \1093 , \3264 );
and \U$3151 ( \4134 , \1085 , \3262 );
nor \U$3152 ( \4135 , \4133 , \4134 );
xnor \U$3153 ( \4136 , \4135 , \3122 );
and \U$3154 ( \4137 , \1167 , \2968 );
and \U$3155 ( \4138 , \1162 , \2966 );
nor \U$3156 ( \4139 , \4137 , \4138 );
xnor \U$3157 ( \4140 , \4139 , \2831 );
and \U$3158 ( \4141 , \4136 , \4140 );
and \U$3159 ( \4142 , \1272 , \2762 );
and \U$3160 ( \4143 , \1221 , \2760 );
nor \U$3161 ( \4144 , \4142 , \4143 );
xnor \U$3162 ( \4145 , \4144 , \2610 );
and \U$3163 ( \4146 , \4140 , \4145 );
and \U$3164 ( \4147 , \4136 , \4145 );
or \U$3165 ( \4148 , \4141 , \4146 , \4147 );
and \U$3166 ( \4149 , \4131 , \4148 );
and \U$3167 ( \4150 , \4113 , \4148 );
or \U$3168 ( \4151 , \4132 , \4149 , \4150 );
and \U$3169 ( \4152 , \3334 , \1076 );
and \U$3170 ( \4153 , \3309 , \1074 );
nor \U$3171 ( \4154 , \4152 , \4153 );
xnor \U$3172 ( \4155 , \4154 , \1046 );
and \U$3173 ( \4156 , \3675 , \1028 );
and \U$3174 ( \4157 , \3508 , \1026 );
nor \U$3175 ( \4158 , \4156 , \4157 );
xnor \U$3176 ( \4159 , \4158 , \1009 );
and \U$3177 ( \4160 , \4155 , \4159 );
and \U$3178 ( \4161 , \3932 , \991 );
and \U$3179 ( \4162 , \3813 , \989 );
nor \U$3180 ( \4163 , \4161 , \4162 );
xnor \U$3181 ( \4164 , \4163 , \996 );
and \U$3182 ( \4165 , \4159 , \4164 );
and \U$3183 ( \4166 , \4155 , \4164 );
or \U$3184 ( \4167 , \4160 , \4165 , \4166 );
and \U$3185 ( \4168 , \1942 , \1828 );
and \U$3186 ( \4169 , \1854 , \1826 );
nor \U$3187 ( \4170 , \4168 , \4169 );
xnor \U$3188 ( \4171 , \4170 , \1750 );
and \U$3189 ( \4172 , \2052 , \1664 );
and \U$3190 ( \4173 , \2047 , \1662 );
nor \U$3191 ( \4174 , \4172 , \4173 );
xnor \U$3192 ( \4175 , \4174 , \1570 );
and \U$3193 ( \4176 , \4171 , \4175 );
and \U$3194 ( \4177 , \2283 , \1494 );
and \U$3195 ( \4178 , \2168 , \1492 );
nor \U$3196 ( \4179 , \4177 , \4178 );
xnor \U$3197 ( \4180 , \4179 , \1422 );
and \U$3198 ( \4181 , \4175 , \4180 );
and \U$3199 ( \4182 , \4171 , \4180 );
or \U$3200 ( \4183 , \4176 , \4181 , \4182 );
and \U$3201 ( \4184 , \4167 , \4183 );
and \U$3202 ( \4185 , \2467 , \1360 );
and \U$3203 ( \4186 , \2459 , \1358 );
nor \U$3204 ( \4187 , \4185 , \4186 );
xnor \U$3205 ( \4188 , \4187 , \1317 );
and \U$3206 ( \4189 , \2715 , \1247 );
and \U$3207 ( \4190 , \2710 , \1245 );
nor \U$3208 ( \4191 , \4189 , \4190 );
xnor \U$3209 ( \4192 , \4191 , \1198 );
and \U$3210 ( \4193 , \4188 , \4192 );
and \U$3211 ( \4194 , \3045 , \1146 );
and \U$3212 ( \4195 , \2901 , \1144 );
nor \U$3213 ( \4196 , \4194 , \4195 );
xnor \U$3214 ( \4197 , \4196 , \1105 );
and \U$3215 ( \4198 , \4192 , \4197 );
and \U$3216 ( \4199 , \4188 , \4197 );
or \U$3217 ( \4200 , \4193 , \4198 , \4199 );
and \U$3218 ( \4201 , \4183 , \4200 );
and \U$3219 ( \4202 , \4167 , \4200 );
or \U$3220 ( \4203 , \4184 , \4201 , \4202 );
and \U$3221 ( \4204 , \4151 , \4203 );
xor \U$3222 ( \4205 , \3926 , \3930 );
xor \U$3223 ( \4206 , \4205 , \3933 );
xor \U$3224 ( \4207 , \3940 , \3944 );
xor \U$3225 ( \4208 , \4207 , \3949 );
or \U$3226 ( \4209 , \4206 , \4208 );
and \U$3227 ( \4210 , \4203 , \4209 );
and \U$3228 ( \4211 , \4151 , \4209 );
or \U$3229 ( \4212 , \4204 , \4210 , \4211 );
xor \U$3230 ( \4213 , \3976 , \3980 );
xor \U$3231 ( \4214 , \4213 , \3985 );
xor \U$3232 ( \4215 , \4012 , \4016 );
xor \U$3233 ( \4216 , \4215 , \4021 );
and \U$3234 ( \4217 , \4214 , \4216 );
xor \U$3235 ( \4218 , \3957 , \3961 );
xor \U$3236 ( \4219 , \4218 , \3966 );
and \U$3237 ( \4220 , \4216 , \4219 );
and \U$3238 ( \4221 , \4214 , \4219 );
or \U$3239 ( \4222 , \4217 , \4220 , \4221 );
xor \U$3240 ( \4223 , \4030 , \4032 );
xor \U$3241 ( \4224 , \4223 , \4035 );
and \U$3242 ( \4225 , \4222 , \4224 );
xor \U$3243 ( \4226 , \4043 , \4045 );
xor \U$3244 ( \4227 , \4226 , \4048 );
and \U$3245 ( \4228 , \4224 , \4227 );
and \U$3246 ( \4229 , \4222 , \4227 );
or \U$3247 ( \4230 , \4225 , \4228 , \4229 );
and \U$3248 ( \4231 , \4212 , \4230 );
xor \U$3249 ( \4232 , \3936 , \3952 );
xor \U$3250 ( \4233 , \4232 , \3969 );
xor \U$3251 ( \4234 , \3988 , \4007 );
xor \U$3252 ( \4235 , \4234 , \4024 );
and \U$3253 ( \4236 , \4233 , \4235 );
and \U$3254 ( \4237 , \4230 , \4236 );
and \U$3255 ( \4238 , \4212 , \4236 );
or \U$3256 ( \4239 , \4231 , \4237 , \4238 );
xor \U$3257 ( \4240 , \3972 , \4027 );
xor \U$3258 ( \4241 , \4240 , \4038 );
xor \U$3259 ( \4242 , \4051 , \4053 );
xor \U$3260 ( \4243 , \4242 , \4056 );
and \U$3261 ( \4244 , \4241 , \4243 );
xor \U$3262 ( \4245 , \4062 , \4064 );
and \U$3263 ( \4246 , \4243 , \4245 );
and \U$3264 ( \4247 , \4241 , \4245 );
or \U$3265 ( \4248 , \4244 , \4246 , \4247 );
and \U$3266 ( \4249 , \4239 , \4248 );
xor \U$3267 ( \4250 , \4070 , \4072 );
xor \U$3268 ( \4251 , \4250 , \4074 );
and \U$3269 ( \4252 , \4248 , \4251 );
and \U$3270 ( \4253 , \4239 , \4251 );
or \U$3271 ( \4254 , \4249 , \4252 , \4253 );
xor \U$3272 ( \4255 , \3866 , \3884 );
xor \U$3273 ( \4256 , \4255 , \3890 );
and \U$3274 ( \4257 , \4254 , \4256 );
xor \U$3275 ( \4258 , \4068 , \4077 );
xor \U$3276 ( \4259 , \4258 , \4080 );
and \U$3277 ( \4260 , \4256 , \4259 );
and \U$3278 ( \4261 , \4254 , \4259 );
or \U$3279 ( \4262 , \4257 , \4260 , \4261 );
xor \U$3280 ( \4263 , \4083 , \4085 );
xor \U$3281 ( \4264 , \4263 , \4088 );
and \U$3282 ( \4265 , \4262 , \4264 );
and \U$3283 ( \4266 , \4097 , \4265 );
xor \U$3284 ( \4267 , \4097 , \4265 );
xor \U$3285 ( \4268 , \4262 , \4264 );
and \U$3286 ( \4269 , \1457 , \2494 );
and \U$3287 ( \4270 , \1377 , \2492 );
nor \U$3288 ( \4271 , \4269 , \4270 );
xnor \U$3289 ( \4272 , \4271 , \2338 );
and \U$3290 ( \4273 , \1593 , \2222 );
and \U$3291 ( \4274 , \1531 , \2220 );
nor \U$3292 ( \4275 , \4273 , \4274 );
xnor \U$3293 ( \4276 , \4275 , \2109 );
and \U$3294 ( \4277 , \4272 , \4276 );
and \U$3295 ( \4278 , \1854 , \2028 );
and \U$3296 ( \4279 , \1656 , \2026 );
nor \U$3297 ( \4280 , \4278 , \4279 );
xnor \U$3298 ( \4281 , \4280 , \1892 );
and \U$3299 ( \4282 , \4276 , \4281 );
and \U$3300 ( \4283 , \4272 , \4281 );
or \U$3301 ( \4284 , \4277 , \4282 , \4283 );
and \U$3302 ( \4285 , \1162 , \3264 );
and \U$3303 ( \4286 , \1093 , \3262 );
nor \U$3304 ( \4287 , \4285 , \4286 );
xnor \U$3305 ( \4288 , \4287 , \3122 );
and \U$3306 ( \4289 , \1221 , \2968 );
and \U$3307 ( \4290 , \1167 , \2966 );
nor \U$3308 ( \4291 , \4289 , \4290 );
xnor \U$3309 ( \4292 , \4291 , \2831 );
and \U$3310 ( \4293 , \4288 , \4292 );
and \U$3311 ( \4294 , \1349 , \2762 );
and \U$3312 ( \4295 , \1272 , \2760 );
nor \U$3313 ( \4296 , \4294 , \4295 );
xnor \U$3314 ( \4297 , \4296 , \2610 );
and \U$3315 ( \4298 , \4292 , \4297 );
and \U$3316 ( \4299 , \4288 , \4297 );
or \U$3317 ( \4300 , \4293 , \4298 , \4299 );
and \U$3318 ( \4301 , \4284 , \4300 );
xor \U$3319 ( \4302 , \3784 , \4114 );
xor \U$3320 ( \4303 , \4114 , \4115 );
not \U$3321 ( \4304 , \4303 );
and \U$3322 ( \4305 , \4302 , \4304 );
and \U$3323 ( \4306 , \984 , \4305 );
not \U$3324 ( \4307 , \4306 );
xnor \U$3325 ( \4308 , \4307 , \4118 );
and \U$3326 ( \4309 , \1016 , \3992 );
and \U$3327 ( \4310 , \998 , \3990 );
nor \U$3328 ( \4311 , \4309 , \4310 );
xnor \U$3329 ( \4312 , \4311 , \3787 );
and \U$3330 ( \4313 , \4308 , \4312 );
and \U$3331 ( \4314 , \1085 , \3586 );
and \U$3332 ( \4315 , \1037 , \3584 );
nor \U$3333 ( \4316 , \4314 , \4315 );
xnor \U$3334 ( \4317 , \4316 , \3437 );
and \U$3335 ( \4318 , \4312 , \4317 );
and \U$3336 ( \4319 , \4308 , \4317 );
or \U$3337 ( \4320 , \4313 , \4318 , \4319 );
and \U$3338 ( \4321 , \4300 , \4320 );
and \U$3339 ( \4322 , \4284 , \4320 );
or \U$3340 ( \4323 , \4301 , \4321 , \4322 );
and \U$3341 ( \4324 , \2047 , \1828 );
and \U$3342 ( \4325 , \1942 , \1826 );
nor \U$3343 ( \4326 , \4324 , \4325 );
xnor \U$3344 ( \4327 , \4326 , \1750 );
and \U$3345 ( \4328 , \2168 , \1664 );
and \U$3346 ( \4329 , \2052 , \1662 );
nor \U$3347 ( \4330 , \4328 , \4329 );
xnor \U$3348 ( \4331 , \4330 , \1570 );
and \U$3349 ( \4332 , \4327 , \4331 );
and \U$3350 ( \4333 , \2459 , \1494 );
and \U$3351 ( \4334 , \2283 , \1492 );
nor \U$3352 ( \4335 , \4333 , \4334 );
xnor \U$3353 ( \4336 , \4335 , \1422 );
and \U$3354 ( \4337 , \4331 , \4336 );
and \U$3355 ( \4338 , \4327 , \4336 );
or \U$3356 ( \4339 , \4332 , \4337 , \4338 );
and \U$3357 ( \4340 , \3508 , \1076 );
and \U$3358 ( \4341 , \3334 , \1074 );
nor \U$3359 ( \4342 , \4340 , \4341 );
xnor \U$3360 ( \4343 , \4342 , \1046 );
and \U$3361 ( \4344 , \3813 , \1028 );
and \U$3362 ( \4345 , \3675 , \1026 );
nor \U$3363 ( \4346 , \4344 , \4345 );
xnor \U$3364 ( \4347 , \4346 , \1009 );
and \U$3365 ( \4348 , \4343 , \4347 );
buf \U$3366 ( \4349 , RIc0da468_99);
and \U$3367 ( \4350 , \4349 , \991 );
and \U$3368 ( \4351 , \3932 , \989 );
nor \U$3369 ( \4352 , \4350 , \4351 );
xnor \U$3370 ( \4353 , \4352 , \996 );
and \U$3371 ( \4354 , \4347 , \4353 );
and \U$3372 ( \4355 , \4343 , \4353 );
or \U$3373 ( \4356 , \4348 , \4354 , \4355 );
and \U$3374 ( \4357 , \4339 , \4356 );
and \U$3375 ( \4358 , \2710 , \1360 );
and \U$3376 ( \4359 , \2467 , \1358 );
nor \U$3377 ( \4360 , \4358 , \4359 );
xnor \U$3378 ( \4361 , \4360 , \1317 );
and \U$3379 ( \4362 , \2901 , \1247 );
and \U$3380 ( \4363 , \2715 , \1245 );
nor \U$3381 ( \4364 , \4362 , \4363 );
xnor \U$3382 ( \4365 , \4364 , \1198 );
and \U$3383 ( \4366 , \4361 , \4365 );
and \U$3384 ( \4367 , \3309 , \1146 );
and \U$3385 ( \4368 , \3045 , \1144 );
nor \U$3386 ( \4369 , \4367 , \4368 );
xnor \U$3387 ( \4370 , \4369 , \1105 );
and \U$3388 ( \4371 , \4365 , \4370 );
and \U$3389 ( \4372 , \4361 , \4370 );
or \U$3390 ( \4373 , \4366 , \4371 , \4372 );
and \U$3391 ( \4374 , \4356 , \4373 );
and \U$3392 ( \4375 , \4339 , \4373 );
or \U$3393 ( \4376 , \4357 , \4374 , \4375 );
and \U$3394 ( \4377 , \4323 , \4376 );
and \U$3395 ( \4378 , \4349 , \985 );
xor \U$3396 ( \4379 , \4155 , \4159 );
xor \U$3397 ( \4380 , \4379 , \4164 );
and \U$3398 ( \4381 , \4378 , \4380 );
xor \U$3399 ( \4382 , \4188 , \4192 );
xor \U$3400 ( \4383 , \4382 , \4197 );
and \U$3401 ( \4384 , \4380 , \4383 );
and \U$3402 ( \4385 , \4378 , \4383 );
or \U$3403 ( \4386 , \4381 , \4384 , \4385 );
and \U$3404 ( \4387 , \4376 , \4386 );
and \U$3405 ( \4388 , \4323 , \4386 );
or \U$3406 ( \4389 , \4377 , \4387 , \4388 );
xor \U$3407 ( \4390 , \4101 , \4105 );
xor \U$3408 ( \4391 , \4390 , \4110 );
xor \U$3409 ( \4392 , \4171 , \4175 );
xor \U$3410 ( \4393 , \4392 , \4180 );
and \U$3411 ( \4394 , \4391 , \4393 );
xor \U$3412 ( \4395 , \4136 , \4140 );
xor \U$3413 ( \4396 , \4395 , \4145 );
and \U$3414 ( \4397 , \4393 , \4396 );
and \U$3415 ( \4398 , \4391 , \4396 );
or \U$3416 ( \4399 , \4394 , \4397 , \4398 );
xor \U$3417 ( \4400 , \3995 , \3999 );
xor \U$3418 ( \4401 , \4400 , \4004 );
and \U$3419 ( \4402 , \4399 , \4401 );
xor \U$3420 ( \4403 , \4214 , \4216 );
xor \U$3421 ( \4404 , \4403 , \4219 );
and \U$3422 ( \4405 , \4401 , \4404 );
and \U$3423 ( \4406 , \4399 , \4404 );
or \U$3424 ( \4407 , \4402 , \4405 , \4406 );
and \U$3425 ( \4408 , \4389 , \4407 );
xor \U$3426 ( \4409 , \4113 , \4131 );
xor \U$3427 ( \4410 , \4409 , \4148 );
xor \U$3428 ( \4411 , \4167 , \4183 );
xor \U$3429 ( \4412 , \4411 , \4200 );
and \U$3430 ( \4413 , \4410 , \4412 );
xnor \U$3431 ( \4414 , \4206 , \4208 );
and \U$3432 ( \4415 , \4412 , \4414 );
and \U$3433 ( \4416 , \4410 , \4414 );
or \U$3434 ( \4417 , \4413 , \4415 , \4416 );
and \U$3435 ( \4418 , \4407 , \4417 );
and \U$3436 ( \4419 , \4389 , \4417 );
or \U$3437 ( \4420 , \4408 , \4418 , \4419 );
xor \U$3438 ( \4421 , \4151 , \4203 );
xor \U$3439 ( \4422 , \4421 , \4209 );
xor \U$3440 ( \4423 , \4222 , \4224 );
xor \U$3441 ( \4424 , \4423 , \4227 );
and \U$3442 ( \4425 , \4422 , \4424 );
xor \U$3443 ( \4426 , \4233 , \4235 );
and \U$3444 ( \4427 , \4424 , \4426 );
and \U$3445 ( \4428 , \4422 , \4426 );
or \U$3446 ( \4429 , \4425 , \4427 , \4428 );
and \U$3447 ( \4430 , \4420 , \4429 );
xor \U$3448 ( \4431 , \4241 , \4243 );
xor \U$3449 ( \4432 , \4431 , \4245 );
and \U$3450 ( \4433 , \4429 , \4432 );
and \U$3451 ( \4434 , \4420 , \4432 );
or \U$3452 ( \4435 , \4430 , \4433 , \4434 );
xor \U$3453 ( \4436 , \4041 , \4059 );
xor \U$3454 ( \4437 , \4436 , \4065 );
and \U$3455 ( \4438 , \4435 , \4437 );
xor \U$3456 ( \4439 , \4239 , \4248 );
xor \U$3457 ( \4440 , \4439 , \4251 );
and \U$3458 ( \4441 , \4437 , \4440 );
and \U$3459 ( \4442 , \4435 , \4440 );
or \U$3460 ( \4443 , \4438 , \4441 , \4442 );
xor \U$3461 ( \4444 , \4254 , \4256 );
xor \U$3462 ( \4445 , \4444 , \4259 );
and \U$3463 ( \4446 , \4443 , \4445 );
and \U$3464 ( \4447 , \4268 , \4446 );
xor \U$3465 ( \4448 , \4268 , \4446 );
xor \U$3466 ( \4449 , \4443 , \4445 );
buf \U$3467 ( \4450 , RIc0d87d0_38);
buf \U$3468 ( \4451 , RIc0d8848_39);
and \U$3469 ( \4452 , \4450 , \4451 );
not \U$3470 ( \4453 , \4452 );
and \U$3471 ( \4454 , \4115 , \4453 );
not \U$3472 ( \4455 , \4454 );
and \U$3473 ( \4456 , \998 , \4305 );
and \U$3474 ( \4457 , \984 , \4303 );
nor \U$3475 ( \4458 , \4456 , \4457 );
xnor \U$3476 ( \4459 , \4458 , \4118 );
and \U$3477 ( \4460 , \4455 , \4459 );
and \U$3478 ( \4461 , \1037 , \3992 );
and \U$3479 ( \4462 , \1016 , \3990 );
nor \U$3480 ( \4463 , \4461 , \4462 );
xnor \U$3481 ( \4464 , \4463 , \3787 );
and \U$3482 ( \4465 , \4459 , \4464 );
and \U$3483 ( \4466 , \4455 , \4464 );
or \U$3484 ( \4467 , \4460 , \4465 , \4466 );
and \U$3485 ( \4468 , \1093 , \3586 );
and \U$3486 ( \4469 , \1085 , \3584 );
nor \U$3487 ( \4470 , \4468 , \4469 );
xnor \U$3488 ( \4471 , \4470 , \3437 );
and \U$3489 ( \4472 , \1167 , \3264 );
and \U$3490 ( \4473 , \1162 , \3262 );
nor \U$3491 ( \4474 , \4472 , \4473 );
xnor \U$3492 ( \4475 , \4474 , \3122 );
and \U$3493 ( \4476 , \4471 , \4475 );
and \U$3494 ( \4477 , \1272 , \2968 );
and \U$3495 ( \4478 , \1221 , \2966 );
nor \U$3496 ( \4479 , \4477 , \4478 );
xnor \U$3497 ( \4480 , \4479 , \2831 );
and \U$3498 ( \4481 , \4475 , \4480 );
and \U$3499 ( \4482 , \4471 , \4480 );
or \U$3500 ( \4483 , \4476 , \4481 , \4482 );
and \U$3501 ( \4484 , \4467 , \4483 );
and \U$3502 ( \4485 , \1377 , \2762 );
and \U$3503 ( \4486 , \1349 , \2760 );
nor \U$3504 ( \4487 , \4485 , \4486 );
xnor \U$3505 ( \4488 , \4487 , \2610 );
and \U$3506 ( \4489 , \1531 , \2494 );
and \U$3507 ( \4490 , \1457 , \2492 );
nor \U$3508 ( \4491 , \4489 , \4490 );
xnor \U$3509 ( \4492 , \4491 , \2338 );
and \U$3510 ( \4493 , \4488 , \4492 );
and \U$3511 ( \4494 , \1656 , \2222 );
and \U$3512 ( \4495 , \1593 , \2220 );
nor \U$3513 ( \4496 , \4494 , \4495 );
xnor \U$3514 ( \4497 , \4496 , \2109 );
and \U$3515 ( \4498 , \4492 , \4497 );
and \U$3516 ( \4499 , \4488 , \4497 );
or \U$3517 ( \4500 , \4493 , \4498 , \4499 );
and \U$3518 ( \4501 , \4483 , \4500 );
and \U$3519 ( \4502 , \4467 , \4500 );
or \U$3520 ( \4503 , \4484 , \4501 , \4502 );
and \U$3521 ( \4504 , \2467 , \1494 );
and \U$3522 ( \4505 , \2459 , \1492 );
nor \U$3523 ( \4506 , \4504 , \4505 );
xnor \U$3524 ( \4507 , \4506 , \1422 );
and \U$3525 ( \4508 , \2715 , \1360 );
and \U$3526 ( \4509 , \2710 , \1358 );
nor \U$3527 ( \4510 , \4508 , \4509 );
xnor \U$3528 ( \4511 , \4510 , \1317 );
and \U$3529 ( \4512 , \4507 , \4511 );
and \U$3530 ( \4513 , \3045 , \1247 );
and \U$3531 ( \4514 , \2901 , \1245 );
nor \U$3532 ( \4515 , \4513 , \4514 );
xnor \U$3533 ( \4516 , \4515 , \1198 );
and \U$3534 ( \4517 , \4511 , \4516 );
and \U$3535 ( \4518 , \4507 , \4516 );
or \U$3536 ( \4519 , \4512 , \4517 , \4518 );
and \U$3537 ( \4520 , \1942 , \2028 );
and \U$3538 ( \4521 , \1854 , \2026 );
nor \U$3539 ( \4522 , \4520 , \4521 );
xnor \U$3540 ( \4523 , \4522 , \1892 );
and \U$3541 ( \4524 , \2052 , \1828 );
and \U$3542 ( \4525 , \2047 , \1826 );
nor \U$3543 ( \4526 , \4524 , \4525 );
xnor \U$3544 ( \4527 , \4526 , \1750 );
and \U$3545 ( \4528 , \4523 , \4527 );
and \U$3546 ( \4529 , \2283 , \1664 );
and \U$3547 ( \4530 , \2168 , \1662 );
nor \U$3548 ( \4531 , \4529 , \4530 );
xnor \U$3549 ( \4532 , \4531 , \1570 );
and \U$3550 ( \4533 , \4527 , \4532 );
and \U$3551 ( \4534 , \4523 , \4532 );
or \U$3552 ( \4535 , \4528 , \4533 , \4534 );
and \U$3553 ( \4536 , \4519 , \4535 );
and \U$3554 ( \4537 , \3334 , \1146 );
and \U$3555 ( \4538 , \3309 , \1144 );
nor \U$3556 ( \4539 , \4537 , \4538 );
xnor \U$3557 ( \4540 , \4539 , \1105 );
and \U$3558 ( \4541 , \3675 , \1076 );
and \U$3559 ( \4542 , \3508 , \1074 );
nor \U$3560 ( \4543 , \4541 , \4542 );
xnor \U$3561 ( \4544 , \4543 , \1046 );
and \U$3562 ( \4545 , \4540 , \4544 );
and \U$3563 ( \4546 , \3932 , \1028 );
and \U$3564 ( \4547 , \3813 , \1026 );
nor \U$3565 ( \4548 , \4546 , \4547 );
xnor \U$3566 ( \4549 , \4548 , \1009 );
and \U$3567 ( \4550 , \4544 , \4549 );
and \U$3568 ( \4551 , \4540 , \4549 );
or \U$3569 ( \4552 , \4545 , \4550 , \4551 );
and \U$3570 ( \4553 , \4535 , \4552 );
and \U$3571 ( \4554 , \4519 , \4552 );
or \U$3572 ( \4555 , \4536 , \4553 , \4554 );
and \U$3573 ( \4556 , \4503 , \4555 );
buf \U$3574 ( \4557 , RIc0da4e0_100);
and \U$3575 ( \4558 , \4557 , \985 );
xor \U$3576 ( \4559 , \4343 , \4347 );
xor \U$3577 ( \4560 , \4559 , \4353 );
or \U$3578 ( \4561 , \4558 , \4560 );
and \U$3579 ( \4562 , \4555 , \4561 );
and \U$3580 ( \4563 , \4503 , \4561 );
or \U$3581 ( \4564 , \4556 , \4562 , \4563 );
xor \U$3582 ( \4565 , \4272 , \4276 );
xor \U$3583 ( \4566 , \4565 , \4281 );
xor \U$3584 ( \4567 , \4327 , \4331 );
xor \U$3585 ( \4568 , \4567 , \4336 );
and \U$3586 ( \4569 , \4566 , \4568 );
xor \U$3587 ( \4570 , \4361 , \4365 );
xor \U$3588 ( \4571 , \4570 , \4370 );
and \U$3589 ( \4572 , \4568 , \4571 );
and \U$3590 ( \4573 , \4566 , \4571 );
or \U$3591 ( \4574 , \4569 , \4572 , \4573 );
xor \U$3592 ( \4575 , \4119 , \4123 );
xor \U$3593 ( \4576 , \4575 , \4128 );
and \U$3594 ( \4577 , \4574 , \4576 );
xor \U$3595 ( \4578 , \4391 , \4393 );
xor \U$3596 ( \4579 , \4578 , \4396 );
and \U$3597 ( \4580 , \4576 , \4579 );
and \U$3598 ( \4581 , \4574 , \4579 );
or \U$3599 ( \4582 , \4577 , \4580 , \4581 );
and \U$3600 ( \4583 , \4564 , \4582 );
xor \U$3601 ( \4584 , \4284 , \4300 );
xor \U$3602 ( \4585 , \4584 , \4320 );
xor \U$3603 ( \4586 , \4339 , \4356 );
xor \U$3604 ( \4587 , \4586 , \4373 );
and \U$3605 ( \4588 , \4585 , \4587 );
xor \U$3606 ( \4589 , \4378 , \4380 );
xor \U$3607 ( \4590 , \4589 , \4383 );
and \U$3608 ( \4591 , \4587 , \4590 );
and \U$3609 ( \4592 , \4585 , \4590 );
or \U$3610 ( \4593 , \4588 , \4591 , \4592 );
and \U$3611 ( \4594 , \4582 , \4593 );
and \U$3612 ( \4595 , \4564 , \4593 );
or \U$3613 ( \4596 , \4583 , \4594 , \4595 );
xor \U$3614 ( \4597 , \4323 , \4376 );
xor \U$3615 ( \4598 , \4597 , \4386 );
xor \U$3616 ( \4599 , \4399 , \4401 );
xor \U$3617 ( \4600 , \4599 , \4404 );
and \U$3618 ( \4601 , \4598 , \4600 );
xor \U$3619 ( \4602 , \4410 , \4412 );
xor \U$3620 ( \4603 , \4602 , \4414 );
and \U$3621 ( \4604 , \4600 , \4603 );
and \U$3622 ( \4605 , \4598 , \4603 );
or \U$3623 ( \4606 , \4601 , \4604 , \4605 );
and \U$3624 ( \4607 , \4596 , \4606 );
xor \U$3625 ( \4608 , \4422 , \4424 );
xor \U$3626 ( \4609 , \4608 , \4426 );
and \U$3627 ( \4610 , \4606 , \4609 );
and \U$3628 ( \4611 , \4596 , \4609 );
or \U$3629 ( \4612 , \4607 , \4610 , \4611 );
xor \U$3630 ( \4613 , \4212 , \4230 );
xor \U$3631 ( \4614 , \4613 , \4236 );
and \U$3632 ( \4615 , \4612 , \4614 );
xor \U$3633 ( \4616 , \4420 , \4429 );
xor \U$3634 ( \4617 , \4616 , \4432 );
and \U$3635 ( \4618 , \4614 , \4617 );
and \U$3636 ( \4619 , \4612 , \4617 );
or \U$3637 ( \4620 , \4615 , \4618 , \4619 );
xor \U$3638 ( \4621 , \4435 , \4437 );
xor \U$3639 ( \4622 , \4621 , \4440 );
and \U$3640 ( \4623 , \4620 , \4622 );
and \U$3641 ( \4624 , \4449 , \4623 );
xor \U$3642 ( \4625 , \4449 , \4623 );
xor \U$3643 ( \4626 , \4620 , \4622 );
and \U$3644 ( \4627 , \2047 , \2028 );
and \U$3645 ( \4628 , \1942 , \2026 );
nor \U$3646 ( \4629 , \4627 , \4628 );
xnor \U$3647 ( \4630 , \4629 , \1892 );
and \U$3648 ( \4631 , \2168 , \1828 );
and \U$3649 ( \4632 , \2052 , \1826 );
nor \U$3650 ( \4633 , \4631 , \4632 );
xnor \U$3651 ( \4634 , \4633 , \1750 );
and \U$3652 ( \4635 , \4630 , \4634 );
and \U$3653 ( \4636 , \2459 , \1664 );
and \U$3654 ( \4637 , \2283 , \1662 );
nor \U$3655 ( \4638 , \4636 , \4637 );
xnor \U$3656 ( \4639 , \4638 , \1570 );
and \U$3657 ( \4640 , \4634 , \4639 );
and \U$3658 ( \4641 , \4630 , \4639 );
or \U$3659 ( \4642 , \4635 , \4640 , \4641 );
and \U$3660 ( \4643 , \2710 , \1494 );
and \U$3661 ( \4644 , \2467 , \1492 );
nor \U$3662 ( \4645 , \4643 , \4644 );
xnor \U$3663 ( \4646 , \4645 , \1422 );
and \U$3664 ( \4647 , \2901 , \1360 );
and \U$3665 ( \4648 , \2715 , \1358 );
nor \U$3666 ( \4649 , \4647 , \4648 );
xnor \U$3667 ( \4650 , \4649 , \1317 );
and \U$3668 ( \4651 , \4646 , \4650 );
and \U$3669 ( \4652 , \3309 , \1247 );
and \U$3670 ( \4653 , \3045 , \1245 );
nor \U$3671 ( \4654 , \4652 , \4653 );
xnor \U$3672 ( \4655 , \4654 , \1198 );
and \U$3673 ( \4656 , \4650 , \4655 );
and \U$3674 ( \4657 , \4646 , \4655 );
or \U$3675 ( \4658 , \4651 , \4656 , \4657 );
and \U$3676 ( \4659 , \4642 , \4658 );
and \U$3677 ( \4660 , \3508 , \1146 );
and \U$3678 ( \4661 , \3334 , \1144 );
nor \U$3679 ( \4662 , \4660 , \4661 );
xnor \U$3680 ( \4663 , \4662 , \1105 );
and \U$3681 ( \4664 , \3813 , \1076 );
and \U$3682 ( \4665 , \3675 , \1074 );
nor \U$3683 ( \4666 , \4664 , \4665 );
xnor \U$3684 ( \4667 , \4666 , \1046 );
and \U$3685 ( \4668 , \4663 , \4667 );
and \U$3686 ( \4669 , \4349 , \1028 );
and \U$3687 ( \4670 , \3932 , \1026 );
nor \U$3688 ( \4671 , \4669 , \4670 );
xnor \U$3689 ( \4672 , \4671 , \1009 );
and \U$3690 ( \4673 , \4667 , \4672 );
and \U$3691 ( \4674 , \4663 , \4672 );
or \U$3692 ( \4675 , \4668 , \4673 , \4674 );
and \U$3693 ( \4676 , \4658 , \4675 );
and \U$3694 ( \4677 , \4642 , \4675 );
or \U$3695 ( \4678 , \4659 , \4676 , \4677 );
buf \U$3696 ( \4679 , RIc0da558_101);
and \U$3697 ( \4680 , \4679 , \991 );
and \U$3698 ( \4681 , \4557 , \989 );
nor \U$3699 ( \4682 , \4680 , \4681 );
xnor \U$3700 ( \4683 , \4682 , \996 );
buf \U$3701 ( \4684 , RIc0da5d0_102);
and \U$3702 ( \4685 , \4684 , \985 );
or \U$3703 ( \4686 , \4683 , \4685 );
and \U$3704 ( \4687 , \4557 , \991 );
and \U$3705 ( \4688 , \4349 , \989 );
nor \U$3706 ( \4689 , \4687 , \4688 );
xnor \U$3707 ( \4690 , \4689 , \996 );
and \U$3708 ( \4691 , \4686 , \4690 );
and \U$3709 ( \4692 , \4679 , \985 );
and \U$3710 ( \4693 , \4690 , \4692 );
and \U$3711 ( \4694 , \4686 , \4692 );
or \U$3712 ( \4695 , \4691 , \4693 , \4694 );
and \U$3713 ( \4696 , \4678 , \4695 );
xor \U$3714 ( \4697 , \4115 , \4450 );
xor \U$3715 ( \4698 , \4450 , \4451 );
not \U$3716 ( \4699 , \4698 );
and \U$3717 ( \4700 , \4697 , \4699 );
and \U$3718 ( \4701 , \984 , \4700 );
not \U$3719 ( \4702 , \4701 );
xnor \U$3720 ( \4703 , \4702 , \4454 );
and \U$3721 ( \4704 , \1016 , \4305 );
and \U$3722 ( \4705 , \998 , \4303 );
nor \U$3723 ( \4706 , \4704 , \4705 );
xnor \U$3724 ( \4707 , \4706 , \4118 );
and \U$3725 ( \4708 , \4703 , \4707 );
and \U$3726 ( \4709 , \1085 , \3992 );
and \U$3727 ( \4710 , \1037 , \3990 );
nor \U$3728 ( \4711 , \4709 , \4710 );
xnor \U$3729 ( \4712 , \4711 , \3787 );
and \U$3730 ( \4713 , \4707 , \4712 );
and \U$3731 ( \4714 , \4703 , \4712 );
or \U$3732 ( \4715 , \4708 , \4713 , \4714 );
and \U$3733 ( \4716 , \1162 , \3586 );
and \U$3734 ( \4717 , \1093 , \3584 );
nor \U$3735 ( \4718 , \4716 , \4717 );
xnor \U$3736 ( \4719 , \4718 , \3437 );
and \U$3737 ( \4720 , \1221 , \3264 );
and \U$3738 ( \4721 , \1167 , \3262 );
nor \U$3739 ( \4722 , \4720 , \4721 );
xnor \U$3740 ( \4723 , \4722 , \3122 );
and \U$3741 ( \4724 , \4719 , \4723 );
and \U$3742 ( \4725 , \1349 , \2968 );
and \U$3743 ( \4726 , \1272 , \2966 );
nor \U$3744 ( \4727 , \4725 , \4726 );
xnor \U$3745 ( \4728 , \4727 , \2831 );
and \U$3746 ( \4729 , \4723 , \4728 );
and \U$3747 ( \4730 , \4719 , \4728 );
or \U$3748 ( \4731 , \4724 , \4729 , \4730 );
and \U$3749 ( \4732 , \4715 , \4731 );
and \U$3750 ( \4733 , \1457 , \2762 );
and \U$3751 ( \4734 , \1377 , \2760 );
nor \U$3752 ( \4735 , \4733 , \4734 );
xnor \U$3753 ( \4736 , \4735 , \2610 );
and \U$3754 ( \4737 , \1593 , \2494 );
and \U$3755 ( \4738 , \1531 , \2492 );
nor \U$3756 ( \4739 , \4737 , \4738 );
xnor \U$3757 ( \4740 , \4739 , \2338 );
and \U$3758 ( \4741 , \4736 , \4740 );
and \U$3759 ( \4742 , \1854 , \2222 );
and \U$3760 ( \4743 , \1656 , \2220 );
nor \U$3761 ( \4744 , \4742 , \4743 );
xnor \U$3762 ( \4745 , \4744 , \2109 );
and \U$3763 ( \4746 , \4740 , \4745 );
and \U$3764 ( \4747 , \4736 , \4745 );
or \U$3765 ( \4748 , \4741 , \4746 , \4747 );
and \U$3766 ( \4749 , \4731 , \4748 );
and \U$3767 ( \4750 , \4715 , \4748 );
or \U$3768 ( \4751 , \4732 , \4749 , \4750 );
and \U$3769 ( \4752 , \4695 , \4751 );
and \U$3770 ( \4753 , \4678 , \4751 );
or \U$3771 ( \4754 , \4696 , \4752 , \4753 );
xor \U$3772 ( \4755 , \4507 , \4511 );
xor \U$3773 ( \4756 , \4755 , \4516 );
xor \U$3774 ( \4757 , \4523 , \4527 );
xor \U$3775 ( \4758 , \4757 , \4532 );
and \U$3776 ( \4759 , \4756 , \4758 );
xor \U$3777 ( \4760 , \4540 , \4544 );
xor \U$3778 ( \4761 , \4760 , \4549 );
and \U$3779 ( \4762 , \4758 , \4761 );
and \U$3780 ( \4763 , \4756 , \4761 );
or \U$3781 ( \4764 , \4759 , \4762 , \4763 );
xor \U$3782 ( \4765 , \4455 , \4459 );
xor \U$3783 ( \4766 , \4765 , \4464 );
xor \U$3784 ( \4767 , \4471 , \4475 );
xor \U$3785 ( \4768 , \4767 , \4480 );
and \U$3786 ( \4769 , \4766 , \4768 );
xor \U$3787 ( \4770 , \4488 , \4492 );
xor \U$3788 ( \4771 , \4770 , \4497 );
and \U$3789 ( \4772 , \4768 , \4771 );
and \U$3790 ( \4773 , \4766 , \4771 );
or \U$3791 ( \4774 , \4769 , \4772 , \4773 );
and \U$3792 ( \4775 , \4764 , \4774 );
xor \U$3793 ( \4776 , \4288 , \4292 );
xor \U$3794 ( \4777 , \4776 , \4297 );
and \U$3795 ( \4778 , \4774 , \4777 );
and \U$3796 ( \4779 , \4764 , \4777 );
or \U$3797 ( \4780 , \4775 , \4778 , \4779 );
and \U$3798 ( \4781 , \4754 , \4780 );
xor \U$3799 ( \4782 , \4308 , \4312 );
xor \U$3800 ( \4783 , \4782 , \4317 );
xor \U$3801 ( \4784 , \4566 , \4568 );
xor \U$3802 ( \4785 , \4784 , \4571 );
and \U$3803 ( \4786 , \4783 , \4785 );
xnor \U$3804 ( \4787 , \4558 , \4560 );
and \U$3805 ( \4788 , \4785 , \4787 );
and \U$3806 ( \4789 , \4783 , \4787 );
or \U$3807 ( \4790 , \4786 , \4788 , \4789 );
and \U$3808 ( \4791 , \4780 , \4790 );
and \U$3809 ( \4792 , \4754 , \4790 );
or \U$3810 ( \4793 , \4781 , \4791 , \4792 );
xor \U$3811 ( \4794 , \4503 , \4555 );
xor \U$3812 ( \4795 , \4794 , \4561 );
xor \U$3813 ( \4796 , \4574 , \4576 );
xor \U$3814 ( \4797 , \4796 , \4579 );
and \U$3815 ( \4798 , \4795 , \4797 );
xor \U$3816 ( \4799 , \4585 , \4587 );
xor \U$3817 ( \4800 , \4799 , \4590 );
and \U$3818 ( \4801 , \4797 , \4800 );
and \U$3819 ( \4802 , \4795 , \4800 );
or \U$3820 ( \4803 , \4798 , \4801 , \4802 );
and \U$3821 ( \4804 , \4793 , \4803 );
xor \U$3822 ( \4805 , \4598 , \4600 );
xor \U$3823 ( \4806 , \4805 , \4603 );
and \U$3824 ( \4807 , \4803 , \4806 );
and \U$3825 ( \4808 , \4793 , \4806 );
or \U$3826 ( \4809 , \4804 , \4807 , \4808 );
xor \U$3827 ( \4810 , \4389 , \4407 );
xor \U$3828 ( \4811 , \4810 , \4417 );
and \U$3829 ( \4812 , \4809 , \4811 );
xor \U$3830 ( \4813 , \4596 , \4606 );
xor \U$3831 ( \4814 , \4813 , \4609 );
and \U$3832 ( \4815 , \4811 , \4814 );
and \U$3833 ( \4816 , \4809 , \4814 );
or \U$3834 ( \4817 , \4812 , \4815 , \4816 );
xor \U$3835 ( \4818 , \4612 , \4614 );
xor \U$3836 ( \4819 , \4818 , \4617 );
and \U$3837 ( \4820 , \4817 , \4819 );
and \U$3838 ( \4821 , \4626 , \4820 );
xor \U$3839 ( \4822 , \4626 , \4820 );
xor \U$3840 ( \4823 , \4817 , \4819 );
and \U$3841 ( \4824 , \2467 , \1664 );
and \U$3842 ( \4825 , \2459 , \1662 );
nor \U$3843 ( \4826 , \4824 , \4825 );
xnor \U$3844 ( \4827 , \4826 , \1570 );
and \U$3845 ( \4828 , \2715 , \1494 );
and \U$3846 ( \4829 , \2710 , \1492 );
nor \U$3847 ( \4830 , \4828 , \4829 );
xnor \U$3848 ( \4831 , \4830 , \1422 );
and \U$3849 ( \4832 , \4827 , \4831 );
and \U$3850 ( \4833 , \3045 , \1360 );
and \U$3851 ( \4834 , \2901 , \1358 );
nor \U$3852 ( \4835 , \4833 , \4834 );
xnor \U$3853 ( \4836 , \4835 , \1317 );
and \U$3854 ( \4837 , \4831 , \4836 );
and \U$3855 ( \4838 , \4827 , \4836 );
or \U$3856 ( \4839 , \4832 , \4837 , \4838 );
and \U$3857 ( \4840 , \1942 , \2222 );
and \U$3858 ( \4841 , \1854 , \2220 );
nor \U$3859 ( \4842 , \4840 , \4841 );
xnor \U$3860 ( \4843 , \4842 , \2109 );
and \U$3861 ( \4844 , \2052 , \2028 );
and \U$3862 ( \4845 , \2047 , \2026 );
nor \U$3863 ( \4846 , \4844 , \4845 );
xnor \U$3864 ( \4847 , \4846 , \1892 );
and \U$3865 ( \4848 , \4843 , \4847 );
and \U$3866 ( \4849 , \2283 , \1828 );
and \U$3867 ( \4850 , \2168 , \1826 );
nor \U$3868 ( \4851 , \4849 , \4850 );
xnor \U$3869 ( \4852 , \4851 , \1750 );
and \U$3870 ( \4853 , \4847 , \4852 );
and \U$3871 ( \4854 , \4843 , \4852 );
or \U$3872 ( \4855 , \4848 , \4853 , \4854 );
and \U$3873 ( \4856 , \4839 , \4855 );
and \U$3874 ( \4857 , \3334 , \1247 );
and \U$3875 ( \4858 , \3309 , \1245 );
nor \U$3876 ( \4859 , \4857 , \4858 );
xnor \U$3877 ( \4860 , \4859 , \1198 );
and \U$3878 ( \4861 , \3675 , \1146 );
and \U$3879 ( \4862 , \3508 , \1144 );
nor \U$3880 ( \4863 , \4861 , \4862 );
xnor \U$3881 ( \4864 , \4863 , \1105 );
and \U$3882 ( \4865 , \4860 , \4864 );
and \U$3883 ( \4866 , \3932 , \1076 );
and \U$3884 ( \4867 , \3813 , \1074 );
nor \U$3885 ( \4868 , \4866 , \4867 );
xnor \U$3886 ( \4869 , \4868 , \1046 );
and \U$3887 ( \4870 , \4864 , \4869 );
and \U$3888 ( \4871 , \4860 , \4869 );
or \U$3889 ( \4872 , \4865 , \4870 , \4871 );
and \U$3890 ( \4873 , \4855 , \4872 );
and \U$3891 ( \4874 , \4839 , \4872 );
or \U$3892 ( \4875 , \4856 , \4873 , \4874 );
buf \U$3893 ( \4876 , RIc0d88c0_40);
buf \U$3894 ( \4877 , RIc0d8938_41);
and \U$3895 ( \4878 , \4876 , \4877 );
not \U$3896 ( \4879 , \4878 );
and \U$3897 ( \4880 , \4451 , \4879 );
not \U$3898 ( \4881 , \4880 );
and \U$3899 ( \4882 , \998 , \4700 );
and \U$3900 ( \4883 , \984 , \4698 );
nor \U$3901 ( \4884 , \4882 , \4883 );
xnor \U$3902 ( \4885 , \4884 , \4454 );
and \U$3903 ( \4886 , \4881 , \4885 );
and \U$3904 ( \4887 , \1037 , \4305 );
and \U$3905 ( \4888 , \1016 , \4303 );
nor \U$3906 ( \4889 , \4887 , \4888 );
xnor \U$3907 ( \4890 , \4889 , \4118 );
and \U$3908 ( \4891 , \4885 , \4890 );
and \U$3909 ( \4892 , \4881 , \4890 );
or \U$3910 ( \4893 , \4886 , \4891 , \4892 );
and \U$3911 ( \4894 , \1093 , \3992 );
and \U$3912 ( \4895 , \1085 , \3990 );
nor \U$3913 ( \4896 , \4894 , \4895 );
xnor \U$3914 ( \4897 , \4896 , \3787 );
and \U$3915 ( \4898 , \1167 , \3586 );
and \U$3916 ( \4899 , \1162 , \3584 );
nor \U$3917 ( \4900 , \4898 , \4899 );
xnor \U$3918 ( \4901 , \4900 , \3437 );
and \U$3919 ( \4902 , \4897 , \4901 );
and \U$3920 ( \4903 , \1272 , \3264 );
and \U$3921 ( \4904 , \1221 , \3262 );
nor \U$3922 ( \4905 , \4903 , \4904 );
xnor \U$3923 ( \4906 , \4905 , \3122 );
and \U$3924 ( \4907 , \4901 , \4906 );
and \U$3925 ( \4908 , \4897 , \4906 );
or \U$3926 ( \4909 , \4902 , \4907 , \4908 );
and \U$3927 ( \4910 , \4893 , \4909 );
and \U$3928 ( \4911 , \1377 , \2968 );
and \U$3929 ( \4912 , \1349 , \2966 );
nor \U$3930 ( \4913 , \4911 , \4912 );
xnor \U$3931 ( \4914 , \4913 , \2831 );
and \U$3932 ( \4915 , \1531 , \2762 );
and \U$3933 ( \4916 , \1457 , \2760 );
nor \U$3934 ( \4917 , \4915 , \4916 );
xnor \U$3935 ( \4918 , \4917 , \2610 );
and \U$3936 ( \4919 , \4914 , \4918 );
and \U$3937 ( \4920 , \1656 , \2494 );
and \U$3938 ( \4921 , \1593 , \2492 );
nor \U$3939 ( \4922 , \4920 , \4921 );
xnor \U$3940 ( \4923 , \4922 , \2338 );
and \U$3941 ( \4924 , \4918 , \4923 );
and \U$3942 ( \4925 , \4914 , \4923 );
or \U$3943 ( \4926 , \4919 , \4924 , \4925 );
and \U$3944 ( \4927 , \4909 , \4926 );
and \U$3945 ( \4928 , \4893 , \4926 );
or \U$3946 ( \4929 , \4910 , \4927 , \4928 );
and \U$3947 ( \4930 , \4875 , \4929 );
and \U$3948 ( \4931 , \4557 , \1028 );
and \U$3949 ( \4932 , \4349 , \1026 );
nor \U$3950 ( \4933 , \4931 , \4932 );
xnor \U$3951 ( \4934 , \4933 , \1009 );
and \U$3952 ( \4935 , \4684 , \991 );
and \U$3953 ( \4936 , \4679 , \989 );
nor \U$3954 ( \4937 , \4935 , \4936 );
xnor \U$3955 ( \4938 , \4937 , \996 );
and \U$3956 ( \4939 , \4934 , \4938 );
buf \U$3957 ( \4940 , RIc0da648_103);
and \U$3958 ( \4941 , \4940 , \985 );
and \U$3959 ( \4942 , \4938 , \4941 );
and \U$3960 ( \4943 , \4934 , \4941 );
or \U$3961 ( \4944 , \4939 , \4942 , \4943 );
xor \U$3962 ( \4945 , \4663 , \4667 );
xor \U$3963 ( \4946 , \4945 , \4672 );
and \U$3964 ( \4947 , \4944 , \4946 );
xnor \U$3965 ( \4948 , \4683 , \4685 );
and \U$3966 ( \4949 , \4946 , \4948 );
and \U$3967 ( \4950 , \4944 , \4948 );
or \U$3968 ( \4951 , \4947 , \4949 , \4950 );
and \U$3969 ( \4952 , \4929 , \4951 );
and \U$3970 ( \4953 , \4875 , \4951 );
or \U$3971 ( \4954 , \4930 , \4952 , \4953 );
xor \U$3972 ( \4955 , \4630 , \4634 );
xor \U$3973 ( \4956 , \4955 , \4639 );
xor \U$3974 ( \4957 , \4646 , \4650 );
xor \U$3975 ( \4958 , \4957 , \4655 );
and \U$3976 ( \4959 , \4956 , \4958 );
xor \U$3977 ( \4960 , \4736 , \4740 );
xor \U$3978 ( \4961 , \4960 , \4745 );
and \U$3979 ( \4962 , \4958 , \4961 );
and \U$3980 ( \4963 , \4956 , \4961 );
or \U$3981 ( \4964 , \4959 , \4962 , \4963 );
xor \U$3982 ( \4965 , \4703 , \4707 );
xor \U$3983 ( \4966 , \4965 , \4712 );
xor \U$3984 ( \4967 , \4719 , \4723 );
xor \U$3985 ( \4968 , \4967 , \4728 );
and \U$3986 ( \4969 , \4966 , \4968 );
and \U$3987 ( \4970 , \4964 , \4969 );
xor \U$3988 ( \4971 , \4766 , \4768 );
xor \U$3989 ( \4972 , \4971 , \4771 );
and \U$3990 ( \4973 , \4969 , \4972 );
and \U$3991 ( \4974 , \4964 , \4972 );
or \U$3992 ( \4975 , \4970 , \4973 , \4974 );
and \U$3993 ( \4976 , \4954 , \4975 );
xor \U$3994 ( \4977 , \4642 , \4658 );
xor \U$3995 ( \4978 , \4977 , \4675 );
xor \U$3996 ( \4979 , \4686 , \4690 );
xor \U$3997 ( \4980 , \4979 , \4692 );
and \U$3998 ( \4981 , \4978 , \4980 );
xor \U$3999 ( \4982 , \4756 , \4758 );
xor \U$4000 ( \4983 , \4982 , \4761 );
and \U$4001 ( \4984 , \4980 , \4983 );
and \U$4002 ( \4985 , \4978 , \4983 );
or \U$4003 ( \4986 , \4981 , \4984 , \4985 );
and \U$4004 ( \4987 , \4975 , \4986 );
and \U$4005 ( \4988 , \4954 , \4986 );
or \U$4006 ( \4989 , \4976 , \4987 , \4988 );
xor \U$4007 ( \4990 , \4467 , \4483 );
xor \U$4008 ( \4991 , \4990 , \4500 );
xor \U$4009 ( \4992 , \4519 , \4535 );
xor \U$4010 ( \4993 , \4992 , \4552 );
and \U$4011 ( \4994 , \4991 , \4993 );
xor \U$4012 ( \4995 , \4783 , \4785 );
xor \U$4013 ( \4996 , \4995 , \4787 );
and \U$4014 ( \4997 , \4993 , \4996 );
and \U$4015 ( \4998 , \4991 , \4996 );
or \U$4016 ( \4999 , \4994 , \4997 , \4998 );
and \U$4017 ( \5000 , \4989 , \4999 );
xor \U$4018 ( \5001 , \4795 , \4797 );
xor \U$4019 ( \5002 , \5001 , \4800 );
and \U$4020 ( \5003 , \4999 , \5002 );
and \U$4021 ( \5004 , \4989 , \5002 );
or \U$4022 ( \5005 , \5000 , \5003 , \5004 );
xor \U$4023 ( \5006 , \4564 , \4582 );
xor \U$4024 ( \5007 , \5006 , \4593 );
and \U$4025 ( \5008 , \5005 , \5007 );
xor \U$4026 ( \5009 , \4793 , \4803 );
xor \U$4027 ( \5010 , \5009 , \4806 );
and \U$4028 ( \5011 , \5007 , \5010 );
and \U$4029 ( \5012 , \5005 , \5010 );
or \U$4030 ( \5013 , \5008 , \5011 , \5012 );
xor \U$4031 ( \5014 , \4809 , \4811 );
xor \U$4032 ( \5015 , \5014 , \4814 );
and \U$4033 ( \5016 , \5013 , \5015 );
and \U$4034 ( \5017 , \4823 , \5016 );
xor \U$4035 ( \5018 , \4823 , \5016 );
xor \U$4036 ( \5019 , \5013 , \5015 );
xor \U$4037 ( \5020 , \4451 , \4876 );
xor \U$4038 ( \5021 , \4876 , \4877 );
not \U$4039 ( \5022 , \5021 );
and \U$4040 ( \5023 , \5020 , \5022 );
and \U$4041 ( \5024 , \984 , \5023 );
not \U$4042 ( \5025 , \5024 );
xnor \U$4043 ( \5026 , \5025 , \4880 );
and \U$4044 ( \5027 , \1016 , \4700 );
and \U$4045 ( \5028 , \998 , \4698 );
nor \U$4046 ( \5029 , \5027 , \5028 );
xnor \U$4047 ( \5030 , \5029 , \4454 );
and \U$4048 ( \5031 , \5026 , \5030 );
and \U$4049 ( \5032 , \1085 , \4305 );
and \U$4050 ( \5033 , \1037 , \4303 );
nor \U$4051 ( \5034 , \5032 , \5033 );
xnor \U$4052 ( \5035 , \5034 , \4118 );
and \U$4053 ( \5036 , \5030 , \5035 );
and \U$4054 ( \5037 , \5026 , \5035 );
or \U$4055 ( \5038 , \5031 , \5036 , \5037 );
and \U$4056 ( \5039 , \1162 , \3992 );
and \U$4057 ( \5040 , \1093 , \3990 );
nor \U$4058 ( \5041 , \5039 , \5040 );
xnor \U$4059 ( \5042 , \5041 , \3787 );
and \U$4060 ( \5043 , \1221 , \3586 );
and \U$4061 ( \5044 , \1167 , \3584 );
nor \U$4062 ( \5045 , \5043 , \5044 );
xnor \U$4063 ( \5046 , \5045 , \3437 );
and \U$4064 ( \5047 , \5042 , \5046 );
and \U$4065 ( \5048 , \1349 , \3264 );
and \U$4066 ( \5049 , \1272 , \3262 );
nor \U$4067 ( \5050 , \5048 , \5049 );
xnor \U$4068 ( \5051 , \5050 , \3122 );
and \U$4069 ( \5052 , \5046 , \5051 );
and \U$4070 ( \5053 , \5042 , \5051 );
or \U$4071 ( \5054 , \5047 , \5052 , \5053 );
and \U$4072 ( \5055 , \5038 , \5054 );
and \U$4073 ( \5056 , \1457 , \2968 );
and \U$4074 ( \5057 , \1377 , \2966 );
nor \U$4075 ( \5058 , \5056 , \5057 );
xnor \U$4076 ( \5059 , \5058 , \2831 );
and \U$4077 ( \5060 , \1593 , \2762 );
and \U$4078 ( \5061 , \1531 , \2760 );
nor \U$4079 ( \5062 , \5060 , \5061 );
xnor \U$4080 ( \5063 , \5062 , \2610 );
and \U$4081 ( \5064 , \5059 , \5063 );
and \U$4082 ( \5065 , \1854 , \2494 );
and \U$4083 ( \5066 , \1656 , \2492 );
nor \U$4084 ( \5067 , \5065 , \5066 );
xnor \U$4085 ( \5068 , \5067 , \2338 );
and \U$4086 ( \5069 , \5063 , \5068 );
and \U$4087 ( \5070 , \5059 , \5068 );
or \U$4088 ( \5071 , \5064 , \5069 , \5070 );
and \U$4089 ( \5072 , \5054 , \5071 );
and \U$4090 ( \5073 , \5038 , \5071 );
or \U$4091 ( \5074 , \5055 , \5072 , \5073 );
and \U$4092 ( \5075 , \3508 , \1247 );
and \U$4093 ( \5076 , \3334 , \1245 );
nor \U$4094 ( \5077 , \5075 , \5076 );
xnor \U$4095 ( \5078 , \5077 , \1198 );
and \U$4096 ( \5079 , \3813 , \1146 );
and \U$4097 ( \5080 , \3675 , \1144 );
nor \U$4098 ( \5081 , \5079 , \5080 );
xnor \U$4099 ( \5082 , \5081 , \1105 );
and \U$4100 ( \5083 , \5078 , \5082 );
and \U$4101 ( \5084 , \4349 , \1076 );
and \U$4102 ( \5085 , \3932 , \1074 );
nor \U$4103 ( \5086 , \5084 , \5085 );
xnor \U$4104 ( \5087 , \5086 , \1046 );
and \U$4105 ( \5088 , \5082 , \5087 );
and \U$4106 ( \5089 , \5078 , \5087 );
or \U$4107 ( \5090 , \5083 , \5088 , \5089 );
and \U$4108 ( \5091 , \2047 , \2222 );
and \U$4109 ( \5092 , \1942 , \2220 );
nor \U$4110 ( \5093 , \5091 , \5092 );
xnor \U$4111 ( \5094 , \5093 , \2109 );
and \U$4112 ( \5095 , \2168 , \2028 );
and \U$4113 ( \5096 , \2052 , \2026 );
nor \U$4114 ( \5097 , \5095 , \5096 );
xnor \U$4115 ( \5098 , \5097 , \1892 );
and \U$4116 ( \5099 , \5094 , \5098 );
and \U$4117 ( \5100 , \2459 , \1828 );
and \U$4118 ( \5101 , \2283 , \1826 );
nor \U$4119 ( \5102 , \5100 , \5101 );
xnor \U$4120 ( \5103 , \5102 , \1750 );
and \U$4121 ( \5104 , \5098 , \5103 );
and \U$4122 ( \5105 , \5094 , \5103 );
or \U$4123 ( \5106 , \5099 , \5104 , \5105 );
and \U$4124 ( \5107 , \5090 , \5106 );
and \U$4125 ( \5108 , \2710 , \1664 );
and \U$4126 ( \5109 , \2467 , \1662 );
nor \U$4127 ( \5110 , \5108 , \5109 );
xnor \U$4128 ( \5111 , \5110 , \1570 );
and \U$4129 ( \5112 , \2901 , \1494 );
and \U$4130 ( \5113 , \2715 , \1492 );
nor \U$4131 ( \5114 , \5112 , \5113 );
xnor \U$4132 ( \5115 , \5114 , \1422 );
and \U$4133 ( \5116 , \5111 , \5115 );
and \U$4134 ( \5117 , \3309 , \1360 );
and \U$4135 ( \5118 , \3045 , \1358 );
nor \U$4136 ( \5119 , \5117 , \5118 );
xnor \U$4137 ( \5120 , \5119 , \1317 );
and \U$4138 ( \5121 , \5115 , \5120 );
and \U$4139 ( \5122 , \5111 , \5120 );
or \U$4140 ( \5123 , \5116 , \5121 , \5122 );
and \U$4141 ( \5124 , \5106 , \5123 );
and \U$4142 ( \5125 , \5090 , \5123 );
or \U$4143 ( \5126 , \5107 , \5124 , \5125 );
and \U$4144 ( \5127 , \5074 , \5126 );
and \U$4145 ( \5128 , \4679 , \1028 );
and \U$4146 ( \5129 , \4557 , \1026 );
nor \U$4147 ( \5130 , \5128 , \5129 );
xnor \U$4148 ( \5131 , \5130 , \1009 );
and \U$4149 ( \5132 , \4940 , \991 );
and \U$4150 ( \5133 , \4684 , \989 );
nor \U$4151 ( \5134 , \5132 , \5133 );
xnor \U$4152 ( \5135 , \5134 , \996 );
and \U$4153 ( \5136 , \5131 , \5135 );
buf \U$4154 ( \5137 , RIc0da6c0_104);
and \U$4155 ( \5138 , \5137 , \985 );
and \U$4156 ( \5139 , \5135 , \5138 );
and \U$4157 ( \5140 , \5131 , \5138 );
or \U$4158 ( \5141 , \5136 , \5139 , \5140 );
xor \U$4159 ( \5142 , \4934 , \4938 );
xor \U$4160 ( \5143 , \5142 , \4941 );
and \U$4161 ( \5144 , \5141 , \5143 );
xor \U$4162 ( \5145 , \4860 , \4864 );
xor \U$4163 ( \5146 , \5145 , \4869 );
and \U$4164 ( \5147 , \5143 , \5146 );
and \U$4165 ( \5148 , \5141 , \5146 );
or \U$4166 ( \5149 , \5144 , \5147 , \5148 );
and \U$4167 ( \5150 , \5126 , \5149 );
and \U$4168 ( \5151 , \5074 , \5149 );
or \U$4169 ( \5152 , \5127 , \5150 , \5151 );
xor \U$4170 ( \5153 , \4839 , \4855 );
xor \U$4171 ( \5154 , \5153 , \4872 );
xor \U$4172 ( \5155 , \4893 , \4909 );
xor \U$4173 ( \5156 , \5155 , \4926 );
and \U$4174 ( \5157 , \5154 , \5156 );
xor \U$4175 ( \5158 , \4944 , \4946 );
xor \U$4176 ( \5159 , \5158 , \4948 );
and \U$4177 ( \5160 , \5156 , \5159 );
and \U$4178 ( \5161 , \5154 , \5159 );
or \U$4179 ( \5162 , \5157 , \5160 , \5161 );
and \U$4180 ( \5163 , \5152 , \5162 );
xor \U$4181 ( \5164 , \4827 , \4831 );
xor \U$4182 ( \5165 , \5164 , \4836 );
xor \U$4183 ( \5166 , \4843 , \4847 );
xor \U$4184 ( \5167 , \5166 , \4852 );
and \U$4185 ( \5168 , \5165 , \5167 );
xor \U$4186 ( \5169 , \4914 , \4918 );
xor \U$4187 ( \5170 , \5169 , \4923 );
and \U$4188 ( \5171 , \5167 , \5170 );
and \U$4189 ( \5172 , \5165 , \5170 );
or \U$4190 ( \5173 , \5168 , \5171 , \5172 );
xor \U$4191 ( \5174 , \4956 , \4958 );
xor \U$4192 ( \5175 , \5174 , \4961 );
and \U$4193 ( \5176 , \5173 , \5175 );
xor \U$4194 ( \5177 , \4966 , \4968 );
and \U$4195 ( \5178 , \5175 , \5177 );
and \U$4196 ( \5179 , \5173 , \5177 );
or \U$4197 ( \5180 , \5176 , \5178 , \5179 );
and \U$4198 ( \5181 , \5162 , \5180 );
and \U$4199 ( \5182 , \5152 , \5180 );
or \U$4200 ( \5183 , \5163 , \5181 , \5182 );
xor \U$4201 ( \5184 , \4715 , \4731 );
xor \U$4202 ( \5185 , \5184 , \4748 );
xor \U$4203 ( \5186 , \4964 , \4969 );
xor \U$4204 ( \5187 , \5186 , \4972 );
and \U$4205 ( \5188 , \5185 , \5187 );
xor \U$4206 ( \5189 , \4978 , \4980 );
xor \U$4207 ( \5190 , \5189 , \4983 );
and \U$4208 ( \5191 , \5187 , \5190 );
and \U$4209 ( \5192 , \5185 , \5190 );
or \U$4210 ( \5193 , \5188 , \5191 , \5192 );
and \U$4211 ( \5194 , \5183 , \5193 );
xor \U$4212 ( \5195 , \4764 , \4774 );
xor \U$4213 ( \5196 , \5195 , \4777 );
and \U$4214 ( \5197 , \5193 , \5196 );
and \U$4215 ( \5198 , \5183 , \5196 );
or \U$4216 ( \5199 , \5194 , \5197 , \5198 );
xor \U$4217 ( \5200 , \4678 , \4695 );
xor \U$4218 ( \5201 , \5200 , \4751 );
xor \U$4219 ( \5202 , \4954 , \4975 );
xor \U$4220 ( \5203 , \5202 , \4986 );
and \U$4221 ( \5204 , \5201 , \5203 );
xor \U$4222 ( \5205 , \4991 , \4993 );
xor \U$4223 ( \5206 , \5205 , \4996 );
and \U$4224 ( \5207 , \5203 , \5206 );
and \U$4225 ( \5208 , \5201 , \5206 );
or \U$4226 ( \5209 , \5204 , \5207 , \5208 );
and \U$4227 ( \5210 , \5199 , \5209 );
xor \U$4228 ( \5211 , \4754 , \4780 );
xor \U$4229 ( \5212 , \5211 , \4790 );
and \U$4230 ( \5213 , \5209 , \5212 );
and \U$4231 ( \5214 , \5199 , \5212 );
or \U$4232 ( \5215 , \5210 , \5213 , \5214 );
xor \U$4233 ( \5216 , \5005 , \5007 );
xor \U$4234 ( \5217 , \5216 , \5010 );
and \U$4235 ( \5218 , \5215 , \5217 );
and \U$4236 ( \5219 , \5019 , \5218 );
xor \U$4237 ( \5220 , \5019 , \5218 );
xor \U$4238 ( \5221 , \5215 , \5217 );
and \U$4239 ( \5222 , \1377 , \3264 );
and \U$4240 ( \5223 , \1349 , \3262 );
nor \U$4241 ( \5224 , \5222 , \5223 );
xnor \U$4242 ( \5225 , \5224 , \3122 );
and \U$4243 ( \5226 , \1531 , \2968 );
and \U$4244 ( \5227 , \1457 , \2966 );
nor \U$4245 ( \5228 , \5226 , \5227 );
xnor \U$4246 ( \5229 , \5228 , \2831 );
and \U$4247 ( \5230 , \5225 , \5229 );
and \U$4248 ( \5231 , \1656 , \2762 );
and \U$4249 ( \5232 , \1593 , \2760 );
nor \U$4250 ( \5233 , \5231 , \5232 );
xnor \U$4251 ( \5234 , \5233 , \2610 );
and \U$4252 ( \5235 , \5229 , \5234 );
and \U$4253 ( \5236 , \5225 , \5234 );
or \U$4254 ( \5237 , \5230 , \5235 , \5236 );
buf \U$4255 ( \5238 , RIc0d89b0_42);
buf \U$4256 ( \5239 , RIc0d8a28_43);
and \U$4257 ( \5240 , \5238 , \5239 );
not \U$4258 ( \5241 , \5240 );
and \U$4259 ( \5242 , \4877 , \5241 );
not \U$4260 ( \5243 , \5242 );
and \U$4261 ( \5244 , \998 , \5023 );
and \U$4262 ( \5245 , \984 , \5021 );
nor \U$4263 ( \5246 , \5244 , \5245 );
xnor \U$4264 ( \5247 , \5246 , \4880 );
and \U$4265 ( \5248 , \5243 , \5247 );
and \U$4266 ( \5249 , \1037 , \4700 );
and \U$4267 ( \5250 , \1016 , \4698 );
nor \U$4268 ( \5251 , \5249 , \5250 );
xnor \U$4269 ( \5252 , \5251 , \4454 );
and \U$4270 ( \5253 , \5247 , \5252 );
and \U$4271 ( \5254 , \5243 , \5252 );
or \U$4272 ( \5255 , \5248 , \5253 , \5254 );
and \U$4273 ( \5256 , \5237 , \5255 );
and \U$4274 ( \5257 , \1093 , \4305 );
and \U$4275 ( \5258 , \1085 , \4303 );
nor \U$4276 ( \5259 , \5257 , \5258 );
xnor \U$4277 ( \5260 , \5259 , \4118 );
and \U$4278 ( \5261 , \1167 , \3992 );
and \U$4279 ( \5262 , \1162 , \3990 );
nor \U$4280 ( \5263 , \5261 , \5262 );
xnor \U$4281 ( \5264 , \5263 , \3787 );
and \U$4282 ( \5265 , \5260 , \5264 );
and \U$4283 ( \5266 , \1272 , \3586 );
and \U$4284 ( \5267 , \1221 , \3584 );
nor \U$4285 ( \5268 , \5266 , \5267 );
xnor \U$4286 ( \5269 , \5268 , \3437 );
and \U$4287 ( \5270 , \5264 , \5269 );
and \U$4288 ( \5271 , \5260 , \5269 );
or \U$4289 ( \5272 , \5265 , \5270 , \5271 );
and \U$4290 ( \5273 , \5255 , \5272 );
and \U$4291 ( \5274 , \5237 , \5272 );
or \U$4292 ( \5275 , \5256 , \5273 , \5274 );
and \U$4293 ( \5276 , \3334 , \1360 );
and \U$4294 ( \5277 , \3309 , \1358 );
nor \U$4295 ( \5278 , \5276 , \5277 );
xnor \U$4296 ( \5279 , \5278 , \1317 );
and \U$4297 ( \5280 , \3675 , \1247 );
and \U$4298 ( \5281 , \3508 , \1245 );
nor \U$4299 ( \5282 , \5280 , \5281 );
xnor \U$4300 ( \5283 , \5282 , \1198 );
and \U$4301 ( \5284 , \5279 , \5283 );
and \U$4302 ( \5285 , \3932 , \1146 );
and \U$4303 ( \5286 , \3813 , \1144 );
nor \U$4304 ( \5287 , \5285 , \5286 );
xnor \U$4305 ( \5288 , \5287 , \1105 );
and \U$4306 ( \5289 , \5283 , \5288 );
and \U$4307 ( \5290 , \5279 , \5288 );
or \U$4308 ( \5291 , \5284 , \5289 , \5290 );
and \U$4309 ( \5292 , \1942 , \2494 );
and \U$4310 ( \5293 , \1854 , \2492 );
nor \U$4311 ( \5294 , \5292 , \5293 );
xnor \U$4312 ( \5295 , \5294 , \2338 );
and \U$4313 ( \5296 , \2052 , \2222 );
and \U$4314 ( \5297 , \2047 , \2220 );
nor \U$4315 ( \5298 , \5296 , \5297 );
xnor \U$4316 ( \5299 , \5298 , \2109 );
and \U$4317 ( \5300 , \5295 , \5299 );
and \U$4318 ( \5301 , \2283 , \2028 );
and \U$4319 ( \5302 , \2168 , \2026 );
nor \U$4320 ( \5303 , \5301 , \5302 );
xnor \U$4321 ( \5304 , \5303 , \1892 );
and \U$4322 ( \5305 , \5299 , \5304 );
and \U$4323 ( \5306 , \5295 , \5304 );
or \U$4324 ( \5307 , \5300 , \5305 , \5306 );
and \U$4325 ( \5308 , \5291 , \5307 );
and \U$4326 ( \5309 , \2467 , \1828 );
and \U$4327 ( \5310 , \2459 , \1826 );
nor \U$4328 ( \5311 , \5309 , \5310 );
xnor \U$4329 ( \5312 , \5311 , \1750 );
and \U$4330 ( \5313 , \2715 , \1664 );
and \U$4331 ( \5314 , \2710 , \1662 );
nor \U$4332 ( \5315 , \5313 , \5314 );
xnor \U$4333 ( \5316 , \5315 , \1570 );
and \U$4334 ( \5317 , \5312 , \5316 );
and \U$4335 ( \5318 , \3045 , \1494 );
and \U$4336 ( \5319 , \2901 , \1492 );
nor \U$4337 ( \5320 , \5318 , \5319 );
xnor \U$4338 ( \5321 , \5320 , \1422 );
and \U$4339 ( \5322 , \5316 , \5321 );
and \U$4340 ( \5323 , \5312 , \5321 );
or \U$4341 ( \5324 , \5317 , \5322 , \5323 );
and \U$4342 ( \5325 , \5307 , \5324 );
and \U$4343 ( \5326 , \5291 , \5324 );
or \U$4344 ( \5327 , \5308 , \5325 , \5326 );
and \U$4345 ( \5328 , \5275 , \5327 );
and \U$4346 ( \5329 , \4557 , \1076 );
and \U$4347 ( \5330 , \4349 , \1074 );
nor \U$4348 ( \5331 , \5329 , \5330 );
xnor \U$4349 ( \5332 , \5331 , \1046 );
and \U$4350 ( \5333 , \4684 , \1028 );
and \U$4351 ( \5334 , \4679 , \1026 );
nor \U$4352 ( \5335 , \5333 , \5334 );
xnor \U$4353 ( \5336 , \5335 , \1009 );
and \U$4354 ( \5337 , \5332 , \5336 );
and \U$4355 ( \5338 , \5137 , \991 );
and \U$4356 ( \5339 , \4940 , \989 );
nor \U$4357 ( \5340 , \5338 , \5339 );
xnor \U$4358 ( \5341 , \5340 , \996 );
and \U$4359 ( \5342 , \5336 , \5341 );
and \U$4360 ( \5343 , \5332 , \5341 );
or \U$4361 ( \5344 , \5337 , \5342 , \5343 );
xor \U$4362 ( \5345 , \5131 , \5135 );
xor \U$4363 ( \5346 , \5345 , \5138 );
or \U$4364 ( \5347 , \5344 , \5346 );
and \U$4365 ( \5348 , \5327 , \5347 );
and \U$4366 ( \5349 , \5275 , \5347 );
or \U$4367 ( \5350 , \5328 , \5348 , \5349 );
xor \U$4368 ( \5351 , \5078 , \5082 );
xor \U$4369 ( \5352 , \5351 , \5087 );
xor \U$4370 ( \5353 , \5094 , \5098 );
xor \U$4371 ( \5354 , \5353 , \5103 );
and \U$4372 ( \5355 , \5352 , \5354 );
xor \U$4373 ( \5356 , \5111 , \5115 );
xor \U$4374 ( \5357 , \5356 , \5120 );
and \U$4375 ( \5358 , \5354 , \5357 );
and \U$4376 ( \5359 , \5352 , \5357 );
or \U$4377 ( \5360 , \5355 , \5358 , \5359 );
xor \U$4378 ( \5361 , \5026 , \5030 );
xor \U$4379 ( \5362 , \5361 , \5035 );
xor \U$4380 ( \5363 , \5042 , \5046 );
xor \U$4381 ( \5364 , \5363 , \5051 );
and \U$4382 ( \5365 , \5362 , \5364 );
xor \U$4383 ( \5366 , \5059 , \5063 );
xor \U$4384 ( \5367 , \5366 , \5068 );
and \U$4385 ( \5368 , \5364 , \5367 );
and \U$4386 ( \5369 , \5362 , \5367 );
or \U$4387 ( \5370 , \5365 , \5368 , \5369 );
and \U$4388 ( \5371 , \5360 , \5370 );
xor \U$4389 ( \5372 , \4897 , \4901 );
xor \U$4390 ( \5373 , \5372 , \4906 );
and \U$4391 ( \5374 , \5370 , \5373 );
and \U$4392 ( \5375 , \5360 , \5373 );
or \U$4393 ( \5376 , \5371 , \5374 , \5375 );
and \U$4394 ( \5377 , \5350 , \5376 );
xor \U$4395 ( \5378 , \4881 , \4885 );
xor \U$4396 ( \5379 , \5378 , \4890 );
xor \U$4397 ( \5380 , \5165 , \5167 );
xor \U$4398 ( \5381 , \5380 , \5170 );
and \U$4399 ( \5382 , \5379 , \5381 );
xor \U$4400 ( \5383 , \5141 , \5143 );
xor \U$4401 ( \5384 , \5383 , \5146 );
and \U$4402 ( \5385 , \5381 , \5384 );
and \U$4403 ( \5386 , \5379 , \5384 );
or \U$4404 ( \5387 , \5382 , \5385 , \5386 );
and \U$4405 ( \5388 , \5376 , \5387 );
and \U$4406 ( \5389 , \5350 , \5387 );
or \U$4407 ( \5390 , \5377 , \5388 , \5389 );
xor \U$4408 ( \5391 , \5074 , \5126 );
xor \U$4409 ( \5392 , \5391 , \5149 );
xor \U$4410 ( \5393 , \5154 , \5156 );
xor \U$4411 ( \5394 , \5393 , \5159 );
and \U$4412 ( \5395 , \5392 , \5394 );
xor \U$4413 ( \5396 , \5173 , \5175 );
xor \U$4414 ( \5397 , \5396 , \5177 );
and \U$4415 ( \5398 , \5394 , \5397 );
and \U$4416 ( \5399 , \5392 , \5397 );
or \U$4417 ( \5400 , \5395 , \5398 , \5399 );
and \U$4418 ( \5401 , \5390 , \5400 );
xor \U$4419 ( \5402 , \4875 , \4929 );
xor \U$4420 ( \5403 , \5402 , \4951 );
and \U$4421 ( \5404 , \5400 , \5403 );
and \U$4422 ( \5405 , \5390 , \5403 );
or \U$4423 ( \5406 , \5401 , \5404 , \5405 );
xor \U$4424 ( \5407 , \5152 , \5162 );
xor \U$4425 ( \5408 , \5407 , \5180 );
xor \U$4426 ( \5409 , \5185 , \5187 );
xor \U$4427 ( \5410 , \5409 , \5190 );
and \U$4428 ( \5411 , \5408 , \5410 );
and \U$4429 ( \5412 , \5406 , \5411 );
xor \U$4430 ( \5413 , \5201 , \5203 );
xor \U$4431 ( \5414 , \5413 , \5206 );
and \U$4432 ( \5415 , \5411 , \5414 );
and \U$4433 ( \5416 , \5406 , \5414 );
or \U$4434 ( \5417 , \5412 , \5415 , \5416 );
xor \U$4435 ( \5418 , \5199 , \5209 );
xor \U$4436 ( \5419 , \5418 , \5212 );
and \U$4437 ( \5420 , \5417 , \5419 );
xor \U$4438 ( \5421 , \4989 , \4999 );
xor \U$4439 ( \5422 , \5421 , \5002 );
and \U$4440 ( \5423 , \5419 , \5422 );
and \U$4441 ( \5424 , \5417 , \5422 );
or \U$4442 ( \5425 , \5420 , \5423 , \5424 );
and \U$4443 ( \5426 , \5221 , \5425 );
xor \U$4444 ( \5427 , \5221 , \5425 );
xor \U$4445 ( \5428 , \5417 , \5419 );
xor \U$4446 ( \5429 , \5428 , \5422 );
and \U$4447 ( \5430 , \4679 , \1076 );
and \U$4448 ( \5431 , \4557 , \1074 );
nor \U$4449 ( \5432 , \5430 , \5431 );
xnor \U$4450 ( \5433 , \5432 , \1046 );
and \U$4451 ( \5434 , \4940 , \1028 );
and \U$4452 ( \5435 , \4684 , \1026 );
nor \U$4453 ( \5436 , \5434 , \5435 );
xnor \U$4454 ( \5437 , \5436 , \1009 );
and \U$4455 ( \5438 , \5433 , \5437 );
buf \U$4456 ( \5439 , RIc0da738_105);
and \U$4457 ( \5440 , \5439 , \991 );
and \U$4458 ( \5441 , \5137 , \989 );
nor \U$4459 ( \5442 , \5440 , \5441 );
xnor \U$4460 ( \5443 , \5442 , \996 );
and \U$4461 ( \5444 , \5437 , \5443 );
and \U$4462 ( \5445 , \5433 , \5443 );
or \U$4463 ( \5446 , \5438 , \5444 , \5445 );
buf \U$4464 ( \5447 , RIc0da7b0_106);
and \U$4465 ( \5448 , \5447 , \985 );
buf \U$4466 ( \5449 , \5448 );
and \U$4467 ( \5450 , \5446 , \5449 );
and \U$4468 ( \5451 , \5439 , \985 );
and \U$4469 ( \5452 , \5449 , \5451 );
and \U$4470 ( \5453 , \5446 , \5451 );
or \U$4471 ( \5454 , \5450 , \5452 , \5453 );
and \U$4472 ( \5455 , \1457 , \3264 );
and \U$4473 ( \5456 , \1377 , \3262 );
nor \U$4474 ( \5457 , \5455 , \5456 );
xnor \U$4475 ( \5458 , \5457 , \3122 );
and \U$4476 ( \5459 , \1593 , \2968 );
and \U$4477 ( \5460 , \1531 , \2966 );
nor \U$4478 ( \5461 , \5459 , \5460 );
xnor \U$4479 ( \5462 , \5461 , \2831 );
and \U$4480 ( \5463 , \5458 , \5462 );
and \U$4481 ( \5464 , \1854 , \2762 );
and \U$4482 ( \5465 , \1656 , \2760 );
nor \U$4483 ( \5466 , \5464 , \5465 );
xnor \U$4484 ( \5467 , \5466 , \2610 );
and \U$4485 ( \5468 , \5462 , \5467 );
and \U$4486 ( \5469 , \5458 , \5467 );
or \U$4487 ( \5470 , \5463 , \5468 , \5469 );
xor \U$4488 ( \5471 , \4877 , \5238 );
xor \U$4489 ( \5472 , \5238 , \5239 );
not \U$4490 ( \5473 , \5472 );
and \U$4491 ( \5474 , \5471 , \5473 );
and \U$4492 ( \5475 , \984 , \5474 );
not \U$4493 ( \5476 , \5475 );
xnor \U$4494 ( \5477 , \5476 , \5242 );
and \U$4495 ( \5478 , \1016 , \5023 );
and \U$4496 ( \5479 , \998 , \5021 );
nor \U$4497 ( \5480 , \5478 , \5479 );
xnor \U$4498 ( \5481 , \5480 , \4880 );
and \U$4499 ( \5482 , \5477 , \5481 );
and \U$4500 ( \5483 , \1085 , \4700 );
and \U$4501 ( \5484 , \1037 , \4698 );
nor \U$4502 ( \5485 , \5483 , \5484 );
xnor \U$4503 ( \5486 , \5485 , \4454 );
and \U$4504 ( \5487 , \5481 , \5486 );
and \U$4505 ( \5488 , \5477 , \5486 );
or \U$4506 ( \5489 , \5482 , \5487 , \5488 );
and \U$4507 ( \5490 , \5470 , \5489 );
and \U$4508 ( \5491 , \1162 , \4305 );
and \U$4509 ( \5492 , \1093 , \4303 );
nor \U$4510 ( \5493 , \5491 , \5492 );
xnor \U$4511 ( \5494 , \5493 , \4118 );
and \U$4512 ( \5495 , \1221 , \3992 );
and \U$4513 ( \5496 , \1167 , \3990 );
nor \U$4514 ( \5497 , \5495 , \5496 );
xnor \U$4515 ( \5498 , \5497 , \3787 );
and \U$4516 ( \5499 , \5494 , \5498 );
and \U$4517 ( \5500 , \1349 , \3586 );
and \U$4518 ( \5501 , \1272 , \3584 );
nor \U$4519 ( \5502 , \5500 , \5501 );
xnor \U$4520 ( \5503 , \5502 , \3437 );
and \U$4521 ( \5504 , \5498 , \5503 );
and \U$4522 ( \5505 , \5494 , \5503 );
or \U$4523 ( \5506 , \5499 , \5504 , \5505 );
and \U$4524 ( \5507 , \5489 , \5506 );
and \U$4525 ( \5508 , \5470 , \5506 );
or \U$4526 ( \5509 , \5490 , \5507 , \5508 );
and \U$4527 ( \5510 , \5454 , \5509 );
and \U$4528 ( \5511 , \3508 , \1360 );
and \U$4529 ( \5512 , \3334 , \1358 );
nor \U$4530 ( \5513 , \5511 , \5512 );
xnor \U$4531 ( \5514 , \5513 , \1317 );
and \U$4532 ( \5515 , \3813 , \1247 );
and \U$4533 ( \5516 , \3675 , \1245 );
nor \U$4534 ( \5517 , \5515 , \5516 );
xnor \U$4535 ( \5518 , \5517 , \1198 );
and \U$4536 ( \5519 , \5514 , \5518 );
and \U$4537 ( \5520 , \4349 , \1146 );
and \U$4538 ( \5521 , \3932 , \1144 );
nor \U$4539 ( \5522 , \5520 , \5521 );
xnor \U$4540 ( \5523 , \5522 , \1105 );
and \U$4541 ( \5524 , \5518 , \5523 );
and \U$4542 ( \5525 , \5514 , \5523 );
or \U$4543 ( \5526 , \5519 , \5524 , \5525 );
and \U$4544 ( \5527 , \2710 , \1828 );
and \U$4545 ( \5528 , \2467 , \1826 );
nor \U$4546 ( \5529 , \5527 , \5528 );
xnor \U$4547 ( \5530 , \5529 , \1750 );
and \U$4548 ( \5531 , \2901 , \1664 );
and \U$4549 ( \5532 , \2715 , \1662 );
nor \U$4550 ( \5533 , \5531 , \5532 );
xnor \U$4551 ( \5534 , \5533 , \1570 );
and \U$4552 ( \5535 , \5530 , \5534 );
and \U$4553 ( \5536 , \3309 , \1494 );
and \U$4554 ( \5537 , \3045 , \1492 );
nor \U$4555 ( \5538 , \5536 , \5537 );
xnor \U$4556 ( \5539 , \5538 , \1422 );
and \U$4557 ( \5540 , \5534 , \5539 );
and \U$4558 ( \5541 , \5530 , \5539 );
or \U$4559 ( \5542 , \5535 , \5540 , \5541 );
and \U$4560 ( \5543 , \5526 , \5542 );
and \U$4561 ( \5544 , \2047 , \2494 );
and \U$4562 ( \5545 , \1942 , \2492 );
nor \U$4563 ( \5546 , \5544 , \5545 );
xnor \U$4564 ( \5547 , \5546 , \2338 );
and \U$4565 ( \5548 , \2168 , \2222 );
and \U$4566 ( \5549 , \2052 , \2220 );
nor \U$4567 ( \5550 , \5548 , \5549 );
xnor \U$4568 ( \5551 , \5550 , \2109 );
and \U$4569 ( \5552 , \5547 , \5551 );
and \U$4570 ( \5553 , \2459 , \2028 );
and \U$4571 ( \5554 , \2283 , \2026 );
nor \U$4572 ( \5555 , \5553 , \5554 );
xnor \U$4573 ( \5556 , \5555 , \1892 );
and \U$4574 ( \5557 , \5551 , \5556 );
and \U$4575 ( \5558 , \5547 , \5556 );
or \U$4576 ( \5559 , \5552 , \5557 , \5558 );
and \U$4577 ( \5560 , \5542 , \5559 );
and \U$4578 ( \5561 , \5526 , \5559 );
or \U$4579 ( \5562 , \5543 , \5560 , \5561 );
and \U$4580 ( \5563 , \5509 , \5562 );
and \U$4581 ( \5564 , \5454 , \5562 );
or \U$4582 ( \5565 , \5510 , \5563 , \5564 );
xor \U$4583 ( \5566 , \5279 , \5283 );
xor \U$4584 ( \5567 , \5566 , \5288 );
xor \U$4585 ( \5568 , \5312 , \5316 );
xor \U$4586 ( \5569 , \5568 , \5321 );
and \U$4587 ( \5570 , \5567 , \5569 );
xor \U$4588 ( \5571 , \5332 , \5336 );
xor \U$4589 ( \5572 , \5571 , \5341 );
and \U$4590 ( \5573 , \5569 , \5572 );
and \U$4591 ( \5574 , \5567 , \5572 );
or \U$4592 ( \5575 , \5570 , \5573 , \5574 );
xor \U$4593 ( \5576 , \5225 , \5229 );
xor \U$4594 ( \5577 , \5576 , \5234 );
xor \U$4595 ( \5578 , \5295 , \5299 );
xor \U$4596 ( \5579 , \5578 , \5304 );
and \U$4597 ( \5580 , \5577 , \5579 );
xor \U$4598 ( \5581 , \5260 , \5264 );
xor \U$4599 ( \5582 , \5581 , \5269 );
and \U$4600 ( \5583 , \5579 , \5582 );
and \U$4601 ( \5584 , \5577 , \5582 );
or \U$4602 ( \5585 , \5580 , \5583 , \5584 );
and \U$4603 ( \5586 , \5575 , \5585 );
xor \U$4604 ( \5587 , \5362 , \5364 );
xor \U$4605 ( \5588 , \5587 , \5367 );
and \U$4606 ( \5589 , \5585 , \5588 );
and \U$4607 ( \5590 , \5575 , \5588 );
or \U$4608 ( \5591 , \5586 , \5589 , \5590 );
and \U$4609 ( \5592 , \5565 , \5591 );
xor \U$4610 ( \5593 , \5291 , \5307 );
xor \U$4611 ( \5594 , \5593 , \5324 );
xor \U$4612 ( \5595 , \5352 , \5354 );
xor \U$4613 ( \5596 , \5595 , \5357 );
and \U$4614 ( \5597 , \5594 , \5596 );
xnor \U$4615 ( \5598 , \5344 , \5346 );
and \U$4616 ( \5599 , \5596 , \5598 );
and \U$4617 ( \5600 , \5594 , \5598 );
or \U$4618 ( \5601 , \5597 , \5599 , \5600 );
and \U$4619 ( \5602 , \5591 , \5601 );
and \U$4620 ( \5603 , \5565 , \5601 );
or \U$4621 ( \5604 , \5592 , \5602 , \5603 );
xor \U$4622 ( \5605 , \5038 , \5054 );
xor \U$4623 ( \5606 , \5605 , \5071 );
xor \U$4624 ( \5607 , \5090 , \5106 );
xor \U$4625 ( \5608 , \5607 , \5123 );
and \U$4626 ( \5609 , \5606 , \5608 );
xor \U$4627 ( \5610 , \5379 , \5381 );
xor \U$4628 ( \5611 , \5610 , \5384 );
and \U$4629 ( \5612 , \5608 , \5611 );
and \U$4630 ( \5613 , \5606 , \5611 );
or \U$4631 ( \5614 , \5609 , \5612 , \5613 );
and \U$4632 ( \5615 , \5604 , \5614 );
xor \U$4633 ( \5616 , \5392 , \5394 );
xor \U$4634 ( \5617 , \5616 , \5397 );
and \U$4635 ( \5618 , \5614 , \5617 );
and \U$4636 ( \5619 , \5604 , \5617 );
or \U$4637 ( \5620 , \5615 , \5618 , \5619 );
xor \U$4638 ( \5621 , \5390 , \5400 );
xor \U$4639 ( \5622 , \5621 , \5403 );
and \U$4640 ( \5623 , \5620 , \5622 );
xor \U$4641 ( \5624 , \5408 , \5410 );
and \U$4642 ( \5625 , \5622 , \5624 );
and \U$4643 ( \5626 , \5620 , \5624 );
or \U$4644 ( \5627 , \5623 , \5625 , \5626 );
xor \U$4645 ( \5628 , \5183 , \5193 );
xor \U$4646 ( \5629 , \5628 , \5196 );
and \U$4647 ( \5630 , \5627 , \5629 );
xor \U$4648 ( \5631 , \5406 , \5411 );
xor \U$4649 ( \5632 , \5631 , \5414 );
and \U$4650 ( \5633 , \5629 , \5632 );
and \U$4651 ( \5634 , \5627 , \5632 );
or \U$4652 ( \5635 , \5630 , \5633 , \5634 );
and \U$4653 ( \5636 , \5429 , \5635 );
xor \U$4654 ( \5637 , \5429 , \5635 );
xor \U$4655 ( \5638 , \5627 , \5629 );
xor \U$4656 ( \5639 , \5638 , \5632 );
and \U$4657 ( \5640 , \1377 , \3586 );
and \U$4658 ( \5641 , \1349 , \3584 );
nor \U$4659 ( \5642 , \5640 , \5641 );
xnor \U$4660 ( \5643 , \5642 , \3437 );
and \U$4661 ( \5644 , \1531 , \3264 );
and \U$4662 ( \5645 , \1457 , \3262 );
nor \U$4663 ( \5646 , \5644 , \5645 );
xnor \U$4664 ( \5647 , \5646 , \3122 );
and \U$4665 ( \5648 , \5643 , \5647 );
and \U$4666 ( \5649 , \1656 , \2968 );
and \U$4667 ( \5650 , \1593 , \2966 );
nor \U$4668 ( \5651 , \5649 , \5650 );
xnor \U$4669 ( \5652 , \5651 , \2831 );
and \U$4670 ( \5653 , \5647 , \5652 );
and \U$4671 ( \5654 , \5643 , \5652 );
or \U$4672 ( \5655 , \5648 , \5653 , \5654 );
buf \U$4673 ( \5656 , RIc0d8aa0_44);
buf \U$4674 ( \5657 , RIc0d8b18_45);
and \U$4675 ( \5658 , \5656 , \5657 );
not \U$4676 ( \5659 , \5658 );
and \U$4677 ( \5660 , \5239 , \5659 );
not \U$4678 ( \5661 , \5660 );
and \U$4679 ( \5662 , \998 , \5474 );
and \U$4680 ( \5663 , \984 , \5472 );
nor \U$4681 ( \5664 , \5662 , \5663 );
xnor \U$4682 ( \5665 , \5664 , \5242 );
and \U$4683 ( \5666 , \5661 , \5665 );
and \U$4684 ( \5667 , \1037 , \5023 );
and \U$4685 ( \5668 , \1016 , \5021 );
nor \U$4686 ( \5669 , \5667 , \5668 );
xnor \U$4687 ( \5670 , \5669 , \4880 );
and \U$4688 ( \5671 , \5665 , \5670 );
and \U$4689 ( \5672 , \5661 , \5670 );
or \U$4690 ( \5673 , \5666 , \5671 , \5672 );
and \U$4691 ( \5674 , \5655 , \5673 );
and \U$4692 ( \5675 , \1093 , \4700 );
and \U$4693 ( \5676 , \1085 , \4698 );
nor \U$4694 ( \5677 , \5675 , \5676 );
xnor \U$4695 ( \5678 , \5677 , \4454 );
and \U$4696 ( \5679 , \1167 , \4305 );
and \U$4697 ( \5680 , \1162 , \4303 );
nor \U$4698 ( \5681 , \5679 , \5680 );
xnor \U$4699 ( \5682 , \5681 , \4118 );
and \U$4700 ( \5683 , \5678 , \5682 );
and \U$4701 ( \5684 , \1272 , \3992 );
and \U$4702 ( \5685 , \1221 , \3990 );
nor \U$4703 ( \5686 , \5684 , \5685 );
xnor \U$4704 ( \5687 , \5686 , \3787 );
and \U$4705 ( \5688 , \5682 , \5687 );
and \U$4706 ( \5689 , \5678 , \5687 );
or \U$4707 ( \5690 , \5683 , \5688 , \5689 );
and \U$4708 ( \5691 , \5673 , \5690 );
and \U$4709 ( \5692 , \5655 , \5690 );
or \U$4710 ( \5693 , \5674 , \5691 , \5692 );
and \U$4711 ( \5694 , \1942 , \2762 );
and \U$4712 ( \5695 , \1854 , \2760 );
nor \U$4713 ( \5696 , \5694 , \5695 );
xnor \U$4714 ( \5697 , \5696 , \2610 );
and \U$4715 ( \5698 , \2052 , \2494 );
and \U$4716 ( \5699 , \2047 , \2492 );
nor \U$4717 ( \5700 , \5698 , \5699 );
xnor \U$4718 ( \5701 , \5700 , \2338 );
and \U$4719 ( \5702 , \5697 , \5701 );
and \U$4720 ( \5703 , \2283 , \2222 );
and \U$4721 ( \5704 , \2168 , \2220 );
nor \U$4722 ( \5705 , \5703 , \5704 );
xnor \U$4723 ( \5706 , \5705 , \2109 );
and \U$4724 ( \5707 , \5701 , \5706 );
and \U$4725 ( \5708 , \5697 , \5706 );
or \U$4726 ( \5709 , \5702 , \5707 , \5708 );
and \U$4727 ( \5710 , \3334 , \1494 );
and \U$4728 ( \5711 , \3309 , \1492 );
nor \U$4729 ( \5712 , \5710 , \5711 );
xnor \U$4730 ( \5713 , \5712 , \1422 );
and \U$4731 ( \5714 , \3675 , \1360 );
and \U$4732 ( \5715 , \3508 , \1358 );
nor \U$4733 ( \5716 , \5714 , \5715 );
xnor \U$4734 ( \5717 , \5716 , \1317 );
and \U$4735 ( \5718 , \5713 , \5717 );
and \U$4736 ( \5719 , \3932 , \1247 );
and \U$4737 ( \5720 , \3813 , \1245 );
nor \U$4738 ( \5721 , \5719 , \5720 );
xnor \U$4739 ( \5722 , \5721 , \1198 );
and \U$4740 ( \5723 , \5717 , \5722 );
and \U$4741 ( \5724 , \5713 , \5722 );
or \U$4742 ( \5725 , \5718 , \5723 , \5724 );
and \U$4743 ( \5726 , \5709 , \5725 );
and \U$4744 ( \5727 , \2467 , \2028 );
and \U$4745 ( \5728 , \2459 , \2026 );
nor \U$4746 ( \5729 , \5727 , \5728 );
xnor \U$4747 ( \5730 , \5729 , \1892 );
and \U$4748 ( \5731 , \2715 , \1828 );
and \U$4749 ( \5732 , \2710 , \1826 );
nor \U$4750 ( \5733 , \5731 , \5732 );
xnor \U$4751 ( \5734 , \5733 , \1750 );
and \U$4752 ( \5735 , \5730 , \5734 );
and \U$4753 ( \5736 , \3045 , \1664 );
and \U$4754 ( \5737 , \2901 , \1662 );
nor \U$4755 ( \5738 , \5736 , \5737 );
xnor \U$4756 ( \5739 , \5738 , \1570 );
and \U$4757 ( \5740 , \5734 , \5739 );
and \U$4758 ( \5741 , \5730 , \5739 );
or \U$4759 ( \5742 , \5735 , \5740 , \5741 );
and \U$4760 ( \5743 , \5725 , \5742 );
and \U$4761 ( \5744 , \5709 , \5742 );
or \U$4762 ( \5745 , \5726 , \5743 , \5744 );
and \U$4763 ( \5746 , \5693 , \5745 );
and \U$4764 ( \5747 , \4557 , \1146 );
and \U$4765 ( \5748 , \4349 , \1144 );
nor \U$4766 ( \5749 , \5747 , \5748 );
xnor \U$4767 ( \5750 , \5749 , \1105 );
and \U$4768 ( \5751 , \4684 , \1076 );
and \U$4769 ( \5752 , \4679 , \1074 );
nor \U$4770 ( \5753 , \5751 , \5752 );
xnor \U$4771 ( \5754 , \5753 , \1046 );
and \U$4772 ( \5755 , \5750 , \5754 );
and \U$4773 ( \5756 , \5137 , \1028 );
and \U$4774 ( \5757 , \4940 , \1026 );
nor \U$4775 ( \5758 , \5756 , \5757 );
xnor \U$4776 ( \5759 , \5758 , \1009 );
and \U$4777 ( \5760 , \5754 , \5759 );
and \U$4778 ( \5761 , \5750 , \5759 );
or \U$4779 ( \5762 , \5755 , \5760 , \5761 );
xor \U$4780 ( \5763 , \5433 , \5437 );
xor \U$4781 ( \5764 , \5763 , \5443 );
and \U$4782 ( \5765 , \5762 , \5764 );
not \U$4783 ( \5766 , \5448 );
and \U$4784 ( \5767 , \5764 , \5766 );
and \U$4785 ( \5768 , \5762 , \5766 );
or \U$4786 ( \5769 , \5765 , \5767 , \5768 );
and \U$4787 ( \5770 , \5745 , \5769 );
and \U$4788 ( \5771 , \5693 , \5769 );
or \U$4789 ( \5772 , \5746 , \5770 , \5771 );
xor \U$4790 ( \5773 , \5514 , \5518 );
xor \U$4791 ( \5774 , \5773 , \5523 );
xor \U$4792 ( \5775 , \5530 , \5534 );
xor \U$4793 ( \5776 , \5775 , \5539 );
and \U$4794 ( \5777 , \5774 , \5776 );
xor \U$4795 ( \5778 , \5547 , \5551 );
xor \U$4796 ( \5779 , \5778 , \5556 );
and \U$4797 ( \5780 , \5776 , \5779 );
and \U$4798 ( \5781 , \5774 , \5779 );
or \U$4799 ( \5782 , \5777 , \5780 , \5781 );
xor \U$4800 ( \5783 , \5458 , \5462 );
xor \U$4801 ( \5784 , \5783 , \5467 );
xor \U$4802 ( \5785 , \5477 , \5481 );
xor \U$4803 ( \5786 , \5785 , \5486 );
and \U$4804 ( \5787 , \5784 , \5786 );
xor \U$4805 ( \5788 , \5494 , \5498 );
xor \U$4806 ( \5789 , \5788 , \5503 );
and \U$4807 ( \5790 , \5786 , \5789 );
and \U$4808 ( \5791 , \5784 , \5789 );
or \U$4809 ( \5792 , \5787 , \5790 , \5791 );
and \U$4810 ( \5793 , \5782 , \5792 );
xor \U$4811 ( \5794 , \5243 , \5247 );
xor \U$4812 ( \5795 , \5794 , \5252 );
and \U$4813 ( \5796 , \5792 , \5795 );
and \U$4814 ( \5797 , \5782 , \5795 );
or \U$4815 ( \5798 , \5793 , \5796 , \5797 );
and \U$4816 ( \5799 , \5772 , \5798 );
xor \U$4817 ( \5800 , \5446 , \5449 );
xor \U$4818 ( \5801 , \5800 , \5451 );
xor \U$4819 ( \5802 , \5567 , \5569 );
xor \U$4820 ( \5803 , \5802 , \5572 );
and \U$4821 ( \5804 , \5801 , \5803 );
xor \U$4822 ( \5805 , \5577 , \5579 );
xor \U$4823 ( \5806 , \5805 , \5582 );
and \U$4824 ( \5807 , \5803 , \5806 );
and \U$4825 ( \5808 , \5801 , \5806 );
or \U$4826 ( \5809 , \5804 , \5807 , \5808 );
and \U$4827 ( \5810 , \5798 , \5809 );
and \U$4828 ( \5811 , \5772 , \5809 );
or \U$4829 ( \5812 , \5799 , \5810 , \5811 );
xor \U$4830 ( \5813 , \5237 , \5255 );
xor \U$4831 ( \5814 , \5813 , \5272 );
xor \U$4832 ( \5815 , \5575 , \5585 );
xor \U$4833 ( \5816 , \5815 , \5588 );
and \U$4834 ( \5817 , \5814 , \5816 );
xor \U$4835 ( \5818 , \5594 , \5596 );
xor \U$4836 ( \5819 , \5818 , \5598 );
and \U$4837 ( \5820 , \5816 , \5819 );
and \U$4838 ( \5821 , \5814 , \5819 );
or \U$4839 ( \5822 , \5817 , \5820 , \5821 );
and \U$4840 ( \5823 , \5812 , \5822 );
xor \U$4841 ( \5824 , \5360 , \5370 );
xor \U$4842 ( \5825 , \5824 , \5373 );
and \U$4843 ( \5826 , \5822 , \5825 );
and \U$4844 ( \5827 , \5812 , \5825 );
or \U$4845 ( \5828 , \5823 , \5826 , \5827 );
xor \U$4846 ( \5829 , \5275 , \5327 );
xor \U$4847 ( \5830 , \5829 , \5347 );
xor \U$4848 ( \5831 , \5565 , \5591 );
xor \U$4849 ( \5832 , \5831 , \5601 );
and \U$4850 ( \5833 , \5830 , \5832 );
xor \U$4851 ( \5834 , \5606 , \5608 );
xor \U$4852 ( \5835 , \5834 , \5611 );
and \U$4853 ( \5836 , \5832 , \5835 );
and \U$4854 ( \5837 , \5830 , \5835 );
or \U$4855 ( \5838 , \5833 , \5836 , \5837 );
and \U$4856 ( \5839 , \5828 , \5838 );
xor \U$4857 ( \5840 , \5350 , \5376 );
xor \U$4858 ( \5841 , \5840 , \5387 );
and \U$4859 ( \5842 , \5838 , \5841 );
and \U$4860 ( \5843 , \5828 , \5841 );
or \U$4861 ( \5844 , \5839 , \5842 , \5843 );
xor \U$4862 ( \5845 , \5239 , \5656 );
xor \U$4863 ( \5846 , \5656 , \5657 );
not \U$4864 ( \5847 , \5846 );
and \U$4865 ( \5848 , \5845 , \5847 );
and \U$4866 ( \5849 , \984 , \5848 );
not \U$4867 ( \5850 , \5849 );
xnor \U$4868 ( \5851 , \5850 , \5660 );
and \U$4869 ( \5852 , \1016 , \5474 );
and \U$4870 ( \5853 , \998 , \5472 );
nor \U$4871 ( \5854 , \5852 , \5853 );
xnor \U$4872 ( \5855 , \5854 , \5242 );
and \U$4873 ( \5856 , \5851 , \5855 );
and \U$4874 ( \5857 , \1085 , \5023 );
and \U$4875 ( \5858 , \1037 , \5021 );
nor \U$4876 ( \5859 , \5857 , \5858 );
xnor \U$4877 ( \5860 , \5859 , \4880 );
and \U$4878 ( \5861 , \5855 , \5860 );
and \U$4879 ( \5862 , \5851 , \5860 );
or \U$4880 ( \5863 , \5856 , \5861 , \5862 );
and \U$4881 ( \5864 , \1457 , \3586 );
and \U$4882 ( \5865 , \1377 , \3584 );
nor \U$4883 ( \5866 , \5864 , \5865 );
xnor \U$4884 ( \5867 , \5866 , \3437 );
and \U$4885 ( \5868 , \1593 , \3264 );
and \U$4886 ( \5869 , \1531 , \3262 );
nor \U$4887 ( \5870 , \5868 , \5869 );
xnor \U$4888 ( \5871 , \5870 , \3122 );
and \U$4889 ( \5872 , \5867 , \5871 );
and \U$4890 ( \5873 , \1854 , \2968 );
and \U$4891 ( \5874 , \1656 , \2966 );
nor \U$4892 ( \5875 , \5873 , \5874 );
xnor \U$4893 ( \5876 , \5875 , \2831 );
and \U$4894 ( \5877 , \5871 , \5876 );
and \U$4895 ( \5878 , \5867 , \5876 );
or \U$4896 ( \5879 , \5872 , \5877 , \5878 );
and \U$4897 ( \5880 , \5863 , \5879 );
and \U$4898 ( \5881 , \1162 , \4700 );
and \U$4899 ( \5882 , \1093 , \4698 );
nor \U$4900 ( \5883 , \5881 , \5882 );
xnor \U$4901 ( \5884 , \5883 , \4454 );
and \U$4902 ( \5885 , \1221 , \4305 );
and \U$4903 ( \5886 , \1167 , \4303 );
nor \U$4904 ( \5887 , \5885 , \5886 );
xnor \U$4905 ( \5888 , \5887 , \4118 );
and \U$4906 ( \5889 , \5884 , \5888 );
and \U$4907 ( \5890 , \1349 , \3992 );
and \U$4908 ( \5891 , \1272 , \3990 );
nor \U$4909 ( \5892 , \5890 , \5891 );
xnor \U$4910 ( \5893 , \5892 , \3787 );
and \U$4911 ( \5894 , \5888 , \5893 );
and \U$4912 ( \5895 , \5884 , \5893 );
or \U$4913 ( \5896 , \5889 , \5894 , \5895 );
and \U$4914 ( \5897 , \5879 , \5896 );
and \U$4915 ( \5898 , \5863 , \5896 );
or \U$4916 ( \5899 , \5880 , \5897 , \5898 );
and \U$4917 ( \5900 , \4679 , \1146 );
and \U$4918 ( \5901 , \4557 , \1144 );
nor \U$4919 ( \5902 , \5900 , \5901 );
xnor \U$4920 ( \5903 , \5902 , \1105 );
and \U$4921 ( \5904 , \4940 , \1076 );
and \U$4922 ( \5905 , \4684 , \1074 );
nor \U$4923 ( \5906 , \5904 , \5905 );
xnor \U$4924 ( \5907 , \5906 , \1046 );
and \U$4925 ( \5908 , \5903 , \5907 );
and \U$4926 ( \5909 , \5439 , \1028 );
and \U$4927 ( \5910 , \5137 , \1026 );
nor \U$4928 ( \5911 , \5909 , \5910 );
xnor \U$4929 ( \5912 , \5911 , \1009 );
and \U$4930 ( \5913 , \5907 , \5912 );
and \U$4931 ( \5914 , \5903 , \5912 );
or \U$4932 ( \5915 , \5908 , \5913 , \5914 );
buf \U$4933 ( \5916 , RIc0da828_107);
and \U$4934 ( \5917 , \5916 , \991 );
and \U$4935 ( \5918 , \5447 , \989 );
nor \U$4936 ( \5919 , \5917 , \5918 );
xnor \U$4937 ( \5920 , \5919 , \996 );
buf \U$4938 ( \5921 , RIc0da8a0_108);
and \U$4939 ( \5922 , \5921 , \985 );
or \U$4940 ( \5923 , \5920 , \5922 );
and \U$4941 ( \5924 , \5915 , \5923 );
and \U$4942 ( \5925 , \5447 , \991 );
and \U$4943 ( \5926 , \5439 , \989 );
nor \U$4944 ( \5927 , \5925 , \5926 );
xnor \U$4945 ( \5928 , \5927 , \996 );
and \U$4946 ( \5929 , \5923 , \5928 );
and \U$4947 ( \5930 , \5915 , \5928 );
or \U$4948 ( \5931 , \5924 , \5929 , \5930 );
and \U$4949 ( \5932 , \5899 , \5931 );
and \U$4950 ( \5933 , \2047 , \2762 );
and \U$4951 ( \5934 , \1942 , \2760 );
nor \U$4952 ( \5935 , \5933 , \5934 );
xnor \U$4953 ( \5936 , \5935 , \2610 );
and \U$4954 ( \5937 , \2168 , \2494 );
and \U$4955 ( \5938 , \2052 , \2492 );
nor \U$4956 ( \5939 , \5937 , \5938 );
xnor \U$4957 ( \5940 , \5939 , \2338 );
and \U$4958 ( \5941 , \5936 , \5940 );
and \U$4959 ( \5942 , \2459 , \2222 );
and \U$4960 ( \5943 , \2283 , \2220 );
nor \U$4961 ( \5944 , \5942 , \5943 );
xnor \U$4962 ( \5945 , \5944 , \2109 );
and \U$4963 ( \5946 , \5940 , \5945 );
and \U$4964 ( \5947 , \5936 , \5945 );
or \U$4965 ( \5948 , \5941 , \5946 , \5947 );
and \U$4966 ( \5949 , \2710 , \2028 );
and \U$4967 ( \5950 , \2467 , \2026 );
nor \U$4968 ( \5951 , \5949 , \5950 );
xnor \U$4969 ( \5952 , \5951 , \1892 );
and \U$4970 ( \5953 , \2901 , \1828 );
and \U$4971 ( \5954 , \2715 , \1826 );
nor \U$4972 ( \5955 , \5953 , \5954 );
xnor \U$4973 ( \5956 , \5955 , \1750 );
and \U$4974 ( \5957 , \5952 , \5956 );
and \U$4975 ( \5958 , \3309 , \1664 );
and \U$4976 ( \5959 , \3045 , \1662 );
nor \U$4977 ( \5960 , \5958 , \5959 );
xnor \U$4978 ( \5961 , \5960 , \1570 );
and \U$4979 ( \5962 , \5956 , \5961 );
and \U$4980 ( \5963 , \5952 , \5961 );
or \U$4981 ( \5964 , \5957 , \5962 , \5963 );
and \U$4982 ( \5965 , \5948 , \5964 );
and \U$4983 ( \5966 , \3508 , \1494 );
and \U$4984 ( \5967 , \3334 , \1492 );
nor \U$4985 ( \5968 , \5966 , \5967 );
xnor \U$4986 ( \5969 , \5968 , \1422 );
and \U$4987 ( \5970 , \3813 , \1360 );
and \U$4988 ( \5971 , \3675 , \1358 );
nor \U$4989 ( \5972 , \5970 , \5971 );
xnor \U$4990 ( \5973 , \5972 , \1317 );
and \U$4991 ( \5974 , \5969 , \5973 );
and \U$4992 ( \5975 , \4349 , \1247 );
and \U$4993 ( \5976 , \3932 , \1245 );
nor \U$4994 ( \5977 , \5975 , \5976 );
xnor \U$4995 ( \5978 , \5977 , \1198 );
and \U$4996 ( \5979 , \5973 , \5978 );
and \U$4997 ( \5980 , \5969 , \5978 );
or \U$4998 ( \5981 , \5974 , \5979 , \5980 );
and \U$4999 ( \5982 , \5964 , \5981 );
and \U$5000 ( \5983 , \5948 , \5981 );
or \U$5001 ( \5984 , \5965 , \5982 , \5983 );
and \U$5002 ( \5985 , \5931 , \5984 );
and \U$5003 ( \5986 , \5899 , \5984 );
or \U$5004 ( \5987 , \5932 , \5985 , \5986 );
and \U$5005 ( \5988 , \5916 , \985 );
xor \U$5006 ( \5989 , \5750 , \5754 );
xor \U$5007 ( \5990 , \5989 , \5759 );
and \U$5008 ( \5991 , \5988 , \5990 );
xor \U$5009 ( \5992 , \5713 , \5717 );
xor \U$5010 ( \5993 , \5992 , \5722 );
and \U$5011 ( \5994 , \5990 , \5993 );
and \U$5012 ( \5995 , \5988 , \5993 );
or \U$5013 ( \5996 , \5991 , \5994 , \5995 );
xor \U$5014 ( \5997 , \5697 , \5701 );
xor \U$5015 ( \5998 , \5997 , \5706 );
xor \U$5016 ( \5999 , \5643 , \5647 );
xor \U$5017 ( \6000 , \5999 , \5652 );
and \U$5018 ( \6001 , \5998 , \6000 );
xor \U$5019 ( \6002 , \5730 , \5734 );
xor \U$5020 ( \6003 , \6002 , \5739 );
and \U$5021 ( \6004 , \6000 , \6003 );
and \U$5022 ( \6005 , \5998 , \6003 );
or \U$5023 ( \6006 , \6001 , \6004 , \6005 );
and \U$5024 ( \6007 , \5996 , \6006 );
xor \U$5025 ( \6008 , \5784 , \5786 );
xor \U$5026 ( \6009 , \6008 , \5789 );
and \U$5027 ( \6010 , \6006 , \6009 );
and \U$5028 ( \6011 , \5996 , \6009 );
or \U$5029 ( \6012 , \6007 , \6010 , \6011 );
and \U$5030 ( \6013 , \5987 , \6012 );
xor \U$5031 ( \6014 , \5709 , \5725 );
xor \U$5032 ( \6015 , \6014 , \5742 );
xor \U$5033 ( \6016 , \5774 , \5776 );
xor \U$5034 ( \6017 , \6016 , \5779 );
and \U$5035 ( \6018 , \6015 , \6017 );
xor \U$5036 ( \6019 , \5762 , \5764 );
xor \U$5037 ( \6020 , \6019 , \5766 );
and \U$5038 ( \6021 , \6017 , \6020 );
and \U$5039 ( \6022 , \6015 , \6020 );
or \U$5040 ( \6023 , \6018 , \6021 , \6022 );
and \U$5041 ( \6024 , \6012 , \6023 );
and \U$5042 ( \6025 , \5987 , \6023 );
or \U$5043 ( \6026 , \6013 , \6024 , \6025 );
xor \U$5044 ( \6027 , \5470 , \5489 );
xor \U$5045 ( \6028 , \6027 , \5506 );
xor \U$5046 ( \6029 , \5526 , \5542 );
xor \U$5047 ( \6030 , \6029 , \5559 );
and \U$5048 ( \6031 , \6028 , \6030 );
xor \U$5049 ( \6032 , \5801 , \5803 );
xor \U$5050 ( \6033 , \6032 , \5806 );
and \U$5051 ( \6034 , \6030 , \6033 );
and \U$5052 ( \6035 , \6028 , \6033 );
or \U$5053 ( \6036 , \6031 , \6034 , \6035 );
and \U$5054 ( \6037 , \6026 , \6036 );
xor \U$5055 ( \6038 , \5454 , \5509 );
xor \U$5056 ( \6039 , \6038 , \5562 );
and \U$5057 ( \6040 , \6036 , \6039 );
and \U$5058 ( \6041 , \6026 , \6039 );
or \U$5059 ( \6042 , \6037 , \6040 , \6041 );
xor \U$5060 ( \6043 , \5812 , \5822 );
xor \U$5061 ( \6044 , \6043 , \5825 );
and \U$5062 ( \6045 , \6042 , \6044 );
xor \U$5063 ( \6046 , \5830 , \5832 );
xor \U$5064 ( \6047 , \6046 , \5835 );
and \U$5065 ( \6048 , \6044 , \6047 );
and \U$5066 ( \6049 , \6042 , \6047 );
or \U$5067 ( \6050 , \6045 , \6048 , \6049 );
xor \U$5068 ( \6051 , \5828 , \5838 );
xor \U$5069 ( \6052 , \6051 , \5841 );
and \U$5070 ( \6053 , \6050 , \6052 );
xor \U$5071 ( \6054 , \5604 , \5614 );
xor \U$5072 ( \6055 , \6054 , \5617 );
and \U$5073 ( \6056 , \6052 , \6055 );
and \U$5074 ( \6057 , \6050 , \6055 );
or \U$5075 ( \6058 , \6053 , \6056 , \6057 );
and \U$5076 ( \6059 , \5844 , \6058 );
xor \U$5077 ( \6060 , \5620 , \5622 );
xor \U$5078 ( \6061 , \6060 , \5624 );
and \U$5079 ( \6062 , \6058 , \6061 );
and \U$5080 ( \6063 , \5844 , \6061 );
or \U$5081 ( \6064 , \6059 , \6062 , \6063 );
and \U$5082 ( \6065 , \5639 , \6064 );
xor \U$5083 ( \6066 , \5639 , \6064 );
xor \U$5084 ( \6067 , \5844 , \6058 );
xor \U$5085 ( \6068 , \6067 , \6061 );
buf \U$5086 ( \6069 , RIc0d8b90_46);
buf \U$5087 ( \6070 , RIc0d8c08_47);
and \U$5088 ( \6071 , \6069 , \6070 );
not \U$5089 ( \6072 , \6071 );
and \U$5090 ( \6073 , \5657 , \6072 );
not \U$5091 ( \6074 , \6073 );
and \U$5092 ( \6075 , \998 , \5848 );
and \U$5093 ( \6076 , \984 , \5846 );
nor \U$5094 ( \6077 , \6075 , \6076 );
xnor \U$5095 ( \6078 , \6077 , \5660 );
and \U$5096 ( \6079 , \6074 , \6078 );
and \U$5097 ( \6080 , \1037 , \5474 );
and \U$5098 ( \6081 , \1016 , \5472 );
nor \U$5099 ( \6082 , \6080 , \6081 );
xnor \U$5100 ( \6083 , \6082 , \5242 );
and \U$5101 ( \6084 , \6078 , \6083 );
and \U$5102 ( \6085 , \6074 , \6083 );
or \U$5103 ( \6086 , \6079 , \6084 , \6085 );
and \U$5104 ( \6087 , \1093 , \5023 );
and \U$5105 ( \6088 , \1085 , \5021 );
nor \U$5106 ( \6089 , \6087 , \6088 );
xnor \U$5107 ( \6090 , \6089 , \4880 );
and \U$5108 ( \6091 , \1167 , \4700 );
and \U$5109 ( \6092 , \1162 , \4698 );
nor \U$5110 ( \6093 , \6091 , \6092 );
xnor \U$5111 ( \6094 , \6093 , \4454 );
and \U$5112 ( \6095 , \6090 , \6094 );
and \U$5113 ( \6096 , \1272 , \4305 );
and \U$5114 ( \6097 , \1221 , \4303 );
nor \U$5115 ( \6098 , \6096 , \6097 );
xnor \U$5116 ( \6099 , \6098 , \4118 );
and \U$5117 ( \6100 , \6094 , \6099 );
and \U$5118 ( \6101 , \6090 , \6099 );
or \U$5119 ( \6102 , \6095 , \6100 , \6101 );
and \U$5120 ( \6103 , \6086 , \6102 );
and \U$5121 ( \6104 , \1377 , \3992 );
and \U$5122 ( \6105 , \1349 , \3990 );
nor \U$5123 ( \6106 , \6104 , \6105 );
xnor \U$5124 ( \6107 , \6106 , \3787 );
and \U$5125 ( \6108 , \1531 , \3586 );
and \U$5126 ( \6109 , \1457 , \3584 );
nor \U$5127 ( \6110 , \6108 , \6109 );
xnor \U$5128 ( \6111 , \6110 , \3437 );
and \U$5129 ( \6112 , \6107 , \6111 );
and \U$5130 ( \6113 , \1656 , \3264 );
and \U$5131 ( \6114 , \1593 , \3262 );
nor \U$5132 ( \6115 , \6113 , \6114 );
xnor \U$5133 ( \6116 , \6115 , \3122 );
and \U$5134 ( \6117 , \6111 , \6116 );
and \U$5135 ( \6118 , \6107 , \6116 );
or \U$5136 ( \6119 , \6112 , \6117 , \6118 );
and \U$5137 ( \6120 , \6102 , \6119 );
and \U$5138 ( \6121 , \6086 , \6119 );
or \U$5139 ( \6122 , \6103 , \6120 , \6121 );
and \U$5140 ( \6123 , \1942 , \2968 );
and \U$5141 ( \6124 , \1854 , \2966 );
nor \U$5142 ( \6125 , \6123 , \6124 );
xnor \U$5143 ( \6126 , \6125 , \2831 );
and \U$5144 ( \6127 , \2052 , \2762 );
and \U$5145 ( \6128 , \2047 , \2760 );
nor \U$5146 ( \6129 , \6127 , \6128 );
xnor \U$5147 ( \6130 , \6129 , \2610 );
and \U$5148 ( \6131 , \6126 , \6130 );
and \U$5149 ( \6132 , \2283 , \2494 );
and \U$5150 ( \6133 , \2168 , \2492 );
nor \U$5151 ( \6134 , \6132 , \6133 );
xnor \U$5152 ( \6135 , \6134 , \2338 );
and \U$5153 ( \6136 , \6130 , \6135 );
and \U$5154 ( \6137 , \6126 , \6135 );
or \U$5155 ( \6138 , \6131 , \6136 , \6137 );
and \U$5156 ( \6139 , \2467 , \2222 );
and \U$5157 ( \6140 , \2459 , \2220 );
nor \U$5158 ( \6141 , \6139 , \6140 );
xnor \U$5159 ( \6142 , \6141 , \2109 );
and \U$5160 ( \6143 , \2715 , \2028 );
and \U$5161 ( \6144 , \2710 , \2026 );
nor \U$5162 ( \6145 , \6143 , \6144 );
xnor \U$5163 ( \6146 , \6145 , \1892 );
and \U$5164 ( \6147 , \6142 , \6146 );
and \U$5165 ( \6148 , \3045 , \1828 );
and \U$5166 ( \6149 , \2901 , \1826 );
nor \U$5167 ( \6150 , \6148 , \6149 );
xnor \U$5168 ( \6151 , \6150 , \1750 );
and \U$5169 ( \6152 , \6146 , \6151 );
and \U$5170 ( \6153 , \6142 , \6151 );
or \U$5171 ( \6154 , \6147 , \6152 , \6153 );
and \U$5172 ( \6155 , \6138 , \6154 );
and \U$5173 ( \6156 , \3334 , \1664 );
and \U$5174 ( \6157 , \3309 , \1662 );
nor \U$5175 ( \6158 , \6156 , \6157 );
xnor \U$5176 ( \6159 , \6158 , \1570 );
and \U$5177 ( \6160 , \3675 , \1494 );
and \U$5178 ( \6161 , \3508 , \1492 );
nor \U$5179 ( \6162 , \6160 , \6161 );
xnor \U$5180 ( \6163 , \6162 , \1422 );
and \U$5181 ( \6164 , \6159 , \6163 );
and \U$5182 ( \6165 , \3932 , \1360 );
and \U$5183 ( \6166 , \3813 , \1358 );
nor \U$5184 ( \6167 , \6165 , \6166 );
xnor \U$5185 ( \6168 , \6167 , \1317 );
and \U$5186 ( \6169 , \6163 , \6168 );
and \U$5187 ( \6170 , \6159 , \6168 );
or \U$5188 ( \6171 , \6164 , \6169 , \6170 );
and \U$5189 ( \6172 , \6154 , \6171 );
and \U$5190 ( \6173 , \6138 , \6171 );
or \U$5191 ( \6174 , \6155 , \6172 , \6173 );
and \U$5192 ( \6175 , \6122 , \6174 );
and \U$5193 ( \6176 , \5447 , \1028 );
and \U$5194 ( \6177 , \5439 , \1026 );
nor \U$5195 ( \6178 , \6176 , \6177 );
xnor \U$5196 ( \6179 , \6178 , \1009 );
and \U$5197 ( \6180 , \5921 , \991 );
and \U$5198 ( \6181 , \5916 , \989 );
nor \U$5199 ( \6182 , \6180 , \6181 );
xnor \U$5200 ( \6183 , \6182 , \996 );
and \U$5201 ( \6184 , \6179 , \6183 );
buf \U$5202 ( \6185 , RIc0da918_109);
and \U$5203 ( \6186 , \6185 , \985 );
and \U$5204 ( \6187 , \6183 , \6186 );
and \U$5205 ( \6188 , \6179 , \6186 );
or \U$5206 ( \6189 , \6184 , \6187 , \6188 );
and \U$5207 ( \6190 , \4557 , \1247 );
and \U$5208 ( \6191 , \4349 , \1245 );
nor \U$5209 ( \6192 , \6190 , \6191 );
xnor \U$5210 ( \6193 , \6192 , \1198 );
and \U$5211 ( \6194 , \4684 , \1146 );
and \U$5212 ( \6195 , \4679 , \1144 );
nor \U$5213 ( \6196 , \6194 , \6195 );
xnor \U$5214 ( \6197 , \6196 , \1105 );
and \U$5215 ( \6198 , \6193 , \6197 );
and \U$5216 ( \6199 , \5137 , \1076 );
and \U$5217 ( \6200 , \4940 , \1074 );
nor \U$5218 ( \6201 , \6199 , \6200 );
xnor \U$5219 ( \6202 , \6201 , \1046 );
and \U$5220 ( \6203 , \6197 , \6202 );
and \U$5221 ( \6204 , \6193 , \6202 );
or \U$5222 ( \6205 , \6198 , \6203 , \6204 );
and \U$5223 ( \6206 , \6189 , \6205 );
xnor \U$5224 ( \6207 , \5920 , \5922 );
and \U$5225 ( \6208 , \6205 , \6207 );
and \U$5226 ( \6209 , \6189 , \6207 );
or \U$5227 ( \6210 , \6206 , \6208 , \6209 );
and \U$5228 ( \6211 , \6174 , \6210 );
and \U$5229 ( \6212 , \6122 , \6210 );
or \U$5230 ( \6213 , \6175 , \6211 , \6212 );
xor \U$5231 ( \6214 , \5903 , \5907 );
xor \U$5232 ( \6215 , \6214 , \5912 );
xor \U$5233 ( \6216 , \5952 , \5956 );
xor \U$5234 ( \6217 , \6216 , \5961 );
and \U$5235 ( \6218 , \6215 , \6217 );
xor \U$5236 ( \6219 , \5969 , \5973 );
xor \U$5237 ( \6220 , \6219 , \5978 );
and \U$5238 ( \6221 , \6217 , \6220 );
and \U$5239 ( \6222 , \6215 , \6220 );
or \U$5240 ( \6223 , \6218 , \6221 , \6222 );
xor \U$5241 ( \6224 , \5936 , \5940 );
xor \U$5242 ( \6225 , \6224 , \5945 );
xor \U$5243 ( \6226 , \5867 , \5871 );
xor \U$5244 ( \6227 , \6226 , \5876 );
and \U$5245 ( \6228 , \6225 , \6227 );
xor \U$5246 ( \6229 , \5884 , \5888 );
xor \U$5247 ( \6230 , \6229 , \5893 );
and \U$5248 ( \6231 , \6227 , \6230 );
and \U$5249 ( \6232 , \6225 , \6230 );
or \U$5250 ( \6233 , \6228 , \6231 , \6232 );
and \U$5251 ( \6234 , \6223 , \6233 );
xor \U$5252 ( \6235 , \5678 , \5682 );
xor \U$5253 ( \6236 , \6235 , \5687 );
and \U$5254 ( \6237 , \6233 , \6236 );
and \U$5255 ( \6238 , \6223 , \6236 );
or \U$5256 ( \6239 , \6234 , \6237 , \6238 );
and \U$5257 ( \6240 , \6213 , \6239 );
xor \U$5258 ( \6241 , \5661 , \5665 );
xor \U$5259 ( \6242 , \6241 , \5670 );
xor \U$5260 ( \6243 , \5988 , \5990 );
xor \U$5261 ( \6244 , \6243 , \5993 );
and \U$5262 ( \6245 , \6242 , \6244 );
xor \U$5263 ( \6246 , \5998 , \6000 );
xor \U$5264 ( \6247 , \6246 , \6003 );
and \U$5265 ( \6248 , \6244 , \6247 );
and \U$5266 ( \6249 , \6242 , \6247 );
or \U$5267 ( \6250 , \6245 , \6248 , \6249 );
and \U$5268 ( \6251 , \6239 , \6250 );
and \U$5269 ( \6252 , \6213 , \6250 );
or \U$5270 ( \6253 , \6240 , \6251 , \6252 );
xor \U$5271 ( \6254 , \5863 , \5879 );
xor \U$5272 ( \6255 , \6254 , \5896 );
xor \U$5273 ( \6256 , \5915 , \5923 );
xor \U$5274 ( \6257 , \6256 , \5928 );
and \U$5275 ( \6258 , \6255 , \6257 );
xor \U$5276 ( \6259 , \5948 , \5964 );
xor \U$5277 ( \6260 , \6259 , \5981 );
and \U$5278 ( \6261 , \6257 , \6260 );
and \U$5279 ( \6262 , \6255 , \6260 );
or \U$5280 ( \6263 , \6258 , \6261 , \6262 );
xor \U$5281 ( \6264 , \5655 , \5673 );
xor \U$5282 ( \6265 , \6264 , \5690 );
and \U$5283 ( \6266 , \6263 , \6265 );
xor \U$5284 ( \6267 , \6015 , \6017 );
xor \U$5285 ( \6268 , \6267 , \6020 );
and \U$5286 ( \6269 , \6265 , \6268 );
and \U$5287 ( \6270 , \6263 , \6268 );
or \U$5288 ( \6271 , \6266 , \6269 , \6270 );
and \U$5289 ( \6272 , \6253 , \6271 );
xor \U$5290 ( \6273 , \5782 , \5792 );
xor \U$5291 ( \6274 , \6273 , \5795 );
and \U$5292 ( \6275 , \6271 , \6274 );
and \U$5293 ( \6276 , \6253 , \6274 );
or \U$5294 ( \6277 , \6272 , \6275 , \6276 );
xor \U$5295 ( \6278 , \5693 , \5745 );
xor \U$5296 ( \6279 , \6278 , \5769 );
xor \U$5297 ( \6280 , \5987 , \6012 );
xor \U$5298 ( \6281 , \6280 , \6023 );
and \U$5299 ( \6282 , \6279 , \6281 );
xor \U$5300 ( \6283 , \6028 , \6030 );
xor \U$5301 ( \6284 , \6283 , \6033 );
and \U$5302 ( \6285 , \6281 , \6284 );
and \U$5303 ( \6286 , \6279 , \6284 );
or \U$5304 ( \6287 , \6282 , \6285 , \6286 );
and \U$5305 ( \6288 , \6277 , \6287 );
xor \U$5306 ( \6289 , \5814 , \5816 );
xor \U$5307 ( \6290 , \6289 , \5819 );
and \U$5308 ( \6291 , \6287 , \6290 );
and \U$5309 ( \6292 , \6277 , \6290 );
or \U$5310 ( \6293 , \6288 , \6291 , \6292 );
xor \U$5311 ( \6294 , \5772 , \5798 );
xor \U$5312 ( \6295 , \6294 , \5809 );
xor \U$5313 ( \6296 , \6026 , \6036 );
xor \U$5314 ( \6297 , \6296 , \6039 );
and \U$5315 ( \6298 , \6295 , \6297 );
and \U$5316 ( \6299 , \6293 , \6298 );
xor \U$5317 ( \6300 , \6042 , \6044 );
xor \U$5318 ( \6301 , \6300 , \6047 );
and \U$5319 ( \6302 , \6298 , \6301 );
and \U$5320 ( \6303 , \6293 , \6301 );
or \U$5321 ( \6304 , \6299 , \6302 , \6303 );
xor \U$5322 ( \6305 , \6050 , \6052 );
xor \U$5323 ( \6306 , \6305 , \6055 );
and \U$5324 ( \6307 , \6304 , \6306 );
and \U$5325 ( \6308 , \6068 , \6307 );
xor \U$5326 ( \6309 , \6068 , \6307 );
xor \U$5327 ( \6310 , \6304 , \6306 );
xor \U$5328 ( \6311 , \5657 , \6069 );
xor \U$5329 ( \6312 , \6069 , \6070 );
not \U$5330 ( \6313 , \6312 );
and \U$5331 ( \6314 , \6311 , \6313 );
and \U$5332 ( \6315 , \984 , \6314 );
not \U$5333 ( \6316 , \6315 );
xnor \U$5334 ( \6317 , \6316 , \6073 );
and \U$5335 ( \6318 , \1016 , \5848 );
and \U$5336 ( \6319 , \998 , \5846 );
nor \U$5337 ( \6320 , \6318 , \6319 );
xnor \U$5338 ( \6321 , \6320 , \5660 );
and \U$5339 ( \6322 , \6317 , \6321 );
and \U$5340 ( \6323 , \1085 , \5474 );
and \U$5341 ( \6324 , \1037 , \5472 );
nor \U$5342 ( \6325 , \6323 , \6324 );
xnor \U$5343 ( \6326 , \6325 , \5242 );
and \U$5344 ( \6327 , \6321 , \6326 );
and \U$5345 ( \6328 , \6317 , \6326 );
or \U$5346 ( \6329 , \6322 , \6327 , \6328 );
and \U$5347 ( \6330 , \1162 , \5023 );
and \U$5348 ( \6331 , \1093 , \5021 );
nor \U$5349 ( \6332 , \6330 , \6331 );
xnor \U$5350 ( \6333 , \6332 , \4880 );
and \U$5351 ( \6334 , \1221 , \4700 );
and \U$5352 ( \6335 , \1167 , \4698 );
nor \U$5353 ( \6336 , \6334 , \6335 );
xnor \U$5354 ( \6337 , \6336 , \4454 );
and \U$5355 ( \6338 , \6333 , \6337 );
and \U$5356 ( \6339 , \1349 , \4305 );
and \U$5357 ( \6340 , \1272 , \4303 );
nor \U$5358 ( \6341 , \6339 , \6340 );
xnor \U$5359 ( \6342 , \6341 , \4118 );
and \U$5360 ( \6343 , \6337 , \6342 );
and \U$5361 ( \6344 , \6333 , \6342 );
or \U$5362 ( \6345 , \6338 , \6343 , \6344 );
and \U$5363 ( \6346 , \6329 , \6345 );
and \U$5364 ( \6347 , \1457 , \3992 );
and \U$5365 ( \6348 , \1377 , \3990 );
nor \U$5366 ( \6349 , \6347 , \6348 );
xnor \U$5367 ( \6350 , \6349 , \3787 );
and \U$5368 ( \6351 , \1593 , \3586 );
and \U$5369 ( \6352 , \1531 , \3584 );
nor \U$5370 ( \6353 , \6351 , \6352 );
xnor \U$5371 ( \6354 , \6353 , \3437 );
and \U$5372 ( \6355 , \6350 , \6354 );
and \U$5373 ( \6356 , \1854 , \3264 );
and \U$5374 ( \6357 , \1656 , \3262 );
nor \U$5375 ( \6358 , \6356 , \6357 );
xnor \U$5376 ( \6359 , \6358 , \3122 );
and \U$5377 ( \6360 , \6354 , \6359 );
and \U$5378 ( \6361 , \6350 , \6359 );
or \U$5379 ( \6362 , \6355 , \6360 , \6361 );
and \U$5380 ( \6363 , \6345 , \6362 );
and \U$5381 ( \6364 , \6329 , \6362 );
or \U$5382 ( \6365 , \6346 , \6363 , \6364 );
and \U$5383 ( \6366 , \2047 , \2968 );
and \U$5384 ( \6367 , \1942 , \2966 );
nor \U$5385 ( \6368 , \6366 , \6367 );
xnor \U$5386 ( \6369 , \6368 , \2831 );
and \U$5387 ( \6370 , \2168 , \2762 );
and \U$5388 ( \6371 , \2052 , \2760 );
nor \U$5389 ( \6372 , \6370 , \6371 );
xnor \U$5390 ( \6373 , \6372 , \2610 );
and \U$5391 ( \6374 , \6369 , \6373 );
and \U$5392 ( \6375 , \2459 , \2494 );
and \U$5393 ( \6376 , \2283 , \2492 );
nor \U$5394 ( \6377 , \6375 , \6376 );
xnor \U$5395 ( \6378 , \6377 , \2338 );
and \U$5396 ( \6379 , \6373 , \6378 );
and \U$5397 ( \6380 , \6369 , \6378 );
or \U$5398 ( \6381 , \6374 , \6379 , \6380 );
and \U$5399 ( \6382 , \2710 , \2222 );
and \U$5400 ( \6383 , \2467 , \2220 );
nor \U$5401 ( \6384 , \6382 , \6383 );
xnor \U$5402 ( \6385 , \6384 , \2109 );
and \U$5403 ( \6386 , \2901 , \2028 );
and \U$5404 ( \6387 , \2715 , \2026 );
nor \U$5405 ( \6388 , \6386 , \6387 );
xnor \U$5406 ( \6389 , \6388 , \1892 );
and \U$5407 ( \6390 , \6385 , \6389 );
and \U$5408 ( \6391 , \3309 , \1828 );
and \U$5409 ( \6392 , \3045 , \1826 );
nor \U$5410 ( \6393 , \6391 , \6392 );
xnor \U$5411 ( \6394 , \6393 , \1750 );
and \U$5412 ( \6395 , \6389 , \6394 );
and \U$5413 ( \6396 , \6385 , \6394 );
or \U$5414 ( \6397 , \6390 , \6395 , \6396 );
and \U$5415 ( \6398 , \6381 , \6397 );
and \U$5416 ( \6399 , \3508 , \1664 );
and \U$5417 ( \6400 , \3334 , \1662 );
nor \U$5418 ( \6401 , \6399 , \6400 );
xnor \U$5419 ( \6402 , \6401 , \1570 );
and \U$5420 ( \6403 , \3813 , \1494 );
and \U$5421 ( \6404 , \3675 , \1492 );
nor \U$5422 ( \6405 , \6403 , \6404 );
xnor \U$5423 ( \6406 , \6405 , \1422 );
and \U$5424 ( \6407 , \6402 , \6406 );
and \U$5425 ( \6408 , \4349 , \1360 );
and \U$5426 ( \6409 , \3932 , \1358 );
nor \U$5427 ( \6410 , \6408 , \6409 );
xnor \U$5428 ( \6411 , \6410 , \1317 );
and \U$5429 ( \6412 , \6406 , \6411 );
and \U$5430 ( \6413 , \6402 , \6411 );
or \U$5431 ( \6414 , \6407 , \6412 , \6413 );
and \U$5432 ( \6415 , \6397 , \6414 );
and \U$5433 ( \6416 , \6381 , \6414 );
or \U$5434 ( \6417 , \6398 , \6415 , \6416 );
and \U$5435 ( \6418 , \6365 , \6417 );
and \U$5436 ( \6419 , \4679 , \1247 );
and \U$5437 ( \6420 , \4557 , \1245 );
nor \U$5438 ( \6421 , \6419 , \6420 );
xnor \U$5439 ( \6422 , \6421 , \1198 );
and \U$5440 ( \6423 , \4940 , \1146 );
and \U$5441 ( \6424 , \4684 , \1144 );
nor \U$5442 ( \6425 , \6423 , \6424 );
xnor \U$5443 ( \6426 , \6425 , \1105 );
and \U$5444 ( \6427 , \6422 , \6426 );
and \U$5445 ( \6428 , \5439 , \1076 );
and \U$5446 ( \6429 , \5137 , \1074 );
nor \U$5447 ( \6430 , \6428 , \6429 );
xnor \U$5448 ( \6431 , \6430 , \1046 );
and \U$5449 ( \6432 , \6426 , \6431 );
and \U$5450 ( \6433 , \6422 , \6431 );
or \U$5451 ( \6434 , \6427 , \6432 , \6433 );
and \U$5452 ( \6435 , \5916 , \1028 );
and \U$5453 ( \6436 , \5447 , \1026 );
nor \U$5454 ( \6437 , \6435 , \6436 );
xnor \U$5455 ( \6438 , \6437 , \1009 );
and \U$5456 ( \6439 , \6185 , \991 );
and \U$5457 ( \6440 , \5921 , \989 );
nor \U$5458 ( \6441 , \6439 , \6440 );
xnor \U$5459 ( \6442 , \6441 , \996 );
and \U$5460 ( \6443 , \6438 , \6442 );
buf \U$5461 ( \6444 , RIc0da990_110);
and \U$5462 ( \6445 , \6444 , \985 );
and \U$5463 ( \6446 , \6442 , \6445 );
and \U$5464 ( \6447 , \6438 , \6445 );
or \U$5465 ( \6448 , \6443 , \6446 , \6447 );
and \U$5466 ( \6449 , \6434 , \6448 );
xor \U$5467 ( \6450 , \6179 , \6183 );
xor \U$5468 ( \6451 , \6450 , \6186 );
and \U$5469 ( \6452 , \6448 , \6451 );
and \U$5470 ( \6453 , \6434 , \6451 );
or \U$5471 ( \6454 , \6449 , \6452 , \6453 );
and \U$5472 ( \6455 , \6417 , \6454 );
and \U$5473 ( \6456 , \6365 , \6454 );
or \U$5474 ( \6457 , \6418 , \6455 , \6456 );
xor \U$5475 ( \6458 , \6126 , \6130 );
xor \U$5476 ( \6459 , \6458 , \6135 );
xor \U$5477 ( \6460 , \6090 , \6094 );
xor \U$5478 ( \6461 , \6460 , \6099 );
and \U$5479 ( \6462 , \6459 , \6461 );
xor \U$5480 ( \6463 , \6107 , \6111 );
xor \U$5481 ( \6464 , \6463 , \6116 );
and \U$5482 ( \6465 , \6461 , \6464 );
and \U$5483 ( \6466 , \6459 , \6464 );
or \U$5484 ( \6467 , \6462 , \6465 , \6466 );
xor \U$5485 ( \6468 , \6142 , \6146 );
xor \U$5486 ( \6469 , \6468 , \6151 );
xor \U$5487 ( \6470 , \6159 , \6163 );
xor \U$5488 ( \6471 , \6470 , \6168 );
and \U$5489 ( \6472 , \6469 , \6471 );
xor \U$5490 ( \6473 , \6193 , \6197 );
xor \U$5491 ( \6474 , \6473 , \6202 );
and \U$5492 ( \6475 , \6471 , \6474 );
and \U$5493 ( \6476 , \6469 , \6474 );
or \U$5494 ( \6477 , \6472 , \6475 , \6476 );
and \U$5495 ( \6478 , \6467 , \6477 );
xor \U$5496 ( \6479 , \5851 , \5855 );
xor \U$5497 ( \6480 , \6479 , \5860 );
and \U$5498 ( \6481 , \6477 , \6480 );
and \U$5499 ( \6482 , \6467 , \6480 );
or \U$5500 ( \6483 , \6478 , \6481 , \6482 );
and \U$5501 ( \6484 , \6457 , \6483 );
xor \U$5502 ( \6485 , \6215 , \6217 );
xor \U$5503 ( \6486 , \6485 , \6220 );
xor \U$5504 ( \6487 , \6225 , \6227 );
xor \U$5505 ( \6488 , \6487 , \6230 );
and \U$5506 ( \6489 , \6486 , \6488 );
xor \U$5507 ( \6490 , \6189 , \6205 );
xor \U$5508 ( \6491 , \6490 , \6207 );
and \U$5509 ( \6492 , \6488 , \6491 );
and \U$5510 ( \6493 , \6486 , \6491 );
or \U$5511 ( \6494 , \6489 , \6492 , \6493 );
and \U$5512 ( \6495 , \6483 , \6494 );
and \U$5513 ( \6496 , \6457 , \6494 );
or \U$5514 ( \6497 , \6484 , \6495 , \6496 );
xor \U$5515 ( \6498 , \6223 , \6233 );
xor \U$5516 ( \6499 , \6498 , \6236 );
xor \U$5517 ( \6500 , \6255 , \6257 );
xor \U$5518 ( \6501 , \6500 , \6260 );
and \U$5519 ( \6502 , \6499 , \6501 );
xor \U$5520 ( \6503 , \6242 , \6244 );
xor \U$5521 ( \6504 , \6503 , \6247 );
and \U$5522 ( \6505 , \6501 , \6504 );
and \U$5523 ( \6506 , \6499 , \6504 );
or \U$5524 ( \6507 , \6502 , \6505 , \6506 );
and \U$5525 ( \6508 , \6497 , \6507 );
xor \U$5526 ( \6509 , \5996 , \6006 );
xor \U$5527 ( \6510 , \6509 , \6009 );
and \U$5528 ( \6511 , \6507 , \6510 );
and \U$5529 ( \6512 , \6497 , \6510 );
or \U$5530 ( \6513 , \6508 , \6511 , \6512 );
xor \U$5531 ( \6514 , \5899 , \5931 );
xor \U$5532 ( \6515 , \6514 , \5984 );
xor \U$5533 ( \6516 , \6213 , \6239 );
xor \U$5534 ( \6517 , \6516 , \6250 );
and \U$5535 ( \6518 , \6515 , \6517 );
xor \U$5536 ( \6519 , \6263 , \6265 );
xor \U$5537 ( \6520 , \6519 , \6268 );
and \U$5538 ( \6521 , \6517 , \6520 );
and \U$5539 ( \6522 , \6515 , \6520 );
or \U$5540 ( \6523 , \6518 , \6521 , \6522 );
and \U$5541 ( \6524 , \6513 , \6523 );
xor \U$5542 ( \6525 , \6279 , \6281 );
xor \U$5543 ( \6526 , \6525 , \6284 );
and \U$5544 ( \6527 , \6523 , \6526 );
and \U$5545 ( \6528 , \6513 , \6526 );
or \U$5546 ( \6529 , \6524 , \6527 , \6528 );
xor \U$5547 ( \6530 , \6277 , \6287 );
xor \U$5548 ( \6531 , \6530 , \6290 );
and \U$5549 ( \6532 , \6529 , \6531 );
xor \U$5550 ( \6533 , \6295 , \6297 );
and \U$5551 ( \6534 , \6531 , \6533 );
and \U$5552 ( \6535 , \6529 , \6533 );
or \U$5553 ( \6536 , \6532 , \6534 , \6535 );
xor \U$5554 ( \6537 , \6293 , \6298 );
xor \U$5555 ( \6538 , \6537 , \6301 );
and \U$5556 ( \6539 , \6536 , \6538 );
and \U$5557 ( \6540 , \6310 , \6539 );
xor \U$5558 ( \6541 , \6310 , \6539 );
xor \U$5559 ( \6542 , \6536 , \6538 );
and \U$5560 ( \6543 , \1093 , \5474 );
and \U$5561 ( \6544 , \1085 , \5472 );
nor \U$5562 ( \6545 , \6543 , \6544 );
xnor \U$5563 ( \6546 , \6545 , \5242 );
and \U$5564 ( \6547 , \1167 , \5023 );
and \U$5565 ( \6548 , \1162 , \5021 );
nor \U$5566 ( \6549 , \6547 , \6548 );
xnor \U$5567 ( \6550 , \6549 , \4880 );
and \U$5568 ( \6551 , \6546 , \6550 );
and \U$5569 ( \6552 , \1272 , \4700 );
and \U$5570 ( \6553 , \1221 , \4698 );
nor \U$5571 ( \6554 , \6552 , \6553 );
xnor \U$5572 ( \6555 , \6554 , \4454 );
and \U$5573 ( \6556 , \6550 , \6555 );
and \U$5574 ( \6557 , \6546 , \6555 );
or \U$5575 ( \6558 , \6551 , \6556 , \6557 );
buf \U$5576 ( \6559 , RIc0d8c80_48);
buf \U$5577 ( \6560 , RIc0d8cf8_49);
and \U$5578 ( \6561 , \6559 , \6560 );
not \U$5579 ( \6562 , \6561 );
and \U$5580 ( \6563 , \6070 , \6562 );
not \U$5581 ( \6564 , \6563 );
and \U$5582 ( \6565 , \998 , \6314 );
and \U$5583 ( \6566 , \984 , \6312 );
nor \U$5584 ( \6567 , \6565 , \6566 );
xnor \U$5585 ( \6568 , \6567 , \6073 );
and \U$5586 ( \6569 , \6564 , \6568 );
and \U$5587 ( \6570 , \1037 , \5848 );
and \U$5588 ( \6571 , \1016 , \5846 );
nor \U$5589 ( \6572 , \6570 , \6571 );
xnor \U$5590 ( \6573 , \6572 , \5660 );
and \U$5591 ( \6574 , \6568 , \6573 );
and \U$5592 ( \6575 , \6564 , \6573 );
or \U$5593 ( \6576 , \6569 , \6574 , \6575 );
and \U$5594 ( \6577 , \6558 , \6576 );
and \U$5595 ( \6578 , \1377 , \4305 );
and \U$5596 ( \6579 , \1349 , \4303 );
nor \U$5597 ( \6580 , \6578 , \6579 );
xnor \U$5598 ( \6581 , \6580 , \4118 );
and \U$5599 ( \6582 , \1531 , \3992 );
and \U$5600 ( \6583 , \1457 , \3990 );
nor \U$5601 ( \6584 , \6582 , \6583 );
xnor \U$5602 ( \6585 , \6584 , \3787 );
and \U$5603 ( \6586 , \6581 , \6585 );
and \U$5604 ( \6587 , \1656 , \3586 );
and \U$5605 ( \6588 , \1593 , \3584 );
nor \U$5606 ( \6589 , \6587 , \6588 );
xnor \U$5607 ( \6590 , \6589 , \3437 );
and \U$5608 ( \6591 , \6585 , \6590 );
and \U$5609 ( \6592 , \6581 , \6590 );
or \U$5610 ( \6593 , \6586 , \6591 , \6592 );
and \U$5611 ( \6594 , \6576 , \6593 );
and \U$5612 ( \6595 , \6558 , \6593 );
or \U$5613 ( \6596 , \6577 , \6594 , \6595 );
and \U$5614 ( \6597 , \3334 , \1828 );
and \U$5615 ( \6598 , \3309 , \1826 );
nor \U$5616 ( \6599 , \6597 , \6598 );
xnor \U$5617 ( \6600 , \6599 , \1750 );
and \U$5618 ( \6601 , \3675 , \1664 );
and \U$5619 ( \6602 , \3508 , \1662 );
nor \U$5620 ( \6603 , \6601 , \6602 );
xnor \U$5621 ( \6604 , \6603 , \1570 );
and \U$5622 ( \6605 , \6600 , \6604 );
and \U$5623 ( \6606 , \3932 , \1494 );
and \U$5624 ( \6607 , \3813 , \1492 );
nor \U$5625 ( \6608 , \6606 , \6607 );
xnor \U$5626 ( \6609 , \6608 , \1422 );
and \U$5627 ( \6610 , \6604 , \6609 );
and \U$5628 ( \6611 , \6600 , \6609 );
or \U$5629 ( \6612 , \6605 , \6610 , \6611 );
and \U$5630 ( \6613 , \2467 , \2494 );
and \U$5631 ( \6614 , \2459 , \2492 );
nor \U$5632 ( \6615 , \6613 , \6614 );
xnor \U$5633 ( \6616 , \6615 , \2338 );
and \U$5634 ( \6617 , \2715 , \2222 );
and \U$5635 ( \6618 , \2710 , \2220 );
nor \U$5636 ( \6619 , \6617 , \6618 );
xnor \U$5637 ( \6620 , \6619 , \2109 );
and \U$5638 ( \6621 , \6616 , \6620 );
and \U$5639 ( \6622 , \3045 , \2028 );
and \U$5640 ( \6623 , \2901 , \2026 );
nor \U$5641 ( \6624 , \6622 , \6623 );
xnor \U$5642 ( \6625 , \6624 , \1892 );
and \U$5643 ( \6626 , \6620 , \6625 );
and \U$5644 ( \6627 , \6616 , \6625 );
or \U$5645 ( \6628 , \6621 , \6626 , \6627 );
and \U$5646 ( \6629 , \6612 , \6628 );
and \U$5647 ( \6630 , \1942 , \3264 );
and \U$5648 ( \6631 , \1854 , \3262 );
nor \U$5649 ( \6632 , \6630 , \6631 );
xnor \U$5650 ( \6633 , \6632 , \3122 );
and \U$5651 ( \6634 , \2052 , \2968 );
and \U$5652 ( \6635 , \2047 , \2966 );
nor \U$5653 ( \6636 , \6634 , \6635 );
xnor \U$5654 ( \6637 , \6636 , \2831 );
and \U$5655 ( \6638 , \6633 , \6637 );
and \U$5656 ( \6639 , \2283 , \2762 );
and \U$5657 ( \6640 , \2168 , \2760 );
nor \U$5658 ( \6641 , \6639 , \6640 );
xnor \U$5659 ( \6642 , \6641 , \2610 );
and \U$5660 ( \6643 , \6637 , \6642 );
and \U$5661 ( \6644 , \6633 , \6642 );
or \U$5662 ( \6645 , \6638 , \6643 , \6644 );
and \U$5663 ( \6646 , \6628 , \6645 );
and \U$5664 ( \6647 , \6612 , \6645 );
or \U$5665 ( \6648 , \6629 , \6646 , \6647 );
and \U$5666 ( \6649 , \6596 , \6648 );
and \U$5667 ( \6650 , \4557 , \1360 );
and \U$5668 ( \6651 , \4349 , \1358 );
nor \U$5669 ( \6652 , \6650 , \6651 );
xnor \U$5670 ( \6653 , \6652 , \1317 );
and \U$5671 ( \6654 , \4684 , \1247 );
and \U$5672 ( \6655 , \4679 , \1245 );
nor \U$5673 ( \6656 , \6654 , \6655 );
xnor \U$5674 ( \6657 , \6656 , \1198 );
and \U$5675 ( \6658 , \6653 , \6657 );
and \U$5676 ( \6659 , \5137 , \1146 );
and \U$5677 ( \6660 , \4940 , \1144 );
nor \U$5678 ( \6661 , \6659 , \6660 );
xnor \U$5679 ( \6662 , \6661 , \1105 );
and \U$5680 ( \6663 , \6657 , \6662 );
and \U$5681 ( \6664 , \6653 , \6662 );
or \U$5682 ( \6665 , \6658 , \6663 , \6664 );
and \U$5683 ( \6666 , \5447 , \1076 );
and \U$5684 ( \6667 , \5439 , \1074 );
nor \U$5685 ( \6668 , \6666 , \6667 );
xnor \U$5686 ( \6669 , \6668 , \1046 );
and \U$5687 ( \6670 , \5921 , \1028 );
and \U$5688 ( \6671 , \5916 , \1026 );
nor \U$5689 ( \6672 , \6670 , \6671 );
xnor \U$5690 ( \6673 , \6672 , \1009 );
and \U$5691 ( \6674 , \6669 , \6673 );
and \U$5692 ( \6675 , \6444 , \991 );
and \U$5693 ( \6676 , \6185 , \989 );
nor \U$5694 ( \6677 , \6675 , \6676 );
xnor \U$5695 ( \6678 , \6677 , \996 );
and \U$5696 ( \6679 , \6673 , \6678 );
and \U$5697 ( \6680 , \6669 , \6678 );
or \U$5698 ( \6681 , \6674 , \6679 , \6680 );
or \U$5699 ( \6682 , \6665 , \6681 );
and \U$5700 ( \6683 , \6648 , \6682 );
and \U$5701 ( \6684 , \6596 , \6682 );
or \U$5702 ( \6685 , \6649 , \6683 , \6684 );
xor \U$5703 ( \6686 , \6369 , \6373 );
xor \U$5704 ( \6687 , \6686 , \6378 );
xor \U$5705 ( \6688 , \6385 , \6389 );
xor \U$5706 ( \6689 , \6688 , \6394 );
and \U$5707 ( \6690 , \6687 , \6689 );
xor \U$5708 ( \6691 , \6350 , \6354 );
xor \U$5709 ( \6692 , \6691 , \6359 );
and \U$5710 ( \6693 , \6689 , \6692 );
and \U$5711 ( \6694 , \6687 , \6692 );
or \U$5712 ( \6695 , \6690 , \6693 , \6694 );
xor \U$5713 ( \6696 , \6402 , \6406 );
xor \U$5714 ( \6697 , \6696 , \6411 );
xor \U$5715 ( \6698 , \6422 , \6426 );
xor \U$5716 ( \6699 , \6698 , \6431 );
and \U$5717 ( \6700 , \6697 , \6699 );
xor \U$5718 ( \6701 , \6438 , \6442 );
xor \U$5719 ( \6702 , \6701 , \6445 );
and \U$5720 ( \6703 , \6699 , \6702 );
and \U$5721 ( \6704 , \6697 , \6702 );
or \U$5722 ( \6705 , \6700 , \6703 , \6704 );
and \U$5723 ( \6706 , \6695 , \6705 );
xor \U$5724 ( \6707 , \6317 , \6321 );
xor \U$5725 ( \6708 , \6707 , \6326 );
xor \U$5726 ( \6709 , \6333 , \6337 );
xor \U$5727 ( \6710 , \6709 , \6342 );
and \U$5728 ( \6711 , \6708 , \6710 );
and \U$5729 ( \6712 , \6705 , \6711 );
and \U$5730 ( \6713 , \6695 , \6711 );
or \U$5731 ( \6714 , \6706 , \6712 , \6713 );
and \U$5732 ( \6715 , \6685 , \6714 );
xor \U$5733 ( \6716 , \6074 , \6078 );
xor \U$5734 ( \6717 , \6716 , \6083 );
xor \U$5735 ( \6718 , \6459 , \6461 );
xor \U$5736 ( \6719 , \6718 , \6464 );
and \U$5737 ( \6720 , \6717 , \6719 );
xor \U$5738 ( \6721 , \6469 , \6471 );
xor \U$5739 ( \6722 , \6721 , \6474 );
and \U$5740 ( \6723 , \6719 , \6722 );
and \U$5741 ( \6724 , \6717 , \6722 );
or \U$5742 ( \6725 , \6720 , \6723 , \6724 );
and \U$5743 ( \6726 , \6714 , \6725 );
and \U$5744 ( \6727 , \6685 , \6725 );
or \U$5745 ( \6728 , \6715 , \6726 , \6727 );
xor \U$5746 ( \6729 , \6329 , \6345 );
xor \U$5747 ( \6730 , \6729 , \6362 );
xor \U$5748 ( \6731 , \6381 , \6397 );
xor \U$5749 ( \6732 , \6731 , \6414 );
and \U$5750 ( \6733 , \6730 , \6732 );
xor \U$5751 ( \6734 , \6434 , \6448 );
xor \U$5752 ( \6735 , \6734 , \6451 );
and \U$5753 ( \6736 , \6732 , \6735 );
and \U$5754 ( \6737 , \6730 , \6735 );
or \U$5755 ( \6738 , \6733 , \6736 , \6737 );
xor \U$5756 ( \6739 , \6086 , \6102 );
xor \U$5757 ( \6740 , \6739 , \6119 );
and \U$5758 ( \6741 , \6738 , \6740 );
xor \U$5759 ( \6742 , \6138 , \6154 );
xor \U$5760 ( \6743 , \6742 , \6171 );
and \U$5761 ( \6744 , \6740 , \6743 );
and \U$5762 ( \6745 , \6738 , \6743 );
or \U$5763 ( \6746 , \6741 , \6744 , \6745 );
and \U$5764 ( \6747 , \6728 , \6746 );
xor \U$5765 ( \6748 , \6365 , \6417 );
xor \U$5766 ( \6749 , \6748 , \6454 );
xor \U$5767 ( \6750 , \6467 , \6477 );
xor \U$5768 ( \6751 , \6750 , \6480 );
and \U$5769 ( \6752 , \6749 , \6751 );
xor \U$5770 ( \6753 , \6486 , \6488 );
xor \U$5771 ( \6754 , \6753 , \6491 );
and \U$5772 ( \6755 , \6751 , \6754 );
and \U$5773 ( \6756 , \6749 , \6754 );
or \U$5774 ( \6757 , \6752 , \6755 , \6756 );
and \U$5775 ( \6758 , \6746 , \6757 );
and \U$5776 ( \6759 , \6728 , \6757 );
or \U$5777 ( \6760 , \6747 , \6758 , \6759 );
xor \U$5778 ( \6761 , \6122 , \6174 );
xor \U$5779 ( \6762 , \6761 , \6210 );
xor \U$5780 ( \6763 , \6457 , \6483 );
xor \U$5781 ( \6764 , \6763 , \6494 );
and \U$5782 ( \6765 , \6762 , \6764 );
xor \U$5783 ( \6766 , \6499 , \6501 );
xor \U$5784 ( \6767 , \6766 , \6504 );
and \U$5785 ( \6768 , \6764 , \6767 );
and \U$5786 ( \6769 , \6762 , \6767 );
or \U$5787 ( \6770 , \6765 , \6768 , \6769 );
and \U$5788 ( \6771 , \6760 , \6770 );
xor \U$5789 ( \6772 , \6515 , \6517 );
xor \U$5790 ( \6773 , \6772 , \6520 );
and \U$5791 ( \6774 , \6770 , \6773 );
and \U$5792 ( \6775 , \6760 , \6773 );
or \U$5793 ( \6776 , \6771 , \6774 , \6775 );
xor \U$5794 ( \6777 , \6253 , \6271 );
xor \U$5795 ( \6778 , \6777 , \6274 );
and \U$5796 ( \6779 , \6776 , \6778 );
xor \U$5797 ( \6780 , \6513 , \6523 );
xor \U$5798 ( \6781 , \6780 , \6526 );
and \U$5799 ( \6782 , \6778 , \6781 );
and \U$5800 ( \6783 , \6776 , \6781 );
or \U$5801 ( \6784 , \6779 , \6782 , \6783 );
xor \U$5802 ( \6785 , \6529 , \6531 );
xor \U$5803 ( \6786 , \6785 , \6533 );
and \U$5804 ( \6787 , \6784 , \6786 );
and \U$5805 ( \6788 , \6542 , \6787 );
xor \U$5806 ( \6789 , \6542 , \6787 );
xor \U$5807 ( \6790 , \6784 , \6786 );
and \U$5808 ( \6791 , \4679 , \1360 );
and \U$5809 ( \6792 , \4557 , \1358 );
nor \U$5810 ( \6793 , \6791 , \6792 );
xnor \U$5811 ( \6794 , \6793 , \1317 );
and \U$5812 ( \6795 , \4940 , \1247 );
and \U$5813 ( \6796 , \4684 , \1245 );
nor \U$5814 ( \6797 , \6795 , \6796 );
xnor \U$5815 ( \6798 , \6797 , \1198 );
and \U$5816 ( \6799 , \6794 , \6798 );
and \U$5817 ( \6800 , \5439 , \1146 );
and \U$5818 ( \6801 , \5137 , \1144 );
nor \U$5819 ( \6802 , \6800 , \6801 );
xnor \U$5820 ( \6803 , \6802 , \1105 );
and \U$5821 ( \6804 , \6798 , \6803 );
and \U$5822 ( \6805 , \6794 , \6803 );
or \U$5823 ( \6806 , \6799 , \6804 , \6805 );
and \U$5824 ( \6807 , \5916 , \1076 );
and \U$5825 ( \6808 , \5447 , \1074 );
nor \U$5826 ( \6809 , \6807 , \6808 );
xnor \U$5827 ( \6810 , \6809 , \1046 );
and \U$5828 ( \6811 , \6185 , \1028 );
and \U$5829 ( \6812 , \5921 , \1026 );
nor \U$5830 ( \6813 , \6811 , \6812 );
xnor \U$5831 ( \6814 , \6813 , \1009 );
and \U$5832 ( \6815 , \6810 , \6814 );
buf \U$5833 ( \6816 , RIc0daa08_111);
and \U$5834 ( \6817 , \6816 , \991 );
and \U$5835 ( \6818 , \6444 , \989 );
nor \U$5836 ( \6819 , \6817 , \6818 );
xnor \U$5837 ( \6820 , \6819 , \996 );
and \U$5838 ( \6821 , \6814 , \6820 );
and \U$5839 ( \6822 , \6810 , \6820 );
or \U$5840 ( \6823 , \6815 , \6821 , \6822 );
and \U$5841 ( \6824 , \6806 , \6823 );
buf \U$5842 ( \6825 , RIc0daa80_112);
and \U$5843 ( \6826 , \6825 , \985 );
buf \U$5844 ( \6827 , \6826 );
and \U$5845 ( \6828 , \6823 , \6827 );
and \U$5846 ( \6829 , \6806 , \6827 );
or \U$5847 ( \6830 , \6824 , \6828 , \6829 );
and \U$5848 ( \6831 , \2710 , \2494 );
and \U$5849 ( \6832 , \2467 , \2492 );
nor \U$5850 ( \6833 , \6831 , \6832 );
xnor \U$5851 ( \6834 , \6833 , \2338 );
and \U$5852 ( \6835 , \2901 , \2222 );
and \U$5853 ( \6836 , \2715 , \2220 );
nor \U$5854 ( \6837 , \6835 , \6836 );
xnor \U$5855 ( \6838 , \6837 , \2109 );
and \U$5856 ( \6839 , \6834 , \6838 );
and \U$5857 ( \6840 , \3309 , \2028 );
and \U$5858 ( \6841 , \3045 , \2026 );
nor \U$5859 ( \6842 , \6840 , \6841 );
xnor \U$5860 ( \6843 , \6842 , \1892 );
and \U$5861 ( \6844 , \6838 , \6843 );
and \U$5862 ( \6845 , \6834 , \6843 );
or \U$5863 ( \6846 , \6839 , \6844 , \6845 );
and \U$5864 ( \6847 , \2047 , \3264 );
and \U$5865 ( \6848 , \1942 , \3262 );
nor \U$5866 ( \6849 , \6847 , \6848 );
xnor \U$5867 ( \6850 , \6849 , \3122 );
and \U$5868 ( \6851 , \2168 , \2968 );
and \U$5869 ( \6852 , \2052 , \2966 );
nor \U$5870 ( \6853 , \6851 , \6852 );
xnor \U$5871 ( \6854 , \6853 , \2831 );
and \U$5872 ( \6855 , \6850 , \6854 );
and \U$5873 ( \6856 , \2459 , \2762 );
and \U$5874 ( \6857 , \2283 , \2760 );
nor \U$5875 ( \6858 , \6856 , \6857 );
xnor \U$5876 ( \6859 , \6858 , \2610 );
and \U$5877 ( \6860 , \6854 , \6859 );
and \U$5878 ( \6861 , \6850 , \6859 );
or \U$5879 ( \6862 , \6855 , \6860 , \6861 );
and \U$5880 ( \6863 , \6846 , \6862 );
and \U$5881 ( \6864 , \3508 , \1828 );
and \U$5882 ( \6865 , \3334 , \1826 );
nor \U$5883 ( \6866 , \6864 , \6865 );
xnor \U$5884 ( \6867 , \6866 , \1750 );
and \U$5885 ( \6868 , \3813 , \1664 );
and \U$5886 ( \6869 , \3675 , \1662 );
nor \U$5887 ( \6870 , \6868 , \6869 );
xnor \U$5888 ( \6871 , \6870 , \1570 );
and \U$5889 ( \6872 , \6867 , \6871 );
and \U$5890 ( \6873 , \4349 , \1494 );
and \U$5891 ( \6874 , \3932 , \1492 );
nor \U$5892 ( \6875 , \6873 , \6874 );
xnor \U$5893 ( \6876 , \6875 , \1422 );
and \U$5894 ( \6877 , \6871 , \6876 );
and \U$5895 ( \6878 , \6867 , \6876 );
or \U$5896 ( \6879 , \6872 , \6877 , \6878 );
and \U$5897 ( \6880 , \6862 , \6879 );
and \U$5898 ( \6881 , \6846 , \6879 );
or \U$5899 ( \6882 , \6863 , \6880 , \6881 );
and \U$5900 ( \6883 , \6830 , \6882 );
and \U$5901 ( \6884 , \1162 , \5474 );
and \U$5902 ( \6885 , \1093 , \5472 );
nor \U$5903 ( \6886 , \6884 , \6885 );
xnor \U$5904 ( \6887 , \6886 , \5242 );
and \U$5905 ( \6888 , \1221 , \5023 );
and \U$5906 ( \6889 , \1167 , \5021 );
nor \U$5907 ( \6890 , \6888 , \6889 );
xnor \U$5908 ( \6891 , \6890 , \4880 );
and \U$5909 ( \6892 , \6887 , \6891 );
and \U$5910 ( \6893 , \1349 , \4700 );
and \U$5911 ( \6894 , \1272 , \4698 );
nor \U$5912 ( \6895 , \6893 , \6894 );
xnor \U$5913 ( \6896 , \6895 , \4454 );
and \U$5914 ( \6897 , \6891 , \6896 );
and \U$5915 ( \6898 , \6887 , \6896 );
or \U$5916 ( \6899 , \6892 , \6897 , \6898 );
xor \U$5917 ( \6900 , \6070 , \6559 );
xor \U$5918 ( \6901 , \6559 , \6560 );
not \U$5919 ( \6902 , \6901 );
and \U$5920 ( \6903 , \6900 , \6902 );
and \U$5921 ( \6904 , \984 , \6903 );
not \U$5922 ( \6905 , \6904 );
xnor \U$5923 ( \6906 , \6905 , \6563 );
and \U$5924 ( \6907 , \1016 , \6314 );
and \U$5925 ( \6908 , \998 , \6312 );
nor \U$5926 ( \6909 , \6907 , \6908 );
xnor \U$5927 ( \6910 , \6909 , \6073 );
and \U$5928 ( \6911 , \6906 , \6910 );
and \U$5929 ( \6912 , \1085 , \5848 );
and \U$5930 ( \6913 , \1037 , \5846 );
nor \U$5931 ( \6914 , \6912 , \6913 );
xnor \U$5932 ( \6915 , \6914 , \5660 );
and \U$5933 ( \6916 , \6910 , \6915 );
and \U$5934 ( \6917 , \6906 , \6915 );
or \U$5935 ( \6918 , \6911 , \6916 , \6917 );
and \U$5936 ( \6919 , \6899 , \6918 );
and \U$5937 ( \6920 , \1457 , \4305 );
and \U$5938 ( \6921 , \1377 , \4303 );
nor \U$5939 ( \6922 , \6920 , \6921 );
xnor \U$5940 ( \6923 , \6922 , \4118 );
and \U$5941 ( \6924 , \1593 , \3992 );
and \U$5942 ( \6925 , \1531 , \3990 );
nor \U$5943 ( \6926 , \6924 , \6925 );
xnor \U$5944 ( \6927 , \6926 , \3787 );
and \U$5945 ( \6928 , \6923 , \6927 );
and \U$5946 ( \6929 , \1854 , \3586 );
and \U$5947 ( \6930 , \1656 , \3584 );
nor \U$5948 ( \6931 , \6929 , \6930 );
xnor \U$5949 ( \6932 , \6931 , \3437 );
and \U$5950 ( \6933 , \6927 , \6932 );
and \U$5951 ( \6934 , \6923 , \6932 );
or \U$5952 ( \6935 , \6928 , \6933 , \6934 );
and \U$5953 ( \6936 , \6918 , \6935 );
and \U$5954 ( \6937 , \6899 , \6935 );
or \U$5955 ( \6938 , \6919 , \6936 , \6937 );
and \U$5956 ( \6939 , \6882 , \6938 );
and \U$5957 ( \6940 , \6830 , \6938 );
or \U$5958 ( \6941 , \6883 , \6939 , \6940 );
xor \U$5959 ( \6942 , \6546 , \6550 );
xor \U$5960 ( \6943 , \6942 , \6555 );
xor \U$5961 ( \6944 , \6564 , \6568 );
xor \U$5962 ( \6945 , \6944 , \6573 );
and \U$5963 ( \6946 , \6943 , \6945 );
xor \U$5964 ( \6947 , \6581 , \6585 );
xor \U$5965 ( \6948 , \6947 , \6590 );
and \U$5966 ( \6949 , \6945 , \6948 );
and \U$5967 ( \6950 , \6943 , \6948 );
or \U$5968 ( \6951 , \6946 , \6949 , \6950 );
xor \U$5969 ( \6952 , \6600 , \6604 );
xor \U$5970 ( \6953 , \6952 , \6609 );
xor \U$5971 ( \6954 , \6616 , \6620 );
xor \U$5972 ( \6955 , \6954 , \6625 );
and \U$5973 ( \6956 , \6953 , \6955 );
xor \U$5974 ( \6957 , \6633 , \6637 );
xor \U$5975 ( \6958 , \6957 , \6642 );
and \U$5976 ( \6959 , \6955 , \6958 );
and \U$5977 ( \6960 , \6953 , \6958 );
or \U$5978 ( \6961 , \6956 , \6959 , \6960 );
and \U$5979 ( \6962 , \6951 , \6961 );
and \U$5980 ( \6963 , \6816 , \985 );
xor \U$5981 ( \6964 , \6653 , \6657 );
xor \U$5982 ( \6965 , \6964 , \6662 );
and \U$5983 ( \6966 , \6963 , \6965 );
xor \U$5984 ( \6967 , \6669 , \6673 );
xor \U$5985 ( \6968 , \6967 , \6678 );
and \U$5986 ( \6969 , \6965 , \6968 );
and \U$5987 ( \6970 , \6963 , \6968 );
or \U$5988 ( \6971 , \6966 , \6969 , \6970 );
and \U$5989 ( \6972 , \6961 , \6971 );
and \U$5990 ( \6973 , \6951 , \6971 );
or \U$5991 ( \6974 , \6962 , \6972 , \6973 );
and \U$5992 ( \6975 , \6941 , \6974 );
xor \U$5993 ( \6976 , \6687 , \6689 );
xor \U$5994 ( \6977 , \6976 , \6692 );
xor \U$5995 ( \6978 , \6697 , \6699 );
xor \U$5996 ( \6979 , \6978 , \6702 );
and \U$5997 ( \6980 , \6977 , \6979 );
xor \U$5998 ( \6981 , \6708 , \6710 );
and \U$5999 ( \6982 , \6979 , \6981 );
and \U$6000 ( \6983 , \6977 , \6981 );
or \U$6001 ( \6984 , \6980 , \6982 , \6983 );
and \U$6002 ( \6985 , \6974 , \6984 );
and \U$6003 ( \6986 , \6941 , \6984 );
or \U$6004 ( \6987 , \6975 , \6985 , \6986 );
xor \U$6005 ( \6988 , \6558 , \6576 );
xor \U$6006 ( \6989 , \6988 , \6593 );
xor \U$6007 ( \6990 , \6612 , \6628 );
xor \U$6008 ( \6991 , \6990 , \6645 );
and \U$6009 ( \6992 , \6989 , \6991 );
xnor \U$6010 ( \6993 , \6665 , \6681 );
and \U$6011 ( \6994 , \6991 , \6993 );
and \U$6012 ( \6995 , \6989 , \6993 );
or \U$6013 ( \6996 , \6992 , \6994 , \6995 );
xor \U$6014 ( \6997 , \6717 , \6719 );
xor \U$6015 ( \6998 , \6997 , \6722 );
and \U$6016 ( \6999 , \6996 , \6998 );
xor \U$6017 ( \7000 , \6730 , \6732 );
xor \U$6018 ( \7001 , \7000 , \6735 );
and \U$6019 ( \7002 , \6998 , \7001 );
and \U$6020 ( \7003 , \6996 , \7001 );
or \U$6021 ( \7004 , \6999 , \7002 , \7003 );
and \U$6022 ( \7005 , \6987 , \7004 );
xor \U$6023 ( \7006 , \6596 , \6648 );
xor \U$6024 ( \7007 , \7006 , \6682 );
xor \U$6025 ( \7008 , \6695 , \6705 );
xor \U$6026 ( \7009 , \7008 , \6711 );
and \U$6027 ( \7010 , \7007 , \7009 );
and \U$6028 ( \7011 , \7004 , \7010 );
and \U$6029 ( \7012 , \6987 , \7010 );
or \U$6030 ( \7013 , \7005 , \7011 , \7012 );
xor \U$6031 ( \7014 , \6685 , \6714 );
xor \U$6032 ( \7015 , \7014 , \6725 );
xor \U$6033 ( \7016 , \6738 , \6740 );
xor \U$6034 ( \7017 , \7016 , \6743 );
and \U$6035 ( \7018 , \7015 , \7017 );
xor \U$6036 ( \7019 , \6749 , \6751 );
xor \U$6037 ( \7020 , \7019 , \6754 );
and \U$6038 ( \7021 , \7017 , \7020 );
and \U$6039 ( \7022 , \7015 , \7020 );
or \U$6040 ( \7023 , \7018 , \7021 , \7022 );
and \U$6041 ( \7024 , \7013 , \7023 );
xor \U$6042 ( \7025 , \6762 , \6764 );
xor \U$6043 ( \7026 , \7025 , \6767 );
and \U$6044 ( \7027 , \7023 , \7026 );
and \U$6045 ( \7028 , \7013 , \7026 );
or \U$6046 ( \7029 , \7024 , \7027 , \7028 );
xor \U$6047 ( \7030 , \6497 , \6507 );
xor \U$6048 ( \7031 , \7030 , \6510 );
and \U$6049 ( \7032 , \7029 , \7031 );
xor \U$6050 ( \7033 , \6760 , \6770 );
xor \U$6051 ( \7034 , \7033 , \6773 );
and \U$6052 ( \7035 , \7031 , \7034 );
and \U$6053 ( \7036 , \7029 , \7034 );
or \U$6054 ( \7037 , \7032 , \7035 , \7036 );
xor \U$6055 ( \7038 , \6776 , \6778 );
xor \U$6056 ( \7039 , \7038 , \6781 );
and \U$6057 ( \7040 , \7037 , \7039 );
and \U$6058 ( \7041 , \6790 , \7040 );
xor \U$6059 ( \7042 , \6790 , \7040 );
xor \U$6060 ( \7043 , \7037 , \7039 );
xor \U$6061 ( \7044 , \6834 , \6838 );
xor \U$6062 ( \7045 , \7044 , \6843 );
xor \U$6063 ( \7046 , \6850 , \6854 );
xor \U$6064 ( \7047 , \7046 , \6859 );
and \U$6065 ( \7048 , \7045 , \7047 );
xor \U$6066 ( \7049 , \6867 , \6871 );
xor \U$6067 ( \7050 , \7049 , \6876 );
and \U$6068 ( \7051 , \7047 , \7050 );
and \U$6069 ( \7052 , \7045 , \7050 );
or \U$6070 ( \7053 , \7048 , \7051 , \7052 );
xor \U$6071 ( \7054 , \6887 , \6891 );
xor \U$6072 ( \7055 , \7054 , \6896 );
xor \U$6073 ( \7056 , \6906 , \6910 );
xor \U$6074 ( \7057 , \7056 , \6915 );
and \U$6075 ( \7058 , \7055 , \7057 );
xor \U$6076 ( \7059 , \6923 , \6927 );
xor \U$6077 ( \7060 , \7059 , \6932 );
and \U$6078 ( \7061 , \7057 , \7060 );
and \U$6079 ( \7062 , \7055 , \7060 );
or \U$6080 ( \7063 , \7058 , \7061 , \7062 );
and \U$6081 ( \7064 , \7053 , \7063 );
xor \U$6082 ( \7065 , \6794 , \6798 );
xor \U$6083 ( \7066 , \7065 , \6803 );
xor \U$6084 ( \7067 , \6810 , \6814 );
xor \U$6085 ( \7068 , \7067 , \6820 );
and \U$6086 ( \7069 , \7066 , \7068 );
not \U$6087 ( \7070 , \6826 );
and \U$6088 ( \7071 , \7068 , \7070 );
and \U$6089 ( \7072 , \7066 , \7070 );
or \U$6090 ( \7073 , \7069 , \7071 , \7072 );
and \U$6091 ( \7074 , \7063 , \7073 );
and \U$6092 ( \7075 , \7053 , \7073 );
or \U$6093 ( \7076 , \7064 , \7074 , \7075 );
and \U$6094 ( \7077 , \1093 , \5848 );
and \U$6095 ( \7078 , \1085 , \5846 );
nor \U$6096 ( \7079 , \7077 , \7078 );
xnor \U$6097 ( \7080 , \7079 , \5660 );
and \U$6098 ( \7081 , \1167 , \5474 );
and \U$6099 ( \7082 , \1162 , \5472 );
nor \U$6100 ( \7083 , \7081 , \7082 );
xnor \U$6101 ( \7084 , \7083 , \5242 );
and \U$6102 ( \7085 , \7080 , \7084 );
and \U$6103 ( \7086 , \1272 , \5023 );
and \U$6104 ( \7087 , \1221 , \5021 );
nor \U$6105 ( \7088 , \7086 , \7087 );
xnor \U$6106 ( \7089 , \7088 , \4880 );
and \U$6107 ( \7090 , \7084 , \7089 );
and \U$6108 ( \7091 , \7080 , \7089 );
or \U$6109 ( \7092 , \7085 , \7090 , \7091 );
buf \U$6110 ( \7093 , RIc0d8d70_50);
buf \U$6111 ( \7094 , RIc0d8de8_51);
and \U$6112 ( \7095 , \7093 , \7094 );
not \U$6113 ( \7096 , \7095 );
and \U$6114 ( \7097 , \6560 , \7096 );
not \U$6115 ( \7098 , \7097 );
and \U$6116 ( \7099 , \998 , \6903 );
and \U$6117 ( \7100 , \984 , \6901 );
nor \U$6118 ( \7101 , \7099 , \7100 );
xnor \U$6119 ( \7102 , \7101 , \6563 );
and \U$6120 ( \7103 , \7098 , \7102 );
and \U$6121 ( \7104 , \1037 , \6314 );
and \U$6122 ( \7105 , \1016 , \6312 );
nor \U$6123 ( \7106 , \7104 , \7105 );
xnor \U$6124 ( \7107 , \7106 , \6073 );
and \U$6125 ( \7108 , \7102 , \7107 );
and \U$6126 ( \7109 , \7098 , \7107 );
or \U$6127 ( \7110 , \7103 , \7108 , \7109 );
and \U$6128 ( \7111 , \7092 , \7110 );
and \U$6129 ( \7112 , \1377 , \4700 );
and \U$6130 ( \7113 , \1349 , \4698 );
nor \U$6131 ( \7114 , \7112 , \7113 );
xnor \U$6132 ( \7115 , \7114 , \4454 );
and \U$6133 ( \7116 , \1531 , \4305 );
and \U$6134 ( \7117 , \1457 , \4303 );
nor \U$6135 ( \7118 , \7116 , \7117 );
xnor \U$6136 ( \7119 , \7118 , \4118 );
and \U$6137 ( \7120 , \7115 , \7119 );
and \U$6138 ( \7121 , \1656 , \3992 );
and \U$6139 ( \7122 , \1593 , \3990 );
nor \U$6140 ( \7123 , \7121 , \7122 );
xnor \U$6141 ( \7124 , \7123 , \3787 );
and \U$6142 ( \7125 , \7119 , \7124 );
and \U$6143 ( \7126 , \7115 , \7124 );
or \U$6144 ( \7127 , \7120 , \7125 , \7126 );
and \U$6145 ( \7128 , \7110 , \7127 );
and \U$6146 ( \7129 , \7092 , \7127 );
or \U$6147 ( \7130 , \7111 , \7128 , \7129 );
and \U$6148 ( \7131 , \4557 , \1494 );
and \U$6149 ( \7132 , \4349 , \1492 );
nor \U$6150 ( \7133 , \7131 , \7132 );
xnor \U$6151 ( \7134 , \7133 , \1422 );
and \U$6152 ( \7135 , \4684 , \1360 );
and \U$6153 ( \7136 , \4679 , \1358 );
nor \U$6154 ( \7137 , \7135 , \7136 );
xnor \U$6155 ( \7138 , \7137 , \1317 );
and \U$6156 ( \7139 , \7134 , \7138 );
and \U$6157 ( \7140 , \5137 , \1247 );
and \U$6158 ( \7141 , \4940 , \1245 );
nor \U$6159 ( \7142 , \7140 , \7141 );
xnor \U$6160 ( \7143 , \7142 , \1198 );
and \U$6161 ( \7144 , \7138 , \7143 );
and \U$6162 ( \7145 , \7134 , \7143 );
or \U$6163 ( \7146 , \7139 , \7144 , \7145 );
and \U$6164 ( \7147 , \5447 , \1146 );
and \U$6165 ( \7148 , \5439 , \1144 );
nor \U$6166 ( \7149 , \7147 , \7148 );
xnor \U$6167 ( \7150 , \7149 , \1105 );
and \U$6168 ( \7151 , \5921 , \1076 );
and \U$6169 ( \7152 , \5916 , \1074 );
nor \U$6170 ( \7153 , \7151 , \7152 );
xnor \U$6171 ( \7154 , \7153 , \1046 );
and \U$6172 ( \7155 , \7150 , \7154 );
and \U$6173 ( \7156 , \6444 , \1028 );
and \U$6174 ( \7157 , \6185 , \1026 );
nor \U$6175 ( \7158 , \7156 , \7157 );
xnor \U$6176 ( \7159 , \7158 , \1009 );
and \U$6177 ( \7160 , \7154 , \7159 );
and \U$6178 ( \7161 , \7150 , \7159 );
or \U$6179 ( \7162 , \7155 , \7160 , \7161 );
and \U$6180 ( \7163 , \7146 , \7162 );
and \U$6181 ( \7164 , \6825 , \991 );
and \U$6182 ( \7165 , \6816 , \989 );
nor \U$6183 ( \7166 , \7164 , \7165 );
xnor \U$6184 ( \7167 , \7166 , \996 );
buf \U$6185 ( \7168 , RIc0daaf8_113);
and \U$6186 ( \7169 , \7168 , \985 );
and \U$6187 ( \7170 , \7167 , \7169 );
and \U$6188 ( \7171 , \7162 , \7170 );
and \U$6189 ( \7172 , \7146 , \7170 );
or \U$6190 ( \7173 , \7163 , \7171 , \7172 );
and \U$6191 ( \7174 , \7130 , \7173 );
and \U$6192 ( \7175 , \1942 , \3586 );
and \U$6193 ( \7176 , \1854 , \3584 );
nor \U$6194 ( \7177 , \7175 , \7176 );
xnor \U$6195 ( \7178 , \7177 , \3437 );
and \U$6196 ( \7179 , \2052 , \3264 );
and \U$6197 ( \7180 , \2047 , \3262 );
nor \U$6198 ( \7181 , \7179 , \7180 );
xnor \U$6199 ( \7182 , \7181 , \3122 );
and \U$6200 ( \7183 , \7178 , \7182 );
and \U$6201 ( \7184 , \2283 , \2968 );
and \U$6202 ( \7185 , \2168 , \2966 );
nor \U$6203 ( \7186 , \7184 , \7185 );
xnor \U$6204 ( \7187 , \7186 , \2831 );
and \U$6205 ( \7188 , \7182 , \7187 );
and \U$6206 ( \7189 , \7178 , \7187 );
or \U$6207 ( \7190 , \7183 , \7188 , \7189 );
and \U$6208 ( \7191 , \2467 , \2762 );
and \U$6209 ( \7192 , \2459 , \2760 );
nor \U$6210 ( \7193 , \7191 , \7192 );
xnor \U$6211 ( \7194 , \7193 , \2610 );
and \U$6212 ( \7195 , \2715 , \2494 );
and \U$6213 ( \7196 , \2710 , \2492 );
nor \U$6214 ( \7197 , \7195 , \7196 );
xnor \U$6215 ( \7198 , \7197 , \2338 );
and \U$6216 ( \7199 , \7194 , \7198 );
and \U$6217 ( \7200 , \3045 , \2222 );
and \U$6218 ( \7201 , \2901 , \2220 );
nor \U$6219 ( \7202 , \7200 , \7201 );
xnor \U$6220 ( \7203 , \7202 , \2109 );
and \U$6221 ( \7204 , \7198 , \7203 );
and \U$6222 ( \7205 , \7194 , \7203 );
or \U$6223 ( \7206 , \7199 , \7204 , \7205 );
and \U$6224 ( \7207 , \7190 , \7206 );
and \U$6225 ( \7208 , \3334 , \2028 );
and \U$6226 ( \7209 , \3309 , \2026 );
nor \U$6227 ( \7210 , \7208 , \7209 );
xnor \U$6228 ( \7211 , \7210 , \1892 );
and \U$6229 ( \7212 , \3675 , \1828 );
and \U$6230 ( \7213 , \3508 , \1826 );
nor \U$6231 ( \7214 , \7212 , \7213 );
xnor \U$6232 ( \7215 , \7214 , \1750 );
and \U$6233 ( \7216 , \7211 , \7215 );
and \U$6234 ( \7217 , \3932 , \1664 );
and \U$6235 ( \7218 , \3813 , \1662 );
nor \U$6236 ( \7219 , \7217 , \7218 );
xnor \U$6237 ( \7220 , \7219 , \1570 );
and \U$6238 ( \7221 , \7215 , \7220 );
and \U$6239 ( \7222 , \7211 , \7220 );
or \U$6240 ( \7223 , \7216 , \7221 , \7222 );
and \U$6241 ( \7224 , \7206 , \7223 );
and \U$6242 ( \7225 , \7190 , \7223 );
or \U$6243 ( \7226 , \7207 , \7224 , \7225 );
and \U$6244 ( \7227 , \7173 , \7226 );
and \U$6245 ( \7228 , \7130 , \7226 );
or \U$6246 ( \7229 , \7174 , \7227 , \7228 );
and \U$6247 ( \7230 , \7076 , \7229 );
xor \U$6248 ( \7231 , \6943 , \6945 );
xor \U$6249 ( \7232 , \7231 , \6948 );
xor \U$6250 ( \7233 , \6953 , \6955 );
xor \U$6251 ( \7234 , \7233 , \6958 );
and \U$6252 ( \7235 , \7232 , \7234 );
xor \U$6253 ( \7236 , \6963 , \6965 );
xor \U$6254 ( \7237 , \7236 , \6968 );
and \U$6255 ( \7238 , \7234 , \7237 );
and \U$6256 ( \7239 , \7232 , \7237 );
or \U$6257 ( \7240 , \7235 , \7238 , \7239 );
and \U$6258 ( \7241 , \7229 , \7240 );
and \U$6259 ( \7242 , \7076 , \7240 );
or \U$6260 ( \7243 , \7230 , \7241 , \7242 );
xor \U$6261 ( \7244 , \6806 , \6823 );
xor \U$6262 ( \7245 , \7244 , \6827 );
xor \U$6263 ( \7246 , \6846 , \6862 );
xor \U$6264 ( \7247 , \7246 , \6879 );
and \U$6265 ( \7248 , \7245 , \7247 );
xor \U$6266 ( \7249 , \6899 , \6918 );
xor \U$6267 ( \7250 , \7249 , \6935 );
and \U$6268 ( \7251 , \7247 , \7250 );
and \U$6269 ( \7252 , \7245 , \7250 );
or \U$6270 ( \7253 , \7248 , \7251 , \7252 );
xor \U$6271 ( \7254 , \6989 , \6991 );
xor \U$6272 ( \7255 , \7254 , \6993 );
and \U$6273 ( \7256 , \7253 , \7255 );
xor \U$6274 ( \7257 , \6977 , \6979 );
xor \U$6275 ( \7258 , \7257 , \6981 );
and \U$6276 ( \7259 , \7255 , \7258 );
and \U$6277 ( \7260 , \7253 , \7258 );
or \U$6278 ( \7261 , \7256 , \7259 , \7260 );
and \U$6279 ( \7262 , \7243 , \7261 );
xor \U$6280 ( \7263 , \6830 , \6882 );
xor \U$6281 ( \7264 , \7263 , \6938 );
xor \U$6282 ( \7265 , \6951 , \6961 );
xor \U$6283 ( \7266 , \7265 , \6971 );
and \U$6284 ( \7267 , \7264 , \7266 );
and \U$6285 ( \7268 , \7261 , \7267 );
and \U$6286 ( \7269 , \7243 , \7267 );
or \U$6287 ( \7270 , \7262 , \7268 , \7269 );
xor \U$6288 ( \7271 , \6941 , \6974 );
xor \U$6289 ( \7272 , \7271 , \6984 );
xor \U$6290 ( \7273 , \6996 , \6998 );
xor \U$6291 ( \7274 , \7273 , \7001 );
and \U$6292 ( \7275 , \7272 , \7274 );
xor \U$6293 ( \7276 , \7007 , \7009 );
and \U$6294 ( \7277 , \7274 , \7276 );
and \U$6295 ( \7278 , \7272 , \7276 );
or \U$6296 ( \7279 , \7275 , \7277 , \7278 );
and \U$6297 ( \7280 , \7270 , \7279 );
xor \U$6298 ( \7281 , \7015 , \7017 );
xor \U$6299 ( \7282 , \7281 , \7020 );
and \U$6300 ( \7283 , \7279 , \7282 );
and \U$6301 ( \7284 , \7270 , \7282 );
or \U$6302 ( \7285 , \7280 , \7283 , \7284 );
xor \U$6303 ( \7286 , \6728 , \6746 );
xor \U$6304 ( \7287 , \7286 , \6757 );
and \U$6305 ( \7288 , \7285 , \7287 );
xor \U$6306 ( \7289 , \7013 , \7023 );
xor \U$6307 ( \7290 , \7289 , \7026 );
and \U$6308 ( \7291 , \7287 , \7290 );
and \U$6309 ( \7292 , \7285 , \7290 );
or \U$6310 ( \7293 , \7288 , \7291 , \7292 );
xor \U$6311 ( \7294 , \7029 , \7031 );
xor \U$6312 ( \7295 , \7294 , \7034 );
and \U$6313 ( \7296 , \7293 , \7295 );
and \U$6314 ( \7297 , \7043 , \7296 );
xor \U$6315 ( \7298 , \7043 , \7296 );
xor \U$6316 ( \7299 , \7293 , \7295 );
xor \U$6317 ( \7300 , \7178 , \7182 );
xor \U$6318 ( \7301 , \7300 , \7187 );
xor \U$6319 ( \7302 , \7194 , \7198 );
xor \U$6320 ( \7303 , \7302 , \7203 );
and \U$6321 ( \7304 , \7301 , \7303 );
xor \U$6322 ( \7305 , \7211 , \7215 );
xor \U$6323 ( \7306 , \7305 , \7220 );
and \U$6324 ( \7307 , \7303 , \7306 );
and \U$6325 ( \7308 , \7301 , \7306 );
or \U$6326 ( \7309 , \7304 , \7307 , \7308 );
xor \U$6327 ( \7310 , \7080 , \7084 );
xor \U$6328 ( \7311 , \7310 , \7089 );
xor \U$6329 ( \7312 , \7098 , \7102 );
xor \U$6330 ( \7313 , \7312 , \7107 );
and \U$6331 ( \7314 , \7311 , \7313 );
xor \U$6332 ( \7315 , \7115 , \7119 );
xor \U$6333 ( \7316 , \7315 , \7124 );
and \U$6334 ( \7317 , \7313 , \7316 );
and \U$6335 ( \7318 , \7311 , \7316 );
or \U$6336 ( \7319 , \7314 , \7317 , \7318 );
and \U$6337 ( \7320 , \7309 , \7319 );
xor \U$6338 ( \7321 , \7134 , \7138 );
xor \U$6339 ( \7322 , \7321 , \7143 );
xor \U$6340 ( \7323 , \7150 , \7154 );
xor \U$6341 ( \7324 , \7323 , \7159 );
and \U$6342 ( \7325 , \7322 , \7324 );
xor \U$6343 ( \7326 , \7167 , \7169 );
and \U$6344 ( \7327 , \7324 , \7326 );
and \U$6345 ( \7328 , \7322 , \7326 );
or \U$6346 ( \7329 , \7325 , \7327 , \7328 );
and \U$6347 ( \7330 , \7319 , \7329 );
and \U$6348 ( \7331 , \7309 , \7329 );
or \U$6349 ( \7332 , \7320 , \7330 , \7331 );
and \U$6350 ( \7333 , \4679 , \1494 );
and \U$6351 ( \7334 , \4557 , \1492 );
nor \U$6352 ( \7335 , \7333 , \7334 );
xnor \U$6353 ( \7336 , \7335 , \1422 );
and \U$6354 ( \7337 , \4940 , \1360 );
and \U$6355 ( \7338 , \4684 , \1358 );
nor \U$6356 ( \7339 , \7337 , \7338 );
xnor \U$6357 ( \7340 , \7339 , \1317 );
and \U$6358 ( \7341 , \7336 , \7340 );
and \U$6359 ( \7342 , \5439 , \1247 );
and \U$6360 ( \7343 , \5137 , \1245 );
nor \U$6361 ( \7344 , \7342 , \7343 );
xnor \U$6362 ( \7345 , \7344 , \1198 );
and \U$6363 ( \7346 , \7340 , \7345 );
and \U$6364 ( \7347 , \7336 , \7345 );
or \U$6365 ( \7348 , \7341 , \7346 , \7347 );
and \U$6366 ( \7349 , \5916 , \1146 );
and \U$6367 ( \7350 , \5447 , \1144 );
nor \U$6368 ( \7351 , \7349 , \7350 );
xnor \U$6369 ( \7352 , \7351 , \1105 );
and \U$6370 ( \7353 , \6185 , \1076 );
and \U$6371 ( \7354 , \5921 , \1074 );
nor \U$6372 ( \7355 , \7353 , \7354 );
xnor \U$6373 ( \7356 , \7355 , \1046 );
and \U$6374 ( \7357 , \7352 , \7356 );
and \U$6375 ( \7358 , \6816 , \1028 );
and \U$6376 ( \7359 , \6444 , \1026 );
nor \U$6377 ( \7360 , \7358 , \7359 );
xnor \U$6378 ( \7361 , \7360 , \1009 );
and \U$6379 ( \7362 , \7356 , \7361 );
and \U$6380 ( \7363 , \7352 , \7361 );
or \U$6381 ( \7364 , \7357 , \7362 , \7363 );
and \U$6382 ( \7365 , \7348 , \7364 );
and \U$6383 ( \7366 , \7168 , \991 );
and \U$6384 ( \7367 , \6825 , \989 );
nor \U$6385 ( \7368 , \7366 , \7367 );
xnor \U$6386 ( \7369 , \7368 , \996 );
buf \U$6387 ( \7370 , RIc0dab70_114);
and \U$6388 ( \7371 , \7370 , \985 );
or \U$6389 ( \7372 , \7369 , \7371 );
and \U$6390 ( \7373 , \7364 , \7372 );
and \U$6391 ( \7374 , \7348 , \7372 );
or \U$6392 ( \7375 , \7365 , \7373 , \7374 );
and \U$6393 ( \7376 , \1457 , \4700 );
and \U$6394 ( \7377 , \1377 , \4698 );
nor \U$6395 ( \7378 , \7376 , \7377 );
xnor \U$6396 ( \7379 , \7378 , \4454 );
and \U$6397 ( \7380 , \1593 , \4305 );
and \U$6398 ( \7381 , \1531 , \4303 );
nor \U$6399 ( \7382 , \7380 , \7381 );
xnor \U$6400 ( \7383 , \7382 , \4118 );
and \U$6401 ( \7384 , \7379 , \7383 );
and \U$6402 ( \7385 , \1854 , \3992 );
and \U$6403 ( \7386 , \1656 , \3990 );
nor \U$6404 ( \7387 , \7385 , \7386 );
xnor \U$6405 ( \7388 , \7387 , \3787 );
and \U$6406 ( \7389 , \7383 , \7388 );
and \U$6407 ( \7390 , \7379 , \7388 );
or \U$6408 ( \7391 , \7384 , \7389 , \7390 );
and \U$6409 ( \7392 , \1162 , \5848 );
and \U$6410 ( \7393 , \1093 , \5846 );
nor \U$6411 ( \7394 , \7392 , \7393 );
xnor \U$6412 ( \7395 , \7394 , \5660 );
and \U$6413 ( \7396 , \1221 , \5474 );
and \U$6414 ( \7397 , \1167 , \5472 );
nor \U$6415 ( \7398 , \7396 , \7397 );
xnor \U$6416 ( \7399 , \7398 , \5242 );
and \U$6417 ( \7400 , \7395 , \7399 );
and \U$6418 ( \7401 , \1349 , \5023 );
and \U$6419 ( \7402 , \1272 , \5021 );
nor \U$6420 ( \7403 , \7401 , \7402 );
xnor \U$6421 ( \7404 , \7403 , \4880 );
and \U$6422 ( \7405 , \7399 , \7404 );
and \U$6423 ( \7406 , \7395 , \7404 );
or \U$6424 ( \7407 , \7400 , \7405 , \7406 );
and \U$6425 ( \7408 , \7391 , \7407 );
xor \U$6426 ( \7409 , \6560 , \7093 );
xor \U$6427 ( \7410 , \7093 , \7094 );
not \U$6428 ( \7411 , \7410 );
and \U$6429 ( \7412 , \7409 , \7411 );
and \U$6430 ( \7413 , \984 , \7412 );
not \U$6431 ( \7414 , \7413 );
xnor \U$6432 ( \7415 , \7414 , \7097 );
and \U$6433 ( \7416 , \1016 , \6903 );
and \U$6434 ( \7417 , \998 , \6901 );
nor \U$6435 ( \7418 , \7416 , \7417 );
xnor \U$6436 ( \7419 , \7418 , \6563 );
and \U$6437 ( \7420 , \7415 , \7419 );
and \U$6438 ( \7421 , \1085 , \6314 );
and \U$6439 ( \7422 , \1037 , \6312 );
nor \U$6440 ( \7423 , \7421 , \7422 );
xnor \U$6441 ( \7424 , \7423 , \6073 );
and \U$6442 ( \7425 , \7419 , \7424 );
and \U$6443 ( \7426 , \7415 , \7424 );
or \U$6444 ( \7427 , \7420 , \7425 , \7426 );
and \U$6445 ( \7428 , \7407 , \7427 );
and \U$6446 ( \7429 , \7391 , \7427 );
or \U$6447 ( \7430 , \7408 , \7428 , \7429 );
and \U$6448 ( \7431 , \7375 , \7430 );
and \U$6449 ( \7432 , \2710 , \2762 );
and \U$6450 ( \7433 , \2467 , \2760 );
nor \U$6451 ( \7434 , \7432 , \7433 );
xnor \U$6452 ( \7435 , \7434 , \2610 );
and \U$6453 ( \7436 , \2901 , \2494 );
and \U$6454 ( \7437 , \2715 , \2492 );
nor \U$6455 ( \7438 , \7436 , \7437 );
xnor \U$6456 ( \7439 , \7438 , \2338 );
and \U$6457 ( \7440 , \7435 , \7439 );
and \U$6458 ( \7441 , \3309 , \2222 );
and \U$6459 ( \7442 , \3045 , \2220 );
nor \U$6460 ( \7443 , \7441 , \7442 );
xnor \U$6461 ( \7444 , \7443 , \2109 );
and \U$6462 ( \7445 , \7439 , \7444 );
and \U$6463 ( \7446 , \7435 , \7444 );
or \U$6464 ( \7447 , \7440 , \7445 , \7446 );
and \U$6465 ( \7448 , \3508 , \2028 );
and \U$6466 ( \7449 , \3334 , \2026 );
nor \U$6467 ( \7450 , \7448 , \7449 );
xnor \U$6468 ( \7451 , \7450 , \1892 );
and \U$6469 ( \7452 , \3813 , \1828 );
and \U$6470 ( \7453 , \3675 , \1826 );
nor \U$6471 ( \7454 , \7452 , \7453 );
xnor \U$6472 ( \7455 , \7454 , \1750 );
and \U$6473 ( \7456 , \7451 , \7455 );
and \U$6474 ( \7457 , \4349 , \1664 );
and \U$6475 ( \7458 , \3932 , \1662 );
nor \U$6476 ( \7459 , \7457 , \7458 );
xnor \U$6477 ( \7460 , \7459 , \1570 );
and \U$6478 ( \7461 , \7455 , \7460 );
and \U$6479 ( \7462 , \7451 , \7460 );
or \U$6480 ( \7463 , \7456 , \7461 , \7462 );
and \U$6481 ( \7464 , \7447 , \7463 );
and \U$6482 ( \7465 , \2047 , \3586 );
and \U$6483 ( \7466 , \1942 , \3584 );
nor \U$6484 ( \7467 , \7465 , \7466 );
xnor \U$6485 ( \7468 , \7467 , \3437 );
and \U$6486 ( \7469 , \2168 , \3264 );
and \U$6487 ( \7470 , \2052 , \3262 );
nor \U$6488 ( \7471 , \7469 , \7470 );
xnor \U$6489 ( \7472 , \7471 , \3122 );
and \U$6490 ( \7473 , \7468 , \7472 );
and \U$6491 ( \7474 , \2459 , \2968 );
and \U$6492 ( \7475 , \2283 , \2966 );
nor \U$6493 ( \7476 , \7474 , \7475 );
xnor \U$6494 ( \7477 , \7476 , \2831 );
and \U$6495 ( \7478 , \7472 , \7477 );
and \U$6496 ( \7479 , \7468 , \7477 );
or \U$6497 ( \7480 , \7473 , \7478 , \7479 );
and \U$6498 ( \7481 , \7463 , \7480 );
and \U$6499 ( \7482 , \7447 , \7480 );
or \U$6500 ( \7483 , \7464 , \7481 , \7482 );
and \U$6501 ( \7484 , \7430 , \7483 );
and \U$6502 ( \7485 , \7375 , \7483 );
or \U$6503 ( \7486 , \7431 , \7484 , \7485 );
and \U$6504 ( \7487 , \7332 , \7486 );
xor \U$6505 ( \7488 , \7045 , \7047 );
xor \U$6506 ( \7489 , \7488 , \7050 );
xor \U$6507 ( \7490 , \7055 , \7057 );
xor \U$6508 ( \7491 , \7490 , \7060 );
and \U$6509 ( \7492 , \7489 , \7491 );
xor \U$6510 ( \7493 , \7066 , \7068 );
xor \U$6511 ( \7494 , \7493 , \7070 );
and \U$6512 ( \7495 , \7491 , \7494 );
and \U$6513 ( \7496 , \7489 , \7494 );
or \U$6514 ( \7497 , \7492 , \7495 , \7496 );
and \U$6515 ( \7498 , \7486 , \7497 );
and \U$6516 ( \7499 , \7332 , \7497 );
or \U$6517 ( \7500 , \7487 , \7498 , \7499 );
xor \U$6518 ( \7501 , \7092 , \7110 );
xor \U$6519 ( \7502 , \7501 , \7127 );
xor \U$6520 ( \7503 , \7146 , \7162 );
xor \U$6521 ( \7504 , \7503 , \7170 );
and \U$6522 ( \7505 , \7502 , \7504 );
xor \U$6523 ( \7506 , \7190 , \7206 );
xor \U$6524 ( \7507 , \7506 , \7223 );
and \U$6525 ( \7508 , \7504 , \7507 );
and \U$6526 ( \7509 , \7502 , \7507 );
or \U$6527 ( \7510 , \7505 , \7508 , \7509 );
xor \U$6528 ( \7511 , \7245 , \7247 );
xor \U$6529 ( \7512 , \7511 , \7250 );
and \U$6530 ( \7513 , \7510 , \7512 );
xor \U$6531 ( \7514 , \7232 , \7234 );
xor \U$6532 ( \7515 , \7514 , \7237 );
and \U$6533 ( \7516 , \7512 , \7515 );
and \U$6534 ( \7517 , \7510 , \7515 );
or \U$6535 ( \7518 , \7513 , \7516 , \7517 );
and \U$6536 ( \7519 , \7500 , \7518 );
xor \U$6537 ( \7520 , \7053 , \7063 );
xor \U$6538 ( \7521 , \7520 , \7073 );
xor \U$6539 ( \7522 , \7130 , \7173 );
xor \U$6540 ( \7523 , \7522 , \7226 );
and \U$6541 ( \7524 , \7521 , \7523 );
and \U$6542 ( \7525 , \7518 , \7524 );
and \U$6543 ( \7526 , \7500 , \7524 );
or \U$6544 ( \7527 , \7519 , \7525 , \7526 );
xor \U$6545 ( \7528 , \7076 , \7229 );
xor \U$6546 ( \7529 , \7528 , \7240 );
xor \U$6547 ( \7530 , \7253 , \7255 );
xor \U$6548 ( \7531 , \7530 , \7258 );
and \U$6549 ( \7532 , \7529 , \7531 );
xor \U$6550 ( \7533 , \7264 , \7266 );
and \U$6551 ( \7534 , \7531 , \7533 );
and \U$6552 ( \7535 , \7529 , \7533 );
or \U$6553 ( \7536 , \7532 , \7534 , \7535 );
and \U$6554 ( \7537 , \7527 , \7536 );
xor \U$6555 ( \7538 , \7272 , \7274 );
xor \U$6556 ( \7539 , \7538 , \7276 );
and \U$6557 ( \7540 , \7536 , \7539 );
and \U$6558 ( \7541 , \7527 , \7539 );
or \U$6559 ( \7542 , \7537 , \7540 , \7541 );
xor \U$6560 ( \7543 , \6987 , \7004 );
xor \U$6561 ( \7544 , \7543 , \7010 );
and \U$6562 ( \7545 , \7542 , \7544 );
xor \U$6563 ( \7546 , \7270 , \7279 );
xor \U$6564 ( \7547 , \7546 , \7282 );
and \U$6565 ( \7548 , \7544 , \7547 );
and \U$6566 ( \7549 , \7542 , \7547 );
or \U$6567 ( \7550 , \7545 , \7548 , \7549 );
xor \U$6568 ( \7551 , \7285 , \7287 );
xor \U$6569 ( \7552 , \7551 , \7290 );
and \U$6570 ( \7553 , \7550 , \7552 );
and \U$6571 ( \7554 , \7299 , \7553 );
xor \U$6572 ( \7555 , \7299 , \7553 );
xor \U$6573 ( \7556 , \7550 , \7552 );
and \U$6574 ( \7557 , \1942 , \3992 );
and \U$6575 ( \7558 , \1854 , \3990 );
nor \U$6576 ( \7559 , \7557 , \7558 );
xnor \U$6577 ( \7560 , \7559 , \3787 );
and \U$6578 ( \7561 , \2052 , \3586 );
and \U$6579 ( \7562 , \2047 , \3584 );
nor \U$6580 ( \7563 , \7561 , \7562 );
xnor \U$6581 ( \7564 , \7563 , \3437 );
and \U$6582 ( \7565 , \7560 , \7564 );
and \U$6583 ( \7566 , \2283 , \3264 );
and \U$6584 ( \7567 , \2168 , \3262 );
nor \U$6585 ( \7568 , \7566 , \7567 );
xnor \U$6586 ( \7569 , \7568 , \3122 );
and \U$6587 ( \7570 , \7564 , \7569 );
and \U$6588 ( \7571 , \7560 , \7569 );
or \U$6589 ( \7572 , \7565 , \7570 , \7571 );
and \U$6590 ( \7573 , \2467 , \2968 );
and \U$6591 ( \7574 , \2459 , \2966 );
nor \U$6592 ( \7575 , \7573 , \7574 );
xnor \U$6593 ( \7576 , \7575 , \2831 );
and \U$6594 ( \7577 , \2715 , \2762 );
and \U$6595 ( \7578 , \2710 , \2760 );
nor \U$6596 ( \7579 , \7577 , \7578 );
xnor \U$6597 ( \7580 , \7579 , \2610 );
and \U$6598 ( \7581 , \7576 , \7580 );
and \U$6599 ( \7582 , \3045 , \2494 );
and \U$6600 ( \7583 , \2901 , \2492 );
nor \U$6601 ( \7584 , \7582 , \7583 );
xnor \U$6602 ( \7585 , \7584 , \2338 );
and \U$6603 ( \7586 , \7580 , \7585 );
and \U$6604 ( \7587 , \7576 , \7585 );
or \U$6605 ( \7588 , \7581 , \7586 , \7587 );
and \U$6606 ( \7589 , \7572 , \7588 );
and \U$6607 ( \7590 , \3334 , \2222 );
and \U$6608 ( \7591 , \3309 , \2220 );
nor \U$6609 ( \7592 , \7590 , \7591 );
xnor \U$6610 ( \7593 , \7592 , \2109 );
and \U$6611 ( \7594 , \3675 , \2028 );
and \U$6612 ( \7595 , \3508 , \2026 );
nor \U$6613 ( \7596 , \7594 , \7595 );
xnor \U$6614 ( \7597 , \7596 , \1892 );
and \U$6615 ( \7598 , \7593 , \7597 );
and \U$6616 ( \7599 , \3932 , \1828 );
and \U$6617 ( \7600 , \3813 , \1826 );
nor \U$6618 ( \7601 , \7599 , \7600 );
xnor \U$6619 ( \7602 , \7601 , \1750 );
and \U$6620 ( \7603 , \7597 , \7602 );
and \U$6621 ( \7604 , \7593 , \7602 );
or \U$6622 ( \7605 , \7598 , \7603 , \7604 );
and \U$6623 ( \7606 , \7588 , \7605 );
and \U$6624 ( \7607 , \7572 , \7605 );
or \U$6625 ( \7608 , \7589 , \7606 , \7607 );
and \U$6626 ( \7609 , \1093 , \6314 );
and \U$6627 ( \7610 , \1085 , \6312 );
nor \U$6628 ( \7611 , \7609 , \7610 );
xnor \U$6629 ( \7612 , \7611 , \6073 );
and \U$6630 ( \7613 , \1167 , \5848 );
and \U$6631 ( \7614 , \1162 , \5846 );
nor \U$6632 ( \7615 , \7613 , \7614 );
xnor \U$6633 ( \7616 , \7615 , \5660 );
and \U$6634 ( \7617 , \7612 , \7616 );
and \U$6635 ( \7618 , \1272 , \5474 );
and \U$6636 ( \7619 , \1221 , \5472 );
nor \U$6637 ( \7620 , \7618 , \7619 );
xnor \U$6638 ( \7621 , \7620 , \5242 );
and \U$6639 ( \7622 , \7616 , \7621 );
and \U$6640 ( \7623 , \7612 , \7621 );
or \U$6641 ( \7624 , \7617 , \7622 , \7623 );
and \U$6642 ( \7625 , \1377 , \5023 );
and \U$6643 ( \7626 , \1349 , \5021 );
nor \U$6644 ( \7627 , \7625 , \7626 );
xnor \U$6645 ( \7628 , \7627 , \4880 );
and \U$6646 ( \7629 , \1531 , \4700 );
and \U$6647 ( \7630 , \1457 , \4698 );
nor \U$6648 ( \7631 , \7629 , \7630 );
xnor \U$6649 ( \7632 , \7631 , \4454 );
and \U$6650 ( \7633 , \7628 , \7632 );
and \U$6651 ( \7634 , \1656 , \4305 );
and \U$6652 ( \7635 , \1593 , \4303 );
nor \U$6653 ( \7636 , \7634 , \7635 );
xnor \U$6654 ( \7637 , \7636 , \4118 );
and \U$6655 ( \7638 , \7632 , \7637 );
and \U$6656 ( \7639 , \7628 , \7637 );
or \U$6657 ( \7640 , \7633 , \7638 , \7639 );
and \U$6658 ( \7641 , \7624 , \7640 );
buf \U$6659 ( \7642 , RIc0d8e60_52);
buf \U$6660 ( \7643 , RIc0d8ed8_53);
and \U$6661 ( \7644 , \7642 , \7643 );
not \U$6662 ( \7645 , \7644 );
and \U$6663 ( \7646 , \7094 , \7645 );
not \U$6664 ( \7647 , \7646 );
and \U$6665 ( \7648 , \998 , \7412 );
and \U$6666 ( \7649 , \984 , \7410 );
nor \U$6667 ( \7650 , \7648 , \7649 );
xnor \U$6668 ( \7651 , \7650 , \7097 );
and \U$6669 ( \7652 , \7647 , \7651 );
and \U$6670 ( \7653 , \1037 , \6903 );
and \U$6671 ( \7654 , \1016 , \6901 );
nor \U$6672 ( \7655 , \7653 , \7654 );
xnor \U$6673 ( \7656 , \7655 , \6563 );
and \U$6674 ( \7657 , \7651 , \7656 );
and \U$6675 ( \7658 , \7647 , \7656 );
or \U$6676 ( \7659 , \7652 , \7657 , \7658 );
and \U$6677 ( \7660 , \7640 , \7659 );
and \U$6678 ( \7661 , \7624 , \7659 );
or \U$6679 ( \7662 , \7641 , \7660 , \7661 );
and \U$6680 ( \7663 , \7608 , \7662 );
and \U$6681 ( \7664 , \6825 , \1028 );
and \U$6682 ( \7665 , \6816 , \1026 );
nor \U$6683 ( \7666 , \7664 , \7665 );
xnor \U$6684 ( \7667 , \7666 , \1009 );
and \U$6685 ( \7668 , \7370 , \991 );
and \U$6686 ( \7669 , \7168 , \989 );
nor \U$6687 ( \7670 , \7668 , \7669 );
xnor \U$6688 ( \7671 , \7670 , \996 );
and \U$6689 ( \7672 , \7667 , \7671 );
buf \U$6690 ( \7673 , RIc0dabe8_115);
and \U$6691 ( \7674 , \7673 , \985 );
and \U$6692 ( \7675 , \7671 , \7674 );
and \U$6693 ( \7676 , \7667 , \7674 );
or \U$6694 ( \7677 , \7672 , \7675 , \7676 );
and \U$6695 ( \7678 , \4557 , \1664 );
and \U$6696 ( \7679 , \4349 , \1662 );
nor \U$6697 ( \7680 , \7678 , \7679 );
xnor \U$6698 ( \7681 , \7680 , \1570 );
and \U$6699 ( \7682 , \4684 , \1494 );
and \U$6700 ( \7683 , \4679 , \1492 );
nor \U$6701 ( \7684 , \7682 , \7683 );
xnor \U$6702 ( \7685 , \7684 , \1422 );
and \U$6703 ( \7686 , \7681 , \7685 );
and \U$6704 ( \7687 , \5137 , \1360 );
and \U$6705 ( \7688 , \4940 , \1358 );
nor \U$6706 ( \7689 , \7687 , \7688 );
xnor \U$6707 ( \7690 , \7689 , \1317 );
and \U$6708 ( \7691 , \7685 , \7690 );
and \U$6709 ( \7692 , \7681 , \7690 );
or \U$6710 ( \7693 , \7686 , \7691 , \7692 );
and \U$6711 ( \7694 , \7677 , \7693 );
and \U$6712 ( \7695 , \5447 , \1247 );
and \U$6713 ( \7696 , \5439 , \1245 );
nor \U$6714 ( \7697 , \7695 , \7696 );
xnor \U$6715 ( \7698 , \7697 , \1198 );
and \U$6716 ( \7699 , \5921 , \1146 );
and \U$6717 ( \7700 , \5916 , \1144 );
nor \U$6718 ( \7701 , \7699 , \7700 );
xnor \U$6719 ( \7702 , \7701 , \1105 );
and \U$6720 ( \7703 , \7698 , \7702 );
and \U$6721 ( \7704 , \6444 , \1076 );
and \U$6722 ( \7705 , \6185 , \1074 );
nor \U$6723 ( \7706 , \7704 , \7705 );
xnor \U$6724 ( \7707 , \7706 , \1046 );
and \U$6725 ( \7708 , \7702 , \7707 );
and \U$6726 ( \7709 , \7698 , \7707 );
or \U$6727 ( \7710 , \7703 , \7708 , \7709 );
and \U$6728 ( \7711 , \7693 , \7710 );
and \U$6729 ( \7712 , \7677 , \7710 );
or \U$6730 ( \7713 , \7694 , \7711 , \7712 );
and \U$6731 ( \7714 , \7662 , \7713 );
and \U$6732 ( \7715 , \7608 , \7713 );
or \U$6733 ( \7716 , \7663 , \7714 , \7715 );
xor \U$6734 ( \7717 , \7435 , \7439 );
xor \U$6735 ( \7718 , \7717 , \7444 );
xor \U$6736 ( \7719 , \7451 , \7455 );
xor \U$6737 ( \7720 , \7719 , \7460 );
and \U$6738 ( \7721 , \7718 , \7720 );
xor \U$6739 ( \7722 , \7468 , \7472 );
xor \U$6740 ( \7723 , \7722 , \7477 );
and \U$6741 ( \7724 , \7720 , \7723 );
and \U$6742 ( \7725 , \7718 , \7723 );
or \U$6743 ( \7726 , \7721 , \7724 , \7725 );
xor \U$6744 ( \7727 , \7379 , \7383 );
xor \U$6745 ( \7728 , \7727 , \7388 );
xor \U$6746 ( \7729 , \7395 , \7399 );
xor \U$6747 ( \7730 , \7729 , \7404 );
and \U$6748 ( \7731 , \7728 , \7730 );
xor \U$6749 ( \7732 , \7415 , \7419 );
xor \U$6750 ( \7733 , \7732 , \7424 );
and \U$6751 ( \7734 , \7730 , \7733 );
and \U$6752 ( \7735 , \7728 , \7733 );
or \U$6753 ( \7736 , \7731 , \7734 , \7735 );
and \U$6754 ( \7737 , \7726 , \7736 );
xor \U$6755 ( \7738 , \7336 , \7340 );
xor \U$6756 ( \7739 , \7738 , \7345 );
xor \U$6757 ( \7740 , \7352 , \7356 );
xor \U$6758 ( \7741 , \7740 , \7361 );
and \U$6759 ( \7742 , \7739 , \7741 );
xnor \U$6760 ( \7743 , \7369 , \7371 );
and \U$6761 ( \7744 , \7741 , \7743 );
and \U$6762 ( \7745 , \7739 , \7743 );
or \U$6763 ( \7746 , \7742 , \7744 , \7745 );
and \U$6764 ( \7747 , \7736 , \7746 );
and \U$6765 ( \7748 , \7726 , \7746 );
or \U$6766 ( \7749 , \7737 , \7747 , \7748 );
and \U$6767 ( \7750 , \7716 , \7749 );
xor \U$6768 ( \7751 , \7301 , \7303 );
xor \U$6769 ( \7752 , \7751 , \7306 );
xor \U$6770 ( \7753 , \7311 , \7313 );
xor \U$6771 ( \7754 , \7753 , \7316 );
and \U$6772 ( \7755 , \7752 , \7754 );
xor \U$6773 ( \7756 , \7322 , \7324 );
xor \U$6774 ( \7757 , \7756 , \7326 );
and \U$6775 ( \7758 , \7754 , \7757 );
and \U$6776 ( \7759 , \7752 , \7757 );
or \U$6777 ( \7760 , \7755 , \7758 , \7759 );
and \U$6778 ( \7761 , \7749 , \7760 );
and \U$6779 ( \7762 , \7716 , \7760 );
or \U$6780 ( \7763 , \7750 , \7761 , \7762 );
xor \U$6781 ( \7764 , \7348 , \7364 );
xor \U$6782 ( \7765 , \7764 , \7372 );
xor \U$6783 ( \7766 , \7391 , \7407 );
xor \U$6784 ( \7767 , \7766 , \7427 );
and \U$6785 ( \7768 , \7765 , \7767 );
xor \U$6786 ( \7769 , \7447 , \7463 );
xor \U$6787 ( \7770 , \7769 , \7480 );
and \U$6788 ( \7771 , \7767 , \7770 );
and \U$6789 ( \7772 , \7765 , \7770 );
or \U$6790 ( \7773 , \7768 , \7771 , \7772 );
xor \U$6791 ( \7774 , \7502 , \7504 );
xor \U$6792 ( \7775 , \7774 , \7507 );
and \U$6793 ( \7776 , \7773 , \7775 );
xor \U$6794 ( \7777 , \7489 , \7491 );
xor \U$6795 ( \7778 , \7777 , \7494 );
and \U$6796 ( \7779 , \7775 , \7778 );
and \U$6797 ( \7780 , \7773 , \7778 );
or \U$6798 ( \7781 , \7776 , \7779 , \7780 );
and \U$6799 ( \7782 , \7763 , \7781 );
xor \U$6800 ( \7783 , \7309 , \7319 );
xor \U$6801 ( \7784 , \7783 , \7329 );
xor \U$6802 ( \7785 , \7375 , \7430 );
xor \U$6803 ( \7786 , \7785 , \7483 );
and \U$6804 ( \7787 , \7784 , \7786 );
and \U$6805 ( \7788 , \7781 , \7787 );
and \U$6806 ( \7789 , \7763 , \7787 );
or \U$6807 ( \7790 , \7782 , \7788 , \7789 );
xor \U$6808 ( \7791 , \7332 , \7486 );
xor \U$6809 ( \7792 , \7791 , \7497 );
xor \U$6810 ( \7793 , \7510 , \7512 );
xor \U$6811 ( \7794 , \7793 , \7515 );
and \U$6812 ( \7795 , \7792 , \7794 );
xor \U$6813 ( \7796 , \7521 , \7523 );
and \U$6814 ( \7797 , \7794 , \7796 );
and \U$6815 ( \7798 , \7792 , \7796 );
or \U$6816 ( \7799 , \7795 , \7797 , \7798 );
and \U$6817 ( \7800 , \7790 , \7799 );
xor \U$6818 ( \7801 , \7529 , \7531 );
xor \U$6819 ( \7802 , \7801 , \7533 );
and \U$6820 ( \7803 , \7799 , \7802 );
and \U$6821 ( \7804 , \7790 , \7802 );
or \U$6822 ( \7805 , \7800 , \7803 , \7804 );
xor \U$6823 ( \7806 , \7243 , \7261 );
xor \U$6824 ( \7807 , \7806 , \7267 );
and \U$6825 ( \7808 , \7805 , \7807 );
xor \U$6826 ( \7809 , \7527 , \7536 );
xor \U$6827 ( \7810 , \7809 , \7539 );
and \U$6828 ( \7811 , \7807 , \7810 );
and \U$6829 ( \7812 , \7805 , \7810 );
or \U$6830 ( \7813 , \7808 , \7811 , \7812 );
xor \U$6831 ( \7814 , \7542 , \7544 );
xor \U$6832 ( \7815 , \7814 , \7547 );
and \U$6833 ( \7816 , \7813 , \7815 );
and \U$6834 ( \7817 , \7556 , \7816 );
xor \U$6835 ( \7818 , \7556 , \7816 );
xor \U$6836 ( \7819 , \7813 , \7815 );
and \U$6837 ( \7820 , \4679 , \1664 );
and \U$6838 ( \7821 , \4557 , \1662 );
nor \U$6839 ( \7822 , \7820 , \7821 );
xnor \U$6840 ( \7823 , \7822 , \1570 );
and \U$6841 ( \7824 , \4940 , \1494 );
and \U$6842 ( \7825 , \4684 , \1492 );
nor \U$6843 ( \7826 , \7824 , \7825 );
xnor \U$6844 ( \7827 , \7826 , \1422 );
and \U$6845 ( \7828 , \7823 , \7827 );
and \U$6846 ( \7829 , \5439 , \1360 );
and \U$6847 ( \7830 , \5137 , \1358 );
nor \U$6848 ( \7831 , \7829 , \7830 );
xnor \U$6849 ( \7832 , \7831 , \1317 );
and \U$6850 ( \7833 , \7827 , \7832 );
and \U$6851 ( \7834 , \7823 , \7832 );
or \U$6852 ( \7835 , \7828 , \7833 , \7834 );
and \U$6853 ( \7836 , \7168 , \1028 );
and \U$6854 ( \7837 , \6825 , \1026 );
nor \U$6855 ( \7838 , \7836 , \7837 );
xnor \U$6856 ( \7839 , \7838 , \1009 );
and \U$6857 ( \7840 , \7673 , \991 );
and \U$6858 ( \7841 , \7370 , \989 );
nor \U$6859 ( \7842 , \7840 , \7841 );
xnor \U$6860 ( \7843 , \7842 , \996 );
and \U$6861 ( \7844 , \7839 , \7843 );
buf \U$6862 ( \7845 , RIc0dac60_116);
and \U$6863 ( \7846 , \7845 , \985 );
and \U$6864 ( \7847 , \7843 , \7846 );
and \U$6865 ( \7848 , \7839 , \7846 );
or \U$6866 ( \7849 , \7844 , \7847 , \7848 );
and \U$6867 ( \7850 , \7835 , \7849 );
and \U$6868 ( \7851 , \5916 , \1247 );
and \U$6869 ( \7852 , \5447 , \1245 );
nor \U$6870 ( \7853 , \7851 , \7852 );
xnor \U$6871 ( \7854 , \7853 , \1198 );
and \U$6872 ( \7855 , \6185 , \1146 );
and \U$6873 ( \7856 , \5921 , \1144 );
nor \U$6874 ( \7857 , \7855 , \7856 );
xnor \U$6875 ( \7858 , \7857 , \1105 );
and \U$6876 ( \7859 , \7854 , \7858 );
and \U$6877 ( \7860 , \6816 , \1076 );
and \U$6878 ( \7861 , \6444 , \1074 );
nor \U$6879 ( \7862 , \7860 , \7861 );
xnor \U$6880 ( \7863 , \7862 , \1046 );
and \U$6881 ( \7864 , \7858 , \7863 );
and \U$6882 ( \7865 , \7854 , \7863 );
or \U$6883 ( \7866 , \7859 , \7864 , \7865 );
and \U$6884 ( \7867 , \7849 , \7866 );
and \U$6885 ( \7868 , \7835 , \7866 );
or \U$6886 ( \7869 , \7850 , \7867 , \7868 );
and \U$6887 ( \7870 , \1162 , \6314 );
and \U$6888 ( \7871 , \1093 , \6312 );
nor \U$6889 ( \7872 , \7870 , \7871 );
xnor \U$6890 ( \7873 , \7872 , \6073 );
and \U$6891 ( \7874 , \1221 , \5848 );
and \U$6892 ( \7875 , \1167 , \5846 );
nor \U$6893 ( \7876 , \7874 , \7875 );
xnor \U$6894 ( \7877 , \7876 , \5660 );
and \U$6895 ( \7878 , \7873 , \7877 );
and \U$6896 ( \7879 , \1349 , \5474 );
and \U$6897 ( \7880 , \1272 , \5472 );
nor \U$6898 ( \7881 , \7879 , \7880 );
xnor \U$6899 ( \7882 , \7881 , \5242 );
and \U$6900 ( \7883 , \7877 , \7882 );
and \U$6901 ( \7884 , \7873 , \7882 );
or \U$6902 ( \7885 , \7878 , \7883 , \7884 );
and \U$6903 ( \7886 , \1457 , \5023 );
and \U$6904 ( \7887 , \1377 , \5021 );
nor \U$6905 ( \7888 , \7886 , \7887 );
xnor \U$6906 ( \7889 , \7888 , \4880 );
and \U$6907 ( \7890 , \1593 , \4700 );
and \U$6908 ( \7891 , \1531 , \4698 );
nor \U$6909 ( \7892 , \7890 , \7891 );
xnor \U$6910 ( \7893 , \7892 , \4454 );
and \U$6911 ( \7894 , \7889 , \7893 );
and \U$6912 ( \7895 , \1854 , \4305 );
and \U$6913 ( \7896 , \1656 , \4303 );
nor \U$6914 ( \7897 , \7895 , \7896 );
xnor \U$6915 ( \7898 , \7897 , \4118 );
and \U$6916 ( \7899 , \7893 , \7898 );
and \U$6917 ( \7900 , \7889 , \7898 );
or \U$6918 ( \7901 , \7894 , \7899 , \7900 );
and \U$6919 ( \7902 , \7885 , \7901 );
xor \U$6920 ( \7903 , \7094 , \7642 );
xor \U$6921 ( \7904 , \7642 , \7643 );
not \U$6922 ( \7905 , \7904 );
and \U$6923 ( \7906 , \7903 , \7905 );
and \U$6924 ( \7907 , \984 , \7906 );
not \U$6925 ( \7908 , \7907 );
xnor \U$6926 ( \7909 , \7908 , \7646 );
and \U$6927 ( \7910 , \1016 , \7412 );
and \U$6928 ( \7911 , \998 , \7410 );
nor \U$6929 ( \7912 , \7910 , \7911 );
xnor \U$6930 ( \7913 , \7912 , \7097 );
and \U$6931 ( \7914 , \7909 , \7913 );
and \U$6932 ( \7915 , \1085 , \6903 );
and \U$6933 ( \7916 , \1037 , \6901 );
nor \U$6934 ( \7917 , \7915 , \7916 );
xnor \U$6935 ( \7918 , \7917 , \6563 );
and \U$6936 ( \7919 , \7913 , \7918 );
and \U$6937 ( \7920 , \7909 , \7918 );
or \U$6938 ( \7921 , \7914 , \7919 , \7920 );
and \U$6939 ( \7922 , \7901 , \7921 );
and \U$6940 ( \7923 , \7885 , \7921 );
or \U$6941 ( \7924 , \7902 , \7922 , \7923 );
and \U$6942 ( \7925 , \7869 , \7924 );
and \U$6943 ( \7926 , \2047 , \3992 );
and \U$6944 ( \7927 , \1942 , \3990 );
nor \U$6945 ( \7928 , \7926 , \7927 );
xnor \U$6946 ( \7929 , \7928 , \3787 );
and \U$6947 ( \7930 , \2168 , \3586 );
and \U$6948 ( \7931 , \2052 , \3584 );
nor \U$6949 ( \7932 , \7930 , \7931 );
xnor \U$6950 ( \7933 , \7932 , \3437 );
and \U$6951 ( \7934 , \7929 , \7933 );
and \U$6952 ( \7935 , \2459 , \3264 );
and \U$6953 ( \7936 , \2283 , \3262 );
nor \U$6954 ( \7937 , \7935 , \7936 );
xnor \U$6955 ( \7938 , \7937 , \3122 );
and \U$6956 ( \7939 , \7933 , \7938 );
and \U$6957 ( \7940 , \7929 , \7938 );
or \U$6958 ( \7941 , \7934 , \7939 , \7940 );
and \U$6959 ( \7942 , \2710 , \2968 );
and \U$6960 ( \7943 , \2467 , \2966 );
nor \U$6961 ( \7944 , \7942 , \7943 );
xnor \U$6962 ( \7945 , \7944 , \2831 );
and \U$6963 ( \7946 , \2901 , \2762 );
and \U$6964 ( \7947 , \2715 , \2760 );
nor \U$6965 ( \7948 , \7946 , \7947 );
xnor \U$6966 ( \7949 , \7948 , \2610 );
and \U$6967 ( \7950 , \7945 , \7949 );
and \U$6968 ( \7951 , \3309 , \2494 );
and \U$6969 ( \7952 , \3045 , \2492 );
nor \U$6970 ( \7953 , \7951 , \7952 );
xnor \U$6971 ( \7954 , \7953 , \2338 );
and \U$6972 ( \7955 , \7949 , \7954 );
and \U$6973 ( \7956 , \7945 , \7954 );
or \U$6974 ( \7957 , \7950 , \7955 , \7956 );
and \U$6975 ( \7958 , \7941 , \7957 );
and \U$6976 ( \7959 , \3508 , \2222 );
and \U$6977 ( \7960 , \3334 , \2220 );
nor \U$6978 ( \7961 , \7959 , \7960 );
xnor \U$6979 ( \7962 , \7961 , \2109 );
and \U$6980 ( \7963 , \3813 , \2028 );
and \U$6981 ( \7964 , \3675 , \2026 );
nor \U$6982 ( \7965 , \7963 , \7964 );
xnor \U$6983 ( \7966 , \7965 , \1892 );
and \U$6984 ( \7967 , \7962 , \7966 );
and \U$6985 ( \7968 , \4349 , \1828 );
and \U$6986 ( \7969 , \3932 , \1826 );
nor \U$6987 ( \7970 , \7968 , \7969 );
xnor \U$6988 ( \7971 , \7970 , \1750 );
and \U$6989 ( \7972 , \7966 , \7971 );
and \U$6990 ( \7973 , \7962 , \7971 );
or \U$6991 ( \7974 , \7967 , \7972 , \7973 );
and \U$6992 ( \7975 , \7957 , \7974 );
and \U$6993 ( \7976 , \7941 , \7974 );
or \U$6994 ( \7977 , \7958 , \7975 , \7976 );
and \U$6995 ( \7978 , \7924 , \7977 );
and \U$6996 ( \7979 , \7869 , \7977 );
or \U$6997 ( \7980 , \7925 , \7978 , \7979 );
xor \U$6998 ( \7981 , \7667 , \7671 );
xor \U$6999 ( \7982 , \7981 , \7674 );
xor \U$7000 ( \7983 , \7681 , \7685 );
xor \U$7001 ( \7984 , \7983 , \7690 );
and \U$7002 ( \7985 , \7982 , \7984 );
xor \U$7003 ( \7986 , \7698 , \7702 );
xor \U$7004 ( \7987 , \7986 , \7707 );
and \U$7005 ( \7988 , \7984 , \7987 );
and \U$7006 ( \7989 , \7982 , \7987 );
or \U$7007 ( \7990 , \7985 , \7988 , \7989 );
xor \U$7008 ( \7991 , \7560 , \7564 );
xor \U$7009 ( \7992 , \7991 , \7569 );
xor \U$7010 ( \7993 , \7576 , \7580 );
xor \U$7011 ( \7994 , \7993 , \7585 );
and \U$7012 ( \7995 , \7992 , \7994 );
xor \U$7013 ( \7996 , \7593 , \7597 );
xor \U$7014 ( \7997 , \7996 , \7602 );
and \U$7015 ( \7998 , \7994 , \7997 );
and \U$7016 ( \7999 , \7992 , \7997 );
or \U$7017 ( \8000 , \7995 , \7998 , \7999 );
and \U$7018 ( \8001 , \7990 , \8000 );
xor \U$7019 ( \8002 , \7612 , \7616 );
xor \U$7020 ( \8003 , \8002 , \7621 );
xor \U$7021 ( \8004 , \7628 , \7632 );
xor \U$7022 ( \8005 , \8004 , \7637 );
and \U$7023 ( \8006 , \8003 , \8005 );
xor \U$7024 ( \8007 , \7647 , \7651 );
xor \U$7025 ( \8008 , \8007 , \7656 );
and \U$7026 ( \8009 , \8005 , \8008 );
and \U$7027 ( \8010 , \8003 , \8008 );
or \U$7028 ( \8011 , \8006 , \8009 , \8010 );
and \U$7029 ( \8012 , \8000 , \8011 );
and \U$7030 ( \8013 , \7990 , \8011 );
or \U$7031 ( \8014 , \8001 , \8012 , \8013 );
and \U$7032 ( \8015 , \7980 , \8014 );
xor \U$7033 ( \8016 , \7718 , \7720 );
xor \U$7034 ( \8017 , \8016 , \7723 );
xor \U$7035 ( \8018 , \7728 , \7730 );
xor \U$7036 ( \8019 , \8018 , \7733 );
and \U$7037 ( \8020 , \8017 , \8019 );
xor \U$7038 ( \8021 , \7739 , \7741 );
xor \U$7039 ( \8022 , \8021 , \7743 );
and \U$7040 ( \8023 , \8019 , \8022 );
and \U$7041 ( \8024 , \8017 , \8022 );
or \U$7042 ( \8025 , \8020 , \8023 , \8024 );
and \U$7043 ( \8026 , \8014 , \8025 );
and \U$7044 ( \8027 , \7980 , \8025 );
or \U$7045 ( \8028 , \8015 , \8026 , \8027 );
xor \U$7046 ( \8029 , \7572 , \7588 );
xor \U$7047 ( \8030 , \8029 , \7605 );
xor \U$7048 ( \8031 , \7624 , \7640 );
xor \U$7049 ( \8032 , \8031 , \7659 );
and \U$7050 ( \8033 , \8030 , \8032 );
xor \U$7051 ( \8034 , \7677 , \7693 );
xor \U$7052 ( \8035 , \8034 , \7710 );
and \U$7053 ( \8036 , \8032 , \8035 );
and \U$7054 ( \8037 , \8030 , \8035 );
or \U$7055 ( \8038 , \8033 , \8036 , \8037 );
xor \U$7056 ( \8039 , \7765 , \7767 );
xor \U$7057 ( \8040 , \8039 , \7770 );
and \U$7058 ( \8041 , \8038 , \8040 );
xor \U$7059 ( \8042 , \7752 , \7754 );
xor \U$7060 ( \8043 , \8042 , \7757 );
and \U$7061 ( \8044 , \8040 , \8043 );
and \U$7062 ( \8045 , \8038 , \8043 );
or \U$7063 ( \8046 , \8041 , \8044 , \8045 );
and \U$7064 ( \8047 , \8028 , \8046 );
xor \U$7065 ( \8048 , \7608 , \7662 );
xor \U$7066 ( \8049 , \8048 , \7713 );
xor \U$7067 ( \8050 , \7726 , \7736 );
xor \U$7068 ( \8051 , \8050 , \7746 );
and \U$7069 ( \8052 , \8049 , \8051 );
and \U$7070 ( \8053 , \8046 , \8052 );
and \U$7071 ( \8054 , \8028 , \8052 );
or \U$7072 ( \8055 , \8047 , \8053 , \8054 );
xor \U$7073 ( \8056 , \7716 , \7749 );
xor \U$7074 ( \8057 , \8056 , \7760 );
xor \U$7075 ( \8058 , \7773 , \7775 );
xor \U$7076 ( \8059 , \8058 , \7778 );
and \U$7077 ( \8060 , \8057 , \8059 );
xor \U$7078 ( \8061 , \7784 , \7786 );
and \U$7079 ( \8062 , \8059 , \8061 );
and \U$7080 ( \8063 , \8057 , \8061 );
or \U$7081 ( \8064 , \8060 , \8062 , \8063 );
and \U$7082 ( \8065 , \8055 , \8064 );
xor \U$7083 ( \8066 , \7792 , \7794 );
xor \U$7084 ( \8067 , \8066 , \7796 );
and \U$7085 ( \8068 , \8064 , \8067 );
and \U$7086 ( \8069 , \8055 , \8067 );
or \U$7087 ( \8070 , \8065 , \8068 , \8069 );
xor \U$7088 ( \8071 , \7500 , \7518 );
xor \U$7089 ( \8072 , \8071 , \7524 );
and \U$7090 ( \8073 , \8070 , \8072 );
xor \U$7091 ( \8074 , \7790 , \7799 );
xor \U$7092 ( \8075 , \8074 , \7802 );
and \U$7093 ( \8076 , \8072 , \8075 );
and \U$7094 ( \8077 , \8070 , \8075 );
or \U$7095 ( \8078 , \8073 , \8076 , \8077 );
xor \U$7096 ( \8079 , \7805 , \7807 );
xor \U$7097 ( \8080 , \8079 , \7810 );
and \U$7098 ( \8081 , \8078 , \8080 );
and \U$7099 ( \8082 , \7819 , \8081 );
xor \U$7100 ( \8083 , \7819 , \8081 );
xor \U$7101 ( \8084 , \8078 , \8080 );
xor \U$7102 ( \8085 , \7873 , \7877 );
xor \U$7103 ( \8086 , \8085 , \7882 );
xor \U$7104 ( \8087 , \7929 , \7933 );
xor \U$7105 ( \8088 , \8087 , \7938 );
and \U$7106 ( \8089 , \8086 , \8088 );
xor \U$7107 ( \8090 , \7889 , \7893 );
xor \U$7108 ( \8091 , \8090 , \7898 );
and \U$7109 ( \8092 , \8088 , \8091 );
and \U$7110 ( \8093 , \8086 , \8091 );
or \U$7111 ( \8094 , \8089 , \8092 , \8093 );
xor \U$7112 ( \8095 , \7945 , \7949 );
xor \U$7113 ( \8096 , \8095 , \7954 );
xor \U$7114 ( \8097 , \7823 , \7827 );
xor \U$7115 ( \8098 , \8097 , \7832 );
and \U$7116 ( \8099 , \8096 , \8098 );
xor \U$7117 ( \8100 , \7962 , \7966 );
xor \U$7118 ( \8101 , \8100 , \7971 );
and \U$7119 ( \8102 , \8098 , \8101 );
and \U$7120 ( \8103 , \8096 , \8101 );
or \U$7121 ( \8104 , \8099 , \8102 , \8103 );
and \U$7122 ( \8105 , \8094 , \8104 );
xor \U$7123 ( \8106 , \7839 , \7843 );
xor \U$7124 ( \8107 , \8106 , \7846 );
xor \U$7125 ( \8108 , \7854 , \7858 );
xor \U$7126 ( \8109 , \8108 , \7863 );
or \U$7127 ( \8110 , \8107 , \8109 );
and \U$7128 ( \8111 , \8104 , \8110 );
and \U$7129 ( \8112 , \8094 , \8110 );
or \U$7130 ( \8113 , \8105 , \8111 , \8112 );
and \U$7131 ( \8114 , \2467 , \3264 );
and \U$7132 ( \8115 , \2459 , \3262 );
nor \U$7133 ( \8116 , \8114 , \8115 );
xnor \U$7134 ( \8117 , \8116 , \3122 );
and \U$7135 ( \8118 , \2715 , \2968 );
and \U$7136 ( \8119 , \2710 , \2966 );
nor \U$7137 ( \8120 , \8118 , \8119 );
xnor \U$7138 ( \8121 , \8120 , \2831 );
and \U$7139 ( \8122 , \8117 , \8121 );
and \U$7140 ( \8123 , \3045 , \2762 );
and \U$7141 ( \8124 , \2901 , \2760 );
nor \U$7142 ( \8125 , \8123 , \8124 );
xnor \U$7143 ( \8126 , \8125 , \2610 );
and \U$7144 ( \8127 , \8121 , \8126 );
and \U$7145 ( \8128 , \8117 , \8126 );
or \U$7146 ( \8129 , \8122 , \8127 , \8128 );
and \U$7147 ( \8130 , \1942 , \4305 );
and \U$7148 ( \8131 , \1854 , \4303 );
nor \U$7149 ( \8132 , \8130 , \8131 );
xnor \U$7150 ( \8133 , \8132 , \4118 );
and \U$7151 ( \8134 , \2052 , \3992 );
and \U$7152 ( \8135 , \2047 , \3990 );
nor \U$7153 ( \8136 , \8134 , \8135 );
xnor \U$7154 ( \8137 , \8136 , \3787 );
and \U$7155 ( \8138 , \8133 , \8137 );
and \U$7156 ( \8139 , \2283 , \3586 );
and \U$7157 ( \8140 , \2168 , \3584 );
nor \U$7158 ( \8141 , \8139 , \8140 );
xnor \U$7159 ( \8142 , \8141 , \3437 );
and \U$7160 ( \8143 , \8137 , \8142 );
and \U$7161 ( \8144 , \8133 , \8142 );
or \U$7162 ( \8145 , \8138 , \8143 , \8144 );
and \U$7163 ( \8146 , \8129 , \8145 );
and \U$7164 ( \8147 , \3334 , \2494 );
and \U$7165 ( \8148 , \3309 , \2492 );
nor \U$7166 ( \8149 , \8147 , \8148 );
xnor \U$7167 ( \8150 , \8149 , \2338 );
and \U$7168 ( \8151 , \3675 , \2222 );
and \U$7169 ( \8152 , \3508 , \2220 );
nor \U$7170 ( \8153 , \8151 , \8152 );
xnor \U$7171 ( \8154 , \8153 , \2109 );
and \U$7172 ( \8155 , \8150 , \8154 );
and \U$7173 ( \8156 , \3932 , \2028 );
and \U$7174 ( \8157 , \3813 , \2026 );
nor \U$7175 ( \8158 , \8156 , \8157 );
xnor \U$7176 ( \8159 , \8158 , \1892 );
and \U$7177 ( \8160 , \8154 , \8159 );
and \U$7178 ( \8161 , \8150 , \8159 );
or \U$7179 ( \8162 , \8155 , \8160 , \8161 );
and \U$7180 ( \8163 , \8145 , \8162 );
and \U$7181 ( \8164 , \8129 , \8162 );
or \U$7182 ( \8165 , \8146 , \8163 , \8164 );
and \U$7183 ( \8166 , \1093 , \6903 );
and \U$7184 ( \8167 , \1085 , \6901 );
nor \U$7185 ( \8168 , \8166 , \8167 );
xnor \U$7186 ( \8169 , \8168 , \6563 );
and \U$7187 ( \8170 , \1167 , \6314 );
and \U$7188 ( \8171 , \1162 , \6312 );
nor \U$7189 ( \8172 , \8170 , \8171 );
xnor \U$7190 ( \8173 , \8172 , \6073 );
and \U$7191 ( \8174 , \8169 , \8173 );
and \U$7192 ( \8175 , \1272 , \5848 );
and \U$7193 ( \8176 , \1221 , \5846 );
nor \U$7194 ( \8177 , \8175 , \8176 );
xnor \U$7195 ( \8178 , \8177 , \5660 );
and \U$7196 ( \8179 , \8173 , \8178 );
and \U$7197 ( \8180 , \8169 , \8178 );
or \U$7198 ( \8181 , \8174 , \8179 , \8180 );
buf \U$7199 ( \8182 , RIc0d8f50_54);
buf \U$7200 ( \8183 , RIc0d8fc8_55);
and \U$7201 ( \8184 , \8182 , \8183 );
not \U$7202 ( \8185 , \8184 );
and \U$7203 ( \8186 , \7643 , \8185 );
not \U$7204 ( \8187 , \8186 );
and \U$7205 ( \8188 , \998 , \7906 );
and \U$7206 ( \8189 , \984 , \7904 );
nor \U$7207 ( \8190 , \8188 , \8189 );
xnor \U$7208 ( \8191 , \8190 , \7646 );
and \U$7209 ( \8192 , \8187 , \8191 );
and \U$7210 ( \8193 , \1037 , \7412 );
and \U$7211 ( \8194 , \1016 , \7410 );
nor \U$7212 ( \8195 , \8193 , \8194 );
xnor \U$7213 ( \8196 , \8195 , \7097 );
and \U$7214 ( \8197 , \8191 , \8196 );
and \U$7215 ( \8198 , \8187 , \8196 );
or \U$7216 ( \8199 , \8192 , \8197 , \8198 );
and \U$7217 ( \8200 , \8181 , \8199 );
and \U$7218 ( \8201 , \1377 , \5474 );
and \U$7219 ( \8202 , \1349 , \5472 );
nor \U$7220 ( \8203 , \8201 , \8202 );
xnor \U$7221 ( \8204 , \8203 , \5242 );
and \U$7222 ( \8205 , \1531 , \5023 );
and \U$7223 ( \8206 , \1457 , \5021 );
nor \U$7224 ( \8207 , \8205 , \8206 );
xnor \U$7225 ( \8208 , \8207 , \4880 );
and \U$7226 ( \8209 , \8204 , \8208 );
and \U$7227 ( \8210 , \1656 , \4700 );
and \U$7228 ( \8211 , \1593 , \4698 );
nor \U$7229 ( \8212 , \8210 , \8211 );
xnor \U$7230 ( \8213 , \8212 , \4454 );
and \U$7231 ( \8214 , \8208 , \8213 );
and \U$7232 ( \8215 , \8204 , \8213 );
or \U$7233 ( \8216 , \8209 , \8214 , \8215 );
and \U$7234 ( \8217 , \8199 , \8216 );
and \U$7235 ( \8218 , \8181 , \8216 );
or \U$7236 ( \8219 , \8200 , \8217 , \8218 );
and \U$7237 ( \8220 , \8165 , \8219 );
and \U$7238 ( \8221 , \4557 , \1828 );
and \U$7239 ( \8222 , \4349 , \1826 );
nor \U$7240 ( \8223 , \8221 , \8222 );
xnor \U$7241 ( \8224 , \8223 , \1750 );
and \U$7242 ( \8225 , \4684 , \1664 );
and \U$7243 ( \8226 , \4679 , \1662 );
nor \U$7244 ( \8227 , \8225 , \8226 );
xnor \U$7245 ( \8228 , \8227 , \1570 );
and \U$7246 ( \8229 , \8224 , \8228 );
and \U$7247 ( \8230 , \5137 , \1494 );
and \U$7248 ( \8231 , \4940 , \1492 );
nor \U$7249 ( \8232 , \8230 , \8231 );
xnor \U$7250 ( \8233 , \8232 , \1422 );
and \U$7251 ( \8234 , \8228 , \8233 );
and \U$7252 ( \8235 , \8224 , \8233 );
or \U$7253 ( \8236 , \8229 , \8234 , \8235 );
and \U$7254 ( \8237 , \5447 , \1360 );
and \U$7255 ( \8238 , \5439 , \1358 );
nor \U$7256 ( \8239 , \8237 , \8238 );
xnor \U$7257 ( \8240 , \8239 , \1317 );
and \U$7258 ( \8241 , \5921 , \1247 );
and \U$7259 ( \8242 , \5916 , \1245 );
nor \U$7260 ( \8243 , \8241 , \8242 );
xnor \U$7261 ( \8244 , \8243 , \1198 );
and \U$7262 ( \8245 , \8240 , \8244 );
and \U$7263 ( \8246 , \6444 , \1146 );
and \U$7264 ( \8247 , \6185 , \1144 );
nor \U$7265 ( \8248 , \8246 , \8247 );
xnor \U$7266 ( \8249 , \8248 , \1105 );
and \U$7267 ( \8250 , \8244 , \8249 );
and \U$7268 ( \8251 , \8240 , \8249 );
or \U$7269 ( \8252 , \8245 , \8250 , \8251 );
and \U$7270 ( \8253 , \8236 , \8252 );
and \U$7271 ( \8254 , \6825 , \1076 );
and \U$7272 ( \8255 , \6816 , \1074 );
nor \U$7273 ( \8256 , \8254 , \8255 );
xnor \U$7274 ( \8257 , \8256 , \1046 );
and \U$7275 ( \8258 , \7370 , \1028 );
and \U$7276 ( \8259 , \7168 , \1026 );
nor \U$7277 ( \8260 , \8258 , \8259 );
xnor \U$7278 ( \8261 , \8260 , \1009 );
and \U$7279 ( \8262 , \8257 , \8261 );
and \U$7280 ( \8263 , \7845 , \991 );
and \U$7281 ( \8264 , \7673 , \989 );
nor \U$7282 ( \8265 , \8263 , \8264 );
xnor \U$7283 ( \8266 , \8265 , \996 );
and \U$7284 ( \8267 , \8261 , \8266 );
and \U$7285 ( \8268 , \8257 , \8266 );
or \U$7286 ( \8269 , \8262 , \8267 , \8268 );
and \U$7287 ( \8270 , \8252 , \8269 );
and \U$7288 ( \8271 , \8236 , \8269 );
or \U$7289 ( \8272 , \8253 , \8270 , \8271 );
and \U$7290 ( \8273 , \8219 , \8272 );
and \U$7291 ( \8274 , \8165 , \8272 );
or \U$7292 ( \8275 , \8220 , \8273 , \8274 );
and \U$7293 ( \8276 , \8113 , \8275 );
xor \U$7294 ( \8277 , \7982 , \7984 );
xor \U$7295 ( \8278 , \8277 , \7987 );
xor \U$7296 ( \8279 , \7992 , \7994 );
xor \U$7297 ( \8280 , \8279 , \7997 );
and \U$7298 ( \8281 , \8278 , \8280 );
xor \U$7299 ( \8282 , \8003 , \8005 );
xor \U$7300 ( \8283 , \8282 , \8008 );
and \U$7301 ( \8284 , \8280 , \8283 );
and \U$7302 ( \8285 , \8278 , \8283 );
or \U$7303 ( \8286 , \8281 , \8284 , \8285 );
and \U$7304 ( \8287 , \8275 , \8286 );
and \U$7305 ( \8288 , \8113 , \8286 );
or \U$7306 ( \8289 , \8276 , \8287 , \8288 );
xor \U$7307 ( \8290 , \7835 , \7849 );
xor \U$7308 ( \8291 , \8290 , \7866 );
xor \U$7309 ( \8292 , \7885 , \7901 );
xor \U$7310 ( \8293 , \8292 , \7921 );
and \U$7311 ( \8294 , \8291 , \8293 );
xor \U$7312 ( \8295 , \7941 , \7957 );
xor \U$7313 ( \8296 , \8295 , \7974 );
and \U$7314 ( \8297 , \8293 , \8296 );
and \U$7315 ( \8298 , \8291 , \8296 );
or \U$7316 ( \8299 , \8294 , \8297 , \8298 );
xor \U$7317 ( \8300 , \8030 , \8032 );
xor \U$7318 ( \8301 , \8300 , \8035 );
and \U$7319 ( \8302 , \8299 , \8301 );
xor \U$7320 ( \8303 , \8017 , \8019 );
xor \U$7321 ( \8304 , \8303 , \8022 );
and \U$7322 ( \8305 , \8301 , \8304 );
and \U$7323 ( \8306 , \8299 , \8304 );
or \U$7324 ( \8307 , \8302 , \8305 , \8306 );
and \U$7325 ( \8308 , \8289 , \8307 );
xor \U$7326 ( \8309 , \7869 , \7924 );
xor \U$7327 ( \8310 , \8309 , \7977 );
xor \U$7328 ( \8311 , \7990 , \8000 );
xor \U$7329 ( \8312 , \8311 , \8011 );
and \U$7330 ( \8313 , \8310 , \8312 );
and \U$7331 ( \8314 , \8307 , \8313 );
and \U$7332 ( \8315 , \8289 , \8313 );
or \U$7333 ( \8316 , \8308 , \8314 , \8315 );
xor \U$7334 ( \8317 , \7980 , \8014 );
xor \U$7335 ( \8318 , \8317 , \8025 );
xor \U$7336 ( \8319 , \8038 , \8040 );
xor \U$7337 ( \8320 , \8319 , \8043 );
and \U$7338 ( \8321 , \8318 , \8320 );
xor \U$7339 ( \8322 , \8049 , \8051 );
and \U$7340 ( \8323 , \8320 , \8322 );
and \U$7341 ( \8324 , \8318 , \8322 );
or \U$7342 ( \8325 , \8321 , \8323 , \8324 );
and \U$7343 ( \8326 , \8316 , \8325 );
xor \U$7344 ( \8327 , \8057 , \8059 );
xor \U$7345 ( \8328 , \8327 , \8061 );
and \U$7346 ( \8329 , \8325 , \8328 );
and \U$7347 ( \8330 , \8316 , \8328 );
or \U$7348 ( \8331 , \8326 , \8329 , \8330 );
xor \U$7349 ( \8332 , \7763 , \7781 );
xor \U$7350 ( \8333 , \8332 , \7787 );
and \U$7351 ( \8334 , \8331 , \8333 );
xor \U$7352 ( \8335 , \8055 , \8064 );
xor \U$7353 ( \8336 , \8335 , \8067 );
and \U$7354 ( \8337 , \8333 , \8336 );
and \U$7355 ( \8338 , \8331 , \8336 );
or \U$7356 ( \8339 , \8334 , \8337 , \8338 );
xor \U$7357 ( \8340 , \8070 , \8072 );
xor \U$7358 ( \8341 , \8340 , \8075 );
and \U$7359 ( \8342 , \8339 , \8341 );
and \U$7360 ( \8343 , \8084 , \8342 );
xor \U$7361 ( \8344 , \8084 , \8342 );
xor \U$7362 ( \8345 , \8339 , \8341 );
and \U$7363 ( \8346 , \4679 , \1828 );
and \U$7364 ( \8347 , \4557 , \1826 );
nor \U$7365 ( \8348 , \8346 , \8347 );
xnor \U$7366 ( \8349 , \8348 , \1750 );
and \U$7367 ( \8350 , \4940 , \1664 );
and \U$7368 ( \8351 , \4684 , \1662 );
nor \U$7369 ( \8352 , \8350 , \8351 );
xnor \U$7370 ( \8353 , \8352 , \1570 );
and \U$7371 ( \8354 , \8349 , \8353 );
and \U$7372 ( \8355 , \5439 , \1494 );
and \U$7373 ( \8356 , \5137 , \1492 );
nor \U$7374 ( \8357 , \8355 , \8356 );
xnor \U$7375 ( \8358 , \8357 , \1422 );
and \U$7376 ( \8359 , \8353 , \8358 );
and \U$7377 ( \8360 , \8349 , \8358 );
or \U$7378 ( \8361 , \8354 , \8359 , \8360 );
and \U$7379 ( \8362 , \7168 , \1076 );
and \U$7380 ( \8363 , \6825 , \1074 );
nor \U$7381 ( \8364 , \8362 , \8363 );
xnor \U$7382 ( \8365 , \8364 , \1046 );
and \U$7383 ( \8366 , \7673 , \1028 );
and \U$7384 ( \8367 , \7370 , \1026 );
nor \U$7385 ( \8368 , \8366 , \8367 );
xnor \U$7386 ( \8369 , \8368 , \1009 );
and \U$7387 ( \8370 , \8365 , \8369 );
buf \U$7388 ( \8371 , RIc0dacd8_117);
and \U$7389 ( \8372 , \8371 , \991 );
and \U$7390 ( \8373 , \7845 , \989 );
nor \U$7391 ( \8374 , \8372 , \8373 );
xnor \U$7392 ( \8375 , \8374 , \996 );
and \U$7393 ( \8376 , \8369 , \8375 );
and \U$7394 ( \8377 , \8365 , \8375 );
or \U$7395 ( \8378 , \8370 , \8376 , \8377 );
and \U$7396 ( \8379 , \8361 , \8378 );
and \U$7397 ( \8380 , \5916 , \1360 );
and \U$7398 ( \8381 , \5447 , \1358 );
nor \U$7399 ( \8382 , \8380 , \8381 );
xnor \U$7400 ( \8383 , \8382 , \1317 );
and \U$7401 ( \8384 , \6185 , \1247 );
and \U$7402 ( \8385 , \5921 , \1245 );
nor \U$7403 ( \8386 , \8384 , \8385 );
xnor \U$7404 ( \8387 , \8386 , \1198 );
and \U$7405 ( \8388 , \8383 , \8387 );
and \U$7406 ( \8389 , \6816 , \1146 );
and \U$7407 ( \8390 , \6444 , \1144 );
nor \U$7408 ( \8391 , \8389 , \8390 );
xnor \U$7409 ( \8392 , \8391 , \1105 );
and \U$7410 ( \8393 , \8387 , \8392 );
and \U$7411 ( \8394 , \8383 , \8392 );
or \U$7412 ( \8395 , \8388 , \8393 , \8394 );
and \U$7413 ( \8396 , \8378 , \8395 );
and \U$7414 ( \8397 , \8361 , \8395 );
or \U$7415 ( \8398 , \8379 , \8396 , \8397 );
and \U$7416 ( \8399 , \1162 , \6903 );
and \U$7417 ( \8400 , \1093 , \6901 );
nor \U$7418 ( \8401 , \8399 , \8400 );
xnor \U$7419 ( \8402 , \8401 , \6563 );
and \U$7420 ( \8403 , \1221 , \6314 );
and \U$7421 ( \8404 , \1167 , \6312 );
nor \U$7422 ( \8405 , \8403 , \8404 );
xnor \U$7423 ( \8406 , \8405 , \6073 );
and \U$7424 ( \8407 , \8402 , \8406 );
and \U$7425 ( \8408 , \1349 , \5848 );
and \U$7426 ( \8409 , \1272 , \5846 );
nor \U$7427 ( \8410 , \8408 , \8409 );
xnor \U$7428 ( \8411 , \8410 , \5660 );
and \U$7429 ( \8412 , \8406 , \8411 );
and \U$7430 ( \8413 , \8402 , \8411 );
or \U$7431 ( \8414 , \8407 , \8412 , \8413 );
and \U$7432 ( \8415 , \1457 , \5474 );
and \U$7433 ( \8416 , \1377 , \5472 );
nor \U$7434 ( \8417 , \8415 , \8416 );
xnor \U$7435 ( \8418 , \8417 , \5242 );
and \U$7436 ( \8419 , \1593 , \5023 );
and \U$7437 ( \8420 , \1531 , \5021 );
nor \U$7438 ( \8421 , \8419 , \8420 );
xnor \U$7439 ( \8422 , \8421 , \4880 );
and \U$7440 ( \8423 , \8418 , \8422 );
and \U$7441 ( \8424 , \1854 , \4700 );
and \U$7442 ( \8425 , \1656 , \4698 );
nor \U$7443 ( \8426 , \8424 , \8425 );
xnor \U$7444 ( \8427 , \8426 , \4454 );
and \U$7445 ( \8428 , \8422 , \8427 );
and \U$7446 ( \8429 , \8418 , \8427 );
or \U$7447 ( \8430 , \8423 , \8428 , \8429 );
and \U$7448 ( \8431 , \8414 , \8430 );
xor \U$7449 ( \8432 , \7643 , \8182 );
xor \U$7450 ( \8433 , \8182 , \8183 );
not \U$7451 ( \8434 , \8433 );
and \U$7452 ( \8435 , \8432 , \8434 );
and \U$7453 ( \8436 , \984 , \8435 );
not \U$7454 ( \8437 , \8436 );
xnor \U$7455 ( \8438 , \8437 , \8186 );
and \U$7456 ( \8439 , \1016 , \7906 );
and \U$7457 ( \8440 , \998 , \7904 );
nor \U$7458 ( \8441 , \8439 , \8440 );
xnor \U$7459 ( \8442 , \8441 , \7646 );
and \U$7460 ( \8443 , \8438 , \8442 );
and \U$7461 ( \8444 , \1085 , \7412 );
and \U$7462 ( \8445 , \1037 , \7410 );
nor \U$7463 ( \8446 , \8444 , \8445 );
xnor \U$7464 ( \8447 , \8446 , \7097 );
and \U$7465 ( \8448 , \8442 , \8447 );
and \U$7466 ( \8449 , \8438 , \8447 );
or \U$7467 ( \8450 , \8443 , \8448 , \8449 );
and \U$7468 ( \8451 , \8430 , \8450 );
and \U$7469 ( \8452 , \8414 , \8450 );
or \U$7470 ( \8453 , \8431 , \8451 , \8452 );
and \U$7471 ( \8454 , \8398 , \8453 );
and \U$7472 ( \8455 , \3508 , \2494 );
and \U$7473 ( \8456 , \3334 , \2492 );
nor \U$7474 ( \8457 , \8455 , \8456 );
xnor \U$7475 ( \8458 , \8457 , \2338 );
and \U$7476 ( \8459 , \3813 , \2222 );
and \U$7477 ( \8460 , \3675 , \2220 );
nor \U$7478 ( \8461 , \8459 , \8460 );
xnor \U$7479 ( \8462 , \8461 , \2109 );
and \U$7480 ( \8463 , \8458 , \8462 );
and \U$7481 ( \8464 , \4349 , \2028 );
and \U$7482 ( \8465 , \3932 , \2026 );
nor \U$7483 ( \8466 , \8464 , \8465 );
xnor \U$7484 ( \8467 , \8466 , \1892 );
and \U$7485 ( \8468 , \8462 , \8467 );
and \U$7486 ( \8469 , \8458 , \8467 );
or \U$7487 ( \8470 , \8463 , \8468 , \8469 );
and \U$7488 ( \8471 , \2047 , \4305 );
and \U$7489 ( \8472 , \1942 , \4303 );
nor \U$7490 ( \8473 , \8471 , \8472 );
xnor \U$7491 ( \8474 , \8473 , \4118 );
and \U$7492 ( \8475 , \2168 , \3992 );
and \U$7493 ( \8476 , \2052 , \3990 );
nor \U$7494 ( \8477 , \8475 , \8476 );
xnor \U$7495 ( \8478 , \8477 , \3787 );
and \U$7496 ( \8479 , \8474 , \8478 );
and \U$7497 ( \8480 , \2459 , \3586 );
and \U$7498 ( \8481 , \2283 , \3584 );
nor \U$7499 ( \8482 , \8480 , \8481 );
xnor \U$7500 ( \8483 , \8482 , \3437 );
and \U$7501 ( \8484 , \8478 , \8483 );
and \U$7502 ( \8485 , \8474 , \8483 );
or \U$7503 ( \8486 , \8479 , \8484 , \8485 );
and \U$7504 ( \8487 , \8470 , \8486 );
and \U$7505 ( \8488 , \2710 , \3264 );
and \U$7506 ( \8489 , \2467 , \3262 );
nor \U$7507 ( \8490 , \8488 , \8489 );
xnor \U$7508 ( \8491 , \8490 , \3122 );
and \U$7509 ( \8492 , \2901 , \2968 );
and \U$7510 ( \8493 , \2715 , \2966 );
nor \U$7511 ( \8494 , \8492 , \8493 );
xnor \U$7512 ( \8495 , \8494 , \2831 );
and \U$7513 ( \8496 , \8491 , \8495 );
and \U$7514 ( \8497 , \3309 , \2762 );
and \U$7515 ( \8498 , \3045 , \2760 );
nor \U$7516 ( \8499 , \8497 , \8498 );
xnor \U$7517 ( \8500 , \8499 , \2610 );
and \U$7518 ( \8501 , \8495 , \8500 );
and \U$7519 ( \8502 , \8491 , \8500 );
or \U$7520 ( \8503 , \8496 , \8501 , \8502 );
and \U$7521 ( \8504 , \8486 , \8503 );
and \U$7522 ( \8505 , \8470 , \8503 );
or \U$7523 ( \8506 , \8487 , \8504 , \8505 );
and \U$7524 ( \8507 , \8453 , \8506 );
and \U$7525 ( \8508 , \8398 , \8506 );
or \U$7526 ( \8509 , \8454 , \8507 , \8508 );
xor \U$7527 ( \8510 , \8169 , \8173 );
xor \U$7528 ( \8511 , \8510 , \8178 );
xor \U$7529 ( \8512 , \8133 , \8137 );
xor \U$7530 ( \8513 , \8512 , \8142 );
and \U$7531 ( \8514 , \8511 , \8513 );
xor \U$7532 ( \8515 , \8204 , \8208 );
xor \U$7533 ( \8516 , \8515 , \8213 );
and \U$7534 ( \8517 , \8513 , \8516 );
and \U$7535 ( \8518 , \8511 , \8516 );
or \U$7536 ( \8519 , \8514 , \8517 , \8518 );
and \U$7537 ( \8520 , \8371 , \985 );
xor \U$7538 ( \8521 , \8240 , \8244 );
xor \U$7539 ( \8522 , \8521 , \8249 );
and \U$7540 ( \8523 , \8520 , \8522 );
xor \U$7541 ( \8524 , \8257 , \8261 );
xor \U$7542 ( \8525 , \8524 , \8266 );
and \U$7543 ( \8526 , \8522 , \8525 );
and \U$7544 ( \8527 , \8520 , \8525 );
or \U$7545 ( \8528 , \8523 , \8526 , \8527 );
and \U$7546 ( \8529 , \8519 , \8528 );
xor \U$7547 ( \8530 , \8224 , \8228 );
xor \U$7548 ( \8531 , \8530 , \8233 );
xor \U$7549 ( \8532 , \8117 , \8121 );
xor \U$7550 ( \8533 , \8532 , \8126 );
and \U$7551 ( \8534 , \8531 , \8533 );
xor \U$7552 ( \8535 , \8150 , \8154 );
xor \U$7553 ( \8536 , \8535 , \8159 );
and \U$7554 ( \8537 , \8533 , \8536 );
and \U$7555 ( \8538 , \8531 , \8536 );
or \U$7556 ( \8539 , \8534 , \8537 , \8538 );
and \U$7557 ( \8540 , \8528 , \8539 );
and \U$7558 ( \8541 , \8519 , \8539 );
or \U$7559 ( \8542 , \8529 , \8540 , \8541 );
and \U$7560 ( \8543 , \8509 , \8542 );
xor \U$7561 ( \8544 , \7909 , \7913 );
xor \U$7562 ( \8545 , \8544 , \7918 );
xor \U$7563 ( \8546 , \8086 , \8088 );
xor \U$7564 ( \8547 , \8546 , \8091 );
and \U$7565 ( \8548 , \8545 , \8547 );
xor \U$7566 ( \8549 , \8096 , \8098 );
xor \U$7567 ( \8550 , \8549 , \8101 );
and \U$7568 ( \8551 , \8547 , \8550 );
and \U$7569 ( \8552 , \8545 , \8550 );
or \U$7570 ( \8553 , \8548 , \8551 , \8552 );
and \U$7571 ( \8554 , \8542 , \8553 );
and \U$7572 ( \8555 , \8509 , \8553 );
or \U$7573 ( \8556 , \8543 , \8554 , \8555 );
xor \U$7574 ( \8557 , \8129 , \8145 );
xor \U$7575 ( \8558 , \8557 , \8162 );
xor \U$7576 ( \8559 , \8236 , \8252 );
xor \U$7577 ( \8560 , \8559 , \8269 );
and \U$7578 ( \8561 , \8558 , \8560 );
xnor \U$7579 ( \8562 , \8107 , \8109 );
and \U$7580 ( \8563 , \8560 , \8562 );
and \U$7581 ( \8564 , \8558 , \8562 );
or \U$7582 ( \8565 , \8561 , \8563 , \8564 );
xor \U$7583 ( \8566 , \8291 , \8293 );
xor \U$7584 ( \8567 , \8566 , \8296 );
and \U$7585 ( \8568 , \8565 , \8567 );
xor \U$7586 ( \8569 , \8278 , \8280 );
xor \U$7587 ( \8570 , \8569 , \8283 );
and \U$7588 ( \8571 , \8567 , \8570 );
and \U$7589 ( \8572 , \8565 , \8570 );
or \U$7590 ( \8573 , \8568 , \8571 , \8572 );
and \U$7591 ( \8574 , \8556 , \8573 );
xor \U$7592 ( \8575 , \8094 , \8104 );
xor \U$7593 ( \8576 , \8575 , \8110 );
xor \U$7594 ( \8577 , \8165 , \8219 );
xor \U$7595 ( \8578 , \8577 , \8272 );
and \U$7596 ( \8579 , \8576 , \8578 );
and \U$7597 ( \8580 , \8573 , \8579 );
and \U$7598 ( \8581 , \8556 , \8579 );
or \U$7599 ( \8582 , \8574 , \8580 , \8581 );
xor \U$7600 ( \8583 , \8113 , \8275 );
xor \U$7601 ( \8584 , \8583 , \8286 );
xor \U$7602 ( \8585 , \8299 , \8301 );
xor \U$7603 ( \8586 , \8585 , \8304 );
and \U$7604 ( \8587 , \8584 , \8586 );
xor \U$7605 ( \8588 , \8310 , \8312 );
and \U$7606 ( \8589 , \8586 , \8588 );
and \U$7607 ( \8590 , \8584 , \8588 );
or \U$7608 ( \8591 , \8587 , \8589 , \8590 );
and \U$7609 ( \8592 , \8582 , \8591 );
xor \U$7610 ( \8593 , \8318 , \8320 );
xor \U$7611 ( \8594 , \8593 , \8322 );
and \U$7612 ( \8595 , \8591 , \8594 );
and \U$7613 ( \8596 , \8582 , \8594 );
or \U$7614 ( \8597 , \8592 , \8595 , \8596 );
xor \U$7615 ( \8598 , \8028 , \8046 );
xor \U$7616 ( \8599 , \8598 , \8052 );
and \U$7617 ( \8600 , \8597 , \8599 );
xor \U$7618 ( \8601 , \8316 , \8325 );
xor \U$7619 ( \8602 , \8601 , \8328 );
and \U$7620 ( \8603 , \8599 , \8602 );
and \U$7621 ( \8604 , \8597 , \8602 );
or \U$7622 ( \8605 , \8600 , \8603 , \8604 );
xor \U$7623 ( \8606 , \8331 , \8333 );
xor \U$7624 ( \8607 , \8606 , \8336 );
and \U$7625 ( \8608 , \8605 , \8607 );
and \U$7626 ( \8609 , \8345 , \8608 );
xor \U$7627 ( \8610 , \8345 , \8608 );
xor \U$7628 ( \8611 , \8605 , \8607 );
and \U$7629 ( \8612 , \3334 , \2762 );
and \U$7630 ( \8613 , \3309 , \2760 );
nor \U$7631 ( \8614 , \8612 , \8613 );
xnor \U$7632 ( \8615 , \8614 , \2610 );
and \U$7633 ( \8616 , \3675 , \2494 );
and \U$7634 ( \8617 , \3508 , \2492 );
nor \U$7635 ( \8618 , \8616 , \8617 );
xnor \U$7636 ( \8619 , \8618 , \2338 );
and \U$7637 ( \8620 , \8615 , \8619 );
and \U$7638 ( \8621 , \3932 , \2222 );
and \U$7639 ( \8622 , \3813 , \2220 );
nor \U$7640 ( \8623 , \8621 , \8622 );
xnor \U$7641 ( \8624 , \8623 , \2109 );
and \U$7642 ( \8625 , \8619 , \8624 );
and \U$7643 ( \8626 , \8615 , \8624 );
or \U$7644 ( \8627 , \8620 , \8625 , \8626 );
and \U$7645 ( \8628 , \1942 , \4700 );
and \U$7646 ( \8629 , \1854 , \4698 );
nor \U$7647 ( \8630 , \8628 , \8629 );
xnor \U$7648 ( \8631 , \8630 , \4454 );
and \U$7649 ( \8632 , \2052 , \4305 );
and \U$7650 ( \8633 , \2047 , \4303 );
nor \U$7651 ( \8634 , \8632 , \8633 );
xnor \U$7652 ( \8635 , \8634 , \4118 );
and \U$7653 ( \8636 , \8631 , \8635 );
and \U$7654 ( \8637 , \2283 , \3992 );
and \U$7655 ( \8638 , \2168 , \3990 );
nor \U$7656 ( \8639 , \8637 , \8638 );
xnor \U$7657 ( \8640 , \8639 , \3787 );
and \U$7658 ( \8641 , \8635 , \8640 );
and \U$7659 ( \8642 , \8631 , \8640 );
or \U$7660 ( \8643 , \8636 , \8641 , \8642 );
and \U$7661 ( \8644 , \8627 , \8643 );
and \U$7662 ( \8645 , \2467 , \3586 );
and \U$7663 ( \8646 , \2459 , \3584 );
nor \U$7664 ( \8647 , \8645 , \8646 );
xnor \U$7665 ( \8648 , \8647 , \3437 );
and \U$7666 ( \8649 , \2715 , \3264 );
and \U$7667 ( \8650 , \2710 , \3262 );
nor \U$7668 ( \8651 , \8649 , \8650 );
xnor \U$7669 ( \8652 , \8651 , \3122 );
and \U$7670 ( \8653 , \8648 , \8652 );
and \U$7671 ( \8654 , \3045 , \2968 );
and \U$7672 ( \8655 , \2901 , \2966 );
nor \U$7673 ( \8656 , \8654 , \8655 );
xnor \U$7674 ( \8657 , \8656 , \2831 );
and \U$7675 ( \8658 , \8652 , \8657 );
and \U$7676 ( \8659 , \8648 , \8657 );
or \U$7677 ( \8660 , \8653 , \8658 , \8659 );
and \U$7678 ( \8661 , \8643 , \8660 );
and \U$7679 ( \8662 , \8627 , \8660 );
or \U$7680 ( \8663 , \8644 , \8661 , \8662 );
and \U$7681 ( \8664 , \1377 , \5848 );
and \U$7682 ( \8665 , \1349 , \5846 );
nor \U$7683 ( \8666 , \8664 , \8665 );
xnor \U$7684 ( \8667 , \8666 , \5660 );
and \U$7685 ( \8668 , \1531 , \5474 );
and \U$7686 ( \8669 , \1457 , \5472 );
nor \U$7687 ( \8670 , \8668 , \8669 );
xnor \U$7688 ( \8671 , \8670 , \5242 );
and \U$7689 ( \8672 , \8667 , \8671 );
and \U$7690 ( \8673 , \1656 , \5023 );
and \U$7691 ( \8674 , \1593 , \5021 );
nor \U$7692 ( \8675 , \8673 , \8674 );
xnor \U$7693 ( \8676 , \8675 , \4880 );
and \U$7694 ( \8677 , \8671 , \8676 );
and \U$7695 ( \8678 , \8667 , \8676 );
or \U$7696 ( \8679 , \8672 , \8677 , \8678 );
buf \U$7697 ( \8680 , RIc0d9040_56);
buf \U$7698 ( \8681 , RIc0d90b8_57);
and \U$7699 ( \8682 , \8680 , \8681 );
not \U$7700 ( \8683 , \8682 );
and \U$7701 ( \8684 , \8183 , \8683 );
not \U$7702 ( \8685 , \8684 );
and \U$7703 ( \8686 , \998 , \8435 );
and \U$7704 ( \8687 , \984 , \8433 );
nor \U$7705 ( \8688 , \8686 , \8687 );
xnor \U$7706 ( \8689 , \8688 , \8186 );
and \U$7707 ( \8690 , \8685 , \8689 );
and \U$7708 ( \8691 , \1037 , \7906 );
and \U$7709 ( \8692 , \1016 , \7904 );
nor \U$7710 ( \8693 , \8691 , \8692 );
xnor \U$7711 ( \8694 , \8693 , \7646 );
and \U$7712 ( \8695 , \8689 , \8694 );
and \U$7713 ( \8696 , \8685 , \8694 );
or \U$7714 ( \8697 , \8690 , \8695 , \8696 );
and \U$7715 ( \8698 , \8679 , \8697 );
and \U$7716 ( \8699 , \1093 , \7412 );
and \U$7717 ( \8700 , \1085 , \7410 );
nor \U$7718 ( \8701 , \8699 , \8700 );
xnor \U$7719 ( \8702 , \8701 , \7097 );
and \U$7720 ( \8703 , \1167 , \6903 );
and \U$7721 ( \8704 , \1162 , \6901 );
nor \U$7722 ( \8705 , \8703 , \8704 );
xnor \U$7723 ( \8706 , \8705 , \6563 );
and \U$7724 ( \8707 , \8702 , \8706 );
and \U$7725 ( \8708 , \1272 , \6314 );
and \U$7726 ( \8709 , \1221 , \6312 );
nor \U$7727 ( \8710 , \8708 , \8709 );
xnor \U$7728 ( \8711 , \8710 , \6073 );
and \U$7729 ( \8712 , \8706 , \8711 );
and \U$7730 ( \8713 , \8702 , \8711 );
or \U$7731 ( \8714 , \8707 , \8712 , \8713 );
and \U$7732 ( \8715 , \8697 , \8714 );
and \U$7733 ( \8716 , \8679 , \8714 );
or \U$7734 ( \8717 , \8698 , \8715 , \8716 );
and \U$7735 ( \8718 , \8663 , \8717 );
and \U$7736 ( \8719 , \5447 , \1494 );
and \U$7737 ( \8720 , \5439 , \1492 );
nor \U$7738 ( \8721 , \8719 , \8720 );
xnor \U$7739 ( \8722 , \8721 , \1422 );
and \U$7740 ( \8723 , \5921 , \1360 );
and \U$7741 ( \8724 , \5916 , \1358 );
nor \U$7742 ( \8725 , \8723 , \8724 );
xnor \U$7743 ( \8726 , \8725 , \1317 );
and \U$7744 ( \8727 , \8722 , \8726 );
and \U$7745 ( \8728 , \6444 , \1247 );
and \U$7746 ( \8729 , \6185 , \1245 );
nor \U$7747 ( \8730 , \8728 , \8729 );
xnor \U$7748 ( \8731 , \8730 , \1198 );
and \U$7749 ( \8732 , \8726 , \8731 );
and \U$7750 ( \8733 , \8722 , \8731 );
or \U$7751 ( \8734 , \8727 , \8732 , \8733 );
and \U$7752 ( \8735 , \6825 , \1146 );
and \U$7753 ( \8736 , \6816 , \1144 );
nor \U$7754 ( \8737 , \8735 , \8736 );
xnor \U$7755 ( \8738 , \8737 , \1105 );
and \U$7756 ( \8739 , \7370 , \1076 );
and \U$7757 ( \8740 , \7168 , \1074 );
nor \U$7758 ( \8741 , \8739 , \8740 );
xnor \U$7759 ( \8742 , \8741 , \1046 );
and \U$7760 ( \8743 , \8738 , \8742 );
and \U$7761 ( \8744 , \7845 , \1028 );
and \U$7762 ( \8745 , \7673 , \1026 );
nor \U$7763 ( \8746 , \8744 , \8745 );
xnor \U$7764 ( \8747 , \8746 , \1009 );
and \U$7765 ( \8748 , \8742 , \8747 );
and \U$7766 ( \8749 , \8738 , \8747 );
or \U$7767 ( \8750 , \8743 , \8748 , \8749 );
and \U$7768 ( \8751 , \8734 , \8750 );
and \U$7769 ( \8752 , \4557 , \2028 );
and \U$7770 ( \8753 , \4349 , \2026 );
nor \U$7771 ( \8754 , \8752 , \8753 );
xnor \U$7772 ( \8755 , \8754 , \1892 );
and \U$7773 ( \8756 , \4684 , \1828 );
and \U$7774 ( \8757 , \4679 , \1826 );
nor \U$7775 ( \8758 , \8756 , \8757 );
xnor \U$7776 ( \8759 , \8758 , \1750 );
and \U$7777 ( \8760 , \8755 , \8759 );
and \U$7778 ( \8761 , \5137 , \1664 );
and \U$7779 ( \8762 , \4940 , \1662 );
nor \U$7780 ( \8763 , \8761 , \8762 );
xnor \U$7781 ( \8764 , \8763 , \1570 );
and \U$7782 ( \8765 , \8759 , \8764 );
and \U$7783 ( \8766 , \8755 , \8764 );
or \U$7784 ( \8767 , \8760 , \8765 , \8766 );
and \U$7785 ( \8768 , \8750 , \8767 );
and \U$7786 ( \8769 , \8734 , \8767 );
or \U$7787 ( \8770 , \8751 , \8768 , \8769 );
and \U$7788 ( \8771 , \8717 , \8770 );
and \U$7789 ( \8772 , \8663 , \8770 );
or \U$7790 ( \8773 , \8718 , \8771 , \8772 );
xor \U$7791 ( \8774 , \8349 , \8353 );
xor \U$7792 ( \8775 , \8774 , \8358 );
xor \U$7793 ( \8776 , \8458 , \8462 );
xor \U$7794 ( \8777 , \8776 , \8467 );
and \U$7795 ( \8778 , \8775 , \8777 );
xor \U$7796 ( \8779 , \8383 , \8387 );
xor \U$7797 ( \8780 , \8779 , \8392 );
and \U$7798 ( \8781 , \8777 , \8780 );
and \U$7799 ( \8782 , \8775 , \8780 );
or \U$7800 ( \8783 , \8778 , \8781 , \8782 );
xor \U$7801 ( \8784 , \8418 , \8422 );
xor \U$7802 ( \8785 , \8784 , \8427 );
xor \U$7803 ( \8786 , \8474 , \8478 );
xor \U$7804 ( \8787 , \8786 , \8483 );
and \U$7805 ( \8788 , \8785 , \8787 );
xor \U$7806 ( \8789 , \8491 , \8495 );
xor \U$7807 ( \8790 , \8789 , \8500 );
and \U$7808 ( \8791 , \8787 , \8790 );
and \U$7809 ( \8792 , \8785 , \8790 );
or \U$7810 ( \8793 , \8788 , \8791 , \8792 );
and \U$7811 ( \8794 , \8783 , \8793 );
buf \U$7812 ( \8795 , RIc0dad50_118);
and \U$7813 ( \8796 , \8795 , \985 );
xor \U$7814 ( \8797 , \8365 , \8369 );
xor \U$7815 ( \8798 , \8797 , \8375 );
or \U$7816 ( \8799 , \8796 , \8798 );
and \U$7817 ( \8800 , \8793 , \8799 );
and \U$7818 ( \8801 , \8783 , \8799 );
or \U$7819 ( \8802 , \8794 , \8800 , \8801 );
and \U$7820 ( \8803 , \8773 , \8802 );
xor \U$7821 ( \8804 , \8187 , \8191 );
xor \U$7822 ( \8805 , \8804 , \8196 );
xor \U$7823 ( \8806 , \8511 , \8513 );
xor \U$7824 ( \8807 , \8806 , \8516 );
and \U$7825 ( \8808 , \8805 , \8807 );
xor \U$7826 ( \8809 , \8531 , \8533 );
xor \U$7827 ( \8810 , \8809 , \8536 );
and \U$7828 ( \8811 , \8807 , \8810 );
and \U$7829 ( \8812 , \8805 , \8810 );
or \U$7830 ( \8813 , \8808 , \8811 , \8812 );
and \U$7831 ( \8814 , \8802 , \8813 );
and \U$7832 ( \8815 , \8773 , \8813 );
or \U$7833 ( \8816 , \8803 , \8814 , \8815 );
xor \U$7834 ( \8817 , \8398 , \8453 );
xor \U$7835 ( \8818 , \8817 , \8506 );
xor \U$7836 ( \8819 , \8519 , \8528 );
xor \U$7837 ( \8820 , \8819 , \8539 );
and \U$7838 ( \8821 , \8818 , \8820 );
xor \U$7839 ( \8822 , \8545 , \8547 );
xor \U$7840 ( \8823 , \8822 , \8550 );
and \U$7841 ( \8824 , \8820 , \8823 );
and \U$7842 ( \8825 , \8818 , \8823 );
or \U$7843 ( \8826 , \8821 , \8824 , \8825 );
and \U$7844 ( \8827 , \8816 , \8826 );
xor \U$7845 ( \8828 , \8361 , \8378 );
xor \U$7846 ( \8829 , \8828 , \8395 );
xor \U$7847 ( \8830 , \8470 , \8486 );
xor \U$7848 ( \8831 , \8830 , \8503 );
and \U$7849 ( \8832 , \8829 , \8831 );
xor \U$7850 ( \8833 , \8520 , \8522 );
xor \U$7851 ( \8834 , \8833 , \8525 );
and \U$7852 ( \8835 , \8831 , \8834 );
and \U$7853 ( \8836 , \8829 , \8834 );
or \U$7854 ( \8837 , \8832 , \8835 , \8836 );
xor \U$7855 ( \8838 , \8181 , \8199 );
xor \U$7856 ( \8839 , \8838 , \8216 );
and \U$7857 ( \8840 , \8837 , \8839 );
xor \U$7858 ( \8841 , \8558 , \8560 );
xor \U$7859 ( \8842 , \8841 , \8562 );
and \U$7860 ( \8843 , \8839 , \8842 );
and \U$7861 ( \8844 , \8837 , \8842 );
or \U$7862 ( \8845 , \8840 , \8843 , \8844 );
and \U$7863 ( \8846 , \8826 , \8845 );
and \U$7864 ( \8847 , \8816 , \8845 );
or \U$7865 ( \8848 , \8827 , \8846 , \8847 );
xor \U$7866 ( \8849 , \8509 , \8542 );
xor \U$7867 ( \8850 , \8849 , \8553 );
xor \U$7868 ( \8851 , \8565 , \8567 );
xor \U$7869 ( \8852 , \8851 , \8570 );
and \U$7870 ( \8853 , \8850 , \8852 );
xor \U$7871 ( \8854 , \8576 , \8578 );
and \U$7872 ( \8855 , \8852 , \8854 );
and \U$7873 ( \8856 , \8850 , \8854 );
or \U$7874 ( \8857 , \8853 , \8855 , \8856 );
and \U$7875 ( \8858 , \8848 , \8857 );
xor \U$7876 ( \8859 , \8584 , \8586 );
xor \U$7877 ( \8860 , \8859 , \8588 );
and \U$7878 ( \8861 , \8857 , \8860 );
and \U$7879 ( \8862 , \8848 , \8860 );
or \U$7880 ( \8863 , \8858 , \8861 , \8862 );
xor \U$7881 ( \8864 , \8289 , \8307 );
xor \U$7882 ( \8865 , \8864 , \8313 );
and \U$7883 ( \8866 , \8863 , \8865 );
xor \U$7884 ( \8867 , \8582 , \8591 );
xor \U$7885 ( \8868 , \8867 , \8594 );
and \U$7886 ( \8869 , \8865 , \8868 );
and \U$7887 ( \8870 , \8863 , \8868 );
or \U$7888 ( \8871 , \8866 , \8869 , \8870 );
xor \U$7889 ( \8872 , \8597 , \8599 );
xor \U$7890 ( \8873 , \8872 , \8602 );
and \U$7891 ( \8874 , \8871 , \8873 );
and \U$7892 ( \8875 , \8611 , \8874 );
xor \U$7893 ( \8876 , \8611 , \8874 );
xor \U$7894 ( \8877 , \8871 , \8873 );
and \U$7895 ( \8878 , \2710 , \3586 );
and \U$7896 ( \8879 , \2467 , \3584 );
nor \U$7897 ( \8880 , \8878 , \8879 );
xnor \U$7898 ( \8881 , \8880 , \3437 );
and \U$7899 ( \8882 , \2901 , \3264 );
and \U$7900 ( \8883 , \2715 , \3262 );
nor \U$7901 ( \8884 , \8882 , \8883 );
xnor \U$7902 ( \8885 , \8884 , \3122 );
and \U$7903 ( \8886 , \8881 , \8885 );
and \U$7904 ( \8887 , \3309 , \2968 );
and \U$7905 ( \8888 , \3045 , \2966 );
nor \U$7906 ( \8889 , \8887 , \8888 );
xnor \U$7907 ( \8890 , \8889 , \2831 );
and \U$7908 ( \8891 , \8885 , \8890 );
and \U$7909 ( \8892 , \8881 , \8890 );
or \U$7910 ( \8893 , \8886 , \8891 , \8892 );
and \U$7911 ( \8894 , \3508 , \2762 );
and \U$7912 ( \8895 , \3334 , \2760 );
nor \U$7913 ( \8896 , \8894 , \8895 );
xnor \U$7914 ( \8897 , \8896 , \2610 );
and \U$7915 ( \8898 , \3813 , \2494 );
and \U$7916 ( \8899 , \3675 , \2492 );
nor \U$7917 ( \8900 , \8898 , \8899 );
xnor \U$7918 ( \8901 , \8900 , \2338 );
and \U$7919 ( \8902 , \8897 , \8901 );
and \U$7920 ( \8903 , \4349 , \2222 );
and \U$7921 ( \8904 , \3932 , \2220 );
nor \U$7922 ( \8905 , \8903 , \8904 );
xnor \U$7923 ( \8906 , \8905 , \2109 );
and \U$7924 ( \8907 , \8901 , \8906 );
and \U$7925 ( \8908 , \8897 , \8906 );
or \U$7926 ( \8909 , \8902 , \8907 , \8908 );
and \U$7927 ( \8910 , \8893 , \8909 );
and \U$7928 ( \8911 , \2047 , \4700 );
and \U$7929 ( \8912 , \1942 , \4698 );
nor \U$7930 ( \8913 , \8911 , \8912 );
xnor \U$7931 ( \8914 , \8913 , \4454 );
and \U$7932 ( \8915 , \2168 , \4305 );
and \U$7933 ( \8916 , \2052 , \4303 );
nor \U$7934 ( \8917 , \8915 , \8916 );
xnor \U$7935 ( \8918 , \8917 , \4118 );
and \U$7936 ( \8919 , \8914 , \8918 );
and \U$7937 ( \8920 , \2459 , \3992 );
and \U$7938 ( \8921 , \2283 , \3990 );
nor \U$7939 ( \8922 , \8920 , \8921 );
xnor \U$7940 ( \8923 , \8922 , \3787 );
and \U$7941 ( \8924 , \8918 , \8923 );
and \U$7942 ( \8925 , \8914 , \8923 );
or \U$7943 ( \8926 , \8919 , \8924 , \8925 );
and \U$7944 ( \8927 , \8909 , \8926 );
and \U$7945 ( \8928 , \8893 , \8926 );
or \U$7946 ( \8929 , \8910 , \8927 , \8928 );
and \U$7947 ( \8930 , \5916 , \1494 );
and \U$7948 ( \8931 , \5447 , \1492 );
nor \U$7949 ( \8932 , \8930 , \8931 );
xnor \U$7950 ( \8933 , \8932 , \1422 );
and \U$7951 ( \8934 , \6185 , \1360 );
and \U$7952 ( \8935 , \5921 , \1358 );
nor \U$7953 ( \8936 , \8934 , \8935 );
xnor \U$7954 ( \8937 , \8936 , \1317 );
and \U$7955 ( \8938 , \8933 , \8937 );
and \U$7956 ( \8939 , \6816 , \1247 );
and \U$7957 ( \8940 , \6444 , \1245 );
nor \U$7958 ( \8941 , \8939 , \8940 );
xnor \U$7959 ( \8942 , \8941 , \1198 );
and \U$7960 ( \8943 , \8937 , \8942 );
and \U$7961 ( \8944 , \8933 , \8942 );
or \U$7962 ( \8945 , \8938 , \8943 , \8944 );
and \U$7963 ( \8946 , \4679 , \2028 );
and \U$7964 ( \8947 , \4557 , \2026 );
nor \U$7965 ( \8948 , \8946 , \8947 );
xnor \U$7966 ( \8949 , \8948 , \1892 );
and \U$7967 ( \8950 , \4940 , \1828 );
and \U$7968 ( \8951 , \4684 , \1826 );
nor \U$7969 ( \8952 , \8950 , \8951 );
xnor \U$7970 ( \8953 , \8952 , \1750 );
and \U$7971 ( \8954 , \8949 , \8953 );
and \U$7972 ( \8955 , \5439 , \1664 );
and \U$7973 ( \8956 , \5137 , \1662 );
nor \U$7974 ( \8957 , \8955 , \8956 );
xnor \U$7975 ( \8958 , \8957 , \1570 );
and \U$7976 ( \8959 , \8953 , \8958 );
and \U$7977 ( \8960 , \8949 , \8958 );
or \U$7978 ( \8961 , \8954 , \8959 , \8960 );
and \U$7979 ( \8962 , \8945 , \8961 );
and \U$7980 ( \8963 , \7168 , \1146 );
and \U$7981 ( \8964 , \6825 , \1144 );
nor \U$7982 ( \8965 , \8963 , \8964 );
xnor \U$7983 ( \8966 , \8965 , \1105 );
and \U$7984 ( \8967 , \7673 , \1076 );
and \U$7985 ( \8968 , \7370 , \1074 );
nor \U$7986 ( \8969 , \8967 , \8968 );
xnor \U$7987 ( \8970 , \8969 , \1046 );
and \U$7988 ( \8971 , \8966 , \8970 );
and \U$7989 ( \8972 , \8371 , \1028 );
and \U$7990 ( \8973 , \7845 , \1026 );
nor \U$7991 ( \8974 , \8972 , \8973 );
xnor \U$7992 ( \8975 , \8974 , \1009 );
and \U$7993 ( \8976 , \8970 , \8975 );
and \U$7994 ( \8977 , \8966 , \8975 );
or \U$7995 ( \8978 , \8971 , \8976 , \8977 );
and \U$7996 ( \8979 , \8961 , \8978 );
and \U$7997 ( \8980 , \8945 , \8978 );
or \U$7998 ( \8981 , \8962 , \8979 , \8980 );
and \U$7999 ( \8982 , \8929 , \8981 );
and \U$8000 ( \8983 , \1457 , \5848 );
and \U$8001 ( \8984 , \1377 , \5846 );
nor \U$8002 ( \8985 , \8983 , \8984 );
xnor \U$8003 ( \8986 , \8985 , \5660 );
and \U$8004 ( \8987 , \1593 , \5474 );
and \U$8005 ( \8988 , \1531 , \5472 );
nor \U$8006 ( \8989 , \8987 , \8988 );
xnor \U$8007 ( \8990 , \8989 , \5242 );
and \U$8008 ( \8991 , \8986 , \8990 );
and \U$8009 ( \8992 , \1854 , \5023 );
and \U$8010 ( \8993 , \1656 , \5021 );
nor \U$8011 ( \8994 , \8992 , \8993 );
xnor \U$8012 ( \8995 , \8994 , \4880 );
and \U$8013 ( \8996 , \8990 , \8995 );
and \U$8014 ( \8997 , \8986 , \8995 );
or \U$8015 ( \8998 , \8991 , \8996 , \8997 );
xor \U$8016 ( \8999 , \8183 , \8680 );
xor \U$8017 ( \9000 , \8680 , \8681 );
not \U$8018 ( \9001 , \9000 );
and \U$8019 ( \9002 , \8999 , \9001 );
and \U$8020 ( \9003 , \984 , \9002 );
not \U$8021 ( \9004 , \9003 );
xnor \U$8022 ( \9005 , \9004 , \8684 );
and \U$8023 ( \9006 , \1016 , \8435 );
and \U$8024 ( \9007 , \998 , \8433 );
nor \U$8025 ( \9008 , \9006 , \9007 );
xnor \U$8026 ( \9009 , \9008 , \8186 );
and \U$8027 ( \9010 , \9005 , \9009 );
and \U$8028 ( \9011 , \1085 , \7906 );
and \U$8029 ( \9012 , \1037 , \7904 );
nor \U$8030 ( \9013 , \9011 , \9012 );
xnor \U$8031 ( \9014 , \9013 , \7646 );
and \U$8032 ( \9015 , \9009 , \9014 );
and \U$8033 ( \9016 , \9005 , \9014 );
or \U$8034 ( \9017 , \9010 , \9015 , \9016 );
and \U$8035 ( \9018 , \8998 , \9017 );
and \U$8036 ( \9019 , \1162 , \7412 );
and \U$8037 ( \9020 , \1093 , \7410 );
nor \U$8038 ( \9021 , \9019 , \9020 );
xnor \U$8039 ( \9022 , \9021 , \7097 );
and \U$8040 ( \9023 , \1221 , \6903 );
and \U$8041 ( \9024 , \1167 , \6901 );
nor \U$8042 ( \9025 , \9023 , \9024 );
xnor \U$8043 ( \9026 , \9025 , \6563 );
and \U$8044 ( \9027 , \9022 , \9026 );
and \U$8045 ( \9028 , \1349 , \6314 );
and \U$8046 ( \9029 , \1272 , \6312 );
nor \U$8047 ( \9030 , \9028 , \9029 );
xnor \U$8048 ( \9031 , \9030 , \6073 );
and \U$8049 ( \9032 , \9026 , \9031 );
and \U$8050 ( \9033 , \9022 , \9031 );
or \U$8051 ( \9034 , \9027 , \9032 , \9033 );
and \U$8052 ( \9035 , \9017 , \9034 );
and \U$8053 ( \9036 , \8998 , \9034 );
or \U$8054 ( \9037 , \9018 , \9035 , \9036 );
and \U$8055 ( \9038 , \8981 , \9037 );
and \U$8056 ( \9039 , \8929 , \9037 );
or \U$8057 ( \9040 , \8982 , \9038 , \9039 );
buf \U$8058 ( \9041 , RIc0dadc8_119);
and \U$8059 ( \9042 , \9041 , \991 );
and \U$8060 ( \9043 , \8795 , \989 );
nor \U$8061 ( \9044 , \9042 , \9043 );
xnor \U$8062 ( \9045 , \9044 , \996 );
buf \U$8063 ( \9046 , RIc0dae40_120);
and \U$8064 ( \9047 , \9046 , \985 );
or \U$8065 ( \9048 , \9045 , \9047 );
and \U$8066 ( \9049 , \8795 , \991 );
and \U$8067 ( \9050 , \8371 , \989 );
nor \U$8068 ( \9051 , \9049 , \9050 );
xnor \U$8069 ( \9052 , \9051 , \996 );
and \U$8070 ( \9053 , \9048 , \9052 );
and \U$8071 ( \9054 , \9041 , \985 );
and \U$8072 ( \9055 , \9052 , \9054 );
and \U$8073 ( \9056 , \9048 , \9054 );
or \U$8074 ( \9057 , \9053 , \9055 , \9056 );
xor \U$8075 ( \9058 , \8722 , \8726 );
xor \U$8076 ( \9059 , \9058 , \8731 );
xor \U$8077 ( \9060 , \8738 , \8742 );
xor \U$8078 ( \9061 , \9060 , \8747 );
and \U$8079 ( \9062 , \9059 , \9061 );
xor \U$8080 ( \9063 , \8755 , \8759 );
xor \U$8081 ( \9064 , \9063 , \8764 );
and \U$8082 ( \9065 , \9061 , \9064 );
and \U$8083 ( \9066 , \9059 , \9064 );
or \U$8084 ( \9067 , \9062 , \9065 , \9066 );
and \U$8085 ( \9068 , \9057 , \9067 );
xor \U$8086 ( \9069 , \8615 , \8619 );
xor \U$8087 ( \9070 , \9069 , \8624 );
xor \U$8088 ( \9071 , \8631 , \8635 );
xor \U$8089 ( \9072 , \9071 , \8640 );
and \U$8090 ( \9073 , \9070 , \9072 );
xor \U$8091 ( \9074 , \8648 , \8652 );
xor \U$8092 ( \9075 , \9074 , \8657 );
and \U$8093 ( \9076 , \9072 , \9075 );
and \U$8094 ( \9077 , \9070 , \9075 );
or \U$8095 ( \9078 , \9073 , \9076 , \9077 );
and \U$8096 ( \9079 , \9067 , \9078 );
and \U$8097 ( \9080 , \9057 , \9078 );
or \U$8098 ( \9081 , \9068 , \9079 , \9080 );
and \U$8099 ( \9082 , \9040 , \9081 );
xor \U$8100 ( \9083 , \8667 , \8671 );
xor \U$8101 ( \9084 , \9083 , \8676 );
xor \U$8102 ( \9085 , \8685 , \8689 );
xor \U$8103 ( \9086 , \9085 , \8694 );
and \U$8104 ( \9087 , \9084 , \9086 );
xor \U$8105 ( \9088 , \8702 , \8706 );
xor \U$8106 ( \9089 , \9088 , \8711 );
and \U$8107 ( \9090 , \9086 , \9089 );
and \U$8108 ( \9091 , \9084 , \9089 );
or \U$8109 ( \9092 , \9087 , \9090 , \9091 );
xor \U$8110 ( \9093 , \8402 , \8406 );
xor \U$8111 ( \9094 , \9093 , \8411 );
and \U$8112 ( \9095 , \9092 , \9094 );
xor \U$8113 ( \9096 , \8438 , \8442 );
xor \U$8114 ( \9097 , \9096 , \8447 );
and \U$8115 ( \9098 , \9094 , \9097 );
and \U$8116 ( \9099 , \9092 , \9097 );
or \U$8117 ( \9100 , \9095 , \9098 , \9099 );
and \U$8118 ( \9101 , \9081 , \9100 );
and \U$8119 ( \9102 , \9040 , \9100 );
or \U$8120 ( \9103 , \9082 , \9101 , \9102 );
xor \U$8121 ( \9104 , \8627 , \8643 );
xor \U$8122 ( \9105 , \9104 , \8660 );
xor \U$8123 ( \9106 , \8679 , \8697 );
xor \U$8124 ( \9107 , \9106 , \8714 );
and \U$8125 ( \9108 , \9105 , \9107 );
xor \U$8126 ( \9109 , \8734 , \8750 );
xor \U$8127 ( \9110 , \9109 , \8767 );
and \U$8128 ( \9111 , \9107 , \9110 );
and \U$8129 ( \9112 , \9105 , \9110 );
or \U$8130 ( \9113 , \9108 , \9111 , \9112 );
xor \U$8131 ( \9114 , \8775 , \8777 );
xor \U$8132 ( \9115 , \9114 , \8780 );
xor \U$8133 ( \9116 , \8785 , \8787 );
xor \U$8134 ( \9117 , \9116 , \8790 );
and \U$8135 ( \9118 , \9115 , \9117 );
xnor \U$8136 ( \9119 , \8796 , \8798 );
and \U$8137 ( \9120 , \9117 , \9119 );
and \U$8138 ( \9121 , \9115 , \9119 );
or \U$8139 ( \9122 , \9118 , \9120 , \9121 );
and \U$8140 ( \9123 , \9113 , \9122 );
xor \U$8141 ( \9124 , \8414 , \8430 );
xor \U$8142 ( \9125 , \9124 , \8450 );
and \U$8143 ( \9126 , \9122 , \9125 );
and \U$8144 ( \9127 , \9113 , \9125 );
or \U$8145 ( \9128 , \9123 , \9126 , \9127 );
and \U$8146 ( \9129 , \9103 , \9128 );
xor \U$8147 ( \9130 , \8783 , \8793 );
xor \U$8148 ( \9131 , \9130 , \8799 );
xor \U$8149 ( \9132 , \8829 , \8831 );
xor \U$8150 ( \9133 , \9132 , \8834 );
and \U$8151 ( \9134 , \9131 , \9133 );
xor \U$8152 ( \9135 , \8805 , \8807 );
xor \U$8153 ( \9136 , \9135 , \8810 );
and \U$8154 ( \9137 , \9133 , \9136 );
and \U$8155 ( \9138 , \9131 , \9136 );
or \U$8156 ( \9139 , \9134 , \9137 , \9138 );
and \U$8157 ( \9140 , \9128 , \9139 );
and \U$8158 ( \9141 , \9103 , \9139 );
or \U$8159 ( \9142 , \9129 , \9140 , \9141 );
xor \U$8160 ( \9143 , \8773 , \8802 );
xor \U$8161 ( \9144 , \9143 , \8813 );
xor \U$8162 ( \9145 , \8818 , \8820 );
xor \U$8163 ( \9146 , \9145 , \8823 );
and \U$8164 ( \9147 , \9144 , \9146 );
xor \U$8165 ( \9148 , \8837 , \8839 );
xor \U$8166 ( \9149 , \9148 , \8842 );
and \U$8167 ( \9150 , \9146 , \9149 );
and \U$8168 ( \9151 , \9144 , \9149 );
or \U$8169 ( \9152 , \9147 , \9150 , \9151 );
and \U$8170 ( \9153 , \9142 , \9152 );
xor \U$8171 ( \9154 , \8850 , \8852 );
xor \U$8172 ( \9155 , \9154 , \8854 );
and \U$8173 ( \9156 , \9152 , \9155 );
and \U$8174 ( \9157 , \9142 , \9155 );
or \U$8175 ( \9158 , \9153 , \9156 , \9157 );
xor \U$8176 ( \9159 , \8556 , \8573 );
xor \U$8177 ( \9160 , \9159 , \8579 );
and \U$8178 ( \9161 , \9158 , \9160 );
xor \U$8179 ( \9162 , \8848 , \8857 );
xor \U$8180 ( \9163 , \9162 , \8860 );
and \U$8181 ( \9164 , \9160 , \9163 );
and \U$8182 ( \9165 , \9158 , \9163 );
or \U$8183 ( \9166 , \9161 , \9164 , \9165 );
xor \U$8184 ( \9167 , \8863 , \8865 );
xor \U$8185 ( \9168 , \9167 , \8868 );
and \U$8186 ( \9169 , \9166 , \9168 );
and \U$8187 ( \9170 , \8877 , \9169 );
xor \U$8188 ( \9171 , \8877 , \9169 );
xor \U$8189 ( \9172 , \9166 , \9168 );
and \U$8190 ( \9173 , \1093 , \7906 );
and \U$8191 ( \9174 , \1085 , \7904 );
nor \U$8192 ( \9175 , \9173 , \9174 );
xnor \U$8193 ( \9176 , \9175 , \7646 );
and \U$8194 ( \9177 , \1167 , \7412 );
and \U$8195 ( \9178 , \1162 , \7410 );
nor \U$8196 ( \9179 , \9177 , \9178 );
xnor \U$8197 ( \9180 , \9179 , \7097 );
and \U$8198 ( \9181 , \9176 , \9180 );
and \U$8199 ( \9182 , \1272 , \6903 );
and \U$8200 ( \9183 , \1221 , \6901 );
nor \U$8201 ( \9184 , \9182 , \9183 );
xnor \U$8202 ( \9185 , \9184 , \6563 );
and \U$8203 ( \9186 , \9180 , \9185 );
and \U$8204 ( \9187 , \9176 , \9185 );
or \U$8205 ( \9188 , \9181 , \9186 , \9187 );
buf \U$8206 ( \9189 , RIc0d9130_58);
buf \U$8207 ( \9190 , RIc0d91a8_59);
and \U$8208 ( \9191 , \9189 , \9190 );
not \U$8209 ( \9192 , \9191 );
and \U$8210 ( \9193 , \8681 , \9192 );
not \U$8211 ( \9194 , \9193 );
and \U$8212 ( \9195 , \998 , \9002 );
and \U$8213 ( \9196 , \984 , \9000 );
nor \U$8214 ( \9197 , \9195 , \9196 );
xnor \U$8215 ( \9198 , \9197 , \8684 );
and \U$8216 ( \9199 , \9194 , \9198 );
and \U$8217 ( \9200 , \1037 , \8435 );
and \U$8218 ( \9201 , \1016 , \8433 );
nor \U$8219 ( \9202 , \9200 , \9201 );
xnor \U$8220 ( \9203 , \9202 , \8186 );
and \U$8221 ( \9204 , \9198 , \9203 );
and \U$8222 ( \9205 , \9194 , \9203 );
or \U$8223 ( \9206 , \9199 , \9204 , \9205 );
and \U$8224 ( \9207 , \9188 , \9206 );
and \U$8225 ( \9208 , \1377 , \6314 );
and \U$8226 ( \9209 , \1349 , \6312 );
nor \U$8227 ( \9210 , \9208 , \9209 );
xnor \U$8228 ( \9211 , \9210 , \6073 );
and \U$8229 ( \9212 , \1531 , \5848 );
and \U$8230 ( \9213 , \1457 , \5846 );
nor \U$8231 ( \9214 , \9212 , \9213 );
xnor \U$8232 ( \9215 , \9214 , \5660 );
and \U$8233 ( \9216 , \9211 , \9215 );
and \U$8234 ( \9217 , \1656 , \5474 );
and \U$8235 ( \9218 , \1593 , \5472 );
nor \U$8236 ( \9219 , \9217 , \9218 );
xnor \U$8237 ( \9220 , \9219 , \5242 );
and \U$8238 ( \9221 , \9215 , \9220 );
and \U$8239 ( \9222 , \9211 , \9220 );
or \U$8240 ( \9223 , \9216 , \9221 , \9222 );
and \U$8241 ( \9224 , \9206 , \9223 );
and \U$8242 ( \9225 , \9188 , \9223 );
or \U$8243 ( \9226 , \9207 , \9224 , \9225 );
and \U$8244 ( \9227 , \3334 , \2968 );
and \U$8245 ( \9228 , \3309 , \2966 );
nor \U$8246 ( \9229 , \9227 , \9228 );
xnor \U$8247 ( \9230 , \9229 , \2831 );
and \U$8248 ( \9231 , \3675 , \2762 );
and \U$8249 ( \9232 , \3508 , \2760 );
nor \U$8250 ( \9233 , \9231 , \9232 );
xnor \U$8251 ( \9234 , \9233 , \2610 );
and \U$8252 ( \9235 , \9230 , \9234 );
and \U$8253 ( \9236 , \3932 , \2494 );
and \U$8254 ( \9237 , \3813 , \2492 );
nor \U$8255 ( \9238 , \9236 , \9237 );
xnor \U$8256 ( \9239 , \9238 , \2338 );
and \U$8257 ( \9240 , \9234 , \9239 );
and \U$8258 ( \9241 , \9230 , \9239 );
or \U$8259 ( \9242 , \9235 , \9240 , \9241 );
and \U$8260 ( \9243 , \2467 , \3992 );
and \U$8261 ( \9244 , \2459 , \3990 );
nor \U$8262 ( \9245 , \9243 , \9244 );
xnor \U$8263 ( \9246 , \9245 , \3787 );
and \U$8264 ( \9247 , \2715 , \3586 );
and \U$8265 ( \9248 , \2710 , \3584 );
nor \U$8266 ( \9249 , \9247 , \9248 );
xnor \U$8267 ( \9250 , \9249 , \3437 );
and \U$8268 ( \9251 , \9246 , \9250 );
and \U$8269 ( \9252 , \3045 , \3264 );
and \U$8270 ( \9253 , \2901 , \3262 );
nor \U$8271 ( \9254 , \9252 , \9253 );
xnor \U$8272 ( \9255 , \9254 , \3122 );
and \U$8273 ( \9256 , \9250 , \9255 );
and \U$8274 ( \9257 , \9246 , \9255 );
or \U$8275 ( \9258 , \9251 , \9256 , \9257 );
and \U$8276 ( \9259 , \9242 , \9258 );
and \U$8277 ( \9260 , \1942 , \5023 );
and \U$8278 ( \9261 , \1854 , \5021 );
nor \U$8279 ( \9262 , \9260 , \9261 );
xnor \U$8280 ( \9263 , \9262 , \4880 );
and \U$8281 ( \9264 , \2052 , \4700 );
and \U$8282 ( \9265 , \2047 , \4698 );
nor \U$8283 ( \9266 , \9264 , \9265 );
xnor \U$8284 ( \9267 , \9266 , \4454 );
and \U$8285 ( \9268 , \9263 , \9267 );
and \U$8286 ( \9269 , \2283 , \4305 );
and \U$8287 ( \9270 , \2168 , \4303 );
nor \U$8288 ( \9271 , \9269 , \9270 );
xnor \U$8289 ( \9272 , \9271 , \4118 );
and \U$8290 ( \9273 , \9267 , \9272 );
and \U$8291 ( \9274 , \9263 , \9272 );
or \U$8292 ( \9275 , \9268 , \9273 , \9274 );
and \U$8293 ( \9276 , \9258 , \9275 );
and \U$8294 ( \9277 , \9242 , \9275 );
or \U$8295 ( \9278 , \9259 , \9276 , \9277 );
and \U$8296 ( \9279 , \9226 , \9278 );
and \U$8297 ( \9280 , \5447 , \1664 );
and \U$8298 ( \9281 , \5439 , \1662 );
nor \U$8299 ( \9282 , \9280 , \9281 );
xnor \U$8300 ( \9283 , \9282 , \1570 );
and \U$8301 ( \9284 , \5921 , \1494 );
and \U$8302 ( \9285 , \5916 , \1492 );
nor \U$8303 ( \9286 , \9284 , \9285 );
xnor \U$8304 ( \9287 , \9286 , \1422 );
and \U$8305 ( \9288 , \9283 , \9287 );
and \U$8306 ( \9289 , \6444 , \1360 );
and \U$8307 ( \9290 , \6185 , \1358 );
nor \U$8308 ( \9291 , \9289 , \9290 );
xnor \U$8309 ( \9292 , \9291 , \1317 );
and \U$8310 ( \9293 , \9287 , \9292 );
and \U$8311 ( \9294 , \9283 , \9292 );
or \U$8312 ( \9295 , \9288 , \9293 , \9294 );
and \U$8313 ( \9296 , \4557 , \2222 );
and \U$8314 ( \9297 , \4349 , \2220 );
nor \U$8315 ( \9298 , \9296 , \9297 );
xnor \U$8316 ( \9299 , \9298 , \2109 );
and \U$8317 ( \9300 , \4684 , \2028 );
and \U$8318 ( \9301 , \4679 , \2026 );
nor \U$8319 ( \9302 , \9300 , \9301 );
xnor \U$8320 ( \9303 , \9302 , \1892 );
and \U$8321 ( \9304 , \9299 , \9303 );
and \U$8322 ( \9305 , \5137 , \1828 );
and \U$8323 ( \9306 , \4940 , \1826 );
nor \U$8324 ( \9307 , \9305 , \9306 );
xnor \U$8325 ( \9308 , \9307 , \1750 );
and \U$8326 ( \9309 , \9303 , \9308 );
and \U$8327 ( \9310 , \9299 , \9308 );
or \U$8328 ( \9311 , \9304 , \9309 , \9310 );
and \U$8329 ( \9312 , \9295 , \9311 );
and \U$8330 ( \9313 , \6825 , \1247 );
and \U$8331 ( \9314 , \6816 , \1245 );
nor \U$8332 ( \9315 , \9313 , \9314 );
xnor \U$8333 ( \9316 , \9315 , \1198 );
and \U$8334 ( \9317 , \7370 , \1146 );
and \U$8335 ( \9318 , \7168 , \1144 );
nor \U$8336 ( \9319 , \9317 , \9318 );
xnor \U$8337 ( \9320 , \9319 , \1105 );
and \U$8338 ( \9321 , \9316 , \9320 );
and \U$8339 ( \9322 , \7845 , \1076 );
and \U$8340 ( \9323 , \7673 , \1074 );
nor \U$8341 ( \9324 , \9322 , \9323 );
xnor \U$8342 ( \9325 , \9324 , \1046 );
and \U$8343 ( \9326 , \9320 , \9325 );
and \U$8344 ( \9327 , \9316 , \9325 );
or \U$8345 ( \9328 , \9321 , \9326 , \9327 );
and \U$8346 ( \9329 , \9311 , \9328 );
and \U$8347 ( \9330 , \9295 , \9328 );
or \U$8348 ( \9331 , \9312 , \9329 , \9330 );
and \U$8349 ( \9332 , \9278 , \9331 );
and \U$8350 ( \9333 , \9226 , \9331 );
or \U$8351 ( \9334 , \9279 , \9332 , \9333 );
xor \U$8352 ( \9335 , \8881 , \8885 );
xor \U$8353 ( \9336 , \9335 , \8890 );
xor \U$8354 ( \9337 , \8986 , \8990 );
xor \U$8355 ( \9338 , \9337 , \8995 );
and \U$8356 ( \9339 , \9336 , \9338 );
xor \U$8357 ( \9340 , \8914 , \8918 );
xor \U$8358 ( \9341 , \9340 , \8923 );
and \U$8359 ( \9342 , \9338 , \9341 );
and \U$8360 ( \9343 , \9336 , \9341 );
or \U$8361 ( \9344 , \9339 , \9342 , \9343 );
xor \U$8362 ( \9345 , \8897 , \8901 );
xor \U$8363 ( \9346 , \9345 , \8906 );
xor \U$8364 ( \9347 , \8933 , \8937 );
xor \U$8365 ( \9348 , \9347 , \8942 );
and \U$8366 ( \9349 , \9346 , \9348 );
xor \U$8367 ( \9350 , \8949 , \8953 );
xor \U$8368 ( \9351 , \9350 , \8958 );
and \U$8369 ( \9352 , \9348 , \9351 );
and \U$8370 ( \9353 , \9346 , \9351 );
or \U$8371 ( \9354 , \9349 , \9352 , \9353 );
and \U$8372 ( \9355 , \9344 , \9354 );
and \U$8373 ( \9356 , \8795 , \1028 );
and \U$8374 ( \9357 , \8371 , \1026 );
nor \U$8375 ( \9358 , \9356 , \9357 );
xnor \U$8376 ( \9359 , \9358 , \1009 );
and \U$8377 ( \9360 , \9046 , \991 );
and \U$8378 ( \9361 , \9041 , \989 );
nor \U$8379 ( \9362 , \9360 , \9361 );
xnor \U$8380 ( \9363 , \9362 , \996 );
and \U$8381 ( \9364 , \9359 , \9363 );
buf \U$8382 ( \9365 , RIc0daeb8_121);
and \U$8383 ( \9366 , \9365 , \985 );
and \U$8384 ( \9367 , \9363 , \9366 );
and \U$8385 ( \9368 , \9359 , \9366 );
or \U$8386 ( \9369 , \9364 , \9367 , \9368 );
xor \U$8387 ( \9370 , \8966 , \8970 );
xor \U$8388 ( \9371 , \9370 , \8975 );
and \U$8389 ( \9372 , \9369 , \9371 );
xnor \U$8390 ( \9373 , \9045 , \9047 );
and \U$8391 ( \9374 , \9371 , \9373 );
and \U$8392 ( \9375 , \9369 , \9373 );
or \U$8393 ( \9376 , \9372 , \9374 , \9375 );
and \U$8394 ( \9377 , \9354 , \9376 );
and \U$8395 ( \9378 , \9344 , \9376 );
or \U$8396 ( \9379 , \9355 , \9377 , \9378 );
and \U$8397 ( \9380 , \9334 , \9379 );
xor \U$8398 ( \9381 , \9059 , \9061 );
xor \U$8399 ( \9382 , \9381 , \9064 );
xor \U$8400 ( \9383 , \9070 , \9072 );
xor \U$8401 ( \9384 , \9383 , \9075 );
and \U$8402 ( \9385 , \9382 , \9384 );
xor \U$8403 ( \9386 , \9084 , \9086 );
xor \U$8404 ( \9387 , \9386 , \9089 );
and \U$8405 ( \9388 , \9384 , \9387 );
and \U$8406 ( \9389 , \9382 , \9387 );
or \U$8407 ( \9390 , \9385 , \9388 , \9389 );
and \U$8408 ( \9391 , \9379 , \9390 );
and \U$8409 ( \9392 , \9334 , \9390 );
or \U$8410 ( \9393 , \9380 , \9391 , \9392 );
xor \U$8411 ( \9394 , \8929 , \8981 );
xor \U$8412 ( \9395 , \9394 , \9037 );
xor \U$8413 ( \9396 , \9057 , \9067 );
xor \U$8414 ( \9397 , \9396 , \9078 );
and \U$8415 ( \9398 , \9395 , \9397 );
xor \U$8416 ( \9399 , \9092 , \9094 );
xor \U$8417 ( \9400 , \9399 , \9097 );
and \U$8418 ( \9401 , \9397 , \9400 );
and \U$8419 ( \9402 , \9395 , \9400 );
or \U$8420 ( \9403 , \9398 , \9401 , \9402 );
and \U$8421 ( \9404 , \9393 , \9403 );
xor \U$8422 ( \9405 , \8893 , \8909 );
xor \U$8423 ( \9406 , \9405 , \8926 );
xor \U$8424 ( \9407 , \8945 , \8961 );
xor \U$8425 ( \9408 , \9407 , \8978 );
and \U$8426 ( \9409 , \9406 , \9408 );
xor \U$8427 ( \9410 , \9048 , \9052 );
xor \U$8428 ( \9411 , \9410 , \9054 );
and \U$8429 ( \9412 , \9408 , \9411 );
and \U$8430 ( \9413 , \9406 , \9411 );
or \U$8431 ( \9414 , \9409 , \9412 , \9413 );
xor \U$8432 ( \9415 , \9105 , \9107 );
xor \U$8433 ( \9416 , \9415 , \9110 );
and \U$8434 ( \9417 , \9414 , \9416 );
xor \U$8435 ( \9418 , \9115 , \9117 );
xor \U$8436 ( \9419 , \9418 , \9119 );
and \U$8437 ( \9420 , \9416 , \9419 );
and \U$8438 ( \9421 , \9414 , \9419 );
or \U$8439 ( \9422 , \9417 , \9420 , \9421 );
and \U$8440 ( \9423 , \9403 , \9422 );
and \U$8441 ( \9424 , \9393 , \9422 );
or \U$8442 ( \9425 , \9404 , \9423 , \9424 );
xor \U$8443 ( \9426 , \8663 , \8717 );
xor \U$8444 ( \9427 , \9426 , \8770 );
xor \U$8445 ( \9428 , \9113 , \9122 );
xor \U$8446 ( \9429 , \9428 , \9125 );
and \U$8447 ( \9430 , \9427 , \9429 );
xor \U$8448 ( \9431 , \9131 , \9133 );
xor \U$8449 ( \9432 , \9431 , \9136 );
and \U$8450 ( \9433 , \9429 , \9432 );
and \U$8451 ( \9434 , \9427 , \9432 );
or \U$8452 ( \9435 , \9430 , \9433 , \9434 );
and \U$8453 ( \9436 , \9425 , \9435 );
xor \U$8454 ( \9437 , \9144 , \9146 );
xor \U$8455 ( \9438 , \9437 , \9149 );
and \U$8456 ( \9439 , \9435 , \9438 );
and \U$8457 ( \9440 , \9425 , \9438 );
or \U$8458 ( \9441 , \9436 , \9439 , \9440 );
xor \U$8459 ( \9442 , \8816 , \8826 );
xor \U$8460 ( \9443 , \9442 , \8845 );
and \U$8461 ( \9444 , \9441 , \9443 );
xor \U$8462 ( \9445 , \9142 , \9152 );
xor \U$8463 ( \9446 , \9445 , \9155 );
and \U$8464 ( \9447 , \9443 , \9446 );
and \U$8465 ( \9448 , \9441 , \9446 );
or \U$8466 ( \9449 , \9444 , \9447 , \9448 );
xor \U$8467 ( \9450 , \9158 , \9160 );
xor \U$8468 ( \9451 , \9450 , \9163 );
and \U$8469 ( \9452 , \9449 , \9451 );
and \U$8470 ( \9453 , \9172 , \9452 );
xor \U$8471 ( \9454 , \9172 , \9452 );
xor \U$8472 ( \9455 , \9449 , \9451 );
and \U$8473 ( \9456 , \3508 , \2968 );
and \U$8474 ( \9457 , \3334 , \2966 );
nor \U$8475 ( \9458 , \9456 , \9457 );
xnor \U$8476 ( \9459 , \9458 , \2831 );
and \U$8477 ( \9460 , \3813 , \2762 );
and \U$8478 ( \9461 , \3675 , \2760 );
nor \U$8479 ( \9462 , \9460 , \9461 );
xnor \U$8480 ( \9463 , \9462 , \2610 );
and \U$8481 ( \9464 , \9459 , \9463 );
and \U$8482 ( \9465 , \4349 , \2494 );
and \U$8483 ( \9466 , \3932 , \2492 );
nor \U$8484 ( \9467 , \9465 , \9466 );
xnor \U$8485 ( \9468 , \9467 , \2338 );
and \U$8486 ( \9469 , \9463 , \9468 );
and \U$8487 ( \9470 , \9459 , \9468 );
or \U$8488 ( \9471 , \9464 , \9469 , \9470 );
and \U$8489 ( \9472 , \2047 , \5023 );
and \U$8490 ( \9473 , \1942 , \5021 );
nor \U$8491 ( \9474 , \9472 , \9473 );
xnor \U$8492 ( \9475 , \9474 , \4880 );
and \U$8493 ( \9476 , \2168 , \4700 );
and \U$8494 ( \9477 , \2052 , \4698 );
nor \U$8495 ( \9478 , \9476 , \9477 );
xnor \U$8496 ( \9479 , \9478 , \4454 );
and \U$8497 ( \9480 , \9475 , \9479 );
and \U$8498 ( \9481 , \2459 , \4305 );
and \U$8499 ( \9482 , \2283 , \4303 );
nor \U$8500 ( \9483 , \9481 , \9482 );
xnor \U$8501 ( \9484 , \9483 , \4118 );
and \U$8502 ( \9485 , \9479 , \9484 );
and \U$8503 ( \9486 , \9475 , \9484 );
or \U$8504 ( \9487 , \9480 , \9485 , \9486 );
and \U$8505 ( \9488 , \9471 , \9487 );
and \U$8506 ( \9489 , \2710 , \3992 );
and \U$8507 ( \9490 , \2467 , \3990 );
nor \U$8508 ( \9491 , \9489 , \9490 );
xnor \U$8509 ( \9492 , \9491 , \3787 );
and \U$8510 ( \9493 , \2901 , \3586 );
and \U$8511 ( \9494 , \2715 , \3584 );
nor \U$8512 ( \9495 , \9493 , \9494 );
xnor \U$8513 ( \9496 , \9495 , \3437 );
and \U$8514 ( \9497 , \9492 , \9496 );
and \U$8515 ( \9498 , \3309 , \3264 );
and \U$8516 ( \9499 , \3045 , \3262 );
nor \U$8517 ( \9500 , \9498 , \9499 );
xnor \U$8518 ( \9501 , \9500 , \3122 );
and \U$8519 ( \9502 , \9496 , \9501 );
and \U$8520 ( \9503 , \9492 , \9501 );
or \U$8521 ( \9504 , \9497 , \9502 , \9503 );
and \U$8522 ( \9505 , \9487 , \9504 );
and \U$8523 ( \9506 , \9471 , \9504 );
or \U$8524 ( \9507 , \9488 , \9505 , \9506 );
and \U$8525 ( \9508 , \7168 , \1247 );
and \U$8526 ( \9509 , \6825 , \1245 );
nor \U$8527 ( \9510 , \9508 , \9509 );
xnor \U$8528 ( \9511 , \9510 , \1198 );
and \U$8529 ( \9512 , \7673 , \1146 );
and \U$8530 ( \9513 , \7370 , \1144 );
nor \U$8531 ( \9514 , \9512 , \9513 );
xnor \U$8532 ( \9515 , \9514 , \1105 );
and \U$8533 ( \9516 , \9511 , \9515 );
and \U$8534 ( \9517 , \8371 , \1076 );
and \U$8535 ( \9518 , \7845 , \1074 );
nor \U$8536 ( \9519 , \9517 , \9518 );
xnor \U$8537 ( \9520 , \9519 , \1046 );
and \U$8538 ( \9521 , \9515 , \9520 );
and \U$8539 ( \9522 , \9511 , \9520 );
or \U$8540 ( \9523 , \9516 , \9521 , \9522 );
and \U$8541 ( \9524 , \5916 , \1664 );
and \U$8542 ( \9525 , \5447 , \1662 );
nor \U$8543 ( \9526 , \9524 , \9525 );
xnor \U$8544 ( \9527 , \9526 , \1570 );
and \U$8545 ( \9528 , \6185 , \1494 );
and \U$8546 ( \9529 , \5921 , \1492 );
nor \U$8547 ( \9530 , \9528 , \9529 );
xnor \U$8548 ( \9531 , \9530 , \1422 );
and \U$8549 ( \9532 , \9527 , \9531 );
and \U$8550 ( \9533 , \6816 , \1360 );
and \U$8551 ( \9534 , \6444 , \1358 );
nor \U$8552 ( \9535 , \9533 , \9534 );
xnor \U$8553 ( \9536 , \9535 , \1317 );
and \U$8554 ( \9537 , \9531 , \9536 );
and \U$8555 ( \9538 , \9527 , \9536 );
or \U$8556 ( \9539 , \9532 , \9537 , \9538 );
and \U$8557 ( \9540 , \9523 , \9539 );
and \U$8558 ( \9541 , \4679 , \2222 );
and \U$8559 ( \9542 , \4557 , \2220 );
nor \U$8560 ( \9543 , \9541 , \9542 );
xnor \U$8561 ( \9544 , \9543 , \2109 );
and \U$8562 ( \9545 , \4940 , \2028 );
and \U$8563 ( \9546 , \4684 , \2026 );
nor \U$8564 ( \9547 , \9545 , \9546 );
xnor \U$8565 ( \9548 , \9547 , \1892 );
and \U$8566 ( \9549 , \9544 , \9548 );
and \U$8567 ( \9550 , \5439 , \1828 );
and \U$8568 ( \9551 , \5137 , \1826 );
nor \U$8569 ( \9552 , \9550 , \9551 );
xnor \U$8570 ( \9553 , \9552 , \1750 );
and \U$8571 ( \9554 , \9548 , \9553 );
and \U$8572 ( \9555 , \9544 , \9553 );
or \U$8573 ( \9556 , \9549 , \9554 , \9555 );
and \U$8574 ( \9557 , \9539 , \9556 );
and \U$8575 ( \9558 , \9523 , \9556 );
or \U$8576 ( \9559 , \9540 , \9557 , \9558 );
and \U$8577 ( \9560 , \9507 , \9559 );
xor \U$8578 ( \9561 , \8681 , \9189 );
xor \U$8579 ( \9562 , \9189 , \9190 );
not \U$8580 ( \9563 , \9562 );
and \U$8581 ( \9564 , \9561 , \9563 );
and \U$8582 ( \9565 , \984 , \9564 );
not \U$8583 ( \9566 , \9565 );
xnor \U$8584 ( \9567 , \9566 , \9193 );
and \U$8585 ( \9568 , \1016 , \9002 );
and \U$8586 ( \9569 , \998 , \9000 );
nor \U$8587 ( \9570 , \9568 , \9569 );
xnor \U$8588 ( \9571 , \9570 , \8684 );
and \U$8589 ( \9572 , \9567 , \9571 );
and \U$8590 ( \9573 , \1085 , \8435 );
and \U$8591 ( \9574 , \1037 , \8433 );
nor \U$8592 ( \9575 , \9573 , \9574 );
xnor \U$8593 ( \9576 , \9575 , \8186 );
and \U$8594 ( \9577 , \9571 , \9576 );
and \U$8595 ( \9578 , \9567 , \9576 );
or \U$8596 ( \9579 , \9572 , \9577 , \9578 );
and \U$8597 ( \9580 , \1457 , \6314 );
and \U$8598 ( \9581 , \1377 , \6312 );
nor \U$8599 ( \9582 , \9580 , \9581 );
xnor \U$8600 ( \9583 , \9582 , \6073 );
and \U$8601 ( \9584 , \1593 , \5848 );
and \U$8602 ( \9585 , \1531 , \5846 );
nor \U$8603 ( \9586 , \9584 , \9585 );
xnor \U$8604 ( \9587 , \9586 , \5660 );
and \U$8605 ( \9588 , \9583 , \9587 );
and \U$8606 ( \9589 , \1854 , \5474 );
and \U$8607 ( \9590 , \1656 , \5472 );
nor \U$8608 ( \9591 , \9589 , \9590 );
xnor \U$8609 ( \9592 , \9591 , \5242 );
and \U$8610 ( \9593 , \9587 , \9592 );
and \U$8611 ( \9594 , \9583 , \9592 );
or \U$8612 ( \9595 , \9588 , \9593 , \9594 );
and \U$8613 ( \9596 , \9579 , \9595 );
and \U$8614 ( \9597 , \1162 , \7906 );
and \U$8615 ( \9598 , \1093 , \7904 );
nor \U$8616 ( \9599 , \9597 , \9598 );
xnor \U$8617 ( \9600 , \9599 , \7646 );
and \U$8618 ( \9601 , \1221 , \7412 );
and \U$8619 ( \9602 , \1167 , \7410 );
nor \U$8620 ( \9603 , \9601 , \9602 );
xnor \U$8621 ( \9604 , \9603 , \7097 );
and \U$8622 ( \9605 , \9600 , \9604 );
and \U$8623 ( \9606 , \1349 , \6903 );
and \U$8624 ( \9607 , \1272 , \6901 );
nor \U$8625 ( \9608 , \9606 , \9607 );
xnor \U$8626 ( \9609 , \9608 , \6563 );
and \U$8627 ( \9610 , \9604 , \9609 );
and \U$8628 ( \9611 , \9600 , \9609 );
or \U$8629 ( \9612 , \9605 , \9610 , \9611 );
and \U$8630 ( \9613 , \9595 , \9612 );
and \U$8631 ( \9614 , \9579 , \9612 );
or \U$8632 ( \9615 , \9596 , \9613 , \9614 );
and \U$8633 ( \9616 , \9559 , \9615 );
and \U$8634 ( \9617 , \9507 , \9615 );
or \U$8635 ( \9618 , \9560 , \9616 , \9617 );
xor \U$8636 ( \9619 , \9211 , \9215 );
xor \U$8637 ( \9620 , \9619 , \9220 );
xor \U$8638 ( \9621 , \9246 , \9250 );
xor \U$8639 ( \9622 , \9621 , \9255 );
and \U$8640 ( \9623 , \9620 , \9622 );
xor \U$8641 ( \9624 , \9263 , \9267 );
xor \U$8642 ( \9625 , \9624 , \9272 );
and \U$8643 ( \9626 , \9622 , \9625 );
and \U$8644 ( \9627 , \9620 , \9625 );
or \U$8645 ( \9628 , \9623 , \9626 , \9627 );
xor \U$8646 ( \9629 , \9230 , \9234 );
xor \U$8647 ( \9630 , \9629 , \9239 );
xor \U$8648 ( \9631 , \9283 , \9287 );
xor \U$8649 ( \9632 , \9631 , \9292 );
and \U$8650 ( \9633 , \9630 , \9632 );
xor \U$8651 ( \9634 , \9299 , \9303 );
xor \U$8652 ( \9635 , \9634 , \9308 );
and \U$8653 ( \9636 , \9632 , \9635 );
and \U$8654 ( \9637 , \9630 , \9635 );
or \U$8655 ( \9638 , \9633 , \9636 , \9637 );
and \U$8656 ( \9639 , \9628 , \9638 );
and \U$8657 ( \9640 , \9041 , \1028 );
and \U$8658 ( \9641 , \8795 , \1026 );
nor \U$8659 ( \9642 , \9640 , \9641 );
xnor \U$8660 ( \9643 , \9642 , \1009 );
and \U$8661 ( \9644 , \9365 , \991 );
and \U$8662 ( \9645 , \9046 , \989 );
nor \U$8663 ( \9646 , \9644 , \9645 );
xnor \U$8664 ( \9647 , \9646 , \996 );
and \U$8665 ( \9648 , \9643 , \9647 );
buf \U$8666 ( \9649 , RIc0daf30_122);
and \U$8667 ( \9650 , \9649 , \985 );
and \U$8668 ( \9651 , \9647 , \9650 );
and \U$8669 ( \9652 , \9643 , \9650 );
or \U$8670 ( \9653 , \9648 , \9651 , \9652 );
xor \U$8671 ( \9654 , \9359 , \9363 );
xor \U$8672 ( \9655 , \9654 , \9366 );
and \U$8673 ( \9656 , \9653 , \9655 );
xor \U$8674 ( \9657 , \9316 , \9320 );
xor \U$8675 ( \9658 , \9657 , \9325 );
and \U$8676 ( \9659 , \9655 , \9658 );
and \U$8677 ( \9660 , \9653 , \9658 );
or \U$8678 ( \9661 , \9656 , \9659 , \9660 );
and \U$8679 ( \9662 , \9638 , \9661 );
and \U$8680 ( \9663 , \9628 , \9661 );
or \U$8681 ( \9664 , \9639 , \9662 , \9663 );
and \U$8682 ( \9665 , \9618 , \9664 );
xor \U$8683 ( \9666 , \9005 , \9009 );
xor \U$8684 ( \9667 , \9666 , \9014 );
xor \U$8685 ( \9668 , \9022 , \9026 );
xor \U$8686 ( \9669 , \9668 , \9031 );
and \U$8687 ( \9670 , \9667 , \9669 );
xor \U$8688 ( \9671 , \9336 , \9338 );
xor \U$8689 ( \9672 , \9671 , \9341 );
and \U$8690 ( \9673 , \9669 , \9672 );
and \U$8691 ( \9674 , \9667 , \9672 );
or \U$8692 ( \9675 , \9670 , \9673 , \9674 );
and \U$8693 ( \9676 , \9664 , \9675 );
and \U$8694 ( \9677 , \9618 , \9675 );
or \U$8695 ( \9678 , \9665 , \9676 , \9677 );
xor \U$8696 ( \9679 , \9295 , \9311 );
xor \U$8697 ( \9680 , \9679 , \9328 );
xor \U$8698 ( \9681 , \9346 , \9348 );
xor \U$8699 ( \9682 , \9681 , \9351 );
and \U$8700 ( \9683 , \9680 , \9682 );
xor \U$8701 ( \9684 , \9369 , \9371 );
xor \U$8702 ( \9685 , \9684 , \9373 );
and \U$8703 ( \9686 , \9682 , \9685 );
and \U$8704 ( \9687 , \9680 , \9685 );
or \U$8705 ( \9688 , \9683 , \9686 , \9687 );
xor \U$8706 ( \9689 , \8998 , \9017 );
xor \U$8707 ( \9690 , \9689 , \9034 );
and \U$8708 ( \9691 , \9688 , \9690 );
xor \U$8709 ( \9692 , \9406 , \9408 );
xor \U$8710 ( \9693 , \9692 , \9411 );
and \U$8711 ( \9694 , \9690 , \9693 );
and \U$8712 ( \9695 , \9688 , \9693 );
or \U$8713 ( \9696 , \9691 , \9694 , \9695 );
and \U$8714 ( \9697 , \9678 , \9696 );
xor \U$8715 ( \9698 , \9226 , \9278 );
xor \U$8716 ( \9699 , \9698 , \9331 );
xor \U$8717 ( \9700 , \9344 , \9354 );
xor \U$8718 ( \9701 , \9700 , \9376 );
and \U$8719 ( \9702 , \9699 , \9701 );
xor \U$8720 ( \9703 , \9382 , \9384 );
xor \U$8721 ( \9704 , \9703 , \9387 );
and \U$8722 ( \9705 , \9701 , \9704 );
and \U$8723 ( \9706 , \9699 , \9704 );
or \U$8724 ( \9707 , \9702 , \9705 , \9706 );
and \U$8725 ( \9708 , \9696 , \9707 );
and \U$8726 ( \9709 , \9678 , \9707 );
or \U$8727 ( \9710 , \9697 , \9708 , \9709 );
xor \U$8728 ( \9711 , \9334 , \9379 );
xor \U$8729 ( \9712 , \9711 , \9390 );
xor \U$8730 ( \9713 , \9395 , \9397 );
xor \U$8731 ( \9714 , \9713 , \9400 );
and \U$8732 ( \9715 , \9712 , \9714 );
xor \U$8733 ( \9716 , \9414 , \9416 );
xor \U$8734 ( \9717 , \9716 , \9419 );
and \U$8735 ( \9718 , \9714 , \9717 );
and \U$8736 ( \9719 , \9712 , \9717 );
or \U$8737 ( \9720 , \9715 , \9718 , \9719 );
and \U$8738 ( \9721 , \9710 , \9720 );
xor \U$8739 ( \9722 , \9040 , \9081 );
xor \U$8740 ( \9723 , \9722 , \9100 );
and \U$8741 ( \9724 , \9720 , \9723 );
and \U$8742 ( \9725 , \9710 , \9723 );
or \U$8743 ( \9726 , \9721 , \9724 , \9725 );
xor \U$8744 ( \9727 , \9393 , \9403 );
xor \U$8745 ( \9728 , \9727 , \9422 );
xor \U$8746 ( \9729 , \9427 , \9429 );
xor \U$8747 ( \9730 , \9729 , \9432 );
and \U$8748 ( \9731 , \9728 , \9730 );
and \U$8749 ( \9732 , \9726 , \9731 );
xor \U$8750 ( \9733 , \9103 , \9128 );
xor \U$8751 ( \9734 , \9733 , \9139 );
and \U$8752 ( \9735 , \9731 , \9734 );
and \U$8753 ( \9736 , \9726 , \9734 );
or \U$8754 ( \9737 , \9732 , \9735 , \9736 );
xor \U$8755 ( \9738 , \9441 , \9443 );
xor \U$8756 ( \9739 , \9738 , \9446 );
and \U$8757 ( \9740 , \9737 , \9739 );
and \U$8758 ( \9741 , \9455 , \9740 );
xor \U$8759 ( \9742 , \9455 , \9740 );
xor \U$8760 ( \9743 , \9737 , \9739 );
xor \U$8761 ( \9744 , \9511 , \9515 );
xor \U$8762 ( \9745 , \9744 , \9520 );
xor \U$8763 ( \9746 , \9527 , \9531 );
xor \U$8764 ( \9747 , \9746 , \9536 );
and \U$8765 ( \9748 , \9745 , \9747 );
xor \U$8766 ( \9749 , \9544 , \9548 );
xor \U$8767 ( \9750 , \9749 , \9553 );
and \U$8768 ( \9751 , \9747 , \9750 );
and \U$8769 ( \9752 , \9745 , \9750 );
or \U$8770 ( \9753 , \9748 , \9751 , \9752 );
xor \U$8771 ( \9754 , \9459 , \9463 );
xor \U$8772 ( \9755 , \9754 , \9468 );
xor \U$8773 ( \9756 , \9475 , \9479 );
xor \U$8774 ( \9757 , \9756 , \9484 );
and \U$8775 ( \9758 , \9755 , \9757 );
xor \U$8776 ( \9759 , \9492 , \9496 );
xor \U$8777 ( \9760 , \9759 , \9501 );
and \U$8778 ( \9761 , \9757 , \9760 );
and \U$8779 ( \9762 , \9755 , \9760 );
or \U$8780 ( \9763 , \9758 , \9761 , \9762 );
and \U$8781 ( \9764 , \9753 , \9763 );
and \U$8782 ( \9765 , \8795 , \1076 );
and \U$8783 ( \9766 , \8371 , \1074 );
nor \U$8784 ( \9767 , \9765 , \9766 );
xnor \U$8785 ( \9768 , \9767 , \1046 );
and \U$8786 ( \9769 , \9046 , \1028 );
and \U$8787 ( \9770 , \9041 , \1026 );
nor \U$8788 ( \9771 , \9769 , \9770 );
xnor \U$8789 ( \9772 , \9771 , \1009 );
and \U$8790 ( \9773 , \9768 , \9772 );
and \U$8791 ( \9774 , \9649 , \991 );
and \U$8792 ( \9775 , \9365 , \989 );
nor \U$8793 ( \9776 , \9774 , \9775 );
xnor \U$8794 ( \9777 , \9776 , \996 );
and \U$8795 ( \9778 , \9772 , \9777 );
and \U$8796 ( \9779 , \9768 , \9777 );
or \U$8797 ( \9780 , \9773 , \9778 , \9779 );
xor \U$8798 ( \9781 , \9643 , \9647 );
xor \U$8799 ( \9782 , \9781 , \9650 );
or \U$8800 ( \9783 , \9780 , \9782 );
and \U$8801 ( \9784 , \9763 , \9783 );
and \U$8802 ( \9785 , \9753 , \9783 );
or \U$8803 ( \9786 , \9764 , \9784 , \9785 );
buf \U$8804 ( \9787 , RIc0d9220_60);
buf \U$8805 ( \9788 , RIc0d9298_61);
and \U$8806 ( \9789 , \9787 , \9788 );
not \U$8807 ( \9790 , \9789 );
and \U$8808 ( \9791 , \9190 , \9790 );
not \U$8809 ( \9792 , \9791 );
and \U$8810 ( \9793 , \998 , \9564 );
and \U$8811 ( \9794 , \984 , \9562 );
nor \U$8812 ( \9795 , \9793 , \9794 );
xnor \U$8813 ( \9796 , \9795 , \9193 );
and \U$8814 ( \9797 , \9792 , \9796 );
and \U$8815 ( \9798 , \1037 , \9002 );
and \U$8816 ( \9799 , \1016 , \9000 );
nor \U$8817 ( \9800 , \9798 , \9799 );
xnor \U$8818 ( \9801 , \9800 , \8684 );
and \U$8819 ( \9802 , \9796 , \9801 );
and \U$8820 ( \9803 , \9792 , \9801 );
or \U$8821 ( \9804 , \9797 , \9802 , \9803 );
and \U$8822 ( \9805 , \1377 , \6903 );
and \U$8823 ( \9806 , \1349 , \6901 );
nor \U$8824 ( \9807 , \9805 , \9806 );
xnor \U$8825 ( \9808 , \9807 , \6563 );
and \U$8826 ( \9809 , \1531 , \6314 );
and \U$8827 ( \9810 , \1457 , \6312 );
nor \U$8828 ( \9811 , \9809 , \9810 );
xnor \U$8829 ( \9812 , \9811 , \6073 );
and \U$8830 ( \9813 , \9808 , \9812 );
and \U$8831 ( \9814 , \1656 , \5848 );
and \U$8832 ( \9815 , \1593 , \5846 );
nor \U$8833 ( \9816 , \9814 , \9815 );
xnor \U$8834 ( \9817 , \9816 , \5660 );
and \U$8835 ( \9818 , \9812 , \9817 );
and \U$8836 ( \9819 , \9808 , \9817 );
or \U$8837 ( \9820 , \9813 , \9818 , \9819 );
and \U$8838 ( \9821 , \9804 , \9820 );
and \U$8839 ( \9822 , \1093 , \8435 );
and \U$8840 ( \9823 , \1085 , \8433 );
nor \U$8841 ( \9824 , \9822 , \9823 );
xnor \U$8842 ( \9825 , \9824 , \8186 );
and \U$8843 ( \9826 , \1167 , \7906 );
and \U$8844 ( \9827 , \1162 , \7904 );
nor \U$8845 ( \9828 , \9826 , \9827 );
xnor \U$8846 ( \9829 , \9828 , \7646 );
and \U$8847 ( \9830 , \9825 , \9829 );
and \U$8848 ( \9831 , \1272 , \7412 );
and \U$8849 ( \9832 , \1221 , \7410 );
nor \U$8850 ( \9833 , \9831 , \9832 );
xnor \U$8851 ( \9834 , \9833 , \7097 );
and \U$8852 ( \9835 , \9829 , \9834 );
and \U$8853 ( \9836 , \9825 , \9834 );
or \U$8854 ( \9837 , \9830 , \9835 , \9836 );
and \U$8855 ( \9838 , \9820 , \9837 );
and \U$8856 ( \9839 , \9804 , \9837 );
or \U$8857 ( \9840 , \9821 , \9838 , \9839 );
and \U$8858 ( \9841 , \2467 , \4305 );
and \U$8859 ( \9842 , \2459 , \4303 );
nor \U$8860 ( \9843 , \9841 , \9842 );
xnor \U$8861 ( \9844 , \9843 , \4118 );
and \U$8862 ( \9845 , \2715 , \3992 );
and \U$8863 ( \9846 , \2710 , \3990 );
nor \U$8864 ( \9847 , \9845 , \9846 );
xnor \U$8865 ( \9848 , \9847 , \3787 );
and \U$8866 ( \9849 , \9844 , \9848 );
and \U$8867 ( \9850 , \3045 , \3586 );
and \U$8868 ( \9851 , \2901 , \3584 );
nor \U$8869 ( \9852 , \9850 , \9851 );
xnor \U$8870 ( \9853 , \9852 , \3437 );
and \U$8871 ( \9854 , \9848 , \9853 );
and \U$8872 ( \9855 , \9844 , \9853 );
or \U$8873 ( \9856 , \9849 , \9854 , \9855 );
and \U$8874 ( \9857 , \3334 , \3264 );
and \U$8875 ( \9858 , \3309 , \3262 );
nor \U$8876 ( \9859 , \9857 , \9858 );
xnor \U$8877 ( \9860 , \9859 , \3122 );
and \U$8878 ( \9861 , \3675 , \2968 );
and \U$8879 ( \9862 , \3508 , \2966 );
nor \U$8880 ( \9863 , \9861 , \9862 );
xnor \U$8881 ( \9864 , \9863 , \2831 );
and \U$8882 ( \9865 , \9860 , \9864 );
and \U$8883 ( \9866 , \3932 , \2762 );
and \U$8884 ( \9867 , \3813 , \2760 );
nor \U$8885 ( \9868 , \9866 , \9867 );
xnor \U$8886 ( \9869 , \9868 , \2610 );
and \U$8887 ( \9870 , \9864 , \9869 );
and \U$8888 ( \9871 , \9860 , \9869 );
or \U$8889 ( \9872 , \9865 , \9870 , \9871 );
and \U$8890 ( \9873 , \9856 , \9872 );
and \U$8891 ( \9874 , \1942 , \5474 );
and \U$8892 ( \9875 , \1854 , \5472 );
nor \U$8893 ( \9876 , \9874 , \9875 );
xnor \U$8894 ( \9877 , \9876 , \5242 );
and \U$8895 ( \9878 , \2052 , \5023 );
and \U$8896 ( \9879 , \2047 , \5021 );
nor \U$8897 ( \9880 , \9878 , \9879 );
xnor \U$8898 ( \9881 , \9880 , \4880 );
and \U$8899 ( \9882 , \9877 , \9881 );
and \U$8900 ( \9883 , \2283 , \4700 );
and \U$8901 ( \9884 , \2168 , \4698 );
nor \U$8902 ( \9885 , \9883 , \9884 );
xnor \U$8903 ( \9886 , \9885 , \4454 );
and \U$8904 ( \9887 , \9881 , \9886 );
and \U$8905 ( \9888 , \9877 , \9886 );
or \U$8906 ( \9889 , \9882 , \9887 , \9888 );
and \U$8907 ( \9890 , \9872 , \9889 );
and \U$8908 ( \9891 , \9856 , \9889 );
or \U$8909 ( \9892 , \9873 , \9890 , \9891 );
and \U$8910 ( \9893 , \9840 , \9892 );
and \U$8911 ( \9894 , \6825 , \1360 );
and \U$8912 ( \9895 , \6816 , \1358 );
nor \U$8913 ( \9896 , \9894 , \9895 );
xnor \U$8914 ( \9897 , \9896 , \1317 );
and \U$8915 ( \9898 , \7370 , \1247 );
and \U$8916 ( \9899 , \7168 , \1245 );
nor \U$8917 ( \9900 , \9898 , \9899 );
xnor \U$8918 ( \9901 , \9900 , \1198 );
and \U$8919 ( \9902 , \9897 , \9901 );
and \U$8920 ( \9903 , \7845 , \1146 );
and \U$8921 ( \9904 , \7673 , \1144 );
nor \U$8922 ( \9905 , \9903 , \9904 );
xnor \U$8923 ( \9906 , \9905 , \1105 );
and \U$8924 ( \9907 , \9901 , \9906 );
and \U$8925 ( \9908 , \9897 , \9906 );
or \U$8926 ( \9909 , \9902 , \9907 , \9908 );
and \U$8927 ( \9910 , \5447 , \1828 );
and \U$8928 ( \9911 , \5439 , \1826 );
nor \U$8929 ( \9912 , \9910 , \9911 );
xnor \U$8930 ( \9913 , \9912 , \1750 );
and \U$8931 ( \9914 , \5921 , \1664 );
and \U$8932 ( \9915 , \5916 , \1662 );
nor \U$8933 ( \9916 , \9914 , \9915 );
xnor \U$8934 ( \9917 , \9916 , \1570 );
and \U$8935 ( \9918 , \9913 , \9917 );
and \U$8936 ( \9919 , \6444 , \1494 );
and \U$8937 ( \9920 , \6185 , \1492 );
nor \U$8938 ( \9921 , \9919 , \9920 );
xnor \U$8939 ( \9922 , \9921 , \1422 );
and \U$8940 ( \9923 , \9917 , \9922 );
and \U$8941 ( \9924 , \9913 , \9922 );
or \U$8942 ( \9925 , \9918 , \9923 , \9924 );
and \U$8943 ( \9926 , \9909 , \9925 );
and \U$8944 ( \9927 , \4557 , \2494 );
and \U$8945 ( \9928 , \4349 , \2492 );
nor \U$8946 ( \9929 , \9927 , \9928 );
xnor \U$8947 ( \9930 , \9929 , \2338 );
and \U$8948 ( \9931 , \4684 , \2222 );
and \U$8949 ( \9932 , \4679 , \2220 );
nor \U$8950 ( \9933 , \9931 , \9932 );
xnor \U$8951 ( \9934 , \9933 , \2109 );
and \U$8952 ( \9935 , \9930 , \9934 );
and \U$8953 ( \9936 , \5137 , \2028 );
and \U$8954 ( \9937 , \4940 , \2026 );
nor \U$8955 ( \9938 , \9936 , \9937 );
xnor \U$8956 ( \9939 , \9938 , \1892 );
and \U$8957 ( \9940 , \9934 , \9939 );
and \U$8958 ( \9941 , \9930 , \9939 );
or \U$8959 ( \9942 , \9935 , \9940 , \9941 );
and \U$8960 ( \9943 , \9925 , \9942 );
and \U$8961 ( \9944 , \9909 , \9942 );
or \U$8962 ( \9945 , \9926 , \9943 , \9944 );
and \U$8963 ( \9946 , \9892 , \9945 );
and \U$8964 ( \9947 , \9840 , \9945 );
or \U$8965 ( \9948 , \9893 , \9946 , \9947 );
and \U$8966 ( \9949 , \9786 , \9948 );
xor \U$8967 ( \9950 , \9567 , \9571 );
xor \U$8968 ( \9951 , \9950 , \9576 );
xor \U$8969 ( \9952 , \9583 , \9587 );
xor \U$8970 ( \9953 , \9952 , \9592 );
and \U$8971 ( \9954 , \9951 , \9953 );
xor \U$8972 ( \9955 , \9600 , \9604 );
xor \U$8973 ( \9956 , \9955 , \9609 );
and \U$8974 ( \9957 , \9953 , \9956 );
and \U$8975 ( \9958 , \9951 , \9956 );
or \U$8976 ( \9959 , \9954 , \9957 , \9958 );
xor \U$8977 ( \9960 , \9176 , \9180 );
xor \U$8978 ( \9961 , \9960 , \9185 );
and \U$8979 ( \9962 , \9959 , \9961 );
xor \U$8980 ( \9963 , \9194 , \9198 );
xor \U$8981 ( \9964 , \9963 , \9203 );
and \U$8982 ( \9965 , \9961 , \9964 );
and \U$8983 ( \9966 , \9959 , \9964 );
or \U$8984 ( \9967 , \9962 , \9965 , \9966 );
and \U$8985 ( \9968 , \9948 , \9967 );
and \U$8986 ( \9969 , \9786 , \9967 );
or \U$8987 ( \9970 , \9949 , \9968 , \9969 );
xor \U$8988 ( \9971 , \9471 , \9487 );
xor \U$8989 ( \9972 , \9971 , \9504 );
xor \U$8990 ( \9973 , \9523 , \9539 );
xor \U$8991 ( \9974 , \9973 , \9556 );
and \U$8992 ( \9975 , \9972 , \9974 );
xor \U$8993 ( \9976 , \9579 , \9595 );
xor \U$8994 ( \9977 , \9976 , \9612 );
and \U$8995 ( \9978 , \9974 , \9977 );
and \U$8996 ( \9979 , \9972 , \9977 );
or \U$8997 ( \9980 , \9975 , \9978 , \9979 );
xor \U$8998 ( \9981 , \9620 , \9622 );
xor \U$8999 ( \9982 , \9981 , \9625 );
xor \U$9000 ( \9983 , \9630 , \9632 );
xor \U$9001 ( \9984 , \9983 , \9635 );
and \U$9002 ( \9985 , \9982 , \9984 );
xor \U$9003 ( \9986 , \9653 , \9655 );
xor \U$9004 ( \9987 , \9986 , \9658 );
and \U$9005 ( \9988 , \9984 , \9987 );
and \U$9006 ( \9989 , \9982 , \9987 );
or \U$9007 ( \9990 , \9985 , \9988 , \9989 );
and \U$9008 ( \9991 , \9980 , \9990 );
xor \U$9009 ( \9992 , \9242 , \9258 );
xor \U$9010 ( \9993 , \9992 , \9275 );
and \U$9011 ( \9994 , \9990 , \9993 );
and \U$9012 ( \9995 , \9980 , \9993 );
or \U$9013 ( \9996 , \9991 , \9994 , \9995 );
and \U$9014 ( \9997 , \9970 , \9996 );
xor \U$9015 ( \9998 , \9188 , \9206 );
xor \U$9016 ( \9999 , \9998 , \9223 );
xor \U$9017 ( \10000 , \9667 , \9669 );
xor \U$9018 ( \10001 , \10000 , \9672 );
and \U$9019 ( \10002 , \9999 , \10001 );
xor \U$9020 ( \10003 , \9680 , \9682 );
xor \U$9021 ( \10004 , \10003 , \9685 );
and \U$9022 ( \10005 , \10001 , \10004 );
and \U$9023 ( \10006 , \9999 , \10004 );
or \U$9024 ( \10007 , \10002 , \10005 , \10006 );
and \U$9025 ( \10008 , \9996 , \10007 );
and \U$9026 ( \10009 , \9970 , \10007 );
or \U$9027 ( \10010 , \9997 , \10008 , \10009 );
xor \U$9028 ( \10011 , \9618 , \9664 );
xor \U$9029 ( \10012 , \10011 , \9675 );
xor \U$9030 ( \10013 , \9688 , \9690 );
xor \U$9031 ( \10014 , \10013 , \9693 );
and \U$9032 ( \10015 , \10012 , \10014 );
xor \U$9033 ( \10016 , \9699 , \9701 );
xor \U$9034 ( \10017 , \10016 , \9704 );
and \U$9035 ( \10018 , \10014 , \10017 );
and \U$9036 ( \10019 , \10012 , \10017 );
or \U$9037 ( \10020 , \10015 , \10018 , \10019 );
and \U$9038 ( \10021 , \10010 , \10020 );
xor \U$9039 ( \10022 , \9712 , \9714 );
xor \U$9040 ( \10023 , \10022 , \9717 );
and \U$9041 ( \10024 , \10020 , \10023 );
and \U$9042 ( \10025 , \10010 , \10023 );
or \U$9043 ( \10026 , \10021 , \10024 , \10025 );
xor \U$9044 ( \10027 , \9710 , \9720 );
xor \U$9045 ( \10028 , \10027 , \9723 );
and \U$9046 ( \10029 , \10026 , \10028 );
xor \U$9047 ( \10030 , \9728 , \9730 );
and \U$9048 ( \10031 , \10028 , \10030 );
and \U$9049 ( \10032 , \10026 , \10030 );
or \U$9050 ( \10033 , \10029 , \10031 , \10032 );
xor \U$9051 ( \10034 , \9726 , \9731 );
xor \U$9052 ( \10035 , \10034 , \9734 );
and \U$9053 ( \10036 , \10033 , \10035 );
xor \U$9054 ( \10037 , \9425 , \9435 );
xor \U$9055 ( \10038 , \10037 , \9438 );
and \U$9056 ( \10039 , \10035 , \10038 );
and \U$9057 ( \10040 , \10033 , \10038 );
or \U$9058 ( \10041 , \10036 , \10039 , \10040 );
and \U$9059 ( \10042 , \9743 , \10041 );
xor \U$9060 ( \10043 , \9743 , \10041 );
xor \U$9061 ( \10044 , \10033 , \10035 );
xor \U$9062 ( \10045 , \10044 , \10038 );
and \U$9063 ( \10046 , \5916 , \1828 );
and \U$9064 ( \10047 , \5447 , \1826 );
nor \U$9065 ( \10048 , \10046 , \10047 );
xnor \U$9066 ( \10049 , \10048 , \1750 );
and \U$9067 ( \10050 , \6185 , \1664 );
and \U$9068 ( \10051 , \5921 , \1662 );
nor \U$9069 ( \10052 , \10050 , \10051 );
xnor \U$9070 ( \10053 , \10052 , \1570 );
and \U$9071 ( \10054 , \10049 , \10053 );
and \U$9072 ( \10055 , \6816 , \1494 );
and \U$9073 ( \10056 , \6444 , \1492 );
nor \U$9074 ( \10057 , \10055 , \10056 );
xnor \U$9075 ( \10058 , \10057 , \1422 );
and \U$9076 ( \10059 , \10053 , \10058 );
and \U$9077 ( \10060 , \10049 , \10058 );
or \U$9078 ( \10061 , \10054 , \10059 , \10060 );
and \U$9079 ( \10062 , \4679 , \2494 );
and \U$9080 ( \10063 , \4557 , \2492 );
nor \U$9081 ( \10064 , \10062 , \10063 );
xnor \U$9082 ( \10065 , \10064 , \2338 );
and \U$9083 ( \10066 , \4940 , \2222 );
and \U$9084 ( \10067 , \4684 , \2220 );
nor \U$9085 ( \10068 , \10066 , \10067 );
xnor \U$9086 ( \10069 , \10068 , \2109 );
and \U$9087 ( \10070 , \10065 , \10069 );
and \U$9088 ( \10071 , \5439 , \2028 );
and \U$9089 ( \10072 , \5137 , \2026 );
nor \U$9090 ( \10073 , \10071 , \10072 );
xnor \U$9091 ( \10074 , \10073 , \1892 );
and \U$9092 ( \10075 , \10069 , \10074 );
and \U$9093 ( \10076 , \10065 , \10074 );
or \U$9094 ( \10077 , \10070 , \10075 , \10076 );
and \U$9095 ( \10078 , \10061 , \10077 );
and \U$9096 ( \10079 , \7168 , \1360 );
and \U$9097 ( \10080 , \6825 , \1358 );
nor \U$9098 ( \10081 , \10079 , \10080 );
xnor \U$9099 ( \10082 , \10081 , \1317 );
and \U$9100 ( \10083 , \7673 , \1247 );
and \U$9101 ( \10084 , \7370 , \1245 );
nor \U$9102 ( \10085 , \10083 , \10084 );
xnor \U$9103 ( \10086 , \10085 , \1198 );
and \U$9104 ( \10087 , \10082 , \10086 );
and \U$9105 ( \10088 , \8371 , \1146 );
and \U$9106 ( \10089 , \7845 , \1144 );
nor \U$9107 ( \10090 , \10088 , \10089 );
xnor \U$9108 ( \10091 , \10090 , \1105 );
and \U$9109 ( \10092 , \10086 , \10091 );
and \U$9110 ( \10093 , \10082 , \10091 );
or \U$9111 ( \10094 , \10087 , \10092 , \10093 );
and \U$9112 ( \10095 , \10077 , \10094 );
and \U$9113 ( \10096 , \10061 , \10094 );
or \U$9114 ( \10097 , \10078 , \10095 , \10096 );
xor \U$9115 ( \10098 , \9190 , \9787 );
xor \U$9116 ( \10099 , \9787 , \9788 );
not \U$9117 ( \10100 , \10099 );
and \U$9118 ( \10101 , \10098 , \10100 );
and \U$9119 ( \10102 , \984 , \10101 );
not \U$9120 ( \10103 , \10102 );
xnor \U$9121 ( \10104 , \10103 , \9791 );
and \U$9122 ( \10105 , \1016 , \9564 );
and \U$9123 ( \10106 , \998 , \9562 );
nor \U$9124 ( \10107 , \10105 , \10106 );
xnor \U$9125 ( \10108 , \10107 , \9193 );
and \U$9126 ( \10109 , \10104 , \10108 );
and \U$9127 ( \10110 , \1085 , \9002 );
and \U$9128 ( \10111 , \1037 , \9000 );
nor \U$9129 ( \10112 , \10110 , \10111 );
xnor \U$9130 ( \10113 , \10112 , \8684 );
and \U$9131 ( \10114 , \10108 , \10113 );
and \U$9132 ( \10115 , \10104 , \10113 );
or \U$9133 ( \10116 , \10109 , \10114 , \10115 );
and \U$9134 ( \10117 , \1457 , \6903 );
and \U$9135 ( \10118 , \1377 , \6901 );
nor \U$9136 ( \10119 , \10117 , \10118 );
xnor \U$9137 ( \10120 , \10119 , \6563 );
and \U$9138 ( \10121 , \1593 , \6314 );
and \U$9139 ( \10122 , \1531 , \6312 );
nor \U$9140 ( \10123 , \10121 , \10122 );
xnor \U$9141 ( \10124 , \10123 , \6073 );
and \U$9142 ( \10125 , \10120 , \10124 );
and \U$9143 ( \10126 , \1854 , \5848 );
and \U$9144 ( \10127 , \1656 , \5846 );
nor \U$9145 ( \10128 , \10126 , \10127 );
xnor \U$9146 ( \10129 , \10128 , \5660 );
and \U$9147 ( \10130 , \10124 , \10129 );
and \U$9148 ( \10131 , \10120 , \10129 );
or \U$9149 ( \10132 , \10125 , \10130 , \10131 );
and \U$9150 ( \10133 , \10116 , \10132 );
and \U$9151 ( \10134 , \1162 , \8435 );
and \U$9152 ( \10135 , \1093 , \8433 );
nor \U$9153 ( \10136 , \10134 , \10135 );
xnor \U$9154 ( \10137 , \10136 , \8186 );
and \U$9155 ( \10138 , \1221 , \7906 );
and \U$9156 ( \10139 , \1167 , \7904 );
nor \U$9157 ( \10140 , \10138 , \10139 );
xnor \U$9158 ( \10141 , \10140 , \7646 );
and \U$9159 ( \10142 , \10137 , \10141 );
and \U$9160 ( \10143 , \1349 , \7412 );
and \U$9161 ( \10144 , \1272 , \7410 );
nor \U$9162 ( \10145 , \10143 , \10144 );
xnor \U$9163 ( \10146 , \10145 , \7097 );
and \U$9164 ( \10147 , \10141 , \10146 );
and \U$9165 ( \10148 , \10137 , \10146 );
or \U$9166 ( \10149 , \10142 , \10147 , \10148 );
and \U$9167 ( \10150 , \10132 , \10149 );
and \U$9168 ( \10151 , \10116 , \10149 );
or \U$9169 ( \10152 , \10133 , \10150 , \10151 );
and \U$9170 ( \10153 , \10097 , \10152 );
and \U$9171 ( \10154 , \2047 , \5474 );
and \U$9172 ( \10155 , \1942 , \5472 );
nor \U$9173 ( \10156 , \10154 , \10155 );
xnor \U$9174 ( \10157 , \10156 , \5242 );
and \U$9175 ( \10158 , \2168 , \5023 );
and \U$9176 ( \10159 , \2052 , \5021 );
nor \U$9177 ( \10160 , \10158 , \10159 );
xnor \U$9178 ( \10161 , \10160 , \4880 );
and \U$9179 ( \10162 , \10157 , \10161 );
and \U$9180 ( \10163 , \2459 , \4700 );
and \U$9181 ( \10164 , \2283 , \4698 );
nor \U$9182 ( \10165 , \10163 , \10164 );
xnor \U$9183 ( \10166 , \10165 , \4454 );
and \U$9184 ( \10167 , \10161 , \10166 );
and \U$9185 ( \10168 , \10157 , \10166 );
or \U$9186 ( \10169 , \10162 , \10167 , \10168 );
and \U$9187 ( \10170 , \3508 , \3264 );
and \U$9188 ( \10171 , \3334 , \3262 );
nor \U$9189 ( \10172 , \10170 , \10171 );
xnor \U$9190 ( \10173 , \10172 , \3122 );
and \U$9191 ( \10174 , \3813 , \2968 );
and \U$9192 ( \10175 , \3675 , \2966 );
nor \U$9193 ( \10176 , \10174 , \10175 );
xnor \U$9194 ( \10177 , \10176 , \2831 );
and \U$9195 ( \10178 , \10173 , \10177 );
and \U$9196 ( \10179 , \4349 , \2762 );
and \U$9197 ( \10180 , \3932 , \2760 );
nor \U$9198 ( \10181 , \10179 , \10180 );
xnor \U$9199 ( \10182 , \10181 , \2610 );
and \U$9200 ( \10183 , \10177 , \10182 );
and \U$9201 ( \10184 , \10173 , \10182 );
or \U$9202 ( \10185 , \10178 , \10183 , \10184 );
and \U$9203 ( \10186 , \10169 , \10185 );
and \U$9204 ( \10187 , \2710 , \4305 );
and \U$9205 ( \10188 , \2467 , \4303 );
nor \U$9206 ( \10189 , \10187 , \10188 );
xnor \U$9207 ( \10190 , \10189 , \4118 );
and \U$9208 ( \10191 , \2901 , \3992 );
and \U$9209 ( \10192 , \2715 , \3990 );
nor \U$9210 ( \10193 , \10191 , \10192 );
xnor \U$9211 ( \10194 , \10193 , \3787 );
and \U$9212 ( \10195 , \10190 , \10194 );
and \U$9213 ( \10196 , \3309 , \3586 );
and \U$9214 ( \10197 , \3045 , \3584 );
nor \U$9215 ( \10198 , \10196 , \10197 );
xnor \U$9216 ( \10199 , \10198 , \3437 );
and \U$9217 ( \10200 , \10194 , \10199 );
and \U$9218 ( \10201 , \10190 , \10199 );
or \U$9219 ( \10202 , \10195 , \10200 , \10201 );
and \U$9220 ( \10203 , \10185 , \10202 );
and \U$9221 ( \10204 , \10169 , \10202 );
or \U$9222 ( \10205 , \10186 , \10203 , \10204 );
and \U$9223 ( \10206 , \10152 , \10205 );
and \U$9224 ( \10207 , \10097 , \10205 );
or \U$9225 ( \10208 , \10153 , \10206 , \10207 );
and \U$9226 ( \10209 , \9041 , \1076 );
and \U$9227 ( \10210 , \8795 , \1074 );
nor \U$9228 ( \10211 , \10209 , \10210 );
xnor \U$9229 ( \10212 , \10211 , \1046 );
and \U$9230 ( \10213 , \9365 , \1028 );
and \U$9231 ( \10214 , \9046 , \1026 );
nor \U$9232 ( \10215 , \10213 , \10214 );
xnor \U$9233 ( \10216 , \10215 , \1009 );
and \U$9234 ( \10217 , \10212 , \10216 );
buf \U$9235 ( \10218 , RIc0dafa8_123);
and \U$9236 ( \10219 , \10218 , \991 );
and \U$9237 ( \10220 , \9649 , \989 );
nor \U$9238 ( \10221 , \10219 , \10220 );
xnor \U$9239 ( \10222 , \10221 , \996 );
and \U$9240 ( \10223 , \10216 , \10222 );
and \U$9241 ( \10224 , \10212 , \10222 );
or \U$9242 ( \10225 , \10217 , \10223 , \10224 );
buf \U$9243 ( \10226 , RIc0db020_124);
and \U$9244 ( \10227 , \10226 , \985 );
buf \U$9245 ( \10228 , \10227 );
and \U$9246 ( \10229 , \10225 , \10228 );
and \U$9247 ( \10230 , \10218 , \985 );
and \U$9248 ( \10231 , \10228 , \10230 );
and \U$9249 ( \10232 , \10225 , \10230 );
or \U$9250 ( \10233 , \10229 , \10231 , \10232 );
xor \U$9251 ( \10234 , \9768 , \9772 );
xor \U$9252 ( \10235 , \10234 , \9777 );
xor \U$9253 ( \10236 , \9897 , \9901 );
xor \U$9254 ( \10237 , \10236 , \9906 );
and \U$9255 ( \10238 , \10235 , \10237 );
xor \U$9256 ( \10239 , \9913 , \9917 );
xor \U$9257 ( \10240 , \10239 , \9922 );
and \U$9258 ( \10241 , \10237 , \10240 );
and \U$9259 ( \10242 , \10235 , \10240 );
or \U$9260 ( \10243 , \10238 , \10241 , \10242 );
and \U$9261 ( \10244 , \10233 , \10243 );
xor \U$9262 ( \10245 , \9930 , \9934 );
xor \U$9263 ( \10246 , \10245 , \9939 );
xor \U$9264 ( \10247 , \9844 , \9848 );
xor \U$9265 ( \10248 , \10247 , \9853 );
and \U$9266 ( \10249 , \10246 , \10248 );
xor \U$9267 ( \10250 , \9860 , \9864 );
xor \U$9268 ( \10251 , \10250 , \9869 );
and \U$9269 ( \10252 , \10248 , \10251 );
and \U$9270 ( \10253 , \10246 , \10251 );
or \U$9271 ( \10254 , \10249 , \10252 , \10253 );
and \U$9272 ( \10255 , \10243 , \10254 );
and \U$9273 ( \10256 , \10233 , \10254 );
or \U$9274 ( \10257 , \10244 , \10255 , \10256 );
and \U$9275 ( \10258 , \10208 , \10257 );
xor \U$9276 ( \10259 , \9808 , \9812 );
xor \U$9277 ( \10260 , \10259 , \9817 );
xor \U$9278 ( \10261 , \9825 , \9829 );
xor \U$9279 ( \10262 , \10261 , \9834 );
and \U$9280 ( \10263 , \10260 , \10262 );
xor \U$9281 ( \10264 , \9877 , \9881 );
xor \U$9282 ( \10265 , \10264 , \9886 );
and \U$9283 ( \10266 , \10262 , \10265 );
and \U$9284 ( \10267 , \10260 , \10265 );
or \U$9285 ( \10268 , \10263 , \10266 , \10267 );
xor \U$9286 ( \10269 , \9951 , \9953 );
xor \U$9287 ( \10270 , \10269 , \9956 );
and \U$9288 ( \10271 , \10268 , \10270 );
xor \U$9289 ( \10272 , \9755 , \9757 );
xor \U$9290 ( \10273 , \10272 , \9760 );
and \U$9291 ( \10274 , \10270 , \10273 );
and \U$9292 ( \10275 , \10268 , \10273 );
or \U$9293 ( \10276 , \10271 , \10274 , \10275 );
and \U$9294 ( \10277 , \10257 , \10276 );
and \U$9295 ( \10278 , \10208 , \10276 );
or \U$9296 ( \10279 , \10258 , \10277 , \10278 );
xor \U$9297 ( \10280 , \9753 , \9763 );
xor \U$9298 ( \10281 , \10280 , \9783 );
xor \U$9299 ( \10282 , \9840 , \9892 );
xor \U$9300 ( \10283 , \10282 , \9945 );
and \U$9301 ( \10284 , \10281 , \10283 );
xor \U$9302 ( \10285 , \9959 , \9961 );
xor \U$9303 ( \10286 , \10285 , \9964 );
and \U$9304 ( \10287 , \10283 , \10286 );
and \U$9305 ( \10288 , \10281 , \10286 );
or \U$9306 ( \10289 , \10284 , \10287 , \10288 );
and \U$9307 ( \10290 , \10279 , \10289 );
xor \U$9308 ( \10291 , \9909 , \9925 );
xor \U$9309 ( \10292 , \10291 , \9942 );
xor \U$9310 ( \10293 , \9745 , \9747 );
xor \U$9311 ( \10294 , \10293 , \9750 );
and \U$9312 ( \10295 , \10292 , \10294 );
xnor \U$9313 ( \10296 , \9780 , \9782 );
and \U$9314 ( \10297 , \10294 , \10296 );
and \U$9315 ( \10298 , \10292 , \10296 );
or \U$9316 ( \10299 , \10295 , \10297 , \10298 );
xor \U$9317 ( \10300 , \9972 , \9974 );
xor \U$9318 ( \10301 , \10300 , \9977 );
and \U$9319 ( \10302 , \10299 , \10301 );
xor \U$9320 ( \10303 , \9982 , \9984 );
xor \U$9321 ( \10304 , \10303 , \9987 );
and \U$9322 ( \10305 , \10301 , \10304 );
and \U$9323 ( \10306 , \10299 , \10304 );
or \U$9324 ( \10307 , \10302 , \10305 , \10306 );
and \U$9325 ( \10308 , \10289 , \10307 );
and \U$9326 ( \10309 , \10279 , \10307 );
or \U$9327 ( \10310 , \10290 , \10308 , \10309 );
xor \U$9328 ( \10311 , \9507 , \9559 );
xor \U$9329 ( \10312 , \10311 , \9615 );
xor \U$9330 ( \10313 , \9628 , \9638 );
xor \U$9331 ( \10314 , \10313 , \9661 );
and \U$9332 ( \10315 , \10312 , \10314 );
xor \U$9333 ( \10316 , \9999 , \10001 );
xor \U$9334 ( \10317 , \10316 , \10004 );
and \U$9335 ( \10318 , \10314 , \10317 );
and \U$9336 ( \10319 , \10312 , \10317 );
or \U$9337 ( \10320 , \10315 , \10318 , \10319 );
and \U$9338 ( \10321 , \10310 , \10320 );
xor \U$9339 ( \10322 , \10012 , \10014 );
xor \U$9340 ( \10323 , \10322 , \10017 );
and \U$9341 ( \10324 , \10320 , \10323 );
and \U$9342 ( \10325 , \10310 , \10323 );
or \U$9343 ( \10326 , \10321 , \10324 , \10325 );
xor \U$9344 ( \10327 , \9678 , \9696 );
xor \U$9345 ( \10328 , \10327 , \9707 );
and \U$9346 ( \10329 , \10326 , \10328 );
xor \U$9347 ( \10330 , \10010 , \10020 );
xor \U$9348 ( \10331 , \10330 , \10023 );
and \U$9349 ( \10332 , \10328 , \10331 );
and \U$9350 ( \10333 , \10326 , \10331 );
or \U$9351 ( \10334 , \10329 , \10332 , \10333 );
xor \U$9352 ( \10335 , \10026 , \10028 );
xor \U$9353 ( \10336 , \10335 , \10030 );
and \U$9354 ( \10337 , \10334 , \10336 );
and \U$9355 ( \10338 , \10045 , \10337 );
xor \U$9356 ( \10339 , \10045 , \10337 );
xor \U$9357 ( \10340 , \10334 , \10336 );
and \U$9358 ( \10341 , \3334 , \3586 );
and \U$9359 ( \10342 , \3309 , \3584 );
nor \U$9360 ( \10343 , \10341 , \10342 );
xnor \U$9361 ( \10344 , \10343 , \3437 );
and \U$9362 ( \10345 , \3675 , \3264 );
and \U$9363 ( \10346 , \3508 , \3262 );
nor \U$9364 ( \10347 , \10345 , \10346 );
xnor \U$9365 ( \10348 , \10347 , \3122 );
and \U$9366 ( \10349 , \10344 , \10348 );
and \U$9367 ( \10350 , \3932 , \2968 );
and \U$9368 ( \10351 , \3813 , \2966 );
nor \U$9369 ( \10352 , \10350 , \10351 );
xnor \U$9370 ( \10353 , \10352 , \2831 );
and \U$9371 ( \10354 , \10348 , \10353 );
and \U$9372 ( \10355 , \10344 , \10353 );
or \U$9373 ( \10356 , \10349 , \10354 , \10355 );
and \U$9374 ( \10357 , \2467 , \4700 );
and \U$9375 ( \10358 , \2459 , \4698 );
nor \U$9376 ( \10359 , \10357 , \10358 );
xnor \U$9377 ( \10360 , \10359 , \4454 );
and \U$9378 ( \10361 , \2715 , \4305 );
and \U$9379 ( \10362 , \2710 , \4303 );
nor \U$9380 ( \10363 , \10361 , \10362 );
xnor \U$9381 ( \10364 , \10363 , \4118 );
and \U$9382 ( \10365 , \10360 , \10364 );
and \U$9383 ( \10366 , \3045 , \3992 );
and \U$9384 ( \10367 , \2901 , \3990 );
nor \U$9385 ( \10368 , \10366 , \10367 );
xnor \U$9386 ( \10369 , \10368 , \3787 );
and \U$9387 ( \10370 , \10364 , \10369 );
and \U$9388 ( \10371 , \10360 , \10369 );
or \U$9389 ( \10372 , \10365 , \10370 , \10371 );
and \U$9390 ( \10373 , \10356 , \10372 );
and \U$9391 ( \10374 , \1942 , \5848 );
and \U$9392 ( \10375 , \1854 , \5846 );
nor \U$9393 ( \10376 , \10374 , \10375 );
xnor \U$9394 ( \10377 , \10376 , \5660 );
and \U$9395 ( \10378 , \2052 , \5474 );
and \U$9396 ( \10379 , \2047 , \5472 );
nor \U$9397 ( \10380 , \10378 , \10379 );
xnor \U$9398 ( \10381 , \10380 , \5242 );
and \U$9399 ( \10382 , \10377 , \10381 );
and \U$9400 ( \10383 , \2283 , \5023 );
and \U$9401 ( \10384 , \2168 , \5021 );
nor \U$9402 ( \10385 , \10383 , \10384 );
xnor \U$9403 ( \10386 , \10385 , \4880 );
and \U$9404 ( \10387 , \10381 , \10386 );
and \U$9405 ( \10388 , \10377 , \10386 );
or \U$9406 ( \10389 , \10382 , \10387 , \10388 );
and \U$9407 ( \10390 , \10372 , \10389 );
and \U$9408 ( \10391 , \10356 , \10389 );
or \U$9409 ( \10392 , \10373 , \10390 , \10391 );
and \U$9410 ( \10393 , \1377 , \7412 );
and \U$9411 ( \10394 , \1349 , \7410 );
nor \U$9412 ( \10395 , \10393 , \10394 );
xnor \U$9413 ( \10396 , \10395 , \7097 );
and \U$9414 ( \10397 , \1531 , \6903 );
and \U$9415 ( \10398 , \1457 , \6901 );
nor \U$9416 ( \10399 , \10397 , \10398 );
xnor \U$9417 ( \10400 , \10399 , \6563 );
and \U$9418 ( \10401 , \10396 , \10400 );
and \U$9419 ( \10402 , \1656 , \6314 );
and \U$9420 ( \10403 , \1593 , \6312 );
nor \U$9421 ( \10404 , \10402 , \10403 );
xnor \U$9422 ( \10405 , \10404 , \6073 );
and \U$9423 ( \10406 , \10400 , \10405 );
and \U$9424 ( \10407 , \10396 , \10405 );
or \U$9425 ( \10408 , \10401 , \10406 , \10407 );
and \U$9426 ( \10409 , \1093 , \9002 );
and \U$9427 ( \10410 , \1085 , \9000 );
nor \U$9428 ( \10411 , \10409 , \10410 );
xnor \U$9429 ( \10412 , \10411 , \8684 );
and \U$9430 ( \10413 , \1167 , \8435 );
and \U$9431 ( \10414 , \1162 , \8433 );
nor \U$9432 ( \10415 , \10413 , \10414 );
xnor \U$9433 ( \10416 , \10415 , \8186 );
and \U$9434 ( \10417 , \10412 , \10416 );
and \U$9435 ( \10418 , \1272 , \7906 );
and \U$9436 ( \10419 , \1221 , \7904 );
nor \U$9437 ( \10420 , \10418 , \10419 );
xnor \U$9438 ( \10421 , \10420 , \7646 );
and \U$9439 ( \10422 , \10416 , \10421 );
and \U$9440 ( \10423 , \10412 , \10421 );
or \U$9441 ( \10424 , \10417 , \10422 , \10423 );
and \U$9442 ( \10425 , \10408 , \10424 );
buf \U$9443 ( \10426 , RIc0d9310_62);
buf \U$9444 ( \10427 , RIc0d9388_63);
and \U$9445 ( \10428 , \10426 , \10427 );
not \U$9446 ( \10429 , \10428 );
and \U$9447 ( \10430 , \9788 , \10429 );
not \U$9448 ( \10431 , \10430 );
and \U$9449 ( \10432 , \998 , \10101 );
and \U$9450 ( \10433 , \984 , \10099 );
nor \U$9451 ( \10434 , \10432 , \10433 );
xnor \U$9452 ( \10435 , \10434 , \9791 );
and \U$9453 ( \10436 , \10431 , \10435 );
and \U$9454 ( \10437 , \1037 , \9564 );
and \U$9455 ( \10438 , \1016 , \9562 );
nor \U$9456 ( \10439 , \10437 , \10438 );
xnor \U$9457 ( \10440 , \10439 , \9193 );
and \U$9458 ( \10441 , \10435 , \10440 );
and \U$9459 ( \10442 , \10431 , \10440 );
or \U$9460 ( \10443 , \10436 , \10441 , \10442 );
and \U$9461 ( \10444 , \10424 , \10443 );
and \U$9462 ( \10445 , \10408 , \10443 );
or \U$9463 ( \10446 , \10425 , \10444 , \10445 );
and \U$9464 ( \10447 , \10392 , \10446 );
and \U$9465 ( \10448 , \6825 , \1494 );
and \U$9466 ( \10449 , \6816 , \1492 );
nor \U$9467 ( \10450 , \10448 , \10449 );
xnor \U$9468 ( \10451 , \10450 , \1422 );
and \U$9469 ( \10452 , \7370 , \1360 );
and \U$9470 ( \10453 , \7168 , \1358 );
nor \U$9471 ( \10454 , \10452 , \10453 );
xnor \U$9472 ( \10455 , \10454 , \1317 );
and \U$9473 ( \10456 , \10451 , \10455 );
and \U$9474 ( \10457 , \7845 , \1247 );
and \U$9475 ( \10458 , \7673 , \1245 );
nor \U$9476 ( \10459 , \10457 , \10458 );
xnor \U$9477 ( \10460 , \10459 , \1198 );
and \U$9478 ( \10461 , \10455 , \10460 );
and \U$9479 ( \10462 , \10451 , \10460 );
or \U$9480 ( \10463 , \10456 , \10461 , \10462 );
and \U$9481 ( \10464 , \5447 , \2028 );
and \U$9482 ( \10465 , \5439 , \2026 );
nor \U$9483 ( \10466 , \10464 , \10465 );
xnor \U$9484 ( \10467 , \10466 , \1892 );
and \U$9485 ( \10468 , \5921 , \1828 );
and \U$9486 ( \10469 , \5916 , \1826 );
nor \U$9487 ( \10470 , \10468 , \10469 );
xnor \U$9488 ( \10471 , \10470 , \1750 );
and \U$9489 ( \10472 , \10467 , \10471 );
and \U$9490 ( \10473 , \6444 , \1664 );
and \U$9491 ( \10474 , \6185 , \1662 );
nor \U$9492 ( \10475 , \10473 , \10474 );
xnor \U$9493 ( \10476 , \10475 , \1570 );
and \U$9494 ( \10477 , \10471 , \10476 );
and \U$9495 ( \10478 , \10467 , \10476 );
or \U$9496 ( \10479 , \10472 , \10477 , \10478 );
and \U$9497 ( \10480 , \10463 , \10479 );
and \U$9498 ( \10481 , \4557 , \2762 );
and \U$9499 ( \10482 , \4349 , \2760 );
nor \U$9500 ( \10483 , \10481 , \10482 );
xnor \U$9501 ( \10484 , \10483 , \2610 );
and \U$9502 ( \10485 , \4684 , \2494 );
and \U$9503 ( \10486 , \4679 , \2492 );
nor \U$9504 ( \10487 , \10485 , \10486 );
xnor \U$9505 ( \10488 , \10487 , \2338 );
and \U$9506 ( \10489 , \10484 , \10488 );
and \U$9507 ( \10490 , \5137 , \2222 );
and \U$9508 ( \10491 , \4940 , \2220 );
nor \U$9509 ( \10492 , \10490 , \10491 );
xnor \U$9510 ( \10493 , \10492 , \2109 );
and \U$9511 ( \10494 , \10488 , \10493 );
and \U$9512 ( \10495 , \10484 , \10493 );
or \U$9513 ( \10496 , \10489 , \10494 , \10495 );
and \U$9514 ( \10497 , \10479 , \10496 );
and \U$9515 ( \10498 , \10463 , \10496 );
or \U$9516 ( \10499 , \10480 , \10497 , \10498 );
and \U$9517 ( \10500 , \10446 , \10499 );
and \U$9518 ( \10501 , \10392 , \10499 );
or \U$9519 ( \10502 , \10447 , \10500 , \10501 );
xor \U$9520 ( \10503 , \10157 , \10161 );
xor \U$9521 ( \10504 , \10503 , \10166 );
xor \U$9522 ( \10505 , \10173 , \10177 );
xor \U$9523 ( \10506 , \10505 , \10182 );
and \U$9524 ( \10507 , \10504 , \10506 );
xor \U$9525 ( \10508 , \10190 , \10194 );
xor \U$9526 ( \10509 , \10508 , \10199 );
and \U$9527 ( \10510 , \10506 , \10509 );
and \U$9528 ( \10511 , \10504 , \10509 );
or \U$9529 ( \10512 , \10507 , \10510 , \10511 );
xor \U$9530 ( \10513 , \10049 , \10053 );
xor \U$9531 ( \10514 , \10513 , \10058 );
xor \U$9532 ( \10515 , \10065 , \10069 );
xor \U$9533 ( \10516 , \10515 , \10074 );
and \U$9534 ( \10517 , \10514 , \10516 );
xor \U$9535 ( \10518 , \10082 , \10086 );
xor \U$9536 ( \10519 , \10518 , \10091 );
and \U$9537 ( \10520 , \10516 , \10519 );
and \U$9538 ( \10521 , \10514 , \10519 );
or \U$9539 ( \10522 , \10517 , \10520 , \10521 );
and \U$9540 ( \10523 , \10512 , \10522 );
and \U$9541 ( \10524 , \8795 , \1146 );
and \U$9542 ( \10525 , \8371 , \1144 );
nor \U$9543 ( \10526 , \10524 , \10525 );
xnor \U$9544 ( \10527 , \10526 , \1105 );
and \U$9545 ( \10528 , \9046 , \1076 );
and \U$9546 ( \10529 , \9041 , \1074 );
nor \U$9547 ( \10530 , \10528 , \10529 );
xnor \U$9548 ( \10531 , \10530 , \1046 );
and \U$9549 ( \10532 , \10527 , \10531 );
and \U$9550 ( \10533 , \9649 , \1028 );
and \U$9551 ( \10534 , \9365 , \1026 );
nor \U$9552 ( \10535 , \10533 , \10534 );
xnor \U$9553 ( \10536 , \10535 , \1009 );
and \U$9554 ( \10537 , \10531 , \10536 );
and \U$9555 ( \10538 , \10527 , \10536 );
or \U$9556 ( \10539 , \10532 , \10537 , \10538 );
xor \U$9557 ( \10540 , \10212 , \10216 );
xor \U$9558 ( \10541 , \10540 , \10222 );
and \U$9559 ( \10542 , \10539 , \10541 );
not \U$9560 ( \10543 , \10227 );
and \U$9561 ( \10544 , \10541 , \10543 );
and \U$9562 ( \10545 , \10539 , \10543 );
or \U$9563 ( \10546 , \10542 , \10544 , \10545 );
and \U$9564 ( \10547 , \10522 , \10546 );
and \U$9565 ( \10548 , \10512 , \10546 );
or \U$9566 ( \10549 , \10523 , \10547 , \10548 );
and \U$9567 ( \10550 , \10502 , \10549 );
xor \U$9568 ( \10551 , \10104 , \10108 );
xor \U$9569 ( \10552 , \10551 , \10113 );
xor \U$9570 ( \10553 , \10120 , \10124 );
xor \U$9571 ( \10554 , \10553 , \10129 );
and \U$9572 ( \10555 , \10552 , \10554 );
xor \U$9573 ( \10556 , \10137 , \10141 );
xor \U$9574 ( \10557 , \10556 , \10146 );
and \U$9575 ( \10558 , \10554 , \10557 );
and \U$9576 ( \10559 , \10552 , \10557 );
or \U$9577 ( \10560 , \10555 , \10558 , \10559 );
xor \U$9578 ( \10561 , \9792 , \9796 );
xor \U$9579 ( \10562 , \10561 , \9801 );
and \U$9580 ( \10563 , \10560 , \10562 );
xor \U$9581 ( \10564 , \10260 , \10262 );
xor \U$9582 ( \10565 , \10564 , \10265 );
and \U$9583 ( \10566 , \10562 , \10565 );
and \U$9584 ( \10567 , \10560 , \10565 );
or \U$9585 ( \10568 , \10563 , \10566 , \10567 );
and \U$9586 ( \10569 , \10549 , \10568 );
and \U$9587 ( \10570 , \10502 , \10568 );
or \U$9588 ( \10571 , \10550 , \10569 , \10570 );
xor \U$9589 ( \10572 , \10061 , \10077 );
xor \U$9590 ( \10573 , \10572 , \10094 );
xor \U$9591 ( \10574 , \10116 , \10132 );
xor \U$9592 ( \10575 , \10574 , \10149 );
and \U$9593 ( \10576 , \10573 , \10575 );
xor \U$9594 ( \10577 , \10169 , \10185 );
xor \U$9595 ( \10578 , \10577 , \10202 );
and \U$9596 ( \10579 , \10575 , \10578 );
and \U$9597 ( \10580 , \10573 , \10578 );
or \U$9598 ( \10581 , \10576 , \10579 , \10580 );
xor \U$9599 ( \10582 , \10225 , \10228 );
xor \U$9600 ( \10583 , \10582 , \10230 );
xor \U$9601 ( \10584 , \10235 , \10237 );
xor \U$9602 ( \10585 , \10584 , \10240 );
and \U$9603 ( \10586 , \10583 , \10585 );
xor \U$9604 ( \10587 , \10246 , \10248 );
xor \U$9605 ( \10588 , \10587 , \10251 );
and \U$9606 ( \10589 , \10585 , \10588 );
and \U$9607 ( \10590 , \10583 , \10588 );
or \U$9608 ( \10591 , \10586 , \10589 , \10590 );
and \U$9609 ( \10592 , \10581 , \10591 );
xor \U$9610 ( \10593 , \9856 , \9872 );
xor \U$9611 ( \10594 , \10593 , \9889 );
and \U$9612 ( \10595 , \10591 , \10594 );
and \U$9613 ( \10596 , \10581 , \10594 );
or \U$9614 ( \10597 , \10592 , \10595 , \10596 );
and \U$9615 ( \10598 , \10571 , \10597 );
xor \U$9616 ( \10599 , \9804 , \9820 );
xor \U$9617 ( \10600 , \10599 , \9837 );
xor \U$9618 ( \10601 , \10268 , \10270 );
xor \U$9619 ( \10602 , \10601 , \10273 );
and \U$9620 ( \10603 , \10600 , \10602 );
xor \U$9621 ( \10604 , \10292 , \10294 );
xor \U$9622 ( \10605 , \10604 , \10296 );
and \U$9623 ( \10606 , \10602 , \10605 );
and \U$9624 ( \10607 , \10600 , \10605 );
or \U$9625 ( \10608 , \10603 , \10606 , \10607 );
and \U$9626 ( \10609 , \10597 , \10608 );
and \U$9627 ( \10610 , \10571 , \10608 );
or \U$9628 ( \10611 , \10598 , \10609 , \10610 );
xor \U$9629 ( \10612 , \10208 , \10257 );
xor \U$9630 ( \10613 , \10612 , \10276 );
xor \U$9631 ( \10614 , \10281 , \10283 );
xor \U$9632 ( \10615 , \10614 , \10286 );
and \U$9633 ( \10616 , \10613 , \10615 );
xor \U$9634 ( \10617 , \10299 , \10301 );
xor \U$9635 ( \10618 , \10617 , \10304 );
and \U$9636 ( \10619 , \10615 , \10618 );
and \U$9637 ( \10620 , \10613 , \10618 );
or \U$9638 ( \10621 , \10616 , \10619 , \10620 );
and \U$9639 ( \10622 , \10611 , \10621 );
xor \U$9640 ( \10623 , \9980 , \9990 );
xor \U$9641 ( \10624 , \10623 , \9993 );
and \U$9642 ( \10625 , \10621 , \10624 );
and \U$9643 ( \10626 , \10611 , \10624 );
or \U$9644 ( \10627 , \10622 , \10625 , \10626 );
xor \U$9645 ( \10628 , \9786 , \9948 );
xor \U$9646 ( \10629 , \10628 , \9967 );
xor \U$9647 ( \10630 , \10279 , \10289 );
xor \U$9648 ( \10631 , \10630 , \10307 );
and \U$9649 ( \10632 , \10629 , \10631 );
xor \U$9650 ( \10633 , \10312 , \10314 );
xor \U$9651 ( \10634 , \10633 , \10317 );
and \U$9652 ( \10635 , \10631 , \10634 );
and \U$9653 ( \10636 , \10629 , \10634 );
or \U$9654 ( \10637 , \10632 , \10635 , \10636 );
and \U$9655 ( \10638 , \10627 , \10637 );
xor \U$9656 ( \10639 , \9970 , \9996 );
xor \U$9657 ( \10640 , \10639 , \10007 );
and \U$9658 ( \10641 , \10637 , \10640 );
and \U$9659 ( \10642 , \10627 , \10640 );
or \U$9660 ( \10643 , \10638 , \10641 , \10642 );
xor \U$9661 ( \10644 , \10326 , \10328 );
xor \U$9662 ( \10645 , \10644 , \10331 );
and \U$9663 ( \10646 , \10643 , \10645 );
and \U$9664 ( \10647 , \10340 , \10646 );
xor \U$9665 ( \10648 , \10340 , \10646 );
xor \U$9666 ( \10649 , \10643 , \10645 );
and \U$9667 ( \10650 , \1457 , \7412 );
and \U$9668 ( \10651 , \1377 , \7410 );
nor \U$9669 ( \10652 , \10650 , \10651 );
xnor \U$9670 ( \10653 , \10652 , \7097 );
and \U$9671 ( \10654 , \1593 , \6903 );
and \U$9672 ( \10655 , \1531 , \6901 );
nor \U$9673 ( \10656 , \10654 , \10655 );
xnor \U$9674 ( \10657 , \10656 , \6563 );
and \U$9675 ( \10658 , \10653 , \10657 );
and \U$9676 ( \10659 , \1854 , \6314 );
and \U$9677 ( \10660 , \1656 , \6312 );
nor \U$9678 ( \10661 , \10659 , \10660 );
xnor \U$9679 ( \10662 , \10661 , \6073 );
and \U$9680 ( \10663 , \10657 , \10662 );
and \U$9681 ( \10664 , \10653 , \10662 );
or \U$9682 ( \10665 , \10658 , \10663 , \10664 );
xor \U$9683 ( \10666 , \9788 , \10426 );
xor \U$9684 ( \10667 , \10426 , \10427 );
not \U$9685 ( \10668 , \10667 );
and \U$9686 ( \10669 , \10666 , \10668 );
and \U$9687 ( \10670 , \984 , \10669 );
not \U$9688 ( \10671 , \10670 );
xnor \U$9689 ( \10672 , \10671 , \10430 );
and \U$9690 ( \10673 , \1016 , \10101 );
and \U$9691 ( \10674 , \998 , \10099 );
nor \U$9692 ( \10675 , \10673 , \10674 );
xnor \U$9693 ( \10676 , \10675 , \9791 );
and \U$9694 ( \10677 , \10672 , \10676 );
and \U$9695 ( \10678 , \1085 , \9564 );
and \U$9696 ( \10679 , \1037 , \9562 );
nor \U$9697 ( \10680 , \10678 , \10679 );
xnor \U$9698 ( \10681 , \10680 , \9193 );
and \U$9699 ( \10682 , \10676 , \10681 );
and \U$9700 ( \10683 , \10672 , \10681 );
or \U$9701 ( \10684 , \10677 , \10682 , \10683 );
and \U$9702 ( \10685 , \10665 , \10684 );
and \U$9703 ( \10686 , \1162 , \9002 );
and \U$9704 ( \10687 , \1093 , \9000 );
nor \U$9705 ( \10688 , \10686 , \10687 );
xnor \U$9706 ( \10689 , \10688 , \8684 );
and \U$9707 ( \10690 , \1221 , \8435 );
and \U$9708 ( \10691 , \1167 , \8433 );
nor \U$9709 ( \10692 , \10690 , \10691 );
xnor \U$9710 ( \10693 , \10692 , \8186 );
and \U$9711 ( \10694 , \10689 , \10693 );
and \U$9712 ( \10695 , \1349 , \7906 );
and \U$9713 ( \10696 , \1272 , \7904 );
nor \U$9714 ( \10697 , \10695 , \10696 );
xnor \U$9715 ( \10698 , \10697 , \7646 );
and \U$9716 ( \10699 , \10693 , \10698 );
and \U$9717 ( \10700 , \10689 , \10698 );
or \U$9718 ( \10701 , \10694 , \10699 , \10700 );
and \U$9719 ( \10702 , \10684 , \10701 );
and \U$9720 ( \10703 , \10665 , \10701 );
or \U$9721 ( \10704 , \10685 , \10702 , \10703 );
and \U$9722 ( \10705 , \7168 , \1494 );
and \U$9723 ( \10706 , \6825 , \1492 );
nor \U$9724 ( \10707 , \10705 , \10706 );
xnor \U$9725 ( \10708 , \10707 , \1422 );
and \U$9726 ( \10709 , \7673 , \1360 );
and \U$9727 ( \10710 , \7370 , \1358 );
nor \U$9728 ( \10711 , \10709 , \10710 );
xnor \U$9729 ( \10712 , \10711 , \1317 );
and \U$9730 ( \10713 , \10708 , \10712 );
and \U$9731 ( \10714 , \8371 , \1247 );
and \U$9732 ( \10715 , \7845 , \1245 );
nor \U$9733 ( \10716 , \10714 , \10715 );
xnor \U$9734 ( \10717 , \10716 , \1198 );
and \U$9735 ( \10718 , \10712 , \10717 );
and \U$9736 ( \10719 , \10708 , \10717 );
or \U$9737 ( \10720 , \10713 , \10718 , \10719 );
and \U$9738 ( \10721 , \4679 , \2762 );
and \U$9739 ( \10722 , \4557 , \2760 );
nor \U$9740 ( \10723 , \10721 , \10722 );
xnor \U$9741 ( \10724 , \10723 , \2610 );
and \U$9742 ( \10725 , \4940 , \2494 );
and \U$9743 ( \10726 , \4684 , \2492 );
nor \U$9744 ( \10727 , \10725 , \10726 );
xnor \U$9745 ( \10728 , \10727 , \2338 );
and \U$9746 ( \10729 , \10724 , \10728 );
and \U$9747 ( \10730 , \5439 , \2222 );
and \U$9748 ( \10731 , \5137 , \2220 );
nor \U$9749 ( \10732 , \10730 , \10731 );
xnor \U$9750 ( \10733 , \10732 , \2109 );
and \U$9751 ( \10734 , \10728 , \10733 );
and \U$9752 ( \10735 , \10724 , \10733 );
or \U$9753 ( \10736 , \10729 , \10734 , \10735 );
and \U$9754 ( \10737 , \10720 , \10736 );
and \U$9755 ( \10738 , \5916 , \2028 );
and \U$9756 ( \10739 , \5447 , \2026 );
nor \U$9757 ( \10740 , \10738 , \10739 );
xnor \U$9758 ( \10741 , \10740 , \1892 );
and \U$9759 ( \10742 , \6185 , \1828 );
and \U$9760 ( \10743 , \5921 , \1826 );
nor \U$9761 ( \10744 , \10742 , \10743 );
xnor \U$9762 ( \10745 , \10744 , \1750 );
and \U$9763 ( \10746 , \10741 , \10745 );
and \U$9764 ( \10747 , \6816 , \1664 );
and \U$9765 ( \10748 , \6444 , \1662 );
nor \U$9766 ( \10749 , \10747 , \10748 );
xnor \U$9767 ( \10750 , \10749 , \1570 );
and \U$9768 ( \10751 , \10745 , \10750 );
and \U$9769 ( \10752 , \10741 , \10750 );
or \U$9770 ( \10753 , \10746 , \10751 , \10752 );
and \U$9771 ( \10754 , \10736 , \10753 );
and \U$9772 ( \10755 , \10720 , \10753 );
or \U$9773 ( \10756 , \10737 , \10754 , \10755 );
and \U$9774 ( \10757 , \10704 , \10756 );
and \U$9775 ( \10758 , \2047 , \5848 );
and \U$9776 ( \10759 , \1942 , \5846 );
nor \U$9777 ( \10760 , \10758 , \10759 );
xnor \U$9778 ( \10761 , \10760 , \5660 );
and \U$9779 ( \10762 , \2168 , \5474 );
and \U$9780 ( \10763 , \2052 , \5472 );
nor \U$9781 ( \10764 , \10762 , \10763 );
xnor \U$9782 ( \10765 , \10764 , \5242 );
and \U$9783 ( \10766 , \10761 , \10765 );
and \U$9784 ( \10767 , \2459 , \5023 );
and \U$9785 ( \10768 , \2283 , \5021 );
nor \U$9786 ( \10769 , \10767 , \10768 );
xnor \U$9787 ( \10770 , \10769 , \4880 );
and \U$9788 ( \10771 , \10765 , \10770 );
and \U$9789 ( \10772 , \10761 , \10770 );
or \U$9790 ( \10773 , \10766 , \10771 , \10772 );
and \U$9791 ( \10774 , \3508 , \3586 );
and \U$9792 ( \10775 , \3334 , \3584 );
nor \U$9793 ( \10776 , \10774 , \10775 );
xnor \U$9794 ( \10777 , \10776 , \3437 );
and \U$9795 ( \10778 , \3813 , \3264 );
and \U$9796 ( \10779 , \3675 , \3262 );
nor \U$9797 ( \10780 , \10778 , \10779 );
xnor \U$9798 ( \10781 , \10780 , \3122 );
and \U$9799 ( \10782 , \10777 , \10781 );
and \U$9800 ( \10783 , \4349 , \2968 );
and \U$9801 ( \10784 , \3932 , \2966 );
nor \U$9802 ( \10785 , \10783 , \10784 );
xnor \U$9803 ( \10786 , \10785 , \2831 );
and \U$9804 ( \10787 , \10781 , \10786 );
and \U$9805 ( \10788 , \10777 , \10786 );
or \U$9806 ( \10789 , \10782 , \10787 , \10788 );
and \U$9807 ( \10790 , \10773 , \10789 );
and \U$9808 ( \10791 , \2710 , \4700 );
and \U$9809 ( \10792 , \2467 , \4698 );
nor \U$9810 ( \10793 , \10791 , \10792 );
xnor \U$9811 ( \10794 , \10793 , \4454 );
and \U$9812 ( \10795 , \2901 , \4305 );
and \U$9813 ( \10796 , \2715 , \4303 );
nor \U$9814 ( \10797 , \10795 , \10796 );
xnor \U$9815 ( \10798 , \10797 , \4118 );
and \U$9816 ( \10799 , \10794 , \10798 );
and \U$9817 ( \10800 , \3309 , \3992 );
and \U$9818 ( \10801 , \3045 , \3990 );
nor \U$9819 ( \10802 , \10800 , \10801 );
xnor \U$9820 ( \10803 , \10802 , \3787 );
and \U$9821 ( \10804 , \10798 , \10803 );
and \U$9822 ( \10805 , \10794 , \10803 );
or \U$9823 ( \10806 , \10799 , \10804 , \10805 );
and \U$9824 ( \10807 , \10789 , \10806 );
and \U$9825 ( \10808 , \10773 , \10806 );
or \U$9826 ( \10809 , \10790 , \10807 , \10808 );
and \U$9827 ( \10810 , \10756 , \10809 );
and \U$9828 ( \10811 , \10704 , \10809 );
or \U$9829 ( \10812 , \10757 , \10810 , \10811 );
and \U$9830 ( \10813 , \9041 , \1146 );
and \U$9831 ( \10814 , \8795 , \1144 );
nor \U$9832 ( \10815 , \10813 , \10814 );
xnor \U$9833 ( \10816 , \10815 , \1105 );
and \U$9834 ( \10817 , \9365 , \1076 );
and \U$9835 ( \10818 , \9046 , \1074 );
nor \U$9836 ( \10819 , \10817 , \10818 );
xnor \U$9837 ( \10820 , \10819 , \1046 );
and \U$9838 ( \10821 , \10816 , \10820 );
and \U$9839 ( \10822 , \10218 , \1028 );
and \U$9840 ( \10823 , \9649 , \1026 );
nor \U$9841 ( \10824 , \10822 , \10823 );
xnor \U$9842 ( \10825 , \10824 , \1009 );
and \U$9843 ( \10826 , \10820 , \10825 );
and \U$9844 ( \10827 , \10816 , \10825 );
or \U$9845 ( \10828 , \10821 , \10826 , \10827 );
buf \U$9846 ( \10829 , RIc0db098_125);
and \U$9847 ( \10830 , \10829 , \991 );
and \U$9848 ( \10831 , \10226 , \989 );
nor \U$9849 ( \10832 , \10830 , \10831 );
xnor \U$9850 ( \10833 , \10832 , \996 );
buf \U$9851 ( \10834 , RIc0db110_126);
and \U$9852 ( \10835 , \10834 , \985 );
or \U$9853 ( \10836 , \10833 , \10835 );
and \U$9854 ( \10837 , \10828 , \10836 );
and \U$9855 ( \10838 , \10226 , \991 );
and \U$9856 ( \10839 , \10218 , \989 );
nor \U$9857 ( \10840 , \10838 , \10839 );
xnor \U$9858 ( \10841 , \10840 , \996 );
and \U$9859 ( \10842 , \10836 , \10841 );
and \U$9860 ( \10843 , \10828 , \10841 );
or \U$9861 ( \10844 , \10837 , \10842 , \10843 );
and \U$9862 ( \10845 , \10829 , \985 );
xor \U$9863 ( \10846 , \10451 , \10455 );
xor \U$9864 ( \10847 , \10846 , \10460 );
and \U$9865 ( \10848 , \10845 , \10847 );
xor \U$9866 ( \10849 , \10527 , \10531 );
xor \U$9867 ( \10850 , \10849 , \10536 );
and \U$9868 ( \10851 , \10847 , \10850 );
and \U$9869 ( \10852 , \10845 , \10850 );
or \U$9870 ( \10853 , \10848 , \10851 , \10852 );
and \U$9871 ( \10854 , \10844 , \10853 );
xor \U$9872 ( \10855 , \10344 , \10348 );
xor \U$9873 ( \10856 , \10855 , \10353 );
xor \U$9874 ( \10857 , \10467 , \10471 );
xor \U$9875 ( \10858 , \10857 , \10476 );
and \U$9876 ( \10859 , \10856 , \10858 );
xor \U$9877 ( \10860 , \10484 , \10488 );
xor \U$9878 ( \10861 , \10860 , \10493 );
and \U$9879 ( \10862 , \10858 , \10861 );
and \U$9880 ( \10863 , \10856 , \10861 );
or \U$9881 ( \10864 , \10859 , \10862 , \10863 );
and \U$9882 ( \10865 , \10853 , \10864 );
and \U$9883 ( \10866 , \10844 , \10864 );
or \U$9884 ( \10867 , \10854 , \10865 , \10866 );
and \U$9885 ( \10868 , \10812 , \10867 );
xor \U$9886 ( \10869 , \10396 , \10400 );
xor \U$9887 ( \10870 , \10869 , \10405 );
xor \U$9888 ( \10871 , \10360 , \10364 );
xor \U$9889 ( \10872 , \10871 , \10369 );
and \U$9890 ( \10873 , \10870 , \10872 );
xor \U$9891 ( \10874 , \10377 , \10381 );
xor \U$9892 ( \10875 , \10874 , \10386 );
and \U$9893 ( \10876 , \10872 , \10875 );
and \U$9894 ( \10877 , \10870 , \10875 );
or \U$9895 ( \10878 , \10873 , \10876 , \10877 );
xor \U$9896 ( \10879 , \10412 , \10416 );
xor \U$9897 ( \10880 , \10879 , \10421 );
xor \U$9898 ( \10881 , \10431 , \10435 );
xor \U$9899 ( \10882 , \10881 , \10440 );
and \U$9900 ( \10883 , \10880 , \10882 );
and \U$9901 ( \10884 , \10878 , \10883 );
xor \U$9902 ( \10885 , \10552 , \10554 );
xor \U$9903 ( \10886 , \10885 , \10557 );
and \U$9904 ( \10887 , \10883 , \10886 );
and \U$9905 ( \10888 , \10878 , \10886 );
or \U$9906 ( \10889 , \10884 , \10887 , \10888 );
and \U$9907 ( \10890 , \10867 , \10889 );
and \U$9908 ( \10891 , \10812 , \10889 );
or \U$9909 ( \10892 , \10868 , \10890 , \10891 );
xor \U$9910 ( \10893 , \10356 , \10372 );
xor \U$9911 ( \10894 , \10893 , \10389 );
xor \U$9912 ( \10895 , \10408 , \10424 );
xor \U$9913 ( \10896 , \10895 , \10443 );
and \U$9914 ( \10897 , \10894 , \10896 );
xor \U$9915 ( \10898 , \10463 , \10479 );
xor \U$9916 ( \10899 , \10898 , \10496 );
and \U$9917 ( \10900 , \10896 , \10899 );
and \U$9918 ( \10901 , \10894 , \10899 );
or \U$9919 ( \10902 , \10897 , \10900 , \10901 );
xor \U$9920 ( \10903 , \10504 , \10506 );
xor \U$9921 ( \10904 , \10903 , \10509 );
xor \U$9922 ( \10905 , \10514 , \10516 );
xor \U$9923 ( \10906 , \10905 , \10519 );
and \U$9924 ( \10907 , \10904 , \10906 );
xor \U$9925 ( \10908 , \10539 , \10541 );
xor \U$9926 ( \10909 , \10908 , \10543 );
and \U$9927 ( \10910 , \10906 , \10909 );
and \U$9928 ( \10911 , \10904 , \10909 );
or \U$9929 ( \10912 , \10907 , \10910 , \10911 );
and \U$9930 ( \10913 , \10902 , \10912 );
xor \U$9931 ( \10914 , \10573 , \10575 );
xor \U$9932 ( \10915 , \10914 , \10578 );
and \U$9933 ( \10916 , \10912 , \10915 );
and \U$9934 ( \10917 , \10902 , \10915 );
or \U$9935 ( \10918 , \10913 , \10916 , \10917 );
and \U$9936 ( \10919 , \10892 , \10918 );
xor \U$9937 ( \10920 , \10512 , \10522 );
xor \U$9938 ( \10921 , \10920 , \10546 );
xor \U$9939 ( \10922 , \10583 , \10585 );
xor \U$9940 ( \10923 , \10922 , \10588 );
and \U$9941 ( \10924 , \10921 , \10923 );
xor \U$9942 ( \10925 , \10560 , \10562 );
xor \U$9943 ( \10926 , \10925 , \10565 );
and \U$9944 ( \10927 , \10923 , \10926 );
and \U$9945 ( \10928 , \10921 , \10926 );
or \U$9946 ( \10929 , \10924 , \10927 , \10928 );
and \U$9947 ( \10930 , \10918 , \10929 );
and \U$9948 ( \10931 , \10892 , \10929 );
or \U$9949 ( \10932 , \10919 , \10930 , \10931 );
xor \U$9950 ( \10933 , \10097 , \10152 );
xor \U$9951 ( \10934 , \10933 , \10205 );
xor \U$9952 ( \10935 , \10233 , \10243 );
xor \U$9953 ( \10936 , \10935 , \10254 );
and \U$9954 ( \10937 , \10934 , \10936 );
xor \U$9955 ( \10938 , \10600 , \10602 );
xor \U$9956 ( \10939 , \10938 , \10605 );
and \U$9957 ( \10940 , \10936 , \10939 );
and \U$9958 ( \10941 , \10934 , \10939 );
or \U$9959 ( \10942 , \10937 , \10940 , \10941 );
and \U$9960 ( \10943 , \10932 , \10942 );
xor \U$9961 ( \10944 , \10613 , \10615 );
xor \U$9962 ( \10945 , \10944 , \10618 );
and \U$9963 ( \10946 , \10942 , \10945 );
and \U$9964 ( \10947 , \10932 , \10945 );
or \U$9965 ( \10948 , \10943 , \10946 , \10947 );
xor \U$9966 ( \10949 , \10611 , \10621 );
xor \U$9967 ( \10950 , \10949 , \10624 );
and \U$9968 ( \10951 , \10948 , \10950 );
xor \U$9969 ( \10952 , \10629 , \10631 );
xor \U$9970 ( \10953 , \10952 , \10634 );
and \U$9971 ( \10954 , \10950 , \10953 );
and \U$9972 ( \10955 , \10948 , \10953 );
or \U$9973 ( \10956 , \10951 , \10954 , \10955 );
xor \U$9974 ( \10957 , \10627 , \10637 );
xor \U$9975 ( \10958 , \10957 , \10640 );
and \U$9976 ( \10959 , \10956 , \10958 );
xor \U$9977 ( \10960 , \10310 , \10320 );
xor \U$9978 ( \10961 , \10960 , \10323 );
and \U$9979 ( \10962 , \10958 , \10961 );
and \U$9980 ( \10963 , \10956 , \10961 );
or \U$9981 ( \10964 , \10959 , \10962 , \10963 );
and \U$9982 ( \10965 , \10649 , \10964 );
xor \U$9983 ( \10966 , \10649 , \10964 );
xor \U$9984 ( \10967 , \10956 , \10958 );
xor \U$9985 ( \10968 , \10967 , \10961 );
xor \U$9986 ( \10969 , \10777 , \10781 );
xor \U$9987 ( \10970 , \10969 , \10786 );
xor \U$9988 ( \10971 , \10794 , \10798 );
xor \U$9989 ( \10972 , \10971 , \10803 );
and \U$9990 ( \10973 , \10970 , \10972 );
xor \U$9991 ( \10974 , \10724 , \10728 );
xor \U$9992 ( \10975 , \10974 , \10733 );
and \U$9993 ( \10976 , \10972 , \10975 );
and \U$9994 ( \10977 , \10970 , \10975 );
or \U$9995 ( \10978 , \10973 , \10976 , \10977 );
xor \U$9996 ( \10979 , \10708 , \10712 );
xor \U$9997 ( \10980 , \10979 , \10717 );
xor \U$9998 ( \10981 , \10816 , \10820 );
xor \U$9999 ( \10982 , \10981 , \10825 );
and \U$10000 ( \10983 , \10980 , \10982 );
xor \U$10001 ( \10984 , \10741 , \10745 );
xor \U$10002 ( \10985 , \10984 , \10750 );
and \U$10003 ( \10986 , \10982 , \10985 );
and \U$10004 ( \10987 , \10980 , \10985 );
or \U$10005 ( \10988 , \10983 , \10986 , \10987 );
and \U$10006 ( \10989 , \10978 , \10988 );
and \U$10007 ( \10990 , \8795 , \1247 );
and \U$10008 ( \10991 , \8371 , \1245 );
nor \U$10009 ( \10992 , \10990 , \10991 );
xnor \U$10010 ( \10993 , \10992 , \1198 );
and \U$10011 ( \10994 , \9046 , \1146 );
and \U$10012 ( \10995 , \9041 , \1144 );
nor \U$10013 ( \10996 , \10994 , \10995 );
xnor \U$10014 ( \10997 , \10996 , \1105 );
and \U$10015 ( \10998 , \10993 , \10997 );
and \U$10016 ( \10999 , \9649 , \1076 );
and \U$10017 ( \11000 , \9365 , \1074 );
nor \U$10018 ( \11001 , \10999 , \11000 );
xnor \U$10019 ( \11002 , \11001 , \1046 );
and \U$10020 ( \11003 , \10997 , \11002 );
and \U$10021 ( \11004 , \10993 , \11002 );
or \U$10022 ( \11005 , \10998 , \11003 , \11004 );
and \U$10023 ( \11006 , \10226 , \1028 );
and \U$10024 ( \11007 , \10218 , \1026 );
nor \U$10025 ( \11008 , \11006 , \11007 );
xnor \U$10026 ( \11009 , \11008 , \1009 );
and \U$10027 ( \11010 , \10834 , \991 );
and \U$10028 ( \11011 , \10829 , \989 );
nor \U$10029 ( \11012 , \11010 , \11011 );
xnor \U$10030 ( \11013 , \11012 , \996 );
and \U$10031 ( \11014 , \11009 , \11013 );
buf \U$10032 ( \11015 , RIc0db188_127);
and \U$10033 ( \11016 , \11015 , \985 );
and \U$10034 ( \11017 , \11013 , \11016 );
and \U$10035 ( \11018 , \11009 , \11016 );
or \U$10036 ( \11019 , \11014 , \11017 , \11018 );
and \U$10037 ( \11020 , \11005 , \11019 );
xnor \U$10038 ( \11021 , \10833 , \10835 );
and \U$10039 ( \11022 , \11019 , \11021 );
and \U$10040 ( \11023 , \11005 , \11021 );
or \U$10041 ( \11024 , \11020 , \11022 , \11023 );
and \U$10042 ( \11025 , \10988 , \11024 );
and \U$10043 ( \11026 , \10978 , \11024 );
or \U$10044 ( \11027 , \10989 , \11025 , \11026 );
not \U$10045 ( \11028 , \10427 );
and \U$10046 ( \11029 , \998 , \10669 );
and \U$10047 ( \11030 , \984 , \10667 );
nor \U$10048 ( \11031 , \11029 , \11030 );
xnor \U$10049 ( \11032 , \11031 , \10430 );
and \U$10050 ( \11033 , \11028 , \11032 );
and \U$10051 ( \11034 , \1037 , \10101 );
and \U$10052 ( \11035 , \1016 , \10099 );
nor \U$10053 ( \11036 , \11034 , \11035 );
xnor \U$10054 ( \11037 , \11036 , \9791 );
and \U$10055 ( \11038 , \11032 , \11037 );
and \U$10056 ( \11039 , \11028 , \11037 );
or \U$10057 ( \11040 , \11033 , \11038 , \11039 );
and \U$10058 ( \11041 , \1093 , \9564 );
and \U$10059 ( \11042 , \1085 , \9562 );
nor \U$10060 ( \11043 , \11041 , \11042 );
xnor \U$10061 ( \11044 , \11043 , \9193 );
and \U$10062 ( \11045 , \1167 , \9002 );
and \U$10063 ( \11046 , \1162 , \9000 );
nor \U$10064 ( \11047 , \11045 , \11046 );
xnor \U$10065 ( \11048 , \11047 , \8684 );
and \U$10066 ( \11049 , \11044 , \11048 );
and \U$10067 ( \11050 , \1272 , \8435 );
and \U$10068 ( \11051 , \1221 , \8433 );
nor \U$10069 ( \11052 , \11050 , \11051 );
xnor \U$10070 ( \11053 , \11052 , \8186 );
and \U$10071 ( \11054 , \11048 , \11053 );
and \U$10072 ( \11055 , \11044 , \11053 );
or \U$10073 ( \11056 , \11049 , \11054 , \11055 );
and \U$10074 ( \11057 , \11040 , \11056 );
and \U$10075 ( \11058 , \1377 , \7906 );
and \U$10076 ( \11059 , \1349 , \7904 );
nor \U$10077 ( \11060 , \11058 , \11059 );
xnor \U$10078 ( \11061 , \11060 , \7646 );
and \U$10079 ( \11062 , \1531 , \7412 );
and \U$10080 ( \11063 , \1457 , \7410 );
nor \U$10081 ( \11064 , \11062 , \11063 );
xnor \U$10082 ( \11065 , \11064 , \7097 );
and \U$10083 ( \11066 , \11061 , \11065 );
and \U$10084 ( \11067 , \1656 , \6903 );
and \U$10085 ( \11068 , \1593 , \6901 );
nor \U$10086 ( \11069 , \11067 , \11068 );
xnor \U$10087 ( \11070 , \11069 , \6563 );
and \U$10088 ( \11071 , \11065 , \11070 );
and \U$10089 ( \11072 , \11061 , \11070 );
or \U$10090 ( \11073 , \11066 , \11071 , \11072 );
and \U$10091 ( \11074 , \11056 , \11073 );
and \U$10092 ( \11075 , \11040 , \11073 );
or \U$10093 ( \11076 , \11057 , \11074 , \11075 );
and \U$10094 ( \11077 , \5447 , \2222 );
and \U$10095 ( \11078 , \5439 , \2220 );
nor \U$10096 ( \11079 , \11077 , \11078 );
xnor \U$10097 ( \11080 , \11079 , \2109 );
and \U$10098 ( \11081 , \5921 , \2028 );
and \U$10099 ( \11082 , \5916 , \2026 );
nor \U$10100 ( \11083 , \11081 , \11082 );
xnor \U$10101 ( \11084 , \11083 , \1892 );
and \U$10102 ( \11085 , \11080 , \11084 );
and \U$10103 ( \11086 , \6444 , \1828 );
and \U$10104 ( \11087 , \6185 , \1826 );
nor \U$10105 ( \11088 , \11086 , \11087 );
xnor \U$10106 ( \11089 , \11088 , \1750 );
and \U$10107 ( \11090 , \11084 , \11089 );
and \U$10108 ( \11091 , \11080 , \11089 );
or \U$10109 ( \11092 , \11085 , \11090 , \11091 );
and \U$10110 ( \11093 , \4557 , \2968 );
and \U$10111 ( \11094 , \4349 , \2966 );
nor \U$10112 ( \11095 , \11093 , \11094 );
xnor \U$10113 ( \11096 , \11095 , \2831 );
and \U$10114 ( \11097 , \4684 , \2762 );
and \U$10115 ( \11098 , \4679 , \2760 );
nor \U$10116 ( \11099 , \11097 , \11098 );
xnor \U$10117 ( \11100 , \11099 , \2610 );
and \U$10118 ( \11101 , \11096 , \11100 );
and \U$10119 ( \11102 , \5137 , \2494 );
and \U$10120 ( \11103 , \4940 , \2492 );
nor \U$10121 ( \11104 , \11102 , \11103 );
xnor \U$10122 ( \11105 , \11104 , \2338 );
and \U$10123 ( \11106 , \11100 , \11105 );
and \U$10124 ( \11107 , \11096 , \11105 );
or \U$10125 ( \11108 , \11101 , \11106 , \11107 );
and \U$10126 ( \11109 , \11092 , \11108 );
and \U$10127 ( \11110 , \6825 , \1664 );
and \U$10128 ( \11111 , \6816 , \1662 );
nor \U$10129 ( \11112 , \11110 , \11111 );
xnor \U$10130 ( \11113 , \11112 , \1570 );
and \U$10131 ( \11114 , \7370 , \1494 );
and \U$10132 ( \11115 , \7168 , \1492 );
nor \U$10133 ( \11116 , \11114 , \11115 );
xnor \U$10134 ( \11117 , \11116 , \1422 );
and \U$10135 ( \11118 , \11113 , \11117 );
and \U$10136 ( \11119 , \7845 , \1360 );
and \U$10137 ( \11120 , \7673 , \1358 );
nor \U$10138 ( \11121 , \11119 , \11120 );
xnor \U$10139 ( \11122 , \11121 , \1317 );
and \U$10140 ( \11123 , \11117 , \11122 );
and \U$10141 ( \11124 , \11113 , \11122 );
or \U$10142 ( \11125 , \11118 , \11123 , \11124 );
and \U$10143 ( \11126 , \11108 , \11125 );
and \U$10144 ( \11127 , \11092 , \11125 );
or \U$10145 ( \11128 , \11109 , \11126 , \11127 );
and \U$10146 ( \11129 , \11076 , \11128 );
and \U$10147 ( \11130 , \2467 , \5023 );
and \U$10148 ( \11131 , \2459 , \5021 );
nor \U$10149 ( \11132 , \11130 , \11131 );
xnor \U$10150 ( \11133 , \11132 , \4880 );
and \U$10151 ( \11134 , \2715 , \4700 );
and \U$10152 ( \11135 , \2710 , \4698 );
nor \U$10153 ( \11136 , \11134 , \11135 );
xnor \U$10154 ( \11137 , \11136 , \4454 );
and \U$10155 ( \11138 , \11133 , \11137 );
and \U$10156 ( \11139 , \3045 , \4305 );
and \U$10157 ( \11140 , \2901 , \4303 );
nor \U$10158 ( \11141 , \11139 , \11140 );
xnor \U$10159 ( \11142 , \11141 , \4118 );
and \U$10160 ( \11143 , \11137 , \11142 );
and \U$10161 ( \11144 , \11133 , \11142 );
or \U$10162 ( \11145 , \11138 , \11143 , \11144 );
and \U$10163 ( \11146 , \3334 , \3992 );
and \U$10164 ( \11147 , \3309 , \3990 );
nor \U$10165 ( \11148 , \11146 , \11147 );
xnor \U$10166 ( \11149 , \11148 , \3787 );
and \U$10167 ( \11150 , \3675 , \3586 );
and \U$10168 ( \11151 , \3508 , \3584 );
nor \U$10169 ( \11152 , \11150 , \11151 );
xnor \U$10170 ( \11153 , \11152 , \3437 );
and \U$10171 ( \11154 , \11149 , \11153 );
and \U$10172 ( \11155 , \3932 , \3264 );
and \U$10173 ( \11156 , \3813 , \3262 );
nor \U$10174 ( \11157 , \11155 , \11156 );
xnor \U$10175 ( \11158 , \11157 , \3122 );
and \U$10176 ( \11159 , \11153 , \11158 );
and \U$10177 ( \11160 , \11149 , \11158 );
or \U$10178 ( \11161 , \11154 , \11159 , \11160 );
and \U$10179 ( \11162 , \11145 , \11161 );
and \U$10180 ( \11163 , \1942 , \6314 );
and \U$10181 ( \11164 , \1854 , \6312 );
nor \U$10182 ( \11165 , \11163 , \11164 );
xnor \U$10183 ( \11166 , \11165 , \6073 );
and \U$10184 ( \11167 , \2052 , \5848 );
and \U$10185 ( \11168 , \2047 , \5846 );
nor \U$10186 ( \11169 , \11167 , \11168 );
xnor \U$10187 ( \11170 , \11169 , \5660 );
and \U$10188 ( \11171 , \11166 , \11170 );
and \U$10189 ( \11172 , \2283 , \5474 );
and \U$10190 ( \11173 , \2168 , \5472 );
nor \U$10191 ( \11174 , \11172 , \11173 );
xnor \U$10192 ( \11175 , \11174 , \5242 );
and \U$10193 ( \11176 , \11170 , \11175 );
and \U$10194 ( \11177 , \11166 , \11175 );
or \U$10195 ( \11178 , \11171 , \11176 , \11177 );
and \U$10196 ( \11179 , \11161 , \11178 );
and \U$10197 ( \11180 , \11145 , \11178 );
or \U$10198 ( \11181 , \11162 , \11179 , \11180 );
and \U$10199 ( \11182 , \11128 , \11181 );
and \U$10200 ( \11183 , \11076 , \11181 );
or \U$10201 ( \11184 , \11129 , \11182 , \11183 );
and \U$10202 ( \11185 , \11027 , \11184 );
xor \U$10203 ( \11186 , \10761 , \10765 );
xor \U$10204 ( \11187 , \11186 , \10770 );
xor \U$10205 ( \11188 , \10653 , \10657 );
xor \U$10206 ( \11189 , \11188 , \10662 );
and \U$10207 ( \11190 , \11187 , \11189 );
xor \U$10208 ( \11191 , \10689 , \10693 );
xor \U$10209 ( \11192 , \11191 , \10698 );
and \U$10210 ( \11193 , \11189 , \11192 );
and \U$10211 ( \11194 , \11187 , \11192 );
or \U$10212 ( \11195 , \11190 , \11193 , \11194 );
xor \U$10213 ( \11196 , \10870 , \10872 );
xor \U$10214 ( \11197 , \11196 , \10875 );
and \U$10215 ( \11198 , \11195 , \11197 );
xor \U$10216 ( \11199 , \10880 , \10882 );
and \U$10217 ( \11200 , \11197 , \11199 );
and \U$10218 ( \11201 , \11195 , \11199 );
or \U$10219 ( \11202 , \11198 , \11200 , \11201 );
and \U$10220 ( \11203 , \11184 , \11202 );
and \U$10221 ( \11204 , \11027 , \11202 );
or \U$10222 ( \11205 , \11185 , \11203 , \11204 );
xor \U$10223 ( \11206 , \10665 , \10684 );
xor \U$10224 ( \11207 , \11206 , \10701 );
xor \U$10225 ( \11208 , \10720 , \10736 );
xor \U$10226 ( \11209 , \11208 , \10753 );
and \U$10227 ( \11210 , \11207 , \11209 );
xor \U$10228 ( \11211 , \10773 , \10789 );
xor \U$10229 ( \11212 , \11211 , \10806 );
and \U$10230 ( \11213 , \11209 , \11212 );
and \U$10231 ( \11214 , \11207 , \11212 );
or \U$10232 ( \11215 , \11210 , \11213 , \11214 );
xor \U$10233 ( \11216 , \10828 , \10836 );
xor \U$10234 ( \11217 , \11216 , \10841 );
xor \U$10235 ( \11218 , \10845 , \10847 );
xor \U$10236 ( \11219 , \11218 , \10850 );
and \U$10237 ( \11220 , \11217 , \11219 );
xor \U$10238 ( \11221 , \10856 , \10858 );
xor \U$10239 ( \11222 , \11221 , \10861 );
and \U$10240 ( \11223 , \11219 , \11222 );
and \U$10241 ( \11224 , \11217 , \11222 );
or \U$10242 ( \11225 , \11220 , \11223 , \11224 );
and \U$10243 ( \11226 , \11215 , \11225 );
xor \U$10244 ( \11227 , \10894 , \10896 );
xor \U$10245 ( \11228 , \11227 , \10899 );
and \U$10246 ( \11229 , \11225 , \11228 );
and \U$10247 ( \11230 , \11215 , \11228 );
or \U$10248 ( \11231 , \11226 , \11229 , \11230 );
and \U$10249 ( \11232 , \11205 , \11231 );
xor \U$10250 ( \11233 , \10844 , \10853 );
xor \U$10251 ( \11234 , \11233 , \10864 );
xor \U$10252 ( \11235 , \10878 , \10883 );
xor \U$10253 ( \11236 , \11235 , \10886 );
and \U$10254 ( \11237 , \11234 , \11236 );
xor \U$10255 ( \11238 , \10904 , \10906 );
xor \U$10256 ( \11239 , \11238 , \10909 );
and \U$10257 ( \11240 , \11236 , \11239 );
and \U$10258 ( \11241 , \11234 , \11239 );
or \U$10259 ( \11242 , \11237 , \11240 , \11241 );
and \U$10260 ( \11243 , \11231 , \11242 );
and \U$10261 ( \11244 , \11205 , \11242 );
or \U$10262 ( \11245 , \11232 , \11243 , \11244 );
xor \U$10263 ( \11246 , \10392 , \10446 );
xor \U$10264 ( \11247 , \11246 , \10499 );
xor \U$10265 ( \11248 , \10902 , \10912 );
xor \U$10266 ( \11249 , \11248 , \10915 );
and \U$10267 ( \11250 , \11247 , \11249 );
xor \U$10268 ( \11251 , \10921 , \10923 );
xor \U$10269 ( \11252 , \11251 , \10926 );
and \U$10270 ( \11253 , \11249 , \11252 );
and \U$10271 ( \11254 , \11247 , \11252 );
or \U$10272 ( \11255 , \11250 , \11253 , \11254 );
and \U$10273 ( \11256 , \11245 , \11255 );
xor \U$10274 ( \11257 , \10581 , \10591 );
xor \U$10275 ( \11258 , \11257 , \10594 );
and \U$10276 ( \11259 , \11255 , \11258 );
and \U$10277 ( \11260 , \11245 , \11258 );
or \U$10278 ( \11261 , \11256 , \11259 , \11260 );
xor \U$10279 ( \11262 , \10502 , \10549 );
xor \U$10280 ( \11263 , \11262 , \10568 );
xor \U$10281 ( \11264 , \10892 , \10918 );
xor \U$10282 ( \11265 , \11264 , \10929 );
and \U$10283 ( \11266 , \11263 , \11265 );
xor \U$10284 ( \11267 , \10934 , \10936 );
xor \U$10285 ( \11268 , \11267 , \10939 );
and \U$10286 ( \11269 , \11265 , \11268 );
and \U$10287 ( \11270 , \11263 , \11268 );
or \U$10288 ( \11271 , \11266 , \11269 , \11270 );
and \U$10289 ( \11272 , \11261 , \11271 );
xor \U$10290 ( \11273 , \10571 , \10597 );
xor \U$10291 ( \11274 , \11273 , \10608 );
and \U$10292 ( \11275 , \11271 , \11274 );
and \U$10293 ( \11276 , \11261 , \11274 );
or \U$10294 ( \11277 , \11272 , \11275 , \11276 );
xor \U$10295 ( \11278 , \10948 , \10950 );
xor \U$10296 ( \11279 , \11278 , \10953 );
and \U$10297 ( \11280 , \11277 , \11279 );
and \U$10298 ( \11281 , \10968 , \11280 );
xor \U$10299 ( \11282 , \10968 , \11280 );
xor \U$10300 ( \11283 , \11277 , \11279 );
xor \U$10301 ( \11284 , \11080 , \11084 );
xor \U$10302 ( \11285 , \11284 , \11089 );
xor \U$10303 ( \11286 , \11096 , \11100 );
xor \U$10304 ( \11287 , \11286 , \11105 );
and \U$10305 ( \11288 , \11285 , \11287 );
xor \U$10306 ( \11289 , \11149 , \11153 );
xor \U$10307 ( \11290 , \11289 , \11158 );
and \U$10308 ( \11291 , \11287 , \11290 );
and \U$10309 ( \11292 , \11285 , \11290 );
or \U$10310 ( \11293 , \11288 , \11291 , \11292 );
xor \U$10311 ( \11294 , \10993 , \10997 );
xor \U$10312 ( \11295 , \11294 , \11002 );
xor \U$10313 ( \11296 , \11009 , \11013 );
xor \U$10314 ( \11297 , \11296 , \11016 );
and \U$10315 ( \11298 , \11295 , \11297 );
xor \U$10316 ( \11299 , \11113 , \11117 );
xor \U$10317 ( \11300 , \11299 , \11122 );
and \U$10318 ( \11301 , \11297 , \11300 );
and \U$10319 ( \11302 , \11295 , \11300 );
or \U$10320 ( \11303 , \11298 , \11301 , \11302 );
and \U$10321 ( \11304 , \11293 , \11303 );
and \U$10322 ( \11305 , \8371 , \1360 );
and \U$10323 ( \11306 , \7845 , \1358 );
nor \U$10324 ( \11307 , \11305 , \11306 );
xnor \U$10325 ( \11308 , \11307 , \1317 );
and \U$10326 ( \11309 , \9041 , \1247 );
and \U$10327 ( \11310 , \8795 , \1245 );
nor \U$10328 ( \11311 , \11309 , \11310 );
xnor \U$10329 ( \11312 , \11311 , \1198 );
and \U$10330 ( \11313 , \11308 , \11312 );
and \U$10331 ( \11314 , \9365 , \1146 );
and \U$10332 ( \11315 , \9046 , \1144 );
nor \U$10333 ( \11316 , \11314 , \11315 );
xnor \U$10334 ( \11317 , \11316 , \1105 );
and \U$10335 ( \11318 , \11312 , \11317 );
and \U$10336 ( \11319 , \11308 , \11317 );
or \U$10337 ( \11320 , \11313 , \11318 , \11319 );
and \U$10338 ( \11321 , \10218 , \1076 );
and \U$10339 ( \11322 , \9649 , \1074 );
nor \U$10340 ( \11323 , \11321 , \11322 );
xnor \U$10341 ( \11324 , \11323 , \1046 );
and \U$10342 ( \11325 , \10829 , \1028 );
and \U$10343 ( \11326 , \10226 , \1026 );
nor \U$10344 ( \11327 , \11325 , \11326 );
xnor \U$10345 ( \11328 , \11327 , \1009 );
and \U$10346 ( \11329 , \11324 , \11328 );
and \U$10347 ( \11330 , \11015 , \991 );
and \U$10348 ( \11331 , \10834 , \989 );
nor \U$10349 ( \11332 , \11330 , \11331 );
xnor \U$10350 ( \11333 , \11332 , \996 );
and \U$10351 ( \11334 , \11328 , \11333 );
and \U$10352 ( \11335 , \11324 , \11333 );
or \U$10353 ( \11336 , \11329 , \11334 , \11335 );
or \U$10354 ( \11337 , \11320 , \11336 );
and \U$10355 ( \11338 , \11303 , \11337 );
and \U$10356 ( \11339 , \11293 , \11337 );
or \U$10357 ( \11340 , \11304 , \11338 , \11339 );
and \U$10358 ( \11341 , \5439 , \2494 );
and \U$10359 ( \11342 , \5137 , \2492 );
nor \U$10360 ( \11343 , \11341 , \11342 );
xnor \U$10361 ( \11344 , \11343 , \2338 );
and \U$10362 ( \11345 , \5916 , \2222 );
and \U$10363 ( \11346 , \5447 , \2220 );
nor \U$10364 ( \11347 , \11345 , \11346 );
xnor \U$10365 ( \11348 , \11347 , \2109 );
and \U$10366 ( \11349 , \11344 , \11348 );
and \U$10367 ( \11350 , \6185 , \2028 );
and \U$10368 ( \11351 , \5921 , \2026 );
nor \U$10369 ( \11352 , \11350 , \11351 );
xnor \U$10370 ( \11353 , \11352 , \1892 );
and \U$10371 ( \11354 , \11348 , \11353 );
and \U$10372 ( \11355 , \11344 , \11353 );
or \U$10373 ( \11356 , \11349 , \11354 , \11355 );
and \U$10374 ( \11357 , \6816 , \1828 );
and \U$10375 ( \11358 , \6444 , \1826 );
nor \U$10376 ( \11359 , \11357 , \11358 );
xnor \U$10377 ( \11360 , \11359 , \1750 );
and \U$10378 ( \11361 , \7168 , \1664 );
and \U$10379 ( \11362 , \6825 , \1662 );
nor \U$10380 ( \11363 , \11361 , \11362 );
xnor \U$10381 ( \11364 , \11363 , \1570 );
and \U$10382 ( \11365 , \11360 , \11364 );
and \U$10383 ( \11366 , \7673 , \1494 );
and \U$10384 ( \11367 , \7370 , \1492 );
nor \U$10385 ( \11368 , \11366 , \11367 );
xnor \U$10386 ( \11369 , \11368 , \1422 );
and \U$10387 ( \11370 , \11364 , \11369 );
and \U$10388 ( \11371 , \11360 , \11369 );
or \U$10389 ( \11372 , \11365 , \11370 , \11371 );
and \U$10390 ( \11373 , \11356 , \11372 );
and \U$10391 ( \11374 , \4349 , \3264 );
and \U$10392 ( \11375 , \3932 , \3262 );
nor \U$10393 ( \11376 , \11374 , \11375 );
xnor \U$10394 ( \11377 , \11376 , \3122 );
and \U$10395 ( \11378 , \4679 , \2968 );
and \U$10396 ( \11379 , \4557 , \2966 );
nor \U$10397 ( \11380 , \11378 , \11379 );
xnor \U$10398 ( \11381 , \11380 , \2831 );
and \U$10399 ( \11382 , \11377 , \11381 );
and \U$10400 ( \11383 , \4940 , \2762 );
and \U$10401 ( \11384 , \4684 , \2760 );
nor \U$10402 ( \11385 , \11383 , \11384 );
xnor \U$10403 ( \11386 , \11385 , \2610 );
and \U$10404 ( \11387 , \11381 , \11386 );
and \U$10405 ( \11388 , \11377 , \11386 );
or \U$10406 ( \11389 , \11382 , \11387 , \11388 );
and \U$10407 ( \11390 , \11372 , \11389 );
and \U$10408 ( \11391 , \11356 , \11389 );
or \U$10409 ( \11392 , \11373 , \11390 , \11391 );
and \U$10410 ( \11393 , \2459 , \5474 );
and \U$10411 ( \11394 , \2283 , \5472 );
nor \U$10412 ( \11395 , \11393 , \11394 );
xnor \U$10413 ( \11396 , \11395 , \5242 );
and \U$10414 ( \11397 , \2710 , \5023 );
and \U$10415 ( \11398 , \2467 , \5021 );
nor \U$10416 ( \11399 , \11397 , \11398 );
xnor \U$10417 ( \11400 , \11399 , \4880 );
and \U$10418 ( \11401 , \11396 , \11400 );
and \U$10419 ( \11402 , \2901 , \4700 );
and \U$10420 ( \11403 , \2715 , \4698 );
nor \U$10421 ( \11404 , \11402 , \11403 );
xnor \U$10422 ( \11405 , \11404 , \4454 );
and \U$10423 ( \11406 , \11400 , \11405 );
and \U$10424 ( \11407 , \11396 , \11405 );
or \U$10425 ( \11408 , \11401 , \11406 , \11407 );
and \U$10426 ( \11409 , \3309 , \4305 );
and \U$10427 ( \11410 , \3045 , \4303 );
nor \U$10428 ( \11411 , \11409 , \11410 );
xnor \U$10429 ( \11412 , \11411 , \4118 );
and \U$10430 ( \11413 , \3508 , \3992 );
and \U$10431 ( \11414 , \3334 , \3990 );
nor \U$10432 ( \11415 , \11413 , \11414 );
xnor \U$10433 ( \11416 , \11415 , \3787 );
and \U$10434 ( \11417 , \11412 , \11416 );
and \U$10435 ( \11418 , \3813 , \3586 );
and \U$10436 ( \11419 , \3675 , \3584 );
nor \U$10437 ( \11420 , \11418 , \11419 );
xnor \U$10438 ( \11421 , \11420 , \3437 );
and \U$10439 ( \11422 , \11416 , \11421 );
and \U$10440 ( \11423 , \11412 , \11421 );
or \U$10441 ( \11424 , \11417 , \11422 , \11423 );
and \U$10442 ( \11425 , \11408 , \11424 );
and \U$10443 ( \11426 , \1854 , \6903 );
and \U$10444 ( \11427 , \1656 , \6901 );
nor \U$10445 ( \11428 , \11426 , \11427 );
xnor \U$10446 ( \11429 , \11428 , \6563 );
and \U$10447 ( \11430 , \2047 , \6314 );
and \U$10448 ( \11431 , \1942 , \6312 );
nor \U$10449 ( \11432 , \11430 , \11431 );
xnor \U$10450 ( \11433 , \11432 , \6073 );
and \U$10451 ( \11434 , \11429 , \11433 );
and \U$10452 ( \11435 , \2168 , \5848 );
and \U$10453 ( \11436 , \2052 , \5846 );
nor \U$10454 ( \11437 , \11435 , \11436 );
xnor \U$10455 ( \11438 , \11437 , \5660 );
and \U$10456 ( \11439 , \11433 , \11438 );
and \U$10457 ( \11440 , \11429 , \11438 );
or \U$10458 ( \11441 , \11434 , \11439 , \11440 );
and \U$10459 ( \11442 , \11424 , \11441 );
and \U$10460 ( \11443 , \11408 , \11441 );
or \U$10461 ( \11444 , \11425 , \11442 , \11443 );
and \U$10462 ( \11445 , \11392 , \11444 );
and \U$10463 ( \11446 , \1085 , \10101 );
and \U$10464 ( \11447 , \1037 , \10099 );
nor \U$10465 ( \11448 , \11446 , \11447 );
xnor \U$10466 ( \11449 , \11448 , \9791 );
and \U$10467 ( \11450 , \1162 , \9564 );
and \U$10468 ( \11451 , \1093 , \9562 );
nor \U$10469 ( \11452 , \11450 , \11451 );
xnor \U$10470 ( \11453 , \11452 , \9193 );
and \U$10471 ( \11454 , \11449 , \11453 );
and \U$10472 ( \11455 , \1221 , \9002 );
and \U$10473 ( \11456 , \1167 , \9000 );
nor \U$10474 ( \11457 , \11455 , \11456 );
xnor \U$10475 ( \11458 , \11457 , \8684 );
and \U$10476 ( \11459 , \11453 , \11458 );
and \U$10477 ( \11460 , \11449 , \11458 );
or \U$10478 ( \11461 , \11454 , \11459 , \11460 );
and \U$10479 ( \11462 , \1349 , \8435 );
and \U$10480 ( \11463 , \1272 , \8433 );
nor \U$10481 ( \11464 , \11462 , \11463 );
xnor \U$10482 ( \11465 , \11464 , \8186 );
and \U$10483 ( \11466 , \1457 , \7906 );
and \U$10484 ( \11467 , \1377 , \7904 );
nor \U$10485 ( \11468 , \11466 , \11467 );
xnor \U$10486 ( \11469 , \11468 , \7646 );
and \U$10487 ( \11470 , \11465 , \11469 );
and \U$10488 ( \11471 , \1593 , \7412 );
and \U$10489 ( \11472 , \1531 , \7410 );
nor \U$10490 ( \11473 , \11471 , \11472 );
xnor \U$10491 ( \11474 , \11473 , \7097 );
and \U$10492 ( \11475 , \11469 , \11474 );
and \U$10493 ( \11476 , \11465 , \11474 );
or \U$10494 ( \11477 , \11470 , \11475 , \11476 );
and \U$10495 ( \11478 , \11461 , \11477 );
buf \U$10496 ( \11479 , RIc0d9400_64);
xor \U$10497 ( \11480 , \10427 , \11479 );
not \U$10498 ( \11481 , \11479 );
and \U$10499 ( \11482 , \11480 , \11481 );
and \U$10500 ( \11483 , \984 , \11482 );
not \U$10501 ( \11484 , \11483 );
xnor \U$10502 ( \11485 , \11484 , \10427 );
and \U$10503 ( \11486 , \1016 , \10669 );
and \U$10504 ( \11487 , \998 , \10667 );
nor \U$10505 ( \11488 , \11486 , \11487 );
xnor \U$10506 ( \11489 , \11488 , \10430 );
and \U$10507 ( \11490 , \11485 , \11489 );
and \U$10508 ( \11491 , \11477 , \11490 );
and \U$10509 ( \11492 , \11461 , \11490 );
or \U$10510 ( \11493 , \11478 , \11491 , \11492 );
and \U$10511 ( \11494 , \11444 , \11493 );
and \U$10512 ( \11495 , \11392 , \11493 );
or \U$10513 ( \11496 , \11445 , \11494 , \11495 );
and \U$10514 ( \11497 , \11340 , \11496 );
xor \U$10515 ( \11498 , \11133 , \11137 );
xor \U$10516 ( \11499 , \11498 , \11142 );
xor \U$10517 ( \11500 , \11061 , \11065 );
xor \U$10518 ( \11501 , \11500 , \11070 );
and \U$10519 ( \11502 , \11499 , \11501 );
xor \U$10520 ( \11503 , \11166 , \11170 );
xor \U$10521 ( \11504 , \11503 , \11175 );
and \U$10522 ( \11505 , \11501 , \11504 );
and \U$10523 ( \11506 , \11499 , \11504 );
or \U$10524 ( \11507 , \11502 , \11505 , \11506 );
xor \U$10525 ( \11508 , \11028 , \11032 );
xor \U$10526 ( \11509 , \11508 , \11037 );
xor \U$10527 ( \11510 , \11044 , \11048 );
xor \U$10528 ( \11511 , \11510 , \11053 );
and \U$10529 ( \11512 , \11509 , \11511 );
and \U$10530 ( \11513 , \11507 , \11512 );
xor \U$10531 ( \11514 , \10672 , \10676 );
xor \U$10532 ( \11515 , \11514 , \10681 );
and \U$10533 ( \11516 , \11512 , \11515 );
and \U$10534 ( \11517 , \11507 , \11515 );
or \U$10535 ( \11518 , \11513 , \11516 , \11517 );
and \U$10536 ( \11519 , \11496 , \11518 );
and \U$10537 ( \11520 , \11340 , \11518 );
or \U$10538 ( \11521 , \11497 , \11519 , \11520 );
xor \U$10539 ( \11522 , \11187 , \11189 );
xor \U$10540 ( \11523 , \11522 , \11192 );
xor \U$10541 ( \11524 , \10970 , \10972 );
xor \U$10542 ( \11525 , \11524 , \10975 );
and \U$10543 ( \11526 , \11523 , \11525 );
xor \U$10544 ( \11527 , \10980 , \10982 );
xor \U$10545 ( \11528 , \11527 , \10985 );
and \U$10546 ( \11529 , \11525 , \11528 );
and \U$10547 ( \11530 , \11523 , \11528 );
or \U$10548 ( \11531 , \11526 , \11529 , \11530 );
xor \U$10549 ( \11532 , \11092 , \11108 );
xor \U$10550 ( \11533 , \11532 , \11125 );
xor \U$10551 ( \11534 , \11145 , \11161 );
xor \U$10552 ( \11535 , \11534 , \11178 );
and \U$10553 ( \11536 , \11533 , \11535 );
xor \U$10554 ( \11537 , \11005 , \11019 );
xor \U$10555 ( \11538 , \11537 , \11021 );
and \U$10556 ( \11539 , \11535 , \11538 );
and \U$10557 ( \11540 , \11533 , \11538 );
or \U$10558 ( \11541 , \11536 , \11539 , \11540 );
and \U$10559 ( \11542 , \11531 , \11541 );
xor \U$10560 ( \11543 , \11207 , \11209 );
xor \U$10561 ( \11544 , \11543 , \11212 );
and \U$10562 ( \11545 , \11541 , \11544 );
and \U$10563 ( \11546 , \11531 , \11544 );
or \U$10564 ( \11547 , \11542 , \11545 , \11546 );
and \U$10565 ( \11548 , \11521 , \11547 );
xor \U$10566 ( \11549 , \10978 , \10988 );
xor \U$10567 ( \11550 , \11549 , \11024 );
xor \U$10568 ( \11551 , \11217 , \11219 );
xor \U$10569 ( \11552 , \11551 , \11222 );
and \U$10570 ( \11553 , \11550 , \11552 );
xor \U$10571 ( \11554 , \11195 , \11197 );
xor \U$10572 ( \11555 , \11554 , \11199 );
and \U$10573 ( \11556 , \11552 , \11555 );
and \U$10574 ( \11557 , \11550 , \11555 );
or \U$10575 ( \11558 , \11553 , \11556 , \11557 );
and \U$10576 ( \11559 , \11547 , \11558 );
and \U$10577 ( \11560 , \11521 , \11558 );
or \U$10578 ( \11561 , \11548 , \11559 , \11560 );
xor \U$10579 ( \11562 , \10704 , \10756 );
xor \U$10580 ( \11563 , \11562 , \10809 );
xor \U$10581 ( \11564 , \11215 , \11225 );
xor \U$10582 ( \11565 , \11564 , \11228 );
and \U$10583 ( \11566 , \11563 , \11565 );
xor \U$10584 ( \11567 , \11234 , \11236 );
xor \U$10585 ( \11568 , \11567 , \11239 );
and \U$10586 ( \11569 , \11565 , \11568 );
and \U$10587 ( \11570 , \11563 , \11568 );
or \U$10588 ( \11571 , \11566 , \11569 , \11570 );
and \U$10589 ( \11572 , \11561 , \11571 );
xor \U$10590 ( \11573 , \10812 , \10867 );
xor \U$10591 ( \11574 , \11573 , \10889 );
and \U$10592 ( \11575 , \11571 , \11574 );
and \U$10593 ( \11576 , \11561 , \11574 );
or \U$10594 ( \11577 , \11572 , \11575 , \11576 );
xor \U$10595 ( \11578 , \11245 , \11255 );
xor \U$10596 ( \11579 , \11578 , \11258 );
and \U$10597 ( \11580 , \11577 , \11579 );
xor \U$10598 ( \11581 , \11263 , \11265 );
xor \U$10599 ( \11582 , \11581 , \11268 );
and \U$10600 ( \11583 , \11579 , \11582 );
and \U$10601 ( \11584 , \11577 , \11582 );
or \U$10602 ( \11585 , \11580 , \11583 , \11584 );
xor \U$10603 ( \11586 , \11261 , \11271 );
xor \U$10604 ( \11587 , \11586 , \11274 );
and \U$10605 ( \11588 , \11585 , \11587 );
xor \U$10606 ( \11589 , \10932 , \10942 );
xor \U$10607 ( \11590 , \11589 , \10945 );
and \U$10608 ( \11591 , \11587 , \11590 );
and \U$10609 ( \11592 , \11585 , \11590 );
or \U$10610 ( \11593 , \11588 , \11591 , \11592 );
and \U$10611 ( \11594 , \11283 , \11593 );
xor \U$10612 ( \11595 , \11283 , \11593 );
xor \U$10613 ( \11596 , \11585 , \11587 );
xor \U$10614 ( \11597 , \11596 , \11590 );
xor \U$10615 ( \11598 , \11344 , \11348 );
xor \U$10616 ( \11599 , \11598 , \11353 );
xor \U$10617 ( \11600 , \11308 , \11312 );
xor \U$10618 ( \11601 , \11600 , \11317 );
and \U$10619 ( \11602 , \11599 , \11601 );
xor \U$10620 ( \11603 , \11360 , \11364 );
xor \U$10621 ( \11604 , \11603 , \11369 );
and \U$10622 ( \11605 , \11601 , \11604 );
and \U$10623 ( \11606 , \11599 , \11604 );
or \U$10624 ( \11607 , \11602 , \11605 , \11606 );
xor \U$10625 ( \11608 , \11396 , \11400 );
xor \U$10626 ( \11609 , \11608 , \11405 );
xor \U$10627 ( \11610 , \11412 , \11416 );
xor \U$10628 ( \11611 , \11610 , \11421 );
and \U$10629 ( \11612 , \11609 , \11611 );
xor \U$10630 ( \11613 , \11377 , \11381 );
xor \U$10631 ( \11614 , \11613 , \11386 );
and \U$10632 ( \11615 , \11611 , \11614 );
and \U$10633 ( \11616 , \11609 , \11614 );
or \U$10634 ( \11617 , \11612 , \11615 , \11616 );
and \U$10635 ( \11618 , \11607 , \11617 );
and \U$10636 ( \11619 , \9046 , \1247 );
and \U$10637 ( \11620 , \9041 , \1245 );
nor \U$10638 ( \11621 , \11619 , \11620 );
xnor \U$10639 ( \11622 , \11621 , \1198 );
and \U$10640 ( \11623 , \9649 , \1146 );
and \U$10641 ( \11624 , \9365 , \1144 );
nor \U$10642 ( \11625 , \11623 , \11624 );
xnor \U$10643 ( \11626 , \11625 , \1105 );
and \U$10644 ( \11627 , \11622 , \11626 );
and \U$10645 ( \11628 , \10226 , \1076 );
and \U$10646 ( \11629 , \10218 , \1074 );
nor \U$10647 ( \11630 , \11628 , \11629 );
xnor \U$10648 ( \11631 , \11630 , \1046 );
and \U$10649 ( \11632 , \11626 , \11631 );
and \U$10650 ( \11633 , \11622 , \11631 );
or \U$10651 ( \11634 , \11627 , \11632 , \11633 );
buf \U$10652 ( \11635 , RIc0db200_128);
nand \U$10653 ( \11636 , \11635 , \985 );
not \U$10654 ( \11637 , \11636 );
and \U$10655 ( \11638 , \11634 , \11637 );
xor \U$10656 ( \11639 , \11324 , \11328 );
xor \U$10657 ( \11640 , \11639 , \11333 );
and \U$10658 ( \11641 , \11637 , \11640 );
and \U$10659 ( \11642 , \11634 , \11640 );
or \U$10660 ( \11643 , \11638 , \11641 , \11642 );
and \U$10661 ( \11644 , \11617 , \11643 );
and \U$10662 ( \11645 , \11607 , \11643 );
or \U$10663 ( \11646 , \11618 , \11644 , \11645 );
and \U$10664 ( \11647 , \2715 , \5023 );
and \U$10665 ( \11648 , \2710 , \5021 );
nor \U$10666 ( \11649 , \11647 , \11648 );
xnor \U$10667 ( \11650 , \11649 , \4880 );
and \U$10668 ( \11651 , \3045 , \4700 );
and \U$10669 ( \11652 , \2901 , \4698 );
nor \U$10670 ( \11653 , \11651 , \11652 );
xnor \U$10671 ( \11654 , \11653 , \4454 );
and \U$10672 ( \11655 , \11650 , \11654 );
and \U$10673 ( \11656 , \3334 , \4305 );
and \U$10674 ( \11657 , \3309 , \4303 );
nor \U$10675 ( \11658 , \11656 , \11657 );
xnor \U$10676 ( \11659 , \11658 , \4118 );
and \U$10677 ( \11660 , \11654 , \11659 );
and \U$10678 ( \11661 , \11650 , \11659 );
or \U$10679 ( \11662 , \11655 , \11660 , \11661 );
and \U$10680 ( \11663 , \2052 , \6314 );
and \U$10681 ( \11664 , \2047 , \6312 );
nor \U$10682 ( \11665 , \11663 , \11664 );
xnor \U$10683 ( \11666 , \11665 , \6073 );
and \U$10684 ( \11667 , \2283 , \5848 );
and \U$10685 ( \11668 , \2168 , \5846 );
nor \U$10686 ( \11669 , \11667 , \11668 );
xnor \U$10687 ( \11670 , \11669 , \5660 );
and \U$10688 ( \11671 , \11666 , \11670 );
and \U$10689 ( \11672 , \2467 , \5474 );
and \U$10690 ( \11673 , \2459 , \5472 );
nor \U$10691 ( \11674 , \11672 , \11673 );
xnor \U$10692 ( \11675 , \11674 , \5242 );
and \U$10693 ( \11676 , \11670 , \11675 );
and \U$10694 ( \11677 , \11666 , \11675 );
or \U$10695 ( \11678 , \11671 , \11676 , \11677 );
and \U$10696 ( \11679 , \11662 , \11678 );
and \U$10697 ( \11680 , \3675 , \3992 );
and \U$10698 ( \11681 , \3508 , \3990 );
nor \U$10699 ( \11682 , \11680 , \11681 );
xnor \U$10700 ( \11683 , \11682 , \3787 );
and \U$10701 ( \11684 , \3932 , \3586 );
and \U$10702 ( \11685 , \3813 , \3584 );
nor \U$10703 ( \11686 , \11684 , \11685 );
xnor \U$10704 ( \11687 , \11686 , \3437 );
and \U$10705 ( \11688 , \11683 , \11687 );
and \U$10706 ( \11689 , \4557 , \3264 );
and \U$10707 ( \11690 , \4349 , \3262 );
nor \U$10708 ( \11691 , \11689 , \11690 );
xnor \U$10709 ( \11692 , \11691 , \3122 );
and \U$10710 ( \11693 , \11687 , \11692 );
and \U$10711 ( \11694 , \11683 , \11692 );
or \U$10712 ( \11695 , \11688 , \11693 , \11694 );
and \U$10713 ( \11696 , \11678 , \11695 );
and \U$10714 ( \11697 , \11662 , \11695 );
or \U$10715 ( \11698 , \11679 , \11696 , \11697 );
and \U$10716 ( \11699 , \1531 , \7906 );
and \U$10717 ( \11700 , \1457 , \7904 );
nor \U$10718 ( \11701 , \11699 , \11700 );
xnor \U$10719 ( \11702 , \11701 , \7646 );
and \U$10720 ( \11703 , \1656 , \7412 );
and \U$10721 ( \11704 , \1593 , \7410 );
nor \U$10722 ( \11705 , \11703 , \11704 );
xnor \U$10723 ( \11706 , \11705 , \7097 );
and \U$10724 ( \11707 , \11702 , \11706 );
and \U$10725 ( \11708 , \1942 , \6903 );
and \U$10726 ( \11709 , \1854 , \6901 );
nor \U$10727 ( \11710 , \11708 , \11709 );
xnor \U$10728 ( \11711 , \11710 , \6563 );
and \U$10729 ( \11712 , \11706 , \11711 );
and \U$10730 ( \11713 , \11702 , \11711 );
or \U$10731 ( \11714 , \11707 , \11712 , \11713 );
and \U$10732 ( \11715 , \1167 , \9564 );
and \U$10733 ( \11716 , \1162 , \9562 );
nor \U$10734 ( \11717 , \11715 , \11716 );
xnor \U$10735 ( \11718 , \11717 , \9193 );
and \U$10736 ( \11719 , \1272 , \9002 );
and \U$10737 ( \11720 , \1221 , \9000 );
nor \U$10738 ( \11721 , \11719 , \11720 );
xnor \U$10739 ( \11722 , \11721 , \8684 );
and \U$10740 ( \11723 , \11718 , \11722 );
and \U$10741 ( \11724 , \1377 , \8435 );
and \U$10742 ( \11725 , \1349 , \8433 );
nor \U$10743 ( \11726 , \11724 , \11725 );
xnor \U$10744 ( \11727 , \11726 , \8186 );
and \U$10745 ( \11728 , \11722 , \11727 );
and \U$10746 ( \11729 , \11718 , \11727 );
or \U$10747 ( \11730 , \11723 , \11728 , \11729 );
and \U$10748 ( \11731 , \11714 , \11730 );
and \U$10749 ( \11732 , \998 , \11482 );
and \U$10750 ( \11733 , \984 , \11479 );
nor \U$10751 ( \11734 , \11732 , \11733 );
xnor \U$10752 ( \11735 , \11734 , \10427 );
and \U$10753 ( \11736 , \1037 , \10669 );
and \U$10754 ( \11737 , \1016 , \10667 );
nor \U$10755 ( \11738 , \11736 , \11737 );
xnor \U$10756 ( \11739 , \11738 , \10430 );
and \U$10757 ( \11740 , \11735 , \11739 );
and \U$10758 ( \11741 , \1093 , \10101 );
and \U$10759 ( \11742 , \1085 , \10099 );
nor \U$10760 ( \11743 , \11741 , \11742 );
xnor \U$10761 ( \11744 , \11743 , \9791 );
and \U$10762 ( \11745 , \11739 , \11744 );
and \U$10763 ( \11746 , \11735 , \11744 );
or \U$10764 ( \11747 , \11740 , \11745 , \11746 );
and \U$10765 ( \11748 , \11730 , \11747 );
and \U$10766 ( \11749 , \11714 , \11747 );
or \U$10767 ( \11750 , \11731 , \11748 , \11749 );
and \U$10768 ( \11751 , \11698 , \11750 );
and \U$10769 ( \11752 , \5921 , \2222 );
and \U$10770 ( \11753 , \5916 , \2220 );
nor \U$10771 ( \11754 , \11752 , \11753 );
xnor \U$10772 ( \11755 , \11754 , \2109 );
and \U$10773 ( \11756 , \6444 , \2028 );
and \U$10774 ( \11757 , \6185 , \2026 );
nor \U$10775 ( \11758 , \11756 , \11757 );
xnor \U$10776 ( \11759 , \11758 , \1892 );
and \U$10777 ( \11760 , \11755 , \11759 );
and \U$10778 ( \11761 , \6825 , \1828 );
and \U$10779 ( \11762 , \6816 , \1826 );
nor \U$10780 ( \11763 , \11761 , \11762 );
xnor \U$10781 ( \11764 , \11763 , \1750 );
and \U$10782 ( \11765 , \11759 , \11764 );
and \U$10783 ( \11766 , \11755 , \11764 );
or \U$10784 ( \11767 , \11760 , \11765 , \11766 );
and \U$10785 ( \11768 , \4684 , \2968 );
and \U$10786 ( \11769 , \4679 , \2966 );
nor \U$10787 ( \11770 , \11768 , \11769 );
xnor \U$10788 ( \11771 , \11770 , \2831 );
and \U$10789 ( \11772 , \5137 , \2762 );
and \U$10790 ( \11773 , \4940 , \2760 );
nor \U$10791 ( \11774 , \11772 , \11773 );
xnor \U$10792 ( \11775 , \11774 , \2610 );
and \U$10793 ( \11776 , \11771 , \11775 );
and \U$10794 ( \11777 , \5447 , \2494 );
and \U$10795 ( \11778 , \5439 , \2492 );
nor \U$10796 ( \11779 , \11777 , \11778 );
xnor \U$10797 ( \11780 , \11779 , \2338 );
and \U$10798 ( \11781 , \11775 , \11780 );
and \U$10799 ( \11782 , \11771 , \11780 );
or \U$10800 ( \11783 , \11776 , \11781 , \11782 );
and \U$10801 ( \11784 , \11767 , \11783 );
and \U$10802 ( \11785 , \7370 , \1664 );
and \U$10803 ( \11786 , \7168 , \1662 );
nor \U$10804 ( \11787 , \11785 , \11786 );
xnor \U$10805 ( \11788 , \11787 , \1570 );
and \U$10806 ( \11789 , \7845 , \1494 );
and \U$10807 ( \11790 , \7673 , \1492 );
nor \U$10808 ( \11791 , \11789 , \11790 );
xnor \U$10809 ( \11792 , \11791 , \1422 );
and \U$10810 ( \11793 , \11788 , \11792 );
and \U$10811 ( \11794 , \8795 , \1360 );
and \U$10812 ( \11795 , \8371 , \1358 );
nor \U$10813 ( \11796 , \11794 , \11795 );
xnor \U$10814 ( \11797 , \11796 , \1317 );
and \U$10815 ( \11798 , \11792 , \11797 );
and \U$10816 ( \11799 , \11788 , \11797 );
or \U$10817 ( \11800 , \11793 , \11798 , \11799 );
and \U$10818 ( \11801 , \11783 , \11800 );
and \U$10819 ( \11802 , \11767 , \11800 );
or \U$10820 ( \11803 , \11784 , \11801 , \11802 );
and \U$10821 ( \11804 , \11750 , \11803 );
and \U$10822 ( \11805 , \11698 , \11803 );
or \U$10823 ( \11806 , \11751 , \11804 , \11805 );
and \U$10824 ( \11807 , \11646 , \11806 );
xor \U$10825 ( \11808 , \11449 , \11453 );
xor \U$10826 ( \11809 , \11808 , \11458 );
xor \U$10827 ( \11810 , \11465 , \11469 );
xor \U$10828 ( \11811 , \11810 , \11474 );
and \U$10829 ( \11812 , \11809 , \11811 );
xor \U$10830 ( \11813 , \11429 , \11433 );
xor \U$10831 ( \11814 , \11813 , \11438 );
and \U$10832 ( \11815 , \11811 , \11814 );
and \U$10833 ( \11816 , \11809 , \11814 );
or \U$10834 ( \11817 , \11812 , \11815 , \11816 );
xor \U$10835 ( \11818 , \11499 , \11501 );
xor \U$10836 ( \11819 , \11818 , \11504 );
and \U$10837 ( \11820 , \11817 , \11819 );
xor \U$10838 ( \11821 , \11509 , \11511 );
and \U$10839 ( \11822 , \11819 , \11821 );
and \U$10840 ( \11823 , \11817 , \11821 );
or \U$10841 ( \11824 , \11820 , \11822 , \11823 );
and \U$10842 ( \11825 , \11806 , \11824 );
and \U$10843 ( \11826 , \11646 , \11824 );
or \U$10844 ( \11827 , \11807 , \11825 , \11826 );
xor \U$10845 ( \11828 , \11356 , \11372 );
xor \U$10846 ( \11829 , \11828 , \11389 );
xor \U$10847 ( \11830 , \11408 , \11424 );
xor \U$10848 ( \11831 , \11830 , \11441 );
and \U$10849 ( \11832 , \11829 , \11831 );
xor \U$10850 ( \11833 , \11461 , \11477 );
xor \U$10851 ( \11834 , \11833 , \11490 );
and \U$10852 ( \11835 , \11831 , \11834 );
and \U$10853 ( \11836 , \11829 , \11834 );
or \U$10854 ( \11837 , \11832 , \11835 , \11836 );
xor \U$10855 ( \11838 , \11285 , \11287 );
xor \U$10856 ( \11839 , \11838 , \11290 );
xor \U$10857 ( \11840 , \11295 , \11297 );
xor \U$10858 ( \11841 , \11840 , \11300 );
and \U$10859 ( \11842 , \11839 , \11841 );
xnor \U$10860 ( \11843 , \11320 , \11336 );
and \U$10861 ( \11844 , \11841 , \11843 );
and \U$10862 ( \11845 , \11839 , \11843 );
or \U$10863 ( \11846 , \11842 , \11844 , \11845 );
and \U$10864 ( \11847 , \11837 , \11846 );
xor \U$10865 ( \11848 , \11040 , \11056 );
xor \U$10866 ( \11849 , \11848 , \11073 );
and \U$10867 ( \11850 , \11846 , \11849 );
and \U$10868 ( \11851 , \11837 , \11849 );
or \U$10869 ( \11852 , \11847 , \11850 , \11851 );
and \U$10870 ( \11853 , \11827 , \11852 );
xor \U$10871 ( \11854 , \11507 , \11512 );
xor \U$10872 ( \11855 , \11854 , \11515 );
xor \U$10873 ( \11856 , \11523 , \11525 );
xor \U$10874 ( \11857 , \11856 , \11528 );
and \U$10875 ( \11858 , \11855 , \11857 );
xor \U$10876 ( \11859 , \11533 , \11535 );
xor \U$10877 ( \11860 , \11859 , \11538 );
and \U$10878 ( \11861 , \11857 , \11860 );
and \U$10879 ( \11862 , \11855 , \11860 );
or \U$10880 ( \11863 , \11858 , \11861 , \11862 );
and \U$10881 ( \11864 , \11852 , \11863 );
and \U$10882 ( \11865 , \11827 , \11863 );
or \U$10883 ( \11866 , \11853 , \11864 , \11865 );
xor \U$10884 ( \11867 , \11076 , \11128 );
xor \U$10885 ( \11868 , \11867 , \11181 );
xor \U$10886 ( \11869 , \11531 , \11541 );
xor \U$10887 ( \11870 , \11869 , \11544 );
and \U$10888 ( \11871 , \11868 , \11870 );
xor \U$10889 ( \11872 , \11550 , \11552 );
xor \U$10890 ( \11873 , \11872 , \11555 );
and \U$10891 ( \11874 , \11870 , \11873 );
and \U$10892 ( \11875 , \11868 , \11873 );
or \U$10893 ( \11876 , \11871 , \11874 , \11875 );
and \U$10894 ( \11877 , \11866 , \11876 );
xor \U$10895 ( \11878 , \11027 , \11184 );
xor \U$10896 ( \11879 , \11878 , \11202 );
and \U$10897 ( \11880 , \11876 , \11879 );
and \U$10898 ( \11881 , \11866 , \11879 );
or \U$10899 ( \11882 , \11877 , \11880 , \11881 );
xor \U$10900 ( \11883 , \11521 , \11547 );
xor \U$10901 ( \11884 , \11883 , \11558 );
xor \U$10902 ( \11885 , \11563 , \11565 );
xor \U$10903 ( \11886 , \11885 , \11568 );
and \U$10904 ( \11887 , \11884 , \11886 );
and \U$10905 ( \11888 , \11882 , \11887 );
xor \U$10906 ( \11889 , \11247 , \11249 );
xor \U$10907 ( \11890 , \11889 , \11252 );
and \U$10908 ( \11891 , \11887 , \11890 );
and \U$10909 ( \11892 , \11882 , \11890 );
or \U$10910 ( \11893 , \11888 , \11891 , \11892 );
xor \U$10911 ( \11894 , \11205 , \11231 );
xor \U$10912 ( \11895 , \11894 , \11242 );
xor \U$10913 ( \11896 , \11561 , \11571 );
xor \U$10914 ( \11897 , \11896 , \11574 );
and \U$10915 ( \11898 , \11895 , \11897 );
and \U$10916 ( \11899 , \11893 , \11898 );
xor \U$10917 ( \11900 , \11577 , \11579 );
xor \U$10918 ( \11901 , \11900 , \11582 );
and \U$10919 ( \11902 , \11898 , \11901 );
and \U$10920 ( \11903 , \11893 , \11901 );
or \U$10921 ( \11904 , \11899 , \11902 , \11903 );
and \U$10922 ( \11905 , \11597 , \11904 );
xor \U$10923 ( \11906 , \11597 , \11904 );
xor \U$10924 ( \11907 , \11893 , \11898 );
xor \U$10925 ( \11908 , \11907 , \11901 );
and \U$10926 ( \11909 , \10829 , \1076 );
and \U$10927 ( \11910 , \10226 , \1074 );
nor \U$10928 ( \11911 , \11909 , \11910 );
xnor \U$10929 ( \11912 , \11911 , \1046 );
and \U$10930 ( \11913 , \11015 , \1028 );
and \U$10931 ( \11914 , \10834 , \1026 );
nor \U$10932 ( \11915 , \11913 , \11914 );
xnor \U$10933 ( \11916 , \11915 , \1009 );
and \U$10934 ( \11917 , \11912 , \11916 );
nand \U$10935 ( \11918 , \11635 , \989 );
xnor \U$10936 ( \11919 , \11918 , \996 );
and \U$10937 ( \11920 , \11916 , \11919 );
and \U$10938 ( \11921 , \11912 , \11919 );
or \U$10939 ( \11922 , \11917 , \11920 , \11921 );
and \U$10940 ( \11923 , \9041 , \1360 );
and \U$10941 ( \11924 , \8795 , \1358 );
nor \U$10942 ( \11925 , \11923 , \11924 );
xnor \U$10943 ( \11926 , \11925 , \1317 );
and \U$10944 ( \11927 , \9365 , \1247 );
and \U$10945 ( \11928 , \9046 , \1245 );
nor \U$10946 ( \11929 , \11927 , \11928 );
xnor \U$10947 ( \11930 , \11929 , \1198 );
and \U$10948 ( \11931 , \11926 , \11930 );
and \U$10949 ( \11932 , \10218 , \1146 );
and \U$10950 ( \11933 , \9649 , \1144 );
nor \U$10951 ( \11934 , \11932 , \11933 );
xnor \U$10952 ( \11935 , \11934 , \1105 );
and \U$10953 ( \11936 , \11930 , \11935 );
and \U$10954 ( \11937 , \11926 , \11935 );
or \U$10955 ( \11938 , \11931 , \11936 , \11937 );
and \U$10956 ( \11939 , \11922 , \11938 );
and \U$10957 ( \11940 , \10834 , \1028 );
and \U$10958 ( \11941 , \10829 , \1026 );
nor \U$10959 ( \11942 , \11940 , \11941 );
xnor \U$10960 ( \11943 , \11942 , \1009 );
and \U$10961 ( \11944 , \11938 , \11943 );
and \U$10962 ( \11945 , \11922 , \11943 );
or \U$10963 ( \11946 , \11939 , \11944 , \11945 );
and \U$10964 ( \11947 , \11635 , \991 );
and \U$10965 ( \11948 , \11015 , \989 );
nor \U$10966 ( \11949 , \11947 , \11948 );
xnor \U$10967 ( \11950 , \11949 , \996 );
xor \U$10968 ( \11951 , \11788 , \11792 );
xor \U$10969 ( \11952 , \11951 , \11797 );
and \U$10970 ( \11953 , \11950 , \11952 );
xor \U$10971 ( \11954 , \11622 , \11626 );
xor \U$10972 ( \11955 , \11954 , \11631 );
and \U$10973 ( \11956 , \11952 , \11955 );
and \U$10974 ( \11957 , \11950 , \11955 );
or \U$10975 ( \11958 , \11953 , \11956 , \11957 );
and \U$10976 ( \11959 , \11946 , \11958 );
xor \U$10977 ( \11960 , \11755 , \11759 );
xor \U$10978 ( \11961 , \11960 , \11764 );
xor \U$10979 ( \11962 , \11771 , \11775 );
xor \U$10980 ( \11963 , \11962 , \11780 );
and \U$10981 ( \11964 , \11961 , \11963 );
xor \U$10982 ( \11965 , \11683 , \11687 );
xor \U$10983 ( \11966 , \11965 , \11692 );
and \U$10984 ( \11967 , \11963 , \11966 );
and \U$10985 ( \11968 , \11961 , \11966 );
or \U$10986 ( \11969 , \11964 , \11967 , \11968 );
and \U$10987 ( \11970 , \11958 , \11969 );
and \U$10988 ( \11971 , \11946 , \11969 );
or \U$10989 ( \11972 , \11959 , \11970 , \11971 );
and \U$10990 ( \11973 , \5916 , \2494 );
and \U$10991 ( \11974 , \5447 , \2492 );
nor \U$10992 ( \11975 , \11973 , \11974 );
xnor \U$10993 ( \11976 , \11975 , \2338 );
and \U$10994 ( \11977 , \6185 , \2222 );
and \U$10995 ( \11978 , \5921 , \2220 );
nor \U$10996 ( \11979 , \11977 , \11978 );
xnor \U$10997 ( \11980 , \11979 , \2109 );
and \U$10998 ( \11981 , \11976 , \11980 );
and \U$10999 ( \11982 , \6816 , \2028 );
and \U$11000 ( \11983 , \6444 , \2026 );
nor \U$11001 ( \11984 , \11982 , \11983 );
xnor \U$11002 ( \11985 , \11984 , \1892 );
and \U$11003 ( \11986 , \11980 , \11985 );
and \U$11004 ( \11987 , \11976 , \11985 );
or \U$11005 ( \11988 , \11981 , \11986 , \11987 );
and \U$11006 ( \11989 , \4679 , \3264 );
and \U$11007 ( \11990 , \4557 , \3262 );
nor \U$11008 ( \11991 , \11989 , \11990 );
xnor \U$11009 ( \11992 , \11991 , \3122 );
and \U$11010 ( \11993 , \4940 , \2968 );
and \U$11011 ( \11994 , \4684 , \2966 );
nor \U$11012 ( \11995 , \11993 , \11994 );
xnor \U$11013 ( \11996 , \11995 , \2831 );
and \U$11014 ( \11997 , \11992 , \11996 );
and \U$11015 ( \11998 , \5439 , \2762 );
and \U$11016 ( \11999 , \5137 , \2760 );
nor \U$11017 ( \12000 , \11998 , \11999 );
xnor \U$11018 ( \12001 , \12000 , \2610 );
and \U$11019 ( \12002 , \11996 , \12001 );
and \U$11020 ( \12003 , \11992 , \12001 );
or \U$11021 ( \12004 , \11997 , \12002 , \12003 );
and \U$11022 ( \12005 , \11988 , \12004 );
and \U$11023 ( \12006 , \7168 , \1828 );
and \U$11024 ( \12007 , \6825 , \1826 );
nor \U$11025 ( \12008 , \12006 , \12007 );
xnor \U$11026 ( \12009 , \12008 , \1750 );
and \U$11027 ( \12010 , \7673 , \1664 );
and \U$11028 ( \12011 , \7370 , \1662 );
nor \U$11029 ( \12012 , \12010 , \12011 );
xnor \U$11030 ( \12013 , \12012 , \1570 );
and \U$11031 ( \12014 , \12009 , \12013 );
and \U$11032 ( \12015 , \8371 , \1494 );
and \U$11033 ( \12016 , \7845 , \1492 );
nor \U$11034 ( \12017 , \12015 , \12016 );
xnor \U$11035 ( \12018 , \12017 , \1422 );
and \U$11036 ( \12019 , \12013 , \12018 );
and \U$11037 ( \12020 , \12009 , \12018 );
or \U$11038 ( \12021 , \12014 , \12019 , \12020 );
and \U$11039 ( \12022 , \12004 , \12021 );
and \U$11040 ( \12023 , \11988 , \12021 );
or \U$11041 ( \12024 , \12005 , \12022 , \12023 );
and \U$11042 ( \12025 , \1457 , \8435 );
and \U$11043 ( \12026 , \1377 , \8433 );
nor \U$11044 ( \12027 , \12025 , \12026 );
xnor \U$11045 ( \12028 , \12027 , \8186 );
and \U$11046 ( \12029 , \1593 , \7906 );
and \U$11047 ( \12030 , \1531 , \7904 );
nor \U$11048 ( \12031 , \12029 , \12030 );
xnor \U$11049 ( \12032 , \12031 , \7646 );
and \U$11050 ( \12033 , \12028 , \12032 );
and \U$11051 ( \12034 , \1854 , \7412 );
and \U$11052 ( \12035 , \1656 , \7410 );
nor \U$11053 ( \12036 , \12034 , \12035 );
xnor \U$11054 ( \12037 , \12036 , \7097 );
and \U$11055 ( \12038 , \12032 , \12037 );
and \U$11056 ( \12039 , \12028 , \12037 );
or \U$11057 ( \12040 , \12033 , \12038 , \12039 );
and \U$11058 ( \12041 , \1016 , \11482 );
and \U$11059 ( \12042 , \998 , \11479 );
nor \U$11060 ( \12043 , \12041 , \12042 );
xnor \U$11061 ( \12044 , \12043 , \10427 );
and \U$11062 ( \12045 , \1085 , \10669 );
and \U$11063 ( \12046 , \1037 , \10667 );
nor \U$11064 ( \12047 , \12045 , \12046 );
xnor \U$11065 ( \12048 , \12047 , \10430 );
and \U$11066 ( \12049 , \12044 , \12048 );
and \U$11067 ( \12050 , \12048 , \996 );
and \U$11068 ( \12051 , \12044 , \996 );
or \U$11069 ( \12052 , \12049 , \12050 , \12051 );
and \U$11070 ( \12053 , \12040 , \12052 );
and \U$11071 ( \12054 , \1162 , \10101 );
and \U$11072 ( \12055 , \1093 , \10099 );
nor \U$11073 ( \12056 , \12054 , \12055 );
xnor \U$11074 ( \12057 , \12056 , \9791 );
and \U$11075 ( \12058 , \1221 , \9564 );
and \U$11076 ( \12059 , \1167 , \9562 );
nor \U$11077 ( \12060 , \12058 , \12059 );
xnor \U$11078 ( \12061 , \12060 , \9193 );
and \U$11079 ( \12062 , \12057 , \12061 );
and \U$11080 ( \12063 , \1349 , \9002 );
and \U$11081 ( \12064 , \1272 , \9000 );
nor \U$11082 ( \12065 , \12063 , \12064 );
xnor \U$11083 ( \12066 , \12065 , \8684 );
and \U$11084 ( \12067 , \12061 , \12066 );
and \U$11085 ( \12068 , \12057 , \12066 );
or \U$11086 ( \12069 , \12062 , \12067 , \12068 );
and \U$11087 ( \12070 , \12052 , \12069 );
and \U$11088 ( \12071 , \12040 , \12069 );
or \U$11089 ( \12072 , \12053 , \12070 , \12071 );
and \U$11090 ( \12073 , \12024 , \12072 );
and \U$11091 ( \12074 , \2710 , \5474 );
and \U$11092 ( \12075 , \2467 , \5472 );
nor \U$11093 ( \12076 , \12074 , \12075 );
xnor \U$11094 ( \12077 , \12076 , \5242 );
and \U$11095 ( \12078 , \2901 , \5023 );
and \U$11096 ( \12079 , \2715 , \5021 );
nor \U$11097 ( \12080 , \12078 , \12079 );
xnor \U$11098 ( \12081 , \12080 , \4880 );
and \U$11099 ( \12082 , \12077 , \12081 );
and \U$11100 ( \12083 , \3309 , \4700 );
and \U$11101 ( \12084 , \3045 , \4698 );
nor \U$11102 ( \12085 , \12083 , \12084 );
xnor \U$11103 ( \12086 , \12085 , \4454 );
and \U$11104 ( \12087 , \12081 , \12086 );
and \U$11105 ( \12088 , \12077 , \12086 );
or \U$11106 ( \12089 , \12082 , \12087 , \12088 );
and \U$11107 ( \12090 , \2047 , \6903 );
and \U$11108 ( \12091 , \1942 , \6901 );
nor \U$11109 ( \12092 , \12090 , \12091 );
xnor \U$11110 ( \12093 , \12092 , \6563 );
and \U$11111 ( \12094 , \2168 , \6314 );
and \U$11112 ( \12095 , \2052 , \6312 );
nor \U$11113 ( \12096 , \12094 , \12095 );
xnor \U$11114 ( \12097 , \12096 , \6073 );
and \U$11115 ( \12098 , \12093 , \12097 );
and \U$11116 ( \12099 , \2459 , \5848 );
and \U$11117 ( \12100 , \2283 , \5846 );
nor \U$11118 ( \12101 , \12099 , \12100 );
xnor \U$11119 ( \12102 , \12101 , \5660 );
and \U$11120 ( \12103 , \12097 , \12102 );
and \U$11121 ( \12104 , \12093 , \12102 );
or \U$11122 ( \12105 , \12098 , \12103 , \12104 );
and \U$11123 ( \12106 , \12089 , \12105 );
and \U$11124 ( \12107 , \3508 , \4305 );
and \U$11125 ( \12108 , \3334 , \4303 );
nor \U$11126 ( \12109 , \12107 , \12108 );
xnor \U$11127 ( \12110 , \12109 , \4118 );
and \U$11128 ( \12111 , \3813 , \3992 );
and \U$11129 ( \12112 , \3675 , \3990 );
nor \U$11130 ( \12113 , \12111 , \12112 );
xnor \U$11131 ( \12114 , \12113 , \3787 );
and \U$11132 ( \12115 , \12110 , \12114 );
and \U$11133 ( \12116 , \4349 , \3586 );
and \U$11134 ( \12117 , \3932 , \3584 );
nor \U$11135 ( \12118 , \12116 , \12117 );
xnor \U$11136 ( \12119 , \12118 , \3437 );
and \U$11137 ( \12120 , \12114 , \12119 );
and \U$11138 ( \12121 , \12110 , \12119 );
or \U$11139 ( \12122 , \12115 , \12120 , \12121 );
and \U$11140 ( \12123 , \12105 , \12122 );
and \U$11141 ( \12124 , \12089 , \12122 );
or \U$11142 ( \12125 , \12106 , \12123 , \12124 );
and \U$11143 ( \12126 , \12072 , \12125 );
and \U$11144 ( \12127 , \12024 , \12125 );
or \U$11145 ( \12128 , \12073 , \12126 , \12127 );
and \U$11146 ( \12129 , \11972 , \12128 );
xor \U$11147 ( \12130 , \11650 , \11654 );
xor \U$11148 ( \12131 , \12130 , \11659 );
xor \U$11149 ( \12132 , \11666 , \11670 );
xor \U$11150 ( \12133 , \12132 , \11675 );
and \U$11151 ( \12134 , \12131 , \12133 );
xor \U$11152 ( \12135 , \11702 , \11706 );
xor \U$11153 ( \12136 , \12135 , \11711 );
and \U$11154 ( \12137 , \12133 , \12136 );
and \U$11155 ( \12138 , \12131 , \12136 );
or \U$11156 ( \12139 , \12134 , \12137 , \12138 );
xor \U$11157 ( \12140 , \11718 , \11722 );
xor \U$11158 ( \12141 , \12140 , \11727 );
xor \U$11159 ( \12142 , \11735 , \11739 );
xor \U$11160 ( \12143 , \12142 , \11744 );
and \U$11161 ( \12144 , \12141 , \12143 );
and \U$11162 ( \12145 , \12139 , \12144 );
xor \U$11163 ( \12146 , \11485 , \11489 );
and \U$11164 ( \12147 , \12144 , \12146 );
and \U$11165 ( \12148 , \12139 , \12146 );
or \U$11166 ( \12149 , \12145 , \12147 , \12148 );
and \U$11167 ( \12150 , \12128 , \12149 );
and \U$11168 ( \12151 , \11972 , \12149 );
or \U$11169 ( \12152 , \12129 , \12150 , \12151 );
xor \U$11170 ( \12153 , \11662 , \11678 );
xor \U$11171 ( \12154 , \12153 , \11695 );
xor \U$11172 ( \12155 , \11767 , \11783 );
xor \U$11173 ( \12156 , \12155 , \11800 );
and \U$11174 ( \12157 , \12154 , \12156 );
xor \U$11175 ( \12158 , \11634 , \11637 );
xor \U$11176 ( \12159 , \12158 , \11640 );
and \U$11177 ( \12160 , \12156 , \12159 );
and \U$11178 ( \12161 , \12154 , \12159 );
or \U$11179 ( \12162 , \12157 , \12160 , \12161 );
xor \U$11180 ( \12163 , \11809 , \11811 );
xor \U$11181 ( \12164 , \12163 , \11814 );
xor \U$11182 ( \12165 , \11599 , \11601 );
xor \U$11183 ( \12166 , \12165 , \11604 );
and \U$11184 ( \12167 , \12164 , \12166 );
xor \U$11185 ( \12168 , \11609 , \11611 );
xor \U$11186 ( \12169 , \12168 , \11614 );
and \U$11187 ( \12170 , \12166 , \12169 );
and \U$11188 ( \12171 , \12164 , \12169 );
or \U$11189 ( \12172 , \12167 , \12170 , \12171 );
and \U$11190 ( \12173 , \12162 , \12172 );
xor \U$11191 ( \12174 , \11829 , \11831 );
xor \U$11192 ( \12175 , \12174 , \11834 );
and \U$11193 ( \12176 , \12172 , \12175 );
and \U$11194 ( \12177 , \12162 , \12175 );
or \U$11195 ( \12178 , \12173 , \12176 , \12177 );
and \U$11196 ( \12179 , \12152 , \12178 );
xor \U$11197 ( \12180 , \11607 , \11617 );
xor \U$11198 ( \12181 , \12180 , \11643 );
xor \U$11199 ( \12182 , \11839 , \11841 );
xor \U$11200 ( \12183 , \12182 , \11843 );
and \U$11201 ( \12184 , \12181 , \12183 );
xor \U$11202 ( \12185 , \11817 , \11819 );
xor \U$11203 ( \12186 , \12185 , \11821 );
and \U$11204 ( \12187 , \12183 , \12186 );
and \U$11205 ( \12188 , \12181 , \12186 );
or \U$11206 ( \12189 , \12184 , \12187 , \12188 );
and \U$11207 ( \12190 , \12178 , \12189 );
and \U$11208 ( \12191 , \12152 , \12189 );
or \U$11209 ( \12192 , \12179 , \12190 , \12191 );
xor \U$11210 ( \12193 , \11293 , \11303 );
xor \U$11211 ( \12194 , \12193 , \11337 );
xor \U$11212 ( \12195 , \11392 , \11444 );
xor \U$11213 ( \12196 , \12195 , \11493 );
and \U$11214 ( \12197 , \12194 , \12196 );
xor \U$11215 ( \12198 , \11855 , \11857 );
xor \U$11216 ( \12199 , \12198 , \11860 );
and \U$11217 ( \12200 , \12196 , \12199 );
and \U$11218 ( \12201 , \12194 , \12199 );
or \U$11219 ( \12202 , \12197 , \12200 , \12201 );
and \U$11220 ( \12203 , \12192 , \12202 );
xor \U$11221 ( \12204 , \11340 , \11496 );
xor \U$11222 ( \12205 , \12204 , \11518 );
and \U$11223 ( \12206 , \12202 , \12205 );
and \U$11224 ( \12207 , \12192 , \12205 );
or \U$11225 ( \12208 , \12203 , \12206 , \12207 );
xor \U$11226 ( \12209 , \11866 , \11876 );
xor \U$11227 ( \12210 , \12209 , \11879 );
and \U$11228 ( \12211 , \12208 , \12210 );
xor \U$11229 ( \12212 , \11884 , \11886 );
and \U$11230 ( \12213 , \12210 , \12212 );
and \U$11231 ( \12214 , \12208 , \12212 );
or \U$11232 ( \12215 , \12211 , \12213 , \12214 );
xor \U$11233 ( \12216 , \11882 , \11887 );
xor \U$11234 ( \12217 , \12216 , \11890 );
and \U$11235 ( \12218 , \12215 , \12217 );
xor \U$11236 ( \12219 , \11895 , \11897 );
and \U$11237 ( \12220 , \12217 , \12219 );
and \U$11238 ( \12221 , \12215 , \12219 );
or \U$11239 ( \12222 , \12218 , \12220 , \12221 );
and \U$11240 ( \12223 , \11908 , \12222 );
xor \U$11241 ( \12224 , \11908 , \12222 );
xor \U$11242 ( \12225 , \12215 , \12217 );
xor \U$11243 ( \12226 , \12225 , \12219 );
and \U$11244 ( \12227 , \1272 , \9564 );
and \U$11245 ( \12228 , \1221 , \9562 );
nor \U$11246 ( \12229 , \12227 , \12228 );
xnor \U$11247 ( \12230 , \12229 , \9193 );
and \U$11248 ( \12231 , \1377 , \9002 );
and \U$11249 ( \12232 , \1349 , \9000 );
nor \U$11250 ( \12233 , \12231 , \12232 );
xnor \U$11251 ( \12234 , \12233 , \8684 );
and \U$11252 ( \12235 , \12230 , \12234 );
and \U$11253 ( \12236 , \1531 , \8435 );
and \U$11254 ( \12237 , \1457 , \8433 );
nor \U$11255 ( \12238 , \12236 , \12237 );
xnor \U$11256 ( \12239 , \12238 , \8186 );
and \U$11257 ( \12240 , \12234 , \12239 );
and \U$11258 ( \12241 , \12230 , \12239 );
or \U$11259 ( \12242 , \12235 , \12240 , \12241 );
and \U$11260 ( \12243 , \1037 , \11482 );
and \U$11261 ( \12244 , \1016 , \11479 );
nor \U$11262 ( \12245 , \12243 , \12244 );
xnor \U$11263 ( \12246 , \12245 , \10427 );
and \U$11264 ( \12247 , \1093 , \10669 );
and \U$11265 ( \12248 , \1085 , \10667 );
nor \U$11266 ( \12249 , \12247 , \12248 );
xnor \U$11267 ( \12250 , \12249 , \10430 );
and \U$11268 ( \12251 , \12246 , \12250 );
and \U$11269 ( \12252 , \1167 , \10101 );
and \U$11270 ( \12253 , \1162 , \10099 );
nor \U$11271 ( \12254 , \12252 , \12253 );
xnor \U$11272 ( \12255 , \12254 , \9791 );
and \U$11273 ( \12256 , \12250 , \12255 );
and \U$11274 ( \12257 , \12246 , \12255 );
or \U$11275 ( \12258 , \12251 , \12256 , \12257 );
and \U$11276 ( \12259 , \12242 , \12258 );
and \U$11277 ( \12260 , \1656 , \7906 );
and \U$11278 ( \12261 , \1593 , \7904 );
nor \U$11279 ( \12262 , \12260 , \12261 );
xnor \U$11280 ( \12263 , \12262 , \7646 );
and \U$11281 ( \12264 , \1942 , \7412 );
and \U$11282 ( \12265 , \1854 , \7410 );
nor \U$11283 ( \12266 , \12264 , \12265 );
xnor \U$11284 ( \12267 , \12266 , \7097 );
and \U$11285 ( \12268 , \12263 , \12267 );
and \U$11286 ( \12269 , \2052 , \6903 );
and \U$11287 ( \12270 , \2047 , \6901 );
nor \U$11288 ( \12271 , \12269 , \12270 );
xnor \U$11289 ( \12272 , \12271 , \6563 );
and \U$11290 ( \12273 , \12267 , \12272 );
and \U$11291 ( \12274 , \12263 , \12272 );
or \U$11292 ( \12275 , \12268 , \12273 , \12274 );
and \U$11293 ( \12276 , \12258 , \12275 );
and \U$11294 ( \12277 , \12242 , \12275 );
or \U$11295 ( \12278 , \12259 , \12276 , \12277 );
and \U$11296 ( \12279 , \6444 , \2222 );
and \U$11297 ( \12280 , \6185 , \2220 );
nor \U$11298 ( \12281 , \12279 , \12280 );
xnor \U$11299 ( \12282 , \12281 , \2109 );
and \U$11300 ( \12283 , \6825 , \2028 );
and \U$11301 ( \12284 , \6816 , \2026 );
nor \U$11302 ( \12285 , \12283 , \12284 );
xnor \U$11303 ( \12286 , \12285 , \1892 );
and \U$11304 ( \12287 , \12282 , \12286 );
and \U$11305 ( \12288 , \7370 , \1828 );
and \U$11306 ( \12289 , \7168 , \1826 );
nor \U$11307 ( \12290 , \12288 , \12289 );
xnor \U$11308 ( \12291 , \12290 , \1750 );
and \U$11309 ( \12292 , \12286 , \12291 );
and \U$11310 ( \12293 , \12282 , \12291 );
or \U$11311 ( \12294 , \12287 , \12292 , \12293 );
and \U$11312 ( \12295 , \7845 , \1664 );
and \U$11313 ( \12296 , \7673 , \1662 );
nor \U$11314 ( \12297 , \12295 , \12296 );
xnor \U$11315 ( \12298 , \12297 , \1570 );
and \U$11316 ( \12299 , \8795 , \1494 );
and \U$11317 ( \12300 , \8371 , \1492 );
nor \U$11318 ( \12301 , \12299 , \12300 );
xnor \U$11319 ( \12302 , \12301 , \1422 );
and \U$11320 ( \12303 , \12298 , \12302 );
and \U$11321 ( \12304 , \9046 , \1360 );
and \U$11322 ( \12305 , \9041 , \1358 );
nor \U$11323 ( \12306 , \12304 , \12305 );
xnor \U$11324 ( \12307 , \12306 , \1317 );
and \U$11325 ( \12308 , \12302 , \12307 );
and \U$11326 ( \12309 , \12298 , \12307 );
or \U$11327 ( \12310 , \12303 , \12308 , \12309 );
and \U$11328 ( \12311 , \12294 , \12310 );
and \U$11329 ( \12312 , \5137 , \2968 );
and \U$11330 ( \12313 , \4940 , \2966 );
nor \U$11331 ( \12314 , \12312 , \12313 );
xnor \U$11332 ( \12315 , \12314 , \2831 );
and \U$11333 ( \12316 , \5447 , \2762 );
and \U$11334 ( \12317 , \5439 , \2760 );
nor \U$11335 ( \12318 , \12316 , \12317 );
xnor \U$11336 ( \12319 , \12318 , \2610 );
and \U$11337 ( \12320 , \12315 , \12319 );
and \U$11338 ( \12321 , \5921 , \2494 );
and \U$11339 ( \12322 , \5916 , \2492 );
nor \U$11340 ( \12323 , \12321 , \12322 );
xnor \U$11341 ( \12324 , \12323 , \2338 );
and \U$11342 ( \12325 , \12319 , \12324 );
and \U$11343 ( \12326 , \12315 , \12324 );
or \U$11344 ( \12327 , \12320 , \12325 , \12326 );
and \U$11345 ( \12328 , \12310 , \12327 );
and \U$11346 ( \12329 , \12294 , \12327 );
or \U$11347 ( \12330 , \12311 , \12328 , \12329 );
and \U$11348 ( \12331 , \12278 , \12330 );
and \U$11349 ( \12332 , \2283 , \6314 );
and \U$11350 ( \12333 , \2168 , \6312 );
nor \U$11351 ( \12334 , \12332 , \12333 );
xnor \U$11352 ( \12335 , \12334 , \6073 );
and \U$11353 ( \12336 , \2467 , \5848 );
and \U$11354 ( \12337 , \2459 , \5846 );
nor \U$11355 ( \12338 , \12336 , \12337 );
xnor \U$11356 ( \12339 , \12338 , \5660 );
and \U$11357 ( \12340 , \12335 , \12339 );
and \U$11358 ( \12341 , \2715 , \5474 );
and \U$11359 ( \12342 , \2710 , \5472 );
nor \U$11360 ( \12343 , \12341 , \12342 );
xnor \U$11361 ( \12344 , \12343 , \5242 );
and \U$11362 ( \12345 , \12339 , \12344 );
and \U$11363 ( \12346 , \12335 , \12344 );
or \U$11364 ( \12347 , \12340 , \12345 , \12346 );
and \U$11365 ( \12348 , \3932 , \3992 );
and \U$11366 ( \12349 , \3813 , \3990 );
nor \U$11367 ( \12350 , \12348 , \12349 );
xnor \U$11368 ( \12351 , \12350 , \3787 );
and \U$11369 ( \12352 , \4557 , \3586 );
and \U$11370 ( \12353 , \4349 , \3584 );
nor \U$11371 ( \12354 , \12352 , \12353 );
xnor \U$11372 ( \12355 , \12354 , \3437 );
and \U$11373 ( \12356 , \12351 , \12355 );
and \U$11374 ( \12357 , \4684 , \3264 );
and \U$11375 ( \12358 , \4679 , \3262 );
nor \U$11376 ( \12359 , \12357 , \12358 );
xnor \U$11377 ( \12360 , \12359 , \3122 );
and \U$11378 ( \12361 , \12355 , \12360 );
and \U$11379 ( \12362 , \12351 , \12360 );
or \U$11380 ( \12363 , \12356 , \12361 , \12362 );
and \U$11381 ( \12364 , \12347 , \12363 );
and \U$11382 ( \12365 , \3045 , \5023 );
and \U$11383 ( \12366 , \2901 , \5021 );
nor \U$11384 ( \12367 , \12365 , \12366 );
xnor \U$11385 ( \12368 , \12367 , \4880 );
and \U$11386 ( \12369 , \3334 , \4700 );
and \U$11387 ( \12370 , \3309 , \4698 );
nor \U$11388 ( \12371 , \12369 , \12370 );
xnor \U$11389 ( \12372 , \12371 , \4454 );
and \U$11390 ( \12373 , \12368 , \12372 );
and \U$11391 ( \12374 , \3675 , \4305 );
and \U$11392 ( \12375 , \3508 , \4303 );
nor \U$11393 ( \12376 , \12374 , \12375 );
xnor \U$11394 ( \12377 , \12376 , \4118 );
and \U$11395 ( \12378 , \12372 , \12377 );
and \U$11396 ( \12379 , \12368 , \12377 );
or \U$11397 ( \12380 , \12373 , \12378 , \12379 );
and \U$11398 ( \12381 , \12363 , \12380 );
and \U$11399 ( \12382 , \12347 , \12380 );
or \U$11400 ( \12383 , \12364 , \12381 , \12382 );
and \U$11401 ( \12384 , \12330 , \12383 );
and \U$11402 ( \12385 , \12278 , \12383 );
or \U$11403 ( \12386 , \12331 , \12384 , \12385 );
xor \U$11404 ( \12387 , \12077 , \12081 );
xor \U$11405 ( \12388 , \12387 , \12086 );
xor \U$11406 ( \12389 , \12093 , \12097 );
xor \U$11407 ( \12390 , \12389 , \12102 );
and \U$11408 ( \12391 , \12388 , \12390 );
xor \U$11409 ( \12392 , \12110 , \12114 );
xor \U$11410 ( \12393 , \12392 , \12119 );
and \U$11411 ( \12394 , \12390 , \12393 );
and \U$11412 ( \12395 , \12388 , \12393 );
or \U$11413 ( \12396 , \12391 , \12394 , \12395 );
and \U$11414 ( \12397 , \9649 , \1247 );
and \U$11415 ( \12398 , \9365 , \1245 );
nor \U$11416 ( \12399 , \12397 , \12398 );
xnor \U$11417 ( \12400 , \12399 , \1198 );
and \U$11418 ( \12401 , \10226 , \1146 );
and \U$11419 ( \12402 , \10218 , \1144 );
nor \U$11420 ( \12403 , \12401 , \12402 );
xnor \U$11421 ( \12404 , \12403 , \1105 );
and \U$11422 ( \12405 , \12400 , \12404 );
and \U$11423 ( \12406 , \10834 , \1076 );
and \U$11424 ( \12407 , \10829 , \1074 );
nor \U$11425 ( \12408 , \12406 , \12407 );
xnor \U$11426 ( \12409 , \12408 , \1046 );
and \U$11427 ( \12410 , \12404 , \12409 );
and \U$11428 ( \12411 , \12400 , \12409 );
or \U$11429 ( \12412 , \12405 , \12410 , \12411 );
xor \U$11430 ( \12413 , \11912 , \11916 );
xor \U$11431 ( \12414 , \12413 , \11919 );
and \U$11432 ( \12415 , \12412 , \12414 );
xor \U$11433 ( \12416 , \11926 , \11930 );
xor \U$11434 ( \12417 , \12416 , \11935 );
and \U$11435 ( \12418 , \12414 , \12417 );
and \U$11436 ( \12419 , \12412 , \12417 );
or \U$11437 ( \12420 , \12415 , \12418 , \12419 );
and \U$11438 ( \12421 , \12396 , \12420 );
xor \U$11439 ( \12422 , \11976 , \11980 );
xor \U$11440 ( \12423 , \12422 , \11985 );
xor \U$11441 ( \12424 , \11992 , \11996 );
xor \U$11442 ( \12425 , \12424 , \12001 );
and \U$11443 ( \12426 , \12423 , \12425 );
xor \U$11444 ( \12427 , \12009 , \12013 );
xor \U$11445 ( \12428 , \12427 , \12018 );
and \U$11446 ( \12429 , \12425 , \12428 );
and \U$11447 ( \12430 , \12423 , \12428 );
or \U$11448 ( \12431 , \12426 , \12429 , \12430 );
and \U$11449 ( \12432 , \12420 , \12431 );
and \U$11450 ( \12433 , \12396 , \12431 );
or \U$11451 ( \12434 , \12421 , \12432 , \12433 );
and \U$11452 ( \12435 , \12386 , \12434 );
xor \U$11453 ( \12436 , \12028 , \12032 );
xor \U$11454 ( \12437 , \12436 , \12037 );
xor \U$11455 ( \12438 , \12044 , \12048 );
xor \U$11456 ( \12439 , \12438 , \996 );
and \U$11457 ( \12440 , \12437 , \12439 );
xor \U$11458 ( \12441 , \12057 , \12061 );
xor \U$11459 ( \12442 , \12441 , \12066 );
and \U$11460 ( \12443 , \12439 , \12442 );
and \U$11461 ( \12444 , \12437 , \12442 );
or \U$11462 ( \12445 , \12440 , \12443 , \12444 );
xor \U$11463 ( \12446 , \12131 , \12133 );
xor \U$11464 ( \12447 , \12446 , \12136 );
and \U$11465 ( \12448 , \12445 , \12447 );
xor \U$11466 ( \12449 , \12141 , \12143 );
and \U$11467 ( \12450 , \12447 , \12449 );
and \U$11468 ( \12451 , \12445 , \12449 );
or \U$11469 ( \12452 , \12448 , \12450 , \12451 );
and \U$11470 ( \12453 , \12434 , \12452 );
and \U$11471 ( \12454 , \12386 , \12452 );
or \U$11472 ( \12455 , \12435 , \12453 , \12454 );
xor \U$11473 ( \12456 , \11988 , \12004 );
xor \U$11474 ( \12457 , \12456 , \12021 );
xor \U$11475 ( \12458 , \12040 , \12052 );
xor \U$11476 ( \12459 , \12458 , \12069 );
and \U$11477 ( \12460 , \12457 , \12459 );
xor \U$11478 ( \12461 , \12089 , \12105 );
xor \U$11479 ( \12462 , \12461 , \12122 );
and \U$11480 ( \12463 , \12459 , \12462 );
and \U$11481 ( \12464 , \12457 , \12462 );
or \U$11482 ( \12465 , \12460 , \12463 , \12464 );
xor \U$11483 ( \12466 , \11922 , \11938 );
xor \U$11484 ( \12467 , \12466 , \11943 );
xor \U$11485 ( \12468 , \11950 , \11952 );
xor \U$11486 ( \12469 , \12468 , \11955 );
and \U$11487 ( \12470 , \12467 , \12469 );
xor \U$11488 ( \12471 , \11961 , \11963 );
xor \U$11489 ( \12472 , \12471 , \11966 );
and \U$11490 ( \12473 , \12469 , \12472 );
and \U$11491 ( \12474 , \12467 , \12472 );
or \U$11492 ( \12475 , \12470 , \12473 , \12474 );
and \U$11493 ( \12476 , \12465 , \12475 );
xor \U$11494 ( \12477 , \11714 , \11730 );
xor \U$11495 ( \12478 , \12477 , \11747 );
and \U$11496 ( \12479 , \12475 , \12478 );
and \U$11497 ( \12480 , \12465 , \12478 );
or \U$11498 ( \12481 , \12476 , \12479 , \12480 );
and \U$11499 ( \12482 , \12455 , \12481 );
xor \U$11500 ( \12483 , \12154 , \12156 );
xor \U$11501 ( \12484 , \12483 , \12159 );
xor \U$11502 ( \12485 , \12164 , \12166 );
xor \U$11503 ( \12486 , \12485 , \12169 );
and \U$11504 ( \12487 , \12484 , \12486 );
xor \U$11505 ( \12488 , \12139 , \12144 );
xor \U$11506 ( \12489 , \12488 , \12146 );
and \U$11507 ( \12490 , \12486 , \12489 );
and \U$11508 ( \12491 , \12484 , \12489 );
or \U$11509 ( \12492 , \12487 , \12490 , \12491 );
and \U$11510 ( \12493 , \12481 , \12492 );
and \U$11511 ( \12494 , \12455 , \12492 );
or \U$11512 ( \12495 , \12482 , \12493 , \12494 );
xor \U$11513 ( \12496 , \11698 , \11750 );
xor \U$11514 ( \12497 , \12496 , \11803 );
xor \U$11515 ( \12498 , \12162 , \12172 );
xor \U$11516 ( \12499 , \12498 , \12175 );
and \U$11517 ( \12500 , \12497 , \12499 );
xor \U$11518 ( \12501 , \12181 , \12183 );
xor \U$11519 ( \12502 , \12501 , \12186 );
and \U$11520 ( \12503 , \12499 , \12502 );
and \U$11521 ( \12504 , \12497 , \12502 );
or \U$11522 ( \12505 , \12500 , \12503 , \12504 );
and \U$11523 ( \12506 , \12495 , \12505 );
xor \U$11524 ( \12507 , \11837 , \11846 );
xor \U$11525 ( \12508 , \12507 , \11849 );
and \U$11526 ( \12509 , \12505 , \12508 );
and \U$11527 ( \12510 , \12495 , \12508 );
or \U$11528 ( \12511 , \12506 , \12509 , \12510 );
xor \U$11529 ( \12512 , \11646 , \11806 );
xor \U$11530 ( \12513 , \12512 , \11824 );
xor \U$11531 ( \12514 , \12152 , \12178 );
xor \U$11532 ( \12515 , \12514 , \12189 );
and \U$11533 ( \12516 , \12513 , \12515 );
xor \U$11534 ( \12517 , \12194 , \12196 );
xor \U$11535 ( \12518 , \12517 , \12199 );
and \U$11536 ( \12519 , \12515 , \12518 );
and \U$11537 ( \12520 , \12513 , \12518 );
or \U$11538 ( \12521 , \12516 , \12519 , \12520 );
and \U$11539 ( \12522 , \12511 , \12521 );
xor \U$11540 ( \12523 , \11868 , \11870 );
xor \U$11541 ( \12524 , \12523 , \11873 );
and \U$11542 ( \12525 , \12521 , \12524 );
and \U$11543 ( \12526 , \12511 , \12524 );
or \U$11544 ( \12527 , \12522 , \12525 , \12526 );
xor \U$11545 ( \12528 , \11827 , \11852 );
xor \U$11546 ( \12529 , \12528 , \11863 );
xor \U$11547 ( \12530 , \12192 , \12202 );
xor \U$11548 ( \12531 , \12530 , \12205 );
and \U$11549 ( \12532 , \12529 , \12531 );
and \U$11550 ( \12533 , \12527 , \12532 );
xor \U$11551 ( \12534 , \12208 , \12210 );
xor \U$11552 ( \12535 , \12534 , \12212 );
and \U$11553 ( \12536 , \12532 , \12535 );
and \U$11554 ( \12537 , \12527 , \12535 );
or \U$11555 ( \12538 , \12533 , \12536 , \12537 );
and \U$11556 ( \12539 , \12226 , \12538 );
xor \U$11557 ( \12540 , \12226 , \12538 );
xor \U$11558 ( \12541 , \12527 , \12532 );
xor \U$11559 ( \12542 , \12541 , \12535 );
and \U$11560 ( \12543 , \7673 , \1828 );
and \U$11561 ( \12544 , \7370 , \1826 );
nor \U$11562 ( \12545 , \12543 , \12544 );
xnor \U$11563 ( \12546 , \12545 , \1750 );
and \U$11564 ( \12547 , \8371 , \1664 );
and \U$11565 ( \12548 , \7845 , \1662 );
nor \U$11566 ( \12549 , \12547 , \12548 );
xnor \U$11567 ( \12550 , \12549 , \1570 );
and \U$11568 ( \12551 , \12546 , \12550 );
and \U$11569 ( \12552 , \9041 , \1494 );
and \U$11570 ( \12553 , \8795 , \1492 );
nor \U$11571 ( \12554 , \12552 , \12553 );
xnor \U$11572 ( \12555 , \12554 , \1422 );
and \U$11573 ( \12556 , \12550 , \12555 );
and \U$11574 ( \12557 , \12546 , \12555 );
or \U$11575 ( \12558 , \12551 , \12556 , \12557 );
and \U$11576 ( \12559 , \4940 , \3264 );
and \U$11577 ( \12560 , \4684 , \3262 );
nor \U$11578 ( \12561 , \12559 , \12560 );
xnor \U$11579 ( \12562 , \12561 , \3122 );
and \U$11580 ( \12563 , \5439 , \2968 );
and \U$11581 ( \12564 , \5137 , \2966 );
nor \U$11582 ( \12565 , \12563 , \12564 );
xnor \U$11583 ( \12566 , \12565 , \2831 );
and \U$11584 ( \12567 , \12562 , \12566 );
and \U$11585 ( \12568 , \5916 , \2762 );
and \U$11586 ( \12569 , \5447 , \2760 );
nor \U$11587 ( \12570 , \12568 , \12569 );
xnor \U$11588 ( \12571 , \12570 , \2610 );
and \U$11589 ( \12572 , \12566 , \12571 );
and \U$11590 ( \12573 , \12562 , \12571 );
or \U$11591 ( \12574 , \12567 , \12572 , \12573 );
and \U$11592 ( \12575 , \12558 , \12574 );
and \U$11593 ( \12576 , \6185 , \2494 );
and \U$11594 ( \12577 , \5921 , \2492 );
nor \U$11595 ( \12578 , \12576 , \12577 );
xnor \U$11596 ( \12579 , \12578 , \2338 );
and \U$11597 ( \12580 , \6816 , \2222 );
and \U$11598 ( \12581 , \6444 , \2220 );
nor \U$11599 ( \12582 , \12580 , \12581 );
xnor \U$11600 ( \12583 , \12582 , \2109 );
and \U$11601 ( \12584 , \12579 , \12583 );
and \U$11602 ( \12585 , \7168 , \2028 );
and \U$11603 ( \12586 , \6825 , \2026 );
nor \U$11604 ( \12587 , \12585 , \12586 );
xnor \U$11605 ( \12588 , \12587 , \1892 );
and \U$11606 ( \12589 , \12583 , \12588 );
and \U$11607 ( \12590 , \12579 , \12588 );
or \U$11608 ( \12591 , \12584 , \12589 , \12590 );
and \U$11609 ( \12592 , \12574 , \12591 );
and \U$11610 ( \12593 , \12558 , \12591 );
or \U$11611 ( \12594 , \12575 , \12592 , \12593 );
and \U$11612 ( \12595 , \1593 , \8435 );
and \U$11613 ( \12596 , \1531 , \8433 );
nor \U$11614 ( \12597 , \12595 , \12596 );
xnor \U$11615 ( \12598 , \12597 , \8186 );
and \U$11616 ( \12599 , \1854 , \7906 );
and \U$11617 ( \12600 , \1656 , \7904 );
nor \U$11618 ( \12601 , \12599 , \12600 );
xnor \U$11619 ( \12602 , \12601 , \7646 );
and \U$11620 ( \12603 , \12598 , \12602 );
and \U$11621 ( \12604 , \2047 , \7412 );
and \U$11622 ( \12605 , \1942 , \7410 );
nor \U$11623 ( \12606 , \12604 , \12605 );
xnor \U$11624 ( \12607 , \12606 , \7097 );
and \U$11625 ( \12608 , \12602 , \12607 );
and \U$11626 ( \12609 , \12598 , \12607 );
or \U$11627 ( \12610 , \12603 , \12608 , \12609 );
and \U$11628 ( \12611 , \1221 , \10101 );
and \U$11629 ( \12612 , \1167 , \10099 );
nor \U$11630 ( \12613 , \12611 , \12612 );
xnor \U$11631 ( \12614 , \12613 , \9791 );
and \U$11632 ( \12615 , \1349 , \9564 );
and \U$11633 ( \12616 , \1272 , \9562 );
nor \U$11634 ( \12617 , \12615 , \12616 );
xnor \U$11635 ( \12618 , \12617 , \9193 );
and \U$11636 ( \12619 , \12614 , \12618 );
and \U$11637 ( \12620 , \1457 , \9002 );
and \U$11638 ( \12621 , \1377 , \9000 );
nor \U$11639 ( \12622 , \12620 , \12621 );
xnor \U$11640 ( \12623 , \12622 , \8684 );
and \U$11641 ( \12624 , \12618 , \12623 );
and \U$11642 ( \12625 , \12614 , \12623 );
or \U$11643 ( \12626 , \12619 , \12624 , \12625 );
and \U$11644 ( \12627 , \12610 , \12626 );
and \U$11645 ( \12628 , \1085 , \11482 );
and \U$11646 ( \12629 , \1037 , \11479 );
nor \U$11647 ( \12630 , \12628 , \12629 );
xnor \U$11648 ( \12631 , \12630 , \10427 );
and \U$11649 ( \12632 , \1162 , \10669 );
and \U$11650 ( \12633 , \1093 , \10667 );
nor \U$11651 ( \12634 , \12632 , \12633 );
xnor \U$11652 ( \12635 , \12634 , \10430 );
and \U$11653 ( \12636 , \12631 , \12635 );
and \U$11654 ( \12637 , \12635 , \1009 );
and \U$11655 ( \12638 , \12631 , \1009 );
or \U$11656 ( \12639 , \12636 , \12637 , \12638 );
and \U$11657 ( \12640 , \12626 , \12639 );
and \U$11658 ( \12641 , \12610 , \12639 );
or \U$11659 ( \12642 , \12627 , \12640 , \12641 );
and \U$11660 ( \12643 , \12594 , \12642 );
and \U$11661 ( \12644 , \2168 , \6903 );
and \U$11662 ( \12645 , \2052 , \6901 );
nor \U$11663 ( \12646 , \12644 , \12645 );
xnor \U$11664 ( \12647 , \12646 , \6563 );
and \U$11665 ( \12648 , \2459 , \6314 );
and \U$11666 ( \12649 , \2283 , \6312 );
nor \U$11667 ( \12650 , \12648 , \12649 );
xnor \U$11668 ( \12651 , \12650 , \6073 );
and \U$11669 ( \12652 , \12647 , \12651 );
and \U$11670 ( \12653 , \2710 , \5848 );
and \U$11671 ( \12654 , \2467 , \5846 );
nor \U$11672 ( \12655 , \12653 , \12654 );
xnor \U$11673 ( \12656 , \12655 , \5660 );
and \U$11674 ( \12657 , \12651 , \12656 );
and \U$11675 ( \12658 , \12647 , \12656 );
or \U$11676 ( \12659 , \12652 , \12657 , \12658 );
and \U$11677 ( \12660 , \2901 , \5474 );
and \U$11678 ( \12661 , \2715 , \5472 );
nor \U$11679 ( \12662 , \12660 , \12661 );
xnor \U$11680 ( \12663 , \12662 , \5242 );
and \U$11681 ( \12664 , \3309 , \5023 );
and \U$11682 ( \12665 , \3045 , \5021 );
nor \U$11683 ( \12666 , \12664 , \12665 );
xnor \U$11684 ( \12667 , \12666 , \4880 );
and \U$11685 ( \12668 , \12663 , \12667 );
and \U$11686 ( \12669 , \3508 , \4700 );
and \U$11687 ( \12670 , \3334 , \4698 );
nor \U$11688 ( \12671 , \12669 , \12670 );
xnor \U$11689 ( \12672 , \12671 , \4454 );
and \U$11690 ( \12673 , \12667 , \12672 );
and \U$11691 ( \12674 , \12663 , \12672 );
or \U$11692 ( \12675 , \12668 , \12673 , \12674 );
and \U$11693 ( \12676 , \12659 , \12675 );
and \U$11694 ( \12677 , \3813 , \4305 );
and \U$11695 ( \12678 , \3675 , \4303 );
nor \U$11696 ( \12679 , \12677 , \12678 );
xnor \U$11697 ( \12680 , \12679 , \4118 );
and \U$11698 ( \12681 , \4349 , \3992 );
and \U$11699 ( \12682 , \3932 , \3990 );
nor \U$11700 ( \12683 , \12681 , \12682 );
xnor \U$11701 ( \12684 , \12683 , \3787 );
and \U$11702 ( \12685 , \12680 , \12684 );
and \U$11703 ( \12686 , \4679 , \3586 );
and \U$11704 ( \12687 , \4557 , \3584 );
nor \U$11705 ( \12688 , \12686 , \12687 );
xnor \U$11706 ( \12689 , \12688 , \3437 );
and \U$11707 ( \12690 , \12684 , \12689 );
and \U$11708 ( \12691 , \12680 , \12689 );
or \U$11709 ( \12692 , \12685 , \12690 , \12691 );
and \U$11710 ( \12693 , \12675 , \12692 );
and \U$11711 ( \12694 , \12659 , \12692 );
or \U$11712 ( \12695 , \12676 , \12693 , \12694 );
and \U$11713 ( \12696 , \12642 , \12695 );
and \U$11714 ( \12697 , \12594 , \12695 );
or \U$11715 ( \12698 , \12643 , \12696 , \12697 );
and \U$11716 ( \12699 , \9365 , \1360 );
and \U$11717 ( \12700 , \9046 , \1358 );
nor \U$11718 ( \12701 , \12699 , \12700 );
xnor \U$11719 ( \12702 , \12701 , \1317 );
and \U$11720 ( \12703 , \10218 , \1247 );
and \U$11721 ( \12704 , \9649 , \1245 );
nor \U$11722 ( \12705 , \12703 , \12704 );
xnor \U$11723 ( \12706 , \12705 , \1198 );
and \U$11724 ( \12707 , \12702 , \12706 );
and \U$11725 ( \12708 , \10829 , \1146 );
and \U$11726 ( \12709 , \10226 , \1144 );
nor \U$11727 ( \12710 , \12708 , \12709 );
xnor \U$11728 ( \12711 , \12710 , \1105 );
and \U$11729 ( \12712 , \12706 , \12711 );
and \U$11730 ( \12713 , \12702 , \12711 );
or \U$11731 ( \12714 , \12707 , \12712 , \12713 );
and \U$11732 ( \12715 , \11015 , \1076 );
and \U$11733 ( \12716 , \10834 , \1074 );
nor \U$11734 ( \12717 , \12715 , \12716 );
xnor \U$11735 ( \12718 , \12717 , \1046 );
nand \U$11736 ( \12719 , \11635 , \1026 );
xnor \U$11737 ( \12720 , \12719 , \1009 );
and \U$11738 ( \12721 , \12718 , \12720 );
and \U$11739 ( \12722 , \12714 , \12721 );
and \U$11740 ( \12723 , \11635 , \1028 );
and \U$11741 ( \12724 , \11015 , \1026 );
nor \U$11742 ( \12725 , \12723 , \12724 );
xnor \U$11743 ( \12726 , \12725 , \1009 );
and \U$11744 ( \12727 , \12721 , \12726 );
and \U$11745 ( \12728 , \12714 , \12726 );
or \U$11746 ( \12729 , \12722 , \12727 , \12728 );
xor \U$11747 ( \12730 , \12315 , \12319 );
xor \U$11748 ( \12731 , \12730 , \12324 );
xor \U$11749 ( \12732 , \12351 , \12355 );
xor \U$11750 ( \12733 , \12732 , \12360 );
and \U$11751 ( \12734 , \12731 , \12733 );
xor \U$11752 ( \12735 , \12368 , \12372 );
xor \U$11753 ( \12736 , \12735 , \12377 );
and \U$11754 ( \12737 , \12733 , \12736 );
and \U$11755 ( \12738 , \12731 , \12736 );
or \U$11756 ( \12739 , \12734 , \12737 , \12738 );
and \U$11757 ( \12740 , \12729 , \12739 );
xor \U$11758 ( \12741 , \12282 , \12286 );
xor \U$11759 ( \12742 , \12741 , \12291 );
xor \U$11760 ( \12743 , \12298 , \12302 );
xor \U$11761 ( \12744 , \12743 , \12307 );
and \U$11762 ( \12745 , \12742 , \12744 );
xor \U$11763 ( \12746 , \12400 , \12404 );
xor \U$11764 ( \12747 , \12746 , \12409 );
and \U$11765 ( \12748 , \12744 , \12747 );
and \U$11766 ( \12749 , \12742 , \12747 );
or \U$11767 ( \12750 , \12745 , \12748 , \12749 );
and \U$11768 ( \12751 , \12739 , \12750 );
and \U$11769 ( \12752 , \12729 , \12750 );
or \U$11770 ( \12753 , \12740 , \12751 , \12752 );
and \U$11771 ( \12754 , \12698 , \12753 );
xor \U$11772 ( \12755 , \12230 , \12234 );
xor \U$11773 ( \12756 , \12755 , \12239 );
xor \U$11774 ( \12757 , \12335 , \12339 );
xor \U$11775 ( \12758 , \12757 , \12344 );
and \U$11776 ( \12759 , \12756 , \12758 );
xor \U$11777 ( \12760 , \12263 , \12267 );
xor \U$11778 ( \12761 , \12760 , \12272 );
and \U$11779 ( \12762 , \12758 , \12761 );
and \U$11780 ( \12763 , \12756 , \12761 );
or \U$11781 ( \12764 , \12759 , \12762 , \12763 );
xor \U$11782 ( \12765 , \12437 , \12439 );
xor \U$11783 ( \12766 , \12765 , \12442 );
and \U$11784 ( \12767 , \12764 , \12766 );
xor \U$11785 ( \12768 , \12388 , \12390 );
xor \U$11786 ( \12769 , \12768 , \12393 );
and \U$11787 ( \12770 , \12766 , \12769 );
and \U$11788 ( \12771 , \12764 , \12769 );
or \U$11789 ( \12772 , \12767 , \12770 , \12771 );
and \U$11790 ( \12773 , \12753 , \12772 );
and \U$11791 ( \12774 , \12698 , \12772 );
or \U$11792 ( \12775 , \12754 , \12773 , \12774 );
xor \U$11793 ( \12776 , \12294 , \12310 );
xor \U$11794 ( \12777 , \12776 , \12327 );
xor \U$11795 ( \12778 , \12412 , \12414 );
xor \U$11796 ( \12779 , \12778 , \12417 );
and \U$11797 ( \12780 , \12777 , \12779 );
xor \U$11798 ( \12781 , \12423 , \12425 );
xor \U$11799 ( \12782 , \12781 , \12428 );
and \U$11800 ( \12783 , \12779 , \12782 );
and \U$11801 ( \12784 , \12777 , \12782 );
or \U$11802 ( \12785 , \12780 , \12783 , \12784 );
xor \U$11803 ( \12786 , \12457 , \12459 );
xor \U$11804 ( \12787 , \12786 , \12462 );
and \U$11805 ( \12788 , \12785 , \12787 );
xor \U$11806 ( \12789 , \12467 , \12469 );
xor \U$11807 ( \12790 , \12789 , \12472 );
and \U$11808 ( \12791 , \12787 , \12790 );
and \U$11809 ( \12792 , \12785 , \12790 );
or \U$11810 ( \12793 , \12788 , \12791 , \12792 );
and \U$11811 ( \12794 , \12775 , \12793 );
xor \U$11812 ( \12795 , \12278 , \12330 );
xor \U$11813 ( \12796 , \12795 , \12383 );
xor \U$11814 ( \12797 , \12396 , \12420 );
xor \U$11815 ( \12798 , \12797 , \12431 );
and \U$11816 ( \12799 , \12796 , \12798 );
xor \U$11817 ( \12800 , \12445 , \12447 );
xor \U$11818 ( \12801 , \12800 , \12449 );
and \U$11819 ( \12802 , \12798 , \12801 );
and \U$11820 ( \12803 , \12796 , \12801 );
or \U$11821 ( \12804 , \12799 , \12802 , \12803 );
and \U$11822 ( \12805 , \12793 , \12804 );
and \U$11823 ( \12806 , \12775 , \12804 );
or \U$11824 ( \12807 , \12794 , \12805 , \12806 );
xor \U$11825 ( \12808 , \11946 , \11958 );
xor \U$11826 ( \12809 , \12808 , \11969 );
xor \U$11827 ( \12810 , \12024 , \12072 );
xor \U$11828 ( \12811 , \12810 , \12125 );
and \U$11829 ( \12812 , \12809 , \12811 );
xor \U$11830 ( \12813 , \12484 , \12486 );
xor \U$11831 ( \12814 , \12813 , \12489 );
and \U$11832 ( \12815 , \12811 , \12814 );
and \U$11833 ( \12816 , \12809 , \12814 );
or \U$11834 ( \12817 , \12812 , \12815 , \12816 );
and \U$11835 ( \12818 , \12807 , \12817 );
xor \U$11836 ( \12819 , \11972 , \12128 );
xor \U$11837 ( \12820 , \12819 , \12149 );
and \U$11838 ( \12821 , \12817 , \12820 );
and \U$11839 ( \12822 , \12807 , \12820 );
or \U$11840 ( \12823 , \12818 , \12821 , \12822 );
xor \U$11841 ( \12824 , \12495 , \12505 );
xor \U$11842 ( \12825 , \12824 , \12508 );
and \U$11843 ( \12826 , \12823 , \12825 );
xor \U$11844 ( \12827 , \12513 , \12515 );
xor \U$11845 ( \12828 , \12827 , \12518 );
and \U$11846 ( \12829 , \12825 , \12828 );
and \U$11847 ( \12830 , \12823 , \12828 );
or \U$11848 ( \12831 , \12826 , \12829 , \12830 );
xor \U$11849 ( \12832 , \12511 , \12521 );
xor \U$11850 ( \12833 , \12832 , \12524 );
and \U$11851 ( \12834 , \12831 , \12833 );
xor \U$11852 ( \12835 , \12529 , \12531 );
and \U$11853 ( \12836 , \12833 , \12835 );
and \U$11854 ( \12837 , \12831 , \12835 );
or \U$11855 ( \12838 , \12834 , \12836 , \12837 );
and \U$11856 ( \12839 , \12542 , \12838 );
xor \U$11857 ( \12840 , \12542 , \12838 );
xor \U$11858 ( \12841 , \12831 , \12833 );
xor \U$11859 ( \12842 , \12841 , \12835 );
xor \U$11860 ( \12843 , \12546 , \12550 );
xor \U$11861 ( \12844 , \12843 , \12555 );
xor \U$11862 ( \12845 , \12562 , \12566 );
xor \U$11863 ( \12846 , \12845 , \12571 );
and \U$11864 ( \12847 , \12844 , \12846 );
xor \U$11865 ( \12848 , \12579 , \12583 );
xor \U$11866 ( \12849 , \12848 , \12588 );
and \U$11867 ( \12850 , \12846 , \12849 );
and \U$11868 ( \12851 , \12844 , \12849 );
or \U$11869 ( \12852 , \12847 , \12850 , \12851 );
xor \U$11870 ( \12853 , \12647 , \12651 );
xor \U$11871 ( \12854 , \12853 , \12656 );
xor \U$11872 ( \12855 , \12663 , \12667 );
xor \U$11873 ( \12856 , \12855 , \12672 );
and \U$11874 ( \12857 , \12854 , \12856 );
xor \U$11875 ( \12858 , \12680 , \12684 );
xor \U$11876 ( \12859 , \12858 , \12689 );
and \U$11877 ( \12860 , \12856 , \12859 );
and \U$11878 ( \12861 , \12854 , \12859 );
or \U$11879 ( \12862 , \12857 , \12860 , \12861 );
and \U$11880 ( \12863 , \12852 , \12862 );
and \U$11881 ( \12864 , \10226 , \1247 );
and \U$11882 ( \12865 , \10218 , \1245 );
nor \U$11883 ( \12866 , \12864 , \12865 );
xnor \U$11884 ( \12867 , \12866 , \1198 );
and \U$11885 ( \12868 , \10834 , \1146 );
and \U$11886 ( \12869 , \10829 , \1144 );
nor \U$11887 ( \12870 , \12868 , \12869 );
xnor \U$11888 ( \12871 , \12870 , \1105 );
and \U$11889 ( \12872 , \12867 , \12871 );
and \U$11890 ( \12873 , \11635 , \1076 );
and \U$11891 ( \12874 , \11015 , \1074 );
nor \U$11892 ( \12875 , \12873 , \12874 );
xnor \U$11893 ( \12876 , \12875 , \1046 );
and \U$11894 ( \12877 , \12871 , \12876 );
and \U$11895 ( \12878 , \12867 , \12876 );
or \U$11896 ( \12879 , \12872 , \12877 , \12878 );
xor \U$11897 ( \12880 , \12702 , \12706 );
xor \U$11898 ( \12881 , \12880 , \12711 );
and \U$11899 ( \12882 , \12879 , \12881 );
xor \U$11900 ( \12883 , \12718 , \12720 );
and \U$11901 ( \12884 , \12881 , \12883 );
and \U$11902 ( \12885 , \12879 , \12883 );
or \U$11903 ( \12886 , \12882 , \12884 , \12885 );
and \U$11904 ( \12887 , \12862 , \12886 );
and \U$11905 ( \12888 , \12852 , \12886 );
or \U$11906 ( \12889 , \12863 , \12887 , \12888 );
and \U$11907 ( \12890 , \4557 , \3992 );
and \U$11908 ( \12891 , \4349 , \3990 );
nor \U$11909 ( \12892 , \12890 , \12891 );
xnor \U$11910 ( \12893 , \12892 , \3787 );
and \U$11911 ( \12894 , \4684 , \3586 );
and \U$11912 ( \12895 , \4679 , \3584 );
nor \U$11913 ( \12896 , \12894 , \12895 );
xnor \U$11914 ( \12897 , \12896 , \3437 );
and \U$11915 ( \12898 , \12893 , \12897 );
and \U$11916 ( \12899 , \5137 , \3264 );
and \U$11917 ( \12900 , \4940 , \3262 );
nor \U$11918 ( \12901 , \12899 , \12900 );
xnor \U$11919 ( \12902 , \12901 , \3122 );
and \U$11920 ( \12903 , \12897 , \12902 );
and \U$11921 ( \12904 , \12893 , \12902 );
or \U$11922 ( \12905 , \12898 , \12903 , \12904 );
and \U$11923 ( \12906 , \2467 , \6314 );
and \U$11924 ( \12907 , \2459 , \6312 );
nor \U$11925 ( \12908 , \12906 , \12907 );
xnor \U$11926 ( \12909 , \12908 , \6073 );
and \U$11927 ( \12910 , \2715 , \5848 );
and \U$11928 ( \12911 , \2710 , \5846 );
nor \U$11929 ( \12912 , \12910 , \12911 );
xnor \U$11930 ( \12913 , \12912 , \5660 );
and \U$11931 ( \12914 , \12909 , \12913 );
and \U$11932 ( \12915 , \3045 , \5474 );
and \U$11933 ( \12916 , \2901 , \5472 );
nor \U$11934 ( \12917 , \12915 , \12916 );
xnor \U$11935 ( \12918 , \12917 , \5242 );
and \U$11936 ( \12919 , \12913 , \12918 );
and \U$11937 ( \12920 , \12909 , \12918 );
or \U$11938 ( \12921 , \12914 , \12919 , \12920 );
and \U$11939 ( \12922 , \12905 , \12921 );
and \U$11940 ( \12923 , \3334 , \5023 );
and \U$11941 ( \12924 , \3309 , \5021 );
nor \U$11942 ( \12925 , \12923 , \12924 );
xnor \U$11943 ( \12926 , \12925 , \4880 );
and \U$11944 ( \12927 , \3675 , \4700 );
and \U$11945 ( \12928 , \3508 , \4698 );
nor \U$11946 ( \12929 , \12927 , \12928 );
xnor \U$11947 ( \12930 , \12929 , \4454 );
and \U$11948 ( \12931 , \12926 , \12930 );
and \U$11949 ( \12932 , \3932 , \4305 );
and \U$11950 ( \12933 , \3813 , \4303 );
nor \U$11951 ( \12934 , \12932 , \12933 );
xnor \U$11952 ( \12935 , \12934 , \4118 );
and \U$11953 ( \12936 , \12930 , \12935 );
and \U$11954 ( \12937 , \12926 , \12935 );
or \U$11955 ( \12938 , \12931 , \12936 , \12937 );
and \U$11956 ( \12939 , \12921 , \12938 );
and \U$11957 ( \12940 , \12905 , \12938 );
or \U$11958 ( \12941 , \12922 , \12939 , \12940 );
and \U$11959 ( \12942 , \1942 , \7906 );
and \U$11960 ( \12943 , \1854 , \7904 );
nor \U$11961 ( \12944 , \12942 , \12943 );
xnor \U$11962 ( \12945 , \12944 , \7646 );
and \U$11963 ( \12946 , \2052 , \7412 );
and \U$11964 ( \12947 , \2047 , \7410 );
nor \U$11965 ( \12948 , \12946 , \12947 );
xnor \U$11966 ( \12949 , \12948 , \7097 );
and \U$11967 ( \12950 , \12945 , \12949 );
and \U$11968 ( \12951 , \2283 , \6903 );
and \U$11969 ( \12952 , \2168 , \6901 );
nor \U$11970 ( \12953 , \12951 , \12952 );
xnor \U$11971 ( \12954 , \12953 , \6563 );
and \U$11972 ( \12955 , \12949 , \12954 );
and \U$11973 ( \12956 , \12945 , \12954 );
or \U$11974 ( \12957 , \12950 , \12955 , \12956 );
and \U$11975 ( \12958 , \1093 , \11482 );
and \U$11976 ( \12959 , \1085 , \11479 );
nor \U$11977 ( \12960 , \12958 , \12959 );
xnor \U$11978 ( \12961 , \12960 , \10427 );
and \U$11979 ( \12962 , \1167 , \10669 );
and \U$11980 ( \12963 , \1162 , \10667 );
nor \U$11981 ( \12964 , \12962 , \12963 );
xnor \U$11982 ( \12965 , \12964 , \10430 );
and \U$11983 ( \12966 , \12961 , \12965 );
and \U$11984 ( \12967 , \1272 , \10101 );
and \U$11985 ( \12968 , \1221 , \10099 );
nor \U$11986 ( \12969 , \12967 , \12968 );
xnor \U$11987 ( \12970 , \12969 , \9791 );
and \U$11988 ( \12971 , \12965 , \12970 );
and \U$11989 ( \12972 , \12961 , \12970 );
or \U$11990 ( \12973 , \12966 , \12971 , \12972 );
and \U$11991 ( \12974 , \12957 , \12973 );
and \U$11992 ( \12975 , \1377 , \9564 );
and \U$11993 ( \12976 , \1349 , \9562 );
nor \U$11994 ( \12977 , \12975 , \12976 );
xnor \U$11995 ( \12978 , \12977 , \9193 );
and \U$11996 ( \12979 , \1531 , \9002 );
and \U$11997 ( \12980 , \1457 , \9000 );
nor \U$11998 ( \12981 , \12979 , \12980 );
xnor \U$11999 ( \12982 , \12981 , \8684 );
and \U$12000 ( \12983 , \12978 , \12982 );
and \U$12001 ( \12984 , \1656 , \8435 );
and \U$12002 ( \12985 , \1593 , \8433 );
nor \U$12003 ( \12986 , \12984 , \12985 );
xnor \U$12004 ( \12987 , \12986 , \8186 );
and \U$12005 ( \12988 , \12982 , \12987 );
and \U$12006 ( \12989 , \12978 , \12987 );
or \U$12007 ( \12990 , \12983 , \12988 , \12989 );
and \U$12008 ( \12991 , \12973 , \12990 );
and \U$12009 ( \12992 , \12957 , \12990 );
or \U$12010 ( \12993 , \12974 , \12991 , \12992 );
and \U$12011 ( \12994 , \12941 , \12993 );
and \U$12012 ( \12995 , \5447 , \2968 );
and \U$12013 ( \12996 , \5439 , \2966 );
nor \U$12014 ( \12997 , \12995 , \12996 );
xnor \U$12015 ( \12998 , \12997 , \2831 );
and \U$12016 ( \12999 , \5921 , \2762 );
and \U$12017 ( \13000 , \5916 , \2760 );
nor \U$12018 ( \13001 , \12999 , \13000 );
xnor \U$12019 ( \13002 , \13001 , \2610 );
and \U$12020 ( \13003 , \12998 , \13002 );
and \U$12021 ( \13004 , \6444 , \2494 );
and \U$12022 ( \13005 , \6185 , \2492 );
nor \U$12023 ( \13006 , \13004 , \13005 );
xnor \U$12024 ( \13007 , \13006 , \2338 );
and \U$12025 ( \13008 , \13002 , \13007 );
and \U$12026 ( \13009 , \12998 , \13007 );
or \U$12027 ( \13010 , \13003 , \13008 , \13009 );
and \U$12028 ( \13011 , \8795 , \1664 );
and \U$12029 ( \13012 , \8371 , \1662 );
nor \U$12030 ( \13013 , \13011 , \13012 );
xnor \U$12031 ( \13014 , \13013 , \1570 );
and \U$12032 ( \13015 , \9046 , \1494 );
and \U$12033 ( \13016 , \9041 , \1492 );
nor \U$12034 ( \13017 , \13015 , \13016 );
xnor \U$12035 ( \13018 , \13017 , \1422 );
and \U$12036 ( \13019 , \13014 , \13018 );
and \U$12037 ( \13020 , \9649 , \1360 );
and \U$12038 ( \13021 , \9365 , \1358 );
nor \U$12039 ( \13022 , \13020 , \13021 );
xnor \U$12040 ( \13023 , \13022 , \1317 );
and \U$12041 ( \13024 , \13018 , \13023 );
and \U$12042 ( \13025 , \13014 , \13023 );
or \U$12043 ( \13026 , \13019 , \13024 , \13025 );
and \U$12044 ( \13027 , \13010 , \13026 );
and \U$12045 ( \13028 , \6825 , \2222 );
and \U$12046 ( \13029 , \6816 , \2220 );
nor \U$12047 ( \13030 , \13028 , \13029 );
xnor \U$12048 ( \13031 , \13030 , \2109 );
and \U$12049 ( \13032 , \7370 , \2028 );
and \U$12050 ( \13033 , \7168 , \2026 );
nor \U$12051 ( \13034 , \13032 , \13033 );
xnor \U$12052 ( \13035 , \13034 , \1892 );
and \U$12053 ( \13036 , \13031 , \13035 );
and \U$12054 ( \13037 , \7845 , \1828 );
and \U$12055 ( \13038 , \7673 , \1826 );
nor \U$12056 ( \13039 , \13037 , \13038 );
xnor \U$12057 ( \13040 , \13039 , \1750 );
and \U$12058 ( \13041 , \13035 , \13040 );
and \U$12059 ( \13042 , \13031 , \13040 );
or \U$12060 ( \13043 , \13036 , \13041 , \13042 );
and \U$12061 ( \13044 , \13026 , \13043 );
and \U$12062 ( \13045 , \13010 , \13043 );
or \U$12063 ( \13046 , \13027 , \13044 , \13045 );
and \U$12064 ( \13047 , \12993 , \13046 );
and \U$12065 ( \13048 , \12941 , \13046 );
or \U$12066 ( \13049 , \12994 , \13047 , \13048 );
and \U$12067 ( \13050 , \12889 , \13049 );
xor \U$12068 ( \13051 , \12598 , \12602 );
xor \U$12069 ( \13052 , \13051 , \12607 );
xor \U$12070 ( \13053 , \12614 , \12618 );
xor \U$12071 ( \13054 , \13053 , \12623 );
and \U$12072 ( \13055 , \13052 , \13054 );
xor \U$12073 ( \13056 , \12631 , \12635 );
xor \U$12074 ( \13057 , \13056 , \1009 );
and \U$12075 ( \13058 , \13054 , \13057 );
and \U$12076 ( \13059 , \13052 , \13057 );
or \U$12077 ( \13060 , \13055 , \13058 , \13059 );
xor \U$12078 ( \13061 , \12246 , \12250 );
xor \U$12079 ( \13062 , \13061 , \12255 );
and \U$12080 ( \13063 , \13060 , \13062 );
xor \U$12081 ( \13064 , \12756 , \12758 );
xor \U$12082 ( \13065 , \13064 , \12761 );
and \U$12083 ( \13066 , \13062 , \13065 );
and \U$12084 ( \13067 , \13060 , \13065 );
or \U$12085 ( \13068 , \13063 , \13066 , \13067 );
and \U$12086 ( \13069 , \13049 , \13068 );
and \U$12087 ( \13070 , \12889 , \13068 );
or \U$12088 ( \13071 , \13050 , \13069 , \13070 );
xor \U$12089 ( \13072 , \12558 , \12574 );
xor \U$12090 ( \13073 , \13072 , \12591 );
xor \U$12091 ( \13074 , \12610 , \12626 );
xor \U$12092 ( \13075 , \13074 , \12639 );
and \U$12093 ( \13076 , \13073 , \13075 );
xor \U$12094 ( \13077 , \12659 , \12675 );
xor \U$12095 ( \13078 , \13077 , \12692 );
and \U$12096 ( \13079 , \13075 , \13078 );
and \U$12097 ( \13080 , \13073 , \13078 );
or \U$12098 ( \13081 , \13076 , \13079 , \13080 );
xor \U$12099 ( \13082 , \12714 , \12721 );
xor \U$12100 ( \13083 , \13082 , \12726 );
xor \U$12101 ( \13084 , \12731 , \12733 );
xor \U$12102 ( \13085 , \13084 , \12736 );
and \U$12103 ( \13086 , \13083 , \13085 );
xor \U$12104 ( \13087 , \12742 , \12744 );
xor \U$12105 ( \13088 , \13087 , \12747 );
and \U$12106 ( \13089 , \13085 , \13088 );
and \U$12107 ( \13090 , \13083 , \13088 );
or \U$12108 ( \13091 , \13086 , \13089 , \13090 );
and \U$12109 ( \13092 , \13081 , \13091 );
xor \U$12110 ( \13093 , \12347 , \12363 );
xor \U$12111 ( \13094 , \13093 , \12380 );
and \U$12112 ( \13095 , \13091 , \13094 );
and \U$12113 ( \13096 , \13081 , \13094 );
or \U$12114 ( \13097 , \13092 , \13095 , \13096 );
and \U$12115 ( \13098 , \13071 , \13097 );
xor \U$12116 ( \13099 , \12242 , \12258 );
xor \U$12117 ( \13100 , \13099 , \12275 );
xor \U$12118 ( \13101 , \12777 , \12779 );
xor \U$12119 ( \13102 , \13101 , \12782 );
and \U$12120 ( \13103 , \13100 , \13102 );
xor \U$12121 ( \13104 , \12764 , \12766 );
xor \U$12122 ( \13105 , \13104 , \12769 );
and \U$12123 ( \13106 , \13102 , \13105 );
and \U$12124 ( \13107 , \13100 , \13105 );
or \U$12125 ( \13108 , \13103 , \13106 , \13107 );
and \U$12126 ( \13109 , \13097 , \13108 );
and \U$12127 ( \13110 , \13071 , \13108 );
or \U$12128 ( \13111 , \13098 , \13109 , \13110 );
xor \U$12129 ( \13112 , \12698 , \12753 );
xor \U$12130 ( \13113 , \13112 , \12772 );
xor \U$12131 ( \13114 , \12785 , \12787 );
xor \U$12132 ( \13115 , \13114 , \12790 );
and \U$12133 ( \13116 , \13113 , \13115 );
xor \U$12134 ( \13117 , \12796 , \12798 );
xor \U$12135 ( \13118 , \13117 , \12801 );
and \U$12136 ( \13119 , \13115 , \13118 );
and \U$12137 ( \13120 , \13113 , \13118 );
or \U$12138 ( \13121 , \13116 , \13119 , \13120 );
and \U$12139 ( \13122 , \13111 , \13121 );
xor \U$12140 ( \13123 , \12465 , \12475 );
xor \U$12141 ( \13124 , \13123 , \12478 );
and \U$12142 ( \13125 , \13121 , \13124 );
and \U$12143 ( \13126 , \13111 , \13124 );
or \U$12144 ( \13127 , \13122 , \13125 , \13126 );
xor \U$12145 ( \13128 , \12386 , \12434 );
xor \U$12146 ( \13129 , \13128 , \12452 );
xor \U$12147 ( \13130 , \12775 , \12793 );
xor \U$12148 ( \13131 , \13130 , \12804 );
and \U$12149 ( \13132 , \13129 , \13131 );
xor \U$12150 ( \13133 , \12809 , \12811 );
xor \U$12151 ( \13134 , \13133 , \12814 );
and \U$12152 ( \13135 , \13131 , \13134 );
and \U$12153 ( \13136 , \13129 , \13134 );
or \U$12154 ( \13137 , \13132 , \13135 , \13136 );
and \U$12155 ( \13138 , \13127 , \13137 );
xor \U$12156 ( \13139 , \12497 , \12499 );
xor \U$12157 ( \13140 , \13139 , \12502 );
and \U$12158 ( \13141 , \13137 , \13140 );
and \U$12159 ( \13142 , \13127 , \13140 );
or \U$12160 ( \13143 , \13138 , \13141 , \13142 );
xor \U$12161 ( \13144 , \12455 , \12481 );
xor \U$12162 ( \13145 , \13144 , \12492 );
xor \U$12163 ( \13146 , \12807 , \12817 );
xor \U$12164 ( \13147 , \13146 , \12820 );
and \U$12165 ( \13148 , \13145 , \13147 );
and \U$12166 ( \13149 , \13143 , \13148 );
xor \U$12167 ( \13150 , \12823 , \12825 );
xor \U$12168 ( \13151 , \13150 , \12828 );
and \U$12169 ( \13152 , \13148 , \13151 );
and \U$12170 ( \13153 , \13143 , \13151 );
or \U$12171 ( \13154 , \13149 , \13152 , \13153 );
and \U$12172 ( \13155 , \12842 , \13154 );
xor \U$12173 ( \13156 , \12842 , \13154 );
xor \U$12174 ( \13157 , \13143 , \13148 );
xor \U$12175 ( \13158 , \13157 , \13151 );
xor \U$12176 ( \13159 , \12893 , \12897 );
xor \U$12177 ( \13160 , \13159 , \12902 );
xor \U$12178 ( \13161 , \12998 , \13002 );
xor \U$12179 ( \13162 , \13161 , \13007 );
and \U$12180 ( \13163 , \13160 , \13162 );
xor \U$12181 ( \13164 , \13031 , \13035 );
xor \U$12182 ( \13165 , \13164 , \13040 );
and \U$12183 ( \13166 , \13162 , \13165 );
and \U$12184 ( \13167 , \13160 , \13165 );
or \U$12185 ( \13168 , \13163 , \13166 , \13167 );
and \U$12186 ( \13169 , \10218 , \1360 );
and \U$12187 ( \13170 , \9649 , \1358 );
nor \U$12188 ( \13171 , \13169 , \13170 );
xnor \U$12189 ( \13172 , \13171 , \1317 );
and \U$12190 ( \13173 , \10829 , \1247 );
and \U$12191 ( \13174 , \10226 , \1245 );
nor \U$12192 ( \13175 , \13173 , \13174 );
xnor \U$12193 ( \13176 , \13175 , \1198 );
and \U$12194 ( \13177 , \13172 , \13176 );
and \U$12195 ( \13178 , \11015 , \1146 );
and \U$12196 ( \13179 , \10834 , \1144 );
nor \U$12197 ( \13180 , \13178 , \13179 );
xnor \U$12198 ( \13181 , \13180 , \1105 );
and \U$12199 ( \13182 , \13176 , \13181 );
and \U$12200 ( \13183 , \13172 , \13181 );
or \U$12201 ( \13184 , \13177 , \13182 , \13183 );
xor \U$12202 ( \13185 , \13014 , \13018 );
xor \U$12203 ( \13186 , \13185 , \13023 );
and \U$12204 ( \13187 , \13184 , \13186 );
xor \U$12205 ( \13188 , \12867 , \12871 );
xor \U$12206 ( \13189 , \13188 , \12876 );
and \U$12207 ( \13190 , \13186 , \13189 );
and \U$12208 ( \13191 , \13184 , \13189 );
or \U$12209 ( \13192 , \13187 , \13190 , \13191 );
and \U$12210 ( \13193 , \13168 , \13192 );
xor \U$12211 ( \13194 , \12945 , \12949 );
xor \U$12212 ( \13195 , \13194 , \12954 );
xor \U$12213 ( \13196 , \12909 , \12913 );
xor \U$12214 ( \13197 , \13196 , \12918 );
and \U$12215 ( \13198 , \13195 , \13197 );
xor \U$12216 ( \13199 , \12926 , \12930 );
xor \U$12217 ( \13200 , \13199 , \12935 );
and \U$12218 ( \13201 , \13197 , \13200 );
and \U$12219 ( \13202 , \13195 , \13200 );
or \U$12220 ( \13203 , \13198 , \13201 , \13202 );
and \U$12221 ( \13204 , \13192 , \13203 );
and \U$12222 ( \13205 , \13168 , \13203 );
or \U$12223 ( \13206 , \13193 , \13204 , \13205 );
and \U$12224 ( \13207 , \1854 , \8435 );
and \U$12225 ( \13208 , \1656 , \8433 );
nor \U$12226 ( \13209 , \13207 , \13208 );
xnor \U$12227 ( \13210 , \13209 , \8186 );
and \U$12228 ( \13211 , \2047 , \7906 );
and \U$12229 ( \13212 , \1942 , \7904 );
nor \U$12230 ( \13213 , \13211 , \13212 );
xnor \U$12231 ( \13214 , \13213 , \7646 );
and \U$12232 ( \13215 , \13210 , \13214 );
and \U$12233 ( \13216 , \2168 , \7412 );
and \U$12234 ( \13217 , \2052 , \7410 );
nor \U$12235 ( \13218 , \13216 , \13217 );
xnor \U$12236 ( \13219 , \13218 , \7097 );
and \U$12237 ( \13220 , \13214 , \13219 );
and \U$12238 ( \13221 , \13210 , \13219 );
or \U$12239 ( \13222 , \13215 , \13220 , \13221 );
and \U$12240 ( \13223 , \1162 , \11482 );
and \U$12241 ( \13224 , \1093 , \11479 );
nor \U$12242 ( \13225 , \13223 , \13224 );
xnor \U$12243 ( \13226 , \13225 , \10427 );
and \U$12244 ( \13227 , \1221 , \10669 );
and \U$12245 ( \13228 , \1167 , \10667 );
nor \U$12246 ( \13229 , \13227 , \13228 );
xnor \U$12247 ( \13230 , \13229 , \10430 );
and \U$12248 ( \13231 , \13226 , \13230 );
and \U$12249 ( \13232 , \13230 , \1046 );
and \U$12250 ( \13233 , \13226 , \1046 );
or \U$12251 ( \13234 , \13231 , \13232 , \13233 );
and \U$12252 ( \13235 , \13222 , \13234 );
and \U$12253 ( \13236 , \1349 , \10101 );
and \U$12254 ( \13237 , \1272 , \10099 );
nor \U$12255 ( \13238 , \13236 , \13237 );
xnor \U$12256 ( \13239 , \13238 , \9791 );
and \U$12257 ( \13240 , \1457 , \9564 );
and \U$12258 ( \13241 , \1377 , \9562 );
nor \U$12259 ( \13242 , \13240 , \13241 );
xnor \U$12260 ( \13243 , \13242 , \9193 );
and \U$12261 ( \13244 , \13239 , \13243 );
and \U$12262 ( \13245 , \1593 , \9002 );
and \U$12263 ( \13246 , \1531 , \9000 );
nor \U$12264 ( \13247 , \13245 , \13246 );
xnor \U$12265 ( \13248 , \13247 , \8684 );
and \U$12266 ( \13249 , \13243 , \13248 );
and \U$12267 ( \13250 , \13239 , \13248 );
or \U$12268 ( \13251 , \13244 , \13249 , \13250 );
and \U$12269 ( \13252 , \13234 , \13251 );
and \U$12270 ( \13253 , \13222 , \13251 );
or \U$12271 ( \13254 , \13235 , \13252 , \13253 );
and \U$12272 ( \13255 , \4349 , \4305 );
and \U$12273 ( \13256 , \3932 , \4303 );
nor \U$12274 ( \13257 , \13255 , \13256 );
xnor \U$12275 ( \13258 , \13257 , \4118 );
and \U$12276 ( \13259 , \4679 , \3992 );
and \U$12277 ( \13260 , \4557 , \3990 );
nor \U$12278 ( \13261 , \13259 , \13260 );
xnor \U$12279 ( \13262 , \13261 , \3787 );
and \U$12280 ( \13263 , \13258 , \13262 );
and \U$12281 ( \13264 , \4940 , \3586 );
and \U$12282 ( \13265 , \4684 , \3584 );
nor \U$12283 ( \13266 , \13264 , \13265 );
xnor \U$12284 ( \13267 , \13266 , \3437 );
and \U$12285 ( \13268 , \13262 , \13267 );
and \U$12286 ( \13269 , \13258 , \13267 );
or \U$12287 ( \13270 , \13263 , \13268 , \13269 );
and \U$12288 ( \13271 , \3309 , \5474 );
and \U$12289 ( \13272 , \3045 , \5472 );
nor \U$12290 ( \13273 , \13271 , \13272 );
xnor \U$12291 ( \13274 , \13273 , \5242 );
and \U$12292 ( \13275 , \3508 , \5023 );
and \U$12293 ( \13276 , \3334 , \5021 );
nor \U$12294 ( \13277 , \13275 , \13276 );
xnor \U$12295 ( \13278 , \13277 , \4880 );
and \U$12296 ( \13279 , \13274 , \13278 );
and \U$12297 ( \13280 , \3813 , \4700 );
and \U$12298 ( \13281 , \3675 , \4698 );
nor \U$12299 ( \13282 , \13280 , \13281 );
xnor \U$12300 ( \13283 , \13282 , \4454 );
and \U$12301 ( \13284 , \13278 , \13283 );
and \U$12302 ( \13285 , \13274 , \13283 );
or \U$12303 ( \13286 , \13279 , \13284 , \13285 );
and \U$12304 ( \13287 , \13270 , \13286 );
and \U$12305 ( \13288 , \2459 , \6903 );
and \U$12306 ( \13289 , \2283 , \6901 );
nor \U$12307 ( \13290 , \13288 , \13289 );
xnor \U$12308 ( \13291 , \13290 , \6563 );
and \U$12309 ( \13292 , \2710 , \6314 );
and \U$12310 ( \13293 , \2467 , \6312 );
nor \U$12311 ( \13294 , \13292 , \13293 );
xnor \U$12312 ( \13295 , \13294 , \6073 );
and \U$12313 ( \13296 , \13291 , \13295 );
and \U$12314 ( \13297 , \2901 , \5848 );
and \U$12315 ( \13298 , \2715 , \5846 );
nor \U$12316 ( \13299 , \13297 , \13298 );
xnor \U$12317 ( \13300 , \13299 , \5660 );
and \U$12318 ( \13301 , \13295 , \13300 );
and \U$12319 ( \13302 , \13291 , \13300 );
or \U$12320 ( \13303 , \13296 , \13301 , \13302 );
and \U$12321 ( \13304 , \13286 , \13303 );
and \U$12322 ( \13305 , \13270 , \13303 );
or \U$12323 ( \13306 , \13287 , \13304 , \13305 );
and \U$12324 ( \13307 , \13254 , \13306 );
and \U$12325 ( \13308 , \5439 , \3264 );
and \U$12326 ( \13309 , \5137 , \3262 );
nor \U$12327 ( \13310 , \13308 , \13309 );
xnor \U$12328 ( \13311 , \13310 , \3122 );
and \U$12329 ( \13312 , \5916 , \2968 );
and \U$12330 ( \13313 , \5447 , \2966 );
nor \U$12331 ( \13314 , \13312 , \13313 );
xnor \U$12332 ( \13315 , \13314 , \2831 );
and \U$12333 ( \13316 , \13311 , \13315 );
and \U$12334 ( \13317 , \6185 , \2762 );
and \U$12335 ( \13318 , \5921 , \2760 );
nor \U$12336 ( \13319 , \13317 , \13318 );
xnor \U$12337 ( \13320 , \13319 , \2610 );
and \U$12338 ( \13321 , \13315 , \13320 );
and \U$12339 ( \13322 , \13311 , \13320 );
or \U$12340 ( \13323 , \13316 , \13321 , \13322 );
and \U$12341 ( \13324 , \6816 , \2494 );
and \U$12342 ( \13325 , \6444 , \2492 );
nor \U$12343 ( \13326 , \13324 , \13325 );
xnor \U$12344 ( \13327 , \13326 , \2338 );
and \U$12345 ( \13328 , \7168 , \2222 );
and \U$12346 ( \13329 , \6825 , \2220 );
nor \U$12347 ( \13330 , \13328 , \13329 );
xnor \U$12348 ( \13331 , \13330 , \2109 );
and \U$12349 ( \13332 , \13327 , \13331 );
and \U$12350 ( \13333 , \7673 , \2028 );
and \U$12351 ( \13334 , \7370 , \2026 );
nor \U$12352 ( \13335 , \13333 , \13334 );
xnor \U$12353 ( \13336 , \13335 , \1892 );
and \U$12354 ( \13337 , \13331 , \13336 );
and \U$12355 ( \13338 , \13327 , \13336 );
or \U$12356 ( \13339 , \13332 , \13337 , \13338 );
and \U$12357 ( \13340 , \13323 , \13339 );
and \U$12358 ( \13341 , \8371 , \1828 );
and \U$12359 ( \13342 , \7845 , \1826 );
nor \U$12360 ( \13343 , \13341 , \13342 );
xnor \U$12361 ( \13344 , \13343 , \1750 );
and \U$12362 ( \13345 , \9041 , \1664 );
and \U$12363 ( \13346 , \8795 , \1662 );
nor \U$12364 ( \13347 , \13345 , \13346 );
xnor \U$12365 ( \13348 , \13347 , \1570 );
and \U$12366 ( \13349 , \13344 , \13348 );
and \U$12367 ( \13350 , \9365 , \1494 );
and \U$12368 ( \13351 , \9046 , \1492 );
nor \U$12369 ( \13352 , \13350 , \13351 );
xnor \U$12370 ( \13353 , \13352 , \1422 );
and \U$12371 ( \13354 , \13348 , \13353 );
and \U$12372 ( \13355 , \13344 , \13353 );
or \U$12373 ( \13356 , \13349 , \13354 , \13355 );
and \U$12374 ( \13357 , \13339 , \13356 );
and \U$12375 ( \13358 , \13323 , \13356 );
or \U$12376 ( \13359 , \13340 , \13357 , \13358 );
and \U$12377 ( \13360 , \13306 , \13359 );
and \U$12378 ( \13361 , \13254 , \13359 );
or \U$12379 ( \13362 , \13307 , \13360 , \13361 );
and \U$12380 ( \13363 , \13206 , \13362 );
xor \U$12381 ( \13364 , \13052 , \13054 );
xor \U$12382 ( \13365 , \13364 , \13057 );
xor \U$12383 ( \13366 , \12844 , \12846 );
xor \U$12384 ( \13367 , \13366 , \12849 );
and \U$12385 ( \13368 , \13365 , \13367 );
xor \U$12386 ( \13369 , \12854 , \12856 );
xor \U$12387 ( \13370 , \13369 , \12859 );
and \U$12388 ( \13371 , \13367 , \13370 );
and \U$12389 ( \13372 , \13365 , \13370 );
or \U$12390 ( \13373 , \13368 , \13371 , \13372 );
and \U$12391 ( \13374 , \13362 , \13373 );
and \U$12392 ( \13375 , \13206 , \13373 );
or \U$12393 ( \13376 , \13363 , \13374 , \13375 );
xor \U$12394 ( \13377 , \12905 , \12921 );
xor \U$12395 ( \13378 , \13377 , \12938 );
xor \U$12396 ( \13379 , \13010 , \13026 );
xor \U$12397 ( \13380 , \13379 , \13043 );
and \U$12398 ( \13381 , \13378 , \13380 );
xor \U$12399 ( \13382 , \12879 , \12881 );
xor \U$12400 ( \13383 , \13382 , \12883 );
and \U$12401 ( \13384 , \13380 , \13383 );
and \U$12402 ( \13385 , \13378 , \13383 );
or \U$12403 ( \13386 , \13381 , \13384 , \13385 );
xor \U$12404 ( \13387 , \13073 , \13075 );
xor \U$12405 ( \13388 , \13387 , \13078 );
and \U$12406 ( \13389 , \13386 , \13388 );
xor \U$12407 ( \13390 , \13083 , \13085 );
xor \U$12408 ( \13391 , \13390 , \13088 );
and \U$12409 ( \13392 , \13388 , \13391 );
and \U$12410 ( \13393 , \13386 , \13391 );
or \U$12411 ( \13394 , \13389 , \13392 , \13393 );
and \U$12412 ( \13395 , \13376 , \13394 );
xor \U$12413 ( \13396 , \12852 , \12862 );
xor \U$12414 ( \13397 , \13396 , \12886 );
xor \U$12415 ( \13398 , \12941 , \12993 );
xor \U$12416 ( \13399 , \13398 , \13046 );
and \U$12417 ( \13400 , \13397 , \13399 );
xor \U$12418 ( \13401 , \13060 , \13062 );
xor \U$12419 ( \13402 , \13401 , \13065 );
and \U$12420 ( \13403 , \13399 , \13402 );
and \U$12421 ( \13404 , \13397 , \13402 );
or \U$12422 ( \13405 , \13400 , \13403 , \13404 );
and \U$12423 ( \13406 , \13394 , \13405 );
and \U$12424 ( \13407 , \13376 , \13405 );
or \U$12425 ( \13408 , \13395 , \13406 , \13407 );
xor \U$12426 ( \13409 , \12594 , \12642 );
xor \U$12427 ( \13410 , \13409 , \12695 );
xor \U$12428 ( \13411 , \12729 , \12739 );
xor \U$12429 ( \13412 , \13411 , \12750 );
and \U$12430 ( \13413 , \13410 , \13412 );
xor \U$12431 ( \13414 , \13100 , \13102 );
xor \U$12432 ( \13415 , \13414 , \13105 );
and \U$12433 ( \13416 , \13412 , \13415 );
and \U$12434 ( \13417 , \13410 , \13415 );
or \U$12435 ( \13418 , \13413 , \13416 , \13417 );
and \U$12436 ( \13419 , \13408 , \13418 );
xor \U$12437 ( \13420 , \13113 , \13115 );
xor \U$12438 ( \13421 , \13420 , \13118 );
and \U$12439 ( \13422 , \13418 , \13421 );
and \U$12440 ( \13423 , \13408 , \13421 );
or \U$12441 ( \13424 , \13419 , \13422 , \13423 );
xor \U$12442 ( \13425 , \13111 , \13121 );
xor \U$12443 ( \13426 , \13425 , \13124 );
and \U$12444 ( \13427 , \13424 , \13426 );
xor \U$12445 ( \13428 , \13129 , \13131 );
xor \U$12446 ( \13429 , \13428 , \13134 );
and \U$12447 ( \13430 , \13426 , \13429 );
and \U$12448 ( \13431 , \13424 , \13429 );
or \U$12449 ( \13432 , \13427 , \13430 , \13431 );
xor \U$12450 ( \13433 , \13127 , \13137 );
xor \U$12451 ( \13434 , \13433 , \13140 );
and \U$12452 ( \13435 , \13432 , \13434 );
xor \U$12453 ( \13436 , \13145 , \13147 );
and \U$12454 ( \13437 , \13434 , \13436 );
and \U$12455 ( \13438 , \13432 , \13436 );
or \U$12456 ( \13439 , \13435 , \13437 , \13438 );
and \U$12457 ( \13440 , \13158 , \13439 );
xor \U$12458 ( \13441 , \13158 , \13439 );
xor \U$12459 ( \13442 , \13432 , \13434 );
xor \U$12460 ( \13443 , \13442 , \13436 );
and \U$12461 ( \13444 , \3675 , \5023 );
and \U$12462 ( \13445 , \3508 , \5021 );
nor \U$12463 ( \13446 , \13444 , \13445 );
xnor \U$12464 ( \13447 , \13446 , \4880 );
and \U$12465 ( \13448 , \3932 , \4700 );
and \U$12466 ( \13449 , \3813 , \4698 );
nor \U$12467 ( \13450 , \13448 , \13449 );
xnor \U$12468 ( \13451 , \13450 , \4454 );
and \U$12469 ( \13452 , \13447 , \13451 );
and \U$12470 ( \13453 , \4557 , \4305 );
and \U$12471 ( \13454 , \4349 , \4303 );
nor \U$12472 ( \13455 , \13453 , \13454 );
xnor \U$12473 ( \13456 , \13455 , \4118 );
and \U$12474 ( \13457 , \13451 , \13456 );
and \U$12475 ( \13458 , \13447 , \13456 );
or \U$12476 ( \13459 , \13452 , \13457 , \13458 );
and \U$12477 ( \13460 , \4684 , \3992 );
and \U$12478 ( \13461 , \4679 , \3990 );
nor \U$12479 ( \13462 , \13460 , \13461 );
xnor \U$12480 ( \13463 , \13462 , \3787 );
and \U$12481 ( \13464 , \5137 , \3586 );
and \U$12482 ( \13465 , \4940 , \3584 );
nor \U$12483 ( \13466 , \13464 , \13465 );
xnor \U$12484 ( \13467 , \13466 , \3437 );
and \U$12485 ( \13468 , \13463 , \13467 );
and \U$12486 ( \13469 , \5447 , \3264 );
and \U$12487 ( \13470 , \5439 , \3262 );
nor \U$12488 ( \13471 , \13469 , \13470 );
xnor \U$12489 ( \13472 , \13471 , \3122 );
and \U$12490 ( \13473 , \13467 , \13472 );
and \U$12491 ( \13474 , \13463 , \13472 );
or \U$12492 ( \13475 , \13468 , \13473 , \13474 );
and \U$12493 ( \13476 , \13459 , \13475 );
and \U$12494 ( \13477 , \2715 , \6314 );
and \U$12495 ( \13478 , \2710 , \6312 );
nor \U$12496 ( \13479 , \13477 , \13478 );
xnor \U$12497 ( \13480 , \13479 , \6073 );
and \U$12498 ( \13481 , \3045 , \5848 );
and \U$12499 ( \13482 , \2901 , \5846 );
nor \U$12500 ( \13483 , \13481 , \13482 );
xnor \U$12501 ( \13484 , \13483 , \5660 );
and \U$12502 ( \13485 , \13480 , \13484 );
and \U$12503 ( \13486 , \3334 , \5474 );
and \U$12504 ( \13487 , \3309 , \5472 );
nor \U$12505 ( \13488 , \13486 , \13487 );
xnor \U$12506 ( \13489 , \13488 , \5242 );
and \U$12507 ( \13490 , \13484 , \13489 );
and \U$12508 ( \13491 , \13480 , \13489 );
or \U$12509 ( \13492 , \13485 , \13490 , \13491 );
and \U$12510 ( \13493 , \13475 , \13492 );
and \U$12511 ( \13494 , \13459 , \13492 );
or \U$12512 ( \13495 , \13476 , \13493 , \13494 );
and \U$12513 ( \13496 , \7370 , \2222 );
and \U$12514 ( \13497 , \7168 , \2220 );
nor \U$12515 ( \13498 , \13496 , \13497 );
xnor \U$12516 ( \13499 , \13498 , \2109 );
and \U$12517 ( \13500 , \7845 , \2028 );
and \U$12518 ( \13501 , \7673 , \2026 );
nor \U$12519 ( \13502 , \13500 , \13501 );
xnor \U$12520 ( \13503 , \13502 , \1892 );
and \U$12521 ( \13504 , \13499 , \13503 );
and \U$12522 ( \13505 , \8795 , \1828 );
and \U$12523 ( \13506 , \8371 , \1826 );
nor \U$12524 ( \13507 , \13505 , \13506 );
xnor \U$12525 ( \13508 , \13507 , \1750 );
and \U$12526 ( \13509 , \13503 , \13508 );
and \U$12527 ( \13510 , \13499 , \13508 );
or \U$12528 ( \13511 , \13504 , \13509 , \13510 );
and \U$12529 ( \13512 , \9046 , \1664 );
and \U$12530 ( \13513 , \9041 , \1662 );
nor \U$12531 ( \13514 , \13512 , \13513 );
xnor \U$12532 ( \13515 , \13514 , \1570 );
and \U$12533 ( \13516 , \9649 , \1494 );
and \U$12534 ( \13517 , \9365 , \1492 );
nor \U$12535 ( \13518 , \13516 , \13517 );
xnor \U$12536 ( \13519 , \13518 , \1422 );
and \U$12537 ( \13520 , \13515 , \13519 );
and \U$12538 ( \13521 , \10226 , \1360 );
and \U$12539 ( \13522 , \10218 , \1358 );
nor \U$12540 ( \13523 , \13521 , \13522 );
xnor \U$12541 ( \13524 , \13523 , \1317 );
and \U$12542 ( \13525 , \13519 , \13524 );
and \U$12543 ( \13526 , \13515 , \13524 );
or \U$12544 ( \13527 , \13520 , \13525 , \13526 );
and \U$12545 ( \13528 , \13511 , \13527 );
and \U$12546 ( \13529 , \5921 , \2968 );
and \U$12547 ( \13530 , \5916 , \2966 );
nor \U$12548 ( \13531 , \13529 , \13530 );
xnor \U$12549 ( \13532 , \13531 , \2831 );
and \U$12550 ( \13533 , \6444 , \2762 );
and \U$12551 ( \13534 , \6185 , \2760 );
nor \U$12552 ( \13535 , \13533 , \13534 );
xnor \U$12553 ( \13536 , \13535 , \2610 );
and \U$12554 ( \13537 , \13532 , \13536 );
and \U$12555 ( \13538 , \6825 , \2494 );
and \U$12556 ( \13539 , \6816 , \2492 );
nor \U$12557 ( \13540 , \13538 , \13539 );
xnor \U$12558 ( \13541 , \13540 , \2338 );
and \U$12559 ( \13542 , \13536 , \13541 );
and \U$12560 ( \13543 , \13532 , \13541 );
or \U$12561 ( \13544 , \13537 , \13542 , \13543 );
and \U$12562 ( \13545 , \13527 , \13544 );
and \U$12563 ( \13546 , \13511 , \13544 );
or \U$12564 ( \13547 , \13528 , \13545 , \13546 );
and \U$12565 ( \13548 , \13495 , \13547 );
and \U$12566 ( \13549 , \1167 , \11482 );
and \U$12567 ( \13550 , \1162 , \11479 );
nor \U$12568 ( \13551 , \13549 , \13550 );
xnor \U$12569 ( \13552 , \13551 , \10427 );
and \U$12570 ( \13553 , \1272 , \10669 );
and \U$12571 ( \13554 , \1221 , \10667 );
nor \U$12572 ( \13555 , \13553 , \13554 );
xnor \U$12573 ( \13556 , \13555 , \10430 );
and \U$12574 ( \13557 , \13552 , \13556 );
and \U$12575 ( \13558 , \1377 , \10101 );
and \U$12576 ( \13559 , \1349 , \10099 );
nor \U$12577 ( \13560 , \13558 , \13559 );
xnor \U$12578 ( \13561 , \13560 , \9791 );
and \U$12579 ( \13562 , \13556 , \13561 );
and \U$12580 ( \13563 , \13552 , \13561 );
or \U$12581 ( \13564 , \13557 , \13562 , \13563 );
and \U$12582 ( \13565 , \1531 , \9564 );
and \U$12583 ( \13566 , \1457 , \9562 );
nor \U$12584 ( \13567 , \13565 , \13566 );
xnor \U$12585 ( \13568 , \13567 , \9193 );
and \U$12586 ( \13569 , \1656 , \9002 );
and \U$12587 ( \13570 , \1593 , \9000 );
nor \U$12588 ( \13571 , \13569 , \13570 );
xnor \U$12589 ( \13572 , \13571 , \8684 );
and \U$12590 ( \13573 , \13568 , \13572 );
and \U$12591 ( \13574 , \1942 , \8435 );
and \U$12592 ( \13575 , \1854 , \8433 );
nor \U$12593 ( \13576 , \13574 , \13575 );
xnor \U$12594 ( \13577 , \13576 , \8186 );
and \U$12595 ( \13578 , \13572 , \13577 );
and \U$12596 ( \13579 , \13568 , \13577 );
or \U$12597 ( \13580 , \13573 , \13578 , \13579 );
and \U$12598 ( \13581 , \13564 , \13580 );
and \U$12599 ( \13582 , \2052 , \7906 );
and \U$12600 ( \13583 , \2047 , \7904 );
nor \U$12601 ( \13584 , \13582 , \13583 );
xnor \U$12602 ( \13585 , \13584 , \7646 );
and \U$12603 ( \13586 , \2283 , \7412 );
and \U$12604 ( \13587 , \2168 , \7410 );
nor \U$12605 ( \13588 , \13586 , \13587 );
xnor \U$12606 ( \13589 , \13588 , \7097 );
and \U$12607 ( \13590 , \13585 , \13589 );
and \U$12608 ( \13591 , \2467 , \6903 );
and \U$12609 ( \13592 , \2459 , \6901 );
nor \U$12610 ( \13593 , \13591 , \13592 );
xnor \U$12611 ( \13594 , \13593 , \6563 );
and \U$12612 ( \13595 , \13589 , \13594 );
and \U$12613 ( \13596 , \13585 , \13594 );
or \U$12614 ( \13597 , \13590 , \13595 , \13596 );
and \U$12615 ( \13598 , \13580 , \13597 );
and \U$12616 ( \13599 , \13564 , \13597 );
or \U$12617 ( \13600 , \13581 , \13598 , \13599 );
and \U$12618 ( \13601 , \13547 , \13600 );
and \U$12619 ( \13602 , \13495 , \13600 );
or \U$12620 ( \13603 , \13548 , \13601 , \13602 );
xor \U$12621 ( \13604 , \13210 , \13214 );
xor \U$12622 ( \13605 , \13604 , \13219 );
xor \U$12623 ( \13606 , \13274 , \13278 );
xor \U$12624 ( \13607 , \13606 , \13283 );
and \U$12625 ( \13608 , \13605 , \13607 );
xor \U$12626 ( \13609 , \13291 , \13295 );
xor \U$12627 ( \13610 , \13609 , \13300 );
and \U$12628 ( \13611 , \13607 , \13610 );
and \U$12629 ( \13612 , \13605 , \13610 );
or \U$12630 ( \13613 , \13608 , \13611 , \13612 );
xor \U$12631 ( \13614 , \13258 , \13262 );
xor \U$12632 ( \13615 , \13614 , \13267 );
xor \U$12633 ( \13616 , \13311 , \13315 );
xor \U$12634 ( \13617 , \13616 , \13320 );
and \U$12635 ( \13618 , \13615 , \13617 );
xor \U$12636 ( \13619 , \13327 , \13331 );
xor \U$12637 ( \13620 , \13619 , \13336 );
and \U$12638 ( \13621 , \13617 , \13620 );
and \U$12639 ( \13622 , \13615 , \13620 );
or \U$12640 ( \13623 , \13618 , \13621 , \13622 );
and \U$12641 ( \13624 , \13613 , \13623 );
nand \U$12642 ( \13625 , \11635 , \1074 );
xnor \U$12643 ( \13626 , \13625 , \1046 );
xor \U$12644 ( \13627 , \13344 , \13348 );
xor \U$12645 ( \13628 , \13627 , \13353 );
and \U$12646 ( \13629 , \13626 , \13628 );
xor \U$12647 ( \13630 , \13172 , \13176 );
xor \U$12648 ( \13631 , \13630 , \13181 );
and \U$12649 ( \13632 , \13628 , \13631 );
and \U$12650 ( \13633 , \13626 , \13631 );
or \U$12651 ( \13634 , \13629 , \13632 , \13633 );
and \U$12652 ( \13635 , \13623 , \13634 );
and \U$12653 ( \13636 , \13613 , \13634 );
or \U$12654 ( \13637 , \13624 , \13635 , \13636 );
and \U$12655 ( \13638 , \13603 , \13637 );
xor \U$12656 ( \13639 , \12961 , \12965 );
xor \U$12657 ( \13640 , \13639 , \12970 );
xor \U$12658 ( \13641 , \12978 , \12982 );
xor \U$12659 ( \13642 , \13641 , \12987 );
and \U$12660 ( \13643 , \13640 , \13642 );
xor \U$12661 ( \13644 , \13195 , \13197 );
xor \U$12662 ( \13645 , \13644 , \13200 );
and \U$12663 ( \13646 , \13642 , \13645 );
and \U$12664 ( \13647 , \13640 , \13645 );
or \U$12665 ( \13648 , \13643 , \13646 , \13647 );
and \U$12666 ( \13649 , \13637 , \13648 );
and \U$12667 ( \13650 , \13603 , \13648 );
or \U$12668 ( \13651 , \13638 , \13649 , \13650 );
xor \U$12669 ( \13652 , \13168 , \13192 );
xor \U$12670 ( \13653 , \13652 , \13203 );
xor \U$12671 ( \13654 , \13254 , \13306 );
xor \U$12672 ( \13655 , \13654 , \13359 );
and \U$12673 ( \13656 , \13653 , \13655 );
xor \U$12674 ( \13657 , \13365 , \13367 );
xor \U$12675 ( \13658 , \13657 , \13370 );
and \U$12676 ( \13659 , \13655 , \13658 );
and \U$12677 ( \13660 , \13653 , \13658 );
or \U$12678 ( \13661 , \13656 , \13659 , \13660 );
and \U$12679 ( \13662 , \13651 , \13661 );
xor \U$12680 ( \13663 , \13323 , \13339 );
xor \U$12681 ( \13664 , \13663 , \13356 );
xor \U$12682 ( \13665 , \13160 , \13162 );
xor \U$12683 ( \13666 , \13665 , \13165 );
and \U$12684 ( \13667 , \13664 , \13666 );
xor \U$12685 ( \13668 , \13184 , \13186 );
xor \U$12686 ( \13669 , \13668 , \13189 );
and \U$12687 ( \13670 , \13666 , \13669 );
and \U$12688 ( \13671 , \13664 , \13669 );
or \U$12689 ( \13672 , \13667 , \13670 , \13671 );
xor \U$12690 ( \13673 , \12957 , \12973 );
xor \U$12691 ( \13674 , \13673 , \12990 );
and \U$12692 ( \13675 , \13672 , \13674 );
xor \U$12693 ( \13676 , \13378 , \13380 );
xor \U$12694 ( \13677 , \13676 , \13383 );
and \U$12695 ( \13678 , \13674 , \13677 );
and \U$12696 ( \13679 , \13672 , \13677 );
or \U$12697 ( \13680 , \13675 , \13678 , \13679 );
and \U$12698 ( \13681 , \13661 , \13680 );
and \U$12699 ( \13682 , \13651 , \13680 );
or \U$12700 ( \13683 , \13662 , \13681 , \13682 );
xor \U$12701 ( \13684 , \13206 , \13362 );
xor \U$12702 ( \13685 , \13684 , \13373 );
xor \U$12703 ( \13686 , \13386 , \13388 );
xor \U$12704 ( \13687 , \13686 , \13391 );
and \U$12705 ( \13688 , \13685 , \13687 );
xor \U$12706 ( \13689 , \13397 , \13399 );
xor \U$12707 ( \13690 , \13689 , \13402 );
and \U$12708 ( \13691 , \13687 , \13690 );
and \U$12709 ( \13692 , \13685 , \13690 );
or \U$12710 ( \13693 , \13688 , \13691 , \13692 );
and \U$12711 ( \13694 , \13683 , \13693 );
xor \U$12712 ( \13695 , \13081 , \13091 );
xor \U$12713 ( \13696 , \13695 , \13094 );
and \U$12714 ( \13697 , \13693 , \13696 );
and \U$12715 ( \13698 , \13683 , \13696 );
or \U$12716 ( \13699 , \13694 , \13697 , \13698 );
xor \U$12717 ( \13700 , \12889 , \13049 );
xor \U$12718 ( \13701 , \13700 , \13068 );
xor \U$12719 ( \13702 , \13376 , \13394 );
xor \U$12720 ( \13703 , \13702 , \13405 );
and \U$12721 ( \13704 , \13701 , \13703 );
xor \U$12722 ( \13705 , \13410 , \13412 );
xor \U$12723 ( \13706 , \13705 , \13415 );
and \U$12724 ( \13707 , \13703 , \13706 );
and \U$12725 ( \13708 , \13701 , \13706 );
or \U$12726 ( \13709 , \13704 , \13707 , \13708 );
and \U$12727 ( \13710 , \13699 , \13709 );
xor \U$12728 ( \13711 , \13071 , \13097 );
xor \U$12729 ( \13712 , \13711 , \13108 );
and \U$12730 ( \13713 , \13709 , \13712 );
and \U$12731 ( \13714 , \13699 , \13712 );
or \U$12732 ( \13715 , \13710 , \13713 , \13714 );
xor \U$12733 ( \13716 , \13424 , \13426 );
xor \U$12734 ( \13717 , \13716 , \13429 );
and \U$12735 ( \13718 , \13715 , \13717 );
and \U$12736 ( \13719 , \13443 , \13718 );
xor \U$12737 ( \13720 , \13443 , \13718 );
xor \U$12738 ( \13721 , \13715 , \13717 );
and \U$12739 ( \13722 , \10829 , \1360 );
and \U$12740 ( \13723 , \10226 , \1358 );
nor \U$12741 ( \13724 , \13722 , \13723 );
xnor \U$12742 ( \13725 , \13724 , \1317 );
and \U$12743 ( \13726 , \11015 , \1247 );
and \U$12744 ( \13727 , \10834 , \1245 );
nor \U$12745 ( \13728 , \13726 , \13727 );
xnor \U$12746 ( \13729 , \13728 , \1198 );
and \U$12747 ( \13730 , \13725 , \13729 );
nand \U$12748 ( \13731 , \11635 , \1144 );
xnor \U$12749 ( \13732 , \13731 , \1105 );
and \U$12750 ( \13733 , \13729 , \13732 );
and \U$12751 ( \13734 , \13725 , \13732 );
or \U$12752 ( \13735 , \13730 , \13733 , \13734 );
and \U$12753 ( \13736 , \10834 , \1247 );
and \U$12754 ( \13737 , \10829 , \1245 );
nor \U$12755 ( \13738 , \13736 , \13737 );
xnor \U$12756 ( \13739 , \13738 , \1198 );
and \U$12757 ( \13740 , \13735 , \13739 );
and \U$12758 ( \13741 , \11635 , \1146 );
and \U$12759 ( \13742 , \11015 , \1144 );
nor \U$12760 ( \13743 , \13741 , \13742 );
xnor \U$12761 ( \13744 , \13743 , \1105 );
and \U$12762 ( \13745 , \13739 , \13744 );
and \U$12763 ( \13746 , \13735 , \13744 );
or \U$12764 ( \13747 , \13740 , \13745 , \13746 );
xor \U$12765 ( \13748 , \13499 , \13503 );
xor \U$12766 ( \13749 , \13748 , \13508 );
xor \U$12767 ( \13750 , \13515 , \13519 );
xor \U$12768 ( \13751 , \13750 , \13524 );
and \U$12769 ( \13752 , \13749 , \13751 );
xor \U$12770 ( \13753 , \13532 , \13536 );
xor \U$12771 ( \13754 , \13753 , \13541 );
and \U$12772 ( \13755 , \13751 , \13754 );
and \U$12773 ( \13756 , \13749 , \13754 );
or \U$12774 ( \13757 , \13752 , \13755 , \13756 );
and \U$12775 ( \13758 , \13747 , \13757 );
xor \U$12776 ( \13759 , \13447 , \13451 );
xor \U$12777 ( \13760 , \13759 , \13456 );
xor \U$12778 ( \13761 , \13463 , \13467 );
xor \U$12779 ( \13762 , \13761 , \13472 );
and \U$12780 ( \13763 , \13760 , \13762 );
xor \U$12781 ( \13764 , \13480 , \13484 );
xor \U$12782 ( \13765 , \13764 , \13489 );
and \U$12783 ( \13766 , \13762 , \13765 );
and \U$12784 ( \13767 , \13760 , \13765 );
or \U$12785 ( \13768 , \13763 , \13766 , \13767 );
and \U$12786 ( \13769 , \13757 , \13768 );
and \U$12787 ( \13770 , \13747 , \13768 );
or \U$12788 ( \13771 , \13758 , \13769 , \13770 );
and \U$12789 ( \13772 , \1457 , \10101 );
and \U$12790 ( \13773 , \1377 , \10099 );
nor \U$12791 ( \13774 , \13772 , \13773 );
xnor \U$12792 ( \13775 , \13774 , \9791 );
and \U$12793 ( \13776 , \1593 , \9564 );
and \U$12794 ( \13777 , \1531 , \9562 );
nor \U$12795 ( \13778 , \13776 , \13777 );
xnor \U$12796 ( \13779 , \13778 , \9193 );
and \U$12797 ( \13780 , \13775 , \13779 );
and \U$12798 ( \13781 , \1854 , \9002 );
and \U$12799 ( \13782 , \1656 , \9000 );
nor \U$12800 ( \13783 , \13781 , \13782 );
xnor \U$12801 ( \13784 , \13783 , \8684 );
and \U$12802 ( \13785 , \13779 , \13784 );
and \U$12803 ( \13786 , \13775 , \13784 );
or \U$12804 ( \13787 , \13780 , \13785 , \13786 );
and \U$12805 ( \13788 , \2047 , \8435 );
and \U$12806 ( \13789 , \1942 , \8433 );
nor \U$12807 ( \13790 , \13788 , \13789 );
xnor \U$12808 ( \13791 , \13790 , \8186 );
and \U$12809 ( \13792 , \2168 , \7906 );
and \U$12810 ( \13793 , \2052 , \7904 );
nor \U$12811 ( \13794 , \13792 , \13793 );
xnor \U$12812 ( \13795 , \13794 , \7646 );
and \U$12813 ( \13796 , \13791 , \13795 );
and \U$12814 ( \13797 , \2459 , \7412 );
and \U$12815 ( \13798 , \2283 , \7410 );
nor \U$12816 ( \13799 , \13797 , \13798 );
xnor \U$12817 ( \13800 , \13799 , \7097 );
and \U$12818 ( \13801 , \13795 , \13800 );
and \U$12819 ( \13802 , \13791 , \13800 );
or \U$12820 ( \13803 , \13796 , \13801 , \13802 );
and \U$12821 ( \13804 , \13787 , \13803 );
and \U$12822 ( \13805 , \1221 , \11482 );
and \U$12823 ( \13806 , \1167 , \11479 );
nor \U$12824 ( \13807 , \13805 , \13806 );
xnor \U$12825 ( \13808 , \13807 , \10427 );
and \U$12826 ( \13809 , \1349 , \10669 );
and \U$12827 ( \13810 , \1272 , \10667 );
nor \U$12828 ( \13811 , \13809 , \13810 );
xnor \U$12829 ( \13812 , \13811 , \10430 );
and \U$12830 ( \13813 , \13808 , \13812 );
and \U$12831 ( \13814 , \13812 , \1105 );
and \U$12832 ( \13815 , \13808 , \1105 );
or \U$12833 ( \13816 , \13813 , \13814 , \13815 );
and \U$12834 ( \13817 , \13803 , \13816 );
and \U$12835 ( \13818 , \13787 , \13816 );
or \U$12836 ( \13819 , \13804 , \13817 , \13818 );
and \U$12837 ( \13820 , \4679 , \4305 );
and \U$12838 ( \13821 , \4557 , \4303 );
nor \U$12839 ( \13822 , \13820 , \13821 );
xnor \U$12840 ( \13823 , \13822 , \4118 );
and \U$12841 ( \13824 , \4940 , \3992 );
and \U$12842 ( \13825 , \4684 , \3990 );
nor \U$12843 ( \13826 , \13824 , \13825 );
xnor \U$12844 ( \13827 , \13826 , \3787 );
and \U$12845 ( \13828 , \13823 , \13827 );
and \U$12846 ( \13829 , \5439 , \3586 );
and \U$12847 ( \13830 , \5137 , \3584 );
nor \U$12848 ( \13831 , \13829 , \13830 );
xnor \U$12849 ( \13832 , \13831 , \3437 );
and \U$12850 ( \13833 , \13827 , \13832 );
and \U$12851 ( \13834 , \13823 , \13832 );
or \U$12852 ( \13835 , \13828 , \13833 , \13834 );
and \U$12853 ( \13836 , \2710 , \6903 );
and \U$12854 ( \13837 , \2467 , \6901 );
nor \U$12855 ( \13838 , \13836 , \13837 );
xnor \U$12856 ( \13839 , \13838 , \6563 );
and \U$12857 ( \13840 , \2901 , \6314 );
and \U$12858 ( \13841 , \2715 , \6312 );
nor \U$12859 ( \13842 , \13840 , \13841 );
xnor \U$12860 ( \13843 , \13842 , \6073 );
and \U$12861 ( \13844 , \13839 , \13843 );
and \U$12862 ( \13845 , \3309 , \5848 );
and \U$12863 ( \13846 , \3045 , \5846 );
nor \U$12864 ( \13847 , \13845 , \13846 );
xnor \U$12865 ( \13848 , \13847 , \5660 );
and \U$12866 ( \13849 , \13843 , \13848 );
and \U$12867 ( \13850 , \13839 , \13848 );
or \U$12868 ( \13851 , \13844 , \13849 , \13850 );
and \U$12869 ( \13852 , \13835 , \13851 );
and \U$12870 ( \13853 , \3508 , \5474 );
and \U$12871 ( \13854 , \3334 , \5472 );
nor \U$12872 ( \13855 , \13853 , \13854 );
xnor \U$12873 ( \13856 , \13855 , \5242 );
and \U$12874 ( \13857 , \3813 , \5023 );
and \U$12875 ( \13858 , \3675 , \5021 );
nor \U$12876 ( \13859 , \13857 , \13858 );
xnor \U$12877 ( \13860 , \13859 , \4880 );
and \U$12878 ( \13861 , \13856 , \13860 );
and \U$12879 ( \13862 , \4349 , \4700 );
and \U$12880 ( \13863 , \3932 , \4698 );
nor \U$12881 ( \13864 , \13862 , \13863 );
xnor \U$12882 ( \13865 , \13864 , \4454 );
and \U$12883 ( \13866 , \13860 , \13865 );
and \U$12884 ( \13867 , \13856 , \13865 );
or \U$12885 ( \13868 , \13861 , \13866 , \13867 );
and \U$12886 ( \13869 , \13851 , \13868 );
and \U$12887 ( \13870 , \13835 , \13868 );
or \U$12888 ( \13871 , \13852 , \13869 , \13870 );
and \U$12889 ( \13872 , \13819 , \13871 );
and \U$12890 ( \13873 , \7168 , \2494 );
and \U$12891 ( \13874 , \6825 , \2492 );
nor \U$12892 ( \13875 , \13873 , \13874 );
xnor \U$12893 ( \13876 , \13875 , \2338 );
and \U$12894 ( \13877 , \7673 , \2222 );
and \U$12895 ( \13878 , \7370 , \2220 );
nor \U$12896 ( \13879 , \13877 , \13878 );
xnor \U$12897 ( \13880 , \13879 , \2109 );
and \U$12898 ( \13881 , \13876 , \13880 );
and \U$12899 ( \13882 , \8371 , \2028 );
and \U$12900 ( \13883 , \7845 , \2026 );
nor \U$12901 ( \13884 , \13882 , \13883 );
xnor \U$12902 ( \13885 , \13884 , \1892 );
and \U$12903 ( \13886 , \13880 , \13885 );
and \U$12904 ( \13887 , \13876 , \13885 );
or \U$12905 ( \13888 , \13881 , \13886 , \13887 );
and \U$12906 ( \13889 , \9041 , \1828 );
and \U$12907 ( \13890 , \8795 , \1826 );
nor \U$12908 ( \13891 , \13889 , \13890 );
xnor \U$12909 ( \13892 , \13891 , \1750 );
and \U$12910 ( \13893 , \9365 , \1664 );
and \U$12911 ( \13894 , \9046 , \1662 );
nor \U$12912 ( \13895 , \13893 , \13894 );
xnor \U$12913 ( \13896 , \13895 , \1570 );
and \U$12914 ( \13897 , \13892 , \13896 );
and \U$12915 ( \13898 , \10218 , \1494 );
and \U$12916 ( \13899 , \9649 , \1492 );
nor \U$12917 ( \13900 , \13898 , \13899 );
xnor \U$12918 ( \13901 , \13900 , \1422 );
and \U$12919 ( \13902 , \13896 , \13901 );
and \U$12920 ( \13903 , \13892 , \13901 );
or \U$12921 ( \13904 , \13897 , \13902 , \13903 );
and \U$12922 ( \13905 , \13888 , \13904 );
and \U$12923 ( \13906 , \5916 , \3264 );
and \U$12924 ( \13907 , \5447 , \3262 );
nor \U$12925 ( \13908 , \13906 , \13907 );
xnor \U$12926 ( \13909 , \13908 , \3122 );
and \U$12927 ( \13910 , \6185 , \2968 );
and \U$12928 ( \13911 , \5921 , \2966 );
nor \U$12929 ( \13912 , \13910 , \13911 );
xnor \U$12930 ( \13913 , \13912 , \2831 );
and \U$12931 ( \13914 , \13909 , \13913 );
and \U$12932 ( \13915 , \6816 , \2762 );
and \U$12933 ( \13916 , \6444 , \2760 );
nor \U$12934 ( \13917 , \13915 , \13916 );
xnor \U$12935 ( \13918 , \13917 , \2610 );
and \U$12936 ( \13919 , \13913 , \13918 );
and \U$12937 ( \13920 , \13909 , \13918 );
or \U$12938 ( \13921 , \13914 , \13919 , \13920 );
and \U$12939 ( \13922 , \13904 , \13921 );
and \U$12940 ( \13923 , \13888 , \13921 );
or \U$12941 ( \13924 , \13905 , \13922 , \13923 );
and \U$12942 ( \13925 , \13871 , \13924 );
and \U$12943 ( \13926 , \13819 , \13924 );
or \U$12944 ( \13927 , \13872 , \13925 , \13926 );
and \U$12945 ( \13928 , \13771 , \13927 );
xor \U$12946 ( \13929 , \13552 , \13556 );
xor \U$12947 ( \13930 , \13929 , \13561 );
xor \U$12948 ( \13931 , \13568 , \13572 );
xor \U$12949 ( \13932 , \13931 , \13577 );
and \U$12950 ( \13933 , \13930 , \13932 );
xor \U$12951 ( \13934 , \13585 , \13589 );
xor \U$12952 ( \13935 , \13934 , \13594 );
and \U$12953 ( \13936 , \13932 , \13935 );
and \U$12954 ( \13937 , \13930 , \13935 );
or \U$12955 ( \13938 , \13933 , \13936 , \13937 );
xor \U$12956 ( \13939 , \13226 , \13230 );
xor \U$12957 ( \13940 , \13939 , \1046 );
and \U$12958 ( \13941 , \13938 , \13940 );
xor \U$12959 ( \13942 , \13239 , \13243 );
xor \U$12960 ( \13943 , \13942 , \13248 );
and \U$12961 ( \13944 , \13940 , \13943 );
and \U$12962 ( \13945 , \13938 , \13943 );
or \U$12963 ( \13946 , \13941 , \13944 , \13945 );
and \U$12964 ( \13947 , \13927 , \13946 );
and \U$12965 ( \13948 , \13771 , \13946 );
or \U$12966 ( \13949 , \13928 , \13947 , \13948 );
xor \U$12967 ( \13950 , \13459 , \13475 );
xor \U$12968 ( \13951 , \13950 , \13492 );
xor \U$12969 ( \13952 , \13511 , \13527 );
xor \U$12970 ( \13953 , \13952 , \13544 );
and \U$12971 ( \13954 , \13951 , \13953 );
xor \U$12972 ( \13955 , \13564 , \13580 );
xor \U$12973 ( \13956 , \13955 , \13597 );
and \U$12974 ( \13957 , \13953 , \13956 );
and \U$12975 ( \13958 , \13951 , \13956 );
or \U$12976 ( \13959 , \13954 , \13957 , \13958 );
xor \U$12977 ( \13960 , \13605 , \13607 );
xor \U$12978 ( \13961 , \13960 , \13610 );
xor \U$12979 ( \13962 , \13615 , \13617 );
xor \U$12980 ( \13963 , \13962 , \13620 );
and \U$12981 ( \13964 , \13961 , \13963 );
xor \U$12982 ( \13965 , \13626 , \13628 );
xor \U$12983 ( \13966 , \13965 , \13631 );
and \U$12984 ( \13967 , \13963 , \13966 );
and \U$12985 ( \13968 , \13961 , \13966 );
or \U$12986 ( \13969 , \13964 , \13967 , \13968 );
and \U$12987 ( \13970 , \13959 , \13969 );
xor \U$12988 ( \13971 , \13270 , \13286 );
xor \U$12989 ( \13972 , \13971 , \13303 );
and \U$12990 ( \13973 , \13969 , \13972 );
and \U$12991 ( \13974 , \13959 , \13972 );
or \U$12992 ( \13975 , \13970 , \13973 , \13974 );
and \U$12993 ( \13976 , \13949 , \13975 );
xor \U$12994 ( \13977 , \13222 , \13234 );
xor \U$12995 ( \13978 , \13977 , \13251 );
xor \U$12996 ( \13979 , \13640 , \13642 );
xor \U$12997 ( \13980 , \13979 , \13645 );
and \U$12998 ( \13981 , \13978 , \13980 );
xor \U$12999 ( \13982 , \13664 , \13666 );
xor \U$13000 ( \13983 , \13982 , \13669 );
and \U$13001 ( \13984 , \13980 , \13983 );
and \U$13002 ( \13985 , \13978 , \13983 );
or \U$13003 ( \13986 , \13981 , \13984 , \13985 );
and \U$13004 ( \13987 , \13975 , \13986 );
and \U$13005 ( \13988 , \13949 , \13986 );
or \U$13006 ( \13989 , \13976 , \13987 , \13988 );
xor \U$13007 ( \13990 , \13603 , \13637 );
xor \U$13008 ( \13991 , \13990 , \13648 );
xor \U$13009 ( \13992 , \13653 , \13655 );
xor \U$13010 ( \13993 , \13992 , \13658 );
and \U$13011 ( \13994 , \13991 , \13993 );
xor \U$13012 ( \13995 , \13672 , \13674 );
xor \U$13013 ( \13996 , \13995 , \13677 );
and \U$13014 ( \13997 , \13993 , \13996 );
and \U$13015 ( \13998 , \13991 , \13996 );
or \U$13016 ( \13999 , \13994 , \13997 , \13998 );
and \U$13017 ( \14000 , \13989 , \13999 );
xor \U$13018 ( \14001 , \13685 , \13687 );
xor \U$13019 ( \14002 , \14001 , \13690 );
and \U$13020 ( \14003 , \13999 , \14002 );
and \U$13021 ( \14004 , \13989 , \14002 );
or \U$13022 ( \14005 , \14000 , \14003 , \14004 );
xor \U$13023 ( \14006 , \13683 , \13693 );
xor \U$13024 ( \14007 , \14006 , \13696 );
and \U$13025 ( \14008 , \14005 , \14007 );
xor \U$13026 ( \14009 , \13701 , \13703 );
xor \U$13027 ( \14010 , \14009 , \13706 );
and \U$13028 ( \14011 , \14007 , \14010 );
and \U$13029 ( \14012 , \14005 , \14010 );
or \U$13030 ( \14013 , \14008 , \14011 , \14012 );
xor \U$13031 ( \14014 , \13699 , \13709 );
xor \U$13032 ( \14015 , \14014 , \13712 );
and \U$13033 ( \14016 , \14013 , \14015 );
xor \U$13034 ( \14017 , \13408 , \13418 );
xor \U$13035 ( \14018 , \14017 , \13421 );
and \U$13036 ( \14019 , \14015 , \14018 );
and \U$13037 ( \14020 , \14013 , \14018 );
or \U$13038 ( \14021 , \14016 , \14019 , \14020 );
and \U$13039 ( \14022 , \13721 , \14021 );
xor \U$13040 ( \14023 , \13721 , \14021 );
xor \U$13041 ( \14024 , \14013 , \14015 );
xor \U$13042 ( \14025 , \14024 , \14018 );
xor \U$13043 ( \14026 , \13775 , \13779 );
xor \U$13044 ( \14027 , \14026 , \13784 );
xor \U$13045 ( \14028 , \13791 , \13795 );
xor \U$13046 ( \14029 , \14028 , \13800 );
and \U$13047 ( \14030 , \14027 , \14029 );
xor \U$13048 ( \14031 , \13839 , \13843 );
xor \U$13049 ( \14032 , \14031 , \13848 );
and \U$13050 ( \14033 , \14029 , \14032 );
and \U$13051 ( \14034 , \14027 , \14032 );
or \U$13052 ( \14035 , \14030 , \14033 , \14034 );
xor \U$13053 ( \14036 , \13823 , \13827 );
xor \U$13054 ( \14037 , \14036 , \13832 );
xor \U$13055 ( \14038 , \13856 , \13860 );
xor \U$13056 ( \14039 , \14038 , \13865 );
and \U$13057 ( \14040 , \14037 , \14039 );
xor \U$13058 ( \14041 , \13909 , \13913 );
xor \U$13059 ( \14042 , \14041 , \13918 );
and \U$13060 ( \14043 , \14039 , \14042 );
and \U$13061 ( \14044 , \14037 , \14042 );
or \U$13062 ( \14045 , \14040 , \14043 , \14044 );
and \U$13063 ( \14046 , \14035 , \14045 );
xor \U$13064 ( \14047 , \13876 , \13880 );
xor \U$13065 ( \14048 , \14047 , \13885 );
xor \U$13066 ( \14049 , \13725 , \13729 );
xor \U$13067 ( \14050 , \14049 , \13732 );
and \U$13068 ( \14051 , \14048 , \14050 );
xor \U$13069 ( \14052 , \13892 , \13896 );
xor \U$13070 ( \14053 , \14052 , \13901 );
and \U$13071 ( \14054 , \14050 , \14053 );
and \U$13072 ( \14055 , \14048 , \14053 );
or \U$13073 ( \14056 , \14051 , \14054 , \14055 );
and \U$13074 ( \14057 , \14045 , \14056 );
and \U$13075 ( \14058 , \14035 , \14056 );
or \U$13076 ( \14059 , \14046 , \14057 , \14058 );
and \U$13077 ( \14060 , \3045 , \6314 );
and \U$13078 ( \14061 , \2901 , \6312 );
nor \U$13079 ( \14062 , \14060 , \14061 );
xnor \U$13080 ( \14063 , \14062 , \6073 );
and \U$13081 ( \14064 , \3334 , \5848 );
and \U$13082 ( \14065 , \3309 , \5846 );
nor \U$13083 ( \14066 , \14064 , \14065 );
xnor \U$13084 ( \14067 , \14066 , \5660 );
and \U$13085 ( \14068 , \14063 , \14067 );
and \U$13086 ( \14069 , \3675 , \5474 );
and \U$13087 ( \14070 , \3508 , \5472 );
nor \U$13088 ( \14071 , \14069 , \14070 );
xnor \U$13089 ( \14072 , \14071 , \5242 );
and \U$13090 ( \14073 , \14067 , \14072 );
and \U$13091 ( \14074 , \14063 , \14072 );
or \U$13092 ( \14075 , \14068 , \14073 , \14074 );
and \U$13093 ( \14076 , \5137 , \3992 );
and \U$13094 ( \14077 , \4940 , \3990 );
nor \U$13095 ( \14078 , \14076 , \14077 );
xnor \U$13096 ( \14079 , \14078 , \3787 );
and \U$13097 ( \14080 , \5447 , \3586 );
and \U$13098 ( \14081 , \5439 , \3584 );
nor \U$13099 ( \14082 , \14080 , \14081 );
xnor \U$13100 ( \14083 , \14082 , \3437 );
and \U$13101 ( \14084 , \14079 , \14083 );
and \U$13102 ( \14085 , \5921 , \3264 );
and \U$13103 ( \14086 , \5916 , \3262 );
nor \U$13104 ( \14087 , \14085 , \14086 );
xnor \U$13105 ( \14088 , \14087 , \3122 );
and \U$13106 ( \14089 , \14083 , \14088 );
and \U$13107 ( \14090 , \14079 , \14088 );
or \U$13108 ( \14091 , \14084 , \14089 , \14090 );
and \U$13109 ( \14092 , \14075 , \14091 );
and \U$13110 ( \14093 , \3932 , \5023 );
and \U$13111 ( \14094 , \3813 , \5021 );
nor \U$13112 ( \14095 , \14093 , \14094 );
xnor \U$13113 ( \14096 , \14095 , \4880 );
and \U$13114 ( \14097 , \4557 , \4700 );
and \U$13115 ( \14098 , \4349 , \4698 );
nor \U$13116 ( \14099 , \14097 , \14098 );
xnor \U$13117 ( \14100 , \14099 , \4454 );
and \U$13118 ( \14101 , \14096 , \14100 );
and \U$13119 ( \14102 , \4684 , \4305 );
and \U$13120 ( \14103 , \4679 , \4303 );
nor \U$13121 ( \14104 , \14102 , \14103 );
xnor \U$13122 ( \14105 , \14104 , \4118 );
and \U$13123 ( \14106 , \14100 , \14105 );
and \U$13124 ( \14107 , \14096 , \14105 );
or \U$13125 ( \14108 , \14101 , \14106 , \14107 );
and \U$13126 ( \14109 , \14091 , \14108 );
and \U$13127 ( \14110 , \14075 , \14108 );
or \U$13128 ( \14111 , \14092 , \14109 , \14110 );
and \U$13129 ( \14112 , \9649 , \1664 );
and \U$13130 ( \14113 , \9365 , \1662 );
nor \U$13131 ( \14114 , \14112 , \14113 );
xnor \U$13132 ( \14115 , \14114 , \1570 );
and \U$13133 ( \14116 , \10226 , \1494 );
and \U$13134 ( \14117 , \10218 , \1492 );
nor \U$13135 ( \14118 , \14116 , \14117 );
xnor \U$13136 ( \14119 , \14118 , \1422 );
and \U$13137 ( \14120 , \14115 , \14119 );
and \U$13138 ( \14121 , \10834 , \1360 );
and \U$13139 ( \14122 , \10829 , \1358 );
nor \U$13140 ( \14123 , \14121 , \14122 );
xnor \U$13141 ( \14124 , \14123 , \1317 );
and \U$13142 ( \14125 , \14119 , \14124 );
and \U$13143 ( \14126 , \14115 , \14124 );
or \U$13144 ( \14127 , \14120 , \14125 , \14126 );
and \U$13145 ( \14128 , \7845 , \2222 );
and \U$13146 ( \14129 , \7673 , \2220 );
nor \U$13147 ( \14130 , \14128 , \14129 );
xnor \U$13148 ( \14131 , \14130 , \2109 );
and \U$13149 ( \14132 , \8795 , \2028 );
and \U$13150 ( \14133 , \8371 , \2026 );
nor \U$13151 ( \14134 , \14132 , \14133 );
xnor \U$13152 ( \14135 , \14134 , \1892 );
and \U$13153 ( \14136 , \14131 , \14135 );
and \U$13154 ( \14137 , \9046 , \1828 );
and \U$13155 ( \14138 , \9041 , \1826 );
nor \U$13156 ( \14139 , \14137 , \14138 );
xnor \U$13157 ( \14140 , \14139 , \1750 );
and \U$13158 ( \14141 , \14135 , \14140 );
and \U$13159 ( \14142 , \14131 , \14140 );
or \U$13160 ( \14143 , \14136 , \14141 , \14142 );
and \U$13161 ( \14144 , \14127 , \14143 );
and \U$13162 ( \14145 , \6444 , \2968 );
and \U$13163 ( \14146 , \6185 , \2966 );
nor \U$13164 ( \14147 , \14145 , \14146 );
xnor \U$13165 ( \14148 , \14147 , \2831 );
and \U$13166 ( \14149 , \6825 , \2762 );
and \U$13167 ( \14150 , \6816 , \2760 );
nor \U$13168 ( \14151 , \14149 , \14150 );
xnor \U$13169 ( \14152 , \14151 , \2610 );
and \U$13170 ( \14153 , \14148 , \14152 );
and \U$13171 ( \14154 , \7370 , \2494 );
and \U$13172 ( \14155 , \7168 , \2492 );
nor \U$13173 ( \14156 , \14154 , \14155 );
xnor \U$13174 ( \14157 , \14156 , \2338 );
and \U$13175 ( \14158 , \14152 , \14157 );
and \U$13176 ( \14159 , \14148 , \14157 );
or \U$13177 ( \14160 , \14153 , \14158 , \14159 );
and \U$13178 ( \14161 , \14143 , \14160 );
and \U$13179 ( \14162 , \14127 , \14160 );
or \U$13180 ( \14163 , \14144 , \14161 , \14162 );
and \U$13181 ( \14164 , \14111 , \14163 );
and \U$13182 ( \14165 , \2283 , \7906 );
and \U$13183 ( \14166 , \2168 , \7904 );
nor \U$13184 ( \14167 , \14165 , \14166 );
xnor \U$13185 ( \14168 , \14167 , \7646 );
and \U$13186 ( \14169 , \2467 , \7412 );
and \U$13187 ( \14170 , \2459 , \7410 );
nor \U$13188 ( \14171 , \14169 , \14170 );
xnor \U$13189 ( \14172 , \14171 , \7097 );
and \U$13190 ( \14173 , \14168 , \14172 );
and \U$13191 ( \14174 , \2715 , \6903 );
and \U$13192 ( \14175 , \2710 , \6901 );
nor \U$13193 ( \14176 , \14174 , \14175 );
xnor \U$13194 ( \14177 , \14176 , \6563 );
and \U$13195 ( \14178 , \14172 , \14177 );
and \U$13196 ( \14179 , \14168 , \14177 );
or \U$13197 ( \14180 , \14173 , \14178 , \14179 );
and \U$13198 ( \14181 , \1272 , \11482 );
and \U$13199 ( \14182 , \1221 , \11479 );
nor \U$13200 ( \14183 , \14181 , \14182 );
xnor \U$13201 ( \14184 , \14183 , \10427 );
and \U$13202 ( \14185 , \1377 , \10669 );
and \U$13203 ( \14186 , \1349 , \10667 );
nor \U$13204 ( \14187 , \14185 , \14186 );
xnor \U$13205 ( \14188 , \14187 , \10430 );
and \U$13206 ( \14189 , \14184 , \14188 );
and \U$13207 ( \14190 , \1531 , \10101 );
and \U$13208 ( \14191 , \1457 , \10099 );
nor \U$13209 ( \14192 , \14190 , \14191 );
xnor \U$13210 ( \14193 , \14192 , \9791 );
and \U$13211 ( \14194 , \14188 , \14193 );
and \U$13212 ( \14195 , \14184 , \14193 );
or \U$13213 ( \14196 , \14189 , \14194 , \14195 );
and \U$13214 ( \14197 , \14180 , \14196 );
and \U$13215 ( \14198 , \1656 , \9564 );
and \U$13216 ( \14199 , \1593 , \9562 );
nor \U$13217 ( \14200 , \14198 , \14199 );
xnor \U$13218 ( \14201 , \14200 , \9193 );
and \U$13219 ( \14202 , \1942 , \9002 );
and \U$13220 ( \14203 , \1854 , \9000 );
nor \U$13221 ( \14204 , \14202 , \14203 );
xnor \U$13222 ( \14205 , \14204 , \8684 );
and \U$13223 ( \14206 , \14201 , \14205 );
and \U$13224 ( \14207 , \2052 , \8435 );
and \U$13225 ( \14208 , \2047 , \8433 );
nor \U$13226 ( \14209 , \14207 , \14208 );
xnor \U$13227 ( \14210 , \14209 , \8186 );
and \U$13228 ( \14211 , \14205 , \14210 );
and \U$13229 ( \14212 , \14201 , \14210 );
or \U$13230 ( \14213 , \14206 , \14211 , \14212 );
and \U$13231 ( \14214 , \14196 , \14213 );
and \U$13232 ( \14215 , \14180 , \14213 );
or \U$13233 ( \14216 , \14197 , \14214 , \14215 );
and \U$13234 ( \14217 , \14163 , \14216 );
and \U$13235 ( \14218 , \14111 , \14216 );
or \U$13236 ( \14219 , \14164 , \14217 , \14218 );
and \U$13237 ( \14220 , \14059 , \14219 );
xor \U$13238 ( \14221 , \13749 , \13751 );
xor \U$13239 ( \14222 , \14221 , \13754 );
xor \U$13240 ( \14223 , \13930 , \13932 );
xor \U$13241 ( \14224 , \14223 , \13935 );
and \U$13242 ( \14225 , \14222 , \14224 );
xor \U$13243 ( \14226 , \13760 , \13762 );
xor \U$13244 ( \14227 , \14226 , \13765 );
and \U$13245 ( \14228 , \14224 , \14227 );
and \U$13246 ( \14229 , \14222 , \14227 );
or \U$13247 ( \14230 , \14225 , \14228 , \14229 );
and \U$13248 ( \14231 , \14219 , \14230 );
and \U$13249 ( \14232 , \14059 , \14230 );
or \U$13250 ( \14233 , \14220 , \14231 , \14232 );
xor \U$13251 ( \14234 , \13747 , \13757 );
xor \U$13252 ( \14235 , \14234 , \13768 );
xor \U$13253 ( \14236 , \13819 , \13871 );
xor \U$13254 ( \14237 , \14236 , \13924 );
and \U$13255 ( \14238 , \14235 , \14237 );
xor \U$13256 ( \14239 , \13938 , \13940 );
xor \U$13257 ( \14240 , \14239 , \13943 );
and \U$13258 ( \14241 , \14237 , \14240 );
and \U$13259 ( \14242 , \14235 , \14240 );
or \U$13260 ( \14243 , \14238 , \14241 , \14242 );
and \U$13261 ( \14244 , \14233 , \14243 );
xor \U$13262 ( \14245 , \13735 , \13739 );
xor \U$13263 ( \14246 , \14245 , \13744 );
xor \U$13264 ( \14247 , \13835 , \13851 );
xor \U$13265 ( \14248 , \14247 , \13868 );
and \U$13266 ( \14249 , \14246 , \14248 );
xor \U$13267 ( \14250 , \13888 , \13904 );
xor \U$13268 ( \14251 , \14250 , \13921 );
and \U$13269 ( \14252 , \14248 , \14251 );
and \U$13270 ( \14253 , \14246 , \14251 );
or \U$13271 ( \14254 , \14249 , \14252 , \14253 );
xor \U$13272 ( \14255 , \13951 , \13953 );
xor \U$13273 ( \14256 , \14255 , \13956 );
and \U$13274 ( \14257 , \14254 , \14256 );
xor \U$13275 ( \14258 , \13961 , \13963 );
xor \U$13276 ( \14259 , \14258 , \13966 );
and \U$13277 ( \14260 , \14256 , \14259 );
and \U$13278 ( \14261 , \14254 , \14259 );
or \U$13279 ( \14262 , \14257 , \14260 , \14261 );
and \U$13280 ( \14263 , \14243 , \14262 );
and \U$13281 ( \14264 , \14233 , \14262 );
or \U$13282 ( \14265 , \14244 , \14263 , \14264 );
xor \U$13283 ( \14266 , \13495 , \13547 );
xor \U$13284 ( \14267 , \14266 , \13600 );
xor \U$13285 ( \14268 , \13613 , \13623 );
xor \U$13286 ( \14269 , \14268 , \13634 );
and \U$13287 ( \14270 , \14267 , \14269 );
xor \U$13288 ( \14271 , \13978 , \13980 );
xor \U$13289 ( \14272 , \14271 , \13983 );
and \U$13290 ( \14273 , \14269 , \14272 );
and \U$13291 ( \14274 , \14267 , \14272 );
or \U$13292 ( \14275 , \14270 , \14273 , \14274 );
and \U$13293 ( \14276 , \14265 , \14275 );
xor \U$13294 ( \14277 , \13991 , \13993 );
xor \U$13295 ( \14278 , \14277 , \13996 );
and \U$13296 ( \14279 , \14275 , \14278 );
and \U$13297 ( \14280 , \14265 , \14278 );
or \U$13298 ( \14281 , \14276 , \14279 , \14280 );
xor \U$13299 ( \14282 , \13651 , \13661 );
xor \U$13300 ( \14283 , \14282 , \13680 );
and \U$13301 ( \14284 , \14281 , \14283 );
xor \U$13302 ( \14285 , \13989 , \13999 );
xor \U$13303 ( \14286 , \14285 , \14002 );
and \U$13304 ( \14287 , \14283 , \14286 );
and \U$13305 ( \14288 , \14281 , \14286 );
or \U$13306 ( \14289 , \14284 , \14287 , \14288 );
xor \U$13307 ( \14290 , \14005 , \14007 );
xor \U$13308 ( \14291 , \14290 , \14010 );
and \U$13309 ( \14292 , \14289 , \14291 );
and \U$13310 ( \14293 , \14025 , \14292 );
xor \U$13311 ( \14294 , \14025 , \14292 );
xor \U$13312 ( \14295 , \14289 , \14291 );
xor \U$13313 ( \14296 , \14079 , \14083 );
xor \U$13314 ( \14297 , \14296 , \14088 );
xor \U$13315 ( \14298 , \14096 , \14100 );
xor \U$13316 ( \14299 , \14298 , \14105 );
and \U$13317 ( \14300 , \14297 , \14299 );
xor \U$13318 ( \14301 , \14148 , \14152 );
xor \U$13319 ( \14302 , \14301 , \14157 );
and \U$13320 ( \14303 , \14299 , \14302 );
and \U$13321 ( \14304 , \14297 , \14302 );
or \U$13322 ( \14305 , \14300 , \14303 , \14304 );
xor \U$13323 ( \14306 , \14063 , \14067 );
xor \U$13324 ( \14307 , \14306 , \14072 );
xor \U$13325 ( \14308 , \14168 , \14172 );
xor \U$13326 ( \14309 , \14308 , \14177 );
and \U$13327 ( \14310 , \14307 , \14309 );
xor \U$13328 ( \14311 , \14201 , \14205 );
xor \U$13329 ( \14312 , \14311 , \14210 );
and \U$13330 ( \14313 , \14309 , \14312 );
and \U$13331 ( \14314 , \14307 , \14312 );
or \U$13332 ( \14315 , \14310 , \14313 , \14314 );
and \U$13333 ( \14316 , \14305 , \14315 );
and \U$13334 ( \14317 , \11635 , \1247 );
and \U$13335 ( \14318 , \11015 , \1245 );
nor \U$13336 ( \14319 , \14317 , \14318 );
xnor \U$13337 ( \14320 , \14319 , \1198 );
xor \U$13338 ( \14321 , \14115 , \14119 );
xor \U$13339 ( \14322 , \14321 , \14124 );
and \U$13340 ( \14323 , \14320 , \14322 );
xor \U$13341 ( \14324 , \14131 , \14135 );
xor \U$13342 ( \14325 , \14324 , \14140 );
and \U$13343 ( \14326 , \14322 , \14325 );
and \U$13344 ( \14327 , \14320 , \14325 );
or \U$13345 ( \14328 , \14323 , \14326 , \14327 );
and \U$13346 ( \14329 , \14315 , \14328 );
and \U$13347 ( \14330 , \14305 , \14328 );
or \U$13348 ( \14331 , \14316 , \14329 , \14330 );
and \U$13349 ( \14332 , \2168 , \8435 );
and \U$13350 ( \14333 , \2052 , \8433 );
nor \U$13351 ( \14334 , \14332 , \14333 );
xnor \U$13352 ( \14335 , \14334 , \8186 );
and \U$13353 ( \14336 , \2459 , \7906 );
and \U$13354 ( \14337 , \2283 , \7904 );
nor \U$13355 ( \14338 , \14336 , \14337 );
xnor \U$13356 ( \14339 , \14338 , \7646 );
and \U$13357 ( \14340 , \14335 , \14339 );
and \U$13358 ( \14341 , \2710 , \7412 );
and \U$13359 ( \14342 , \2467 , \7410 );
nor \U$13360 ( \14343 , \14341 , \14342 );
xnor \U$13361 ( \14344 , \14343 , \7097 );
and \U$13362 ( \14345 , \14339 , \14344 );
and \U$13363 ( \14346 , \14335 , \14344 );
or \U$13364 ( \14347 , \14340 , \14345 , \14346 );
and \U$13365 ( \14348 , \1593 , \10101 );
and \U$13366 ( \14349 , \1531 , \10099 );
nor \U$13367 ( \14350 , \14348 , \14349 );
xnor \U$13368 ( \14351 , \14350 , \9791 );
and \U$13369 ( \14352 , \1854 , \9564 );
and \U$13370 ( \14353 , \1656 , \9562 );
nor \U$13371 ( \14354 , \14352 , \14353 );
xnor \U$13372 ( \14355 , \14354 , \9193 );
and \U$13373 ( \14356 , \14351 , \14355 );
and \U$13374 ( \14357 , \2047 , \9002 );
and \U$13375 ( \14358 , \1942 , \9000 );
nor \U$13376 ( \14359 , \14357 , \14358 );
xnor \U$13377 ( \14360 , \14359 , \8684 );
and \U$13378 ( \14361 , \14355 , \14360 );
and \U$13379 ( \14362 , \14351 , \14360 );
or \U$13380 ( \14363 , \14356 , \14361 , \14362 );
and \U$13381 ( \14364 , \14347 , \14363 );
and \U$13382 ( \14365 , \1349 , \11482 );
and \U$13383 ( \14366 , \1272 , \11479 );
nor \U$13384 ( \14367 , \14365 , \14366 );
xnor \U$13385 ( \14368 , \14367 , \10427 );
and \U$13386 ( \14369 , \1457 , \10669 );
and \U$13387 ( \14370 , \1377 , \10667 );
nor \U$13388 ( \14371 , \14369 , \14370 );
xnor \U$13389 ( \14372 , \14371 , \10430 );
and \U$13390 ( \14373 , \14368 , \14372 );
and \U$13391 ( \14374 , \14372 , \1198 );
and \U$13392 ( \14375 , \14368 , \1198 );
or \U$13393 ( \14376 , \14373 , \14374 , \14375 );
and \U$13394 ( \14377 , \14363 , \14376 );
and \U$13395 ( \14378 , \14347 , \14376 );
or \U$13396 ( \14379 , \14364 , \14377 , \14378 );
and \U$13397 ( \14380 , \9365 , \1828 );
and \U$13398 ( \14381 , \9046 , \1826 );
nor \U$13399 ( \14382 , \14380 , \14381 );
xnor \U$13400 ( \14383 , \14382 , \1750 );
and \U$13401 ( \14384 , \10218 , \1664 );
and \U$13402 ( \14385 , \9649 , \1662 );
nor \U$13403 ( \14386 , \14384 , \14385 );
xnor \U$13404 ( \14387 , \14386 , \1570 );
and \U$13405 ( \14388 , \14383 , \14387 );
and \U$13406 ( \14389 , \10829 , \1494 );
and \U$13407 ( \14390 , \10226 , \1492 );
nor \U$13408 ( \14391 , \14389 , \14390 );
xnor \U$13409 ( \14392 , \14391 , \1422 );
and \U$13410 ( \14393 , \14387 , \14392 );
and \U$13411 ( \14394 , \14383 , \14392 );
or \U$13412 ( \14395 , \14388 , \14393 , \14394 );
and \U$13413 ( \14396 , \6185 , \3264 );
and \U$13414 ( \14397 , \5921 , \3262 );
nor \U$13415 ( \14398 , \14396 , \14397 );
xnor \U$13416 ( \14399 , \14398 , \3122 );
and \U$13417 ( \14400 , \6816 , \2968 );
and \U$13418 ( \14401 , \6444 , \2966 );
nor \U$13419 ( \14402 , \14400 , \14401 );
xnor \U$13420 ( \14403 , \14402 , \2831 );
and \U$13421 ( \14404 , \14399 , \14403 );
and \U$13422 ( \14405 , \7168 , \2762 );
and \U$13423 ( \14406 , \6825 , \2760 );
nor \U$13424 ( \14407 , \14405 , \14406 );
xnor \U$13425 ( \14408 , \14407 , \2610 );
and \U$13426 ( \14409 , \14403 , \14408 );
and \U$13427 ( \14410 , \14399 , \14408 );
or \U$13428 ( \14411 , \14404 , \14409 , \14410 );
and \U$13429 ( \14412 , \14395 , \14411 );
and \U$13430 ( \14413 , \7673 , \2494 );
and \U$13431 ( \14414 , \7370 , \2492 );
nor \U$13432 ( \14415 , \14413 , \14414 );
xnor \U$13433 ( \14416 , \14415 , \2338 );
and \U$13434 ( \14417 , \8371 , \2222 );
and \U$13435 ( \14418 , \7845 , \2220 );
nor \U$13436 ( \14419 , \14417 , \14418 );
xnor \U$13437 ( \14420 , \14419 , \2109 );
and \U$13438 ( \14421 , \14416 , \14420 );
and \U$13439 ( \14422 , \9041 , \2028 );
and \U$13440 ( \14423 , \8795 , \2026 );
nor \U$13441 ( \14424 , \14422 , \14423 );
xnor \U$13442 ( \14425 , \14424 , \1892 );
and \U$13443 ( \14426 , \14420 , \14425 );
and \U$13444 ( \14427 , \14416 , \14425 );
or \U$13445 ( \14428 , \14421 , \14426 , \14427 );
and \U$13446 ( \14429 , \14411 , \14428 );
and \U$13447 ( \14430 , \14395 , \14428 );
or \U$13448 ( \14431 , \14412 , \14429 , \14430 );
and \U$13449 ( \14432 , \14379 , \14431 );
and \U$13450 ( \14433 , \4940 , \4305 );
and \U$13451 ( \14434 , \4684 , \4303 );
nor \U$13452 ( \14435 , \14433 , \14434 );
xnor \U$13453 ( \14436 , \14435 , \4118 );
and \U$13454 ( \14437 , \5439 , \3992 );
and \U$13455 ( \14438 , \5137 , \3990 );
nor \U$13456 ( \14439 , \14437 , \14438 );
xnor \U$13457 ( \14440 , \14439 , \3787 );
and \U$13458 ( \14441 , \14436 , \14440 );
and \U$13459 ( \14442 , \5916 , \3586 );
and \U$13460 ( \14443 , \5447 , \3584 );
nor \U$13461 ( \14444 , \14442 , \14443 );
xnor \U$13462 ( \14445 , \14444 , \3437 );
and \U$13463 ( \14446 , \14440 , \14445 );
and \U$13464 ( \14447 , \14436 , \14445 );
or \U$13465 ( \14448 , \14441 , \14446 , \14447 );
and \U$13466 ( \14449 , \3813 , \5474 );
and \U$13467 ( \14450 , \3675 , \5472 );
nor \U$13468 ( \14451 , \14449 , \14450 );
xnor \U$13469 ( \14452 , \14451 , \5242 );
and \U$13470 ( \14453 , \4349 , \5023 );
and \U$13471 ( \14454 , \3932 , \5021 );
nor \U$13472 ( \14455 , \14453 , \14454 );
xnor \U$13473 ( \14456 , \14455 , \4880 );
and \U$13474 ( \14457 , \14452 , \14456 );
and \U$13475 ( \14458 , \4679 , \4700 );
and \U$13476 ( \14459 , \4557 , \4698 );
nor \U$13477 ( \14460 , \14458 , \14459 );
xnor \U$13478 ( \14461 , \14460 , \4454 );
and \U$13479 ( \14462 , \14456 , \14461 );
and \U$13480 ( \14463 , \14452 , \14461 );
or \U$13481 ( \14464 , \14457 , \14462 , \14463 );
and \U$13482 ( \14465 , \14448 , \14464 );
and \U$13483 ( \14466 , \2901 , \6903 );
and \U$13484 ( \14467 , \2715 , \6901 );
nor \U$13485 ( \14468 , \14466 , \14467 );
xnor \U$13486 ( \14469 , \14468 , \6563 );
and \U$13487 ( \14470 , \3309 , \6314 );
and \U$13488 ( \14471 , \3045 , \6312 );
nor \U$13489 ( \14472 , \14470 , \14471 );
xnor \U$13490 ( \14473 , \14472 , \6073 );
and \U$13491 ( \14474 , \14469 , \14473 );
and \U$13492 ( \14475 , \3508 , \5848 );
and \U$13493 ( \14476 , \3334 , \5846 );
nor \U$13494 ( \14477 , \14475 , \14476 );
xnor \U$13495 ( \14478 , \14477 , \5660 );
and \U$13496 ( \14479 , \14473 , \14478 );
and \U$13497 ( \14480 , \14469 , \14478 );
or \U$13498 ( \14481 , \14474 , \14479 , \14480 );
and \U$13499 ( \14482 , \14464 , \14481 );
and \U$13500 ( \14483 , \14448 , \14481 );
or \U$13501 ( \14484 , \14465 , \14482 , \14483 );
and \U$13502 ( \14485 , \14431 , \14484 );
and \U$13503 ( \14486 , \14379 , \14484 );
or \U$13504 ( \14487 , \14432 , \14485 , \14486 );
and \U$13505 ( \14488 , \14331 , \14487 );
xor \U$13506 ( \14489 , \13808 , \13812 );
xor \U$13507 ( \14490 , \14489 , \1105 );
xor \U$13508 ( \14491 , \14027 , \14029 );
xor \U$13509 ( \14492 , \14491 , \14032 );
and \U$13510 ( \14493 , \14490 , \14492 );
xor \U$13511 ( \14494 , \14037 , \14039 );
xor \U$13512 ( \14495 , \14494 , \14042 );
and \U$13513 ( \14496 , \14492 , \14495 );
and \U$13514 ( \14497 , \14490 , \14495 );
or \U$13515 ( \14498 , \14493 , \14496 , \14497 );
and \U$13516 ( \14499 , \14487 , \14498 );
and \U$13517 ( \14500 , \14331 , \14498 );
or \U$13518 ( \14501 , \14488 , \14499 , \14500 );
xor \U$13519 ( \14502 , \14075 , \14091 );
xor \U$13520 ( \14503 , \14502 , \14108 );
xor \U$13521 ( \14504 , \14127 , \14143 );
xor \U$13522 ( \14505 , \14504 , \14160 );
and \U$13523 ( \14506 , \14503 , \14505 );
xor \U$13524 ( \14507 , \14048 , \14050 );
xor \U$13525 ( \14508 , \14507 , \14053 );
and \U$13526 ( \14509 , \14505 , \14508 );
and \U$13527 ( \14510 , \14503 , \14508 );
or \U$13528 ( \14511 , \14506 , \14509 , \14510 );
xor \U$13529 ( \14512 , \13787 , \13803 );
xor \U$13530 ( \14513 , \14512 , \13816 );
and \U$13531 ( \14514 , \14511 , \14513 );
xor \U$13532 ( \14515 , \14246 , \14248 );
xor \U$13533 ( \14516 , \14515 , \14251 );
and \U$13534 ( \14517 , \14513 , \14516 );
and \U$13535 ( \14518 , \14511 , \14516 );
or \U$13536 ( \14519 , \14514 , \14517 , \14518 );
and \U$13537 ( \14520 , \14501 , \14519 );
xor \U$13538 ( \14521 , \14035 , \14045 );
xor \U$13539 ( \14522 , \14521 , \14056 );
xor \U$13540 ( \14523 , \14111 , \14163 );
xor \U$13541 ( \14524 , \14523 , \14216 );
and \U$13542 ( \14525 , \14522 , \14524 );
xor \U$13543 ( \14526 , \14222 , \14224 );
xor \U$13544 ( \14527 , \14526 , \14227 );
and \U$13545 ( \14528 , \14524 , \14527 );
and \U$13546 ( \14529 , \14522 , \14527 );
or \U$13547 ( \14530 , \14525 , \14528 , \14529 );
and \U$13548 ( \14531 , \14519 , \14530 );
and \U$13549 ( \14532 , \14501 , \14530 );
or \U$13550 ( \14533 , \14520 , \14531 , \14532 );
xor \U$13551 ( \14534 , \14059 , \14219 );
xor \U$13552 ( \14535 , \14534 , \14230 );
xor \U$13553 ( \14536 , \14235 , \14237 );
xor \U$13554 ( \14537 , \14536 , \14240 );
and \U$13555 ( \14538 , \14535 , \14537 );
xor \U$13556 ( \14539 , \14254 , \14256 );
xor \U$13557 ( \14540 , \14539 , \14259 );
and \U$13558 ( \14541 , \14537 , \14540 );
and \U$13559 ( \14542 , \14535 , \14540 );
or \U$13560 ( \14543 , \14538 , \14541 , \14542 );
and \U$13561 ( \14544 , \14533 , \14543 );
xor \U$13562 ( \14545 , \13959 , \13969 );
xor \U$13563 ( \14546 , \14545 , \13972 );
and \U$13564 ( \14547 , \14543 , \14546 );
and \U$13565 ( \14548 , \14533 , \14546 );
or \U$13566 ( \14549 , \14544 , \14547 , \14548 );
xor \U$13567 ( \14550 , \13771 , \13927 );
xor \U$13568 ( \14551 , \14550 , \13946 );
xor \U$13569 ( \14552 , \14233 , \14243 );
xor \U$13570 ( \14553 , \14552 , \14262 );
and \U$13571 ( \14554 , \14551 , \14553 );
xor \U$13572 ( \14555 , \14267 , \14269 );
xor \U$13573 ( \14556 , \14555 , \14272 );
and \U$13574 ( \14557 , \14553 , \14556 );
and \U$13575 ( \14558 , \14551 , \14556 );
or \U$13576 ( \14559 , \14554 , \14557 , \14558 );
and \U$13577 ( \14560 , \14549 , \14559 );
xor \U$13578 ( \14561 , \13949 , \13975 );
xor \U$13579 ( \14562 , \14561 , \13986 );
and \U$13580 ( \14563 , \14559 , \14562 );
and \U$13581 ( \14564 , \14549 , \14562 );
or \U$13582 ( \14565 , \14560 , \14563 , \14564 );
xor \U$13583 ( \14566 , \14281 , \14283 );
xor \U$13584 ( \14567 , \14566 , \14286 );
and \U$13585 ( \14568 , \14565 , \14567 );
and \U$13586 ( \14569 , \14295 , \14568 );
xor \U$13587 ( \14570 , \14295 , \14568 );
xor \U$13588 ( \14571 , \14565 , \14567 );
xor \U$13589 ( \14572 , \14436 , \14440 );
xor \U$13590 ( \14573 , \14572 , \14445 );
xor \U$13591 ( \14574 , \14399 , \14403 );
xor \U$13592 ( \14575 , \14574 , \14408 );
and \U$13593 ( \14576 , \14573 , \14575 );
xor \U$13594 ( \14577 , \14416 , \14420 );
xor \U$13595 ( \14578 , \14577 , \14425 );
and \U$13596 ( \14579 , \14575 , \14578 );
and \U$13597 ( \14580 , \14573 , \14578 );
or \U$13598 ( \14581 , \14576 , \14579 , \14580 );
and \U$13599 ( \14582 , \11015 , \1360 );
and \U$13600 ( \14583 , \10834 , \1358 );
nor \U$13601 ( \14584 , \14582 , \14583 );
xnor \U$13602 ( \14585 , \14584 , \1317 );
nand \U$13603 ( \14586 , \11635 , \1245 );
xnor \U$13604 ( \14587 , \14586 , \1198 );
and \U$13605 ( \14588 , \14585 , \14587 );
xor \U$13606 ( \14589 , \14383 , \14387 );
xor \U$13607 ( \14590 , \14589 , \14392 );
and \U$13608 ( \14591 , \14587 , \14590 );
and \U$13609 ( \14592 , \14585 , \14590 );
or \U$13610 ( \14593 , \14588 , \14591 , \14592 );
and \U$13611 ( \14594 , \14581 , \14593 );
xor \U$13612 ( \14595 , \14335 , \14339 );
xor \U$13613 ( \14596 , \14595 , \14344 );
xor \U$13614 ( \14597 , \14452 , \14456 );
xor \U$13615 ( \14598 , \14597 , \14461 );
and \U$13616 ( \14599 , \14596 , \14598 );
xor \U$13617 ( \14600 , \14469 , \14473 );
xor \U$13618 ( \14601 , \14600 , \14478 );
and \U$13619 ( \14602 , \14598 , \14601 );
and \U$13620 ( \14603 , \14596 , \14601 );
or \U$13621 ( \14604 , \14599 , \14602 , \14603 );
and \U$13622 ( \14605 , \14593 , \14604 );
and \U$13623 ( \14606 , \14581 , \14604 );
or \U$13624 ( \14607 , \14594 , \14605 , \14606 );
and \U$13625 ( \14608 , \10226 , \1664 );
and \U$13626 ( \14609 , \10218 , \1662 );
nor \U$13627 ( \14610 , \14608 , \14609 );
xnor \U$13628 ( \14611 , \14610 , \1570 );
and \U$13629 ( \14612 , \10834 , \1494 );
and \U$13630 ( \14613 , \10829 , \1492 );
nor \U$13631 ( \14614 , \14612 , \14613 );
xnor \U$13632 ( \14615 , \14614 , \1422 );
and \U$13633 ( \14616 , \14611 , \14615 );
and \U$13634 ( \14617 , \11635 , \1360 );
and \U$13635 ( \14618 , \11015 , \1358 );
nor \U$13636 ( \14619 , \14617 , \14618 );
xnor \U$13637 ( \14620 , \14619 , \1317 );
and \U$13638 ( \14621 , \14615 , \14620 );
and \U$13639 ( \14622 , \14611 , \14620 );
or \U$13640 ( \14623 , \14616 , \14621 , \14622 );
and \U$13641 ( \14624 , \6825 , \2968 );
and \U$13642 ( \14625 , \6816 , \2966 );
nor \U$13643 ( \14626 , \14624 , \14625 );
xnor \U$13644 ( \14627 , \14626 , \2831 );
and \U$13645 ( \14628 , \7370 , \2762 );
and \U$13646 ( \14629 , \7168 , \2760 );
nor \U$13647 ( \14630 , \14628 , \14629 );
xnor \U$13648 ( \14631 , \14630 , \2610 );
and \U$13649 ( \14632 , \14627 , \14631 );
and \U$13650 ( \14633 , \7845 , \2494 );
and \U$13651 ( \14634 , \7673 , \2492 );
nor \U$13652 ( \14635 , \14633 , \14634 );
xnor \U$13653 ( \14636 , \14635 , \2338 );
and \U$13654 ( \14637 , \14631 , \14636 );
and \U$13655 ( \14638 , \14627 , \14636 );
or \U$13656 ( \14639 , \14632 , \14637 , \14638 );
and \U$13657 ( \14640 , \14623 , \14639 );
and \U$13658 ( \14641 , \8795 , \2222 );
and \U$13659 ( \14642 , \8371 , \2220 );
nor \U$13660 ( \14643 , \14641 , \14642 );
xnor \U$13661 ( \14644 , \14643 , \2109 );
and \U$13662 ( \14645 , \9046 , \2028 );
and \U$13663 ( \14646 , \9041 , \2026 );
nor \U$13664 ( \14647 , \14645 , \14646 );
xnor \U$13665 ( \14648 , \14647 , \1892 );
and \U$13666 ( \14649 , \14644 , \14648 );
and \U$13667 ( \14650 , \9649 , \1828 );
and \U$13668 ( \14651 , \9365 , \1826 );
nor \U$13669 ( \14652 , \14650 , \14651 );
xnor \U$13670 ( \14653 , \14652 , \1750 );
and \U$13671 ( \14654 , \14648 , \14653 );
and \U$13672 ( \14655 , \14644 , \14653 );
or \U$13673 ( \14656 , \14649 , \14654 , \14655 );
and \U$13674 ( \14657 , \14639 , \14656 );
and \U$13675 ( \14658 , \14623 , \14656 );
or \U$13676 ( \14659 , \14640 , \14657 , \14658 );
and \U$13677 ( \14660 , \1942 , \9564 );
and \U$13678 ( \14661 , \1854 , \9562 );
nor \U$13679 ( \14662 , \14660 , \14661 );
xnor \U$13680 ( \14663 , \14662 , \9193 );
and \U$13681 ( \14664 , \2052 , \9002 );
and \U$13682 ( \14665 , \2047 , \9000 );
nor \U$13683 ( \14666 , \14664 , \14665 );
xnor \U$13684 ( \14667 , \14666 , \8684 );
and \U$13685 ( \14668 , \14663 , \14667 );
and \U$13686 ( \14669 , \2283 , \8435 );
and \U$13687 ( \14670 , \2168 , \8433 );
nor \U$13688 ( \14671 , \14669 , \14670 );
xnor \U$13689 ( \14672 , \14671 , \8186 );
and \U$13690 ( \14673 , \14667 , \14672 );
and \U$13691 ( \14674 , \14663 , \14672 );
or \U$13692 ( \14675 , \14668 , \14673 , \14674 );
and \U$13693 ( \14676 , \2467 , \7906 );
and \U$13694 ( \14677 , \2459 , \7904 );
nor \U$13695 ( \14678 , \14676 , \14677 );
xnor \U$13696 ( \14679 , \14678 , \7646 );
and \U$13697 ( \14680 , \2715 , \7412 );
and \U$13698 ( \14681 , \2710 , \7410 );
nor \U$13699 ( \14682 , \14680 , \14681 );
xnor \U$13700 ( \14683 , \14682 , \7097 );
and \U$13701 ( \14684 , \14679 , \14683 );
and \U$13702 ( \14685 , \3045 , \6903 );
and \U$13703 ( \14686 , \2901 , \6901 );
nor \U$13704 ( \14687 , \14685 , \14686 );
xnor \U$13705 ( \14688 , \14687 , \6563 );
and \U$13706 ( \14689 , \14683 , \14688 );
and \U$13707 ( \14690 , \14679 , \14688 );
or \U$13708 ( \14691 , \14684 , \14689 , \14690 );
and \U$13709 ( \14692 , \14675 , \14691 );
and \U$13710 ( \14693 , \1377 , \11482 );
and \U$13711 ( \14694 , \1349 , \11479 );
nor \U$13712 ( \14695 , \14693 , \14694 );
xnor \U$13713 ( \14696 , \14695 , \10427 );
and \U$13714 ( \14697 , \1531 , \10669 );
and \U$13715 ( \14698 , \1457 , \10667 );
nor \U$13716 ( \14699 , \14697 , \14698 );
xnor \U$13717 ( \14700 , \14699 , \10430 );
and \U$13718 ( \14701 , \14696 , \14700 );
and \U$13719 ( \14702 , \1656 , \10101 );
and \U$13720 ( \14703 , \1593 , \10099 );
nor \U$13721 ( \14704 , \14702 , \14703 );
xnor \U$13722 ( \14705 , \14704 , \9791 );
and \U$13723 ( \14706 , \14700 , \14705 );
and \U$13724 ( \14707 , \14696 , \14705 );
or \U$13725 ( \14708 , \14701 , \14706 , \14707 );
and \U$13726 ( \14709 , \14691 , \14708 );
and \U$13727 ( \14710 , \14675 , \14708 );
or \U$13728 ( \14711 , \14692 , \14709 , \14710 );
and \U$13729 ( \14712 , \14659 , \14711 );
and \U$13730 ( \14713 , \5447 , \3992 );
and \U$13731 ( \14714 , \5439 , \3990 );
nor \U$13732 ( \14715 , \14713 , \14714 );
xnor \U$13733 ( \14716 , \14715 , \3787 );
and \U$13734 ( \14717 , \5921 , \3586 );
and \U$13735 ( \14718 , \5916 , \3584 );
nor \U$13736 ( \14719 , \14717 , \14718 );
xnor \U$13737 ( \14720 , \14719 , \3437 );
and \U$13738 ( \14721 , \14716 , \14720 );
and \U$13739 ( \14722 , \6444 , \3264 );
and \U$13740 ( \14723 , \6185 , \3262 );
nor \U$13741 ( \14724 , \14722 , \14723 );
xnor \U$13742 ( \14725 , \14724 , \3122 );
and \U$13743 ( \14726 , \14720 , \14725 );
and \U$13744 ( \14727 , \14716 , \14725 );
or \U$13745 ( \14728 , \14721 , \14726 , \14727 );
and \U$13746 ( \14729 , \4557 , \5023 );
and \U$13747 ( \14730 , \4349 , \5021 );
nor \U$13748 ( \14731 , \14729 , \14730 );
xnor \U$13749 ( \14732 , \14731 , \4880 );
and \U$13750 ( \14733 , \4684 , \4700 );
and \U$13751 ( \14734 , \4679 , \4698 );
nor \U$13752 ( \14735 , \14733 , \14734 );
xnor \U$13753 ( \14736 , \14735 , \4454 );
and \U$13754 ( \14737 , \14732 , \14736 );
and \U$13755 ( \14738 , \5137 , \4305 );
and \U$13756 ( \14739 , \4940 , \4303 );
nor \U$13757 ( \14740 , \14738 , \14739 );
xnor \U$13758 ( \14741 , \14740 , \4118 );
and \U$13759 ( \14742 , \14736 , \14741 );
and \U$13760 ( \14743 , \14732 , \14741 );
or \U$13761 ( \14744 , \14737 , \14742 , \14743 );
and \U$13762 ( \14745 , \14728 , \14744 );
and \U$13763 ( \14746 , \3334 , \6314 );
and \U$13764 ( \14747 , \3309 , \6312 );
nor \U$13765 ( \14748 , \14746 , \14747 );
xnor \U$13766 ( \14749 , \14748 , \6073 );
and \U$13767 ( \14750 , \3675 , \5848 );
and \U$13768 ( \14751 , \3508 , \5846 );
nor \U$13769 ( \14752 , \14750 , \14751 );
xnor \U$13770 ( \14753 , \14752 , \5660 );
and \U$13771 ( \14754 , \14749 , \14753 );
and \U$13772 ( \14755 , \3932 , \5474 );
and \U$13773 ( \14756 , \3813 , \5472 );
nor \U$13774 ( \14757 , \14755 , \14756 );
xnor \U$13775 ( \14758 , \14757 , \5242 );
and \U$13776 ( \14759 , \14753 , \14758 );
and \U$13777 ( \14760 , \14749 , \14758 );
or \U$13778 ( \14761 , \14754 , \14759 , \14760 );
and \U$13779 ( \14762 , \14744 , \14761 );
and \U$13780 ( \14763 , \14728 , \14761 );
or \U$13781 ( \14764 , \14745 , \14762 , \14763 );
and \U$13782 ( \14765 , \14711 , \14764 );
and \U$13783 ( \14766 , \14659 , \14764 );
or \U$13784 ( \14767 , \14712 , \14765 , \14766 );
and \U$13785 ( \14768 , \14607 , \14767 );
xor \U$13786 ( \14769 , \14184 , \14188 );
xor \U$13787 ( \14770 , \14769 , \14193 );
xor \U$13788 ( \14771 , \14297 , \14299 );
xor \U$13789 ( \14772 , \14771 , \14302 );
and \U$13790 ( \14773 , \14770 , \14772 );
xor \U$13791 ( \14774 , \14307 , \14309 );
xor \U$13792 ( \14775 , \14774 , \14312 );
and \U$13793 ( \14776 , \14772 , \14775 );
and \U$13794 ( \14777 , \14770 , \14775 );
or \U$13795 ( \14778 , \14773 , \14776 , \14777 );
and \U$13796 ( \14779 , \14767 , \14778 );
and \U$13797 ( \14780 , \14607 , \14778 );
or \U$13798 ( \14781 , \14768 , \14779 , \14780 );
xor \U$13799 ( \14782 , \14395 , \14411 );
xor \U$13800 ( \14783 , \14782 , \14428 );
xor \U$13801 ( \14784 , \14448 , \14464 );
xor \U$13802 ( \14785 , \14784 , \14481 );
and \U$13803 ( \14786 , \14783 , \14785 );
xor \U$13804 ( \14787 , \14320 , \14322 );
xor \U$13805 ( \14788 , \14787 , \14325 );
and \U$13806 ( \14789 , \14785 , \14788 );
and \U$13807 ( \14790 , \14783 , \14788 );
or \U$13808 ( \14791 , \14786 , \14789 , \14790 );
xor \U$13809 ( \14792 , \14180 , \14196 );
xor \U$13810 ( \14793 , \14792 , \14213 );
and \U$13811 ( \14794 , \14791 , \14793 );
xor \U$13812 ( \14795 , \14503 , \14505 );
xor \U$13813 ( \14796 , \14795 , \14508 );
and \U$13814 ( \14797 , \14793 , \14796 );
and \U$13815 ( \14798 , \14791 , \14796 );
or \U$13816 ( \14799 , \14794 , \14797 , \14798 );
and \U$13817 ( \14800 , \14781 , \14799 );
xor \U$13818 ( \14801 , \14305 , \14315 );
xor \U$13819 ( \14802 , \14801 , \14328 );
xor \U$13820 ( \14803 , \14379 , \14431 );
xor \U$13821 ( \14804 , \14803 , \14484 );
and \U$13822 ( \14805 , \14802 , \14804 );
xor \U$13823 ( \14806 , \14490 , \14492 );
xor \U$13824 ( \14807 , \14806 , \14495 );
and \U$13825 ( \14808 , \14804 , \14807 );
and \U$13826 ( \14809 , \14802 , \14807 );
or \U$13827 ( \14810 , \14805 , \14808 , \14809 );
and \U$13828 ( \14811 , \14799 , \14810 );
and \U$13829 ( \14812 , \14781 , \14810 );
or \U$13830 ( \14813 , \14800 , \14811 , \14812 );
xor \U$13831 ( \14814 , \14331 , \14487 );
xor \U$13832 ( \14815 , \14814 , \14498 );
xor \U$13833 ( \14816 , \14511 , \14513 );
xor \U$13834 ( \14817 , \14816 , \14516 );
and \U$13835 ( \14818 , \14815 , \14817 );
xor \U$13836 ( \14819 , \14522 , \14524 );
xor \U$13837 ( \14820 , \14819 , \14527 );
and \U$13838 ( \14821 , \14817 , \14820 );
and \U$13839 ( \14822 , \14815 , \14820 );
or \U$13840 ( \14823 , \14818 , \14821 , \14822 );
and \U$13841 ( \14824 , \14813 , \14823 );
xor \U$13842 ( \14825 , \14535 , \14537 );
xor \U$13843 ( \14826 , \14825 , \14540 );
and \U$13844 ( \14827 , \14823 , \14826 );
and \U$13845 ( \14828 , \14813 , \14826 );
or \U$13846 ( \14829 , \14824 , \14827 , \14828 );
xor \U$13847 ( \14830 , \14533 , \14543 );
xor \U$13848 ( \14831 , \14830 , \14546 );
and \U$13849 ( \14832 , \14829 , \14831 );
xor \U$13850 ( \14833 , \14551 , \14553 );
xor \U$13851 ( \14834 , \14833 , \14556 );
and \U$13852 ( \14835 , \14831 , \14834 );
and \U$13853 ( \14836 , \14829 , \14834 );
or \U$13854 ( \14837 , \14832 , \14835 , \14836 );
xor \U$13855 ( \14838 , \14549 , \14559 );
xor \U$13856 ( \14839 , \14838 , \14562 );
and \U$13857 ( \14840 , \14837 , \14839 );
xor \U$13858 ( \14841 , \14265 , \14275 );
xor \U$13859 ( \14842 , \14841 , \14278 );
and \U$13860 ( \14843 , \14839 , \14842 );
and \U$13861 ( \14844 , \14837 , \14842 );
or \U$13862 ( \14845 , \14840 , \14843 , \14844 );
and \U$13863 ( \14846 , \14571 , \14845 );
xor \U$13864 ( \14847 , \14571 , \14845 );
xor \U$13865 ( \14848 , \14837 , \14839 );
xor \U$13866 ( \14849 , \14848 , \14842 );
xor \U$13867 ( \14850 , \14716 , \14720 );
xor \U$13868 ( \14851 , \14850 , \14725 );
xor \U$13869 ( \14852 , \14732 , \14736 );
xor \U$13870 ( \14853 , \14852 , \14741 );
and \U$13871 ( \14854 , \14851 , \14853 );
xor \U$13872 ( \14855 , \14749 , \14753 );
xor \U$13873 ( \14856 , \14855 , \14758 );
and \U$13874 ( \14857 , \14853 , \14856 );
and \U$13875 ( \14858 , \14851 , \14856 );
or \U$13876 ( \14859 , \14854 , \14857 , \14858 );
xor \U$13877 ( \14860 , \14611 , \14615 );
xor \U$13878 ( \14861 , \14860 , \14620 );
xor \U$13879 ( \14862 , \14627 , \14631 );
xor \U$13880 ( \14863 , \14862 , \14636 );
and \U$13881 ( \14864 , \14861 , \14863 );
xor \U$13882 ( \14865 , \14644 , \14648 );
xor \U$13883 ( \14866 , \14865 , \14653 );
and \U$13884 ( \14867 , \14863 , \14866 );
and \U$13885 ( \14868 , \14861 , \14866 );
or \U$13886 ( \14869 , \14864 , \14867 , \14868 );
and \U$13887 ( \14870 , \14859 , \14869 );
xor \U$13888 ( \14871 , \14663 , \14667 );
xor \U$13889 ( \14872 , \14871 , \14672 );
xor \U$13890 ( \14873 , \14679 , \14683 );
xor \U$13891 ( \14874 , \14873 , \14688 );
and \U$13892 ( \14875 , \14872 , \14874 );
xor \U$13893 ( \14876 , \14696 , \14700 );
xor \U$13894 ( \14877 , \14876 , \14705 );
and \U$13895 ( \14878 , \14874 , \14877 );
and \U$13896 ( \14879 , \14872 , \14877 );
or \U$13897 ( \14880 , \14875 , \14878 , \14879 );
and \U$13898 ( \14881 , \14869 , \14880 );
and \U$13899 ( \14882 , \14859 , \14880 );
or \U$13900 ( \14883 , \14870 , \14881 , \14882 );
and \U$13901 ( \14884 , \5439 , \4305 );
and \U$13902 ( \14885 , \5137 , \4303 );
nor \U$13903 ( \14886 , \14884 , \14885 );
xnor \U$13904 ( \14887 , \14886 , \4118 );
and \U$13905 ( \14888 , \5916 , \3992 );
and \U$13906 ( \14889 , \5447 , \3990 );
nor \U$13907 ( \14890 , \14888 , \14889 );
xnor \U$13908 ( \14891 , \14890 , \3787 );
and \U$13909 ( \14892 , \14887 , \14891 );
and \U$13910 ( \14893 , \6185 , \3586 );
and \U$13911 ( \14894 , \5921 , \3584 );
nor \U$13912 ( \14895 , \14893 , \14894 );
xnor \U$13913 ( \14896 , \14895 , \3437 );
and \U$13914 ( \14897 , \14891 , \14896 );
and \U$13915 ( \14898 , \14887 , \14896 );
or \U$13916 ( \14899 , \14892 , \14897 , \14898 );
and \U$13917 ( \14900 , \3309 , \6903 );
and \U$13918 ( \14901 , \3045 , \6901 );
nor \U$13919 ( \14902 , \14900 , \14901 );
xnor \U$13920 ( \14903 , \14902 , \6563 );
and \U$13921 ( \14904 , \3508 , \6314 );
and \U$13922 ( \14905 , \3334 , \6312 );
nor \U$13923 ( \14906 , \14904 , \14905 );
xnor \U$13924 ( \14907 , \14906 , \6073 );
and \U$13925 ( \14908 , \14903 , \14907 );
and \U$13926 ( \14909 , \3813 , \5848 );
and \U$13927 ( \14910 , \3675 , \5846 );
nor \U$13928 ( \14911 , \14909 , \14910 );
xnor \U$13929 ( \14912 , \14911 , \5660 );
and \U$13930 ( \14913 , \14907 , \14912 );
and \U$13931 ( \14914 , \14903 , \14912 );
or \U$13932 ( \14915 , \14908 , \14913 , \14914 );
and \U$13933 ( \14916 , \14899 , \14915 );
and \U$13934 ( \14917 , \4349 , \5474 );
and \U$13935 ( \14918 , \3932 , \5472 );
nor \U$13936 ( \14919 , \14917 , \14918 );
xnor \U$13937 ( \14920 , \14919 , \5242 );
and \U$13938 ( \14921 , \4679 , \5023 );
and \U$13939 ( \14922 , \4557 , \5021 );
nor \U$13940 ( \14923 , \14921 , \14922 );
xnor \U$13941 ( \14924 , \14923 , \4880 );
and \U$13942 ( \14925 , \14920 , \14924 );
and \U$13943 ( \14926 , \4940 , \4700 );
and \U$13944 ( \14927 , \4684 , \4698 );
nor \U$13945 ( \14928 , \14926 , \14927 );
xnor \U$13946 ( \14929 , \14928 , \4454 );
and \U$13947 ( \14930 , \14924 , \14929 );
and \U$13948 ( \14931 , \14920 , \14929 );
or \U$13949 ( \14932 , \14925 , \14930 , \14931 );
and \U$13950 ( \14933 , \14915 , \14932 );
and \U$13951 ( \14934 , \14899 , \14932 );
or \U$13952 ( \14935 , \14916 , \14933 , \14934 );
and \U$13953 ( \14936 , \1854 , \10101 );
and \U$13954 ( \14937 , \1656 , \10099 );
nor \U$13955 ( \14938 , \14936 , \14937 );
xnor \U$13956 ( \14939 , \14938 , \9791 );
and \U$13957 ( \14940 , \2047 , \9564 );
and \U$13958 ( \14941 , \1942 , \9562 );
nor \U$13959 ( \14942 , \14940 , \14941 );
xnor \U$13960 ( \14943 , \14942 , \9193 );
and \U$13961 ( \14944 , \14939 , \14943 );
and \U$13962 ( \14945 , \2168 , \9002 );
and \U$13963 ( \14946 , \2052 , \9000 );
nor \U$13964 ( \14947 , \14945 , \14946 );
xnor \U$13965 ( \14948 , \14947 , \8684 );
and \U$13966 ( \14949 , \14943 , \14948 );
and \U$13967 ( \14950 , \14939 , \14948 );
or \U$13968 ( \14951 , \14944 , \14949 , \14950 );
and \U$13969 ( \14952 , \1457 , \11482 );
and \U$13970 ( \14953 , \1377 , \11479 );
nor \U$13971 ( \14954 , \14952 , \14953 );
xnor \U$13972 ( \14955 , \14954 , \10427 );
and \U$13973 ( \14956 , \1593 , \10669 );
and \U$13974 ( \14957 , \1531 , \10667 );
nor \U$13975 ( \14958 , \14956 , \14957 );
xnor \U$13976 ( \14959 , \14958 , \10430 );
and \U$13977 ( \14960 , \14955 , \14959 );
and \U$13978 ( \14961 , \14959 , \1317 );
and \U$13979 ( \14962 , \14955 , \1317 );
or \U$13980 ( \14963 , \14960 , \14961 , \14962 );
and \U$13981 ( \14964 , \14951 , \14963 );
and \U$13982 ( \14965 , \2459 , \8435 );
and \U$13983 ( \14966 , \2283 , \8433 );
nor \U$13984 ( \14967 , \14965 , \14966 );
xnor \U$13985 ( \14968 , \14967 , \8186 );
and \U$13986 ( \14969 , \2710 , \7906 );
and \U$13987 ( \14970 , \2467 , \7904 );
nor \U$13988 ( \14971 , \14969 , \14970 );
xnor \U$13989 ( \14972 , \14971 , \7646 );
and \U$13990 ( \14973 , \14968 , \14972 );
and \U$13991 ( \14974 , \2901 , \7412 );
and \U$13992 ( \14975 , \2715 , \7410 );
nor \U$13993 ( \14976 , \14974 , \14975 );
xnor \U$13994 ( \14977 , \14976 , \7097 );
and \U$13995 ( \14978 , \14972 , \14977 );
and \U$13996 ( \14979 , \14968 , \14977 );
or \U$13997 ( \14980 , \14973 , \14978 , \14979 );
and \U$13998 ( \14981 , \14963 , \14980 );
and \U$13999 ( \14982 , \14951 , \14980 );
or \U$14000 ( \14983 , \14964 , \14981 , \14982 );
and \U$14001 ( \14984 , \14935 , \14983 );
and \U$14002 ( \14985 , \10218 , \1828 );
and \U$14003 ( \14986 , \9649 , \1826 );
nor \U$14004 ( \14987 , \14985 , \14986 );
xnor \U$14005 ( \14988 , \14987 , \1750 );
and \U$14006 ( \14989 , \10829 , \1664 );
and \U$14007 ( \14990 , \10226 , \1662 );
nor \U$14008 ( \14991 , \14989 , \14990 );
xnor \U$14009 ( \14992 , \14991 , \1570 );
and \U$14010 ( \14993 , \14988 , \14992 );
and \U$14011 ( \14994 , \11015 , \1494 );
and \U$14012 ( \14995 , \10834 , \1492 );
nor \U$14013 ( \14996 , \14994 , \14995 );
xnor \U$14014 ( \14997 , \14996 , \1422 );
and \U$14015 ( \14998 , \14992 , \14997 );
and \U$14016 ( \14999 , \14988 , \14997 );
or \U$14017 ( \15000 , \14993 , \14998 , \14999 );
and \U$14018 ( \15001 , \6816 , \3264 );
and \U$14019 ( \15002 , \6444 , \3262 );
nor \U$14020 ( \15003 , \15001 , \15002 );
xnor \U$14021 ( \15004 , \15003 , \3122 );
and \U$14022 ( \15005 , \7168 , \2968 );
and \U$14023 ( \15006 , \6825 , \2966 );
nor \U$14024 ( \15007 , \15005 , \15006 );
xnor \U$14025 ( \15008 , \15007 , \2831 );
and \U$14026 ( \15009 , \15004 , \15008 );
and \U$14027 ( \15010 , \7673 , \2762 );
and \U$14028 ( \15011 , \7370 , \2760 );
nor \U$14029 ( \15012 , \15010 , \15011 );
xnor \U$14030 ( \15013 , \15012 , \2610 );
and \U$14031 ( \15014 , \15008 , \15013 );
and \U$14032 ( \15015 , \15004 , \15013 );
or \U$14033 ( \15016 , \15009 , \15014 , \15015 );
and \U$14034 ( \15017 , \15000 , \15016 );
and \U$14035 ( \15018 , \8371 , \2494 );
and \U$14036 ( \15019 , \7845 , \2492 );
nor \U$14037 ( \15020 , \15018 , \15019 );
xnor \U$14038 ( \15021 , \15020 , \2338 );
and \U$14039 ( \15022 , \9041 , \2222 );
and \U$14040 ( \15023 , \8795 , \2220 );
nor \U$14041 ( \15024 , \15022 , \15023 );
xnor \U$14042 ( \15025 , \15024 , \2109 );
and \U$14043 ( \15026 , \15021 , \15025 );
and \U$14044 ( \15027 , \9365 , \2028 );
and \U$14045 ( \15028 , \9046 , \2026 );
nor \U$14046 ( \15029 , \15027 , \15028 );
xnor \U$14047 ( \15030 , \15029 , \1892 );
and \U$14048 ( \15031 , \15025 , \15030 );
and \U$14049 ( \15032 , \15021 , \15030 );
or \U$14050 ( \15033 , \15026 , \15031 , \15032 );
and \U$14051 ( \15034 , \15016 , \15033 );
and \U$14052 ( \15035 , \15000 , \15033 );
or \U$14053 ( \15036 , \15017 , \15034 , \15035 );
and \U$14054 ( \15037 , \14983 , \15036 );
and \U$14055 ( \15038 , \14935 , \15036 );
or \U$14056 ( \15039 , \14984 , \15037 , \15038 );
and \U$14057 ( \15040 , \14883 , \15039 );
xor \U$14058 ( \15041 , \14351 , \14355 );
xor \U$14059 ( \15042 , \15041 , \14360 );
xor \U$14060 ( \15043 , \14368 , \14372 );
xor \U$14061 ( \15044 , \15043 , \1198 );
and \U$14062 ( \15045 , \15042 , \15044 );
xor \U$14063 ( \15046 , \14596 , \14598 );
xor \U$14064 ( \15047 , \15046 , \14601 );
and \U$14065 ( \15048 , \15044 , \15047 );
and \U$14066 ( \15049 , \15042 , \15047 );
or \U$14067 ( \15050 , \15045 , \15048 , \15049 );
and \U$14068 ( \15051 , \15039 , \15050 );
and \U$14069 ( \15052 , \14883 , \15050 );
or \U$14070 ( \15053 , \15040 , \15051 , \15052 );
xor \U$14071 ( \15054 , \14623 , \14639 );
xor \U$14072 ( \15055 , \15054 , \14656 );
xor \U$14073 ( \15056 , \14573 , \14575 );
xor \U$14074 ( \15057 , \15056 , \14578 );
and \U$14075 ( \15058 , \15055 , \15057 );
xor \U$14076 ( \15059 , \14585 , \14587 );
xor \U$14077 ( \15060 , \15059 , \14590 );
and \U$14078 ( \15061 , \15057 , \15060 );
and \U$14079 ( \15062 , \15055 , \15060 );
or \U$14080 ( \15063 , \15058 , \15061 , \15062 );
xor \U$14081 ( \15064 , \14675 , \14691 );
xor \U$14082 ( \15065 , \15064 , \14708 );
xor \U$14083 ( \15066 , \14728 , \14744 );
xor \U$14084 ( \15067 , \15066 , \14761 );
and \U$14085 ( \15068 , \15065 , \15067 );
and \U$14086 ( \15069 , \15063 , \15068 );
xor \U$14087 ( \15070 , \14347 , \14363 );
xor \U$14088 ( \15071 , \15070 , \14376 );
and \U$14089 ( \15072 , \15068 , \15071 );
and \U$14090 ( \15073 , \15063 , \15071 );
or \U$14091 ( \15074 , \15069 , \15072 , \15073 );
and \U$14092 ( \15075 , \15053 , \15074 );
xor \U$14093 ( \15076 , \14581 , \14593 );
xor \U$14094 ( \15077 , \15076 , \14604 );
xor \U$14095 ( \15078 , \14783 , \14785 );
xor \U$14096 ( \15079 , \15078 , \14788 );
and \U$14097 ( \15080 , \15077 , \15079 );
xor \U$14098 ( \15081 , \14770 , \14772 );
xor \U$14099 ( \15082 , \15081 , \14775 );
and \U$14100 ( \15083 , \15079 , \15082 );
and \U$14101 ( \15084 , \15077 , \15082 );
or \U$14102 ( \15085 , \15080 , \15083 , \15084 );
and \U$14103 ( \15086 , \15074 , \15085 );
and \U$14104 ( \15087 , \15053 , \15085 );
or \U$14105 ( \15088 , \15075 , \15086 , \15087 );
xor \U$14106 ( \15089 , \14607 , \14767 );
xor \U$14107 ( \15090 , \15089 , \14778 );
xor \U$14108 ( \15091 , \14791 , \14793 );
xor \U$14109 ( \15092 , \15091 , \14796 );
and \U$14110 ( \15093 , \15090 , \15092 );
xor \U$14111 ( \15094 , \14802 , \14804 );
xor \U$14112 ( \15095 , \15094 , \14807 );
and \U$14113 ( \15096 , \15092 , \15095 );
and \U$14114 ( \15097 , \15090 , \15095 );
or \U$14115 ( \15098 , \15093 , \15096 , \15097 );
and \U$14116 ( \15099 , \15088 , \15098 );
xor \U$14117 ( \15100 , \14815 , \14817 );
xor \U$14118 ( \15101 , \15100 , \14820 );
and \U$14119 ( \15102 , \15098 , \15101 );
and \U$14120 ( \15103 , \15088 , \15101 );
or \U$14121 ( \15104 , \15099 , \15102 , \15103 );
xor \U$14122 ( \15105 , \14501 , \14519 );
xor \U$14123 ( \15106 , \15105 , \14530 );
and \U$14124 ( \15107 , \15104 , \15106 );
xor \U$14125 ( \15108 , \14813 , \14823 );
xor \U$14126 ( \15109 , \15108 , \14826 );
and \U$14127 ( \15110 , \15106 , \15109 );
and \U$14128 ( \15111 , \15104 , \15109 );
or \U$14129 ( \15112 , \15107 , \15110 , \15111 );
xor \U$14130 ( \15113 , \14829 , \14831 );
xor \U$14131 ( \15114 , \15113 , \14834 );
and \U$14132 ( \15115 , \15112 , \15114 );
and \U$14133 ( \15116 , \14849 , \15115 );
xor \U$14134 ( \15117 , \14849 , \15115 );
xor \U$14135 ( \15118 , \15112 , \15114 );
and \U$14136 ( \15119 , \4684 , \5023 );
and \U$14137 ( \15120 , \4679 , \5021 );
nor \U$14138 ( \15121 , \15119 , \15120 );
xnor \U$14139 ( \15122 , \15121 , \4880 );
and \U$14140 ( \15123 , \5137 , \4700 );
and \U$14141 ( \15124 , \4940 , \4698 );
nor \U$14142 ( \15125 , \15123 , \15124 );
xnor \U$14143 ( \15126 , \15125 , \4454 );
and \U$14144 ( \15127 , \15122 , \15126 );
and \U$14145 ( \15128 , \5447 , \4305 );
and \U$14146 ( \15129 , \5439 , \4303 );
nor \U$14147 ( \15130 , \15128 , \15129 );
xnor \U$14148 ( \15131 , \15130 , \4118 );
and \U$14149 ( \15132 , \15126 , \15131 );
and \U$14150 ( \15133 , \15122 , \15131 );
or \U$14151 ( \15134 , \15127 , \15132 , \15133 );
and \U$14152 ( \15135 , \3675 , \6314 );
and \U$14153 ( \15136 , \3508 , \6312 );
nor \U$14154 ( \15137 , \15135 , \15136 );
xnor \U$14155 ( \15138 , \15137 , \6073 );
and \U$14156 ( \15139 , \3932 , \5848 );
and \U$14157 ( \15140 , \3813 , \5846 );
nor \U$14158 ( \15141 , \15139 , \15140 );
xnor \U$14159 ( \15142 , \15141 , \5660 );
and \U$14160 ( \15143 , \15138 , \15142 );
and \U$14161 ( \15144 , \4557 , \5474 );
and \U$14162 ( \15145 , \4349 , \5472 );
nor \U$14163 ( \15146 , \15144 , \15145 );
xnor \U$14164 ( \15147 , \15146 , \5242 );
and \U$14165 ( \15148 , \15142 , \15147 );
and \U$14166 ( \15149 , \15138 , \15147 );
or \U$14167 ( \15150 , \15143 , \15148 , \15149 );
and \U$14168 ( \15151 , \15134 , \15150 );
and \U$14169 ( \15152 , \5921 , \3992 );
and \U$14170 ( \15153 , \5916 , \3990 );
nor \U$14171 ( \15154 , \15152 , \15153 );
xnor \U$14172 ( \15155 , \15154 , \3787 );
and \U$14173 ( \15156 , \6444 , \3586 );
and \U$14174 ( \15157 , \6185 , \3584 );
nor \U$14175 ( \15158 , \15156 , \15157 );
xnor \U$14176 ( \15159 , \15158 , \3437 );
and \U$14177 ( \15160 , \15155 , \15159 );
and \U$14178 ( \15161 , \6825 , \3264 );
and \U$14179 ( \15162 , \6816 , \3262 );
nor \U$14180 ( \15163 , \15161 , \15162 );
xnor \U$14181 ( \15164 , \15163 , \3122 );
and \U$14182 ( \15165 , \15159 , \15164 );
and \U$14183 ( \15166 , \15155 , \15164 );
or \U$14184 ( \15167 , \15160 , \15165 , \15166 );
and \U$14185 ( \15168 , \15150 , \15167 );
and \U$14186 ( \15169 , \15134 , \15167 );
or \U$14187 ( \15170 , \15151 , \15168 , \15169 );
and \U$14188 ( \15171 , \9046 , \2222 );
and \U$14189 ( \15172 , \9041 , \2220 );
nor \U$14190 ( \15173 , \15171 , \15172 );
xnor \U$14191 ( \15174 , \15173 , \2109 );
and \U$14192 ( \15175 , \9649 , \2028 );
and \U$14193 ( \15176 , \9365 , \2026 );
nor \U$14194 ( \15177 , \15175 , \15176 );
xnor \U$14195 ( \15178 , \15177 , \1892 );
and \U$14196 ( \15179 , \15174 , \15178 );
and \U$14197 ( \15180 , \10226 , \1828 );
and \U$14198 ( \15181 , \10218 , \1826 );
nor \U$14199 ( \15182 , \15180 , \15181 );
xnor \U$14200 ( \15183 , \15182 , \1750 );
and \U$14201 ( \15184 , \15178 , \15183 );
and \U$14202 ( \15185 , \15174 , \15183 );
or \U$14203 ( \15186 , \15179 , \15184 , \15185 );
and \U$14204 ( \15187 , \7370 , \2968 );
and \U$14205 ( \15188 , \7168 , \2966 );
nor \U$14206 ( \15189 , \15187 , \15188 );
xnor \U$14207 ( \15190 , \15189 , \2831 );
and \U$14208 ( \15191 , \7845 , \2762 );
and \U$14209 ( \15192 , \7673 , \2760 );
nor \U$14210 ( \15193 , \15191 , \15192 );
xnor \U$14211 ( \15194 , \15193 , \2610 );
and \U$14212 ( \15195 , \15190 , \15194 );
and \U$14213 ( \15196 , \8795 , \2494 );
and \U$14214 ( \15197 , \8371 , \2492 );
nor \U$14215 ( \15198 , \15196 , \15197 );
xnor \U$14216 ( \15199 , \15198 , \2338 );
and \U$14217 ( \15200 , \15194 , \15199 );
and \U$14218 ( \15201 , \15190 , \15199 );
or \U$14219 ( \15202 , \15195 , \15200 , \15201 );
and \U$14220 ( \15203 , \15186 , \15202 );
and \U$14221 ( \15204 , \10834 , \1664 );
and \U$14222 ( \15205 , \10829 , \1662 );
nor \U$14223 ( \15206 , \15204 , \15205 );
xnor \U$14224 ( \15207 , \15206 , \1570 );
and \U$14225 ( \15208 , \11635 , \1494 );
and \U$14226 ( \15209 , \11015 , \1492 );
nor \U$14227 ( \15210 , \15208 , \15209 );
xnor \U$14228 ( \15211 , \15210 , \1422 );
and \U$14229 ( \15212 , \15207 , \15211 );
and \U$14230 ( \15213 , \15202 , \15212 );
and \U$14231 ( \15214 , \15186 , \15212 );
or \U$14232 ( \15215 , \15203 , \15213 , \15214 );
and \U$14233 ( \15216 , \15170 , \15215 );
and \U$14234 ( \15217 , \2715 , \7906 );
and \U$14235 ( \15218 , \2710 , \7904 );
nor \U$14236 ( \15219 , \15217 , \15218 );
xnor \U$14237 ( \15220 , \15219 , \7646 );
and \U$14238 ( \15221 , \3045 , \7412 );
and \U$14239 ( \15222 , \2901 , \7410 );
nor \U$14240 ( \15223 , \15221 , \15222 );
xnor \U$14241 ( \15224 , \15223 , \7097 );
and \U$14242 ( \15225 , \15220 , \15224 );
and \U$14243 ( \15226 , \3334 , \6903 );
and \U$14244 ( \15227 , \3309 , \6901 );
nor \U$14245 ( \15228 , \15226 , \15227 );
xnor \U$14246 ( \15229 , \15228 , \6563 );
and \U$14247 ( \15230 , \15224 , \15229 );
and \U$14248 ( \15231 , \15220 , \15229 );
or \U$14249 ( \15232 , \15225 , \15230 , \15231 );
and \U$14250 ( \15233 , \1531 , \11482 );
and \U$14251 ( \15234 , \1457 , \11479 );
nor \U$14252 ( \15235 , \15233 , \15234 );
xnor \U$14253 ( \15236 , \15235 , \10427 );
and \U$14254 ( \15237 , \1656 , \10669 );
and \U$14255 ( \15238 , \1593 , \10667 );
nor \U$14256 ( \15239 , \15237 , \15238 );
xnor \U$14257 ( \15240 , \15239 , \10430 );
and \U$14258 ( \15241 , \15236 , \15240 );
and \U$14259 ( \15242 , \1942 , \10101 );
and \U$14260 ( \15243 , \1854 , \10099 );
nor \U$14261 ( \15244 , \15242 , \15243 );
xnor \U$14262 ( \15245 , \15244 , \9791 );
and \U$14263 ( \15246 , \15240 , \15245 );
and \U$14264 ( \15247 , \15236 , \15245 );
or \U$14265 ( \15248 , \15241 , \15246 , \15247 );
and \U$14266 ( \15249 , \15232 , \15248 );
and \U$14267 ( \15250 , \2052 , \9564 );
and \U$14268 ( \15251 , \2047 , \9562 );
nor \U$14269 ( \15252 , \15250 , \15251 );
xnor \U$14270 ( \15253 , \15252 , \9193 );
and \U$14271 ( \15254 , \2283 , \9002 );
and \U$14272 ( \15255 , \2168 , \9000 );
nor \U$14273 ( \15256 , \15254 , \15255 );
xnor \U$14274 ( \15257 , \15256 , \8684 );
and \U$14275 ( \15258 , \15253 , \15257 );
and \U$14276 ( \15259 , \2467 , \8435 );
and \U$14277 ( \15260 , \2459 , \8433 );
nor \U$14278 ( \15261 , \15259 , \15260 );
xnor \U$14279 ( \15262 , \15261 , \8186 );
and \U$14280 ( \15263 , \15257 , \15262 );
and \U$14281 ( \15264 , \15253 , \15262 );
or \U$14282 ( \15265 , \15258 , \15263 , \15264 );
and \U$14283 ( \15266 , \15248 , \15265 );
and \U$14284 ( \15267 , \15232 , \15265 );
or \U$14285 ( \15268 , \15249 , \15266 , \15267 );
and \U$14286 ( \15269 , \15215 , \15268 );
and \U$14287 ( \15270 , \15170 , \15268 );
or \U$14288 ( \15271 , \15216 , \15269 , \15270 );
xor \U$14289 ( \15272 , \14939 , \14943 );
xor \U$14290 ( \15273 , \15272 , \14948 );
xor \U$14291 ( \15274 , \14968 , \14972 );
xor \U$14292 ( \15275 , \15274 , \14977 );
and \U$14293 ( \15276 , \15273 , \15275 );
xor \U$14294 ( \15277 , \14903 , \14907 );
xor \U$14295 ( \15278 , \15277 , \14912 );
and \U$14296 ( \15279 , \15275 , \15278 );
and \U$14297 ( \15280 , \15273 , \15278 );
or \U$14298 ( \15281 , \15276 , \15279 , \15280 );
nand \U$14299 ( \15282 , \11635 , \1358 );
xnor \U$14300 ( \15283 , \15282 , \1317 );
xor \U$14301 ( \15284 , \14988 , \14992 );
xor \U$14302 ( \15285 , \15284 , \14997 );
and \U$14303 ( \15286 , \15283 , \15285 );
xor \U$14304 ( \15287 , \15021 , \15025 );
xor \U$14305 ( \15288 , \15287 , \15030 );
and \U$14306 ( \15289 , \15285 , \15288 );
and \U$14307 ( \15290 , \15283 , \15288 );
or \U$14308 ( \15291 , \15286 , \15289 , \15290 );
and \U$14309 ( \15292 , \15281 , \15291 );
xor \U$14310 ( \15293 , \15004 , \15008 );
xor \U$14311 ( \15294 , \15293 , \15013 );
xor \U$14312 ( \15295 , \14887 , \14891 );
xor \U$14313 ( \15296 , \15295 , \14896 );
and \U$14314 ( \15297 , \15294 , \15296 );
xor \U$14315 ( \15298 , \14920 , \14924 );
xor \U$14316 ( \15299 , \15298 , \14929 );
and \U$14317 ( \15300 , \15296 , \15299 );
and \U$14318 ( \15301 , \15294 , \15299 );
or \U$14319 ( \15302 , \15297 , \15300 , \15301 );
and \U$14320 ( \15303 , \15291 , \15302 );
and \U$14321 ( \15304 , \15281 , \15302 );
or \U$14322 ( \15305 , \15292 , \15303 , \15304 );
and \U$14323 ( \15306 , \15271 , \15305 );
xor \U$14324 ( \15307 , \14851 , \14853 );
xor \U$14325 ( \15308 , \15307 , \14856 );
xor \U$14326 ( \15309 , \14861 , \14863 );
xor \U$14327 ( \15310 , \15309 , \14866 );
and \U$14328 ( \15311 , \15308 , \15310 );
xor \U$14329 ( \15312 , \14872 , \14874 );
xor \U$14330 ( \15313 , \15312 , \14877 );
and \U$14331 ( \15314 , \15310 , \15313 );
and \U$14332 ( \15315 , \15308 , \15313 );
or \U$14333 ( \15316 , \15311 , \15314 , \15315 );
and \U$14334 ( \15317 , \15305 , \15316 );
and \U$14335 ( \15318 , \15271 , \15316 );
or \U$14336 ( \15319 , \15306 , \15317 , \15318 );
xor \U$14337 ( \15320 , \14859 , \14869 );
xor \U$14338 ( \15321 , \15320 , \14880 );
xor \U$14339 ( \15322 , \14935 , \14983 );
xor \U$14340 ( \15323 , \15322 , \15036 );
and \U$14341 ( \15324 , \15321 , \15323 );
xor \U$14342 ( \15325 , \15042 , \15044 );
xor \U$14343 ( \15326 , \15325 , \15047 );
and \U$14344 ( \15327 , \15323 , \15326 );
and \U$14345 ( \15328 , \15321 , \15326 );
or \U$14346 ( \15329 , \15324 , \15327 , \15328 );
and \U$14347 ( \15330 , \15319 , \15329 );
xor \U$14348 ( \15331 , \14899 , \14915 );
xor \U$14349 ( \15332 , \15331 , \14932 );
xor \U$14350 ( \15333 , \14951 , \14963 );
xor \U$14351 ( \15334 , \15333 , \14980 );
and \U$14352 ( \15335 , \15332 , \15334 );
xor \U$14353 ( \15336 , \15000 , \15016 );
xor \U$14354 ( \15337 , \15336 , \15033 );
and \U$14355 ( \15338 , \15334 , \15337 );
and \U$14356 ( \15339 , \15332 , \15337 );
or \U$14357 ( \15340 , \15335 , \15338 , \15339 );
xor \U$14358 ( \15341 , \15055 , \15057 );
xor \U$14359 ( \15342 , \15341 , \15060 );
and \U$14360 ( \15343 , \15340 , \15342 );
xor \U$14361 ( \15344 , \15065 , \15067 );
and \U$14362 ( \15345 , \15342 , \15344 );
and \U$14363 ( \15346 , \15340 , \15344 );
or \U$14364 ( \15347 , \15343 , \15345 , \15346 );
and \U$14365 ( \15348 , \15329 , \15347 );
and \U$14366 ( \15349 , \15319 , \15347 );
or \U$14367 ( \15350 , \15330 , \15348 , \15349 );
xor \U$14368 ( \15351 , \14659 , \14711 );
xor \U$14369 ( \15352 , \15351 , \14764 );
xor \U$14370 ( \15353 , \15063 , \15068 );
xor \U$14371 ( \15354 , \15353 , \15071 );
and \U$14372 ( \15355 , \15352 , \15354 );
xor \U$14373 ( \15356 , \15077 , \15079 );
xor \U$14374 ( \15357 , \15356 , \15082 );
and \U$14375 ( \15358 , \15354 , \15357 );
and \U$14376 ( \15359 , \15352 , \15357 );
or \U$14377 ( \15360 , \15355 , \15358 , \15359 );
and \U$14378 ( \15361 , \15350 , \15360 );
xor \U$14379 ( \15362 , \15090 , \15092 );
xor \U$14380 ( \15363 , \15362 , \15095 );
and \U$14381 ( \15364 , \15360 , \15363 );
and \U$14382 ( \15365 , \15350 , \15363 );
or \U$14383 ( \15366 , \15361 , \15364 , \15365 );
xor \U$14384 ( \15367 , \14781 , \14799 );
xor \U$14385 ( \15368 , \15367 , \14810 );
and \U$14386 ( \15369 , \15366 , \15368 );
xor \U$14387 ( \15370 , \15088 , \15098 );
xor \U$14388 ( \15371 , \15370 , \15101 );
and \U$14389 ( \15372 , \15368 , \15371 );
and \U$14390 ( \15373 , \15366 , \15371 );
or \U$14391 ( \15374 , \15369 , \15372 , \15373 );
xor \U$14392 ( \15375 , \15104 , \15106 );
xor \U$14393 ( \15376 , \15375 , \15109 );
and \U$14394 ( \15377 , \15374 , \15376 );
and \U$14395 ( \15378 , \15118 , \15377 );
xor \U$14396 ( \15379 , \15118 , \15377 );
xor \U$14397 ( \15380 , \15374 , \15376 );
and \U$14398 ( \15381 , \4679 , \5474 );
and \U$14399 ( \15382 , \4557 , \5472 );
nor \U$14400 ( \15383 , \15381 , \15382 );
xnor \U$14401 ( \15384 , \15383 , \5242 );
and \U$14402 ( \15385 , \4940 , \5023 );
and \U$14403 ( \15386 , \4684 , \5021 );
nor \U$14404 ( \15387 , \15385 , \15386 );
xnor \U$14405 ( \15388 , \15387 , \4880 );
and \U$14406 ( \15389 , \15384 , \15388 );
and \U$14407 ( \15390 , \5439 , \4700 );
and \U$14408 ( \15391 , \5137 , \4698 );
nor \U$14409 ( \15392 , \15390 , \15391 );
xnor \U$14410 ( \15393 , \15392 , \4454 );
and \U$14411 ( \15394 , \15388 , \15393 );
and \U$14412 ( \15395 , \15384 , \15393 );
or \U$14413 ( \15396 , \15389 , \15394 , \15395 );
and \U$14414 ( \15397 , \3508 , \6903 );
and \U$14415 ( \15398 , \3334 , \6901 );
nor \U$14416 ( \15399 , \15397 , \15398 );
xnor \U$14417 ( \15400 , \15399 , \6563 );
and \U$14418 ( \15401 , \3813 , \6314 );
and \U$14419 ( \15402 , \3675 , \6312 );
nor \U$14420 ( \15403 , \15401 , \15402 );
xnor \U$14421 ( \15404 , \15403 , \6073 );
and \U$14422 ( \15405 , \15400 , \15404 );
and \U$14423 ( \15406 , \4349 , \5848 );
and \U$14424 ( \15407 , \3932 , \5846 );
nor \U$14425 ( \15408 , \15406 , \15407 );
xnor \U$14426 ( \15409 , \15408 , \5660 );
and \U$14427 ( \15410 , \15404 , \15409 );
and \U$14428 ( \15411 , \15400 , \15409 );
or \U$14429 ( \15412 , \15405 , \15410 , \15411 );
and \U$14430 ( \15413 , \15396 , \15412 );
and \U$14431 ( \15414 , \5916 , \4305 );
and \U$14432 ( \15415 , \5447 , \4303 );
nor \U$14433 ( \15416 , \15414 , \15415 );
xnor \U$14434 ( \15417 , \15416 , \4118 );
and \U$14435 ( \15418 , \6185 , \3992 );
and \U$14436 ( \15419 , \5921 , \3990 );
nor \U$14437 ( \15420 , \15418 , \15419 );
xnor \U$14438 ( \15421 , \15420 , \3787 );
and \U$14439 ( \15422 , \15417 , \15421 );
and \U$14440 ( \15423 , \6816 , \3586 );
and \U$14441 ( \15424 , \6444 , \3584 );
nor \U$14442 ( \15425 , \15423 , \15424 );
xnor \U$14443 ( \15426 , \15425 , \3437 );
and \U$14444 ( \15427 , \15421 , \15426 );
and \U$14445 ( \15428 , \15417 , \15426 );
or \U$14446 ( \15429 , \15422 , \15427 , \15428 );
and \U$14447 ( \15430 , \15412 , \15429 );
and \U$14448 ( \15431 , \15396 , \15429 );
or \U$14449 ( \15432 , \15413 , \15430 , \15431 );
and \U$14450 ( \15433 , \2710 , \8435 );
and \U$14451 ( \15434 , \2467 , \8433 );
nor \U$14452 ( \15435 , \15433 , \15434 );
xnor \U$14453 ( \15436 , \15435 , \8186 );
and \U$14454 ( \15437 , \2901 , \7906 );
and \U$14455 ( \15438 , \2715 , \7904 );
nor \U$14456 ( \15439 , \15437 , \15438 );
xnor \U$14457 ( \15440 , \15439 , \7646 );
and \U$14458 ( \15441 , \15436 , \15440 );
and \U$14459 ( \15442 , \3309 , \7412 );
and \U$14460 ( \15443 , \3045 , \7410 );
nor \U$14461 ( \15444 , \15442 , \15443 );
xnor \U$14462 ( \15445 , \15444 , \7097 );
and \U$14463 ( \15446 , \15440 , \15445 );
and \U$14464 ( \15447 , \15436 , \15445 );
or \U$14465 ( \15448 , \15441 , \15446 , \15447 );
and \U$14466 ( \15449 , \2047 , \10101 );
and \U$14467 ( \15450 , \1942 , \10099 );
nor \U$14468 ( \15451 , \15449 , \15450 );
xnor \U$14469 ( \15452 , \15451 , \9791 );
and \U$14470 ( \15453 , \2168 , \9564 );
and \U$14471 ( \15454 , \2052 , \9562 );
nor \U$14472 ( \15455 , \15453 , \15454 );
xnor \U$14473 ( \15456 , \15455 , \9193 );
and \U$14474 ( \15457 , \15452 , \15456 );
and \U$14475 ( \15458 , \2459 , \9002 );
and \U$14476 ( \15459 , \2283 , \9000 );
nor \U$14477 ( \15460 , \15458 , \15459 );
xnor \U$14478 ( \15461 , \15460 , \8684 );
and \U$14479 ( \15462 , \15456 , \15461 );
and \U$14480 ( \15463 , \15452 , \15461 );
or \U$14481 ( \15464 , \15457 , \15462 , \15463 );
and \U$14482 ( \15465 , \15448 , \15464 );
and \U$14483 ( \15466 , \1593 , \11482 );
and \U$14484 ( \15467 , \1531 , \11479 );
nor \U$14485 ( \15468 , \15466 , \15467 );
xnor \U$14486 ( \15469 , \15468 , \10427 );
and \U$14487 ( \15470 , \1854 , \10669 );
and \U$14488 ( \15471 , \1656 , \10667 );
nor \U$14489 ( \15472 , \15470 , \15471 );
xnor \U$14490 ( \15473 , \15472 , \10430 );
and \U$14491 ( \15474 , \15469 , \15473 );
and \U$14492 ( \15475 , \15473 , \1422 );
and \U$14493 ( \15476 , \15469 , \1422 );
or \U$14494 ( \15477 , \15474 , \15475 , \15476 );
and \U$14495 ( \15478 , \15464 , \15477 );
and \U$14496 ( \15479 , \15448 , \15477 );
or \U$14497 ( \15480 , \15465 , \15478 , \15479 );
and \U$14498 ( \15481 , \15432 , \15480 );
and \U$14499 ( \15482 , \7168 , \3264 );
and \U$14500 ( \15483 , \6825 , \3262 );
nor \U$14501 ( \15484 , \15482 , \15483 );
xnor \U$14502 ( \15485 , \15484 , \3122 );
and \U$14503 ( \15486 , \7673 , \2968 );
and \U$14504 ( \15487 , \7370 , \2966 );
nor \U$14505 ( \15488 , \15486 , \15487 );
xnor \U$14506 ( \15489 , \15488 , \2831 );
and \U$14507 ( \15490 , \15485 , \15489 );
and \U$14508 ( \15491 , \8371 , \2762 );
and \U$14509 ( \15492 , \7845 , \2760 );
nor \U$14510 ( \15493 , \15491 , \15492 );
xnor \U$14511 ( \15494 , \15493 , \2610 );
and \U$14512 ( \15495 , \15489 , \15494 );
and \U$14513 ( \15496 , \15485 , \15494 );
or \U$14514 ( \15497 , \15490 , \15495 , \15496 );
and \U$14515 ( \15498 , \10829 , \1828 );
and \U$14516 ( \15499 , \10226 , \1826 );
nor \U$14517 ( \15500 , \15498 , \15499 );
xnor \U$14518 ( \15501 , \15500 , \1750 );
and \U$14519 ( \15502 , \11015 , \1664 );
and \U$14520 ( \15503 , \10834 , \1662 );
nor \U$14521 ( \15504 , \15502 , \15503 );
xnor \U$14522 ( \15505 , \15504 , \1570 );
and \U$14523 ( \15506 , \15501 , \15505 );
nand \U$14524 ( \15507 , \11635 , \1492 );
xnor \U$14525 ( \15508 , \15507 , \1422 );
and \U$14526 ( \15509 , \15505 , \15508 );
and \U$14527 ( \15510 , \15501 , \15508 );
or \U$14528 ( \15511 , \15506 , \15509 , \15510 );
and \U$14529 ( \15512 , \15497 , \15511 );
and \U$14530 ( \15513 , \9041 , \2494 );
and \U$14531 ( \15514 , \8795 , \2492 );
nor \U$14532 ( \15515 , \15513 , \15514 );
xnor \U$14533 ( \15516 , \15515 , \2338 );
and \U$14534 ( \15517 , \9365 , \2222 );
and \U$14535 ( \15518 , \9046 , \2220 );
nor \U$14536 ( \15519 , \15517 , \15518 );
xnor \U$14537 ( \15520 , \15519 , \2109 );
and \U$14538 ( \15521 , \15516 , \15520 );
and \U$14539 ( \15522 , \10218 , \2028 );
and \U$14540 ( \15523 , \9649 , \2026 );
nor \U$14541 ( \15524 , \15522 , \15523 );
xnor \U$14542 ( \15525 , \15524 , \1892 );
and \U$14543 ( \15526 , \15520 , \15525 );
and \U$14544 ( \15527 , \15516 , \15525 );
or \U$14545 ( \15528 , \15521 , \15526 , \15527 );
and \U$14546 ( \15529 , \15511 , \15528 );
and \U$14547 ( \15530 , \15497 , \15528 );
or \U$14548 ( \15531 , \15512 , \15529 , \15530 );
and \U$14549 ( \15532 , \15480 , \15531 );
and \U$14550 ( \15533 , \15432 , \15531 );
or \U$14551 ( \15534 , \15481 , \15532 , \15533 );
xor \U$14552 ( \15535 , \15220 , \15224 );
xor \U$14553 ( \15536 , \15535 , \15229 );
xor \U$14554 ( \15537 , \15236 , \15240 );
xor \U$14555 ( \15538 , \15537 , \15245 );
and \U$14556 ( \15539 , \15536 , \15538 );
xor \U$14557 ( \15540 , \15253 , \15257 );
xor \U$14558 ( \15541 , \15540 , \15262 );
and \U$14559 ( \15542 , \15538 , \15541 );
and \U$14560 ( \15543 , \15536 , \15541 );
or \U$14561 ( \15544 , \15539 , \15542 , \15543 );
xor \U$14562 ( \15545 , \15122 , \15126 );
xor \U$14563 ( \15546 , \15545 , \15131 );
xor \U$14564 ( \15547 , \15138 , \15142 );
xor \U$14565 ( \15548 , \15547 , \15147 );
and \U$14566 ( \15549 , \15546 , \15548 );
xor \U$14567 ( \15550 , \15155 , \15159 );
xor \U$14568 ( \15551 , \15550 , \15164 );
and \U$14569 ( \15552 , \15548 , \15551 );
and \U$14570 ( \15553 , \15546 , \15551 );
or \U$14571 ( \15554 , \15549 , \15552 , \15553 );
and \U$14572 ( \15555 , \15544 , \15554 );
xor \U$14573 ( \15556 , \15174 , \15178 );
xor \U$14574 ( \15557 , \15556 , \15183 );
xor \U$14575 ( \15558 , \15190 , \15194 );
xor \U$14576 ( \15559 , \15558 , \15199 );
and \U$14577 ( \15560 , \15557 , \15559 );
xor \U$14578 ( \15561 , \15207 , \15211 );
and \U$14579 ( \15562 , \15559 , \15561 );
and \U$14580 ( \15563 , \15557 , \15561 );
or \U$14581 ( \15564 , \15560 , \15562 , \15563 );
and \U$14582 ( \15565 , \15554 , \15564 );
and \U$14583 ( \15566 , \15544 , \15564 );
or \U$14584 ( \15567 , \15555 , \15565 , \15566 );
and \U$14585 ( \15568 , \15534 , \15567 );
xor \U$14586 ( \15569 , \14955 , \14959 );
xor \U$14587 ( \15570 , \15569 , \1317 );
xor \U$14588 ( \15571 , \15273 , \15275 );
xor \U$14589 ( \15572 , \15571 , \15278 );
and \U$14590 ( \15573 , \15570 , \15572 );
xor \U$14591 ( \15574 , \15294 , \15296 );
xor \U$14592 ( \15575 , \15574 , \15299 );
and \U$14593 ( \15576 , \15572 , \15575 );
and \U$14594 ( \15577 , \15570 , \15575 );
or \U$14595 ( \15578 , \15573 , \15576 , \15577 );
and \U$14596 ( \15579 , \15567 , \15578 );
and \U$14597 ( \15580 , \15534 , \15578 );
or \U$14598 ( \15581 , \15568 , \15579 , \15580 );
xor \U$14599 ( \15582 , \15134 , \15150 );
xor \U$14600 ( \15583 , \15582 , \15167 );
xor \U$14601 ( \15584 , \15186 , \15202 );
xor \U$14602 ( \15585 , \15584 , \15212 );
and \U$14603 ( \15586 , \15583 , \15585 );
xor \U$14604 ( \15587 , \15283 , \15285 );
xor \U$14605 ( \15588 , \15587 , \15288 );
and \U$14606 ( \15589 , \15585 , \15588 );
and \U$14607 ( \15590 , \15583 , \15588 );
or \U$14608 ( \15591 , \15586 , \15589 , \15590 );
xor \U$14609 ( \15592 , \15332 , \15334 );
xor \U$14610 ( \15593 , \15592 , \15337 );
and \U$14611 ( \15594 , \15591 , \15593 );
xor \U$14612 ( \15595 , \15308 , \15310 );
xor \U$14613 ( \15596 , \15595 , \15313 );
and \U$14614 ( \15597 , \15593 , \15596 );
and \U$14615 ( \15598 , \15591 , \15596 );
or \U$14616 ( \15599 , \15594 , \15597 , \15598 );
and \U$14617 ( \15600 , \15581 , \15599 );
xor \U$14618 ( \15601 , \15170 , \15215 );
xor \U$14619 ( \15602 , \15601 , \15268 );
xor \U$14620 ( \15603 , \15281 , \15291 );
xor \U$14621 ( \15604 , \15603 , \15302 );
and \U$14622 ( \15605 , \15602 , \15604 );
and \U$14623 ( \15606 , \15599 , \15605 );
and \U$14624 ( \15607 , \15581 , \15605 );
or \U$14625 ( \15608 , \15600 , \15606 , \15607 );
xor \U$14626 ( \15609 , \15271 , \15305 );
xor \U$14627 ( \15610 , \15609 , \15316 );
xor \U$14628 ( \15611 , \15321 , \15323 );
xor \U$14629 ( \15612 , \15611 , \15326 );
and \U$14630 ( \15613 , \15610 , \15612 );
xor \U$14631 ( \15614 , \15340 , \15342 );
xor \U$14632 ( \15615 , \15614 , \15344 );
and \U$14633 ( \15616 , \15612 , \15615 );
and \U$14634 ( \15617 , \15610 , \15615 );
or \U$14635 ( \15618 , \15613 , \15616 , \15617 );
and \U$14636 ( \15619 , \15608 , \15618 );
xor \U$14637 ( \15620 , \14883 , \15039 );
xor \U$14638 ( \15621 , \15620 , \15050 );
and \U$14639 ( \15622 , \15618 , \15621 );
and \U$14640 ( \15623 , \15608 , \15621 );
or \U$14641 ( \15624 , \15619 , \15622 , \15623 );
xor \U$14642 ( \15625 , \15319 , \15329 );
xor \U$14643 ( \15626 , \15625 , \15347 );
xor \U$14644 ( \15627 , \15352 , \15354 );
xor \U$14645 ( \15628 , \15627 , \15357 );
and \U$14646 ( \15629 , \15626 , \15628 );
and \U$14647 ( \15630 , \15624 , \15629 );
xor \U$14648 ( \15631 , \15053 , \15074 );
xor \U$14649 ( \15632 , \15631 , \15085 );
and \U$14650 ( \15633 , \15629 , \15632 );
and \U$14651 ( \15634 , \15624 , \15632 );
or \U$14652 ( \15635 , \15630 , \15633 , \15634 );
xor \U$14653 ( \15636 , \15366 , \15368 );
xor \U$14654 ( \15637 , \15636 , \15371 );
and \U$14655 ( \15638 , \15635 , \15637 );
and \U$14656 ( \15639 , \15380 , \15638 );
xor \U$14657 ( \15640 , \15380 , \15638 );
xor \U$14658 ( \15641 , \15635 , \15637 );
xor \U$14659 ( \15642 , \15624 , \15629 );
xor \U$14660 ( \15643 , \15642 , \15632 );
xor \U$14661 ( \15644 , \15350 , \15360 );
xor \U$14662 ( \15645 , \15644 , \15363 );
and \U$14663 ( \15646 , \15643 , \15645 );
and \U$14664 ( \15647 , \15641 , \15646 );
xor \U$14665 ( \15648 , \15641 , \15646 );
xor \U$14666 ( \15649 , \15643 , \15645 );
and \U$14667 ( \15650 , \3045 , \7906 );
and \U$14668 ( \15651 , \2901 , \7904 );
nor \U$14669 ( \15652 , \15650 , \15651 );
xnor \U$14670 ( \15653 , \15652 , \7646 );
and \U$14671 ( \15654 , \3334 , \7412 );
and \U$14672 ( \15655 , \3309 , \7410 );
nor \U$14673 ( \15656 , \15654 , \15655 );
xnor \U$14674 ( \15657 , \15656 , \7097 );
and \U$14675 ( \15658 , \15653 , \15657 );
and \U$14676 ( \15659 , \3675 , \6903 );
and \U$14677 ( \15660 , \3508 , \6901 );
nor \U$14678 ( \15661 , \15659 , \15660 );
xnor \U$14679 ( \15662 , \15661 , \6563 );
and \U$14680 ( \15663 , \15657 , \15662 );
and \U$14681 ( \15664 , \15653 , \15662 );
or \U$14682 ( \15665 , \15658 , \15663 , \15664 );
and \U$14683 ( \15666 , \1656 , \11482 );
and \U$14684 ( \15667 , \1593 , \11479 );
nor \U$14685 ( \15668 , \15666 , \15667 );
xnor \U$14686 ( \15669 , \15668 , \10427 );
and \U$14687 ( \15670 , \1942 , \10669 );
and \U$14688 ( \15671 , \1854 , \10667 );
nor \U$14689 ( \15672 , \15670 , \15671 );
xnor \U$14690 ( \15673 , \15672 , \10430 );
and \U$14691 ( \15674 , \15669 , \15673 );
and \U$14692 ( \15675 , \2052 , \10101 );
and \U$14693 ( \15676 , \2047 , \10099 );
nor \U$14694 ( \15677 , \15675 , \15676 );
xnor \U$14695 ( \15678 , \15677 , \9791 );
and \U$14696 ( \15679 , \15673 , \15678 );
and \U$14697 ( \15680 , \15669 , \15678 );
or \U$14698 ( \15681 , \15674 , \15679 , \15680 );
and \U$14699 ( \15682 , \15665 , \15681 );
and \U$14700 ( \15683 , \2283 , \9564 );
and \U$14701 ( \15684 , \2168 , \9562 );
nor \U$14702 ( \15685 , \15683 , \15684 );
xnor \U$14703 ( \15686 , \15685 , \9193 );
and \U$14704 ( \15687 , \2467 , \9002 );
and \U$14705 ( \15688 , \2459 , \9000 );
nor \U$14706 ( \15689 , \15687 , \15688 );
xnor \U$14707 ( \15690 , \15689 , \8684 );
and \U$14708 ( \15691 , \15686 , \15690 );
and \U$14709 ( \15692 , \2715 , \8435 );
and \U$14710 ( \15693 , \2710 , \8433 );
nor \U$14711 ( \15694 , \15692 , \15693 );
xnor \U$14712 ( \15695 , \15694 , \8186 );
and \U$14713 ( \15696 , \15690 , \15695 );
and \U$14714 ( \15697 , \15686 , \15695 );
or \U$14715 ( \15698 , \15691 , \15696 , \15697 );
and \U$14716 ( \15699 , \15681 , \15698 );
and \U$14717 ( \15700 , \15665 , \15698 );
or \U$14718 ( \15701 , \15682 , \15699 , \15700 );
and \U$14719 ( \15702 , \5137 , \5023 );
and \U$14720 ( \15703 , \4940 , \5021 );
nor \U$14721 ( \15704 , \15702 , \15703 );
xnor \U$14722 ( \15705 , \15704 , \4880 );
and \U$14723 ( \15706 , \5447 , \4700 );
and \U$14724 ( \15707 , \5439 , \4698 );
nor \U$14725 ( \15708 , \15706 , \15707 );
xnor \U$14726 ( \15709 , \15708 , \4454 );
and \U$14727 ( \15710 , \15705 , \15709 );
and \U$14728 ( \15711 , \5921 , \4305 );
and \U$14729 ( \15712 , \5916 , \4303 );
nor \U$14730 ( \15713 , \15711 , \15712 );
xnor \U$14731 ( \15714 , \15713 , \4118 );
and \U$14732 ( \15715 , \15709 , \15714 );
and \U$14733 ( \15716 , \15705 , \15714 );
or \U$14734 ( \15717 , \15710 , \15715 , \15716 );
and \U$14735 ( \15718 , \3932 , \6314 );
and \U$14736 ( \15719 , \3813 , \6312 );
nor \U$14737 ( \15720 , \15718 , \15719 );
xnor \U$14738 ( \15721 , \15720 , \6073 );
and \U$14739 ( \15722 , \4557 , \5848 );
and \U$14740 ( \15723 , \4349 , \5846 );
nor \U$14741 ( \15724 , \15722 , \15723 );
xnor \U$14742 ( \15725 , \15724 , \5660 );
and \U$14743 ( \15726 , \15721 , \15725 );
and \U$14744 ( \15727 , \4684 , \5474 );
and \U$14745 ( \15728 , \4679 , \5472 );
nor \U$14746 ( \15729 , \15727 , \15728 );
xnor \U$14747 ( \15730 , \15729 , \5242 );
and \U$14748 ( \15731 , \15725 , \15730 );
and \U$14749 ( \15732 , \15721 , \15730 );
or \U$14750 ( \15733 , \15726 , \15731 , \15732 );
and \U$14751 ( \15734 , \15717 , \15733 );
and \U$14752 ( \15735 , \6444 , \3992 );
and \U$14753 ( \15736 , \6185 , \3990 );
nor \U$14754 ( \15737 , \15735 , \15736 );
xnor \U$14755 ( \15738 , \15737 , \3787 );
and \U$14756 ( \15739 , \6825 , \3586 );
and \U$14757 ( \15740 , \6816 , \3584 );
nor \U$14758 ( \15741 , \15739 , \15740 );
xnor \U$14759 ( \15742 , \15741 , \3437 );
and \U$14760 ( \15743 , \15738 , \15742 );
and \U$14761 ( \15744 , \7370 , \3264 );
and \U$14762 ( \15745 , \7168 , \3262 );
nor \U$14763 ( \15746 , \15744 , \15745 );
xnor \U$14764 ( \15747 , \15746 , \3122 );
and \U$14765 ( \15748 , \15742 , \15747 );
and \U$14766 ( \15749 , \15738 , \15747 );
or \U$14767 ( \15750 , \15743 , \15748 , \15749 );
and \U$14768 ( \15751 , \15733 , \15750 );
and \U$14769 ( \15752 , \15717 , \15750 );
or \U$14770 ( \15753 , \15734 , \15751 , \15752 );
and \U$14771 ( \15754 , \15701 , \15753 );
and \U$14772 ( \15755 , \9649 , \2222 );
and \U$14773 ( \15756 , \9365 , \2220 );
nor \U$14774 ( \15757 , \15755 , \15756 );
xnor \U$14775 ( \15758 , \15757 , \2109 );
and \U$14776 ( \15759 , \10226 , \2028 );
and \U$14777 ( \15760 , \10218 , \2026 );
nor \U$14778 ( \15761 , \15759 , \15760 );
xnor \U$14779 ( \15762 , \15761 , \1892 );
and \U$14780 ( \15763 , \15758 , \15762 );
and \U$14781 ( \15764 , \10834 , \1828 );
and \U$14782 ( \15765 , \10829 , \1826 );
nor \U$14783 ( \15766 , \15764 , \15765 );
xnor \U$14784 ( \15767 , \15766 , \1750 );
and \U$14785 ( \15768 , \15762 , \15767 );
and \U$14786 ( \15769 , \15758 , \15767 );
or \U$14787 ( \15770 , \15763 , \15768 , \15769 );
and \U$14788 ( \15771 , \7845 , \2968 );
and \U$14789 ( \15772 , \7673 , \2966 );
nor \U$14790 ( \15773 , \15771 , \15772 );
xnor \U$14791 ( \15774 , \15773 , \2831 );
and \U$14792 ( \15775 , \8795 , \2762 );
and \U$14793 ( \15776 , \8371 , \2760 );
nor \U$14794 ( \15777 , \15775 , \15776 );
xnor \U$14795 ( \15778 , \15777 , \2610 );
and \U$14796 ( \15779 , \15774 , \15778 );
and \U$14797 ( \15780 , \9046 , \2494 );
and \U$14798 ( \15781 , \9041 , \2492 );
nor \U$14799 ( \15782 , \15780 , \15781 );
xnor \U$14800 ( \15783 , \15782 , \2338 );
and \U$14801 ( \15784 , \15778 , \15783 );
and \U$14802 ( \15785 , \15774 , \15783 );
or \U$14803 ( \15786 , \15779 , \15784 , \15785 );
and \U$14804 ( \15787 , \15770 , \15786 );
xor \U$14805 ( \15788 , \15501 , \15505 );
xor \U$14806 ( \15789 , \15788 , \15508 );
and \U$14807 ( \15790 , \15786 , \15789 );
and \U$14808 ( \15791 , \15770 , \15789 );
or \U$14809 ( \15792 , \15787 , \15790 , \15791 );
and \U$14810 ( \15793 , \15753 , \15792 );
and \U$14811 ( \15794 , \15701 , \15792 );
or \U$14812 ( \15795 , \15754 , \15793 , \15794 );
xor \U$14813 ( \15796 , \15485 , \15489 );
xor \U$14814 ( \15797 , \15796 , \15494 );
xor \U$14815 ( \15798 , \15417 , \15421 );
xor \U$14816 ( \15799 , \15798 , \15426 );
and \U$14817 ( \15800 , \15797 , \15799 );
xor \U$14818 ( \15801 , \15516 , \15520 );
xor \U$14819 ( \15802 , \15801 , \15525 );
and \U$14820 ( \15803 , \15799 , \15802 );
and \U$14821 ( \15804 , \15797 , \15802 );
or \U$14822 ( \15805 , \15800 , \15803 , \15804 );
xor \U$14823 ( \15806 , \15384 , \15388 );
xor \U$14824 ( \15807 , \15806 , \15393 );
xor \U$14825 ( \15808 , \15400 , \15404 );
xor \U$14826 ( \15809 , \15808 , \15409 );
and \U$14827 ( \15810 , \15807 , \15809 );
xor \U$14828 ( \15811 , \15436 , \15440 );
xor \U$14829 ( \15812 , \15811 , \15445 );
and \U$14830 ( \15813 , \15809 , \15812 );
and \U$14831 ( \15814 , \15807 , \15812 );
or \U$14832 ( \15815 , \15810 , \15813 , \15814 );
and \U$14833 ( \15816 , \15805 , \15815 );
xor \U$14834 ( \15817 , \15452 , \15456 );
xor \U$14835 ( \15818 , \15817 , \15461 );
xor \U$14836 ( \15819 , \15469 , \15473 );
xor \U$14837 ( \15820 , \15819 , \1422 );
and \U$14838 ( \15821 , \15818 , \15820 );
and \U$14839 ( \15822 , \15815 , \15821 );
and \U$14840 ( \15823 , \15805 , \15821 );
or \U$14841 ( \15824 , \15816 , \15822 , \15823 );
and \U$14842 ( \15825 , \15795 , \15824 );
xor \U$14843 ( \15826 , \15536 , \15538 );
xor \U$14844 ( \15827 , \15826 , \15541 );
xor \U$14845 ( \15828 , \15546 , \15548 );
xor \U$14846 ( \15829 , \15828 , \15551 );
and \U$14847 ( \15830 , \15827 , \15829 );
xor \U$14848 ( \15831 , \15557 , \15559 );
xor \U$14849 ( \15832 , \15831 , \15561 );
and \U$14850 ( \15833 , \15829 , \15832 );
and \U$14851 ( \15834 , \15827 , \15832 );
or \U$14852 ( \15835 , \15830 , \15833 , \15834 );
and \U$14853 ( \15836 , \15824 , \15835 );
and \U$14854 ( \15837 , \15795 , \15835 );
or \U$14855 ( \15838 , \15825 , \15836 , \15837 );
xor \U$14856 ( \15839 , \15396 , \15412 );
xor \U$14857 ( \15840 , \15839 , \15429 );
xor \U$14858 ( \15841 , \15448 , \15464 );
xor \U$14859 ( \15842 , \15841 , \15477 );
and \U$14860 ( \15843 , \15840 , \15842 );
xor \U$14861 ( \15844 , \15497 , \15511 );
xor \U$14862 ( \15845 , \15844 , \15528 );
and \U$14863 ( \15846 , \15842 , \15845 );
and \U$14864 ( \15847 , \15840 , \15845 );
or \U$14865 ( \15848 , \15843 , \15846 , \15847 );
xor \U$14866 ( \15849 , \15232 , \15248 );
xor \U$14867 ( \15850 , \15849 , \15265 );
and \U$14868 ( \15851 , \15848 , \15850 );
xor \U$14869 ( \15852 , \15583 , \15585 );
xor \U$14870 ( \15853 , \15852 , \15588 );
and \U$14871 ( \15854 , \15850 , \15853 );
and \U$14872 ( \15855 , \15848 , \15853 );
or \U$14873 ( \15856 , \15851 , \15854 , \15855 );
and \U$14874 ( \15857 , \15838 , \15856 );
xor \U$14875 ( \15858 , \15432 , \15480 );
xor \U$14876 ( \15859 , \15858 , \15531 );
xor \U$14877 ( \15860 , \15544 , \15554 );
xor \U$14878 ( \15861 , \15860 , \15564 );
and \U$14879 ( \15862 , \15859 , \15861 );
xor \U$14880 ( \15863 , \15570 , \15572 );
xor \U$14881 ( \15864 , \15863 , \15575 );
and \U$14882 ( \15865 , \15861 , \15864 );
and \U$14883 ( \15866 , \15859 , \15864 );
or \U$14884 ( \15867 , \15862 , \15865 , \15866 );
and \U$14885 ( \15868 , \15856 , \15867 );
and \U$14886 ( \15869 , \15838 , \15867 );
or \U$14887 ( \15870 , \15857 , \15868 , \15869 );
xor \U$14888 ( \15871 , \15534 , \15567 );
xor \U$14889 ( \15872 , \15871 , \15578 );
xor \U$14890 ( \15873 , \15591 , \15593 );
xor \U$14891 ( \15874 , \15873 , \15596 );
and \U$14892 ( \15875 , \15872 , \15874 );
xor \U$14893 ( \15876 , \15602 , \15604 );
and \U$14894 ( \15877 , \15874 , \15876 );
and \U$14895 ( \15878 , \15872 , \15876 );
or \U$14896 ( \15879 , \15875 , \15877 , \15878 );
and \U$14897 ( \15880 , \15870 , \15879 );
xor \U$14898 ( \15881 , \15610 , \15612 );
xor \U$14899 ( \15882 , \15881 , \15615 );
and \U$14900 ( \15883 , \15879 , \15882 );
and \U$14901 ( \15884 , \15870 , \15882 );
or \U$14902 ( \15885 , \15880 , \15883 , \15884 );
xor \U$14903 ( \15886 , \15608 , \15618 );
xor \U$14904 ( \15887 , \15886 , \15621 );
and \U$14905 ( \15888 , \15885 , \15887 );
xor \U$14906 ( \15889 , \15626 , \15628 );
and \U$14907 ( \15890 , \15887 , \15889 );
and \U$14908 ( \15891 , \15885 , \15889 );
or \U$14909 ( \15892 , \15888 , \15890 , \15891 );
and \U$14910 ( \15893 , \15649 , \15892 );
xor \U$14911 ( \15894 , \15649 , \15892 );
xor \U$14912 ( \15895 , \15885 , \15887 );
xor \U$14913 ( \15896 , \15895 , \15889 );
and \U$14914 ( \15897 , \2901 , \8435 );
and \U$14915 ( \15898 , \2715 , \8433 );
nor \U$14916 ( \15899 , \15897 , \15898 );
xnor \U$14917 ( \15900 , \15899 , \8186 );
and \U$14918 ( \15901 , \3309 , \7906 );
and \U$14919 ( \15902 , \3045 , \7904 );
nor \U$14920 ( \15903 , \15901 , \15902 );
xnor \U$14921 ( \15904 , \15903 , \7646 );
and \U$14922 ( \15905 , \15900 , \15904 );
and \U$14923 ( \15906 , \3508 , \7412 );
and \U$14924 ( \15907 , \3334 , \7410 );
nor \U$14925 ( \15908 , \15906 , \15907 );
xnor \U$14926 ( \15909 , \15908 , \7097 );
and \U$14927 ( \15910 , \15904 , \15909 );
and \U$14928 ( \15911 , \15900 , \15909 );
or \U$14929 ( \15912 , \15905 , \15910 , \15911 );
and \U$14930 ( \15913 , \2168 , \10101 );
and \U$14931 ( \15914 , \2052 , \10099 );
nor \U$14932 ( \15915 , \15913 , \15914 );
xnor \U$14933 ( \15916 , \15915 , \9791 );
and \U$14934 ( \15917 , \2459 , \9564 );
and \U$14935 ( \15918 , \2283 , \9562 );
nor \U$14936 ( \15919 , \15917 , \15918 );
xnor \U$14937 ( \15920 , \15919 , \9193 );
and \U$14938 ( \15921 , \15916 , \15920 );
and \U$14939 ( \15922 , \2710 , \9002 );
and \U$14940 ( \15923 , \2467 , \9000 );
nor \U$14941 ( \15924 , \15922 , \15923 );
xnor \U$14942 ( \15925 , \15924 , \8684 );
and \U$14943 ( \15926 , \15920 , \15925 );
and \U$14944 ( \15927 , \15916 , \15925 );
or \U$14945 ( \15928 , \15921 , \15926 , \15927 );
and \U$14946 ( \15929 , \15912 , \15928 );
and \U$14947 ( \15930 , \1854 , \11482 );
and \U$14948 ( \15931 , \1656 , \11479 );
nor \U$14949 ( \15932 , \15930 , \15931 );
xnor \U$14950 ( \15933 , \15932 , \10427 );
and \U$14951 ( \15934 , \2047 , \10669 );
and \U$14952 ( \15935 , \1942 , \10667 );
nor \U$14953 ( \15936 , \15934 , \15935 );
xnor \U$14954 ( \15937 , \15936 , \10430 );
and \U$14955 ( \15938 , \15933 , \15937 );
and \U$14956 ( \15939 , \15937 , \1570 );
and \U$14957 ( \15940 , \15933 , \1570 );
or \U$14958 ( \15941 , \15938 , \15939 , \15940 );
and \U$14959 ( \15942 , \15928 , \15941 );
and \U$14960 ( \15943 , \15912 , \15941 );
or \U$14961 ( \15944 , \15929 , \15942 , \15943 );
and \U$14962 ( \15945 , \7673 , \3264 );
and \U$14963 ( \15946 , \7370 , \3262 );
nor \U$14964 ( \15947 , \15945 , \15946 );
xnor \U$14965 ( \15948 , \15947 , \3122 );
and \U$14966 ( \15949 , \8371 , \2968 );
and \U$14967 ( \15950 , \7845 , \2966 );
nor \U$14968 ( \15951 , \15949 , \15950 );
xnor \U$14969 ( \15952 , \15951 , \2831 );
and \U$14970 ( \15953 , \15948 , \15952 );
and \U$14971 ( \15954 , \9041 , \2762 );
and \U$14972 ( \15955 , \8795 , \2760 );
nor \U$14973 ( \15956 , \15954 , \15955 );
xnor \U$14974 ( \15957 , \15956 , \2610 );
and \U$14975 ( \15958 , \15952 , \15957 );
and \U$14976 ( \15959 , \15948 , \15957 );
or \U$14977 ( \15960 , \15953 , \15958 , \15959 );
and \U$14978 ( \15961 , \9365 , \2494 );
and \U$14979 ( \15962 , \9046 , \2492 );
nor \U$14980 ( \15963 , \15961 , \15962 );
xnor \U$14981 ( \15964 , \15963 , \2338 );
and \U$14982 ( \15965 , \10218 , \2222 );
and \U$14983 ( \15966 , \9649 , \2220 );
nor \U$14984 ( \15967 , \15965 , \15966 );
xnor \U$14985 ( \15968 , \15967 , \2109 );
and \U$14986 ( \15969 , \15964 , \15968 );
and \U$14987 ( \15970 , \10829 , \2028 );
and \U$14988 ( \15971 , \10226 , \2026 );
nor \U$14989 ( \15972 , \15970 , \15971 );
xnor \U$14990 ( \15973 , \15972 , \1892 );
and \U$14991 ( \15974 , \15968 , \15973 );
and \U$14992 ( \15975 , \15964 , \15973 );
or \U$14993 ( \15976 , \15969 , \15974 , \15975 );
and \U$14994 ( \15977 , \15960 , \15976 );
and \U$14995 ( \15978 , \11635 , \1664 );
and \U$14996 ( \15979 , \11015 , \1662 );
nor \U$14997 ( \15980 , \15978 , \15979 );
xnor \U$14998 ( \15981 , \15980 , \1570 );
and \U$14999 ( \15982 , \15976 , \15981 );
and \U$15000 ( \15983 , \15960 , \15981 );
or \U$15001 ( \15984 , \15977 , \15982 , \15983 );
and \U$15002 ( \15985 , \15944 , \15984 );
and \U$15003 ( \15986 , \4940 , \5474 );
and \U$15004 ( \15987 , \4684 , \5472 );
nor \U$15005 ( \15988 , \15986 , \15987 );
xnor \U$15006 ( \15989 , \15988 , \5242 );
and \U$15007 ( \15990 , \5439 , \5023 );
and \U$15008 ( \15991 , \5137 , \5021 );
nor \U$15009 ( \15992 , \15990 , \15991 );
xnor \U$15010 ( \15993 , \15992 , \4880 );
and \U$15011 ( \15994 , \15989 , \15993 );
and \U$15012 ( \15995 , \5916 , \4700 );
and \U$15013 ( \15996 , \5447 , \4698 );
nor \U$15014 ( \15997 , \15995 , \15996 );
xnor \U$15015 ( \15998 , \15997 , \4454 );
and \U$15016 ( \15999 , \15993 , \15998 );
and \U$15017 ( \16000 , \15989 , \15998 );
or \U$15018 ( \16001 , \15994 , \15999 , \16000 );
and \U$15019 ( \16002 , \3813 , \6903 );
and \U$15020 ( \16003 , \3675 , \6901 );
nor \U$15021 ( \16004 , \16002 , \16003 );
xnor \U$15022 ( \16005 , \16004 , \6563 );
and \U$15023 ( \16006 , \4349 , \6314 );
and \U$15024 ( \16007 , \3932 , \6312 );
nor \U$15025 ( \16008 , \16006 , \16007 );
xnor \U$15026 ( \16009 , \16008 , \6073 );
and \U$15027 ( \16010 , \16005 , \16009 );
and \U$15028 ( \16011 , \4679 , \5848 );
and \U$15029 ( \16012 , \4557 , \5846 );
nor \U$15030 ( \16013 , \16011 , \16012 );
xnor \U$15031 ( \16014 , \16013 , \5660 );
and \U$15032 ( \16015 , \16009 , \16014 );
and \U$15033 ( \16016 , \16005 , \16014 );
or \U$15034 ( \16017 , \16010 , \16015 , \16016 );
and \U$15035 ( \16018 , \16001 , \16017 );
and \U$15036 ( \16019 , \6185 , \4305 );
and \U$15037 ( \16020 , \5921 , \4303 );
nor \U$15038 ( \16021 , \16019 , \16020 );
xnor \U$15039 ( \16022 , \16021 , \4118 );
and \U$15040 ( \16023 , \6816 , \3992 );
and \U$15041 ( \16024 , \6444 , \3990 );
nor \U$15042 ( \16025 , \16023 , \16024 );
xnor \U$15043 ( \16026 , \16025 , \3787 );
and \U$15044 ( \16027 , \16022 , \16026 );
and \U$15045 ( \16028 , \7168 , \3586 );
and \U$15046 ( \16029 , \6825 , \3584 );
nor \U$15047 ( \16030 , \16028 , \16029 );
xnor \U$15048 ( \16031 , \16030 , \3437 );
and \U$15049 ( \16032 , \16026 , \16031 );
and \U$15050 ( \16033 , \16022 , \16031 );
or \U$15051 ( \16034 , \16027 , \16032 , \16033 );
and \U$15052 ( \16035 , \16017 , \16034 );
and \U$15053 ( \16036 , \16001 , \16034 );
or \U$15054 ( \16037 , \16018 , \16035 , \16036 );
and \U$15055 ( \16038 , \15984 , \16037 );
and \U$15056 ( \16039 , \15944 , \16037 );
or \U$15057 ( \16040 , \15985 , \16038 , \16039 );
xor \U$15058 ( \16041 , \15758 , \15762 );
xor \U$15059 ( \16042 , \16041 , \15767 );
xor \U$15060 ( \16043 , \15738 , \15742 );
xor \U$15061 ( \16044 , \16043 , \15747 );
and \U$15062 ( \16045 , \16042 , \16044 );
xor \U$15063 ( \16046 , \15774 , \15778 );
xor \U$15064 ( \16047 , \16046 , \15783 );
and \U$15065 ( \16048 , \16044 , \16047 );
and \U$15066 ( \16049 , \16042 , \16047 );
or \U$15067 ( \16050 , \16045 , \16048 , \16049 );
xor \U$15068 ( \16051 , \15705 , \15709 );
xor \U$15069 ( \16052 , \16051 , \15714 );
xor \U$15070 ( \16053 , \15721 , \15725 );
xor \U$15071 ( \16054 , \16053 , \15730 );
and \U$15072 ( \16055 , \16052 , \16054 );
xor \U$15073 ( \16056 , \15653 , \15657 );
xor \U$15074 ( \16057 , \16056 , \15662 );
and \U$15075 ( \16058 , \16054 , \16057 );
and \U$15076 ( \16059 , \16052 , \16057 );
or \U$15077 ( \16060 , \16055 , \16058 , \16059 );
and \U$15078 ( \16061 , \16050 , \16060 );
xor \U$15079 ( \16062 , \15669 , \15673 );
xor \U$15080 ( \16063 , \16062 , \15678 );
xor \U$15081 ( \16064 , \15686 , \15690 );
xor \U$15082 ( \16065 , \16064 , \15695 );
and \U$15083 ( \16066 , \16063 , \16065 );
and \U$15084 ( \16067 , \16060 , \16066 );
and \U$15085 ( \16068 , \16050 , \16066 );
or \U$15086 ( \16069 , \16061 , \16067 , \16068 );
and \U$15087 ( \16070 , \16040 , \16069 );
xor \U$15088 ( \16071 , \15797 , \15799 );
xor \U$15089 ( \16072 , \16071 , \15802 );
xor \U$15090 ( \16073 , \15807 , \15809 );
xor \U$15091 ( \16074 , \16073 , \15812 );
and \U$15092 ( \16075 , \16072 , \16074 );
xor \U$15093 ( \16076 , \15818 , \15820 );
and \U$15094 ( \16077 , \16074 , \16076 );
and \U$15095 ( \16078 , \16072 , \16076 );
or \U$15096 ( \16079 , \16075 , \16077 , \16078 );
and \U$15097 ( \16080 , \16069 , \16079 );
and \U$15098 ( \16081 , \16040 , \16079 );
or \U$15099 ( \16082 , \16070 , \16080 , \16081 );
xor \U$15100 ( \16083 , \15665 , \15681 );
xor \U$15101 ( \16084 , \16083 , \15698 );
xor \U$15102 ( \16085 , \15717 , \15733 );
xor \U$15103 ( \16086 , \16085 , \15750 );
and \U$15104 ( \16087 , \16084 , \16086 );
xor \U$15105 ( \16088 , \15770 , \15786 );
xor \U$15106 ( \16089 , \16088 , \15789 );
and \U$15107 ( \16090 , \16086 , \16089 );
and \U$15108 ( \16091 , \16084 , \16089 );
or \U$15109 ( \16092 , \16087 , \16090 , \16091 );
xor \U$15110 ( \16093 , \15840 , \15842 );
xor \U$15111 ( \16094 , \16093 , \15845 );
and \U$15112 ( \16095 , \16092 , \16094 );
xor \U$15113 ( \16096 , \15827 , \15829 );
xor \U$15114 ( \16097 , \16096 , \15832 );
and \U$15115 ( \16098 , \16094 , \16097 );
and \U$15116 ( \16099 , \16092 , \16097 );
or \U$15117 ( \16100 , \16095 , \16098 , \16099 );
and \U$15118 ( \16101 , \16082 , \16100 );
xor \U$15119 ( \16102 , \15859 , \15861 );
xor \U$15120 ( \16103 , \16102 , \15864 );
and \U$15121 ( \16104 , \16100 , \16103 );
and \U$15122 ( \16105 , \16082 , \16103 );
or \U$15123 ( \16106 , \16101 , \16104 , \16105 );
xor \U$15124 ( \16107 , \15838 , \15856 );
xor \U$15125 ( \16108 , \16107 , \15867 );
and \U$15126 ( \16109 , \16106 , \16108 );
xor \U$15127 ( \16110 , \15872 , \15874 );
xor \U$15128 ( \16111 , \16110 , \15876 );
and \U$15129 ( \16112 , \16108 , \16111 );
and \U$15130 ( \16113 , \16106 , \16111 );
or \U$15131 ( \16114 , \16109 , \16112 , \16113 );
xor \U$15132 ( \16115 , \15581 , \15599 );
xor \U$15133 ( \16116 , \16115 , \15605 );
and \U$15134 ( \16117 , \16114 , \16116 );
xor \U$15135 ( \16118 , \15870 , \15879 );
xor \U$15136 ( \16119 , \16118 , \15882 );
and \U$15137 ( \16120 , \16116 , \16119 );
and \U$15138 ( \16121 , \16114 , \16119 );
or \U$15139 ( \16122 , \16117 , \16120 , \16121 );
and \U$15140 ( \16123 , \15896 , \16122 );
xor \U$15141 ( \16124 , \15896 , \16122 );
xor \U$15142 ( \16125 , \16114 , \16116 );
xor \U$15143 ( \16126 , \16125 , \16119 );
xor \U$15144 ( \16127 , \15900 , \15904 );
xor \U$15145 ( \16128 , \16127 , \15909 );
xor \U$15146 ( \16129 , \15916 , \15920 );
xor \U$15147 ( \16130 , \16129 , \15925 );
and \U$15148 ( \16131 , \16128 , \16130 );
xor \U$15149 ( \16132 , \15933 , \15937 );
xor \U$15150 ( \16133 , \16132 , \1570 );
and \U$15151 ( \16134 , \16130 , \16133 );
and \U$15152 ( \16135 , \16128 , \16133 );
or \U$15153 ( \16136 , \16131 , \16134 , \16135 );
nand \U$15154 ( \16137 , \11635 , \1662 );
xnor \U$15155 ( \16138 , \16137 , \1570 );
xor \U$15156 ( \16139 , \15948 , \15952 );
xor \U$15157 ( \16140 , \16139 , \15957 );
and \U$15158 ( \16141 , \16138 , \16140 );
xor \U$15159 ( \16142 , \15964 , \15968 );
xor \U$15160 ( \16143 , \16142 , \15973 );
and \U$15161 ( \16144 , \16140 , \16143 );
and \U$15162 ( \16145 , \16138 , \16143 );
or \U$15163 ( \16146 , \16141 , \16144 , \16145 );
and \U$15164 ( \16147 , \16136 , \16146 );
xor \U$15165 ( \16148 , \15989 , \15993 );
xor \U$15166 ( \16149 , \16148 , \15998 );
xor \U$15167 ( \16150 , \16005 , \16009 );
xor \U$15168 ( \16151 , \16150 , \16014 );
and \U$15169 ( \16152 , \16149 , \16151 );
xor \U$15170 ( \16153 , \16022 , \16026 );
xor \U$15171 ( \16154 , \16153 , \16031 );
and \U$15172 ( \16155 , \16151 , \16154 );
and \U$15173 ( \16156 , \16149 , \16154 );
or \U$15174 ( \16157 , \16152 , \16155 , \16156 );
and \U$15175 ( \16158 , \16146 , \16157 );
and \U$15176 ( \16159 , \16136 , \16157 );
or \U$15177 ( \16160 , \16147 , \16158 , \16159 );
and \U$15178 ( \16161 , \8795 , \2968 );
and \U$15179 ( \16162 , \8371 , \2966 );
nor \U$15180 ( \16163 , \16161 , \16162 );
xnor \U$15181 ( \16164 , \16163 , \2831 );
and \U$15182 ( \16165 , \9046 , \2762 );
and \U$15183 ( \16166 , \9041 , \2760 );
nor \U$15184 ( \16167 , \16165 , \16166 );
xnor \U$15185 ( \16168 , \16167 , \2610 );
and \U$15186 ( \16169 , \16164 , \16168 );
and \U$15187 ( \16170 , \9649 , \2494 );
and \U$15188 ( \16171 , \9365 , \2492 );
nor \U$15189 ( \16172 , \16170 , \16171 );
xnor \U$15190 ( \16173 , \16172 , \2338 );
and \U$15191 ( \16174 , \16168 , \16173 );
and \U$15192 ( \16175 , \16164 , \16173 );
or \U$15193 ( \16176 , \16169 , \16174 , \16175 );
and \U$15194 ( \16177 , \10226 , \2222 );
and \U$15195 ( \16178 , \10218 , \2220 );
nor \U$15196 ( \16179 , \16177 , \16178 );
xnor \U$15197 ( \16180 , \16179 , \2109 );
and \U$15198 ( \16181 , \10834 , \2028 );
and \U$15199 ( \16182 , \10829 , \2026 );
nor \U$15200 ( \16183 , \16181 , \16182 );
xnor \U$15201 ( \16184 , \16183 , \1892 );
and \U$15202 ( \16185 , \16180 , \16184 );
and \U$15203 ( \16186 , \11635 , \1828 );
and \U$15204 ( \16187 , \11015 , \1826 );
nor \U$15205 ( \16188 , \16186 , \16187 );
xnor \U$15206 ( \16189 , \16188 , \1750 );
and \U$15207 ( \16190 , \16184 , \16189 );
and \U$15208 ( \16191 , \16180 , \16189 );
or \U$15209 ( \16192 , \16185 , \16190 , \16191 );
and \U$15210 ( \16193 , \16176 , \16192 );
and \U$15211 ( \16194 , \11015 , \1828 );
and \U$15212 ( \16195 , \10834 , \1826 );
nor \U$15213 ( \16196 , \16194 , \16195 );
xnor \U$15214 ( \16197 , \16196 , \1750 );
and \U$15215 ( \16198 , \16192 , \16197 );
and \U$15216 ( \16199 , \16176 , \16197 );
or \U$15217 ( \16200 , \16193 , \16198 , \16199 );
and \U$15218 ( \16201 , \1942 , \11482 );
and \U$15219 ( \16202 , \1854 , \11479 );
nor \U$15220 ( \16203 , \16201 , \16202 );
xnor \U$15221 ( \16204 , \16203 , \10427 );
and \U$15222 ( \16205 , \2052 , \10669 );
and \U$15223 ( \16206 , \2047 , \10667 );
nor \U$15224 ( \16207 , \16205 , \16206 );
xnor \U$15225 ( \16208 , \16207 , \10430 );
and \U$15226 ( \16209 , \16204 , \16208 );
and \U$15227 ( \16210 , \2283 , \10101 );
and \U$15228 ( \16211 , \2168 , \10099 );
nor \U$15229 ( \16212 , \16210 , \16211 );
xnor \U$15230 ( \16213 , \16212 , \9791 );
and \U$15231 ( \16214 , \16208 , \16213 );
and \U$15232 ( \16215 , \16204 , \16213 );
or \U$15233 ( \16216 , \16209 , \16214 , \16215 );
and \U$15234 ( \16217 , \2467 , \9564 );
and \U$15235 ( \16218 , \2459 , \9562 );
nor \U$15236 ( \16219 , \16217 , \16218 );
xnor \U$15237 ( \16220 , \16219 , \9193 );
and \U$15238 ( \16221 , \2715 , \9002 );
and \U$15239 ( \16222 , \2710 , \9000 );
nor \U$15240 ( \16223 , \16221 , \16222 );
xnor \U$15241 ( \16224 , \16223 , \8684 );
and \U$15242 ( \16225 , \16220 , \16224 );
and \U$15243 ( \16226 , \3045 , \8435 );
and \U$15244 ( \16227 , \2901 , \8433 );
nor \U$15245 ( \16228 , \16226 , \16227 );
xnor \U$15246 ( \16229 , \16228 , \8186 );
and \U$15247 ( \16230 , \16224 , \16229 );
and \U$15248 ( \16231 , \16220 , \16229 );
or \U$15249 ( \16232 , \16225 , \16230 , \16231 );
and \U$15250 ( \16233 , \16216 , \16232 );
and \U$15251 ( \16234 , \3334 , \7906 );
and \U$15252 ( \16235 , \3309 , \7904 );
nor \U$15253 ( \16236 , \16234 , \16235 );
xnor \U$15254 ( \16237 , \16236 , \7646 );
and \U$15255 ( \16238 , \3675 , \7412 );
and \U$15256 ( \16239 , \3508 , \7410 );
nor \U$15257 ( \16240 , \16238 , \16239 );
xnor \U$15258 ( \16241 , \16240 , \7097 );
and \U$15259 ( \16242 , \16237 , \16241 );
and \U$15260 ( \16243 , \3932 , \6903 );
and \U$15261 ( \16244 , \3813 , \6901 );
nor \U$15262 ( \16245 , \16243 , \16244 );
xnor \U$15263 ( \16246 , \16245 , \6563 );
and \U$15264 ( \16247 , \16241 , \16246 );
and \U$15265 ( \16248 , \16237 , \16246 );
or \U$15266 ( \16249 , \16242 , \16247 , \16248 );
and \U$15267 ( \16250 , \16232 , \16249 );
and \U$15268 ( \16251 , \16216 , \16249 );
or \U$15269 ( \16252 , \16233 , \16250 , \16251 );
and \U$15270 ( \16253 , \16200 , \16252 );
and \U$15271 ( \16254 , \5447 , \5023 );
and \U$15272 ( \16255 , \5439 , \5021 );
nor \U$15273 ( \16256 , \16254 , \16255 );
xnor \U$15274 ( \16257 , \16256 , \4880 );
and \U$15275 ( \16258 , \5921 , \4700 );
and \U$15276 ( \16259 , \5916 , \4698 );
nor \U$15277 ( \16260 , \16258 , \16259 );
xnor \U$15278 ( \16261 , \16260 , \4454 );
and \U$15279 ( \16262 , \16257 , \16261 );
and \U$15280 ( \16263 , \6444 , \4305 );
and \U$15281 ( \16264 , \6185 , \4303 );
nor \U$15282 ( \16265 , \16263 , \16264 );
xnor \U$15283 ( \16266 , \16265 , \4118 );
and \U$15284 ( \16267 , \16261 , \16266 );
and \U$15285 ( \16268 , \16257 , \16266 );
or \U$15286 ( \16269 , \16262 , \16267 , \16268 );
and \U$15287 ( \16270 , \6825 , \3992 );
and \U$15288 ( \16271 , \6816 , \3990 );
nor \U$15289 ( \16272 , \16270 , \16271 );
xnor \U$15290 ( \16273 , \16272 , \3787 );
and \U$15291 ( \16274 , \7370 , \3586 );
and \U$15292 ( \16275 , \7168 , \3584 );
nor \U$15293 ( \16276 , \16274 , \16275 );
xnor \U$15294 ( \16277 , \16276 , \3437 );
and \U$15295 ( \16278 , \16273 , \16277 );
and \U$15296 ( \16279 , \7845 , \3264 );
and \U$15297 ( \16280 , \7673 , \3262 );
nor \U$15298 ( \16281 , \16279 , \16280 );
xnor \U$15299 ( \16282 , \16281 , \3122 );
and \U$15300 ( \16283 , \16277 , \16282 );
and \U$15301 ( \16284 , \16273 , \16282 );
or \U$15302 ( \16285 , \16278 , \16283 , \16284 );
and \U$15303 ( \16286 , \16269 , \16285 );
and \U$15304 ( \16287 , \4557 , \6314 );
and \U$15305 ( \16288 , \4349 , \6312 );
nor \U$15306 ( \16289 , \16287 , \16288 );
xnor \U$15307 ( \16290 , \16289 , \6073 );
and \U$15308 ( \16291 , \4684 , \5848 );
and \U$15309 ( \16292 , \4679 , \5846 );
nor \U$15310 ( \16293 , \16291 , \16292 );
xnor \U$15311 ( \16294 , \16293 , \5660 );
and \U$15312 ( \16295 , \16290 , \16294 );
and \U$15313 ( \16296 , \5137 , \5474 );
and \U$15314 ( \16297 , \4940 , \5472 );
nor \U$15315 ( \16298 , \16296 , \16297 );
xnor \U$15316 ( \16299 , \16298 , \5242 );
and \U$15317 ( \16300 , \16294 , \16299 );
and \U$15318 ( \16301 , \16290 , \16299 );
or \U$15319 ( \16302 , \16295 , \16300 , \16301 );
and \U$15320 ( \16303 , \16285 , \16302 );
and \U$15321 ( \16304 , \16269 , \16302 );
or \U$15322 ( \16305 , \16286 , \16303 , \16304 );
and \U$15323 ( \16306 , \16252 , \16305 );
and \U$15324 ( \16307 , \16200 , \16305 );
or \U$15325 ( \16308 , \16253 , \16306 , \16307 );
and \U$15326 ( \16309 , \16160 , \16308 );
xor \U$15327 ( \16310 , \16042 , \16044 );
xor \U$15328 ( \16311 , \16310 , \16047 );
xor \U$15329 ( \16312 , \16052 , \16054 );
xor \U$15330 ( \16313 , \16312 , \16057 );
and \U$15331 ( \16314 , \16311 , \16313 );
xor \U$15332 ( \16315 , \16063 , \16065 );
and \U$15333 ( \16316 , \16313 , \16315 );
and \U$15334 ( \16317 , \16311 , \16315 );
or \U$15335 ( \16318 , \16314 , \16316 , \16317 );
and \U$15336 ( \16319 , \16308 , \16318 );
and \U$15337 ( \16320 , \16160 , \16318 );
or \U$15338 ( \16321 , \16309 , \16319 , \16320 );
xor \U$15339 ( \16322 , \15912 , \15928 );
xor \U$15340 ( \16323 , \16322 , \15941 );
xor \U$15341 ( \16324 , \15960 , \15976 );
xor \U$15342 ( \16325 , \16324 , \15981 );
and \U$15343 ( \16326 , \16323 , \16325 );
xor \U$15344 ( \16327 , \16001 , \16017 );
xor \U$15345 ( \16328 , \16327 , \16034 );
and \U$15346 ( \16329 , \16325 , \16328 );
and \U$15347 ( \16330 , \16323 , \16328 );
or \U$15348 ( \16331 , \16326 , \16329 , \16330 );
xor \U$15349 ( \16332 , \16084 , \16086 );
xor \U$15350 ( \16333 , \16332 , \16089 );
and \U$15351 ( \16334 , \16331 , \16333 );
xor \U$15352 ( \16335 , \16072 , \16074 );
xor \U$15353 ( \16336 , \16335 , \16076 );
and \U$15354 ( \16337 , \16333 , \16336 );
and \U$15355 ( \16338 , \16331 , \16336 );
or \U$15356 ( \16339 , \16334 , \16337 , \16338 );
and \U$15357 ( \16340 , \16321 , \16339 );
xor \U$15358 ( \16341 , \15805 , \15815 );
xor \U$15359 ( \16342 , \16341 , \15821 );
and \U$15360 ( \16343 , \16339 , \16342 );
and \U$15361 ( \16344 , \16321 , \16342 );
or \U$15362 ( \16345 , \16340 , \16343 , \16344 );
xor \U$15363 ( \16346 , \15701 , \15753 );
xor \U$15364 ( \16347 , \16346 , \15792 );
xor \U$15365 ( \16348 , \16040 , \16069 );
xor \U$15366 ( \16349 , \16348 , \16079 );
and \U$15367 ( \16350 , \16347 , \16349 );
xor \U$15368 ( \16351 , \16092 , \16094 );
xor \U$15369 ( \16352 , \16351 , \16097 );
and \U$15370 ( \16353 , \16349 , \16352 );
and \U$15371 ( \16354 , \16347 , \16352 );
or \U$15372 ( \16355 , \16350 , \16353 , \16354 );
and \U$15373 ( \16356 , \16345 , \16355 );
xor \U$15374 ( \16357 , \15848 , \15850 );
xor \U$15375 ( \16358 , \16357 , \15853 );
and \U$15376 ( \16359 , \16355 , \16358 );
and \U$15377 ( \16360 , \16345 , \16358 );
or \U$15378 ( \16361 , \16356 , \16359 , \16360 );
xor \U$15379 ( \16362 , \15795 , \15824 );
xor \U$15380 ( \16363 , \16362 , \15835 );
xor \U$15381 ( \16364 , \16082 , \16100 );
xor \U$15382 ( \16365 , \16364 , \16103 );
and \U$15383 ( \16366 , \16363 , \16365 );
and \U$15384 ( \16367 , \16361 , \16366 );
xor \U$15385 ( \16368 , \16106 , \16108 );
xor \U$15386 ( \16369 , \16368 , \16111 );
and \U$15387 ( \16370 , \16366 , \16369 );
and \U$15388 ( \16371 , \16361 , \16369 );
or \U$15389 ( \16372 , \16367 , \16370 , \16371 );
and \U$15390 ( \16373 , \16126 , \16372 );
xor \U$15391 ( \16374 , \16126 , \16372 );
xor \U$15392 ( \16375 , \16361 , \16366 );
xor \U$15393 ( \16376 , \16375 , \16369 );
and \U$15394 ( \16377 , \6816 , \4305 );
and \U$15395 ( \16378 , \6444 , \4303 );
nor \U$15396 ( \16379 , \16377 , \16378 );
xnor \U$15397 ( \16380 , \16379 , \4118 );
and \U$15398 ( \16381 , \7168 , \3992 );
and \U$15399 ( \16382 , \6825 , \3990 );
nor \U$15400 ( \16383 , \16381 , \16382 );
xnor \U$15401 ( \16384 , \16383 , \3787 );
and \U$15402 ( \16385 , \16380 , \16384 );
and \U$15403 ( \16386 , \7673 , \3586 );
and \U$15404 ( \16387 , \7370 , \3584 );
nor \U$15405 ( \16388 , \16386 , \16387 );
xnor \U$15406 ( \16389 , \16388 , \3437 );
and \U$15407 ( \16390 , \16384 , \16389 );
and \U$15408 ( \16391 , \16380 , \16389 );
or \U$15409 ( \16392 , \16385 , \16390 , \16391 );
and \U$15410 ( \16393 , \5439 , \5474 );
and \U$15411 ( \16394 , \5137 , \5472 );
nor \U$15412 ( \16395 , \16393 , \16394 );
xnor \U$15413 ( \16396 , \16395 , \5242 );
and \U$15414 ( \16397 , \5916 , \5023 );
and \U$15415 ( \16398 , \5447 , \5021 );
nor \U$15416 ( \16399 , \16397 , \16398 );
xnor \U$15417 ( \16400 , \16399 , \4880 );
and \U$15418 ( \16401 , \16396 , \16400 );
and \U$15419 ( \16402 , \6185 , \4700 );
and \U$15420 ( \16403 , \5921 , \4698 );
nor \U$15421 ( \16404 , \16402 , \16403 );
xnor \U$15422 ( \16405 , \16404 , \4454 );
and \U$15423 ( \16406 , \16400 , \16405 );
and \U$15424 ( \16407 , \16396 , \16405 );
or \U$15425 ( \16408 , \16401 , \16406 , \16407 );
and \U$15426 ( \16409 , \16392 , \16408 );
and \U$15427 ( \16410 , \4349 , \6903 );
and \U$15428 ( \16411 , \3932 , \6901 );
nor \U$15429 ( \16412 , \16410 , \16411 );
xnor \U$15430 ( \16413 , \16412 , \6563 );
and \U$15431 ( \16414 , \4679 , \6314 );
and \U$15432 ( \16415 , \4557 , \6312 );
nor \U$15433 ( \16416 , \16414 , \16415 );
xnor \U$15434 ( \16417 , \16416 , \6073 );
and \U$15435 ( \16418 , \16413 , \16417 );
and \U$15436 ( \16419 , \4940 , \5848 );
and \U$15437 ( \16420 , \4684 , \5846 );
nor \U$15438 ( \16421 , \16419 , \16420 );
xnor \U$15439 ( \16422 , \16421 , \5660 );
and \U$15440 ( \16423 , \16417 , \16422 );
and \U$15441 ( \16424 , \16413 , \16422 );
or \U$15442 ( \16425 , \16418 , \16423 , \16424 );
and \U$15443 ( \16426 , \16408 , \16425 );
and \U$15444 ( \16427 , \16392 , \16425 );
or \U$15445 ( \16428 , \16409 , \16426 , \16427 );
and \U$15446 ( \16429 , \2459 , \10101 );
and \U$15447 ( \16430 , \2283 , \10099 );
nor \U$15448 ( \16431 , \16429 , \16430 );
xnor \U$15449 ( \16432 , \16431 , \9791 );
and \U$15450 ( \16433 , \2710 , \9564 );
and \U$15451 ( \16434 , \2467 , \9562 );
nor \U$15452 ( \16435 , \16433 , \16434 );
xnor \U$15453 ( \16436 , \16435 , \9193 );
and \U$15454 ( \16437 , \16432 , \16436 );
and \U$15455 ( \16438 , \2901 , \9002 );
and \U$15456 ( \16439 , \2715 , \9000 );
nor \U$15457 ( \16440 , \16438 , \16439 );
xnor \U$15458 ( \16441 , \16440 , \8684 );
and \U$15459 ( \16442 , \16436 , \16441 );
and \U$15460 ( \16443 , \16432 , \16441 );
or \U$15461 ( \16444 , \16437 , \16442 , \16443 );
and \U$15462 ( \16445 , \2047 , \11482 );
and \U$15463 ( \16446 , \1942 , \11479 );
nor \U$15464 ( \16447 , \16445 , \16446 );
xnor \U$15465 ( \16448 , \16447 , \10427 );
and \U$15466 ( \16449 , \2168 , \10669 );
and \U$15467 ( \16450 , \2052 , \10667 );
nor \U$15468 ( \16451 , \16449 , \16450 );
xnor \U$15469 ( \16452 , \16451 , \10430 );
and \U$15470 ( \16453 , \16448 , \16452 );
and \U$15471 ( \16454 , \16452 , \1750 );
and \U$15472 ( \16455 , \16448 , \1750 );
or \U$15473 ( \16456 , \16453 , \16454 , \16455 );
and \U$15474 ( \16457 , \16444 , \16456 );
and \U$15475 ( \16458 , \3309 , \8435 );
and \U$15476 ( \16459 , \3045 , \8433 );
nor \U$15477 ( \16460 , \16458 , \16459 );
xnor \U$15478 ( \16461 , \16460 , \8186 );
and \U$15479 ( \16462 , \3508 , \7906 );
and \U$15480 ( \16463 , \3334 , \7904 );
nor \U$15481 ( \16464 , \16462 , \16463 );
xnor \U$15482 ( \16465 , \16464 , \7646 );
and \U$15483 ( \16466 , \16461 , \16465 );
and \U$15484 ( \16467 , \3813 , \7412 );
and \U$15485 ( \16468 , \3675 , \7410 );
nor \U$15486 ( \16469 , \16467 , \16468 );
xnor \U$15487 ( \16470 , \16469 , \7097 );
and \U$15488 ( \16471 , \16465 , \16470 );
and \U$15489 ( \16472 , \16461 , \16470 );
or \U$15490 ( \16473 , \16466 , \16471 , \16472 );
and \U$15491 ( \16474 , \16456 , \16473 );
and \U$15492 ( \16475 , \16444 , \16473 );
or \U$15493 ( \16476 , \16457 , \16474 , \16475 );
and \U$15494 ( \16477 , \16428 , \16476 );
and \U$15495 ( \16478 , \8371 , \3264 );
and \U$15496 ( \16479 , \7845 , \3262 );
nor \U$15497 ( \16480 , \16478 , \16479 );
xnor \U$15498 ( \16481 , \16480 , \3122 );
and \U$15499 ( \16482 , \9041 , \2968 );
and \U$15500 ( \16483 , \8795 , \2966 );
nor \U$15501 ( \16484 , \16482 , \16483 );
xnor \U$15502 ( \16485 , \16484 , \2831 );
and \U$15503 ( \16486 , \16481 , \16485 );
and \U$15504 ( \16487 , \9365 , \2762 );
and \U$15505 ( \16488 , \9046 , \2760 );
nor \U$15506 ( \16489 , \16487 , \16488 );
xnor \U$15507 ( \16490 , \16489 , \2610 );
and \U$15508 ( \16491 , \16485 , \16490 );
and \U$15509 ( \16492 , \16481 , \16490 );
or \U$15510 ( \16493 , \16486 , \16491 , \16492 );
and \U$15511 ( \16494 , \10218 , \2494 );
and \U$15512 ( \16495 , \9649 , \2492 );
nor \U$15513 ( \16496 , \16494 , \16495 );
xnor \U$15514 ( \16497 , \16496 , \2338 );
and \U$15515 ( \16498 , \10829 , \2222 );
and \U$15516 ( \16499 , \10226 , \2220 );
nor \U$15517 ( \16500 , \16498 , \16499 );
xnor \U$15518 ( \16501 , \16500 , \2109 );
and \U$15519 ( \16502 , \16497 , \16501 );
and \U$15520 ( \16503 , \11015 , \2028 );
and \U$15521 ( \16504 , \10834 , \2026 );
nor \U$15522 ( \16505 , \16503 , \16504 );
xnor \U$15523 ( \16506 , \16505 , \1892 );
and \U$15524 ( \16507 , \16501 , \16506 );
and \U$15525 ( \16508 , \16497 , \16506 );
or \U$15526 ( \16509 , \16502 , \16507 , \16508 );
and \U$15527 ( \16510 , \16493 , \16509 );
xor \U$15528 ( \16511 , \16180 , \16184 );
xor \U$15529 ( \16512 , \16511 , \16189 );
and \U$15530 ( \16513 , \16509 , \16512 );
and \U$15531 ( \16514 , \16493 , \16512 );
or \U$15532 ( \16515 , \16510 , \16513 , \16514 );
and \U$15533 ( \16516 , \16476 , \16515 );
and \U$15534 ( \16517 , \16428 , \16515 );
or \U$15535 ( \16518 , \16477 , \16516 , \16517 );
xor \U$15536 ( \16519 , \16164 , \16168 );
xor \U$15537 ( \16520 , \16519 , \16173 );
xor \U$15538 ( \16521 , \16257 , \16261 );
xor \U$15539 ( \16522 , \16521 , \16266 );
and \U$15540 ( \16523 , \16520 , \16522 );
xor \U$15541 ( \16524 , \16273 , \16277 );
xor \U$15542 ( \16525 , \16524 , \16282 );
and \U$15543 ( \16526 , \16522 , \16525 );
and \U$15544 ( \16527 , \16520 , \16525 );
or \U$15545 ( \16528 , \16523 , \16526 , \16527 );
xor \U$15546 ( \16529 , \16220 , \16224 );
xor \U$15547 ( \16530 , \16529 , \16229 );
xor \U$15548 ( \16531 , \16290 , \16294 );
xor \U$15549 ( \16532 , \16531 , \16299 );
and \U$15550 ( \16533 , \16530 , \16532 );
xor \U$15551 ( \16534 , \16237 , \16241 );
xor \U$15552 ( \16535 , \16534 , \16246 );
and \U$15553 ( \16536 , \16532 , \16535 );
and \U$15554 ( \16537 , \16530 , \16535 );
or \U$15555 ( \16538 , \16533 , \16536 , \16537 );
and \U$15556 ( \16539 , \16528 , \16538 );
xor \U$15557 ( \16540 , \16128 , \16130 );
xor \U$15558 ( \16541 , \16540 , \16133 );
and \U$15559 ( \16542 , \16538 , \16541 );
and \U$15560 ( \16543 , \16528 , \16541 );
or \U$15561 ( \16544 , \16539 , \16542 , \16543 );
and \U$15562 ( \16545 , \16518 , \16544 );
xor \U$15563 ( \16546 , \16176 , \16192 );
xor \U$15564 ( \16547 , \16546 , \16197 );
xor \U$15565 ( \16548 , \16138 , \16140 );
xor \U$15566 ( \16549 , \16548 , \16143 );
and \U$15567 ( \16550 , \16547 , \16549 );
xor \U$15568 ( \16551 , \16149 , \16151 );
xor \U$15569 ( \16552 , \16551 , \16154 );
and \U$15570 ( \16553 , \16549 , \16552 );
and \U$15571 ( \16554 , \16547 , \16552 );
or \U$15572 ( \16555 , \16550 , \16553 , \16554 );
and \U$15573 ( \16556 , \16544 , \16555 );
and \U$15574 ( \16557 , \16518 , \16555 );
or \U$15575 ( \16558 , \16545 , \16556 , \16557 );
xor \U$15576 ( \16559 , \16136 , \16146 );
xor \U$15577 ( \16560 , \16559 , \16157 );
xor \U$15578 ( \16561 , \16323 , \16325 );
xor \U$15579 ( \16562 , \16561 , \16328 );
and \U$15580 ( \16563 , \16560 , \16562 );
xor \U$15581 ( \16564 , \16311 , \16313 );
xor \U$15582 ( \16565 , \16564 , \16315 );
and \U$15583 ( \16566 , \16562 , \16565 );
and \U$15584 ( \16567 , \16560 , \16565 );
or \U$15585 ( \16568 , \16563 , \16566 , \16567 );
and \U$15586 ( \16569 , \16558 , \16568 );
xor \U$15587 ( \16570 , \16050 , \16060 );
xor \U$15588 ( \16571 , \16570 , \16066 );
and \U$15589 ( \16572 , \16568 , \16571 );
and \U$15590 ( \16573 , \16558 , \16571 );
or \U$15591 ( \16574 , \16569 , \16572 , \16573 );
xor \U$15592 ( \16575 , \15944 , \15984 );
xor \U$15593 ( \16576 , \16575 , \16037 );
xor \U$15594 ( \16577 , \16160 , \16308 );
xor \U$15595 ( \16578 , \16577 , \16318 );
and \U$15596 ( \16579 , \16576 , \16578 );
xor \U$15597 ( \16580 , \16331 , \16333 );
xor \U$15598 ( \16581 , \16580 , \16336 );
and \U$15599 ( \16582 , \16578 , \16581 );
and \U$15600 ( \16583 , \16576 , \16581 );
or \U$15601 ( \16584 , \16579 , \16582 , \16583 );
and \U$15602 ( \16585 , \16574 , \16584 );
xor \U$15603 ( \16586 , \16347 , \16349 );
xor \U$15604 ( \16587 , \16586 , \16352 );
and \U$15605 ( \16588 , \16584 , \16587 );
and \U$15606 ( \16589 , \16574 , \16587 );
or \U$15607 ( \16590 , \16585 , \16588 , \16589 );
xor \U$15608 ( \16591 , \16345 , \16355 );
xor \U$15609 ( \16592 , \16591 , \16358 );
and \U$15610 ( \16593 , \16590 , \16592 );
xor \U$15611 ( \16594 , \16363 , \16365 );
and \U$15612 ( \16595 , \16592 , \16594 );
and \U$15613 ( \16596 , \16590 , \16594 );
or \U$15614 ( \16597 , \16593 , \16595 , \16596 );
and \U$15615 ( \16598 , \16376 , \16597 );
xor \U$15616 ( \16599 , \16376 , \16597 );
xor \U$15617 ( \16600 , \16590 , \16592 );
xor \U$15618 ( \16601 , \16600 , \16594 );
and \U$15619 ( \16602 , \4684 , \6314 );
and \U$15620 ( \16603 , \4679 , \6312 );
nor \U$15621 ( \16604 , \16602 , \16603 );
xnor \U$15622 ( \16605 , \16604 , \6073 );
and \U$15623 ( \16606 , \5137 , \5848 );
and \U$15624 ( \16607 , \4940 , \5846 );
nor \U$15625 ( \16608 , \16606 , \16607 );
xnor \U$15626 ( \16609 , \16608 , \5660 );
and \U$15627 ( \16610 , \16605 , \16609 );
and \U$15628 ( \16611 , \5447 , \5474 );
and \U$15629 ( \16612 , \5439 , \5472 );
nor \U$15630 ( \16613 , \16611 , \16612 );
xnor \U$15631 ( \16614 , \16613 , \5242 );
and \U$15632 ( \16615 , \16609 , \16614 );
and \U$15633 ( \16616 , \16605 , \16614 );
or \U$15634 ( \16617 , \16610 , \16615 , \16616 );
and \U$15635 ( \16618 , \5921 , \5023 );
and \U$15636 ( \16619 , \5916 , \5021 );
nor \U$15637 ( \16620 , \16618 , \16619 );
xnor \U$15638 ( \16621 , \16620 , \4880 );
and \U$15639 ( \16622 , \6444 , \4700 );
and \U$15640 ( \16623 , \6185 , \4698 );
nor \U$15641 ( \16624 , \16622 , \16623 );
xnor \U$15642 ( \16625 , \16624 , \4454 );
and \U$15643 ( \16626 , \16621 , \16625 );
and \U$15644 ( \16627 , \6825 , \4305 );
and \U$15645 ( \16628 , \6816 , \4303 );
nor \U$15646 ( \16629 , \16627 , \16628 );
xnor \U$15647 ( \16630 , \16629 , \4118 );
and \U$15648 ( \16631 , \16625 , \16630 );
and \U$15649 ( \16632 , \16621 , \16630 );
or \U$15650 ( \16633 , \16626 , \16631 , \16632 );
and \U$15651 ( \16634 , \16617 , \16633 );
and \U$15652 ( \16635 , \7370 , \3992 );
and \U$15653 ( \16636 , \7168 , \3990 );
nor \U$15654 ( \16637 , \16635 , \16636 );
xnor \U$15655 ( \16638 , \16637 , \3787 );
and \U$15656 ( \16639 , \7845 , \3586 );
and \U$15657 ( \16640 , \7673 , \3584 );
nor \U$15658 ( \16641 , \16639 , \16640 );
xnor \U$15659 ( \16642 , \16641 , \3437 );
and \U$15660 ( \16643 , \16638 , \16642 );
and \U$15661 ( \16644 , \8795 , \3264 );
and \U$15662 ( \16645 , \8371 , \3262 );
nor \U$15663 ( \16646 , \16644 , \16645 );
xnor \U$15664 ( \16647 , \16646 , \3122 );
and \U$15665 ( \16648 , \16642 , \16647 );
and \U$15666 ( \16649 , \16638 , \16647 );
or \U$15667 ( \16650 , \16643 , \16648 , \16649 );
and \U$15668 ( \16651 , \16633 , \16650 );
and \U$15669 ( \16652 , \16617 , \16650 );
or \U$15670 ( \16653 , \16634 , \16651 , \16652 );
and \U$15671 ( \16654 , \2715 , \9564 );
and \U$15672 ( \16655 , \2710 , \9562 );
nor \U$15673 ( \16656 , \16654 , \16655 );
xnor \U$15674 ( \16657 , \16656 , \9193 );
and \U$15675 ( \16658 , \3045 , \9002 );
and \U$15676 ( \16659 , \2901 , \9000 );
nor \U$15677 ( \16660 , \16658 , \16659 );
xnor \U$15678 ( \16661 , \16660 , \8684 );
and \U$15679 ( \16662 , \16657 , \16661 );
and \U$15680 ( \16663 , \3334 , \8435 );
and \U$15681 ( \16664 , \3309 , \8433 );
nor \U$15682 ( \16665 , \16663 , \16664 );
xnor \U$15683 ( \16666 , \16665 , \8186 );
and \U$15684 ( \16667 , \16661 , \16666 );
and \U$15685 ( \16668 , \16657 , \16666 );
or \U$15686 ( \16669 , \16662 , \16667 , \16668 );
and \U$15687 ( \16670 , \3675 , \7906 );
and \U$15688 ( \16671 , \3508 , \7904 );
nor \U$15689 ( \16672 , \16670 , \16671 );
xnor \U$15690 ( \16673 , \16672 , \7646 );
and \U$15691 ( \16674 , \3932 , \7412 );
and \U$15692 ( \16675 , \3813 , \7410 );
nor \U$15693 ( \16676 , \16674 , \16675 );
xnor \U$15694 ( \16677 , \16676 , \7097 );
and \U$15695 ( \16678 , \16673 , \16677 );
and \U$15696 ( \16679 , \4557 , \6903 );
and \U$15697 ( \16680 , \4349 , \6901 );
nor \U$15698 ( \16681 , \16679 , \16680 );
xnor \U$15699 ( \16682 , \16681 , \6563 );
and \U$15700 ( \16683 , \16677 , \16682 );
and \U$15701 ( \16684 , \16673 , \16682 );
or \U$15702 ( \16685 , \16678 , \16683 , \16684 );
and \U$15703 ( \16686 , \16669 , \16685 );
and \U$15704 ( \16687 , \2052 , \11482 );
and \U$15705 ( \16688 , \2047 , \11479 );
nor \U$15706 ( \16689 , \16687 , \16688 );
xnor \U$15707 ( \16690 , \16689 , \10427 );
and \U$15708 ( \16691 , \2283 , \10669 );
and \U$15709 ( \16692 , \2168 , \10667 );
nor \U$15710 ( \16693 , \16691 , \16692 );
xnor \U$15711 ( \16694 , \16693 , \10430 );
and \U$15712 ( \16695 , \16690 , \16694 );
and \U$15713 ( \16696 , \2467 , \10101 );
and \U$15714 ( \16697 , \2459 , \10099 );
nor \U$15715 ( \16698 , \16696 , \16697 );
xnor \U$15716 ( \16699 , \16698 , \9791 );
and \U$15717 ( \16700 , \16694 , \16699 );
and \U$15718 ( \16701 , \16690 , \16699 );
or \U$15719 ( \16702 , \16695 , \16700 , \16701 );
and \U$15720 ( \16703 , \16685 , \16702 );
and \U$15721 ( \16704 , \16669 , \16702 );
or \U$15722 ( \16705 , \16686 , \16703 , \16704 );
and \U$15723 ( \16706 , \16653 , \16705 );
and \U$15724 ( \16707 , \9046 , \2968 );
and \U$15725 ( \16708 , \9041 , \2966 );
nor \U$15726 ( \16709 , \16707 , \16708 );
xnor \U$15727 ( \16710 , \16709 , \2831 );
and \U$15728 ( \16711 , \9649 , \2762 );
and \U$15729 ( \16712 , \9365 , \2760 );
nor \U$15730 ( \16713 , \16711 , \16712 );
xnor \U$15731 ( \16714 , \16713 , \2610 );
and \U$15732 ( \16715 , \16710 , \16714 );
and \U$15733 ( \16716 , \10226 , \2494 );
and \U$15734 ( \16717 , \10218 , \2492 );
nor \U$15735 ( \16718 , \16716 , \16717 );
xnor \U$15736 ( \16719 , \16718 , \2338 );
and \U$15737 ( \16720 , \16714 , \16719 );
and \U$15738 ( \16721 , \16710 , \16719 );
or \U$15739 ( \16722 , \16715 , \16720 , \16721 );
nand \U$15740 ( \16723 , \11635 , \1826 );
xnor \U$15741 ( \16724 , \16723 , \1750 );
and \U$15742 ( \16725 , \16722 , \16724 );
xor \U$15743 ( \16726 , \16497 , \16501 );
xor \U$15744 ( \16727 , \16726 , \16506 );
and \U$15745 ( \16728 , \16724 , \16727 );
and \U$15746 ( \16729 , \16722 , \16727 );
or \U$15747 ( \16730 , \16725 , \16728 , \16729 );
and \U$15748 ( \16731 , \16705 , \16730 );
and \U$15749 ( \16732 , \16653 , \16730 );
or \U$15750 ( \16733 , \16706 , \16731 , \16732 );
xor \U$15751 ( \16734 , \16380 , \16384 );
xor \U$15752 ( \16735 , \16734 , \16389 );
xor \U$15753 ( \16736 , \16481 , \16485 );
xor \U$15754 ( \16737 , \16736 , \16490 );
and \U$15755 ( \16738 , \16735 , \16737 );
xor \U$15756 ( \16739 , \16396 , \16400 );
xor \U$15757 ( \16740 , \16739 , \16405 );
and \U$15758 ( \16741 , \16737 , \16740 );
and \U$15759 ( \16742 , \16735 , \16740 );
or \U$15760 ( \16743 , \16738 , \16741 , \16742 );
xor \U$15761 ( \16744 , \16432 , \16436 );
xor \U$15762 ( \16745 , \16744 , \16441 );
xor \U$15763 ( \16746 , \16413 , \16417 );
xor \U$15764 ( \16747 , \16746 , \16422 );
and \U$15765 ( \16748 , \16745 , \16747 );
xor \U$15766 ( \16749 , \16461 , \16465 );
xor \U$15767 ( \16750 , \16749 , \16470 );
and \U$15768 ( \16751 , \16747 , \16750 );
and \U$15769 ( \16752 , \16745 , \16750 );
or \U$15770 ( \16753 , \16748 , \16751 , \16752 );
and \U$15771 ( \16754 , \16743 , \16753 );
xor \U$15772 ( \16755 , \16204 , \16208 );
xor \U$15773 ( \16756 , \16755 , \16213 );
and \U$15774 ( \16757 , \16753 , \16756 );
and \U$15775 ( \16758 , \16743 , \16756 );
or \U$15776 ( \16759 , \16754 , \16757 , \16758 );
and \U$15777 ( \16760 , \16733 , \16759 );
xor \U$15778 ( \16761 , \16520 , \16522 );
xor \U$15779 ( \16762 , \16761 , \16525 );
xor \U$15780 ( \16763 , \16530 , \16532 );
xor \U$15781 ( \16764 , \16763 , \16535 );
and \U$15782 ( \16765 , \16762 , \16764 );
xor \U$15783 ( \16766 , \16493 , \16509 );
xor \U$15784 ( \16767 , \16766 , \16512 );
and \U$15785 ( \16768 , \16764 , \16767 );
and \U$15786 ( \16769 , \16762 , \16767 );
or \U$15787 ( \16770 , \16765 , \16768 , \16769 );
and \U$15788 ( \16771 , \16759 , \16770 );
and \U$15789 ( \16772 , \16733 , \16770 );
or \U$15790 ( \16773 , \16760 , \16771 , \16772 );
xor \U$15791 ( \16774 , \16216 , \16232 );
xor \U$15792 ( \16775 , \16774 , \16249 );
xor \U$15793 ( \16776 , \16269 , \16285 );
xor \U$15794 ( \16777 , \16776 , \16302 );
and \U$15795 ( \16778 , \16775 , \16777 );
xor \U$15796 ( \16779 , \16547 , \16549 );
xor \U$15797 ( \16780 , \16779 , \16552 );
and \U$15798 ( \16781 , \16777 , \16780 );
and \U$15799 ( \16782 , \16775 , \16780 );
or \U$15800 ( \16783 , \16778 , \16781 , \16782 );
and \U$15801 ( \16784 , \16773 , \16783 );
xor \U$15802 ( \16785 , \16428 , \16476 );
xor \U$15803 ( \16786 , \16785 , \16515 );
xor \U$15804 ( \16787 , \16528 , \16538 );
xor \U$15805 ( \16788 , \16787 , \16541 );
and \U$15806 ( \16789 , \16786 , \16788 );
and \U$15807 ( \16790 , \16783 , \16789 );
and \U$15808 ( \16791 , \16773 , \16789 );
or \U$15809 ( \16792 , \16784 , \16790 , \16791 );
xor \U$15810 ( \16793 , \16200 , \16252 );
xor \U$15811 ( \16794 , \16793 , \16305 );
xor \U$15812 ( \16795 , \16518 , \16544 );
xor \U$15813 ( \16796 , \16795 , \16555 );
and \U$15814 ( \16797 , \16794 , \16796 );
xor \U$15815 ( \16798 , \16560 , \16562 );
xor \U$15816 ( \16799 , \16798 , \16565 );
and \U$15817 ( \16800 , \16796 , \16799 );
and \U$15818 ( \16801 , \16794 , \16799 );
or \U$15819 ( \16802 , \16797 , \16800 , \16801 );
and \U$15820 ( \16803 , \16792 , \16802 );
xor \U$15821 ( \16804 , \16576 , \16578 );
xor \U$15822 ( \16805 , \16804 , \16581 );
and \U$15823 ( \16806 , \16802 , \16805 );
and \U$15824 ( \16807 , \16792 , \16805 );
or \U$15825 ( \16808 , \16803 , \16806 , \16807 );
xor \U$15826 ( \16809 , \16321 , \16339 );
xor \U$15827 ( \16810 , \16809 , \16342 );
and \U$15828 ( \16811 , \16808 , \16810 );
xor \U$15829 ( \16812 , \16574 , \16584 );
xor \U$15830 ( \16813 , \16812 , \16587 );
and \U$15831 ( \16814 , \16810 , \16813 );
and \U$15832 ( \16815 , \16808 , \16813 );
or \U$15833 ( \16816 , \16811 , \16814 , \16815 );
and \U$15834 ( \16817 , \16601 , \16816 );
xor \U$15835 ( \16818 , \16601 , \16816 );
xor \U$15836 ( \16819 , \16808 , \16810 );
xor \U$15837 ( \16820 , \16819 , \16813 );
and \U$15838 ( \16821 , \2168 , \11482 );
and \U$15839 ( \16822 , \2052 , \11479 );
nor \U$15840 ( \16823 , \16821 , \16822 );
xnor \U$15841 ( \16824 , \16823 , \10427 );
and \U$15842 ( \16825 , \2459 , \10669 );
and \U$15843 ( \16826 , \2283 , \10667 );
nor \U$15844 ( \16827 , \16825 , \16826 );
xnor \U$15845 ( \16828 , \16827 , \10430 );
and \U$15846 ( \16829 , \16824 , \16828 );
and \U$15847 ( \16830 , \16828 , \1892 );
and \U$15848 ( \16831 , \16824 , \1892 );
or \U$15849 ( \16832 , \16829 , \16830 , \16831 );
and \U$15850 ( \16833 , \3508 , \8435 );
and \U$15851 ( \16834 , \3334 , \8433 );
nor \U$15852 ( \16835 , \16833 , \16834 );
xnor \U$15853 ( \16836 , \16835 , \8186 );
and \U$15854 ( \16837 , \3813 , \7906 );
and \U$15855 ( \16838 , \3675 , \7904 );
nor \U$15856 ( \16839 , \16837 , \16838 );
xnor \U$15857 ( \16840 , \16839 , \7646 );
and \U$15858 ( \16841 , \16836 , \16840 );
and \U$15859 ( \16842 , \4349 , \7412 );
and \U$15860 ( \16843 , \3932 , \7410 );
nor \U$15861 ( \16844 , \16842 , \16843 );
xnor \U$15862 ( \16845 , \16844 , \7097 );
and \U$15863 ( \16846 , \16840 , \16845 );
and \U$15864 ( \16847 , \16836 , \16845 );
or \U$15865 ( \16848 , \16841 , \16846 , \16847 );
and \U$15866 ( \16849 , \16832 , \16848 );
and \U$15867 ( \16850 , \2710 , \10101 );
and \U$15868 ( \16851 , \2467 , \10099 );
nor \U$15869 ( \16852 , \16850 , \16851 );
xnor \U$15870 ( \16853 , \16852 , \9791 );
and \U$15871 ( \16854 , \2901 , \9564 );
and \U$15872 ( \16855 , \2715 , \9562 );
nor \U$15873 ( \16856 , \16854 , \16855 );
xnor \U$15874 ( \16857 , \16856 , \9193 );
and \U$15875 ( \16858 , \16853 , \16857 );
and \U$15876 ( \16859 , \3309 , \9002 );
and \U$15877 ( \16860 , \3045 , \9000 );
nor \U$15878 ( \16861 , \16859 , \16860 );
xnor \U$15879 ( \16862 , \16861 , \8684 );
and \U$15880 ( \16863 , \16857 , \16862 );
and \U$15881 ( \16864 , \16853 , \16862 );
or \U$15882 ( \16865 , \16858 , \16863 , \16864 );
and \U$15883 ( \16866 , \16848 , \16865 );
and \U$15884 ( \16867 , \16832 , \16865 );
or \U$15885 ( \16868 , \16849 , \16866 , \16867 );
and \U$15886 ( \16869 , \4679 , \6903 );
and \U$15887 ( \16870 , \4557 , \6901 );
nor \U$15888 ( \16871 , \16869 , \16870 );
xnor \U$15889 ( \16872 , \16871 , \6563 );
and \U$15890 ( \16873 , \4940 , \6314 );
and \U$15891 ( \16874 , \4684 , \6312 );
nor \U$15892 ( \16875 , \16873 , \16874 );
xnor \U$15893 ( \16876 , \16875 , \6073 );
and \U$15894 ( \16877 , \16872 , \16876 );
and \U$15895 ( \16878 , \5439 , \5848 );
and \U$15896 ( \16879 , \5137 , \5846 );
nor \U$15897 ( \16880 , \16878 , \16879 );
xnor \U$15898 ( \16881 , \16880 , \5660 );
and \U$15899 ( \16882 , \16876 , \16881 );
and \U$15900 ( \16883 , \16872 , \16881 );
or \U$15901 ( \16884 , \16877 , \16882 , \16883 );
and \U$15902 ( \16885 , \5916 , \5474 );
and \U$15903 ( \16886 , \5447 , \5472 );
nor \U$15904 ( \16887 , \16885 , \16886 );
xnor \U$15905 ( \16888 , \16887 , \5242 );
and \U$15906 ( \16889 , \6185 , \5023 );
and \U$15907 ( \16890 , \5921 , \5021 );
nor \U$15908 ( \16891 , \16889 , \16890 );
xnor \U$15909 ( \16892 , \16891 , \4880 );
and \U$15910 ( \16893 , \16888 , \16892 );
and \U$15911 ( \16894 , \6816 , \4700 );
and \U$15912 ( \16895 , \6444 , \4698 );
nor \U$15913 ( \16896 , \16894 , \16895 );
xnor \U$15914 ( \16897 , \16896 , \4454 );
and \U$15915 ( \16898 , \16892 , \16897 );
and \U$15916 ( \16899 , \16888 , \16897 );
or \U$15917 ( \16900 , \16893 , \16898 , \16899 );
and \U$15918 ( \16901 , \16884 , \16900 );
and \U$15919 ( \16902 , \7168 , \4305 );
and \U$15920 ( \16903 , \6825 , \4303 );
nor \U$15921 ( \16904 , \16902 , \16903 );
xnor \U$15922 ( \16905 , \16904 , \4118 );
and \U$15923 ( \16906 , \7673 , \3992 );
and \U$15924 ( \16907 , \7370 , \3990 );
nor \U$15925 ( \16908 , \16906 , \16907 );
xnor \U$15926 ( \16909 , \16908 , \3787 );
and \U$15927 ( \16910 , \16905 , \16909 );
and \U$15928 ( \16911 , \8371 , \3586 );
and \U$15929 ( \16912 , \7845 , \3584 );
nor \U$15930 ( \16913 , \16911 , \16912 );
xnor \U$15931 ( \16914 , \16913 , \3437 );
and \U$15932 ( \16915 , \16909 , \16914 );
and \U$15933 ( \16916 , \16905 , \16914 );
or \U$15934 ( \16917 , \16910 , \16915 , \16916 );
and \U$15935 ( \16918 , \16900 , \16917 );
and \U$15936 ( \16919 , \16884 , \16917 );
or \U$15937 ( \16920 , \16901 , \16918 , \16919 );
and \U$15938 ( \16921 , \16868 , \16920 );
and \U$15939 ( \16922 , \10829 , \2494 );
and \U$15940 ( \16923 , \10226 , \2492 );
nor \U$15941 ( \16924 , \16922 , \16923 );
xnor \U$15942 ( \16925 , \16924 , \2338 );
and \U$15943 ( \16926 , \11015 , \2222 );
and \U$15944 ( \16927 , \10834 , \2220 );
nor \U$15945 ( \16928 , \16926 , \16927 );
xnor \U$15946 ( \16929 , \16928 , \2109 );
and \U$15947 ( \16930 , \16925 , \16929 );
nand \U$15948 ( \16931 , \11635 , \2026 );
xnor \U$15949 ( \16932 , \16931 , \1892 );
and \U$15950 ( \16933 , \16929 , \16932 );
and \U$15951 ( \16934 , \16925 , \16932 );
or \U$15952 ( \16935 , \16930 , \16933 , \16934 );
and \U$15953 ( \16936 , \9041 , \3264 );
and \U$15954 ( \16937 , \8795 , \3262 );
nor \U$15955 ( \16938 , \16936 , \16937 );
xnor \U$15956 ( \16939 , \16938 , \3122 );
and \U$15957 ( \16940 , \9365 , \2968 );
and \U$15958 ( \16941 , \9046 , \2966 );
nor \U$15959 ( \16942 , \16940 , \16941 );
xnor \U$15960 ( \16943 , \16942 , \2831 );
and \U$15961 ( \16944 , \16939 , \16943 );
and \U$15962 ( \16945 , \10218 , \2762 );
and \U$15963 ( \16946 , \9649 , \2760 );
nor \U$15964 ( \16947 , \16945 , \16946 );
xnor \U$15965 ( \16948 , \16947 , \2610 );
and \U$15966 ( \16949 , \16943 , \16948 );
and \U$15967 ( \16950 , \16939 , \16948 );
or \U$15968 ( \16951 , \16944 , \16949 , \16950 );
and \U$15969 ( \16952 , \16935 , \16951 );
and \U$15970 ( \16953 , \10834 , \2222 );
and \U$15971 ( \16954 , \10829 , \2220 );
nor \U$15972 ( \16955 , \16953 , \16954 );
xnor \U$15973 ( \16956 , \16955 , \2109 );
and \U$15974 ( \16957 , \16951 , \16956 );
and \U$15975 ( \16958 , \16935 , \16956 );
or \U$15976 ( \16959 , \16952 , \16957 , \16958 );
and \U$15977 ( \16960 , \16920 , \16959 );
and \U$15978 ( \16961 , \16868 , \16959 );
or \U$15979 ( \16962 , \16921 , \16960 , \16961 );
and \U$15980 ( \16963 , \11635 , \2028 );
and \U$15981 ( \16964 , \11015 , \2026 );
nor \U$15982 ( \16965 , \16963 , \16964 );
xnor \U$15983 ( \16966 , \16965 , \1892 );
xor \U$15984 ( \16967 , \16638 , \16642 );
xor \U$15985 ( \16968 , \16967 , \16647 );
and \U$15986 ( \16969 , \16966 , \16968 );
xor \U$15987 ( \16970 , \16710 , \16714 );
xor \U$15988 ( \16971 , \16970 , \16719 );
and \U$15989 ( \16972 , \16968 , \16971 );
and \U$15990 ( \16973 , \16966 , \16971 );
or \U$15991 ( \16974 , \16969 , \16972 , \16973 );
xor \U$15992 ( \16975 , \16605 , \16609 );
xor \U$15993 ( \16976 , \16975 , \16614 );
xor \U$15994 ( \16977 , \16621 , \16625 );
xor \U$15995 ( \16978 , \16977 , \16630 );
and \U$15996 ( \16979 , \16976 , \16978 );
xor \U$15997 ( \16980 , \16673 , \16677 );
xor \U$15998 ( \16981 , \16980 , \16682 );
and \U$15999 ( \16982 , \16978 , \16981 );
and \U$16000 ( \16983 , \16976 , \16981 );
or \U$16001 ( \16984 , \16979 , \16982 , \16983 );
and \U$16002 ( \16985 , \16974 , \16984 );
xor \U$16003 ( \16986 , \16448 , \16452 );
xor \U$16004 ( \16987 , \16986 , \1750 );
and \U$16005 ( \16988 , \16984 , \16987 );
and \U$16006 ( \16989 , \16974 , \16987 );
or \U$16007 ( \16990 , \16985 , \16988 , \16989 );
and \U$16008 ( \16991 , \16962 , \16990 );
xor \U$16009 ( \16992 , \16722 , \16724 );
xor \U$16010 ( \16993 , \16992 , \16727 );
xor \U$16011 ( \16994 , \16735 , \16737 );
xor \U$16012 ( \16995 , \16994 , \16740 );
and \U$16013 ( \16996 , \16993 , \16995 );
xor \U$16014 ( \16997 , \16745 , \16747 );
xor \U$16015 ( \16998 , \16997 , \16750 );
and \U$16016 ( \16999 , \16995 , \16998 );
and \U$16017 ( \17000 , \16993 , \16998 );
or \U$16018 ( \17001 , \16996 , \16999 , \17000 );
and \U$16019 ( \17002 , \16990 , \17001 );
and \U$16020 ( \17003 , \16962 , \17001 );
or \U$16021 ( \17004 , \16991 , \17002 , \17003 );
xor \U$16022 ( \17005 , \16392 , \16408 );
xor \U$16023 ( \17006 , \17005 , \16425 );
xor \U$16024 ( \17007 , \16444 , \16456 );
xor \U$16025 ( \17008 , \17007 , \16473 );
and \U$16026 ( \17009 , \17006 , \17008 );
xor \U$16027 ( \17010 , \16762 , \16764 );
xor \U$16028 ( \17011 , \17010 , \16767 );
and \U$16029 ( \17012 , \17008 , \17011 );
and \U$16030 ( \17013 , \17006 , \17011 );
or \U$16031 ( \17014 , \17009 , \17012 , \17013 );
and \U$16032 ( \17015 , \17004 , \17014 );
xor \U$16033 ( \17016 , \16653 , \16705 );
xor \U$16034 ( \17017 , \17016 , \16730 );
xor \U$16035 ( \17018 , \16743 , \16753 );
xor \U$16036 ( \17019 , \17018 , \16756 );
and \U$16037 ( \17020 , \17017 , \17019 );
and \U$16038 ( \17021 , \17014 , \17020 );
and \U$16039 ( \17022 , \17004 , \17020 );
or \U$16040 ( \17023 , \17015 , \17021 , \17022 );
xor \U$16041 ( \17024 , \16733 , \16759 );
xor \U$16042 ( \17025 , \17024 , \16770 );
xor \U$16043 ( \17026 , \16775 , \16777 );
xor \U$16044 ( \17027 , \17026 , \16780 );
and \U$16045 ( \17028 , \17025 , \17027 );
xor \U$16046 ( \17029 , \16786 , \16788 );
and \U$16047 ( \17030 , \17027 , \17029 );
and \U$16048 ( \17031 , \17025 , \17029 );
or \U$16049 ( \17032 , \17028 , \17030 , \17031 );
and \U$16050 ( \17033 , \17023 , \17032 );
xor \U$16051 ( \17034 , \16794 , \16796 );
xor \U$16052 ( \17035 , \17034 , \16799 );
and \U$16053 ( \17036 , \17032 , \17035 );
and \U$16054 ( \17037 , \17023 , \17035 );
or \U$16055 ( \17038 , \17033 , \17036 , \17037 );
xor \U$16056 ( \17039 , \16558 , \16568 );
xor \U$16057 ( \17040 , \17039 , \16571 );
and \U$16058 ( \17041 , \17038 , \17040 );
xor \U$16059 ( \17042 , \16792 , \16802 );
xor \U$16060 ( \17043 , \17042 , \16805 );
and \U$16061 ( \17044 , \17040 , \17043 );
and \U$16062 ( \17045 , \17038 , \17043 );
or \U$16063 ( \17046 , \17041 , \17044 , \17045 );
and \U$16064 ( \17047 , \16820 , \17046 );
xor \U$16065 ( \17048 , \16820 , \17046 );
xor \U$16066 ( \17049 , \17038 , \17040 );
xor \U$16067 ( \17050 , \17049 , \17043 );
and \U$16068 ( \17051 , \2283 , \11482 );
and \U$16069 ( \17052 , \2168 , \11479 );
nor \U$16070 ( \17053 , \17051 , \17052 );
xnor \U$16071 ( \17054 , \17053 , \10427 );
and \U$16072 ( \17055 , \2467 , \10669 );
and \U$16073 ( \17056 , \2459 , \10667 );
nor \U$16074 ( \17057 , \17055 , \17056 );
xnor \U$16075 ( \17058 , \17057 , \10430 );
and \U$16076 ( \17059 , \17054 , \17058 );
and \U$16077 ( \17060 , \2715 , \10101 );
and \U$16078 ( \17061 , \2710 , \10099 );
nor \U$16079 ( \17062 , \17060 , \17061 );
xnor \U$16080 ( \17063 , \17062 , \9791 );
and \U$16081 ( \17064 , \17058 , \17063 );
and \U$16082 ( \17065 , \17054 , \17063 );
or \U$16083 ( \17066 , \17059 , \17064 , \17065 );
and \U$16084 ( \17067 , \3045 , \9564 );
and \U$16085 ( \17068 , \2901 , \9562 );
nor \U$16086 ( \17069 , \17067 , \17068 );
xnor \U$16087 ( \17070 , \17069 , \9193 );
and \U$16088 ( \17071 , \3334 , \9002 );
and \U$16089 ( \17072 , \3309 , \9000 );
nor \U$16090 ( \17073 , \17071 , \17072 );
xnor \U$16091 ( \17074 , \17073 , \8684 );
and \U$16092 ( \17075 , \17070 , \17074 );
and \U$16093 ( \17076 , \3675 , \8435 );
and \U$16094 ( \17077 , \3508 , \8433 );
nor \U$16095 ( \17078 , \17076 , \17077 );
xnor \U$16096 ( \17079 , \17078 , \8186 );
and \U$16097 ( \17080 , \17074 , \17079 );
and \U$16098 ( \17081 , \17070 , \17079 );
or \U$16099 ( \17082 , \17075 , \17080 , \17081 );
and \U$16100 ( \17083 , \17066 , \17082 );
and \U$16101 ( \17084 , \3932 , \7906 );
and \U$16102 ( \17085 , \3813 , \7904 );
nor \U$16103 ( \17086 , \17084 , \17085 );
xnor \U$16104 ( \17087 , \17086 , \7646 );
and \U$16105 ( \17088 , \4557 , \7412 );
and \U$16106 ( \17089 , \4349 , \7410 );
nor \U$16107 ( \17090 , \17088 , \17089 );
xnor \U$16108 ( \17091 , \17090 , \7097 );
and \U$16109 ( \17092 , \17087 , \17091 );
and \U$16110 ( \17093 , \4684 , \6903 );
and \U$16111 ( \17094 , \4679 , \6901 );
nor \U$16112 ( \17095 , \17093 , \17094 );
xnor \U$16113 ( \17096 , \17095 , \6563 );
and \U$16114 ( \17097 , \17091 , \17096 );
and \U$16115 ( \17098 , \17087 , \17096 );
or \U$16116 ( \17099 , \17092 , \17097 , \17098 );
and \U$16117 ( \17100 , \17082 , \17099 );
and \U$16118 ( \17101 , \17066 , \17099 );
or \U$16119 ( \17102 , \17083 , \17100 , \17101 );
and \U$16120 ( \17103 , \6444 , \5023 );
and \U$16121 ( \17104 , \6185 , \5021 );
nor \U$16122 ( \17105 , \17103 , \17104 );
xnor \U$16123 ( \17106 , \17105 , \4880 );
and \U$16124 ( \17107 , \6825 , \4700 );
and \U$16125 ( \17108 , \6816 , \4698 );
nor \U$16126 ( \17109 , \17107 , \17108 );
xnor \U$16127 ( \17110 , \17109 , \4454 );
and \U$16128 ( \17111 , \17106 , \17110 );
and \U$16129 ( \17112 , \7370 , \4305 );
and \U$16130 ( \17113 , \7168 , \4303 );
nor \U$16131 ( \17114 , \17112 , \17113 );
xnor \U$16132 ( \17115 , \17114 , \4118 );
and \U$16133 ( \17116 , \17110 , \17115 );
and \U$16134 ( \17117 , \17106 , \17115 );
or \U$16135 ( \17118 , \17111 , \17116 , \17117 );
and \U$16136 ( \17119 , \7845 , \3992 );
and \U$16137 ( \17120 , \7673 , \3990 );
nor \U$16138 ( \17121 , \17119 , \17120 );
xnor \U$16139 ( \17122 , \17121 , \3787 );
and \U$16140 ( \17123 , \8795 , \3586 );
and \U$16141 ( \17124 , \8371 , \3584 );
nor \U$16142 ( \17125 , \17123 , \17124 );
xnor \U$16143 ( \17126 , \17125 , \3437 );
and \U$16144 ( \17127 , \17122 , \17126 );
and \U$16145 ( \17128 , \9046 , \3264 );
and \U$16146 ( \17129 , \9041 , \3262 );
nor \U$16147 ( \17130 , \17128 , \17129 );
xnor \U$16148 ( \17131 , \17130 , \3122 );
and \U$16149 ( \17132 , \17126 , \17131 );
and \U$16150 ( \17133 , \17122 , \17131 );
or \U$16151 ( \17134 , \17127 , \17132 , \17133 );
and \U$16152 ( \17135 , \17118 , \17134 );
and \U$16153 ( \17136 , \5137 , \6314 );
and \U$16154 ( \17137 , \4940 , \6312 );
nor \U$16155 ( \17138 , \17136 , \17137 );
xnor \U$16156 ( \17139 , \17138 , \6073 );
and \U$16157 ( \17140 , \5447 , \5848 );
and \U$16158 ( \17141 , \5439 , \5846 );
nor \U$16159 ( \17142 , \17140 , \17141 );
xnor \U$16160 ( \17143 , \17142 , \5660 );
and \U$16161 ( \17144 , \17139 , \17143 );
and \U$16162 ( \17145 , \5921 , \5474 );
and \U$16163 ( \17146 , \5916 , \5472 );
nor \U$16164 ( \17147 , \17145 , \17146 );
xnor \U$16165 ( \17148 , \17147 , \5242 );
and \U$16166 ( \17149 , \17143 , \17148 );
and \U$16167 ( \17150 , \17139 , \17148 );
or \U$16168 ( \17151 , \17144 , \17149 , \17150 );
and \U$16169 ( \17152 , \17134 , \17151 );
and \U$16170 ( \17153 , \17118 , \17151 );
or \U$16171 ( \17154 , \17135 , \17152 , \17153 );
and \U$16172 ( \17155 , \17102 , \17154 );
and \U$16173 ( \17156 , \9649 , \2968 );
and \U$16174 ( \17157 , \9365 , \2966 );
nor \U$16175 ( \17158 , \17156 , \17157 );
xnor \U$16176 ( \17159 , \17158 , \2831 );
and \U$16177 ( \17160 , \10226 , \2762 );
and \U$16178 ( \17161 , \10218 , \2760 );
nor \U$16179 ( \17162 , \17160 , \17161 );
xnor \U$16180 ( \17163 , \17162 , \2610 );
and \U$16181 ( \17164 , \17159 , \17163 );
and \U$16182 ( \17165 , \10834 , \2494 );
and \U$16183 ( \17166 , \10829 , \2492 );
nor \U$16184 ( \17167 , \17165 , \17166 );
xnor \U$16185 ( \17168 , \17167 , \2338 );
and \U$16186 ( \17169 , \17163 , \17168 );
and \U$16187 ( \17170 , \17159 , \17168 );
or \U$16188 ( \17171 , \17164 , \17169 , \17170 );
xor \U$16189 ( \17172 , \16925 , \16929 );
xor \U$16190 ( \17173 , \17172 , \16932 );
and \U$16191 ( \17174 , \17171 , \17173 );
xor \U$16192 ( \17175 , \16939 , \16943 );
xor \U$16193 ( \17176 , \17175 , \16948 );
and \U$16194 ( \17177 , \17173 , \17176 );
and \U$16195 ( \17178 , \17171 , \17176 );
or \U$16196 ( \17179 , \17174 , \17177 , \17178 );
and \U$16197 ( \17180 , \17154 , \17179 );
and \U$16198 ( \17181 , \17102 , \17179 );
or \U$16199 ( \17182 , \17155 , \17180 , \17181 );
xor \U$16200 ( \17183 , \16872 , \16876 );
xor \U$16201 ( \17184 , \17183 , \16881 );
xor \U$16202 ( \17185 , \16888 , \16892 );
xor \U$16203 ( \17186 , \17185 , \16897 );
and \U$16204 ( \17187 , \17184 , \17186 );
xor \U$16205 ( \17188 , \16905 , \16909 );
xor \U$16206 ( \17189 , \17188 , \16914 );
and \U$16207 ( \17190 , \17186 , \17189 );
and \U$16208 ( \17191 , \17184 , \17189 );
or \U$16209 ( \17192 , \17187 , \17190 , \17191 );
xor \U$16210 ( \17193 , \16824 , \16828 );
xor \U$16211 ( \17194 , \17193 , \1892 );
xor \U$16212 ( \17195 , \16836 , \16840 );
xor \U$16213 ( \17196 , \17195 , \16845 );
and \U$16214 ( \17197 , \17194 , \17196 );
xor \U$16215 ( \17198 , \16853 , \16857 );
xor \U$16216 ( \17199 , \17198 , \16862 );
and \U$16217 ( \17200 , \17196 , \17199 );
and \U$16218 ( \17201 , \17194 , \17199 );
or \U$16219 ( \17202 , \17197 , \17200 , \17201 );
and \U$16220 ( \17203 , \17192 , \17202 );
xor \U$16221 ( \17204 , \16657 , \16661 );
xor \U$16222 ( \17205 , \17204 , \16666 );
and \U$16223 ( \17206 , \17202 , \17205 );
and \U$16224 ( \17207 , \17192 , \17205 );
or \U$16225 ( \17208 , \17203 , \17206 , \17207 );
and \U$16226 ( \17209 , \17182 , \17208 );
xor \U$16227 ( \17210 , \16690 , \16694 );
xor \U$16228 ( \17211 , \17210 , \16699 );
xor \U$16229 ( \17212 , \16966 , \16968 );
xor \U$16230 ( \17213 , \17212 , \16971 );
and \U$16231 ( \17214 , \17211 , \17213 );
xor \U$16232 ( \17215 , \16976 , \16978 );
xor \U$16233 ( \17216 , \17215 , \16981 );
and \U$16234 ( \17217 , \17213 , \17216 );
and \U$16235 ( \17218 , \17211 , \17216 );
or \U$16236 ( \17219 , \17214 , \17217 , \17218 );
and \U$16237 ( \17220 , \17208 , \17219 );
and \U$16238 ( \17221 , \17182 , \17219 );
or \U$16239 ( \17222 , \17209 , \17220 , \17221 );
xor \U$16240 ( \17223 , \16832 , \16848 );
xor \U$16241 ( \17224 , \17223 , \16865 );
xor \U$16242 ( \17225 , \16884 , \16900 );
xor \U$16243 ( \17226 , \17225 , \16917 );
and \U$16244 ( \17227 , \17224 , \17226 );
xor \U$16245 ( \17228 , \16935 , \16951 );
xor \U$16246 ( \17229 , \17228 , \16956 );
and \U$16247 ( \17230 , \17226 , \17229 );
and \U$16248 ( \17231 , \17224 , \17229 );
or \U$16249 ( \17232 , \17227 , \17230 , \17231 );
xor \U$16250 ( \17233 , \16617 , \16633 );
xor \U$16251 ( \17234 , \17233 , \16650 );
and \U$16252 ( \17235 , \17232 , \17234 );
xor \U$16253 ( \17236 , \16669 , \16685 );
xor \U$16254 ( \17237 , \17236 , \16702 );
and \U$16255 ( \17238 , \17234 , \17237 );
and \U$16256 ( \17239 , \17232 , \17237 );
or \U$16257 ( \17240 , \17235 , \17238 , \17239 );
and \U$16258 ( \17241 , \17222 , \17240 );
xor \U$16259 ( \17242 , \16868 , \16920 );
xor \U$16260 ( \17243 , \17242 , \16959 );
xor \U$16261 ( \17244 , \16974 , \16984 );
xor \U$16262 ( \17245 , \17244 , \16987 );
and \U$16263 ( \17246 , \17243 , \17245 );
xor \U$16264 ( \17247 , \16993 , \16995 );
xor \U$16265 ( \17248 , \17247 , \16998 );
and \U$16266 ( \17249 , \17245 , \17248 );
and \U$16267 ( \17250 , \17243 , \17248 );
or \U$16268 ( \17251 , \17246 , \17249 , \17250 );
and \U$16269 ( \17252 , \17240 , \17251 );
and \U$16270 ( \17253 , \17222 , \17251 );
or \U$16271 ( \17254 , \17241 , \17252 , \17253 );
xor \U$16272 ( \17255 , \16962 , \16990 );
xor \U$16273 ( \17256 , \17255 , \17001 );
xor \U$16274 ( \17257 , \17006 , \17008 );
xor \U$16275 ( \17258 , \17257 , \17011 );
and \U$16276 ( \17259 , \17256 , \17258 );
xor \U$16277 ( \17260 , \17017 , \17019 );
and \U$16278 ( \17261 , \17258 , \17260 );
and \U$16279 ( \17262 , \17256 , \17260 );
or \U$16280 ( \17263 , \17259 , \17261 , \17262 );
and \U$16281 ( \17264 , \17254 , \17263 );
xor \U$16282 ( \17265 , \17025 , \17027 );
xor \U$16283 ( \17266 , \17265 , \17029 );
and \U$16284 ( \17267 , \17263 , \17266 );
and \U$16285 ( \17268 , \17254 , \17266 );
or \U$16286 ( \17269 , \17264 , \17267 , \17268 );
xor \U$16287 ( \17270 , \16773 , \16783 );
xor \U$16288 ( \17271 , \17270 , \16789 );
and \U$16289 ( \17272 , \17269 , \17271 );
xor \U$16290 ( \17273 , \17023 , \17032 );
xor \U$16291 ( \17274 , \17273 , \17035 );
and \U$16292 ( \17275 , \17271 , \17274 );
and \U$16293 ( \17276 , \17269 , \17274 );
or \U$16294 ( \17277 , \17272 , \17275 , \17276 );
and \U$16295 ( \17278 , \17050 , \17277 );
xor \U$16296 ( \17279 , \17050 , \17277 );
xor \U$16297 ( \17280 , \17269 , \17271 );
xor \U$16298 ( \17281 , \17280 , \17274 );
and \U$16299 ( \17282 , \7673 , \4305 );
and \U$16300 ( \17283 , \7370 , \4303 );
nor \U$16301 ( \17284 , \17282 , \17283 );
xnor \U$16302 ( \17285 , \17284 , \4118 );
and \U$16303 ( \17286 , \8371 , \3992 );
and \U$16304 ( \17287 , \7845 , \3990 );
nor \U$16305 ( \17288 , \17286 , \17287 );
xnor \U$16306 ( \17289 , \17288 , \3787 );
and \U$16307 ( \17290 , \17285 , \17289 );
and \U$16308 ( \17291 , \9041 , \3586 );
and \U$16309 ( \17292 , \8795 , \3584 );
nor \U$16310 ( \17293 , \17291 , \17292 );
xnor \U$16311 ( \17294 , \17293 , \3437 );
and \U$16312 ( \17295 , \17289 , \17294 );
and \U$16313 ( \17296 , \17285 , \17294 );
or \U$16314 ( \17297 , \17290 , \17295 , \17296 );
and \U$16315 ( \17298 , \4940 , \6903 );
and \U$16316 ( \17299 , \4684 , \6901 );
nor \U$16317 ( \17300 , \17298 , \17299 );
xnor \U$16318 ( \17301 , \17300 , \6563 );
and \U$16319 ( \17302 , \5439 , \6314 );
and \U$16320 ( \17303 , \5137 , \6312 );
nor \U$16321 ( \17304 , \17302 , \17303 );
xnor \U$16322 ( \17305 , \17304 , \6073 );
and \U$16323 ( \17306 , \17301 , \17305 );
and \U$16324 ( \17307 , \5916 , \5848 );
and \U$16325 ( \17308 , \5447 , \5846 );
nor \U$16326 ( \17309 , \17307 , \17308 );
xnor \U$16327 ( \17310 , \17309 , \5660 );
and \U$16328 ( \17311 , \17305 , \17310 );
and \U$16329 ( \17312 , \17301 , \17310 );
or \U$16330 ( \17313 , \17306 , \17311 , \17312 );
and \U$16331 ( \17314 , \17297 , \17313 );
and \U$16332 ( \17315 , \6185 , \5474 );
and \U$16333 ( \17316 , \5921 , \5472 );
nor \U$16334 ( \17317 , \17315 , \17316 );
xnor \U$16335 ( \17318 , \17317 , \5242 );
and \U$16336 ( \17319 , \6816 , \5023 );
and \U$16337 ( \17320 , \6444 , \5021 );
nor \U$16338 ( \17321 , \17319 , \17320 );
xnor \U$16339 ( \17322 , \17321 , \4880 );
and \U$16340 ( \17323 , \17318 , \17322 );
and \U$16341 ( \17324 , \7168 , \4700 );
and \U$16342 ( \17325 , \6825 , \4698 );
nor \U$16343 ( \17326 , \17324 , \17325 );
xnor \U$16344 ( \17327 , \17326 , \4454 );
and \U$16345 ( \17328 , \17322 , \17327 );
and \U$16346 ( \17329 , \17318 , \17327 );
or \U$16347 ( \17330 , \17323 , \17328 , \17329 );
and \U$16348 ( \17331 , \17313 , \17330 );
and \U$16349 ( \17332 , \17297 , \17330 );
or \U$16350 ( \17333 , \17314 , \17331 , \17332 );
and \U$16351 ( \17334 , \2459 , \11482 );
and \U$16352 ( \17335 , \2283 , \11479 );
nor \U$16353 ( \17336 , \17334 , \17335 );
xnor \U$16354 ( \17337 , \17336 , \10427 );
and \U$16355 ( \17338 , \2710 , \10669 );
and \U$16356 ( \17339 , \2467 , \10667 );
nor \U$16357 ( \17340 , \17338 , \17339 );
xnor \U$16358 ( \17341 , \17340 , \10430 );
and \U$16359 ( \17342 , \17337 , \17341 );
and \U$16360 ( \17343 , \17341 , \2109 );
and \U$16361 ( \17344 , \17337 , \2109 );
or \U$16362 ( \17345 , \17342 , \17343 , \17344 );
and \U$16363 ( \17346 , \3813 , \8435 );
and \U$16364 ( \17347 , \3675 , \8433 );
nor \U$16365 ( \17348 , \17346 , \17347 );
xnor \U$16366 ( \17349 , \17348 , \8186 );
and \U$16367 ( \17350 , \4349 , \7906 );
and \U$16368 ( \17351 , \3932 , \7904 );
nor \U$16369 ( \17352 , \17350 , \17351 );
xnor \U$16370 ( \17353 , \17352 , \7646 );
and \U$16371 ( \17354 , \17349 , \17353 );
and \U$16372 ( \17355 , \4679 , \7412 );
and \U$16373 ( \17356 , \4557 , \7410 );
nor \U$16374 ( \17357 , \17355 , \17356 );
xnor \U$16375 ( \17358 , \17357 , \7097 );
and \U$16376 ( \17359 , \17353 , \17358 );
and \U$16377 ( \17360 , \17349 , \17358 );
or \U$16378 ( \17361 , \17354 , \17359 , \17360 );
and \U$16379 ( \17362 , \17345 , \17361 );
and \U$16380 ( \17363 , \2901 , \10101 );
and \U$16381 ( \17364 , \2715 , \10099 );
nor \U$16382 ( \17365 , \17363 , \17364 );
xnor \U$16383 ( \17366 , \17365 , \9791 );
and \U$16384 ( \17367 , \3309 , \9564 );
and \U$16385 ( \17368 , \3045 , \9562 );
nor \U$16386 ( \17369 , \17367 , \17368 );
xnor \U$16387 ( \17370 , \17369 , \9193 );
and \U$16388 ( \17371 , \17366 , \17370 );
and \U$16389 ( \17372 , \3508 , \9002 );
and \U$16390 ( \17373 , \3334 , \9000 );
nor \U$16391 ( \17374 , \17372 , \17373 );
xnor \U$16392 ( \17375 , \17374 , \8684 );
and \U$16393 ( \17376 , \17370 , \17375 );
and \U$16394 ( \17377 , \17366 , \17375 );
or \U$16395 ( \17378 , \17371 , \17376 , \17377 );
and \U$16396 ( \17379 , \17361 , \17378 );
and \U$16397 ( \17380 , \17345 , \17378 );
or \U$16398 ( \17381 , \17362 , \17379 , \17380 );
and \U$16399 ( \17382 , \17333 , \17381 );
and \U$16400 ( \17383 , \9365 , \3264 );
and \U$16401 ( \17384 , \9046 , \3262 );
nor \U$16402 ( \17385 , \17383 , \17384 );
xnor \U$16403 ( \17386 , \17385 , \3122 );
and \U$16404 ( \17387 , \10218 , \2968 );
and \U$16405 ( \17388 , \9649 , \2966 );
nor \U$16406 ( \17389 , \17387 , \17388 );
xnor \U$16407 ( \17390 , \17389 , \2831 );
and \U$16408 ( \17391 , \17386 , \17390 );
and \U$16409 ( \17392 , \10829 , \2762 );
and \U$16410 ( \17393 , \10226 , \2760 );
nor \U$16411 ( \17394 , \17392 , \17393 );
xnor \U$16412 ( \17395 , \17394 , \2610 );
and \U$16413 ( \17396 , \17390 , \17395 );
and \U$16414 ( \17397 , \17386 , \17395 );
or \U$16415 ( \17398 , \17391 , \17396 , \17397 );
and \U$16416 ( \17399 , \11015 , \2494 );
and \U$16417 ( \17400 , \10834 , \2492 );
nor \U$16418 ( \17401 , \17399 , \17400 );
xnor \U$16419 ( \17402 , \17401 , \2338 );
nand \U$16420 ( \17403 , \11635 , \2220 );
xnor \U$16421 ( \17404 , \17403 , \2109 );
and \U$16422 ( \17405 , \17402 , \17404 );
and \U$16423 ( \17406 , \17398 , \17405 );
and \U$16424 ( \17407 , \11635 , \2222 );
and \U$16425 ( \17408 , \11015 , \2220 );
nor \U$16426 ( \17409 , \17407 , \17408 );
xnor \U$16427 ( \17410 , \17409 , \2109 );
and \U$16428 ( \17411 , \17405 , \17410 );
and \U$16429 ( \17412 , \17398 , \17410 );
or \U$16430 ( \17413 , \17406 , \17411 , \17412 );
and \U$16431 ( \17414 , \17381 , \17413 );
and \U$16432 ( \17415 , \17333 , \17413 );
or \U$16433 ( \17416 , \17382 , \17414 , \17415 );
xor \U$16434 ( \17417 , \17070 , \17074 );
xor \U$16435 ( \17418 , \17417 , \17079 );
xor \U$16436 ( \17419 , \17139 , \17143 );
xor \U$16437 ( \17420 , \17419 , \17148 );
and \U$16438 ( \17421 , \17418 , \17420 );
xor \U$16439 ( \17422 , \17087 , \17091 );
xor \U$16440 ( \17423 , \17422 , \17096 );
and \U$16441 ( \17424 , \17420 , \17423 );
and \U$16442 ( \17425 , \17418 , \17423 );
or \U$16443 ( \17426 , \17421 , \17424 , \17425 );
xor \U$16444 ( \17427 , \17106 , \17110 );
xor \U$16445 ( \17428 , \17427 , \17115 );
xor \U$16446 ( \17429 , \17159 , \17163 );
xor \U$16447 ( \17430 , \17429 , \17168 );
and \U$16448 ( \17431 , \17428 , \17430 );
xor \U$16449 ( \17432 , \17122 , \17126 );
xor \U$16450 ( \17433 , \17432 , \17131 );
and \U$16451 ( \17434 , \17430 , \17433 );
and \U$16452 ( \17435 , \17428 , \17433 );
or \U$16453 ( \17436 , \17431 , \17434 , \17435 );
and \U$16454 ( \17437 , \17426 , \17436 );
xor \U$16455 ( \17438 , \17194 , \17196 );
xor \U$16456 ( \17439 , \17438 , \17199 );
and \U$16457 ( \17440 , \17436 , \17439 );
and \U$16458 ( \17441 , \17426 , \17439 );
or \U$16459 ( \17442 , \17437 , \17440 , \17441 );
and \U$16460 ( \17443 , \17416 , \17442 );
xor \U$16461 ( \17444 , \17118 , \17134 );
xor \U$16462 ( \17445 , \17444 , \17151 );
xor \U$16463 ( \17446 , \17184 , \17186 );
xor \U$16464 ( \17447 , \17446 , \17189 );
and \U$16465 ( \17448 , \17445 , \17447 );
xor \U$16466 ( \17449 , \17171 , \17173 );
xor \U$16467 ( \17450 , \17449 , \17176 );
and \U$16468 ( \17451 , \17447 , \17450 );
and \U$16469 ( \17452 , \17445 , \17450 );
or \U$16470 ( \17453 , \17448 , \17451 , \17452 );
and \U$16471 ( \17454 , \17442 , \17453 );
and \U$16472 ( \17455 , \17416 , \17453 );
or \U$16473 ( \17456 , \17443 , \17454 , \17455 );
xor \U$16474 ( \17457 , \17224 , \17226 );
xor \U$16475 ( \17458 , \17457 , \17229 );
xor \U$16476 ( \17459 , \17192 , \17202 );
xor \U$16477 ( \17460 , \17459 , \17205 );
and \U$16478 ( \17461 , \17458 , \17460 );
xor \U$16479 ( \17462 , \17211 , \17213 );
xor \U$16480 ( \17463 , \17462 , \17216 );
and \U$16481 ( \17464 , \17460 , \17463 );
and \U$16482 ( \17465 , \17458 , \17463 );
or \U$16483 ( \17466 , \17461 , \17464 , \17465 );
and \U$16484 ( \17467 , \17456 , \17466 );
xor \U$16485 ( \17468 , \17243 , \17245 );
xor \U$16486 ( \17469 , \17468 , \17248 );
and \U$16487 ( \17470 , \17466 , \17469 );
and \U$16488 ( \17471 , \17456 , \17469 );
or \U$16489 ( \17472 , \17467 , \17470 , \17471 );
xor \U$16490 ( \17473 , \17222 , \17240 );
xor \U$16491 ( \17474 , \17473 , \17251 );
and \U$16492 ( \17475 , \17472 , \17474 );
xor \U$16493 ( \17476 , \17256 , \17258 );
xor \U$16494 ( \17477 , \17476 , \17260 );
and \U$16495 ( \17478 , \17474 , \17477 );
and \U$16496 ( \17479 , \17472 , \17477 );
or \U$16497 ( \17480 , \17475 , \17478 , \17479 );
xor \U$16498 ( \17481 , \17004 , \17014 );
xor \U$16499 ( \17482 , \17481 , \17020 );
and \U$16500 ( \17483 , \17480 , \17482 );
xor \U$16501 ( \17484 , \17254 , \17263 );
xor \U$16502 ( \17485 , \17484 , \17266 );
and \U$16503 ( \17486 , \17482 , \17485 );
and \U$16504 ( \17487 , \17480 , \17485 );
or \U$16505 ( \17488 , \17483 , \17486 , \17487 );
and \U$16506 ( \17489 , \17281 , \17488 );
xor \U$16507 ( \17490 , \17281 , \17488 );
xor \U$16508 ( \17491 , \17480 , \17482 );
xor \U$16509 ( \17492 , \17491 , \17485 );
and \U$16510 ( \17493 , \6825 , \5023 );
and \U$16511 ( \17494 , \6816 , \5021 );
nor \U$16512 ( \17495 , \17493 , \17494 );
xnor \U$16513 ( \17496 , \17495 , \4880 );
and \U$16514 ( \17497 , \7370 , \4700 );
and \U$16515 ( \17498 , \7168 , \4698 );
nor \U$16516 ( \17499 , \17497 , \17498 );
xnor \U$16517 ( \17500 , \17499 , \4454 );
and \U$16518 ( \17501 , \17496 , \17500 );
and \U$16519 ( \17502 , \7845 , \4305 );
and \U$16520 ( \17503 , \7673 , \4303 );
nor \U$16521 ( \17504 , \17502 , \17503 );
xnor \U$16522 ( \17505 , \17504 , \4118 );
and \U$16523 ( \17506 , \17500 , \17505 );
and \U$16524 ( \17507 , \17496 , \17505 );
or \U$16525 ( \17508 , \17501 , \17506 , \17507 );
and \U$16526 ( \17509 , \8795 , \3992 );
and \U$16527 ( \17510 , \8371 , \3990 );
nor \U$16528 ( \17511 , \17509 , \17510 );
xnor \U$16529 ( \17512 , \17511 , \3787 );
and \U$16530 ( \17513 , \9046 , \3586 );
and \U$16531 ( \17514 , \9041 , \3584 );
nor \U$16532 ( \17515 , \17513 , \17514 );
xnor \U$16533 ( \17516 , \17515 , \3437 );
and \U$16534 ( \17517 , \17512 , \17516 );
and \U$16535 ( \17518 , \9649 , \3264 );
and \U$16536 ( \17519 , \9365 , \3262 );
nor \U$16537 ( \17520 , \17518 , \17519 );
xnor \U$16538 ( \17521 , \17520 , \3122 );
and \U$16539 ( \17522 , \17516 , \17521 );
and \U$16540 ( \17523 , \17512 , \17521 );
or \U$16541 ( \17524 , \17517 , \17522 , \17523 );
and \U$16542 ( \17525 , \17508 , \17524 );
and \U$16543 ( \17526 , \5447 , \6314 );
and \U$16544 ( \17527 , \5439 , \6312 );
nor \U$16545 ( \17528 , \17526 , \17527 );
xnor \U$16546 ( \17529 , \17528 , \6073 );
and \U$16547 ( \17530 , \5921 , \5848 );
and \U$16548 ( \17531 , \5916 , \5846 );
nor \U$16549 ( \17532 , \17530 , \17531 );
xnor \U$16550 ( \17533 , \17532 , \5660 );
and \U$16551 ( \17534 , \17529 , \17533 );
and \U$16552 ( \17535 , \6444 , \5474 );
and \U$16553 ( \17536 , \6185 , \5472 );
nor \U$16554 ( \17537 , \17535 , \17536 );
xnor \U$16555 ( \17538 , \17537 , \5242 );
and \U$16556 ( \17539 , \17533 , \17538 );
and \U$16557 ( \17540 , \17529 , \17538 );
or \U$16558 ( \17541 , \17534 , \17539 , \17540 );
and \U$16559 ( \17542 , \17524 , \17541 );
and \U$16560 ( \17543 , \17508 , \17541 );
or \U$16561 ( \17544 , \17525 , \17542 , \17543 );
and \U$16562 ( \17545 , \4557 , \7906 );
and \U$16563 ( \17546 , \4349 , \7904 );
nor \U$16564 ( \17547 , \17545 , \17546 );
xnor \U$16565 ( \17548 , \17547 , \7646 );
and \U$16566 ( \17549 , \4684 , \7412 );
and \U$16567 ( \17550 , \4679 , \7410 );
nor \U$16568 ( \17551 , \17549 , \17550 );
xnor \U$16569 ( \17552 , \17551 , \7097 );
and \U$16570 ( \17553 , \17548 , \17552 );
and \U$16571 ( \17554 , \5137 , \6903 );
and \U$16572 ( \17555 , \4940 , \6901 );
nor \U$16573 ( \17556 , \17554 , \17555 );
xnor \U$16574 ( \17557 , \17556 , \6563 );
and \U$16575 ( \17558 , \17552 , \17557 );
and \U$16576 ( \17559 , \17548 , \17557 );
or \U$16577 ( \17560 , \17553 , \17558 , \17559 );
and \U$16578 ( \17561 , \3334 , \9564 );
and \U$16579 ( \17562 , \3309 , \9562 );
nor \U$16580 ( \17563 , \17561 , \17562 );
xnor \U$16581 ( \17564 , \17563 , \9193 );
and \U$16582 ( \17565 , \3675 , \9002 );
and \U$16583 ( \17566 , \3508 , \9000 );
nor \U$16584 ( \17567 , \17565 , \17566 );
xnor \U$16585 ( \17568 , \17567 , \8684 );
and \U$16586 ( \17569 , \17564 , \17568 );
and \U$16587 ( \17570 , \3932 , \8435 );
and \U$16588 ( \17571 , \3813 , \8433 );
nor \U$16589 ( \17572 , \17570 , \17571 );
xnor \U$16590 ( \17573 , \17572 , \8186 );
and \U$16591 ( \17574 , \17568 , \17573 );
and \U$16592 ( \17575 , \17564 , \17573 );
or \U$16593 ( \17576 , \17569 , \17574 , \17575 );
and \U$16594 ( \17577 , \17560 , \17576 );
and \U$16595 ( \17578 , \2467 , \11482 );
and \U$16596 ( \17579 , \2459 , \11479 );
nor \U$16597 ( \17580 , \17578 , \17579 );
xnor \U$16598 ( \17581 , \17580 , \10427 );
and \U$16599 ( \17582 , \2715 , \10669 );
and \U$16600 ( \17583 , \2710 , \10667 );
nor \U$16601 ( \17584 , \17582 , \17583 );
xnor \U$16602 ( \17585 , \17584 , \10430 );
and \U$16603 ( \17586 , \17581 , \17585 );
and \U$16604 ( \17587 , \3045 , \10101 );
and \U$16605 ( \17588 , \2901 , \10099 );
nor \U$16606 ( \17589 , \17587 , \17588 );
xnor \U$16607 ( \17590 , \17589 , \9791 );
and \U$16608 ( \17591 , \17585 , \17590 );
and \U$16609 ( \17592 , \17581 , \17590 );
or \U$16610 ( \17593 , \17586 , \17591 , \17592 );
and \U$16611 ( \17594 , \17576 , \17593 );
and \U$16612 ( \17595 , \17560 , \17593 );
or \U$16613 ( \17596 , \17577 , \17594 , \17595 );
and \U$16614 ( \17597 , \17544 , \17596 );
and \U$16615 ( \17598 , \10226 , \2968 );
and \U$16616 ( \17599 , \10218 , \2966 );
nor \U$16617 ( \17600 , \17598 , \17599 );
xnor \U$16618 ( \17601 , \17600 , \2831 );
and \U$16619 ( \17602 , \10834 , \2762 );
and \U$16620 ( \17603 , \10829 , \2760 );
nor \U$16621 ( \17604 , \17602 , \17603 );
xnor \U$16622 ( \17605 , \17604 , \2610 );
and \U$16623 ( \17606 , \17601 , \17605 );
and \U$16624 ( \17607 , \11635 , \2494 );
and \U$16625 ( \17608 , \11015 , \2492 );
nor \U$16626 ( \17609 , \17607 , \17608 );
xnor \U$16627 ( \17610 , \17609 , \2338 );
and \U$16628 ( \17611 , \17605 , \17610 );
and \U$16629 ( \17612 , \17601 , \17610 );
or \U$16630 ( \17613 , \17606 , \17611 , \17612 );
xor \U$16631 ( \17614 , \17386 , \17390 );
xor \U$16632 ( \17615 , \17614 , \17395 );
and \U$16633 ( \17616 , \17613 , \17615 );
xor \U$16634 ( \17617 , \17402 , \17404 );
and \U$16635 ( \17618 , \17615 , \17617 );
and \U$16636 ( \17619 , \17613 , \17617 );
or \U$16637 ( \17620 , \17616 , \17618 , \17619 );
and \U$16638 ( \17621 , \17596 , \17620 );
and \U$16639 ( \17622 , \17544 , \17620 );
or \U$16640 ( \17623 , \17597 , \17621 , \17622 );
xor \U$16641 ( \17624 , \17337 , \17341 );
xor \U$16642 ( \17625 , \17624 , \2109 );
xor \U$16643 ( \17626 , \17349 , \17353 );
xor \U$16644 ( \17627 , \17626 , \17358 );
and \U$16645 ( \17628 , \17625 , \17627 );
xor \U$16646 ( \17629 , \17366 , \17370 );
xor \U$16647 ( \17630 , \17629 , \17375 );
and \U$16648 ( \17631 , \17627 , \17630 );
and \U$16649 ( \17632 , \17625 , \17630 );
or \U$16650 ( \17633 , \17628 , \17631 , \17632 );
xor \U$16651 ( \17634 , \17285 , \17289 );
xor \U$16652 ( \17635 , \17634 , \17294 );
xor \U$16653 ( \17636 , \17301 , \17305 );
xor \U$16654 ( \17637 , \17636 , \17310 );
and \U$16655 ( \17638 , \17635 , \17637 );
xor \U$16656 ( \17639 , \17318 , \17322 );
xor \U$16657 ( \17640 , \17639 , \17327 );
and \U$16658 ( \17641 , \17637 , \17640 );
and \U$16659 ( \17642 , \17635 , \17640 );
or \U$16660 ( \17643 , \17638 , \17641 , \17642 );
and \U$16661 ( \17644 , \17633 , \17643 );
xor \U$16662 ( \17645 , \17054 , \17058 );
xor \U$16663 ( \17646 , \17645 , \17063 );
and \U$16664 ( \17647 , \17643 , \17646 );
and \U$16665 ( \17648 , \17633 , \17646 );
or \U$16666 ( \17649 , \17644 , \17647 , \17648 );
and \U$16667 ( \17650 , \17623 , \17649 );
xor \U$16668 ( \17651 , \17398 , \17405 );
xor \U$16669 ( \17652 , \17651 , \17410 );
xor \U$16670 ( \17653 , \17418 , \17420 );
xor \U$16671 ( \17654 , \17653 , \17423 );
and \U$16672 ( \17655 , \17652 , \17654 );
xor \U$16673 ( \17656 , \17428 , \17430 );
xor \U$16674 ( \17657 , \17656 , \17433 );
and \U$16675 ( \17658 , \17654 , \17657 );
and \U$16676 ( \17659 , \17652 , \17657 );
or \U$16677 ( \17660 , \17655 , \17658 , \17659 );
and \U$16678 ( \17661 , \17649 , \17660 );
and \U$16679 ( \17662 , \17623 , \17660 );
or \U$16680 ( \17663 , \17650 , \17661 , \17662 );
xor \U$16681 ( \17664 , \17066 , \17082 );
xor \U$16682 ( \17665 , \17664 , \17099 );
xor \U$16683 ( \17666 , \17426 , \17436 );
xor \U$16684 ( \17667 , \17666 , \17439 );
and \U$16685 ( \17668 , \17665 , \17667 );
xor \U$16686 ( \17669 , \17445 , \17447 );
xor \U$16687 ( \17670 , \17669 , \17450 );
and \U$16688 ( \17671 , \17667 , \17670 );
and \U$16689 ( \17672 , \17665 , \17670 );
or \U$16690 ( \17673 , \17668 , \17671 , \17672 );
and \U$16691 ( \17674 , \17663 , \17673 );
xor \U$16692 ( \17675 , \17102 , \17154 );
xor \U$16693 ( \17676 , \17675 , \17179 );
and \U$16694 ( \17677 , \17673 , \17676 );
and \U$16695 ( \17678 , \17663 , \17676 );
or \U$16696 ( \17679 , \17674 , \17677 , \17678 );
xor \U$16697 ( \17680 , \17416 , \17442 );
xor \U$16698 ( \17681 , \17680 , \17453 );
xor \U$16699 ( \17682 , \17458 , \17460 );
xor \U$16700 ( \17683 , \17682 , \17463 );
and \U$16701 ( \17684 , \17681 , \17683 );
and \U$16702 ( \17685 , \17679 , \17684 );
xor \U$16703 ( \17686 , \17232 , \17234 );
xor \U$16704 ( \17687 , \17686 , \17237 );
and \U$16705 ( \17688 , \17684 , \17687 );
and \U$16706 ( \17689 , \17679 , \17687 );
or \U$16707 ( \17690 , \17685 , \17688 , \17689 );
xor \U$16708 ( \17691 , \17182 , \17208 );
xor \U$16709 ( \17692 , \17691 , \17219 );
xor \U$16710 ( \17693 , \17456 , \17466 );
xor \U$16711 ( \17694 , \17693 , \17469 );
and \U$16712 ( \17695 , \17692 , \17694 );
and \U$16713 ( \17696 , \17690 , \17695 );
xor \U$16714 ( \17697 , \17472 , \17474 );
xor \U$16715 ( \17698 , \17697 , \17477 );
and \U$16716 ( \17699 , \17695 , \17698 );
and \U$16717 ( \17700 , \17690 , \17698 );
or \U$16718 ( \17701 , \17696 , \17699 , \17700 );
and \U$16719 ( \17702 , \17492 , \17701 );
xor \U$16720 ( \17703 , \17492 , \17701 );
xor \U$16721 ( \17704 , \17690 , \17695 );
xor \U$16722 ( \17705 , \17704 , \17698 );
and \U$16723 ( \17706 , \4349 , \8435 );
and \U$16724 ( \17707 , \3932 , \8433 );
nor \U$16725 ( \17708 , \17706 , \17707 );
xnor \U$16726 ( \17709 , \17708 , \8186 );
and \U$16727 ( \17710 , \4679 , \7906 );
and \U$16728 ( \17711 , \4557 , \7904 );
nor \U$16729 ( \17712 , \17710 , \17711 );
xnor \U$16730 ( \17713 , \17712 , \7646 );
and \U$16731 ( \17714 , \17709 , \17713 );
and \U$16732 ( \17715 , \4940 , \7412 );
and \U$16733 ( \17716 , \4684 , \7410 );
nor \U$16734 ( \17717 , \17715 , \17716 );
xnor \U$16735 ( \17718 , \17717 , \7097 );
and \U$16736 ( \17719 , \17713 , \17718 );
and \U$16737 ( \17720 , \17709 , \17718 );
or \U$16738 ( \17721 , \17714 , \17719 , \17720 );
and \U$16739 ( \17722 , \3309 , \10101 );
and \U$16740 ( \17723 , \3045 , \10099 );
nor \U$16741 ( \17724 , \17722 , \17723 );
xnor \U$16742 ( \17725 , \17724 , \9791 );
and \U$16743 ( \17726 , \3508 , \9564 );
and \U$16744 ( \17727 , \3334 , \9562 );
nor \U$16745 ( \17728 , \17726 , \17727 );
xnor \U$16746 ( \17729 , \17728 , \9193 );
and \U$16747 ( \17730 , \17725 , \17729 );
and \U$16748 ( \17731 , \3813 , \9002 );
and \U$16749 ( \17732 , \3675 , \9000 );
nor \U$16750 ( \17733 , \17731 , \17732 );
xnor \U$16751 ( \17734 , \17733 , \8684 );
and \U$16752 ( \17735 , \17729 , \17734 );
and \U$16753 ( \17736 , \17725 , \17734 );
or \U$16754 ( \17737 , \17730 , \17735 , \17736 );
and \U$16755 ( \17738 , \17721 , \17737 );
and \U$16756 ( \17739 , \2710 , \11482 );
and \U$16757 ( \17740 , \2467 , \11479 );
nor \U$16758 ( \17741 , \17739 , \17740 );
xnor \U$16759 ( \17742 , \17741 , \10427 );
and \U$16760 ( \17743 , \2901 , \10669 );
and \U$16761 ( \17744 , \2715 , \10667 );
nor \U$16762 ( \17745 , \17743 , \17744 );
xnor \U$16763 ( \17746 , \17745 , \10430 );
and \U$16764 ( \17747 , \17742 , \17746 );
and \U$16765 ( \17748 , \17746 , \2338 );
and \U$16766 ( \17749 , \17742 , \2338 );
or \U$16767 ( \17750 , \17747 , \17748 , \17749 );
and \U$16768 ( \17751 , \17737 , \17750 );
and \U$16769 ( \17752 , \17721 , \17750 );
or \U$16770 ( \17753 , \17738 , \17751 , \17752 );
and \U$16771 ( \17754 , \8371 , \4305 );
and \U$16772 ( \17755 , \7845 , \4303 );
nor \U$16773 ( \17756 , \17754 , \17755 );
xnor \U$16774 ( \17757 , \17756 , \4118 );
and \U$16775 ( \17758 , \9041 , \3992 );
and \U$16776 ( \17759 , \8795 , \3990 );
nor \U$16777 ( \17760 , \17758 , \17759 );
xnor \U$16778 ( \17761 , \17760 , \3787 );
and \U$16779 ( \17762 , \17757 , \17761 );
and \U$16780 ( \17763 , \9365 , \3586 );
and \U$16781 ( \17764 , \9046 , \3584 );
nor \U$16782 ( \17765 , \17763 , \17764 );
xnor \U$16783 ( \17766 , \17765 , \3437 );
and \U$16784 ( \17767 , \17761 , \17766 );
and \U$16785 ( \17768 , \17757 , \17766 );
or \U$16786 ( \17769 , \17762 , \17767 , \17768 );
and \U$16787 ( \17770 , \5439 , \6903 );
and \U$16788 ( \17771 , \5137 , \6901 );
nor \U$16789 ( \17772 , \17770 , \17771 );
xnor \U$16790 ( \17773 , \17772 , \6563 );
and \U$16791 ( \17774 , \5916 , \6314 );
and \U$16792 ( \17775 , \5447 , \6312 );
nor \U$16793 ( \17776 , \17774 , \17775 );
xnor \U$16794 ( \17777 , \17776 , \6073 );
and \U$16795 ( \17778 , \17773 , \17777 );
and \U$16796 ( \17779 , \6185 , \5848 );
and \U$16797 ( \17780 , \5921 , \5846 );
nor \U$16798 ( \17781 , \17779 , \17780 );
xnor \U$16799 ( \17782 , \17781 , \5660 );
and \U$16800 ( \17783 , \17777 , \17782 );
and \U$16801 ( \17784 , \17773 , \17782 );
or \U$16802 ( \17785 , \17778 , \17783 , \17784 );
and \U$16803 ( \17786 , \17769 , \17785 );
and \U$16804 ( \17787 , \6816 , \5474 );
and \U$16805 ( \17788 , \6444 , \5472 );
nor \U$16806 ( \17789 , \17787 , \17788 );
xnor \U$16807 ( \17790 , \17789 , \5242 );
and \U$16808 ( \17791 , \7168 , \5023 );
and \U$16809 ( \17792 , \6825 , \5021 );
nor \U$16810 ( \17793 , \17791 , \17792 );
xnor \U$16811 ( \17794 , \17793 , \4880 );
and \U$16812 ( \17795 , \17790 , \17794 );
and \U$16813 ( \17796 , \7673 , \4700 );
and \U$16814 ( \17797 , \7370 , \4698 );
nor \U$16815 ( \17798 , \17796 , \17797 );
xnor \U$16816 ( \17799 , \17798 , \4454 );
and \U$16817 ( \17800 , \17794 , \17799 );
and \U$16818 ( \17801 , \17790 , \17799 );
or \U$16819 ( \17802 , \17795 , \17800 , \17801 );
and \U$16820 ( \17803 , \17785 , \17802 );
and \U$16821 ( \17804 , \17769 , \17802 );
or \U$16822 ( \17805 , \17786 , \17803 , \17804 );
and \U$16823 ( \17806 , \17753 , \17805 );
and \U$16824 ( \17807 , \10218 , \3264 );
and \U$16825 ( \17808 , \9649 , \3262 );
nor \U$16826 ( \17809 , \17807 , \17808 );
xnor \U$16827 ( \17810 , \17809 , \3122 );
and \U$16828 ( \17811 , \10829 , \2968 );
and \U$16829 ( \17812 , \10226 , \2966 );
nor \U$16830 ( \17813 , \17811 , \17812 );
xnor \U$16831 ( \17814 , \17813 , \2831 );
and \U$16832 ( \17815 , \17810 , \17814 );
and \U$16833 ( \17816 , \11015 , \2762 );
and \U$16834 ( \17817 , \10834 , \2760 );
nor \U$16835 ( \17818 , \17816 , \17817 );
xnor \U$16836 ( \17819 , \17818 , \2610 );
and \U$16837 ( \17820 , \17814 , \17819 );
and \U$16838 ( \17821 , \17810 , \17819 );
or \U$16839 ( \17822 , \17815 , \17820 , \17821 );
xor \U$16840 ( \17823 , \17512 , \17516 );
xor \U$16841 ( \17824 , \17823 , \17521 );
and \U$16842 ( \17825 , \17822 , \17824 );
xor \U$16843 ( \17826 , \17601 , \17605 );
xor \U$16844 ( \17827 , \17826 , \17610 );
and \U$16845 ( \17828 , \17824 , \17827 );
and \U$16846 ( \17829 , \17822 , \17827 );
or \U$16847 ( \17830 , \17825 , \17828 , \17829 );
and \U$16848 ( \17831 , \17805 , \17830 );
and \U$16849 ( \17832 , \17753 , \17830 );
or \U$16850 ( \17833 , \17806 , \17831 , \17832 );
xor \U$16851 ( \17834 , \17496 , \17500 );
xor \U$16852 ( \17835 , \17834 , \17505 );
xor \U$16853 ( \17836 , \17548 , \17552 );
xor \U$16854 ( \17837 , \17836 , \17557 );
and \U$16855 ( \17838 , \17835 , \17837 );
xor \U$16856 ( \17839 , \17529 , \17533 );
xor \U$16857 ( \17840 , \17839 , \17538 );
and \U$16858 ( \17841 , \17837 , \17840 );
and \U$16859 ( \17842 , \17835 , \17840 );
or \U$16860 ( \17843 , \17838 , \17841 , \17842 );
xor \U$16861 ( \17844 , \17564 , \17568 );
xor \U$16862 ( \17845 , \17844 , \17573 );
xor \U$16863 ( \17846 , \17581 , \17585 );
xor \U$16864 ( \17847 , \17846 , \17590 );
and \U$16865 ( \17848 , \17845 , \17847 );
and \U$16866 ( \17849 , \17843 , \17848 );
xor \U$16867 ( \17850 , \17625 , \17627 );
xor \U$16868 ( \17851 , \17850 , \17630 );
and \U$16869 ( \17852 , \17848 , \17851 );
and \U$16870 ( \17853 , \17843 , \17851 );
or \U$16871 ( \17854 , \17849 , \17852 , \17853 );
and \U$16872 ( \17855 , \17833 , \17854 );
xor \U$16873 ( \17856 , \17508 , \17524 );
xor \U$16874 ( \17857 , \17856 , \17541 );
xor \U$16875 ( \17858 , \17635 , \17637 );
xor \U$16876 ( \17859 , \17858 , \17640 );
and \U$16877 ( \17860 , \17857 , \17859 );
xor \U$16878 ( \17861 , \17613 , \17615 );
xor \U$16879 ( \17862 , \17861 , \17617 );
and \U$16880 ( \17863 , \17859 , \17862 );
and \U$16881 ( \17864 , \17857 , \17862 );
or \U$16882 ( \17865 , \17860 , \17863 , \17864 );
and \U$16883 ( \17866 , \17854 , \17865 );
and \U$16884 ( \17867 , \17833 , \17865 );
or \U$16885 ( \17868 , \17855 , \17866 , \17867 );
xor \U$16886 ( \17869 , \17297 , \17313 );
xor \U$16887 ( \17870 , \17869 , \17330 );
xor \U$16888 ( \17871 , \17345 , \17361 );
xor \U$16889 ( \17872 , \17871 , \17378 );
and \U$16890 ( \17873 , \17870 , \17872 );
xor \U$16891 ( \17874 , \17652 , \17654 );
xor \U$16892 ( \17875 , \17874 , \17657 );
and \U$16893 ( \17876 , \17872 , \17875 );
and \U$16894 ( \17877 , \17870 , \17875 );
or \U$16895 ( \17878 , \17873 , \17876 , \17877 );
and \U$16896 ( \17879 , \17868 , \17878 );
xor \U$16897 ( \17880 , \17333 , \17381 );
xor \U$16898 ( \17881 , \17880 , \17413 );
and \U$16899 ( \17882 , \17878 , \17881 );
and \U$16900 ( \17883 , \17868 , \17881 );
or \U$16901 ( \17884 , \17879 , \17882 , \17883 );
xor \U$16902 ( \17885 , \17663 , \17673 );
xor \U$16903 ( \17886 , \17885 , \17676 );
and \U$16904 ( \17887 , \17884 , \17886 );
xor \U$16905 ( \17888 , \17681 , \17683 );
and \U$16906 ( \17889 , \17886 , \17888 );
and \U$16907 ( \17890 , \17884 , \17888 );
or \U$16908 ( \17891 , \17887 , \17889 , \17890 );
xor \U$16909 ( \17892 , \17679 , \17684 );
xor \U$16910 ( \17893 , \17892 , \17687 );
and \U$16911 ( \17894 , \17891 , \17893 );
xor \U$16912 ( \17895 , \17692 , \17694 );
and \U$16913 ( \17896 , \17893 , \17895 );
and \U$16914 ( \17897 , \17891 , \17895 );
or \U$16915 ( \17898 , \17894 , \17896 , \17897 );
and \U$16916 ( \17899 , \17705 , \17898 );
xor \U$16917 ( \17900 , \17705 , \17898 );
xor \U$16918 ( \17901 , \17891 , \17893 );
xor \U$16919 ( \17902 , \17901 , \17895 );
and \U$16920 ( \17903 , \2715 , \11482 );
and \U$16921 ( \17904 , \2710 , \11479 );
nor \U$16922 ( \17905 , \17903 , \17904 );
xnor \U$16923 ( \17906 , \17905 , \10427 );
and \U$16924 ( \17907 , \3045 , \10669 );
and \U$16925 ( \17908 , \2901 , \10667 );
nor \U$16926 ( \17909 , \17907 , \17908 );
xnor \U$16927 ( \17910 , \17909 , \10430 );
and \U$16928 ( \17911 , \17906 , \17910 );
and \U$16929 ( \17912 , \3334 , \10101 );
and \U$16930 ( \17913 , \3309 , \10099 );
nor \U$16931 ( \17914 , \17912 , \17913 );
xnor \U$16932 ( \17915 , \17914 , \9791 );
and \U$16933 ( \17916 , \17910 , \17915 );
and \U$16934 ( \17917 , \17906 , \17915 );
or \U$16935 ( \17918 , \17911 , \17916 , \17917 );
and \U$16936 ( \17919 , \3675 , \9564 );
and \U$16937 ( \17920 , \3508 , \9562 );
nor \U$16938 ( \17921 , \17919 , \17920 );
xnor \U$16939 ( \17922 , \17921 , \9193 );
and \U$16940 ( \17923 , \3932 , \9002 );
and \U$16941 ( \17924 , \3813 , \9000 );
nor \U$16942 ( \17925 , \17923 , \17924 );
xnor \U$16943 ( \17926 , \17925 , \8684 );
and \U$16944 ( \17927 , \17922 , \17926 );
and \U$16945 ( \17928 , \4557 , \8435 );
and \U$16946 ( \17929 , \4349 , \8433 );
nor \U$16947 ( \17930 , \17928 , \17929 );
xnor \U$16948 ( \17931 , \17930 , \8186 );
and \U$16949 ( \17932 , \17926 , \17931 );
and \U$16950 ( \17933 , \17922 , \17931 );
or \U$16951 ( \17934 , \17927 , \17932 , \17933 );
and \U$16952 ( \17935 , \17918 , \17934 );
and \U$16953 ( \17936 , \4684 , \7906 );
and \U$16954 ( \17937 , \4679 , \7904 );
nor \U$16955 ( \17938 , \17936 , \17937 );
xnor \U$16956 ( \17939 , \17938 , \7646 );
and \U$16957 ( \17940 , \5137 , \7412 );
and \U$16958 ( \17941 , \4940 , \7410 );
nor \U$16959 ( \17942 , \17940 , \17941 );
xnor \U$16960 ( \17943 , \17942 , \7097 );
and \U$16961 ( \17944 , \17939 , \17943 );
and \U$16962 ( \17945 , \5447 , \6903 );
and \U$16963 ( \17946 , \5439 , \6901 );
nor \U$16964 ( \17947 , \17945 , \17946 );
xnor \U$16965 ( \17948 , \17947 , \6563 );
and \U$16966 ( \17949 , \17943 , \17948 );
and \U$16967 ( \17950 , \17939 , \17948 );
or \U$16968 ( \17951 , \17944 , \17949 , \17950 );
and \U$16969 ( \17952 , \17934 , \17951 );
and \U$16970 ( \17953 , \17918 , \17951 );
or \U$16971 ( \17954 , \17935 , \17952 , \17953 );
and \U$16972 ( \17955 , \7370 , \5023 );
and \U$16973 ( \17956 , \7168 , \5021 );
nor \U$16974 ( \17957 , \17955 , \17956 );
xnor \U$16975 ( \17958 , \17957 , \4880 );
and \U$16976 ( \17959 , \7845 , \4700 );
and \U$16977 ( \17960 , \7673 , \4698 );
nor \U$16978 ( \17961 , \17959 , \17960 );
xnor \U$16979 ( \17962 , \17961 , \4454 );
and \U$16980 ( \17963 , \17958 , \17962 );
and \U$16981 ( \17964 , \8795 , \4305 );
and \U$16982 ( \17965 , \8371 , \4303 );
nor \U$16983 ( \17966 , \17964 , \17965 );
xnor \U$16984 ( \17967 , \17966 , \4118 );
and \U$16985 ( \17968 , \17962 , \17967 );
and \U$16986 ( \17969 , \17958 , \17967 );
or \U$16987 ( \17970 , \17963 , \17968 , \17969 );
and \U$16988 ( \17971 , \5921 , \6314 );
and \U$16989 ( \17972 , \5916 , \6312 );
nor \U$16990 ( \17973 , \17971 , \17972 );
xnor \U$16991 ( \17974 , \17973 , \6073 );
and \U$16992 ( \17975 , \6444 , \5848 );
and \U$16993 ( \17976 , \6185 , \5846 );
nor \U$16994 ( \17977 , \17975 , \17976 );
xnor \U$16995 ( \17978 , \17977 , \5660 );
and \U$16996 ( \17979 , \17974 , \17978 );
and \U$16997 ( \17980 , \6825 , \5474 );
and \U$16998 ( \17981 , \6816 , \5472 );
nor \U$16999 ( \17982 , \17980 , \17981 );
xnor \U$17000 ( \17983 , \17982 , \5242 );
and \U$17001 ( \17984 , \17978 , \17983 );
and \U$17002 ( \17985 , \17974 , \17983 );
or \U$17003 ( \17986 , \17979 , \17984 , \17985 );
and \U$17004 ( \17987 , \17970 , \17986 );
and \U$17005 ( \17988 , \9046 , \3992 );
and \U$17006 ( \17989 , \9041 , \3990 );
nor \U$17007 ( \17990 , \17988 , \17989 );
xnor \U$17008 ( \17991 , \17990 , \3787 );
and \U$17009 ( \17992 , \9649 , \3586 );
and \U$17010 ( \17993 , \9365 , \3584 );
nor \U$17011 ( \17994 , \17992 , \17993 );
xnor \U$17012 ( \17995 , \17994 , \3437 );
and \U$17013 ( \17996 , \17991 , \17995 );
and \U$17014 ( \17997 , \10226 , \3264 );
and \U$17015 ( \17998 , \10218 , \3262 );
nor \U$17016 ( \17999 , \17997 , \17998 );
xnor \U$17017 ( \18000 , \17999 , \3122 );
and \U$17018 ( \18001 , \17995 , \18000 );
and \U$17019 ( \18002 , \17991 , \18000 );
or \U$17020 ( \18003 , \17996 , \18001 , \18002 );
and \U$17021 ( \18004 , \17986 , \18003 );
and \U$17022 ( \18005 , \17970 , \18003 );
or \U$17023 ( \18006 , \17987 , \18004 , \18005 );
and \U$17024 ( \18007 , \17954 , \18006 );
nand \U$17025 ( \18008 , \11635 , \2492 );
xnor \U$17026 ( \18009 , \18008 , \2338 );
xor \U$17027 ( \18010 , \17757 , \17761 );
xor \U$17028 ( \18011 , \18010 , \17766 );
and \U$17029 ( \18012 , \18009 , \18011 );
xor \U$17030 ( \18013 , \17810 , \17814 );
xor \U$17031 ( \18014 , \18013 , \17819 );
and \U$17032 ( \18015 , \18011 , \18014 );
and \U$17033 ( \18016 , \18009 , \18014 );
or \U$17034 ( \18017 , \18012 , \18015 , \18016 );
and \U$17035 ( \18018 , \18006 , \18017 );
and \U$17036 ( \18019 , \17954 , \18017 );
or \U$17037 ( \18020 , \18007 , \18018 , \18019 );
xor \U$17038 ( \18021 , \17721 , \17737 );
xor \U$17039 ( \18022 , \18021 , \17750 );
xor \U$17040 ( \18023 , \17769 , \17785 );
xor \U$17041 ( \18024 , \18023 , \17802 );
and \U$17042 ( \18025 , \18022 , \18024 );
xor \U$17043 ( \18026 , \17822 , \17824 );
xor \U$17044 ( \18027 , \18026 , \17827 );
and \U$17045 ( \18028 , \18024 , \18027 );
and \U$17046 ( \18029 , \18022 , \18027 );
or \U$17047 ( \18030 , \18025 , \18028 , \18029 );
and \U$17048 ( \18031 , \18020 , \18030 );
xor \U$17049 ( \18032 , \17709 , \17713 );
xor \U$17050 ( \18033 , \18032 , \17718 );
xor \U$17051 ( \18034 , \17773 , \17777 );
xor \U$17052 ( \18035 , \18034 , \17782 );
and \U$17053 ( \18036 , \18033 , \18035 );
xor \U$17054 ( \18037 , \17790 , \17794 );
xor \U$17055 ( \18038 , \18037 , \17799 );
and \U$17056 ( \18039 , \18035 , \18038 );
and \U$17057 ( \18040 , \18033 , \18038 );
or \U$17058 ( \18041 , \18036 , \18039 , \18040 );
xor \U$17059 ( \18042 , \17835 , \17837 );
xor \U$17060 ( \18043 , \18042 , \17840 );
and \U$17061 ( \18044 , \18041 , \18043 );
xor \U$17062 ( \18045 , \17845 , \17847 );
and \U$17063 ( \18046 , \18043 , \18045 );
and \U$17064 ( \18047 , \18041 , \18045 );
or \U$17065 ( \18048 , \18044 , \18046 , \18047 );
and \U$17066 ( \18049 , \18030 , \18048 );
and \U$17067 ( \18050 , \18020 , \18048 );
or \U$17068 ( \18051 , \18031 , \18049 , \18050 );
xor \U$17069 ( \18052 , \17560 , \17576 );
xor \U$17070 ( \18053 , \18052 , \17593 );
xor \U$17071 ( \18054 , \17843 , \17848 );
xor \U$17072 ( \18055 , \18054 , \17851 );
and \U$17073 ( \18056 , \18053 , \18055 );
xor \U$17074 ( \18057 , \17857 , \17859 );
xor \U$17075 ( \18058 , \18057 , \17862 );
and \U$17076 ( \18059 , \18055 , \18058 );
and \U$17077 ( \18060 , \18053 , \18058 );
or \U$17078 ( \18061 , \18056 , \18059 , \18060 );
and \U$17079 ( \18062 , \18051 , \18061 );
xor \U$17080 ( \18063 , \17633 , \17643 );
xor \U$17081 ( \18064 , \18063 , \17646 );
and \U$17082 ( \18065 , \18061 , \18064 );
and \U$17083 ( \18066 , \18051 , \18064 );
or \U$17084 ( \18067 , \18062 , \18065 , \18066 );
xor \U$17085 ( \18068 , \17544 , \17596 );
xor \U$17086 ( \18069 , \18068 , \17620 );
xor \U$17087 ( \18070 , \17833 , \17854 );
xor \U$17088 ( \18071 , \18070 , \17865 );
and \U$17089 ( \18072 , \18069 , \18071 );
xor \U$17090 ( \18073 , \17870 , \17872 );
xor \U$17091 ( \18074 , \18073 , \17875 );
and \U$17092 ( \18075 , \18071 , \18074 );
and \U$17093 ( \18076 , \18069 , \18074 );
or \U$17094 ( \18077 , \18072 , \18075 , \18076 );
and \U$17095 ( \18078 , \18067 , \18077 );
xor \U$17096 ( \18079 , \17665 , \17667 );
xor \U$17097 ( \18080 , \18079 , \17670 );
and \U$17098 ( \18081 , \18077 , \18080 );
and \U$17099 ( \18082 , \18067 , \18080 );
or \U$17100 ( \18083 , \18078 , \18081 , \18082 );
xor \U$17101 ( \18084 , \17623 , \17649 );
xor \U$17102 ( \18085 , \18084 , \17660 );
xor \U$17103 ( \18086 , \17868 , \17878 );
xor \U$17104 ( \18087 , \18086 , \17881 );
and \U$17105 ( \18088 , \18085 , \18087 );
and \U$17106 ( \18089 , \18083 , \18088 );
xor \U$17107 ( \18090 , \17884 , \17886 );
xor \U$17108 ( \18091 , \18090 , \17888 );
and \U$17109 ( \18092 , \18088 , \18091 );
and \U$17110 ( \18093 , \18083 , \18091 );
or \U$17111 ( \18094 , \18089 , \18092 , \18093 );
and \U$17112 ( \18095 , \17902 , \18094 );
xor \U$17113 ( \18096 , \17902 , \18094 );
xor \U$17114 ( \18097 , \18083 , \18088 );
xor \U$17115 ( \18098 , \18097 , \18091 );
and \U$17116 ( \18099 , \2901 , \11482 );
and \U$17117 ( \18100 , \2715 , \11479 );
nor \U$17118 ( \18101 , \18099 , \18100 );
xnor \U$17119 ( \18102 , \18101 , \10427 );
and \U$17120 ( \18103 , \3309 , \10669 );
and \U$17121 ( \18104 , \3045 , \10667 );
nor \U$17122 ( \18105 , \18103 , \18104 );
xnor \U$17123 ( \18106 , \18105 , \10430 );
and \U$17124 ( \18107 , \18102 , \18106 );
and \U$17125 ( \18108 , \18106 , \2610 );
and \U$17126 ( \18109 , \18102 , \2610 );
or \U$17127 ( \18110 , \18107 , \18108 , \18109 );
and \U$17128 ( \18111 , \4679 , \8435 );
and \U$17129 ( \18112 , \4557 , \8433 );
nor \U$17130 ( \18113 , \18111 , \18112 );
xnor \U$17131 ( \18114 , \18113 , \8186 );
and \U$17132 ( \18115 , \4940 , \7906 );
and \U$17133 ( \18116 , \4684 , \7904 );
nor \U$17134 ( \18117 , \18115 , \18116 );
xnor \U$17135 ( \18118 , \18117 , \7646 );
and \U$17136 ( \18119 , \18114 , \18118 );
and \U$17137 ( \18120 , \5439 , \7412 );
and \U$17138 ( \18121 , \5137 , \7410 );
nor \U$17139 ( \18122 , \18120 , \18121 );
xnor \U$17140 ( \18123 , \18122 , \7097 );
and \U$17141 ( \18124 , \18118 , \18123 );
and \U$17142 ( \18125 , \18114 , \18123 );
or \U$17143 ( \18126 , \18119 , \18124 , \18125 );
and \U$17144 ( \18127 , \18110 , \18126 );
and \U$17145 ( \18128 , \3508 , \10101 );
and \U$17146 ( \18129 , \3334 , \10099 );
nor \U$17147 ( \18130 , \18128 , \18129 );
xnor \U$17148 ( \18131 , \18130 , \9791 );
and \U$17149 ( \18132 , \3813 , \9564 );
and \U$17150 ( \18133 , \3675 , \9562 );
nor \U$17151 ( \18134 , \18132 , \18133 );
xnor \U$17152 ( \18135 , \18134 , \9193 );
and \U$17153 ( \18136 , \18131 , \18135 );
and \U$17154 ( \18137 , \4349 , \9002 );
and \U$17155 ( \18138 , \3932 , \9000 );
nor \U$17156 ( \18139 , \18137 , \18138 );
xnor \U$17157 ( \18140 , \18139 , \8684 );
and \U$17158 ( \18141 , \18135 , \18140 );
and \U$17159 ( \18142 , \18131 , \18140 );
or \U$17160 ( \18143 , \18136 , \18141 , \18142 );
and \U$17161 ( \18144 , \18126 , \18143 );
and \U$17162 ( \18145 , \18110 , \18143 );
or \U$17163 ( \18146 , \18127 , \18144 , \18145 );
and \U$17164 ( \18147 , \10829 , \3264 );
and \U$17165 ( \18148 , \10226 , \3262 );
nor \U$17166 ( \18149 , \18147 , \18148 );
xnor \U$17167 ( \18150 , \18149 , \3122 );
and \U$17168 ( \18151 , \11015 , \2968 );
and \U$17169 ( \18152 , \10834 , \2966 );
nor \U$17170 ( \18153 , \18151 , \18152 );
xnor \U$17171 ( \18154 , \18153 , \2831 );
and \U$17172 ( \18155 , \18150 , \18154 );
nand \U$17173 ( \18156 , \11635 , \2760 );
xnor \U$17174 ( \18157 , \18156 , \2610 );
and \U$17175 ( \18158 , \18154 , \18157 );
and \U$17176 ( \18159 , \18150 , \18157 );
or \U$17177 ( \18160 , \18155 , \18158 , \18159 );
and \U$17178 ( \18161 , \10834 , \2968 );
and \U$17179 ( \18162 , \10829 , \2966 );
nor \U$17180 ( \18163 , \18161 , \18162 );
xnor \U$17181 ( \18164 , \18163 , \2831 );
and \U$17182 ( \18165 , \18160 , \18164 );
and \U$17183 ( \18166 , \11635 , \2762 );
and \U$17184 ( \18167 , \11015 , \2760 );
nor \U$17185 ( \18168 , \18166 , \18167 );
xnor \U$17186 ( \18169 , \18168 , \2610 );
and \U$17187 ( \18170 , \18164 , \18169 );
and \U$17188 ( \18171 , \18160 , \18169 );
or \U$17189 ( \18172 , \18165 , \18170 , \18171 );
and \U$17190 ( \18173 , \18146 , \18172 );
and \U$17191 ( \18174 , \5916 , \6903 );
and \U$17192 ( \18175 , \5447 , \6901 );
nor \U$17193 ( \18176 , \18174 , \18175 );
xnor \U$17194 ( \18177 , \18176 , \6563 );
and \U$17195 ( \18178 , \6185 , \6314 );
and \U$17196 ( \18179 , \5921 , \6312 );
nor \U$17197 ( \18180 , \18178 , \18179 );
xnor \U$17198 ( \18181 , \18180 , \6073 );
and \U$17199 ( \18182 , \18177 , \18181 );
and \U$17200 ( \18183 , \6816 , \5848 );
and \U$17201 ( \18184 , \6444 , \5846 );
nor \U$17202 ( \18185 , \18183 , \18184 );
xnor \U$17203 ( \18186 , \18185 , \5660 );
and \U$17204 ( \18187 , \18181 , \18186 );
and \U$17205 ( \18188 , \18177 , \18186 );
or \U$17206 ( \18189 , \18182 , \18187 , \18188 );
and \U$17207 ( \18190 , \9041 , \4305 );
and \U$17208 ( \18191 , \8795 , \4303 );
nor \U$17209 ( \18192 , \18190 , \18191 );
xnor \U$17210 ( \18193 , \18192 , \4118 );
and \U$17211 ( \18194 , \9365 , \3992 );
and \U$17212 ( \18195 , \9046 , \3990 );
nor \U$17213 ( \18196 , \18194 , \18195 );
xnor \U$17214 ( \18197 , \18196 , \3787 );
and \U$17215 ( \18198 , \18193 , \18197 );
and \U$17216 ( \18199 , \10218 , \3586 );
and \U$17217 ( \18200 , \9649 , \3584 );
nor \U$17218 ( \18201 , \18199 , \18200 );
xnor \U$17219 ( \18202 , \18201 , \3437 );
and \U$17220 ( \18203 , \18197 , \18202 );
and \U$17221 ( \18204 , \18193 , \18202 );
or \U$17222 ( \18205 , \18198 , \18203 , \18204 );
and \U$17223 ( \18206 , \18189 , \18205 );
and \U$17224 ( \18207 , \7168 , \5474 );
and \U$17225 ( \18208 , \6825 , \5472 );
nor \U$17226 ( \18209 , \18207 , \18208 );
xnor \U$17227 ( \18210 , \18209 , \5242 );
and \U$17228 ( \18211 , \7673 , \5023 );
and \U$17229 ( \18212 , \7370 , \5021 );
nor \U$17230 ( \18213 , \18211 , \18212 );
xnor \U$17231 ( \18214 , \18213 , \4880 );
and \U$17232 ( \18215 , \18210 , \18214 );
and \U$17233 ( \18216 , \8371 , \4700 );
and \U$17234 ( \18217 , \7845 , \4698 );
nor \U$17235 ( \18218 , \18216 , \18217 );
xnor \U$17236 ( \18219 , \18218 , \4454 );
and \U$17237 ( \18220 , \18214 , \18219 );
and \U$17238 ( \18221 , \18210 , \18219 );
or \U$17239 ( \18222 , \18215 , \18220 , \18221 );
and \U$17240 ( \18223 , \18205 , \18222 );
and \U$17241 ( \18224 , \18189 , \18222 );
or \U$17242 ( \18225 , \18206 , \18223 , \18224 );
and \U$17243 ( \18226 , \18172 , \18225 );
and \U$17244 ( \18227 , \18146 , \18225 );
or \U$17245 ( \18228 , \18173 , \18226 , \18227 );
xor \U$17246 ( \18229 , \17906 , \17910 );
xor \U$17247 ( \18230 , \18229 , \17915 );
xor \U$17248 ( \18231 , \17922 , \17926 );
xor \U$17249 ( \18232 , \18231 , \17931 );
and \U$17250 ( \18233 , \18230 , \18232 );
xor \U$17251 ( \18234 , \17939 , \17943 );
xor \U$17252 ( \18235 , \18234 , \17948 );
and \U$17253 ( \18236 , \18232 , \18235 );
and \U$17254 ( \18237 , \18230 , \18235 );
or \U$17255 ( \18238 , \18233 , \18236 , \18237 );
xor \U$17256 ( \18239 , \17958 , \17962 );
xor \U$17257 ( \18240 , \18239 , \17967 );
xor \U$17258 ( \18241 , \17974 , \17978 );
xor \U$17259 ( \18242 , \18241 , \17983 );
and \U$17260 ( \18243 , \18240 , \18242 );
xor \U$17261 ( \18244 , \17991 , \17995 );
xor \U$17262 ( \18245 , \18244 , \18000 );
and \U$17263 ( \18246 , \18242 , \18245 );
and \U$17264 ( \18247 , \18240 , \18245 );
or \U$17265 ( \18248 , \18243 , \18246 , \18247 );
and \U$17266 ( \18249 , \18238 , \18248 );
xor \U$17267 ( \18250 , \17725 , \17729 );
xor \U$17268 ( \18251 , \18250 , \17734 );
and \U$17269 ( \18252 , \18248 , \18251 );
and \U$17270 ( \18253 , \18238 , \18251 );
or \U$17271 ( \18254 , \18249 , \18252 , \18253 );
and \U$17272 ( \18255 , \18228 , \18254 );
xor \U$17273 ( \18256 , \17742 , \17746 );
xor \U$17274 ( \18257 , \18256 , \2338 );
xor \U$17275 ( \18258 , \18033 , \18035 );
xor \U$17276 ( \18259 , \18258 , \18038 );
and \U$17277 ( \18260 , \18257 , \18259 );
xor \U$17278 ( \18261 , \18009 , \18011 );
xor \U$17279 ( \18262 , \18261 , \18014 );
and \U$17280 ( \18263 , \18259 , \18262 );
and \U$17281 ( \18264 , \18257 , \18262 );
or \U$17282 ( \18265 , \18260 , \18263 , \18264 );
and \U$17283 ( \18266 , \18254 , \18265 );
and \U$17284 ( \18267 , \18228 , \18265 );
or \U$17285 ( \18268 , \18255 , \18266 , \18267 );
xor \U$17286 ( \18269 , \17954 , \18006 );
xor \U$17287 ( \18270 , \18269 , \18017 );
xor \U$17288 ( \18271 , \18022 , \18024 );
xor \U$17289 ( \18272 , \18271 , \18027 );
and \U$17290 ( \18273 , \18270 , \18272 );
xor \U$17291 ( \18274 , \18041 , \18043 );
xor \U$17292 ( \18275 , \18274 , \18045 );
and \U$17293 ( \18276 , \18272 , \18275 );
and \U$17294 ( \18277 , \18270 , \18275 );
or \U$17295 ( \18278 , \18273 , \18276 , \18277 );
and \U$17296 ( \18279 , \18268 , \18278 );
xor \U$17297 ( \18280 , \17753 , \17805 );
xor \U$17298 ( \18281 , \18280 , \17830 );
and \U$17299 ( \18282 , \18278 , \18281 );
and \U$17300 ( \18283 , \18268 , \18281 );
or \U$17301 ( \18284 , \18279 , \18282 , \18283 );
xor \U$17302 ( \18285 , \18020 , \18030 );
xor \U$17303 ( \18286 , \18285 , \18048 );
xor \U$17304 ( \18287 , \18053 , \18055 );
xor \U$17305 ( \18288 , \18287 , \18058 );
and \U$17306 ( \18289 , \18286 , \18288 );
and \U$17307 ( \18290 , \18284 , \18289 );
xor \U$17308 ( \18291 , \18069 , \18071 );
xor \U$17309 ( \18292 , \18291 , \18074 );
and \U$17310 ( \18293 , \18289 , \18292 );
and \U$17311 ( \18294 , \18284 , \18292 );
or \U$17312 ( \18295 , \18290 , \18293 , \18294 );
xor \U$17313 ( \18296 , \18067 , \18077 );
xor \U$17314 ( \18297 , \18296 , \18080 );
and \U$17315 ( \18298 , \18295 , \18297 );
xor \U$17316 ( \18299 , \18085 , \18087 );
and \U$17317 ( \18300 , \18297 , \18299 );
and \U$17318 ( \18301 , \18295 , \18299 );
or \U$17319 ( \18302 , \18298 , \18300 , \18301 );
and \U$17320 ( \18303 , \18098 , \18302 );
xor \U$17321 ( \18304 , \18098 , \18302 );
xor \U$17322 ( \18305 , \18295 , \18297 );
xor \U$17323 ( \18306 , \18305 , \18299 );
and \U$17324 ( \18307 , \9649 , \3992 );
and \U$17325 ( \18308 , \9365 , \3990 );
nor \U$17326 ( \18309 , \18307 , \18308 );
xnor \U$17327 ( \18310 , \18309 , \3787 );
and \U$17328 ( \18311 , \10226 , \3586 );
and \U$17329 ( \18312 , \10218 , \3584 );
nor \U$17330 ( \18313 , \18311 , \18312 );
xnor \U$17331 ( \18314 , \18313 , \3437 );
and \U$17332 ( \18315 , \18310 , \18314 );
and \U$17333 ( \18316 , \10834 , \3264 );
and \U$17334 ( \18317 , \10829 , \3262 );
nor \U$17335 ( \18318 , \18316 , \18317 );
xnor \U$17336 ( \18319 , \18318 , \3122 );
and \U$17337 ( \18320 , \18314 , \18319 );
and \U$17338 ( \18321 , \18310 , \18319 );
or \U$17339 ( \18322 , \18315 , \18320 , \18321 );
and \U$17340 ( \18323 , \6444 , \6314 );
and \U$17341 ( \18324 , \6185 , \6312 );
nor \U$17342 ( \18325 , \18323 , \18324 );
xnor \U$17343 ( \18326 , \18325 , \6073 );
and \U$17344 ( \18327 , \6825 , \5848 );
and \U$17345 ( \18328 , \6816 , \5846 );
nor \U$17346 ( \18329 , \18327 , \18328 );
xnor \U$17347 ( \18330 , \18329 , \5660 );
and \U$17348 ( \18331 , \18326 , \18330 );
and \U$17349 ( \18332 , \7370 , \5474 );
and \U$17350 ( \18333 , \7168 , \5472 );
nor \U$17351 ( \18334 , \18332 , \18333 );
xnor \U$17352 ( \18335 , \18334 , \5242 );
and \U$17353 ( \18336 , \18330 , \18335 );
and \U$17354 ( \18337 , \18326 , \18335 );
or \U$17355 ( \18338 , \18331 , \18336 , \18337 );
and \U$17356 ( \18339 , \18322 , \18338 );
and \U$17357 ( \18340 , \7845 , \5023 );
and \U$17358 ( \18341 , \7673 , \5021 );
nor \U$17359 ( \18342 , \18340 , \18341 );
xnor \U$17360 ( \18343 , \18342 , \4880 );
and \U$17361 ( \18344 , \8795 , \4700 );
and \U$17362 ( \18345 , \8371 , \4698 );
nor \U$17363 ( \18346 , \18344 , \18345 );
xnor \U$17364 ( \18347 , \18346 , \4454 );
and \U$17365 ( \18348 , \18343 , \18347 );
and \U$17366 ( \18349 , \9046 , \4305 );
and \U$17367 ( \18350 , \9041 , \4303 );
nor \U$17368 ( \18351 , \18349 , \18350 );
xnor \U$17369 ( \18352 , \18351 , \4118 );
and \U$17370 ( \18353 , \18347 , \18352 );
and \U$17371 ( \18354 , \18343 , \18352 );
or \U$17372 ( \18355 , \18348 , \18353 , \18354 );
and \U$17373 ( \18356 , \18338 , \18355 );
and \U$17374 ( \18357 , \18322 , \18355 );
or \U$17375 ( \18358 , \18339 , \18356 , \18357 );
and \U$17376 ( \18359 , \5137 , \7906 );
and \U$17377 ( \18360 , \4940 , \7904 );
nor \U$17378 ( \18361 , \18359 , \18360 );
xnor \U$17379 ( \18362 , \18361 , \7646 );
and \U$17380 ( \18363 , \5447 , \7412 );
and \U$17381 ( \18364 , \5439 , \7410 );
nor \U$17382 ( \18365 , \18363 , \18364 );
xnor \U$17383 ( \18366 , \18365 , \7097 );
and \U$17384 ( \18367 , \18362 , \18366 );
and \U$17385 ( \18368 , \5921 , \6903 );
and \U$17386 ( \18369 , \5916 , \6901 );
nor \U$17387 ( \18370 , \18368 , \18369 );
xnor \U$17388 ( \18371 , \18370 , \6563 );
and \U$17389 ( \18372 , \18366 , \18371 );
and \U$17390 ( \18373 , \18362 , \18371 );
or \U$17391 ( \18374 , \18367 , \18372 , \18373 );
and \U$17392 ( \18375 , \3932 , \9564 );
and \U$17393 ( \18376 , \3813 , \9562 );
nor \U$17394 ( \18377 , \18375 , \18376 );
xnor \U$17395 ( \18378 , \18377 , \9193 );
and \U$17396 ( \18379 , \4557 , \9002 );
and \U$17397 ( \18380 , \4349 , \9000 );
nor \U$17398 ( \18381 , \18379 , \18380 );
xnor \U$17399 ( \18382 , \18381 , \8684 );
and \U$17400 ( \18383 , \18378 , \18382 );
and \U$17401 ( \18384 , \4684 , \8435 );
and \U$17402 ( \18385 , \4679 , \8433 );
nor \U$17403 ( \18386 , \18384 , \18385 );
xnor \U$17404 ( \18387 , \18386 , \8186 );
and \U$17405 ( \18388 , \18382 , \18387 );
and \U$17406 ( \18389 , \18378 , \18387 );
or \U$17407 ( \18390 , \18383 , \18388 , \18389 );
and \U$17408 ( \18391 , \18374 , \18390 );
and \U$17409 ( \18392 , \3045 , \11482 );
and \U$17410 ( \18393 , \2901 , \11479 );
nor \U$17411 ( \18394 , \18392 , \18393 );
xnor \U$17412 ( \18395 , \18394 , \10427 );
and \U$17413 ( \18396 , \3334 , \10669 );
and \U$17414 ( \18397 , \3309 , \10667 );
nor \U$17415 ( \18398 , \18396 , \18397 );
xnor \U$17416 ( \18399 , \18398 , \10430 );
and \U$17417 ( \18400 , \18395 , \18399 );
and \U$17418 ( \18401 , \3675 , \10101 );
and \U$17419 ( \18402 , \3508 , \10099 );
nor \U$17420 ( \18403 , \18401 , \18402 );
xnor \U$17421 ( \18404 , \18403 , \9791 );
and \U$17422 ( \18405 , \18399 , \18404 );
and \U$17423 ( \18406 , \18395 , \18404 );
or \U$17424 ( \18407 , \18400 , \18405 , \18406 );
and \U$17425 ( \18408 , \18390 , \18407 );
and \U$17426 ( \18409 , \18374 , \18407 );
or \U$17427 ( \18410 , \18391 , \18408 , \18409 );
and \U$17428 ( \18411 , \18358 , \18410 );
xor \U$17429 ( \18412 , \18150 , \18154 );
xor \U$17430 ( \18413 , \18412 , \18157 );
xor \U$17431 ( \18414 , \18193 , \18197 );
xor \U$17432 ( \18415 , \18414 , \18202 );
and \U$17433 ( \18416 , \18413 , \18415 );
xor \U$17434 ( \18417 , \18210 , \18214 );
xor \U$17435 ( \18418 , \18417 , \18219 );
and \U$17436 ( \18419 , \18415 , \18418 );
and \U$17437 ( \18420 , \18413 , \18418 );
or \U$17438 ( \18421 , \18416 , \18419 , \18420 );
and \U$17439 ( \18422 , \18410 , \18421 );
and \U$17440 ( \18423 , \18358 , \18421 );
or \U$17441 ( \18424 , \18411 , \18422 , \18423 );
xor \U$17442 ( \18425 , \18110 , \18126 );
xor \U$17443 ( \18426 , \18425 , \18143 );
xor \U$17444 ( \18427 , \18160 , \18164 );
xor \U$17445 ( \18428 , \18427 , \18169 );
and \U$17446 ( \18429 , \18426 , \18428 );
xor \U$17447 ( \18430 , \18189 , \18205 );
xor \U$17448 ( \18431 , \18430 , \18222 );
and \U$17449 ( \18432 , \18428 , \18431 );
and \U$17450 ( \18433 , \18426 , \18431 );
or \U$17451 ( \18434 , \18429 , \18432 , \18433 );
and \U$17452 ( \18435 , \18424 , \18434 );
xor \U$17453 ( \18436 , \18177 , \18181 );
xor \U$17454 ( \18437 , \18436 , \18186 );
xor \U$17455 ( \18438 , \18114 , \18118 );
xor \U$17456 ( \18439 , \18438 , \18123 );
and \U$17457 ( \18440 , \18437 , \18439 );
xor \U$17458 ( \18441 , \18131 , \18135 );
xor \U$17459 ( \18442 , \18441 , \18140 );
and \U$17460 ( \18443 , \18439 , \18442 );
and \U$17461 ( \18444 , \18437 , \18442 );
or \U$17462 ( \18445 , \18440 , \18443 , \18444 );
xor \U$17463 ( \18446 , \18230 , \18232 );
xor \U$17464 ( \18447 , \18446 , \18235 );
and \U$17465 ( \18448 , \18445 , \18447 );
xor \U$17466 ( \18449 , \18240 , \18242 );
xor \U$17467 ( \18450 , \18449 , \18245 );
and \U$17468 ( \18451 , \18447 , \18450 );
and \U$17469 ( \18452 , \18445 , \18450 );
or \U$17470 ( \18453 , \18448 , \18451 , \18452 );
and \U$17471 ( \18454 , \18434 , \18453 );
and \U$17472 ( \18455 , \18424 , \18453 );
or \U$17473 ( \18456 , \18435 , \18454 , \18455 );
xor \U$17474 ( \18457 , \17918 , \17934 );
xor \U$17475 ( \18458 , \18457 , \17951 );
xor \U$17476 ( \18459 , \17970 , \17986 );
xor \U$17477 ( \18460 , \18459 , \18003 );
and \U$17478 ( \18461 , \18458 , \18460 );
xor \U$17479 ( \18462 , \18257 , \18259 );
xor \U$17480 ( \18463 , \18462 , \18262 );
and \U$17481 ( \18464 , \18460 , \18463 );
and \U$17482 ( \18465 , \18458 , \18463 );
or \U$17483 ( \18466 , \18461 , \18464 , \18465 );
and \U$17484 ( \18467 , \18456 , \18466 );
xor \U$17485 ( \18468 , \18270 , \18272 );
xor \U$17486 ( \18469 , \18468 , \18275 );
and \U$17487 ( \18470 , \18466 , \18469 );
and \U$17488 ( \18471 , \18456 , \18469 );
or \U$17489 ( \18472 , \18467 , \18470 , \18471 );
xor \U$17490 ( \18473 , \18268 , \18278 );
xor \U$17491 ( \18474 , \18473 , \18281 );
and \U$17492 ( \18475 , \18472 , \18474 );
xor \U$17493 ( \18476 , \18286 , \18288 );
and \U$17494 ( \18477 , \18474 , \18476 );
and \U$17495 ( \18478 , \18472 , \18476 );
or \U$17496 ( \18479 , \18475 , \18477 , \18478 );
xor \U$17497 ( \18480 , \18051 , \18061 );
xor \U$17498 ( \18481 , \18480 , \18064 );
and \U$17499 ( \18482 , \18479 , \18481 );
xor \U$17500 ( \18483 , \18284 , \18289 );
xor \U$17501 ( \18484 , \18483 , \18292 );
and \U$17502 ( \18485 , \18481 , \18484 );
and \U$17503 ( \18486 , \18479 , \18484 );
or \U$17504 ( \18487 , \18482 , \18485 , \18486 );
and \U$17505 ( \18488 , \18306 , \18487 );
xor \U$17506 ( \18489 , \18306 , \18487 );
xor \U$17507 ( \18490 , \18479 , \18481 );
xor \U$17508 ( \18491 , \18490 , \18484 );
and \U$17509 ( \18492 , \4940 , \8435 );
and \U$17510 ( \18493 , \4684 , \8433 );
nor \U$17511 ( \18494 , \18492 , \18493 );
xnor \U$17512 ( \18495 , \18494 , \8186 );
and \U$17513 ( \18496 , \5439 , \7906 );
and \U$17514 ( \18497 , \5137 , \7904 );
nor \U$17515 ( \18498 , \18496 , \18497 );
xnor \U$17516 ( \18499 , \18498 , \7646 );
and \U$17517 ( \18500 , \18495 , \18499 );
and \U$17518 ( \18501 , \5916 , \7412 );
and \U$17519 ( \18502 , \5447 , \7410 );
nor \U$17520 ( \18503 , \18501 , \18502 );
xnor \U$17521 ( \18504 , \18503 , \7097 );
and \U$17522 ( \18505 , \18499 , \18504 );
and \U$17523 ( \18506 , \18495 , \18504 );
or \U$17524 ( \18507 , \18500 , \18505 , \18506 );
and \U$17525 ( \18508 , \3813 , \10101 );
and \U$17526 ( \18509 , \3675 , \10099 );
nor \U$17527 ( \18510 , \18508 , \18509 );
xnor \U$17528 ( \18511 , \18510 , \9791 );
and \U$17529 ( \18512 , \4349 , \9564 );
and \U$17530 ( \18513 , \3932 , \9562 );
nor \U$17531 ( \18514 , \18512 , \18513 );
xnor \U$17532 ( \18515 , \18514 , \9193 );
and \U$17533 ( \18516 , \18511 , \18515 );
and \U$17534 ( \18517 , \4679 , \9002 );
and \U$17535 ( \18518 , \4557 , \9000 );
nor \U$17536 ( \18519 , \18517 , \18518 );
xnor \U$17537 ( \18520 , \18519 , \8684 );
and \U$17538 ( \18521 , \18515 , \18520 );
and \U$17539 ( \18522 , \18511 , \18520 );
or \U$17540 ( \18523 , \18516 , \18521 , \18522 );
and \U$17541 ( \18524 , \18507 , \18523 );
and \U$17542 ( \18525 , \3309 , \11482 );
and \U$17543 ( \18526 , \3045 , \11479 );
nor \U$17544 ( \18527 , \18525 , \18526 );
xnor \U$17545 ( \18528 , \18527 , \10427 );
and \U$17546 ( \18529 , \3508 , \10669 );
and \U$17547 ( \18530 , \3334 , \10667 );
nor \U$17548 ( \18531 , \18529 , \18530 );
xnor \U$17549 ( \18532 , \18531 , \10430 );
and \U$17550 ( \18533 , \18528 , \18532 );
and \U$17551 ( \18534 , \18532 , \2831 );
and \U$17552 ( \18535 , \18528 , \2831 );
or \U$17553 ( \18536 , \18533 , \18534 , \18535 );
and \U$17554 ( \18537 , \18523 , \18536 );
and \U$17555 ( \18538 , \18507 , \18536 );
or \U$17556 ( \18539 , \18524 , \18537 , \18538 );
and \U$17557 ( \18540 , \9365 , \4305 );
and \U$17558 ( \18541 , \9046 , \4303 );
nor \U$17559 ( \18542 , \18540 , \18541 );
xnor \U$17560 ( \18543 , \18542 , \4118 );
and \U$17561 ( \18544 , \10218 , \3992 );
and \U$17562 ( \18545 , \9649 , \3990 );
nor \U$17563 ( \18546 , \18544 , \18545 );
xnor \U$17564 ( \18547 , \18546 , \3787 );
and \U$17565 ( \18548 , \18543 , \18547 );
and \U$17566 ( \18549 , \10829 , \3586 );
and \U$17567 ( \18550 , \10226 , \3584 );
nor \U$17568 ( \18551 , \18549 , \18550 );
xnor \U$17569 ( \18552 , \18551 , \3437 );
and \U$17570 ( \18553 , \18547 , \18552 );
and \U$17571 ( \18554 , \18543 , \18552 );
or \U$17572 ( \18555 , \18548 , \18553 , \18554 );
and \U$17573 ( \18556 , \6185 , \6903 );
and \U$17574 ( \18557 , \5921 , \6901 );
nor \U$17575 ( \18558 , \18556 , \18557 );
xnor \U$17576 ( \18559 , \18558 , \6563 );
and \U$17577 ( \18560 , \6816 , \6314 );
and \U$17578 ( \18561 , \6444 , \6312 );
nor \U$17579 ( \18562 , \18560 , \18561 );
xnor \U$17580 ( \18563 , \18562 , \6073 );
and \U$17581 ( \18564 , \18559 , \18563 );
and \U$17582 ( \18565 , \7168 , \5848 );
and \U$17583 ( \18566 , \6825 , \5846 );
nor \U$17584 ( \18567 , \18565 , \18566 );
xnor \U$17585 ( \18568 , \18567 , \5660 );
and \U$17586 ( \18569 , \18563 , \18568 );
and \U$17587 ( \18570 , \18559 , \18568 );
or \U$17588 ( \18571 , \18564 , \18569 , \18570 );
and \U$17589 ( \18572 , \18555 , \18571 );
and \U$17590 ( \18573 , \7673 , \5474 );
and \U$17591 ( \18574 , \7370 , \5472 );
nor \U$17592 ( \18575 , \18573 , \18574 );
xnor \U$17593 ( \18576 , \18575 , \5242 );
and \U$17594 ( \18577 , \8371 , \5023 );
and \U$17595 ( \18578 , \7845 , \5021 );
nor \U$17596 ( \18579 , \18577 , \18578 );
xnor \U$17597 ( \18580 , \18579 , \4880 );
and \U$17598 ( \18581 , \18576 , \18580 );
and \U$17599 ( \18582 , \9041 , \4700 );
and \U$17600 ( \18583 , \8795 , \4698 );
nor \U$17601 ( \18584 , \18582 , \18583 );
xnor \U$17602 ( \18585 , \18584 , \4454 );
and \U$17603 ( \18586 , \18580 , \18585 );
and \U$17604 ( \18587 , \18576 , \18585 );
or \U$17605 ( \18588 , \18581 , \18586 , \18587 );
and \U$17606 ( \18589 , \18571 , \18588 );
and \U$17607 ( \18590 , \18555 , \18588 );
or \U$17608 ( \18591 , \18572 , \18589 , \18590 );
and \U$17609 ( \18592 , \18539 , \18591 );
and \U$17610 ( \18593 , \11635 , \2968 );
and \U$17611 ( \18594 , \11015 , \2966 );
nor \U$17612 ( \18595 , \18593 , \18594 );
xnor \U$17613 ( \18596 , \18595 , \2831 );
xor \U$17614 ( \18597 , \18310 , \18314 );
xor \U$17615 ( \18598 , \18597 , \18319 );
and \U$17616 ( \18599 , \18596 , \18598 );
xor \U$17617 ( \18600 , \18343 , \18347 );
xor \U$17618 ( \18601 , \18600 , \18352 );
and \U$17619 ( \18602 , \18598 , \18601 );
and \U$17620 ( \18603 , \18596 , \18601 );
or \U$17621 ( \18604 , \18599 , \18602 , \18603 );
and \U$17622 ( \18605 , \18591 , \18604 );
and \U$17623 ( \18606 , \18539 , \18604 );
or \U$17624 ( \18607 , \18592 , \18605 , \18606 );
xor \U$17625 ( \18608 , \18362 , \18366 );
xor \U$17626 ( \18609 , \18608 , \18371 );
xor \U$17627 ( \18610 , \18326 , \18330 );
xor \U$17628 ( \18611 , \18610 , \18335 );
and \U$17629 ( \18612 , \18609 , \18611 );
xor \U$17630 ( \18613 , \18378 , \18382 );
xor \U$17631 ( \18614 , \18613 , \18387 );
and \U$17632 ( \18615 , \18611 , \18614 );
and \U$17633 ( \18616 , \18609 , \18614 );
or \U$17634 ( \18617 , \18612 , \18615 , \18616 );
xor \U$17635 ( \18618 , \18102 , \18106 );
xor \U$17636 ( \18619 , \18618 , \2610 );
and \U$17637 ( \18620 , \18617 , \18619 );
xor \U$17638 ( \18621 , \18437 , \18439 );
xor \U$17639 ( \18622 , \18621 , \18442 );
and \U$17640 ( \18623 , \18619 , \18622 );
and \U$17641 ( \18624 , \18617 , \18622 );
or \U$17642 ( \18625 , \18620 , \18623 , \18624 );
and \U$17643 ( \18626 , \18607 , \18625 );
xor \U$17644 ( \18627 , \18322 , \18338 );
xor \U$17645 ( \18628 , \18627 , \18355 );
xor \U$17646 ( \18629 , \18374 , \18390 );
xor \U$17647 ( \18630 , \18629 , \18407 );
and \U$17648 ( \18631 , \18628 , \18630 );
xor \U$17649 ( \18632 , \18413 , \18415 );
xor \U$17650 ( \18633 , \18632 , \18418 );
and \U$17651 ( \18634 , \18630 , \18633 );
and \U$17652 ( \18635 , \18628 , \18633 );
or \U$17653 ( \18636 , \18631 , \18634 , \18635 );
and \U$17654 ( \18637 , \18625 , \18636 );
and \U$17655 ( \18638 , \18607 , \18636 );
or \U$17656 ( \18639 , \18626 , \18637 , \18638 );
xor \U$17657 ( \18640 , \18358 , \18410 );
xor \U$17658 ( \18641 , \18640 , \18421 );
xor \U$17659 ( \18642 , \18426 , \18428 );
xor \U$17660 ( \18643 , \18642 , \18431 );
and \U$17661 ( \18644 , \18641 , \18643 );
xor \U$17662 ( \18645 , \18445 , \18447 );
xor \U$17663 ( \18646 , \18645 , \18450 );
and \U$17664 ( \18647 , \18643 , \18646 );
and \U$17665 ( \18648 , \18641 , \18646 );
or \U$17666 ( \18649 , \18644 , \18647 , \18648 );
and \U$17667 ( \18650 , \18639 , \18649 );
xor \U$17668 ( \18651 , \18238 , \18248 );
xor \U$17669 ( \18652 , \18651 , \18251 );
and \U$17670 ( \18653 , \18649 , \18652 );
and \U$17671 ( \18654 , \18639 , \18652 );
or \U$17672 ( \18655 , \18650 , \18653 , \18654 );
xor \U$17673 ( \18656 , \18146 , \18172 );
xor \U$17674 ( \18657 , \18656 , \18225 );
xor \U$17675 ( \18658 , \18424 , \18434 );
xor \U$17676 ( \18659 , \18658 , \18453 );
and \U$17677 ( \18660 , \18657 , \18659 );
xor \U$17678 ( \18661 , \18458 , \18460 );
xor \U$17679 ( \18662 , \18661 , \18463 );
and \U$17680 ( \18663 , \18659 , \18662 );
and \U$17681 ( \18664 , \18657 , \18662 );
or \U$17682 ( \18665 , \18660 , \18663 , \18664 );
and \U$17683 ( \18666 , \18655 , \18665 );
xor \U$17684 ( \18667 , \18228 , \18254 );
xor \U$17685 ( \18668 , \18667 , \18265 );
and \U$17686 ( \18669 , \18665 , \18668 );
and \U$17687 ( \18670 , \18655 , \18668 );
or \U$17688 ( \18671 , \18666 , \18669 , \18670 );
xor \U$17689 ( \18672 , \18472 , \18474 );
xor \U$17690 ( \18673 , \18672 , \18476 );
and \U$17691 ( \18674 , \18671 , \18673 );
and \U$17692 ( \18675 , \18491 , \18674 );
xor \U$17693 ( \18676 , \18491 , \18674 );
xor \U$17694 ( \18677 , \18671 , \18673 );
and \U$17695 ( \18678 , \3334 , \11482 );
and \U$17696 ( \18679 , \3309 , \11479 );
nor \U$17697 ( \18680 , \18678 , \18679 );
xnor \U$17698 ( \18681 , \18680 , \10427 );
and \U$17699 ( \18682 , \3675 , \10669 );
and \U$17700 ( \18683 , \3508 , \10667 );
nor \U$17701 ( \18684 , \18682 , \18683 );
xnor \U$17702 ( \18685 , \18684 , \10430 );
and \U$17703 ( \18686 , \18681 , \18685 );
and \U$17704 ( \18687 , \3932 , \10101 );
and \U$17705 ( \18688 , \3813 , \10099 );
nor \U$17706 ( \18689 , \18687 , \18688 );
xnor \U$17707 ( \18690 , \18689 , \9791 );
and \U$17708 ( \18691 , \18685 , \18690 );
and \U$17709 ( \18692 , \18681 , \18690 );
or \U$17710 ( \18693 , \18686 , \18691 , \18692 );
and \U$17711 ( \18694 , \4557 , \9564 );
and \U$17712 ( \18695 , \4349 , \9562 );
nor \U$17713 ( \18696 , \18694 , \18695 );
xnor \U$17714 ( \18697 , \18696 , \9193 );
and \U$17715 ( \18698 , \4684 , \9002 );
and \U$17716 ( \18699 , \4679 , \9000 );
nor \U$17717 ( \18700 , \18698 , \18699 );
xnor \U$17718 ( \18701 , \18700 , \8684 );
and \U$17719 ( \18702 , \18697 , \18701 );
and \U$17720 ( \18703 , \5137 , \8435 );
and \U$17721 ( \18704 , \4940 , \8433 );
nor \U$17722 ( \18705 , \18703 , \18704 );
xnor \U$17723 ( \18706 , \18705 , \8186 );
and \U$17724 ( \18707 , \18701 , \18706 );
and \U$17725 ( \18708 , \18697 , \18706 );
or \U$17726 ( \18709 , \18702 , \18707 , \18708 );
and \U$17727 ( \18710 , \18693 , \18709 );
and \U$17728 ( \18711 , \5447 , \7906 );
and \U$17729 ( \18712 , \5439 , \7904 );
nor \U$17730 ( \18713 , \18711 , \18712 );
xnor \U$17731 ( \18714 , \18713 , \7646 );
and \U$17732 ( \18715 , \5921 , \7412 );
and \U$17733 ( \18716 , \5916 , \7410 );
nor \U$17734 ( \18717 , \18715 , \18716 );
xnor \U$17735 ( \18718 , \18717 , \7097 );
and \U$17736 ( \18719 , \18714 , \18718 );
and \U$17737 ( \18720 , \6444 , \6903 );
and \U$17738 ( \18721 , \6185 , \6901 );
nor \U$17739 ( \18722 , \18720 , \18721 );
xnor \U$17740 ( \18723 , \18722 , \6563 );
and \U$17741 ( \18724 , \18718 , \18723 );
and \U$17742 ( \18725 , \18714 , \18723 );
or \U$17743 ( \18726 , \18719 , \18724 , \18725 );
and \U$17744 ( \18727 , \18709 , \18726 );
and \U$17745 ( \18728 , \18693 , \18726 );
or \U$17746 ( \18729 , \18710 , \18727 , \18728 );
and \U$17747 ( \18730 , \10226 , \3992 );
and \U$17748 ( \18731 , \10218 , \3990 );
nor \U$17749 ( \18732 , \18730 , \18731 );
xnor \U$17750 ( \18733 , \18732 , \3787 );
and \U$17751 ( \18734 , \10834 , \3586 );
and \U$17752 ( \18735 , \10829 , \3584 );
nor \U$17753 ( \18736 , \18734 , \18735 );
xnor \U$17754 ( \18737 , \18736 , \3437 );
and \U$17755 ( \18738 , \18733 , \18737 );
and \U$17756 ( \18739 , \11635 , \3264 );
and \U$17757 ( \18740 , \11015 , \3262 );
nor \U$17758 ( \18741 , \18739 , \18740 );
xnor \U$17759 ( \18742 , \18741 , \3122 );
and \U$17760 ( \18743 , \18737 , \18742 );
and \U$17761 ( \18744 , \18733 , \18742 );
or \U$17762 ( \18745 , \18738 , \18743 , \18744 );
and \U$17763 ( \18746 , \8795 , \5023 );
and \U$17764 ( \18747 , \8371 , \5021 );
nor \U$17765 ( \18748 , \18746 , \18747 );
xnor \U$17766 ( \18749 , \18748 , \4880 );
and \U$17767 ( \18750 , \9046 , \4700 );
and \U$17768 ( \18751 , \9041 , \4698 );
nor \U$17769 ( \18752 , \18750 , \18751 );
xnor \U$17770 ( \18753 , \18752 , \4454 );
and \U$17771 ( \18754 , \18749 , \18753 );
and \U$17772 ( \18755 , \9649 , \4305 );
and \U$17773 ( \18756 , \9365 , \4303 );
nor \U$17774 ( \18757 , \18755 , \18756 );
xnor \U$17775 ( \18758 , \18757 , \4118 );
and \U$17776 ( \18759 , \18753 , \18758 );
and \U$17777 ( \18760 , \18749 , \18758 );
or \U$17778 ( \18761 , \18754 , \18759 , \18760 );
and \U$17779 ( \18762 , \18745 , \18761 );
and \U$17780 ( \18763 , \6825 , \6314 );
and \U$17781 ( \18764 , \6816 , \6312 );
nor \U$17782 ( \18765 , \18763 , \18764 );
xnor \U$17783 ( \18766 , \18765 , \6073 );
and \U$17784 ( \18767 , \7370 , \5848 );
and \U$17785 ( \18768 , \7168 , \5846 );
nor \U$17786 ( \18769 , \18767 , \18768 );
xnor \U$17787 ( \18770 , \18769 , \5660 );
and \U$17788 ( \18771 , \18766 , \18770 );
and \U$17789 ( \18772 , \7845 , \5474 );
and \U$17790 ( \18773 , \7673 , \5472 );
nor \U$17791 ( \18774 , \18772 , \18773 );
xnor \U$17792 ( \18775 , \18774 , \5242 );
and \U$17793 ( \18776 , \18770 , \18775 );
and \U$17794 ( \18777 , \18766 , \18775 );
or \U$17795 ( \18778 , \18771 , \18776 , \18777 );
and \U$17796 ( \18779 , \18761 , \18778 );
and \U$17797 ( \18780 , \18745 , \18778 );
or \U$17798 ( \18781 , \18762 , \18779 , \18780 );
and \U$17799 ( \18782 , \18729 , \18781 );
and \U$17800 ( \18783 , \11015 , \3264 );
and \U$17801 ( \18784 , \10834 , \3262 );
nor \U$17802 ( \18785 , \18783 , \18784 );
xnor \U$17803 ( \18786 , \18785 , \3122 );
nand \U$17804 ( \18787 , \11635 , \2966 );
xnor \U$17805 ( \18788 , \18787 , \2831 );
and \U$17806 ( \18789 , \18786 , \18788 );
xor \U$17807 ( \18790 , \18543 , \18547 );
xor \U$17808 ( \18791 , \18790 , \18552 );
and \U$17809 ( \18792 , \18788 , \18791 );
and \U$17810 ( \18793 , \18786 , \18791 );
or \U$17811 ( \18794 , \18789 , \18792 , \18793 );
and \U$17812 ( \18795 , \18781 , \18794 );
and \U$17813 ( \18796 , \18729 , \18794 );
or \U$17814 ( \18797 , \18782 , \18795 , \18796 );
xor \U$17815 ( \18798 , \18495 , \18499 );
xor \U$17816 ( \18799 , \18798 , \18504 );
xor \U$17817 ( \18800 , \18559 , \18563 );
xor \U$17818 ( \18801 , \18800 , \18568 );
and \U$17819 ( \18802 , \18799 , \18801 );
xor \U$17820 ( \18803 , \18576 , \18580 );
xor \U$17821 ( \18804 , \18803 , \18585 );
and \U$17822 ( \18805 , \18801 , \18804 );
and \U$17823 ( \18806 , \18799 , \18804 );
or \U$17824 ( \18807 , \18802 , \18805 , \18806 );
xor \U$17825 ( \18808 , \18511 , \18515 );
xor \U$17826 ( \18809 , \18808 , \18520 );
xor \U$17827 ( \18810 , \18528 , \18532 );
xor \U$17828 ( \18811 , \18810 , \2831 );
and \U$17829 ( \18812 , \18809 , \18811 );
and \U$17830 ( \18813 , \18807 , \18812 );
xor \U$17831 ( \18814 , \18395 , \18399 );
xor \U$17832 ( \18815 , \18814 , \18404 );
and \U$17833 ( \18816 , \18812 , \18815 );
and \U$17834 ( \18817 , \18807 , \18815 );
or \U$17835 ( \18818 , \18813 , \18816 , \18817 );
and \U$17836 ( \18819 , \18797 , \18818 );
xor \U$17837 ( \18820 , \18555 , \18571 );
xor \U$17838 ( \18821 , \18820 , \18588 );
xor \U$17839 ( \18822 , \18609 , \18611 );
xor \U$17840 ( \18823 , \18822 , \18614 );
and \U$17841 ( \18824 , \18821 , \18823 );
xor \U$17842 ( \18825 , \18596 , \18598 );
xor \U$17843 ( \18826 , \18825 , \18601 );
and \U$17844 ( \18827 , \18823 , \18826 );
and \U$17845 ( \18828 , \18821 , \18826 );
or \U$17846 ( \18829 , \18824 , \18827 , \18828 );
and \U$17847 ( \18830 , \18818 , \18829 );
and \U$17848 ( \18831 , \18797 , \18829 );
or \U$17849 ( \18832 , \18819 , \18830 , \18831 );
xor \U$17850 ( \18833 , \18539 , \18591 );
xor \U$17851 ( \18834 , \18833 , \18604 );
xor \U$17852 ( \18835 , \18617 , \18619 );
xor \U$17853 ( \18836 , \18835 , \18622 );
and \U$17854 ( \18837 , \18834 , \18836 );
xor \U$17855 ( \18838 , \18628 , \18630 );
xor \U$17856 ( \18839 , \18838 , \18633 );
and \U$17857 ( \18840 , \18836 , \18839 );
and \U$17858 ( \18841 , \18834 , \18839 );
or \U$17859 ( \18842 , \18837 , \18840 , \18841 );
and \U$17860 ( \18843 , \18832 , \18842 );
xor \U$17861 ( \18844 , \18641 , \18643 );
xor \U$17862 ( \18845 , \18844 , \18646 );
and \U$17863 ( \18846 , \18842 , \18845 );
and \U$17864 ( \18847 , \18832 , \18845 );
or \U$17865 ( \18848 , \18843 , \18846 , \18847 );
xor \U$17866 ( \18849 , \18639 , \18649 );
xor \U$17867 ( \18850 , \18849 , \18652 );
and \U$17868 ( \18851 , \18848 , \18850 );
xor \U$17869 ( \18852 , \18657 , \18659 );
xor \U$17870 ( \18853 , \18852 , \18662 );
and \U$17871 ( \18854 , \18850 , \18853 );
and \U$17872 ( \18855 , \18848 , \18853 );
or \U$17873 ( \18856 , \18851 , \18854 , \18855 );
xor \U$17874 ( \18857 , \18655 , \18665 );
xor \U$17875 ( \18858 , \18857 , \18668 );
and \U$17876 ( \18859 , \18856 , \18858 );
xor \U$17877 ( \18860 , \18456 , \18466 );
xor \U$17878 ( \18861 , \18860 , \18469 );
and \U$17879 ( \18862 , \18858 , \18861 );
and \U$17880 ( \18863 , \18856 , \18861 );
or \U$17881 ( \18864 , \18859 , \18862 , \18863 );
and \U$17882 ( \18865 , \18677 , \18864 );
xor \U$17883 ( \18866 , \18677 , \18864 );
xor \U$17884 ( \18867 , \18856 , \18858 );
xor \U$17885 ( \18868 , \18867 , \18861 );
and \U$17886 ( \18869 , \3508 , \11482 );
and \U$17887 ( \18870 , \3334 , \11479 );
nor \U$17888 ( \18871 , \18869 , \18870 );
xnor \U$17889 ( \18872 , \18871 , \10427 );
and \U$17890 ( \18873 , \3813 , \10669 );
and \U$17891 ( \18874 , \3675 , \10667 );
nor \U$17892 ( \18875 , \18873 , \18874 );
xnor \U$17893 ( \18876 , \18875 , \10430 );
and \U$17894 ( \18877 , \18872 , \18876 );
and \U$17895 ( \18878 , \18876 , \3122 );
and \U$17896 ( \18879 , \18872 , \3122 );
or \U$17897 ( \18880 , \18877 , \18878 , \18879 );
and \U$17898 ( \18881 , \4349 , \10101 );
and \U$17899 ( \18882 , \3932 , \10099 );
nor \U$17900 ( \18883 , \18881 , \18882 );
xnor \U$17901 ( \18884 , \18883 , \9791 );
and \U$17902 ( \18885 , \4679 , \9564 );
and \U$17903 ( \18886 , \4557 , \9562 );
nor \U$17904 ( \18887 , \18885 , \18886 );
xnor \U$17905 ( \18888 , \18887 , \9193 );
and \U$17906 ( \18889 , \18884 , \18888 );
and \U$17907 ( \18890 , \4940 , \9002 );
and \U$17908 ( \18891 , \4684 , \9000 );
nor \U$17909 ( \18892 , \18890 , \18891 );
xnor \U$17910 ( \18893 , \18892 , \8684 );
and \U$17911 ( \18894 , \18888 , \18893 );
and \U$17912 ( \18895 , \18884 , \18893 );
or \U$17913 ( \18896 , \18889 , \18894 , \18895 );
and \U$17914 ( \18897 , \18880 , \18896 );
and \U$17915 ( \18898 , \5439 , \8435 );
and \U$17916 ( \18899 , \5137 , \8433 );
nor \U$17917 ( \18900 , \18898 , \18899 );
xnor \U$17918 ( \18901 , \18900 , \8186 );
and \U$17919 ( \18902 , \5916 , \7906 );
and \U$17920 ( \18903 , \5447 , \7904 );
nor \U$17921 ( \18904 , \18902 , \18903 );
xnor \U$17922 ( \18905 , \18904 , \7646 );
and \U$17923 ( \18906 , \18901 , \18905 );
and \U$17924 ( \18907 , \6185 , \7412 );
and \U$17925 ( \18908 , \5921 , \7410 );
nor \U$17926 ( \18909 , \18907 , \18908 );
xnor \U$17927 ( \18910 , \18909 , \7097 );
and \U$17928 ( \18911 , \18905 , \18910 );
and \U$17929 ( \18912 , \18901 , \18910 );
or \U$17930 ( \18913 , \18906 , \18911 , \18912 );
and \U$17931 ( \18914 , \18896 , \18913 );
and \U$17932 ( \18915 , \18880 , \18913 );
or \U$17933 ( \18916 , \18897 , \18914 , \18915 );
and \U$17934 ( \18917 , \6816 , \6903 );
and \U$17935 ( \18918 , \6444 , \6901 );
nor \U$17936 ( \18919 , \18917 , \18918 );
xnor \U$17937 ( \18920 , \18919 , \6563 );
and \U$17938 ( \18921 , \7168 , \6314 );
and \U$17939 ( \18922 , \6825 , \6312 );
nor \U$17940 ( \18923 , \18921 , \18922 );
xnor \U$17941 ( \18924 , \18923 , \6073 );
and \U$17942 ( \18925 , \18920 , \18924 );
and \U$17943 ( \18926 , \7673 , \5848 );
and \U$17944 ( \18927 , \7370 , \5846 );
nor \U$17945 ( \18928 , \18926 , \18927 );
xnor \U$17946 ( \18929 , \18928 , \5660 );
and \U$17947 ( \18930 , \18924 , \18929 );
and \U$17948 ( \18931 , \18920 , \18929 );
or \U$17949 ( \18932 , \18925 , \18930 , \18931 );
and \U$17950 ( \18933 , \8371 , \5474 );
and \U$17951 ( \18934 , \7845 , \5472 );
nor \U$17952 ( \18935 , \18933 , \18934 );
xnor \U$17953 ( \18936 , \18935 , \5242 );
and \U$17954 ( \18937 , \9041 , \5023 );
and \U$17955 ( \18938 , \8795 , \5021 );
nor \U$17956 ( \18939 , \18937 , \18938 );
xnor \U$17957 ( \18940 , \18939 , \4880 );
and \U$17958 ( \18941 , \18936 , \18940 );
and \U$17959 ( \18942 , \9365 , \4700 );
and \U$17960 ( \18943 , \9046 , \4698 );
nor \U$17961 ( \18944 , \18942 , \18943 );
xnor \U$17962 ( \18945 , \18944 , \4454 );
and \U$17963 ( \18946 , \18940 , \18945 );
and \U$17964 ( \18947 , \18936 , \18945 );
or \U$17965 ( \18948 , \18941 , \18946 , \18947 );
and \U$17966 ( \18949 , \18932 , \18948 );
and \U$17967 ( \18950 , \10218 , \4305 );
and \U$17968 ( \18951 , \9649 , \4303 );
nor \U$17969 ( \18952 , \18950 , \18951 );
xnor \U$17970 ( \18953 , \18952 , \4118 );
and \U$17971 ( \18954 , \10829 , \3992 );
and \U$17972 ( \18955 , \10226 , \3990 );
nor \U$17973 ( \18956 , \18954 , \18955 );
xnor \U$17974 ( \18957 , \18956 , \3787 );
and \U$17975 ( \18958 , \18953 , \18957 );
and \U$17976 ( \18959 , \11015 , \3586 );
and \U$17977 ( \18960 , \10834 , \3584 );
nor \U$17978 ( \18961 , \18959 , \18960 );
xnor \U$17979 ( \18962 , \18961 , \3437 );
and \U$17980 ( \18963 , \18957 , \18962 );
and \U$17981 ( \18964 , \18953 , \18962 );
or \U$17982 ( \18965 , \18958 , \18963 , \18964 );
and \U$17983 ( \18966 , \18948 , \18965 );
and \U$17984 ( \18967 , \18932 , \18965 );
or \U$17985 ( \18968 , \18949 , \18966 , \18967 );
and \U$17986 ( \18969 , \18916 , \18968 );
xor \U$17987 ( \18970 , \18733 , \18737 );
xor \U$17988 ( \18971 , \18970 , \18742 );
xor \U$17989 ( \18972 , \18749 , \18753 );
xor \U$17990 ( \18973 , \18972 , \18758 );
and \U$17991 ( \18974 , \18971 , \18973 );
xor \U$17992 ( \18975 , \18766 , \18770 );
xor \U$17993 ( \18976 , \18975 , \18775 );
and \U$17994 ( \18977 , \18973 , \18976 );
and \U$17995 ( \18978 , \18971 , \18976 );
or \U$17996 ( \18979 , \18974 , \18977 , \18978 );
and \U$17997 ( \18980 , \18968 , \18979 );
and \U$17998 ( \18981 , \18916 , \18979 );
or \U$17999 ( \18982 , \18969 , \18980 , \18981 );
xor \U$18000 ( \18983 , \18693 , \18709 );
xor \U$18001 ( \18984 , \18983 , \18726 );
xor \U$18002 ( \18985 , \18745 , \18761 );
xor \U$18003 ( \18986 , \18985 , \18778 );
and \U$18004 ( \18987 , \18984 , \18986 );
xor \U$18005 ( \18988 , \18786 , \18788 );
xor \U$18006 ( \18989 , \18988 , \18791 );
and \U$18007 ( \18990 , \18986 , \18989 );
and \U$18008 ( \18991 , \18984 , \18989 );
or \U$18009 ( \18992 , \18987 , \18990 , \18991 );
and \U$18010 ( \18993 , \18982 , \18992 );
xor \U$18011 ( \18994 , \18681 , \18685 );
xor \U$18012 ( \18995 , \18994 , \18690 );
xor \U$18013 ( \18996 , \18697 , \18701 );
xor \U$18014 ( \18997 , \18996 , \18706 );
and \U$18015 ( \18998 , \18995 , \18997 );
xor \U$18016 ( \18999 , \18714 , \18718 );
xor \U$18017 ( \19000 , \18999 , \18723 );
and \U$18018 ( \19001 , \18997 , \19000 );
and \U$18019 ( \19002 , \18995 , \19000 );
or \U$18020 ( \19003 , \18998 , \19001 , \19002 );
xor \U$18021 ( \19004 , \18799 , \18801 );
xor \U$18022 ( \19005 , \19004 , \18804 );
and \U$18023 ( \19006 , \19003 , \19005 );
xor \U$18024 ( \19007 , \18809 , \18811 );
and \U$18025 ( \19008 , \19005 , \19007 );
and \U$18026 ( \19009 , \19003 , \19007 );
or \U$18027 ( \19010 , \19006 , \19008 , \19009 );
and \U$18028 ( \19011 , \18992 , \19010 );
and \U$18029 ( \19012 , \18982 , \19010 );
or \U$18030 ( \19013 , \18993 , \19011 , \19012 );
xor \U$18031 ( \19014 , \18507 , \18523 );
xor \U$18032 ( \19015 , \19014 , \18536 );
xor \U$18033 ( \19016 , \18807 , \18812 );
xor \U$18034 ( \19017 , \19016 , \18815 );
and \U$18035 ( \19018 , \19015 , \19017 );
xor \U$18036 ( \19019 , \18821 , \18823 );
xor \U$18037 ( \19020 , \19019 , \18826 );
and \U$18038 ( \19021 , \19017 , \19020 );
and \U$18039 ( \19022 , \19015 , \19020 );
or \U$18040 ( \19023 , \19018 , \19021 , \19022 );
and \U$18041 ( \19024 , \19013 , \19023 );
xor \U$18042 ( \19025 , \18834 , \18836 );
xor \U$18043 ( \19026 , \19025 , \18839 );
and \U$18044 ( \19027 , \19023 , \19026 );
and \U$18045 ( \19028 , \19013 , \19026 );
or \U$18046 ( \19029 , \19024 , \19027 , \19028 );
xor \U$18047 ( \19030 , \18607 , \18625 );
xor \U$18048 ( \19031 , \19030 , \18636 );
and \U$18049 ( \19032 , \19029 , \19031 );
xor \U$18050 ( \19033 , \18832 , \18842 );
xor \U$18051 ( \19034 , \19033 , \18845 );
and \U$18052 ( \19035 , \19031 , \19034 );
and \U$18053 ( \19036 , \19029 , \19034 );
or \U$18054 ( \19037 , \19032 , \19035 , \19036 );
xor \U$18055 ( \19038 , \18848 , \18850 );
xor \U$18056 ( \19039 , \19038 , \18853 );
and \U$18057 ( \19040 , \19037 , \19039 );
and \U$18058 ( \19041 , \18868 , \19040 );
xor \U$18059 ( \19042 , \18868 , \19040 );
xor \U$18060 ( \19043 , \19037 , \19039 );
and \U$18061 ( \19044 , \5921 , \7906 );
and \U$18062 ( \19045 , \5916 , \7904 );
nor \U$18063 ( \19046 , \19044 , \19045 );
xnor \U$18064 ( \19047 , \19046 , \7646 );
and \U$18065 ( \19048 , \6444 , \7412 );
and \U$18066 ( \19049 , \6185 , \7410 );
nor \U$18067 ( \19050 , \19048 , \19049 );
xnor \U$18068 ( \19051 , \19050 , \7097 );
and \U$18069 ( \19052 , \19047 , \19051 );
and \U$18070 ( \19053 , \6825 , \6903 );
and \U$18071 ( \19054 , \6816 , \6901 );
nor \U$18072 ( \19055 , \19053 , \19054 );
xnor \U$18073 ( \19056 , \19055 , \6563 );
and \U$18074 ( \19057 , \19051 , \19056 );
and \U$18075 ( \19058 , \19047 , \19056 );
or \U$18076 ( \19059 , \19052 , \19057 , \19058 );
and \U$18077 ( \19060 , \3675 , \11482 );
and \U$18078 ( \19061 , \3508 , \11479 );
nor \U$18079 ( \19062 , \19060 , \19061 );
xnor \U$18080 ( \19063 , \19062 , \10427 );
and \U$18081 ( \19064 , \3932 , \10669 );
and \U$18082 ( \19065 , \3813 , \10667 );
nor \U$18083 ( \19066 , \19064 , \19065 );
xnor \U$18084 ( \19067 , \19066 , \10430 );
and \U$18085 ( \19068 , \19063 , \19067 );
and \U$18086 ( \19069 , \4557 , \10101 );
and \U$18087 ( \19070 , \4349 , \10099 );
nor \U$18088 ( \19071 , \19069 , \19070 );
xnor \U$18089 ( \19072 , \19071 , \9791 );
and \U$18090 ( \19073 , \19067 , \19072 );
and \U$18091 ( \19074 , \19063 , \19072 );
or \U$18092 ( \19075 , \19068 , \19073 , \19074 );
and \U$18093 ( \19076 , \19059 , \19075 );
and \U$18094 ( \19077 , \4684 , \9564 );
and \U$18095 ( \19078 , \4679 , \9562 );
nor \U$18096 ( \19079 , \19077 , \19078 );
xnor \U$18097 ( \19080 , \19079 , \9193 );
and \U$18098 ( \19081 , \5137 , \9002 );
and \U$18099 ( \19082 , \4940 , \9000 );
nor \U$18100 ( \19083 , \19081 , \19082 );
xnor \U$18101 ( \19084 , \19083 , \8684 );
and \U$18102 ( \19085 , \19080 , \19084 );
and \U$18103 ( \19086 , \5447 , \8435 );
and \U$18104 ( \19087 , \5439 , \8433 );
nor \U$18105 ( \19088 , \19086 , \19087 );
xnor \U$18106 ( \19089 , \19088 , \8186 );
and \U$18107 ( \19090 , \19084 , \19089 );
and \U$18108 ( \19091 , \19080 , \19089 );
or \U$18109 ( \19092 , \19085 , \19090 , \19091 );
and \U$18110 ( \19093 , \19075 , \19092 );
and \U$18111 ( \19094 , \19059 , \19092 );
or \U$18112 ( \19095 , \19076 , \19093 , \19094 );
and \U$18113 ( \19096 , \9046 , \5023 );
and \U$18114 ( \19097 , \9041 , \5021 );
nor \U$18115 ( \19098 , \19096 , \19097 );
xnor \U$18116 ( \19099 , \19098 , \4880 );
and \U$18117 ( \19100 , \9649 , \4700 );
and \U$18118 ( \19101 , \9365 , \4698 );
nor \U$18119 ( \19102 , \19100 , \19101 );
xnor \U$18120 ( \19103 , \19102 , \4454 );
and \U$18121 ( \19104 , \19099 , \19103 );
and \U$18122 ( \19105 , \10226 , \4305 );
and \U$18123 ( \19106 , \10218 , \4303 );
nor \U$18124 ( \19107 , \19105 , \19106 );
xnor \U$18125 ( \19108 , \19107 , \4118 );
and \U$18126 ( \19109 , \19103 , \19108 );
and \U$18127 ( \19110 , \19099 , \19108 );
or \U$18128 ( \19111 , \19104 , \19109 , \19110 );
and \U$18129 ( \19112 , \7370 , \6314 );
and \U$18130 ( \19113 , \7168 , \6312 );
nor \U$18131 ( \19114 , \19112 , \19113 );
xnor \U$18132 ( \19115 , \19114 , \6073 );
and \U$18133 ( \19116 , \7845 , \5848 );
and \U$18134 ( \19117 , \7673 , \5846 );
nor \U$18135 ( \19118 , \19116 , \19117 );
xnor \U$18136 ( \19119 , \19118 , \5660 );
and \U$18137 ( \19120 , \19115 , \19119 );
and \U$18138 ( \19121 , \8795 , \5474 );
and \U$18139 ( \19122 , \8371 , \5472 );
nor \U$18140 ( \19123 , \19121 , \19122 );
xnor \U$18141 ( \19124 , \19123 , \5242 );
and \U$18142 ( \19125 , \19119 , \19124 );
and \U$18143 ( \19126 , \19115 , \19124 );
or \U$18144 ( \19127 , \19120 , \19125 , \19126 );
and \U$18145 ( \19128 , \19111 , \19127 );
and \U$18146 ( \19129 , \10834 , \3992 );
and \U$18147 ( \19130 , \10829 , \3990 );
nor \U$18148 ( \19131 , \19129 , \19130 );
xnor \U$18149 ( \19132 , \19131 , \3787 );
and \U$18150 ( \19133 , \11635 , \3586 );
and \U$18151 ( \19134 , \11015 , \3584 );
nor \U$18152 ( \19135 , \19133 , \19134 );
xnor \U$18153 ( \19136 , \19135 , \3437 );
and \U$18154 ( \19137 , \19132 , \19136 );
and \U$18155 ( \19138 , \19127 , \19137 );
and \U$18156 ( \19139 , \19111 , \19137 );
or \U$18157 ( \19140 , \19128 , \19138 , \19139 );
and \U$18158 ( \19141 , \19095 , \19140 );
nand \U$18159 ( \19142 , \11635 , \3262 );
xnor \U$18160 ( \19143 , \19142 , \3122 );
xor \U$18161 ( \19144 , \18936 , \18940 );
xor \U$18162 ( \19145 , \19144 , \18945 );
and \U$18163 ( \19146 , \19143 , \19145 );
xor \U$18164 ( \19147 , \18953 , \18957 );
xor \U$18165 ( \19148 , \19147 , \18962 );
and \U$18166 ( \19149 , \19145 , \19148 );
and \U$18167 ( \19150 , \19143 , \19148 );
or \U$18168 ( \19151 , \19146 , \19149 , \19150 );
and \U$18169 ( \19152 , \19140 , \19151 );
and \U$18170 ( \19153 , \19095 , \19151 );
or \U$18171 ( \19154 , \19141 , \19152 , \19153 );
xor \U$18172 ( \19155 , \18884 , \18888 );
xor \U$18173 ( \19156 , \19155 , \18893 );
xor \U$18174 ( \19157 , \18920 , \18924 );
xor \U$18175 ( \19158 , \19157 , \18929 );
and \U$18176 ( \19159 , \19156 , \19158 );
xor \U$18177 ( \19160 , \18901 , \18905 );
xor \U$18178 ( \19161 , \19160 , \18910 );
and \U$18179 ( \19162 , \19158 , \19161 );
and \U$18180 ( \19163 , \19156 , \19161 );
or \U$18181 ( \19164 , \19159 , \19162 , \19163 );
xor \U$18182 ( \19165 , \18971 , \18973 );
xor \U$18183 ( \19166 , \19165 , \18976 );
and \U$18184 ( \19167 , \19164 , \19166 );
xor \U$18185 ( \19168 , \18995 , \18997 );
xor \U$18186 ( \19169 , \19168 , \19000 );
and \U$18187 ( \19170 , \19166 , \19169 );
and \U$18188 ( \19171 , \19164 , \19169 );
or \U$18189 ( \19172 , \19167 , \19170 , \19171 );
and \U$18190 ( \19173 , \19154 , \19172 );
xor \U$18191 ( \19174 , \18880 , \18896 );
xor \U$18192 ( \19175 , \19174 , \18913 );
xor \U$18193 ( \19176 , \18932 , \18948 );
xor \U$18194 ( \19177 , \19176 , \18965 );
and \U$18195 ( \19178 , \19175 , \19177 );
and \U$18196 ( \19179 , \19172 , \19178 );
and \U$18197 ( \19180 , \19154 , \19178 );
or \U$18198 ( \19181 , \19173 , \19179 , \19180 );
xor \U$18199 ( \19182 , \18916 , \18968 );
xor \U$18200 ( \19183 , \19182 , \18979 );
xor \U$18201 ( \19184 , \18984 , \18986 );
xor \U$18202 ( \19185 , \19184 , \18989 );
and \U$18203 ( \19186 , \19183 , \19185 );
xor \U$18204 ( \19187 , \19003 , \19005 );
xor \U$18205 ( \19188 , \19187 , \19007 );
and \U$18206 ( \19189 , \19185 , \19188 );
and \U$18207 ( \19190 , \19183 , \19188 );
or \U$18208 ( \19191 , \19186 , \19189 , \19190 );
and \U$18209 ( \19192 , \19181 , \19191 );
xor \U$18210 ( \19193 , \18729 , \18781 );
xor \U$18211 ( \19194 , \19193 , \18794 );
and \U$18212 ( \19195 , \19191 , \19194 );
and \U$18213 ( \19196 , \19181 , \19194 );
or \U$18214 ( \19197 , \19192 , \19195 , \19196 );
xor \U$18215 ( \19198 , \18982 , \18992 );
xor \U$18216 ( \19199 , \19198 , \19010 );
xor \U$18217 ( \19200 , \19015 , \19017 );
xor \U$18218 ( \19201 , \19200 , \19020 );
and \U$18219 ( \19202 , \19199 , \19201 );
and \U$18220 ( \19203 , \19197 , \19202 );
xor \U$18221 ( \19204 , \18797 , \18818 );
xor \U$18222 ( \19205 , \19204 , \18829 );
and \U$18223 ( \19206 , \19202 , \19205 );
and \U$18224 ( \19207 , \19197 , \19205 );
or \U$18225 ( \19208 , \19203 , \19206 , \19207 );
xor \U$18226 ( \19209 , \19029 , \19031 );
xor \U$18227 ( \19210 , \19209 , \19034 );
and \U$18228 ( \19211 , \19208 , \19210 );
and \U$18229 ( \19212 , \19043 , \19211 );
xor \U$18230 ( \19213 , \19043 , \19211 );
xor \U$18231 ( \19214 , \19208 , \19210 );
xor \U$18232 ( \19215 , \19197 , \19202 );
xor \U$18233 ( \19216 , \19215 , \19205 );
xor \U$18234 ( \19217 , \19013 , \19023 );
xor \U$18235 ( \19218 , \19217 , \19026 );
and \U$18236 ( \19219 , \19216 , \19218 );
and \U$18237 ( \19220 , \19214 , \19219 );
xor \U$18238 ( \19221 , \19214 , \19219 );
xor \U$18239 ( \19222 , \19216 , \19218 );
and \U$18240 ( \19223 , \9041 , \5474 );
and \U$18241 ( \19224 , \8795 , \5472 );
nor \U$18242 ( \19225 , \19223 , \19224 );
xnor \U$18243 ( \19226 , \19225 , \5242 );
and \U$18244 ( \19227 , \9365 , \5023 );
and \U$18245 ( \19228 , \9046 , \5021 );
nor \U$18246 ( \19229 , \19227 , \19228 );
xnor \U$18247 ( \19230 , \19229 , \4880 );
and \U$18248 ( \19231 , \19226 , \19230 );
and \U$18249 ( \19232 , \10218 , \4700 );
and \U$18250 ( \19233 , \9649 , \4698 );
nor \U$18251 ( \19234 , \19232 , \19233 );
xnor \U$18252 ( \19235 , \19234 , \4454 );
and \U$18253 ( \19236 , \19230 , \19235 );
and \U$18254 ( \19237 , \19226 , \19235 );
or \U$18255 ( \19238 , \19231 , \19236 , \19237 );
and \U$18256 ( \19239 , \10829 , \4305 );
and \U$18257 ( \19240 , \10226 , \4303 );
nor \U$18258 ( \19241 , \19239 , \19240 );
xnor \U$18259 ( \19242 , \19241 , \4118 );
and \U$18260 ( \19243 , \11015 , \3992 );
and \U$18261 ( \19244 , \10834 , \3990 );
nor \U$18262 ( \19245 , \19243 , \19244 );
xnor \U$18263 ( \19246 , \19245 , \3787 );
and \U$18264 ( \19247 , \19242 , \19246 );
nand \U$18265 ( \19248 , \11635 , \3584 );
xnor \U$18266 ( \19249 , \19248 , \3437 );
and \U$18267 ( \19250 , \19246 , \19249 );
and \U$18268 ( \19251 , \19242 , \19249 );
or \U$18269 ( \19252 , \19247 , \19250 , \19251 );
and \U$18270 ( \19253 , \19238 , \19252 );
and \U$18271 ( \19254 , \7168 , \6903 );
and \U$18272 ( \19255 , \6825 , \6901 );
nor \U$18273 ( \19256 , \19254 , \19255 );
xnor \U$18274 ( \19257 , \19256 , \6563 );
and \U$18275 ( \19258 , \7673 , \6314 );
and \U$18276 ( \19259 , \7370 , \6312 );
nor \U$18277 ( \19260 , \19258 , \19259 );
xnor \U$18278 ( \19261 , \19260 , \6073 );
and \U$18279 ( \19262 , \19257 , \19261 );
and \U$18280 ( \19263 , \8371 , \5848 );
and \U$18281 ( \19264 , \7845 , \5846 );
nor \U$18282 ( \19265 , \19263 , \19264 );
xnor \U$18283 ( \19266 , \19265 , \5660 );
and \U$18284 ( \19267 , \19261 , \19266 );
and \U$18285 ( \19268 , \19257 , \19266 );
or \U$18286 ( \19269 , \19262 , \19267 , \19268 );
and \U$18287 ( \19270 , \19252 , \19269 );
and \U$18288 ( \19271 , \19238 , \19269 );
or \U$18289 ( \19272 , \19253 , \19270 , \19271 );
and \U$18290 ( \19273 , \5916 , \8435 );
and \U$18291 ( \19274 , \5447 , \8433 );
nor \U$18292 ( \19275 , \19273 , \19274 );
xnor \U$18293 ( \19276 , \19275 , \8186 );
and \U$18294 ( \19277 , \6185 , \7906 );
and \U$18295 ( \19278 , \5921 , \7904 );
nor \U$18296 ( \19279 , \19277 , \19278 );
xnor \U$18297 ( \19280 , \19279 , \7646 );
and \U$18298 ( \19281 , \19276 , \19280 );
and \U$18299 ( \19282 , \6816 , \7412 );
and \U$18300 ( \19283 , \6444 , \7410 );
nor \U$18301 ( \19284 , \19282 , \19283 );
xnor \U$18302 ( \19285 , \19284 , \7097 );
and \U$18303 ( \19286 , \19280 , \19285 );
and \U$18304 ( \19287 , \19276 , \19285 );
or \U$18305 ( \19288 , \19281 , \19286 , \19287 );
and \U$18306 ( \19289 , \3813 , \11482 );
and \U$18307 ( \19290 , \3675 , \11479 );
nor \U$18308 ( \19291 , \19289 , \19290 );
xnor \U$18309 ( \19292 , \19291 , \10427 );
and \U$18310 ( \19293 , \4349 , \10669 );
and \U$18311 ( \19294 , \3932 , \10667 );
nor \U$18312 ( \19295 , \19293 , \19294 );
xnor \U$18313 ( \19296 , \19295 , \10430 );
and \U$18314 ( \19297 , \19292 , \19296 );
and \U$18315 ( \19298 , \19296 , \3437 );
and \U$18316 ( \19299 , \19292 , \3437 );
or \U$18317 ( \19300 , \19297 , \19298 , \19299 );
and \U$18318 ( \19301 , \19288 , \19300 );
and \U$18319 ( \19302 , \4679 , \10101 );
and \U$18320 ( \19303 , \4557 , \10099 );
nor \U$18321 ( \19304 , \19302 , \19303 );
xnor \U$18322 ( \19305 , \19304 , \9791 );
and \U$18323 ( \19306 , \4940 , \9564 );
and \U$18324 ( \19307 , \4684 , \9562 );
nor \U$18325 ( \19308 , \19306 , \19307 );
xnor \U$18326 ( \19309 , \19308 , \9193 );
and \U$18327 ( \19310 , \19305 , \19309 );
and \U$18328 ( \19311 , \5439 , \9002 );
and \U$18329 ( \19312 , \5137 , \9000 );
nor \U$18330 ( \19313 , \19311 , \19312 );
xnor \U$18331 ( \19314 , \19313 , \8684 );
and \U$18332 ( \19315 , \19309 , \19314 );
and \U$18333 ( \19316 , \19305 , \19314 );
or \U$18334 ( \19317 , \19310 , \19315 , \19316 );
and \U$18335 ( \19318 , \19300 , \19317 );
and \U$18336 ( \19319 , \19288 , \19317 );
or \U$18337 ( \19320 , \19301 , \19318 , \19319 );
and \U$18338 ( \19321 , \19272 , \19320 );
xor \U$18339 ( \19322 , \19099 , \19103 );
xor \U$18340 ( \19323 , \19322 , \19108 );
xor \U$18341 ( \19324 , \19115 , \19119 );
xor \U$18342 ( \19325 , \19324 , \19124 );
and \U$18343 ( \19326 , \19323 , \19325 );
xor \U$18344 ( \19327 , \19132 , \19136 );
and \U$18345 ( \19328 , \19325 , \19327 );
and \U$18346 ( \19329 , \19323 , \19327 );
or \U$18347 ( \19330 , \19326 , \19328 , \19329 );
and \U$18348 ( \19331 , \19320 , \19330 );
and \U$18349 ( \19332 , \19272 , \19330 );
or \U$18350 ( \19333 , \19321 , \19331 , \19332 );
xor \U$18351 ( \19334 , \19047 , \19051 );
xor \U$18352 ( \19335 , \19334 , \19056 );
xor \U$18353 ( \19336 , \19063 , \19067 );
xor \U$18354 ( \19337 , \19336 , \19072 );
and \U$18355 ( \19338 , \19335 , \19337 );
xor \U$18356 ( \19339 , \19080 , \19084 );
xor \U$18357 ( \19340 , \19339 , \19089 );
and \U$18358 ( \19341 , \19337 , \19340 );
and \U$18359 ( \19342 , \19335 , \19340 );
or \U$18360 ( \19343 , \19338 , \19341 , \19342 );
xor \U$18361 ( \19344 , \18872 , \18876 );
xor \U$18362 ( \19345 , \19344 , \3122 );
and \U$18363 ( \19346 , \19343 , \19345 );
xor \U$18364 ( \19347 , \19156 , \19158 );
xor \U$18365 ( \19348 , \19347 , \19161 );
and \U$18366 ( \19349 , \19345 , \19348 );
and \U$18367 ( \19350 , \19343 , \19348 );
or \U$18368 ( \19351 , \19346 , \19349 , \19350 );
and \U$18369 ( \19352 , \19333 , \19351 );
xor \U$18370 ( \19353 , \19059 , \19075 );
xor \U$18371 ( \19354 , \19353 , \19092 );
xor \U$18372 ( \19355 , \19111 , \19127 );
xor \U$18373 ( \19356 , \19355 , \19137 );
and \U$18374 ( \19357 , \19354 , \19356 );
xor \U$18375 ( \19358 , \19143 , \19145 );
xor \U$18376 ( \19359 , \19358 , \19148 );
and \U$18377 ( \19360 , \19356 , \19359 );
and \U$18378 ( \19361 , \19354 , \19359 );
or \U$18379 ( \19362 , \19357 , \19360 , \19361 );
and \U$18380 ( \19363 , \19351 , \19362 );
and \U$18381 ( \19364 , \19333 , \19362 );
or \U$18382 ( \19365 , \19352 , \19363 , \19364 );
xor \U$18383 ( \19366 , \19095 , \19140 );
xor \U$18384 ( \19367 , \19366 , \19151 );
xor \U$18385 ( \19368 , \19164 , \19166 );
xor \U$18386 ( \19369 , \19368 , \19169 );
and \U$18387 ( \19370 , \19367 , \19369 );
xor \U$18388 ( \19371 , \19175 , \19177 );
and \U$18389 ( \19372 , \19369 , \19371 );
and \U$18390 ( \19373 , \19367 , \19371 );
or \U$18391 ( \19374 , \19370 , \19372 , \19373 );
and \U$18392 ( \19375 , \19365 , \19374 );
xor \U$18393 ( \19376 , \19183 , \19185 );
xor \U$18394 ( \19377 , \19376 , \19188 );
and \U$18395 ( \19378 , \19374 , \19377 );
and \U$18396 ( \19379 , \19365 , \19377 );
or \U$18397 ( \19380 , \19375 , \19378 , \19379 );
xor \U$18398 ( \19381 , \19181 , \19191 );
xor \U$18399 ( \19382 , \19381 , \19194 );
and \U$18400 ( \19383 , \19380 , \19382 );
xor \U$18401 ( \19384 , \19199 , \19201 );
and \U$18402 ( \19385 , \19382 , \19384 );
and \U$18403 ( \19386 , \19380 , \19384 );
or \U$18404 ( \19387 , \19383 , \19385 , \19386 );
and \U$18405 ( \19388 , \19222 , \19387 );
xor \U$18406 ( \19389 , \19222 , \19387 );
xor \U$18407 ( \19390 , \19380 , \19382 );
xor \U$18408 ( \19391 , \19390 , \19384 );
and \U$18409 ( \19392 , \5137 , \9564 );
and \U$18410 ( \19393 , \4940 , \9562 );
nor \U$18411 ( \19394 , \19392 , \19393 );
xnor \U$18412 ( \19395 , \19394 , \9193 );
and \U$18413 ( \19396 , \5447 , \9002 );
and \U$18414 ( \19397 , \5439 , \9000 );
nor \U$18415 ( \19398 , \19396 , \19397 );
xnor \U$18416 ( \19399 , \19398 , \8684 );
and \U$18417 ( \19400 , \19395 , \19399 );
and \U$18418 ( \19401 , \5921 , \8435 );
and \U$18419 ( \19402 , \5916 , \8433 );
nor \U$18420 ( \19403 , \19401 , \19402 );
xnor \U$18421 ( \19404 , \19403 , \8186 );
and \U$18422 ( \19405 , \19399 , \19404 );
and \U$18423 ( \19406 , \19395 , \19404 );
or \U$18424 ( \19407 , \19400 , \19405 , \19406 );
and \U$18425 ( \19408 , \3932 , \11482 );
and \U$18426 ( \19409 , \3813 , \11479 );
nor \U$18427 ( \19410 , \19408 , \19409 );
xnor \U$18428 ( \19411 , \19410 , \10427 );
and \U$18429 ( \19412 , \4557 , \10669 );
and \U$18430 ( \19413 , \4349 , \10667 );
nor \U$18431 ( \19414 , \19412 , \19413 );
xnor \U$18432 ( \19415 , \19414 , \10430 );
and \U$18433 ( \19416 , \19411 , \19415 );
and \U$18434 ( \19417 , \4684 , \10101 );
and \U$18435 ( \19418 , \4679 , \10099 );
nor \U$18436 ( \19419 , \19417 , \19418 );
xnor \U$18437 ( \19420 , \19419 , \9791 );
and \U$18438 ( \19421 , \19415 , \19420 );
and \U$18439 ( \19422 , \19411 , \19420 );
or \U$18440 ( \19423 , \19416 , \19421 , \19422 );
and \U$18441 ( \19424 , \19407 , \19423 );
and \U$18442 ( \19425 , \6444 , \7906 );
and \U$18443 ( \19426 , \6185 , \7904 );
nor \U$18444 ( \19427 , \19425 , \19426 );
xnor \U$18445 ( \19428 , \19427 , \7646 );
and \U$18446 ( \19429 , \6825 , \7412 );
and \U$18447 ( \19430 , \6816 , \7410 );
nor \U$18448 ( \19431 , \19429 , \19430 );
xnor \U$18449 ( \19432 , \19431 , \7097 );
and \U$18450 ( \19433 , \19428 , \19432 );
and \U$18451 ( \19434 , \7370 , \6903 );
and \U$18452 ( \19435 , \7168 , \6901 );
nor \U$18453 ( \19436 , \19434 , \19435 );
xnor \U$18454 ( \19437 , \19436 , \6563 );
and \U$18455 ( \19438 , \19432 , \19437 );
and \U$18456 ( \19439 , \19428 , \19437 );
or \U$18457 ( \19440 , \19433 , \19438 , \19439 );
and \U$18458 ( \19441 , \19423 , \19440 );
and \U$18459 ( \19442 , \19407 , \19440 );
or \U$18460 ( \19443 , \19424 , \19441 , \19442 );
xor \U$18461 ( \19444 , \19226 , \19230 );
xor \U$18462 ( \19445 , \19444 , \19235 );
xor \U$18463 ( \19446 , \19276 , \19280 );
xor \U$18464 ( \19447 , \19446 , \19285 );
and \U$18465 ( \19448 , \19445 , \19447 );
xor \U$18466 ( \19449 , \19257 , \19261 );
xor \U$18467 ( \19450 , \19449 , \19266 );
and \U$18468 ( \19451 , \19447 , \19450 );
and \U$18469 ( \19452 , \19445 , \19450 );
or \U$18470 ( \19453 , \19448 , \19451 , \19452 );
and \U$18471 ( \19454 , \19443 , \19453 );
and \U$18472 ( \19455 , \7845 , \6314 );
and \U$18473 ( \19456 , \7673 , \6312 );
nor \U$18474 ( \19457 , \19455 , \19456 );
xnor \U$18475 ( \19458 , \19457 , \6073 );
and \U$18476 ( \19459 , \8795 , \5848 );
and \U$18477 ( \19460 , \8371 , \5846 );
nor \U$18478 ( \19461 , \19459 , \19460 );
xnor \U$18479 ( \19462 , \19461 , \5660 );
and \U$18480 ( \19463 , \19458 , \19462 );
and \U$18481 ( \19464 , \9046 , \5474 );
and \U$18482 ( \19465 , \9041 , \5472 );
nor \U$18483 ( \19466 , \19464 , \19465 );
xnor \U$18484 ( \19467 , \19466 , \5242 );
and \U$18485 ( \19468 , \19462 , \19467 );
and \U$18486 ( \19469 , \19458 , \19467 );
or \U$18487 ( \19470 , \19463 , \19468 , \19469 );
and \U$18488 ( \19471 , \9649 , \5023 );
and \U$18489 ( \19472 , \9365 , \5021 );
nor \U$18490 ( \19473 , \19471 , \19472 );
xnor \U$18491 ( \19474 , \19473 , \4880 );
and \U$18492 ( \19475 , \10226 , \4700 );
and \U$18493 ( \19476 , \10218 , \4698 );
nor \U$18494 ( \19477 , \19475 , \19476 );
xnor \U$18495 ( \19478 , \19477 , \4454 );
and \U$18496 ( \19479 , \19474 , \19478 );
and \U$18497 ( \19480 , \10834 , \4305 );
and \U$18498 ( \19481 , \10829 , \4303 );
nor \U$18499 ( \19482 , \19480 , \19481 );
xnor \U$18500 ( \19483 , \19482 , \4118 );
and \U$18501 ( \19484 , \19478 , \19483 );
and \U$18502 ( \19485 , \19474 , \19483 );
or \U$18503 ( \19486 , \19479 , \19484 , \19485 );
and \U$18504 ( \19487 , \19470 , \19486 );
xor \U$18505 ( \19488 , \19242 , \19246 );
xor \U$18506 ( \19489 , \19488 , \19249 );
and \U$18507 ( \19490 , \19486 , \19489 );
and \U$18508 ( \19491 , \19470 , \19489 );
or \U$18509 ( \19492 , \19487 , \19490 , \19491 );
and \U$18510 ( \19493 , \19453 , \19492 );
and \U$18511 ( \19494 , \19443 , \19492 );
or \U$18512 ( \19495 , \19454 , \19493 , \19494 );
xor \U$18513 ( \19496 , \19238 , \19252 );
xor \U$18514 ( \19497 , \19496 , \19269 );
xor \U$18515 ( \19498 , \19335 , \19337 );
xor \U$18516 ( \19499 , \19498 , \19340 );
and \U$18517 ( \19500 , \19497 , \19499 );
xor \U$18518 ( \19501 , \19323 , \19325 );
xor \U$18519 ( \19502 , \19501 , \19327 );
and \U$18520 ( \19503 , \19499 , \19502 );
and \U$18521 ( \19504 , \19497 , \19502 );
or \U$18522 ( \19505 , \19500 , \19503 , \19504 );
and \U$18523 ( \19506 , \19495 , \19505 );
xor \U$18524 ( \19507 , \19354 , \19356 );
xor \U$18525 ( \19508 , \19507 , \19359 );
and \U$18526 ( \19509 , \19505 , \19508 );
and \U$18527 ( \19510 , \19495 , \19508 );
or \U$18528 ( \19511 , \19506 , \19509 , \19510 );
xor \U$18529 ( \19512 , \19333 , \19351 );
xor \U$18530 ( \19513 , \19512 , \19362 );
and \U$18531 ( \19514 , \19511 , \19513 );
xor \U$18532 ( \19515 , \19367 , \19369 );
xor \U$18533 ( \19516 , \19515 , \19371 );
and \U$18534 ( \19517 , \19513 , \19516 );
and \U$18535 ( \19518 , \19511 , \19516 );
or \U$18536 ( \19519 , \19514 , \19517 , \19518 );
xor \U$18537 ( \19520 , \19154 , \19172 );
xor \U$18538 ( \19521 , \19520 , \19178 );
and \U$18539 ( \19522 , \19519 , \19521 );
xor \U$18540 ( \19523 , \19365 , \19374 );
xor \U$18541 ( \19524 , \19523 , \19377 );
and \U$18542 ( \19525 , \19521 , \19524 );
and \U$18543 ( \19526 , \19519 , \19524 );
or \U$18544 ( \19527 , \19522 , \19525 , \19526 );
and \U$18545 ( \19528 , \19391 , \19527 );
xor \U$18546 ( \19529 , \19391 , \19527 );
xor \U$18547 ( \19530 , \19519 , \19521 );
xor \U$18548 ( \19531 , \19530 , \19524 );
and \U$18549 ( \19532 , \4940 , \10101 );
and \U$18550 ( \19533 , \4684 , \10099 );
nor \U$18551 ( \19534 , \19532 , \19533 );
xnor \U$18552 ( \19535 , \19534 , \9791 );
and \U$18553 ( \19536 , \5439 , \9564 );
and \U$18554 ( \19537 , \5137 , \9562 );
nor \U$18555 ( \19538 , \19536 , \19537 );
xnor \U$18556 ( \19539 , \19538 , \9193 );
and \U$18557 ( \19540 , \19535 , \19539 );
and \U$18558 ( \19541 , \5916 , \9002 );
and \U$18559 ( \19542 , \5447 , \9000 );
nor \U$18560 ( \19543 , \19541 , \19542 );
xnor \U$18561 ( \19544 , \19543 , \8684 );
and \U$18562 ( \19545 , \19539 , \19544 );
and \U$18563 ( \19546 , \19535 , \19544 );
or \U$18564 ( \19547 , \19540 , \19545 , \19546 );
and \U$18565 ( \19548 , \6185 , \8435 );
and \U$18566 ( \19549 , \5921 , \8433 );
nor \U$18567 ( \19550 , \19548 , \19549 );
xnor \U$18568 ( \19551 , \19550 , \8186 );
and \U$18569 ( \19552 , \6816 , \7906 );
and \U$18570 ( \19553 , \6444 , \7904 );
nor \U$18571 ( \19554 , \19552 , \19553 );
xnor \U$18572 ( \19555 , \19554 , \7646 );
and \U$18573 ( \19556 , \19551 , \19555 );
and \U$18574 ( \19557 , \7168 , \7412 );
and \U$18575 ( \19558 , \6825 , \7410 );
nor \U$18576 ( \19559 , \19557 , \19558 );
xnor \U$18577 ( \19560 , \19559 , \7097 );
and \U$18578 ( \19561 , \19555 , \19560 );
and \U$18579 ( \19562 , \19551 , \19560 );
or \U$18580 ( \19563 , \19556 , \19561 , \19562 );
and \U$18581 ( \19564 , \19547 , \19563 );
and \U$18582 ( \19565 , \4349 , \11482 );
and \U$18583 ( \19566 , \3932 , \11479 );
nor \U$18584 ( \19567 , \19565 , \19566 );
xnor \U$18585 ( \19568 , \19567 , \10427 );
and \U$18586 ( \19569 , \4679 , \10669 );
and \U$18587 ( \19570 , \4557 , \10667 );
nor \U$18588 ( \19571 , \19569 , \19570 );
xnor \U$18589 ( \19572 , \19571 , \10430 );
and \U$18590 ( \19573 , \19568 , \19572 );
and \U$18591 ( \19574 , \19572 , \3787 );
and \U$18592 ( \19575 , \19568 , \3787 );
or \U$18593 ( \19576 , \19573 , \19574 , \19575 );
and \U$18594 ( \19577 , \19563 , \19576 );
and \U$18595 ( \19578 , \19547 , \19576 );
or \U$18596 ( \19579 , \19564 , \19577 , \19578 );
and \U$18597 ( \19580 , \9365 , \5474 );
and \U$18598 ( \19581 , \9046 , \5472 );
nor \U$18599 ( \19582 , \19580 , \19581 );
xnor \U$18600 ( \19583 , \19582 , \5242 );
and \U$18601 ( \19584 , \10218 , \5023 );
and \U$18602 ( \19585 , \9649 , \5021 );
nor \U$18603 ( \19586 , \19584 , \19585 );
xnor \U$18604 ( \19587 , \19586 , \4880 );
and \U$18605 ( \19588 , \19583 , \19587 );
and \U$18606 ( \19589 , \10829 , \4700 );
and \U$18607 ( \19590 , \10226 , \4698 );
nor \U$18608 ( \19591 , \19589 , \19590 );
xnor \U$18609 ( \19592 , \19591 , \4454 );
and \U$18610 ( \19593 , \19587 , \19592 );
and \U$18611 ( \19594 , \19583 , \19592 );
or \U$18612 ( \19595 , \19588 , \19593 , \19594 );
and \U$18613 ( \19596 , \7673 , \6903 );
and \U$18614 ( \19597 , \7370 , \6901 );
nor \U$18615 ( \19598 , \19596 , \19597 );
xnor \U$18616 ( \19599 , \19598 , \6563 );
and \U$18617 ( \19600 , \8371 , \6314 );
and \U$18618 ( \19601 , \7845 , \6312 );
nor \U$18619 ( \19602 , \19600 , \19601 );
xnor \U$18620 ( \19603 , \19602 , \6073 );
and \U$18621 ( \19604 , \19599 , \19603 );
and \U$18622 ( \19605 , \9041 , \5848 );
and \U$18623 ( \19606 , \8795 , \5846 );
nor \U$18624 ( \19607 , \19605 , \19606 );
xnor \U$18625 ( \19608 , \19607 , \5660 );
and \U$18626 ( \19609 , \19603 , \19608 );
and \U$18627 ( \19610 , \19599 , \19608 );
or \U$18628 ( \19611 , \19604 , \19609 , \19610 );
and \U$18629 ( \19612 , \19595 , \19611 );
and \U$18630 ( \19613 , \11635 , \3992 );
and \U$18631 ( \19614 , \11015 , \3990 );
nor \U$18632 ( \19615 , \19613 , \19614 );
xnor \U$18633 ( \19616 , \19615 , \3787 );
and \U$18634 ( \19617 , \19611 , \19616 );
and \U$18635 ( \19618 , \19595 , \19616 );
or \U$18636 ( \19619 , \19612 , \19617 , \19618 );
and \U$18637 ( \19620 , \19579 , \19619 );
xor \U$18638 ( \19621 , \19458 , \19462 );
xor \U$18639 ( \19622 , \19621 , \19467 );
xor \U$18640 ( \19623 , \19474 , \19478 );
xor \U$18641 ( \19624 , \19623 , \19483 );
and \U$18642 ( \19625 , \19622 , \19624 );
xor \U$18643 ( \19626 , \19428 , \19432 );
xor \U$18644 ( \19627 , \19626 , \19437 );
and \U$18645 ( \19628 , \19624 , \19627 );
and \U$18646 ( \19629 , \19622 , \19627 );
or \U$18647 ( \19630 , \19625 , \19628 , \19629 );
and \U$18648 ( \19631 , \19619 , \19630 );
and \U$18649 ( \19632 , \19579 , \19630 );
or \U$18650 ( \19633 , \19620 , \19631 , \19632 );
xor \U$18651 ( \19634 , \19292 , \19296 );
xor \U$18652 ( \19635 , \19634 , \3437 );
xor \U$18653 ( \19636 , \19305 , \19309 );
xor \U$18654 ( \19637 , \19636 , \19314 );
and \U$18655 ( \19638 , \19635 , \19637 );
xor \U$18656 ( \19639 , \19445 , \19447 );
xor \U$18657 ( \19640 , \19639 , \19450 );
and \U$18658 ( \19641 , \19637 , \19640 );
and \U$18659 ( \19642 , \19635 , \19640 );
or \U$18660 ( \19643 , \19638 , \19641 , \19642 );
and \U$18661 ( \19644 , \19633 , \19643 );
xor \U$18662 ( \19645 , \19407 , \19423 );
xor \U$18663 ( \19646 , \19645 , \19440 );
xor \U$18664 ( \19647 , \19470 , \19486 );
xor \U$18665 ( \19648 , \19647 , \19489 );
and \U$18666 ( \19649 , \19646 , \19648 );
and \U$18667 ( \19650 , \19643 , \19649 );
and \U$18668 ( \19651 , \19633 , \19649 );
or \U$18669 ( \19652 , \19644 , \19650 , \19651 );
xor \U$18670 ( \19653 , \19288 , \19300 );
xor \U$18671 ( \19654 , \19653 , \19317 );
xor \U$18672 ( \19655 , \19443 , \19453 );
xor \U$18673 ( \19656 , \19655 , \19492 );
and \U$18674 ( \19657 , \19654 , \19656 );
xor \U$18675 ( \19658 , \19497 , \19499 );
xor \U$18676 ( \19659 , \19658 , \19502 );
and \U$18677 ( \19660 , \19656 , \19659 );
and \U$18678 ( \19661 , \19654 , \19659 );
or \U$18679 ( \19662 , \19657 , \19660 , \19661 );
and \U$18680 ( \19663 , \19652 , \19662 );
xor \U$18681 ( \19664 , \19343 , \19345 );
xor \U$18682 ( \19665 , \19664 , \19348 );
and \U$18683 ( \19666 , \19662 , \19665 );
and \U$18684 ( \19667 , \19652 , \19665 );
or \U$18685 ( \19668 , \19663 , \19666 , \19667 );
xor \U$18686 ( \19669 , \19272 , \19320 );
xor \U$18687 ( \19670 , \19669 , \19330 );
xor \U$18688 ( \19671 , \19495 , \19505 );
xor \U$18689 ( \19672 , \19671 , \19508 );
and \U$18690 ( \19673 , \19670 , \19672 );
and \U$18691 ( \19674 , \19668 , \19673 );
xor \U$18692 ( \19675 , \19511 , \19513 );
xor \U$18693 ( \19676 , \19675 , \19516 );
and \U$18694 ( \19677 , \19673 , \19676 );
and \U$18695 ( \19678 , \19668 , \19676 );
or \U$18696 ( \19679 , \19674 , \19677 , \19678 );
and \U$18697 ( \19680 , \19531 , \19679 );
xor \U$18698 ( \19681 , \19531 , \19679 );
xor \U$18699 ( \19682 , \19668 , \19673 );
xor \U$18700 ( \19683 , \19682 , \19676 );
and \U$18701 ( \19684 , \6825 , \7906 );
and \U$18702 ( \19685 , \6816 , \7904 );
nor \U$18703 ( \19686 , \19684 , \19685 );
xnor \U$18704 ( \19687 , \19686 , \7646 );
and \U$18705 ( \19688 , \7370 , \7412 );
and \U$18706 ( \19689 , \7168 , \7410 );
nor \U$18707 ( \19690 , \19688 , \19689 );
xnor \U$18708 ( \19691 , \19690 , \7097 );
and \U$18709 ( \19692 , \19687 , \19691 );
and \U$18710 ( \19693 , \7845 , \6903 );
and \U$18711 ( \19694 , \7673 , \6901 );
nor \U$18712 ( \19695 , \19693 , \19694 );
xnor \U$18713 ( \19696 , \19695 , \6563 );
and \U$18714 ( \19697 , \19691 , \19696 );
and \U$18715 ( \19698 , \19687 , \19696 );
or \U$18716 ( \19699 , \19692 , \19697 , \19698 );
and \U$18717 ( \19700 , \5447 , \9564 );
and \U$18718 ( \19701 , \5439 , \9562 );
nor \U$18719 ( \19702 , \19700 , \19701 );
xnor \U$18720 ( \19703 , \19702 , \9193 );
and \U$18721 ( \19704 , \5921 , \9002 );
and \U$18722 ( \19705 , \5916 , \9000 );
nor \U$18723 ( \19706 , \19704 , \19705 );
xnor \U$18724 ( \19707 , \19706 , \8684 );
and \U$18725 ( \19708 , \19703 , \19707 );
and \U$18726 ( \19709 , \6444 , \8435 );
and \U$18727 ( \19710 , \6185 , \8433 );
nor \U$18728 ( \19711 , \19709 , \19710 );
xnor \U$18729 ( \19712 , \19711 , \8186 );
and \U$18730 ( \19713 , \19707 , \19712 );
and \U$18731 ( \19714 , \19703 , \19712 );
or \U$18732 ( \19715 , \19708 , \19713 , \19714 );
and \U$18733 ( \19716 , \19699 , \19715 );
and \U$18734 ( \19717 , \4557 , \11482 );
and \U$18735 ( \19718 , \4349 , \11479 );
nor \U$18736 ( \19719 , \19717 , \19718 );
xnor \U$18737 ( \19720 , \19719 , \10427 );
and \U$18738 ( \19721 , \4684 , \10669 );
and \U$18739 ( \19722 , \4679 , \10667 );
nor \U$18740 ( \19723 , \19721 , \19722 );
xnor \U$18741 ( \19724 , \19723 , \10430 );
and \U$18742 ( \19725 , \19720 , \19724 );
and \U$18743 ( \19726 , \5137 , \10101 );
and \U$18744 ( \19727 , \4940 , \10099 );
nor \U$18745 ( \19728 , \19726 , \19727 );
xnor \U$18746 ( \19729 , \19728 , \9791 );
and \U$18747 ( \19730 , \19724 , \19729 );
and \U$18748 ( \19731 , \19720 , \19729 );
or \U$18749 ( \19732 , \19725 , \19730 , \19731 );
and \U$18750 ( \19733 , \19715 , \19732 );
and \U$18751 ( \19734 , \19699 , \19732 );
or \U$18752 ( \19735 , \19716 , \19733 , \19734 );
and \U$18753 ( \19736 , \10226 , \5023 );
and \U$18754 ( \19737 , \10218 , \5021 );
nor \U$18755 ( \19738 , \19736 , \19737 );
xnor \U$18756 ( \19739 , \19738 , \4880 );
and \U$18757 ( \19740 , \10834 , \4700 );
and \U$18758 ( \19741 , \10829 , \4698 );
nor \U$18759 ( \19742 , \19740 , \19741 );
xnor \U$18760 ( \19743 , \19742 , \4454 );
and \U$18761 ( \19744 , \19739 , \19743 );
and \U$18762 ( \19745 , \11635 , \4305 );
and \U$18763 ( \19746 , \11015 , \4303 );
nor \U$18764 ( \19747 , \19745 , \19746 );
xnor \U$18765 ( \19748 , \19747 , \4118 );
and \U$18766 ( \19749 , \19743 , \19748 );
and \U$18767 ( \19750 , \19739 , \19748 );
or \U$18768 ( \19751 , \19744 , \19749 , \19750 );
and \U$18769 ( \19752 , \8795 , \6314 );
and \U$18770 ( \19753 , \8371 , \6312 );
nor \U$18771 ( \19754 , \19752 , \19753 );
xnor \U$18772 ( \19755 , \19754 , \6073 );
and \U$18773 ( \19756 , \9046 , \5848 );
and \U$18774 ( \19757 , \9041 , \5846 );
nor \U$18775 ( \19758 , \19756 , \19757 );
xnor \U$18776 ( \19759 , \19758 , \5660 );
and \U$18777 ( \19760 , \19755 , \19759 );
and \U$18778 ( \19761 , \9649 , \5474 );
and \U$18779 ( \19762 , \9365 , \5472 );
nor \U$18780 ( \19763 , \19761 , \19762 );
xnor \U$18781 ( \19764 , \19763 , \5242 );
and \U$18782 ( \19765 , \19759 , \19764 );
and \U$18783 ( \19766 , \19755 , \19764 );
or \U$18784 ( \19767 , \19760 , \19765 , \19766 );
and \U$18785 ( \19768 , \19751 , \19767 );
and \U$18786 ( \19769 , \11015 , \4305 );
and \U$18787 ( \19770 , \10834 , \4303 );
nor \U$18788 ( \19771 , \19769 , \19770 );
xnor \U$18789 ( \19772 , \19771 , \4118 );
and \U$18790 ( \19773 , \19767 , \19772 );
and \U$18791 ( \19774 , \19751 , \19772 );
or \U$18792 ( \19775 , \19768 , \19773 , \19774 );
and \U$18793 ( \19776 , \19735 , \19775 );
nand \U$18794 ( \19777 , \11635 , \3990 );
xnor \U$18795 ( \19778 , \19777 , \3787 );
xor \U$18796 ( \19779 , \19583 , \19587 );
xor \U$18797 ( \19780 , \19779 , \19592 );
and \U$18798 ( \19781 , \19778 , \19780 );
xor \U$18799 ( \19782 , \19599 , \19603 );
xor \U$18800 ( \19783 , \19782 , \19608 );
and \U$18801 ( \19784 , \19780 , \19783 );
and \U$18802 ( \19785 , \19778 , \19783 );
or \U$18803 ( \19786 , \19781 , \19784 , \19785 );
and \U$18804 ( \19787 , \19775 , \19786 );
and \U$18805 ( \19788 , \19735 , \19786 );
or \U$18806 ( \19789 , \19776 , \19787 , \19788 );
xor \U$18807 ( \19790 , \19535 , \19539 );
xor \U$18808 ( \19791 , \19790 , \19544 );
xor \U$18809 ( \19792 , \19551 , \19555 );
xor \U$18810 ( \19793 , \19792 , \19560 );
and \U$18811 ( \19794 , \19791 , \19793 );
xor \U$18812 ( \19795 , \19568 , \19572 );
xor \U$18813 ( \19796 , \19795 , \3787 );
and \U$18814 ( \19797 , \19793 , \19796 );
and \U$18815 ( \19798 , \19791 , \19796 );
or \U$18816 ( \19799 , \19794 , \19797 , \19798 );
xor \U$18817 ( \19800 , \19395 , \19399 );
xor \U$18818 ( \19801 , \19800 , \19404 );
and \U$18819 ( \19802 , \19799 , \19801 );
xor \U$18820 ( \19803 , \19411 , \19415 );
xor \U$18821 ( \19804 , \19803 , \19420 );
and \U$18822 ( \19805 , \19801 , \19804 );
and \U$18823 ( \19806 , \19799 , \19804 );
or \U$18824 ( \19807 , \19802 , \19805 , \19806 );
and \U$18825 ( \19808 , \19789 , \19807 );
xor \U$18826 ( \19809 , \19547 , \19563 );
xor \U$18827 ( \19810 , \19809 , \19576 );
xor \U$18828 ( \19811 , \19595 , \19611 );
xor \U$18829 ( \19812 , \19811 , \19616 );
and \U$18830 ( \19813 , \19810 , \19812 );
xor \U$18831 ( \19814 , \19622 , \19624 );
xor \U$18832 ( \19815 , \19814 , \19627 );
and \U$18833 ( \19816 , \19812 , \19815 );
and \U$18834 ( \19817 , \19810 , \19815 );
or \U$18835 ( \19818 , \19813 , \19816 , \19817 );
and \U$18836 ( \19819 , \19807 , \19818 );
and \U$18837 ( \19820 , \19789 , \19818 );
or \U$18838 ( \19821 , \19808 , \19819 , \19820 );
xor \U$18839 ( \19822 , \19579 , \19619 );
xor \U$18840 ( \19823 , \19822 , \19630 );
xor \U$18841 ( \19824 , \19635 , \19637 );
xor \U$18842 ( \19825 , \19824 , \19640 );
and \U$18843 ( \19826 , \19823 , \19825 );
xor \U$18844 ( \19827 , \19646 , \19648 );
and \U$18845 ( \19828 , \19825 , \19827 );
and \U$18846 ( \19829 , \19823 , \19827 );
or \U$18847 ( \19830 , \19826 , \19828 , \19829 );
and \U$18848 ( \19831 , \19821 , \19830 );
xor \U$18849 ( \19832 , \19654 , \19656 );
xor \U$18850 ( \19833 , \19832 , \19659 );
and \U$18851 ( \19834 , \19830 , \19833 );
and \U$18852 ( \19835 , \19821 , \19833 );
or \U$18853 ( \19836 , \19831 , \19834 , \19835 );
xor \U$18854 ( \19837 , \19652 , \19662 );
xor \U$18855 ( \19838 , \19837 , \19665 );
and \U$18856 ( \19839 , \19836 , \19838 );
xor \U$18857 ( \19840 , \19670 , \19672 );
and \U$18858 ( \19841 , \19838 , \19840 );
and \U$18859 ( \19842 , \19836 , \19840 );
or \U$18860 ( \19843 , \19839 , \19841 , \19842 );
and \U$18861 ( \19844 , \19683 , \19843 );
xor \U$18862 ( \19845 , \19683 , \19843 );
xor \U$18863 ( \19846 , \19836 , \19838 );
xor \U$18864 ( \19847 , \19846 , \19840 );
and \U$18865 ( \19848 , \6816 , \8435 );
and \U$18866 ( \19849 , \6444 , \8433 );
nor \U$18867 ( \19850 , \19848 , \19849 );
xnor \U$18868 ( \19851 , \19850 , \8186 );
and \U$18869 ( \19852 , \7168 , \7906 );
and \U$18870 ( \19853 , \6825 , \7904 );
nor \U$18871 ( \19854 , \19852 , \19853 );
xnor \U$18872 ( \19855 , \19854 , \7646 );
and \U$18873 ( \19856 , \19851 , \19855 );
and \U$18874 ( \19857 , \7673 , \7412 );
and \U$18875 ( \19858 , \7370 , \7410 );
nor \U$18876 ( \19859 , \19857 , \19858 );
xnor \U$18877 ( \19860 , \19859 , \7097 );
and \U$18878 ( \19861 , \19855 , \19860 );
and \U$18879 ( \19862 , \19851 , \19860 );
or \U$18880 ( \19863 , \19856 , \19861 , \19862 );
and \U$18881 ( \19864 , \5439 , \10101 );
and \U$18882 ( \19865 , \5137 , \10099 );
nor \U$18883 ( \19866 , \19864 , \19865 );
xnor \U$18884 ( \19867 , \19866 , \9791 );
and \U$18885 ( \19868 , \5916 , \9564 );
and \U$18886 ( \19869 , \5447 , \9562 );
nor \U$18887 ( \19870 , \19868 , \19869 );
xnor \U$18888 ( \19871 , \19870 , \9193 );
and \U$18889 ( \19872 , \19867 , \19871 );
and \U$18890 ( \19873 , \6185 , \9002 );
and \U$18891 ( \19874 , \5921 , \9000 );
nor \U$18892 ( \19875 , \19873 , \19874 );
xnor \U$18893 ( \19876 , \19875 , \8684 );
and \U$18894 ( \19877 , \19871 , \19876 );
and \U$18895 ( \19878 , \19867 , \19876 );
or \U$18896 ( \19879 , \19872 , \19877 , \19878 );
and \U$18897 ( \19880 , \19863 , \19879 );
and \U$18898 ( \19881 , \4679 , \11482 );
and \U$18899 ( \19882 , \4557 , \11479 );
nor \U$18900 ( \19883 , \19881 , \19882 );
xnor \U$18901 ( \19884 , \19883 , \10427 );
and \U$18902 ( \19885 , \4940 , \10669 );
and \U$18903 ( \19886 , \4684 , \10667 );
nor \U$18904 ( \19887 , \19885 , \19886 );
xnor \U$18905 ( \19888 , \19887 , \10430 );
and \U$18906 ( \19889 , \19884 , \19888 );
and \U$18907 ( \19890 , \19888 , \4118 );
and \U$18908 ( \19891 , \19884 , \4118 );
or \U$18909 ( \19892 , \19889 , \19890 , \19891 );
and \U$18910 ( \19893 , \19879 , \19892 );
and \U$18911 ( \19894 , \19863 , \19892 );
or \U$18912 ( \19895 , \19880 , \19893 , \19894 );
and \U$18913 ( \19896 , \8371 , \6903 );
and \U$18914 ( \19897 , \7845 , \6901 );
nor \U$18915 ( \19898 , \19896 , \19897 );
xnor \U$18916 ( \19899 , \19898 , \6563 );
and \U$18917 ( \19900 , \9041 , \6314 );
and \U$18918 ( \19901 , \8795 , \6312 );
nor \U$18919 ( \19902 , \19900 , \19901 );
xnor \U$18920 ( \19903 , \19902 , \6073 );
and \U$18921 ( \19904 , \19899 , \19903 );
and \U$18922 ( \19905 , \9365 , \5848 );
and \U$18923 ( \19906 , \9046 , \5846 );
nor \U$18924 ( \19907 , \19905 , \19906 );
xnor \U$18925 ( \19908 , \19907 , \5660 );
and \U$18926 ( \19909 , \19903 , \19908 );
and \U$18927 ( \19910 , \19899 , \19908 );
or \U$18928 ( \19911 , \19904 , \19909 , \19910 );
and \U$18929 ( \19912 , \10218 , \5474 );
and \U$18930 ( \19913 , \9649 , \5472 );
nor \U$18931 ( \19914 , \19912 , \19913 );
xnor \U$18932 ( \19915 , \19914 , \5242 );
and \U$18933 ( \19916 , \10829 , \5023 );
and \U$18934 ( \19917 , \10226 , \5021 );
nor \U$18935 ( \19918 , \19916 , \19917 );
xnor \U$18936 ( \19919 , \19918 , \4880 );
and \U$18937 ( \19920 , \19915 , \19919 );
and \U$18938 ( \19921 , \11015 , \4700 );
and \U$18939 ( \19922 , \10834 , \4698 );
nor \U$18940 ( \19923 , \19921 , \19922 );
xnor \U$18941 ( \19924 , \19923 , \4454 );
and \U$18942 ( \19925 , \19919 , \19924 );
and \U$18943 ( \19926 , \19915 , \19924 );
or \U$18944 ( \19927 , \19920 , \19925 , \19926 );
and \U$18945 ( \19928 , \19911 , \19927 );
xor \U$18946 ( \19929 , \19739 , \19743 );
xor \U$18947 ( \19930 , \19929 , \19748 );
and \U$18948 ( \19931 , \19927 , \19930 );
and \U$18949 ( \19932 , \19911 , \19930 );
or \U$18950 ( \19933 , \19928 , \19931 , \19932 );
and \U$18951 ( \19934 , \19895 , \19933 );
xor \U$18952 ( \19935 , \19687 , \19691 );
xor \U$18953 ( \19936 , \19935 , \19696 );
xor \U$18954 ( \19937 , \19703 , \19707 );
xor \U$18955 ( \19938 , \19937 , \19712 );
and \U$18956 ( \19939 , \19936 , \19938 );
xor \U$18957 ( \19940 , \19755 , \19759 );
xor \U$18958 ( \19941 , \19940 , \19764 );
and \U$18959 ( \19942 , \19938 , \19941 );
and \U$18960 ( \19943 , \19936 , \19941 );
or \U$18961 ( \19944 , \19939 , \19942 , \19943 );
and \U$18962 ( \19945 , \19933 , \19944 );
and \U$18963 ( \19946 , \19895 , \19944 );
or \U$18964 ( \19947 , \19934 , \19945 , \19946 );
xor \U$18965 ( \19948 , \19751 , \19767 );
xor \U$18966 ( \19949 , \19948 , \19772 );
xor \U$18967 ( \19950 , \19791 , \19793 );
xor \U$18968 ( \19951 , \19950 , \19796 );
and \U$18969 ( \19952 , \19949 , \19951 );
xor \U$18970 ( \19953 , \19778 , \19780 );
xor \U$18971 ( \19954 , \19953 , \19783 );
and \U$18972 ( \19955 , \19951 , \19954 );
and \U$18973 ( \19956 , \19949 , \19954 );
or \U$18974 ( \19957 , \19952 , \19955 , \19956 );
and \U$18975 ( \19958 , \19947 , \19957 );
xor \U$18976 ( \19959 , \19810 , \19812 );
xor \U$18977 ( \19960 , \19959 , \19815 );
and \U$18978 ( \19961 , \19957 , \19960 );
and \U$18979 ( \19962 , \19947 , \19960 );
or \U$18980 ( \19963 , \19958 , \19961 , \19962 );
xor \U$18981 ( \19964 , \19735 , \19775 );
xor \U$18982 ( \19965 , \19964 , \19786 );
xor \U$18983 ( \19966 , \19799 , \19801 );
xor \U$18984 ( \19967 , \19966 , \19804 );
and \U$18985 ( \19968 , \19965 , \19967 );
and \U$18986 ( \19969 , \19963 , \19968 );
xor \U$18987 ( \19970 , \19823 , \19825 );
xor \U$18988 ( \19971 , \19970 , \19827 );
and \U$18989 ( \19972 , \19968 , \19971 );
and \U$18990 ( \19973 , \19963 , \19971 );
or \U$18991 ( \19974 , \19969 , \19972 , \19973 );
xor \U$18992 ( \19975 , \19633 , \19643 );
xor \U$18993 ( \19976 , \19975 , \19649 );
and \U$18994 ( \19977 , \19974 , \19976 );
xor \U$18995 ( \19978 , \19821 , \19830 );
xor \U$18996 ( \19979 , \19978 , \19833 );
and \U$18997 ( \19980 , \19976 , \19979 );
and \U$18998 ( \19981 , \19974 , \19979 );
or \U$18999 ( \19982 , \19977 , \19980 , \19981 );
and \U$19000 ( \19983 , \19847 , \19982 );
xor \U$19001 ( \19984 , \19847 , \19982 );
xor \U$19002 ( \19985 , \19974 , \19976 );
xor \U$19003 ( \19986 , \19985 , \19979 );
and \U$19004 ( \19987 , \4684 , \11482 );
and \U$19005 ( \19988 , \4679 , \11479 );
nor \U$19006 ( \19989 , \19987 , \19988 );
xnor \U$19007 ( \19990 , \19989 , \10427 );
and \U$19008 ( \19991 , \5137 , \10669 );
and \U$19009 ( \19992 , \4940 , \10667 );
nor \U$19010 ( \19993 , \19991 , \19992 );
xnor \U$19011 ( \19994 , \19993 , \10430 );
and \U$19012 ( \19995 , \19990 , \19994 );
and \U$19013 ( \19996 , \5447 , \10101 );
and \U$19014 ( \19997 , \5439 , \10099 );
nor \U$19015 ( \19998 , \19996 , \19997 );
xnor \U$19016 ( \19999 , \19998 , \9791 );
and \U$19017 ( \20000 , \19994 , \19999 );
and \U$19018 ( \20001 , \19990 , \19999 );
or \U$19019 ( \20002 , \19995 , \20000 , \20001 );
and \U$19020 ( \20003 , \7370 , \7906 );
and \U$19021 ( \20004 , \7168 , \7904 );
nor \U$19022 ( \20005 , \20003 , \20004 );
xnor \U$19023 ( \20006 , \20005 , \7646 );
and \U$19024 ( \20007 , \7845 , \7412 );
and \U$19025 ( \20008 , \7673 , \7410 );
nor \U$19026 ( \20009 , \20007 , \20008 );
xnor \U$19027 ( \20010 , \20009 , \7097 );
and \U$19028 ( \20011 , \20006 , \20010 );
and \U$19029 ( \20012 , \8795 , \6903 );
and \U$19030 ( \20013 , \8371 , \6901 );
nor \U$19031 ( \20014 , \20012 , \20013 );
xnor \U$19032 ( \20015 , \20014 , \6563 );
and \U$19033 ( \20016 , \20010 , \20015 );
and \U$19034 ( \20017 , \20006 , \20015 );
or \U$19035 ( \20018 , \20011 , \20016 , \20017 );
and \U$19036 ( \20019 , \20002 , \20018 );
and \U$19037 ( \20020 , \5921 , \9564 );
and \U$19038 ( \20021 , \5916 , \9562 );
nor \U$19039 ( \20022 , \20020 , \20021 );
xnor \U$19040 ( \20023 , \20022 , \9193 );
and \U$19041 ( \20024 , \6444 , \9002 );
and \U$19042 ( \20025 , \6185 , \9000 );
nor \U$19043 ( \20026 , \20024 , \20025 );
xnor \U$19044 ( \20027 , \20026 , \8684 );
and \U$19045 ( \20028 , \20023 , \20027 );
and \U$19046 ( \20029 , \6825 , \8435 );
and \U$19047 ( \20030 , \6816 , \8433 );
nor \U$19048 ( \20031 , \20029 , \20030 );
xnor \U$19049 ( \20032 , \20031 , \8186 );
and \U$19050 ( \20033 , \20027 , \20032 );
and \U$19051 ( \20034 , \20023 , \20032 );
or \U$19052 ( \20035 , \20028 , \20033 , \20034 );
and \U$19053 ( \20036 , \20018 , \20035 );
and \U$19054 ( \20037 , \20002 , \20035 );
or \U$19055 ( \20038 , \20019 , \20036 , \20037 );
xor \U$19056 ( \20039 , \19851 , \19855 );
xor \U$19057 ( \20040 , \20039 , \19860 );
xor \U$19058 ( \20041 , \19867 , \19871 );
xor \U$19059 ( \20042 , \20041 , \19876 );
and \U$19060 ( \20043 , \20040 , \20042 );
xor \U$19061 ( \20044 , \19899 , \19903 );
xor \U$19062 ( \20045 , \20044 , \19908 );
and \U$19063 ( \20046 , \20042 , \20045 );
and \U$19064 ( \20047 , \20040 , \20045 );
or \U$19065 ( \20048 , \20043 , \20046 , \20047 );
and \U$19066 ( \20049 , \20038 , \20048 );
and \U$19067 ( \20050 , \9046 , \6314 );
and \U$19068 ( \20051 , \9041 , \6312 );
nor \U$19069 ( \20052 , \20050 , \20051 );
xnor \U$19070 ( \20053 , \20052 , \6073 );
and \U$19071 ( \20054 , \9649 , \5848 );
and \U$19072 ( \20055 , \9365 , \5846 );
nor \U$19073 ( \20056 , \20054 , \20055 );
xnor \U$19074 ( \20057 , \20056 , \5660 );
and \U$19075 ( \20058 , \20053 , \20057 );
and \U$19076 ( \20059 , \10226 , \5474 );
and \U$19077 ( \20060 , \10218 , \5472 );
nor \U$19078 ( \20061 , \20059 , \20060 );
xnor \U$19079 ( \20062 , \20061 , \5242 );
and \U$19080 ( \20063 , \20057 , \20062 );
and \U$19081 ( \20064 , \20053 , \20062 );
or \U$19082 ( \20065 , \20058 , \20063 , \20064 );
nand \U$19083 ( \20066 , \11635 , \4303 );
xnor \U$19084 ( \20067 , \20066 , \4118 );
and \U$19085 ( \20068 , \20065 , \20067 );
xor \U$19086 ( \20069 , \19915 , \19919 );
xor \U$19087 ( \20070 , \20069 , \19924 );
and \U$19088 ( \20071 , \20067 , \20070 );
and \U$19089 ( \20072 , \20065 , \20070 );
or \U$19090 ( \20073 , \20068 , \20071 , \20072 );
and \U$19091 ( \20074 , \20048 , \20073 );
and \U$19092 ( \20075 , \20038 , \20073 );
or \U$19093 ( \20076 , \20049 , \20074 , \20075 );
xor \U$19094 ( \20077 , \19720 , \19724 );
xor \U$19095 ( \20078 , \20077 , \19729 );
xor \U$19096 ( \20079 , \19911 , \19927 );
xor \U$19097 ( \20080 , \20079 , \19930 );
and \U$19098 ( \20081 , \20078 , \20080 );
xor \U$19099 ( \20082 , \19936 , \19938 );
xor \U$19100 ( \20083 , \20082 , \19941 );
and \U$19101 ( \20084 , \20080 , \20083 );
and \U$19102 ( \20085 , \20078 , \20083 );
or \U$19103 ( \20086 , \20081 , \20084 , \20085 );
and \U$19104 ( \20087 , \20076 , \20086 );
xor \U$19105 ( \20088 , \19699 , \19715 );
xor \U$19106 ( \20089 , \20088 , \19732 );
and \U$19107 ( \20090 , \20086 , \20089 );
and \U$19108 ( \20091 , \20076 , \20089 );
or \U$19109 ( \20092 , \20087 , \20090 , \20091 );
xor \U$19110 ( \20093 , \19947 , \19957 );
xor \U$19111 ( \20094 , \20093 , \19960 );
and \U$19112 ( \20095 , \20092 , \20094 );
xor \U$19113 ( \20096 , \19965 , \19967 );
and \U$19114 ( \20097 , \20094 , \20096 );
and \U$19115 ( \20098 , \20092 , \20096 );
or \U$19116 ( \20099 , \20095 , \20097 , \20098 );
xor \U$19117 ( \20100 , \19789 , \19807 );
xor \U$19118 ( \20101 , \20100 , \19818 );
and \U$19119 ( \20102 , \20099 , \20101 );
xor \U$19120 ( \20103 , \19963 , \19968 );
xor \U$19121 ( \20104 , \20103 , \19971 );
and \U$19122 ( \20105 , \20101 , \20104 );
and \U$19123 ( \20106 , \20099 , \20104 );
or \U$19124 ( \20107 , \20102 , \20105 , \20106 );
and \U$19125 ( \20108 , \19986 , \20107 );
xor \U$19126 ( \20109 , \19986 , \20107 );
xor \U$19127 ( \20110 , \20099 , \20101 );
xor \U$19128 ( \20111 , \20110 , \20104 );
and \U$19129 ( \20112 , \9041 , \6903 );
and \U$19130 ( \20113 , \8795 , \6901 );
nor \U$19131 ( \20114 , \20112 , \20113 );
xnor \U$19132 ( \20115 , \20114 , \6563 );
and \U$19133 ( \20116 , \9365 , \6314 );
and \U$19134 ( \20117 , \9046 , \6312 );
nor \U$19135 ( \20118 , \20116 , \20117 );
xnor \U$19136 ( \20119 , \20118 , \6073 );
and \U$19137 ( \20120 , \20115 , \20119 );
and \U$19138 ( \20121 , \10218 , \5848 );
and \U$19139 ( \20122 , \9649 , \5846 );
nor \U$19140 ( \20123 , \20121 , \20122 );
xnor \U$19141 ( \20124 , \20123 , \5660 );
and \U$19142 ( \20125 , \20119 , \20124 );
and \U$19143 ( \20126 , \20115 , \20124 );
or \U$19144 ( \20127 , \20120 , \20125 , \20126 );
and \U$19145 ( \20128 , \10829 , \5474 );
and \U$19146 ( \20129 , \10226 , \5472 );
nor \U$19147 ( \20130 , \20128 , \20129 );
xnor \U$19148 ( \20131 , \20130 , \5242 );
and \U$19149 ( \20132 , \11015 , \5023 );
and \U$19150 ( \20133 , \10834 , \5021 );
nor \U$19151 ( \20134 , \20132 , \20133 );
xnor \U$19152 ( \20135 , \20134 , \4880 );
and \U$19153 ( \20136 , \20131 , \20135 );
nand \U$19154 ( \20137 , \11635 , \4698 );
xnor \U$19155 ( \20138 , \20137 , \4454 );
and \U$19156 ( \20139 , \20135 , \20138 );
and \U$19157 ( \20140 , \20131 , \20138 );
or \U$19158 ( \20141 , \20136 , \20139 , \20140 );
and \U$19159 ( \20142 , \20127 , \20141 );
and \U$19160 ( \20143 , \10834 , \5023 );
and \U$19161 ( \20144 , \10829 , \5021 );
nor \U$19162 ( \20145 , \20143 , \20144 );
xnor \U$19163 ( \20146 , \20145 , \4880 );
and \U$19164 ( \20147 , \20141 , \20146 );
and \U$19165 ( \20148 , \20127 , \20146 );
or \U$19166 ( \20149 , \20142 , \20147 , \20148 );
and \U$19167 ( \20150 , \7168 , \8435 );
and \U$19168 ( \20151 , \6825 , \8433 );
nor \U$19169 ( \20152 , \20150 , \20151 );
xnor \U$19170 ( \20153 , \20152 , \8186 );
and \U$19171 ( \20154 , \7673 , \7906 );
and \U$19172 ( \20155 , \7370 , \7904 );
nor \U$19173 ( \20156 , \20154 , \20155 );
xnor \U$19174 ( \20157 , \20156 , \7646 );
and \U$19175 ( \20158 , \20153 , \20157 );
and \U$19176 ( \20159 , \8371 , \7412 );
and \U$19177 ( \20160 , \7845 , \7410 );
nor \U$19178 ( \20161 , \20159 , \20160 );
xnor \U$19179 ( \20162 , \20161 , \7097 );
and \U$19180 ( \20163 , \20157 , \20162 );
and \U$19181 ( \20164 , \20153 , \20162 );
or \U$19182 ( \20165 , \20158 , \20163 , \20164 );
and \U$19183 ( \20166 , \4940 , \11482 );
and \U$19184 ( \20167 , \4684 , \11479 );
nor \U$19185 ( \20168 , \20166 , \20167 );
xnor \U$19186 ( \20169 , \20168 , \10427 );
and \U$19187 ( \20170 , \5439 , \10669 );
and \U$19188 ( \20171 , \5137 , \10667 );
nor \U$19189 ( \20172 , \20170 , \20171 );
xnor \U$19190 ( \20173 , \20172 , \10430 );
and \U$19191 ( \20174 , \20169 , \20173 );
and \U$19192 ( \20175 , \20173 , \4454 );
and \U$19193 ( \20176 , \20169 , \4454 );
or \U$19194 ( \20177 , \20174 , \20175 , \20176 );
and \U$19195 ( \20178 , \20165 , \20177 );
and \U$19196 ( \20179 , \5916 , \10101 );
and \U$19197 ( \20180 , \5447 , \10099 );
nor \U$19198 ( \20181 , \20179 , \20180 );
xnor \U$19199 ( \20182 , \20181 , \9791 );
and \U$19200 ( \20183 , \6185 , \9564 );
and \U$19201 ( \20184 , \5921 , \9562 );
nor \U$19202 ( \20185 , \20183 , \20184 );
xnor \U$19203 ( \20186 , \20185 , \9193 );
and \U$19204 ( \20187 , \20182 , \20186 );
and \U$19205 ( \20188 , \6816 , \9002 );
and \U$19206 ( \20189 , \6444 , \9000 );
nor \U$19207 ( \20190 , \20188 , \20189 );
xnor \U$19208 ( \20191 , \20190 , \8684 );
and \U$19209 ( \20192 , \20186 , \20191 );
and \U$19210 ( \20193 , \20182 , \20191 );
or \U$19211 ( \20194 , \20187 , \20192 , \20193 );
and \U$19212 ( \20195 , \20177 , \20194 );
and \U$19213 ( \20196 , \20165 , \20194 );
or \U$19214 ( \20197 , \20178 , \20195 , \20196 );
and \U$19215 ( \20198 , \20149 , \20197 );
and \U$19216 ( \20199 , \11635 , \4700 );
and \U$19217 ( \20200 , \11015 , \4698 );
nor \U$19218 ( \20201 , \20199 , \20200 );
xnor \U$19219 ( \20202 , \20201 , \4454 );
xor \U$19220 ( \20203 , \20053 , \20057 );
xor \U$19221 ( \20204 , \20203 , \20062 );
and \U$19222 ( \20205 , \20202 , \20204 );
xor \U$19223 ( \20206 , \20006 , \20010 );
xor \U$19224 ( \20207 , \20206 , \20015 );
and \U$19225 ( \20208 , \20204 , \20207 );
and \U$19226 ( \20209 , \20202 , \20207 );
or \U$19227 ( \20210 , \20205 , \20208 , \20209 );
and \U$19228 ( \20211 , \20197 , \20210 );
and \U$19229 ( \20212 , \20149 , \20210 );
or \U$19230 ( \20213 , \20198 , \20211 , \20212 );
xor \U$19231 ( \20214 , \19884 , \19888 );
xor \U$19232 ( \20215 , \20214 , \4118 );
xor \U$19233 ( \20216 , \20040 , \20042 );
xor \U$19234 ( \20217 , \20216 , \20045 );
and \U$19235 ( \20218 , \20215 , \20217 );
xor \U$19236 ( \20219 , \20065 , \20067 );
xor \U$19237 ( \20220 , \20219 , \20070 );
and \U$19238 ( \20221 , \20217 , \20220 );
and \U$19239 ( \20222 , \20215 , \20220 );
or \U$19240 ( \20223 , \20218 , \20221 , \20222 );
and \U$19241 ( \20224 , \20213 , \20223 );
xor \U$19242 ( \20225 , \19863 , \19879 );
xor \U$19243 ( \20226 , \20225 , \19892 );
and \U$19244 ( \20227 , \20223 , \20226 );
and \U$19245 ( \20228 , \20213 , \20226 );
or \U$19246 ( \20229 , \20224 , \20227 , \20228 );
xor \U$19247 ( \20230 , \20038 , \20048 );
xor \U$19248 ( \20231 , \20230 , \20073 );
xor \U$19249 ( \20232 , \20078 , \20080 );
xor \U$19250 ( \20233 , \20232 , \20083 );
and \U$19251 ( \20234 , \20231 , \20233 );
and \U$19252 ( \20235 , \20229 , \20234 );
xor \U$19253 ( \20236 , \19949 , \19951 );
xor \U$19254 ( \20237 , \20236 , \19954 );
and \U$19255 ( \20238 , \20234 , \20237 );
and \U$19256 ( \20239 , \20229 , \20237 );
or \U$19257 ( \20240 , \20235 , \20238 , \20239 );
xor \U$19258 ( \20241 , \19895 , \19933 );
xor \U$19259 ( \20242 , \20241 , \19944 );
xor \U$19260 ( \20243 , \20076 , \20086 );
xor \U$19261 ( \20244 , \20243 , \20089 );
and \U$19262 ( \20245 , \20242 , \20244 );
and \U$19263 ( \20246 , \20240 , \20245 );
xor \U$19264 ( \20247 , \20092 , \20094 );
xor \U$19265 ( \20248 , \20247 , \20096 );
and \U$19266 ( \20249 , \20245 , \20248 );
and \U$19267 ( \20250 , \20240 , \20248 );
or \U$19268 ( \20251 , \20246 , \20249 , \20250 );
and \U$19269 ( \20252 , \20111 , \20251 );
xor \U$19270 ( \20253 , \20111 , \20251 );
xor \U$19271 ( \20254 , \20240 , \20245 );
xor \U$19272 ( \20255 , \20254 , \20248 );
and \U$19273 ( \20256 , \6444 , \9564 );
and \U$19274 ( \20257 , \6185 , \9562 );
nor \U$19275 ( \20258 , \20256 , \20257 );
xnor \U$19276 ( \20259 , \20258 , \9193 );
and \U$19277 ( \20260 , \6825 , \9002 );
and \U$19278 ( \20261 , \6816 , \9000 );
nor \U$19279 ( \20262 , \20260 , \20261 );
xnor \U$19280 ( \20263 , \20262 , \8684 );
and \U$19281 ( \20264 , \20259 , \20263 );
and \U$19282 ( \20265 , \7370 , \8435 );
and \U$19283 ( \20266 , \7168 , \8433 );
nor \U$19284 ( \20267 , \20265 , \20266 );
xnor \U$19285 ( \20268 , \20267 , \8186 );
and \U$19286 ( \20269 , \20263 , \20268 );
and \U$19287 ( \20270 , \20259 , \20268 );
or \U$19288 ( \20271 , \20264 , \20269 , \20270 );
and \U$19289 ( \20272 , \5137 , \11482 );
and \U$19290 ( \20273 , \4940 , \11479 );
nor \U$19291 ( \20274 , \20272 , \20273 );
xnor \U$19292 ( \20275 , \20274 , \10427 );
and \U$19293 ( \20276 , \5447 , \10669 );
and \U$19294 ( \20277 , \5439 , \10667 );
nor \U$19295 ( \20278 , \20276 , \20277 );
xnor \U$19296 ( \20279 , \20278 , \10430 );
and \U$19297 ( \20280 , \20275 , \20279 );
and \U$19298 ( \20281 , \5921 , \10101 );
and \U$19299 ( \20282 , \5916 , \10099 );
nor \U$19300 ( \20283 , \20281 , \20282 );
xnor \U$19301 ( \20284 , \20283 , \9791 );
and \U$19302 ( \20285 , \20279 , \20284 );
and \U$19303 ( \20286 , \20275 , \20284 );
or \U$19304 ( \20287 , \20280 , \20285 , \20286 );
and \U$19305 ( \20288 , \20271 , \20287 );
and \U$19306 ( \20289 , \7845 , \7906 );
and \U$19307 ( \20290 , \7673 , \7904 );
nor \U$19308 ( \20291 , \20289 , \20290 );
xnor \U$19309 ( \20292 , \20291 , \7646 );
and \U$19310 ( \20293 , \8795 , \7412 );
and \U$19311 ( \20294 , \8371 , \7410 );
nor \U$19312 ( \20295 , \20293 , \20294 );
xnor \U$19313 ( \20296 , \20295 , \7097 );
and \U$19314 ( \20297 , \20292 , \20296 );
and \U$19315 ( \20298 , \9046 , \6903 );
and \U$19316 ( \20299 , \9041 , \6901 );
nor \U$19317 ( \20300 , \20298 , \20299 );
xnor \U$19318 ( \20301 , \20300 , \6563 );
and \U$19319 ( \20302 , \20296 , \20301 );
and \U$19320 ( \20303 , \20292 , \20301 );
or \U$19321 ( \20304 , \20297 , \20302 , \20303 );
and \U$19322 ( \20305 , \20287 , \20304 );
and \U$19323 ( \20306 , \20271 , \20304 );
or \U$19324 ( \20307 , \20288 , \20305 , \20306 );
xor \U$19325 ( \20308 , \20153 , \20157 );
xor \U$19326 ( \20309 , \20308 , \20162 );
xor \U$19327 ( \20310 , \20169 , \20173 );
xor \U$19328 ( \20311 , \20310 , \4454 );
and \U$19329 ( \20312 , \20309 , \20311 );
xor \U$19330 ( \20313 , \20182 , \20186 );
xor \U$19331 ( \20314 , \20313 , \20191 );
and \U$19332 ( \20315 , \20311 , \20314 );
and \U$19333 ( \20316 , \20309 , \20314 );
or \U$19334 ( \20317 , \20312 , \20315 , \20316 );
and \U$19335 ( \20318 , \20307 , \20317 );
and \U$19336 ( \20319 , \9649 , \6314 );
and \U$19337 ( \20320 , \9365 , \6312 );
nor \U$19338 ( \20321 , \20319 , \20320 );
xnor \U$19339 ( \20322 , \20321 , \6073 );
and \U$19340 ( \20323 , \10226 , \5848 );
and \U$19341 ( \20324 , \10218 , \5846 );
nor \U$19342 ( \20325 , \20323 , \20324 );
xnor \U$19343 ( \20326 , \20325 , \5660 );
and \U$19344 ( \20327 , \20322 , \20326 );
and \U$19345 ( \20328 , \10834 , \5474 );
and \U$19346 ( \20329 , \10829 , \5472 );
nor \U$19347 ( \20330 , \20328 , \20329 );
xnor \U$19348 ( \20331 , \20330 , \5242 );
and \U$19349 ( \20332 , \20326 , \20331 );
and \U$19350 ( \20333 , \20322 , \20331 );
or \U$19351 ( \20334 , \20327 , \20332 , \20333 );
xor \U$19352 ( \20335 , \20115 , \20119 );
xor \U$19353 ( \20336 , \20335 , \20124 );
and \U$19354 ( \20337 , \20334 , \20336 );
xor \U$19355 ( \20338 , \20131 , \20135 );
xor \U$19356 ( \20339 , \20338 , \20138 );
and \U$19357 ( \20340 , \20336 , \20339 );
and \U$19358 ( \20341 , \20334 , \20339 );
or \U$19359 ( \20342 , \20337 , \20340 , \20341 );
and \U$19360 ( \20343 , \20317 , \20342 );
and \U$19361 ( \20344 , \20307 , \20342 );
or \U$19362 ( \20345 , \20318 , \20343 , \20344 );
xor \U$19363 ( \20346 , \19990 , \19994 );
xor \U$19364 ( \20347 , \20346 , \19999 );
xor \U$19365 ( \20348 , \20023 , \20027 );
xor \U$19366 ( \20349 , \20348 , \20032 );
and \U$19367 ( \20350 , \20347 , \20349 );
xor \U$19368 ( \20351 , \20202 , \20204 );
xor \U$19369 ( \20352 , \20351 , \20207 );
and \U$19370 ( \20353 , \20349 , \20352 );
and \U$19371 ( \20354 , \20347 , \20352 );
or \U$19372 ( \20355 , \20350 , \20353 , \20354 );
and \U$19373 ( \20356 , \20345 , \20355 );
xor \U$19374 ( \20357 , \20002 , \20018 );
xor \U$19375 ( \20358 , \20357 , \20035 );
and \U$19376 ( \20359 , \20355 , \20358 );
and \U$19377 ( \20360 , \20345 , \20358 );
or \U$19378 ( \20361 , \20356 , \20359 , \20360 );
xor \U$19379 ( \20362 , \20213 , \20223 );
xor \U$19380 ( \20363 , \20362 , \20226 );
and \U$19381 ( \20364 , \20361 , \20363 );
xor \U$19382 ( \20365 , \20231 , \20233 );
and \U$19383 ( \20366 , \20363 , \20365 );
and \U$19384 ( \20367 , \20361 , \20365 );
or \U$19385 ( \20368 , \20364 , \20366 , \20367 );
xor \U$19386 ( \20369 , \20229 , \20234 );
xor \U$19387 ( \20370 , \20369 , \20237 );
and \U$19388 ( \20371 , \20368 , \20370 );
xor \U$19389 ( \20372 , \20242 , \20244 );
and \U$19390 ( \20373 , \20370 , \20372 );
and \U$19391 ( \20374 , \20368 , \20372 );
or \U$19392 ( \20375 , \20371 , \20373 , \20374 );
and \U$19393 ( \20376 , \20255 , \20375 );
xor \U$19394 ( \20377 , \20255 , \20375 );
xor \U$19395 ( \20378 , \20368 , \20370 );
xor \U$19396 ( \20379 , \20378 , \20372 );
and \U$19397 ( \20380 , \6185 , \10101 );
and \U$19398 ( \20381 , \5921 , \10099 );
nor \U$19399 ( \20382 , \20380 , \20381 );
xnor \U$19400 ( \20383 , \20382 , \9791 );
and \U$19401 ( \20384 , \6816 , \9564 );
and \U$19402 ( \20385 , \6444 , \9562 );
nor \U$19403 ( \20386 , \20384 , \20385 );
xnor \U$19404 ( \20387 , \20386 , \9193 );
and \U$19405 ( \20388 , \20383 , \20387 );
and \U$19406 ( \20389 , \7168 , \9002 );
and \U$19407 ( \20390 , \6825 , \9000 );
nor \U$19408 ( \20391 , \20389 , \20390 );
xnor \U$19409 ( \20392 , \20391 , \8684 );
and \U$19410 ( \20393 , \20387 , \20392 );
and \U$19411 ( \20394 , \20383 , \20392 );
or \U$19412 ( \20395 , \20388 , \20393 , \20394 );
and \U$19413 ( \20396 , \5439 , \11482 );
and \U$19414 ( \20397 , \5137 , \11479 );
nor \U$19415 ( \20398 , \20396 , \20397 );
xnor \U$19416 ( \20399 , \20398 , \10427 );
and \U$19417 ( \20400 , \5916 , \10669 );
and \U$19418 ( \20401 , \5447 , \10667 );
nor \U$19419 ( \20402 , \20400 , \20401 );
xnor \U$19420 ( \20403 , \20402 , \10430 );
and \U$19421 ( \20404 , \20399 , \20403 );
and \U$19422 ( \20405 , \20403 , \4880 );
and \U$19423 ( \20406 , \20399 , \4880 );
or \U$19424 ( \20407 , \20404 , \20405 , \20406 );
and \U$19425 ( \20408 , \20395 , \20407 );
and \U$19426 ( \20409 , \7673 , \8435 );
and \U$19427 ( \20410 , \7370 , \8433 );
nor \U$19428 ( \20411 , \20409 , \20410 );
xnor \U$19429 ( \20412 , \20411 , \8186 );
and \U$19430 ( \20413 , \8371 , \7906 );
and \U$19431 ( \20414 , \7845 , \7904 );
nor \U$19432 ( \20415 , \20413 , \20414 );
xnor \U$19433 ( \20416 , \20415 , \7646 );
and \U$19434 ( \20417 , \20412 , \20416 );
and \U$19435 ( \20418 , \9041 , \7412 );
and \U$19436 ( \20419 , \8795 , \7410 );
nor \U$19437 ( \20420 , \20418 , \20419 );
xnor \U$19438 ( \20421 , \20420 , \7097 );
and \U$19439 ( \20422 , \20416 , \20421 );
and \U$19440 ( \20423 , \20412 , \20421 );
or \U$19441 ( \20424 , \20417 , \20422 , \20423 );
and \U$19442 ( \20425 , \20407 , \20424 );
and \U$19443 ( \20426 , \20395 , \20424 );
or \U$19444 ( \20427 , \20408 , \20425 , \20426 );
and \U$19445 ( \20428 , \9365 , \6903 );
and \U$19446 ( \20429 , \9046 , \6901 );
nor \U$19447 ( \20430 , \20428 , \20429 );
xnor \U$19448 ( \20431 , \20430 , \6563 );
and \U$19449 ( \20432 , \10218 , \6314 );
and \U$19450 ( \20433 , \9649 , \6312 );
nor \U$19451 ( \20434 , \20432 , \20433 );
xnor \U$19452 ( \20435 , \20434 , \6073 );
and \U$19453 ( \20436 , \20431 , \20435 );
and \U$19454 ( \20437 , \10829 , \5848 );
and \U$19455 ( \20438 , \10226 , \5846 );
nor \U$19456 ( \20439 , \20437 , \20438 );
xnor \U$19457 ( \20440 , \20439 , \5660 );
and \U$19458 ( \20441 , \20435 , \20440 );
and \U$19459 ( \20442 , \20431 , \20440 );
or \U$19460 ( \20443 , \20436 , \20441 , \20442 );
and \U$19461 ( \20444 , \11015 , \5474 );
and \U$19462 ( \20445 , \10834 , \5472 );
nor \U$19463 ( \20446 , \20444 , \20445 );
xnor \U$19464 ( \20447 , \20446 , \5242 );
nand \U$19465 ( \20448 , \11635 , \5021 );
xnor \U$19466 ( \20449 , \20448 , \4880 );
and \U$19467 ( \20450 , \20447 , \20449 );
and \U$19468 ( \20451 , \20443 , \20450 );
and \U$19469 ( \20452 , \11635 , \5023 );
and \U$19470 ( \20453 , \11015 , \5021 );
nor \U$19471 ( \20454 , \20452 , \20453 );
xnor \U$19472 ( \20455 , \20454 , \4880 );
and \U$19473 ( \20456 , \20450 , \20455 );
and \U$19474 ( \20457 , \20443 , \20455 );
or \U$19475 ( \20458 , \20451 , \20456 , \20457 );
and \U$19476 ( \20459 , \20427 , \20458 );
xor \U$19477 ( \20460 , \20259 , \20263 );
xor \U$19478 ( \20461 , \20460 , \20268 );
xor \U$19479 ( \20462 , \20322 , \20326 );
xor \U$19480 ( \20463 , \20462 , \20331 );
and \U$19481 ( \20464 , \20461 , \20463 );
xor \U$19482 ( \20465 , \20292 , \20296 );
xor \U$19483 ( \20466 , \20465 , \20301 );
and \U$19484 ( \20467 , \20463 , \20466 );
and \U$19485 ( \20468 , \20461 , \20466 );
or \U$19486 ( \20469 , \20464 , \20467 , \20468 );
and \U$19487 ( \20470 , \20458 , \20469 );
and \U$19488 ( \20471 , \20427 , \20469 );
or \U$19489 ( \20472 , \20459 , \20470 , \20471 );
xor \U$19490 ( \20473 , \20271 , \20287 );
xor \U$19491 ( \20474 , \20473 , \20304 );
xor \U$19492 ( \20475 , \20309 , \20311 );
xor \U$19493 ( \20476 , \20475 , \20314 );
and \U$19494 ( \20477 , \20474 , \20476 );
xor \U$19495 ( \20478 , \20334 , \20336 );
xor \U$19496 ( \20479 , \20478 , \20339 );
and \U$19497 ( \20480 , \20476 , \20479 );
and \U$19498 ( \20481 , \20474 , \20479 );
or \U$19499 ( \20482 , \20477 , \20480 , \20481 );
and \U$19500 ( \20483 , \20472 , \20482 );
xor \U$19501 ( \20484 , \20127 , \20141 );
xor \U$19502 ( \20485 , \20484 , \20146 );
and \U$19503 ( \20486 , \20482 , \20485 );
and \U$19504 ( \20487 , \20472 , \20485 );
or \U$19505 ( \20488 , \20483 , \20486 , \20487 );
xor \U$19506 ( \20489 , \20165 , \20177 );
xor \U$19507 ( \20490 , \20489 , \20194 );
xor \U$19508 ( \20491 , \20307 , \20317 );
xor \U$19509 ( \20492 , \20491 , \20342 );
and \U$19510 ( \20493 , \20490 , \20492 );
xor \U$19511 ( \20494 , \20347 , \20349 );
xor \U$19512 ( \20495 , \20494 , \20352 );
and \U$19513 ( \20496 , \20492 , \20495 );
and \U$19514 ( \20497 , \20490 , \20495 );
or \U$19515 ( \20498 , \20493 , \20496 , \20497 );
and \U$19516 ( \20499 , \20488 , \20498 );
xor \U$19517 ( \20500 , \20215 , \20217 );
xor \U$19518 ( \20501 , \20500 , \20220 );
and \U$19519 ( \20502 , \20498 , \20501 );
and \U$19520 ( \20503 , \20488 , \20501 );
or \U$19521 ( \20504 , \20499 , \20502 , \20503 );
xor \U$19522 ( \20505 , \20149 , \20197 );
xor \U$19523 ( \20506 , \20505 , \20210 );
xor \U$19524 ( \20507 , \20345 , \20355 );
xor \U$19525 ( \20508 , \20507 , \20358 );
and \U$19526 ( \20509 , \20506 , \20508 );
and \U$19527 ( \20510 , \20504 , \20509 );
xor \U$19528 ( \20511 , \20361 , \20363 );
xor \U$19529 ( \20512 , \20511 , \20365 );
and \U$19530 ( \20513 , \20509 , \20512 );
and \U$19531 ( \20514 , \20504 , \20512 );
or \U$19532 ( \20515 , \20510 , \20513 , \20514 );
and \U$19533 ( \20516 , \20379 , \20515 );
xor \U$19534 ( \20517 , \20379 , \20515 );
xor \U$19535 ( \20518 , \20504 , \20509 );
xor \U$19536 ( \20519 , \20518 , \20512 );
and \U$19537 ( \20520 , \6825 , \9564 );
and \U$19538 ( \20521 , \6816 , \9562 );
nor \U$19539 ( \20522 , \20520 , \20521 );
xnor \U$19540 ( \20523 , \20522 , \9193 );
and \U$19541 ( \20524 , \7370 , \9002 );
and \U$19542 ( \20525 , \7168 , \9000 );
nor \U$19543 ( \20526 , \20524 , \20525 );
xnor \U$19544 ( \20527 , \20526 , \8684 );
and \U$19545 ( \20528 , \20523 , \20527 );
and \U$19546 ( \20529 , \7845 , \8435 );
and \U$19547 ( \20530 , \7673 , \8433 );
nor \U$19548 ( \20531 , \20529 , \20530 );
xnor \U$19549 ( \20532 , \20531 , \8186 );
and \U$19550 ( \20533 , \20527 , \20532 );
and \U$19551 ( \20534 , \20523 , \20532 );
or \U$19552 ( \20535 , \20528 , \20533 , \20534 );
and \U$19553 ( \20536 , \8795 , \7906 );
and \U$19554 ( \20537 , \8371 , \7904 );
nor \U$19555 ( \20538 , \20536 , \20537 );
xnor \U$19556 ( \20539 , \20538 , \7646 );
and \U$19557 ( \20540 , \9046 , \7412 );
and \U$19558 ( \20541 , \9041 , \7410 );
nor \U$19559 ( \20542 , \20540 , \20541 );
xnor \U$19560 ( \20543 , \20542 , \7097 );
and \U$19561 ( \20544 , \20539 , \20543 );
and \U$19562 ( \20545 , \9649 , \6903 );
and \U$19563 ( \20546 , \9365 , \6901 );
nor \U$19564 ( \20547 , \20545 , \20546 );
xnor \U$19565 ( \20548 , \20547 , \6563 );
and \U$19566 ( \20549 , \20543 , \20548 );
and \U$19567 ( \20550 , \20539 , \20548 );
or \U$19568 ( \20551 , \20544 , \20549 , \20550 );
and \U$19569 ( \20552 , \20535 , \20551 );
and \U$19570 ( \20553 , \5447 , \11482 );
and \U$19571 ( \20554 , \5439 , \11479 );
nor \U$19572 ( \20555 , \20553 , \20554 );
xnor \U$19573 ( \20556 , \20555 , \10427 );
and \U$19574 ( \20557 , \5921 , \10669 );
and \U$19575 ( \20558 , \5916 , \10667 );
nor \U$19576 ( \20559 , \20557 , \20558 );
xnor \U$19577 ( \20560 , \20559 , \10430 );
and \U$19578 ( \20561 , \20556 , \20560 );
and \U$19579 ( \20562 , \6444 , \10101 );
and \U$19580 ( \20563 , \6185 , \10099 );
nor \U$19581 ( \20564 , \20562 , \20563 );
xnor \U$19582 ( \20565 , \20564 , \9791 );
and \U$19583 ( \20566 , \20560 , \20565 );
and \U$19584 ( \20567 , \20556 , \20565 );
or \U$19585 ( \20568 , \20561 , \20566 , \20567 );
and \U$19586 ( \20569 , \20551 , \20568 );
and \U$19587 ( \20570 , \20535 , \20568 );
or \U$19588 ( \20571 , \20552 , \20569 , \20570 );
xor \U$19589 ( \20572 , \20383 , \20387 );
xor \U$19590 ( \20573 , \20572 , \20392 );
xor \U$19591 ( \20574 , \20399 , \20403 );
xor \U$19592 ( \20575 , \20574 , \4880 );
and \U$19593 ( \20576 , \20573 , \20575 );
xor \U$19594 ( \20577 , \20412 , \20416 );
xor \U$19595 ( \20578 , \20577 , \20421 );
and \U$19596 ( \20579 , \20575 , \20578 );
and \U$19597 ( \20580 , \20573 , \20578 );
or \U$19598 ( \20581 , \20576 , \20579 , \20580 );
and \U$19599 ( \20582 , \20571 , \20581 );
and \U$19600 ( \20583 , \10226 , \6314 );
and \U$19601 ( \20584 , \10218 , \6312 );
nor \U$19602 ( \20585 , \20583 , \20584 );
xnor \U$19603 ( \20586 , \20585 , \6073 );
and \U$19604 ( \20587 , \10834 , \5848 );
and \U$19605 ( \20588 , \10829 , \5846 );
nor \U$19606 ( \20589 , \20587 , \20588 );
xnor \U$19607 ( \20590 , \20589 , \5660 );
and \U$19608 ( \20591 , \20586 , \20590 );
and \U$19609 ( \20592 , \11635 , \5474 );
and \U$19610 ( \20593 , \11015 , \5472 );
nor \U$19611 ( \20594 , \20592 , \20593 );
xnor \U$19612 ( \20595 , \20594 , \5242 );
and \U$19613 ( \20596 , \20590 , \20595 );
and \U$19614 ( \20597 , \20586 , \20595 );
or \U$19615 ( \20598 , \20591 , \20596 , \20597 );
xor \U$19616 ( \20599 , \20431 , \20435 );
xor \U$19617 ( \20600 , \20599 , \20440 );
and \U$19618 ( \20601 , \20598 , \20600 );
xor \U$19619 ( \20602 , \20447 , \20449 );
and \U$19620 ( \20603 , \20600 , \20602 );
and \U$19621 ( \20604 , \20598 , \20602 );
or \U$19622 ( \20605 , \20601 , \20603 , \20604 );
and \U$19623 ( \20606 , \20581 , \20605 );
and \U$19624 ( \20607 , \20571 , \20605 );
or \U$19625 ( \20608 , \20582 , \20606 , \20607 );
xor \U$19626 ( \20609 , \20275 , \20279 );
xor \U$19627 ( \20610 , \20609 , \20284 );
xor \U$19628 ( \20611 , \20443 , \20450 );
xor \U$19629 ( \20612 , \20611 , \20455 );
and \U$19630 ( \20613 , \20610 , \20612 );
xor \U$19631 ( \20614 , \20461 , \20463 );
xor \U$19632 ( \20615 , \20614 , \20466 );
and \U$19633 ( \20616 , \20612 , \20615 );
and \U$19634 ( \20617 , \20610 , \20615 );
or \U$19635 ( \20618 , \20613 , \20616 , \20617 );
and \U$19636 ( \20619 , \20608 , \20618 );
xor \U$19637 ( \20620 , \20474 , \20476 );
xor \U$19638 ( \20621 , \20620 , \20479 );
and \U$19639 ( \20622 , \20618 , \20621 );
and \U$19640 ( \20623 , \20608 , \20621 );
or \U$19641 ( \20624 , \20619 , \20622 , \20623 );
xor \U$19642 ( \20625 , \20472 , \20482 );
xor \U$19643 ( \20626 , \20625 , \20485 );
and \U$19644 ( \20627 , \20624 , \20626 );
xor \U$19645 ( \20628 , \20490 , \20492 );
xor \U$19646 ( \20629 , \20628 , \20495 );
and \U$19647 ( \20630 , \20626 , \20629 );
and \U$19648 ( \20631 , \20624 , \20629 );
or \U$19649 ( \20632 , \20627 , \20630 , \20631 );
xor \U$19650 ( \20633 , \20488 , \20498 );
xor \U$19651 ( \20634 , \20633 , \20501 );
and \U$19652 ( \20635 , \20632 , \20634 );
xor \U$19653 ( \20636 , \20506 , \20508 );
and \U$19654 ( \20637 , \20634 , \20636 );
and \U$19655 ( \20638 , \20632 , \20636 );
or \U$19656 ( \20639 , \20635 , \20637 , \20638 );
and \U$19657 ( \20640 , \20519 , \20639 );
xor \U$19658 ( \20641 , \20519 , \20639 );
xor \U$19659 ( \20642 , \20632 , \20634 );
xor \U$19660 ( \20643 , \20642 , \20636 );
and \U$19661 ( \20644 , \6816 , \10101 );
and \U$19662 ( \20645 , \6444 , \10099 );
nor \U$19663 ( \20646 , \20644 , \20645 );
xnor \U$19664 ( \20647 , \20646 , \9791 );
and \U$19665 ( \20648 , \7168 , \9564 );
and \U$19666 ( \20649 , \6825 , \9562 );
nor \U$19667 ( \20650 , \20648 , \20649 );
xnor \U$19668 ( \20651 , \20650 , \9193 );
and \U$19669 ( \20652 , \20647 , \20651 );
and \U$19670 ( \20653 , \7673 , \9002 );
and \U$19671 ( \20654 , \7370 , \9000 );
nor \U$19672 ( \20655 , \20653 , \20654 );
xnor \U$19673 ( \20656 , \20655 , \8684 );
and \U$19674 ( \20657 , \20651 , \20656 );
and \U$19675 ( \20658 , \20647 , \20656 );
or \U$19676 ( \20659 , \20652 , \20657 , \20658 );
and \U$19677 ( \20660 , \8371 , \8435 );
and \U$19678 ( \20661 , \7845 , \8433 );
nor \U$19679 ( \20662 , \20660 , \20661 );
xnor \U$19680 ( \20663 , \20662 , \8186 );
and \U$19681 ( \20664 , \9041 , \7906 );
and \U$19682 ( \20665 , \8795 , \7904 );
nor \U$19683 ( \20666 , \20664 , \20665 );
xnor \U$19684 ( \20667 , \20666 , \7646 );
and \U$19685 ( \20668 , \20663 , \20667 );
and \U$19686 ( \20669 , \9365 , \7412 );
and \U$19687 ( \20670 , \9046 , \7410 );
nor \U$19688 ( \20671 , \20669 , \20670 );
xnor \U$19689 ( \20672 , \20671 , \7097 );
and \U$19690 ( \20673 , \20667 , \20672 );
and \U$19691 ( \20674 , \20663 , \20672 );
or \U$19692 ( \20675 , \20668 , \20673 , \20674 );
and \U$19693 ( \20676 , \20659 , \20675 );
and \U$19694 ( \20677 , \5916 , \11482 );
and \U$19695 ( \20678 , \5447 , \11479 );
nor \U$19696 ( \20679 , \20677 , \20678 );
xnor \U$19697 ( \20680 , \20679 , \10427 );
and \U$19698 ( \20681 , \6185 , \10669 );
and \U$19699 ( \20682 , \5921 , \10667 );
nor \U$19700 ( \20683 , \20681 , \20682 );
xnor \U$19701 ( \20684 , \20683 , \10430 );
and \U$19702 ( \20685 , \20680 , \20684 );
and \U$19703 ( \20686 , \20684 , \5242 );
and \U$19704 ( \20687 , \20680 , \5242 );
or \U$19705 ( \20688 , \20685 , \20686 , \20687 );
and \U$19706 ( \20689 , \20675 , \20688 );
and \U$19707 ( \20690 , \20659 , \20688 );
or \U$19708 ( \20691 , \20676 , \20689 , \20690 );
and \U$19709 ( \20692 , \10218 , \6903 );
and \U$19710 ( \20693 , \9649 , \6901 );
nor \U$19711 ( \20694 , \20692 , \20693 );
xnor \U$19712 ( \20695 , \20694 , \6563 );
and \U$19713 ( \20696 , \10829 , \6314 );
and \U$19714 ( \20697 , \10226 , \6312 );
nor \U$19715 ( \20698 , \20696 , \20697 );
xnor \U$19716 ( \20699 , \20698 , \6073 );
and \U$19717 ( \20700 , \20695 , \20699 );
and \U$19718 ( \20701 , \11015 , \5848 );
and \U$19719 ( \20702 , \10834 , \5846 );
nor \U$19720 ( \20703 , \20701 , \20702 );
xnor \U$19721 ( \20704 , \20703 , \5660 );
and \U$19722 ( \20705 , \20699 , \20704 );
and \U$19723 ( \20706 , \20695 , \20704 );
or \U$19724 ( \20707 , \20700 , \20705 , \20706 );
xor \U$19725 ( \20708 , \20539 , \20543 );
xor \U$19726 ( \20709 , \20708 , \20548 );
and \U$19727 ( \20710 , \20707 , \20709 );
xor \U$19728 ( \20711 , \20586 , \20590 );
xor \U$19729 ( \20712 , \20711 , \20595 );
and \U$19730 ( \20713 , \20709 , \20712 );
and \U$19731 ( \20714 , \20707 , \20712 );
or \U$19732 ( \20715 , \20710 , \20713 , \20714 );
and \U$19733 ( \20716 , \20691 , \20715 );
xor \U$19734 ( \20717 , \20523 , \20527 );
xor \U$19735 ( \20718 , \20717 , \20532 );
xor \U$19736 ( \20719 , \20556 , \20560 );
xor \U$19737 ( \20720 , \20719 , \20565 );
and \U$19738 ( \20721 , \20718 , \20720 );
and \U$19739 ( \20722 , \20715 , \20721 );
and \U$19740 ( \20723 , \20691 , \20721 );
or \U$19741 ( \20724 , \20716 , \20722 , \20723 );
xor \U$19742 ( \20725 , \20535 , \20551 );
xor \U$19743 ( \20726 , \20725 , \20568 );
xor \U$19744 ( \20727 , \20573 , \20575 );
xor \U$19745 ( \20728 , \20727 , \20578 );
and \U$19746 ( \20729 , \20726 , \20728 );
xor \U$19747 ( \20730 , \20598 , \20600 );
xor \U$19748 ( \20731 , \20730 , \20602 );
and \U$19749 ( \20732 , \20728 , \20731 );
and \U$19750 ( \20733 , \20726 , \20731 );
or \U$19751 ( \20734 , \20729 , \20732 , \20733 );
and \U$19752 ( \20735 , \20724 , \20734 );
xor \U$19753 ( \20736 , \20395 , \20407 );
xor \U$19754 ( \20737 , \20736 , \20424 );
and \U$19755 ( \20738 , \20734 , \20737 );
and \U$19756 ( \20739 , \20724 , \20737 );
or \U$19757 ( \20740 , \20735 , \20738 , \20739 );
xor \U$19758 ( \20741 , \20571 , \20581 );
xor \U$19759 ( \20742 , \20741 , \20605 );
xor \U$19760 ( \20743 , \20610 , \20612 );
xor \U$19761 ( \20744 , \20743 , \20615 );
and \U$19762 ( \20745 , \20742 , \20744 );
and \U$19763 ( \20746 , \20740 , \20745 );
xor \U$19764 ( \20747 , \20427 , \20458 );
xor \U$19765 ( \20748 , \20747 , \20469 );
and \U$19766 ( \20749 , \20745 , \20748 );
and \U$19767 ( \20750 , \20740 , \20748 );
or \U$19768 ( \20751 , \20746 , \20749 , \20750 );
xor \U$19769 ( \20752 , \20624 , \20626 );
xor \U$19770 ( \20753 , \20752 , \20629 );
and \U$19771 ( \20754 , \20751 , \20753 );
and \U$19772 ( \20755 , \20643 , \20754 );
xor \U$19773 ( \20756 , \20643 , \20754 );
xor \U$19774 ( \20757 , \20751 , \20753 );
xor \U$19775 ( \20758 , \20740 , \20745 );
xor \U$19776 ( \20759 , \20758 , \20748 );
xor \U$19777 ( \20760 , \20608 , \20618 );
xor \U$19778 ( \20761 , \20760 , \20621 );
and \U$19779 ( \20762 , \20759 , \20761 );
and \U$19780 ( \20763 , \20757 , \20762 );
xor \U$19781 ( \20764 , \20757 , \20762 );
xor \U$19782 ( \20765 , \20759 , \20761 );
and \U$19783 ( \20766 , \5921 , \11482 );
and \U$19784 ( \20767 , \5916 , \11479 );
nor \U$19785 ( \20768 , \20766 , \20767 );
xnor \U$19786 ( \20769 , \20768 , \10427 );
and \U$19787 ( \20770 , \6444 , \10669 );
and \U$19788 ( \20771 , \6185 , \10667 );
nor \U$19789 ( \20772 , \20770 , \20771 );
xnor \U$19790 ( \20773 , \20772 , \10430 );
and \U$19791 ( \20774 , \20769 , \20773 );
and \U$19792 ( \20775 , \6825 , \10101 );
and \U$19793 ( \20776 , \6816 , \10099 );
nor \U$19794 ( \20777 , \20775 , \20776 );
xnor \U$19795 ( \20778 , \20777 , \9791 );
and \U$19796 ( \20779 , \20773 , \20778 );
and \U$19797 ( \20780 , \20769 , \20778 );
or \U$19798 ( \20781 , \20774 , \20779 , \20780 );
and \U$19799 ( \20782 , \9046 , \7906 );
and \U$19800 ( \20783 , \9041 , \7904 );
nor \U$19801 ( \20784 , \20782 , \20783 );
xnor \U$19802 ( \20785 , \20784 , \7646 );
and \U$19803 ( \20786 , \9649 , \7412 );
and \U$19804 ( \20787 , \9365 , \7410 );
nor \U$19805 ( \20788 , \20786 , \20787 );
xnor \U$19806 ( \20789 , \20788 , \7097 );
and \U$19807 ( \20790 , \20785 , \20789 );
and \U$19808 ( \20791 , \10226 , \6903 );
and \U$19809 ( \20792 , \10218 , \6901 );
nor \U$19810 ( \20793 , \20791 , \20792 );
xnor \U$19811 ( \20794 , \20793 , \6563 );
and \U$19812 ( \20795 , \20789 , \20794 );
and \U$19813 ( \20796 , \20785 , \20794 );
or \U$19814 ( \20797 , \20790 , \20795 , \20796 );
and \U$19815 ( \20798 , \20781 , \20797 );
and \U$19816 ( \20799 , \7370 , \9564 );
and \U$19817 ( \20800 , \7168 , \9562 );
nor \U$19818 ( \20801 , \20799 , \20800 );
xnor \U$19819 ( \20802 , \20801 , \9193 );
and \U$19820 ( \20803 , \7845 , \9002 );
and \U$19821 ( \20804 , \7673 , \9000 );
nor \U$19822 ( \20805 , \20803 , \20804 );
xnor \U$19823 ( \20806 , \20805 , \8684 );
and \U$19824 ( \20807 , \20802 , \20806 );
and \U$19825 ( \20808 , \8795 , \8435 );
and \U$19826 ( \20809 , \8371 , \8433 );
nor \U$19827 ( \20810 , \20808 , \20809 );
xnor \U$19828 ( \20811 , \20810 , \8186 );
and \U$19829 ( \20812 , \20806 , \20811 );
and \U$19830 ( \20813 , \20802 , \20811 );
or \U$19831 ( \20814 , \20807 , \20812 , \20813 );
and \U$19832 ( \20815 , \20797 , \20814 );
and \U$19833 ( \20816 , \20781 , \20814 );
or \U$19834 ( \20817 , \20798 , \20815 , \20816 );
nand \U$19835 ( \20818 , \11635 , \5472 );
xnor \U$19836 ( \20819 , \20818 , \5242 );
xor \U$19837 ( \20820 , \20663 , \20667 );
xor \U$19838 ( \20821 , \20820 , \20672 );
and \U$19839 ( \20822 , \20819 , \20821 );
xor \U$19840 ( \20823 , \20695 , \20699 );
xor \U$19841 ( \20824 , \20823 , \20704 );
and \U$19842 ( \20825 , \20821 , \20824 );
and \U$19843 ( \20826 , \20819 , \20824 );
or \U$19844 ( \20827 , \20822 , \20825 , \20826 );
and \U$19845 ( \20828 , \20817 , \20827 );
xor \U$19846 ( \20829 , \20647 , \20651 );
xor \U$19847 ( \20830 , \20829 , \20656 );
xor \U$19848 ( \20831 , \20680 , \20684 );
xor \U$19849 ( \20832 , \20831 , \5242 );
and \U$19850 ( \20833 , \20830 , \20832 );
and \U$19851 ( \20834 , \20827 , \20833 );
and \U$19852 ( \20835 , \20817 , \20833 );
or \U$19853 ( \20836 , \20828 , \20834 , \20835 );
xor \U$19854 ( \20837 , \20659 , \20675 );
xor \U$19855 ( \20838 , \20837 , \20688 );
xor \U$19856 ( \20839 , \20707 , \20709 );
xor \U$19857 ( \20840 , \20839 , \20712 );
and \U$19858 ( \20841 , \20838 , \20840 );
xor \U$19859 ( \20842 , \20718 , \20720 );
and \U$19860 ( \20843 , \20840 , \20842 );
and \U$19861 ( \20844 , \20838 , \20842 );
or \U$19862 ( \20845 , \20841 , \20843 , \20844 );
and \U$19863 ( \20846 , \20836 , \20845 );
xor \U$19864 ( \20847 , \20726 , \20728 );
xor \U$19865 ( \20848 , \20847 , \20731 );
and \U$19866 ( \20849 , \20845 , \20848 );
and \U$19867 ( \20850 , \20836 , \20848 );
or \U$19868 ( \20851 , \20846 , \20849 , \20850 );
xor \U$19869 ( \20852 , \20724 , \20734 );
xor \U$19870 ( \20853 , \20852 , \20737 );
and \U$19871 ( \20854 , \20851 , \20853 );
xor \U$19872 ( \20855 , \20742 , \20744 );
and \U$19873 ( \20856 , \20853 , \20855 );
and \U$19874 ( \20857 , \20851 , \20855 );
or \U$19875 ( \20858 , \20854 , \20856 , \20857 );
and \U$19876 ( \20859 , \20765 , \20858 );
xor \U$19877 ( \20860 , \20765 , \20858 );
xor \U$19878 ( \20861 , \20851 , \20853 );
xor \U$19879 ( \20862 , \20861 , \20855 );
and \U$19880 ( \20863 , \10829 , \6903 );
and \U$19881 ( \20864 , \10226 , \6901 );
nor \U$19882 ( \20865 , \20863 , \20864 );
xnor \U$19883 ( \20866 , \20865 , \6563 );
and \U$19884 ( \20867 , \11015 , \6314 );
and \U$19885 ( \20868 , \10834 , \6312 );
nor \U$19886 ( \20869 , \20867 , \20868 );
xnor \U$19887 ( \20870 , \20869 , \6073 );
and \U$19888 ( \20871 , \20866 , \20870 );
nand \U$19889 ( \20872 , \11635 , \5846 );
xnor \U$19890 ( \20873 , \20872 , \5660 );
and \U$19891 ( \20874 , \20870 , \20873 );
and \U$19892 ( \20875 , \20866 , \20873 );
or \U$19893 ( \20876 , \20871 , \20874 , \20875 );
and \U$19894 ( \20877 , \10834 , \6314 );
and \U$19895 ( \20878 , \10829 , \6312 );
nor \U$19896 ( \20879 , \20877 , \20878 );
xnor \U$19897 ( \20880 , \20879 , \6073 );
and \U$19898 ( \20881 , \20876 , \20880 );
and \U$19899 ( \20882 , \11635 , \5848 );
and \U$19900 ( \20883 , \11015 , \5846 );
nor \U$19901 ( \20884 , \20882 , \20883 );
xnor \U$19902 ( \20885 , \20884 , \5660 );
and \U$19903 ( \20886 , \20880 , \20885 );
and \U$19904 ( \20887 , \20876 , \20885 );
or \U$19905 ( \20888 , \20881 , \20886 , \20887 );
and \U$19906 ( \20889 , \6185 , \11482 );
and \U$19907 ( \20890 , \5921 , \11479 );
nor \U$19908 ( \20891 , \20889 , \20890 );
xnor \U$19909 ( \20892 , \20891 , \10427 );
and \U$19910 ( \20893 , \6816 , \10669 );
and \U$19911 ( \20894 , \6444 , \10667 );
nor \U$19912 ( \20895 , \20893 , \20894 );
xnor \U$19913 ( \20896 , \20895 , \10430 );
and \U$19914 ( \20897 , \20892 , \20896 );
and \U$19915 ( \20898 , \20896 , \5660 );
and \U$19916 ( \20899 , \20892 , \5660 );
or \U$19917 ( \20900 , \20897 , \20898 , \20899 );
and \U$19918 ( \20901 , \7168 , \10101 );
and \U$19919 ( \20902 , \6825 , \10099 );
nor \U$19920 ( \20903 , \20901 , \20902 );
xnor \U$19921 ( \20904 , \20903 , \9791 );
and \U$19922 ( \20905 , \7673 , \9564 );
and \U$19923 ( \20906 , \7370 , \9562 );
nor \U$19924 ( \20907 , \20905 , \20906 );
xnor \U$19925 ( \20908 , \20907 , \9193 );
and \U$19926 ( \20909 , \20904 , \20908 );
and \U$19927 ( \20910 , \8371 , \9002 );
and \U$19928 ( \20911 , \7845 , \9000 );
nor \U$19929 ( \20912 , \20910 , \20911 );
xnor \U$19930 ( \20913 , \20912 , \8684 );
and \U$19931 ( \20914 , \20908 , \20913 );
and \U$19932 ( \20915 , \20904 , \20913 );
or \U$19933 ( \20916 , \20909 , \20914 , \20915 );
and \U$19934 ( \20917 , \20900 , \20916 );
and \U$19935 ( \20918 , \9041 , \8435 );
and \U$19936 ( \20919 , \8795 , \8433 );
nor \U$19937 ( \20920 , \20918 , \20919 );
xnor \U$19938 ( \20921 , \20920 , \8186 );
and \U$19939 ( \20922 , \9365 , \7906 );
and \U$19940 ( \20923 , \9046 , \7904 );
nor \U$19941 ( \20924 , \20922 , \20923 );
xnor \U$19942 ( \20925 , \20924 , \7646 );
and \U$19943 ( \20926 , \20921 , \20925 );
and \U$19944 ( \20927 , \10218 , \7412 );
and \U$19945 ( \20928 , \9649 , \7410 );
nor \U$19946 ( \20929 , \20927 , \20928 );
xnor \U$19947 ( \20930 , \20929 , \7097 );
and \U$19948 ( \20931 , \20925 , \20930 );
and \U$19949 ( \20932 , \20921 , \20930 );
or \U$19950 ( \20933 , \20926 , \20931 , \20932 );
and \U$19951 ( \20934 , \20916 , \20933 );
and \U$19952 ( \20935 , \20900 , \20933 );
or \U$19953 ( \20936 , \20917 , \20934 , \20935 );
and \U$19954 ( \20937 , \20888 , \20936 );
xor \U$19955 ( \20938 , \20769 , \20773 );
xor \U$19956 ( \20939 , \20938 , \20778 );
xor \U$19957 ( \20940 , \20785 , \20789 );
xor \U$19958 ( \20941 , \20940 , \20794 );
and \U$19959 ( \20942 , \20939 , \20941 );
xor \U$19960 ( \20943 , \20802 , \20806 );
xor \U$19961 ( \20944 , \20943 , \20811 );
and \U$19962 ( \20945 , \20941 , \20944 );
and \U$19963 ( \20946 , \20939 , \20944 );
or \U$19964 ( \20947 , \20942 , \20945 , \20946 );
and \U$19965 ( \20948 , \20936 , \20947 );
and \U$19966 ( \20949 , \20888 , \20947 );
or \U$19967 ( \20950 , \20937 , \20948 , \20949 );
xor \U$19968 ( \20951 , \20781 , \20797 );
xor \U$19969 ( \20952 , \20951 , \20814 );
xor \U$19970 ( \20953 , \20819 , \20821 );
xor \U$19971 ( \20954 , \20953 , \20824 );
and \U$19972 ( \20955 , \20952 , \20954 );
xor \U$19973 ( \20956 , \20830 , \20832 );
and \U$19974 ( \20957 , \20954 , \20956 );
and \U$19975 ( \20958 , \20952 , \20956 );
or \U$19976 ( \20959 , \20955 , \20957 , \20958 );
and \U$19977 ( \20960 , \20950 , \20959 );
xor \U$19978 ( \20961 , \20838 , \20840 );
xor \U$19979 ( \20962 , \20961 , \20842 );
and \U$19980 ( \20963 , \20959 , \20962 );
and \U$19981 ( \20964 , \20950 , \20962 );
or \U$19982 ( \20965 , \20960 , \20963 , \20964 );
xor \U$19983 ( \20966 , \20691 , \20715 );
xor \U$19984 ( \20967 , \20966 , \20721 );
and \U$19985 ( \20968 , \20965 , \20967 );
xor \U$19986 ( \20969 , \20836 , \20845 );
xor \U$19987 ( \20970 , \20969 , \20848 );
and \U$19988 ( \20971 , \20967 , \20970 );
and \U$19989 ( \20972 , \20965 , \20970 );
or \U$19990 ( \20973 , \20968 , \20971 , \20972 );
and \U$19991 ( \20974 , \20862 , \20973 );
xor \U$19992 ( \20975 , \20862 , \20973 );
xor \U$19993 ( \20976 , \20965 , \20967 );
xor \U$19994 ( \20977 , \20976 , \20970 );
and \U$19995 ( \20978 , \9649 , \7906 );
and \U$19996 ( \20979 , \9365 , \7904 );
nor \U$19997 ( \20980 , \20978 , \20979 );
xnor \U$19998 ( \20981 , \20980 , \7646 );
and \U$19999 ( \20982 , \10226 , \7412 );
and \U$20000 ( \20983 , \10218 , \7410 );
nor \U$20001 ( \20984 , \20982 , \20983 );
xnor \U$20002 ( \20985 , \20984 , \7097 );
and \U$20003 ( \20986 , \20981 , \20985 );
and \U$20004 ( \20987 , \10834 , \6903 );
and \U$20005 ( \20988 , \10829 , \6901 );
nor \U$20006 ( \20989 , \20987 , \20988 );
xnor \U$20007 ( \20990 , \20989 , \6563 );
and \U$20008 ( \20991 , \20985 , \20990 );
and \U$20009 ( \20992 , \20981 , \20990 );
or \U$20010 ( \20993 , \20986 , \20991 , \20992 );
and \U$20011 ( \20994 , \6444 , \11482 );
and \U$20012 ( \20995 , \6185 , \11479 );
nor \U$20013 ( \20996 , \20994 , \20995 );
xnor \U$20014 ( \20997 , \20996 , \10427 );
and \U$20015 ( \20998 , \6825 , \10669 );
and \U$20016 ( \20999 , \6816 , \10667 );
nor \U$20017 ( \21000 , \20998 , \20999 );
xnor \U$20018 ( \21001 , \21000 , \10430 );
and \U$20019 ( \21002 , \20997 , \21001 );
and \U$20020 ( \21003 , \7370 , \10101 );
and \U$20021 ( \21004 , \7168 , \10099 );
nor \U$20022 ( \21005 , \21003 , \21004 );
xnor \U$20023 ( \21006 , \21005 , \9791 );
and \U$20024 ( \21007 , \21001 , \21006 );
and \U$20025 ( \21008 , \20997 , \21006 );
or \U$20026 ( \21009 , \21002 , \21007 , \21008 );
and \U$20027 ( \21010 , \20993 , \21009 );
and \U$20028 ( \21011 , \7845 , \9564 );
and \U$20029 ( \21012 , \7673 , \9562 );
nor \U$20030 ( \21013 , \21011 , \21012 );
xnor \U$20031 ( \21014 , \21013 , \9193 );
and \U$20032 ( \21015 , \8795 , \9002 );
and \U$20033 ( \21016 , \8371 , \9000 );
nor \U$20034 ( \21017 , \21015 , \21016 );
xnor \U$20035 ( \21018 , \21017 , \8684 );
and \U$20036 ( \21019 , \21014 , \21018 );
and \U$20037 ( \21020 , \9046 , \8435 );
and \U$20038 ( \21021 , \9041 , \8433 );
nor \U$20039 ( \21022 , \21020 , \21021 );
xnor \U$20040 ( \21023 , \21022 , \8186 );
and \U$20041 ( \21024 , \21018 , \21023 );
and \U$20042 ( \21025 , \21014 , \21023 );
or \U$20043 ( \21026 , \21019 , \21024 , \21025 );
and \U$20044 ( \21027 , \21009 , \21026 );
and \U$20045 ( \21028 , \20993 , \21026 );
or \U$20046 ( \21029 , \21010 , \21027 , \21028 );
xor \U$20047 ( \21030 , \20904 , \20908 );
xor \U$20048 ( \21031 , \21030 , \20913 );
xor \U$20049 ( \21032 , \20866 , \20870 );
xor \U$20050 ( \21033 , \21032 , \20873 );
and \U$20051 ( \21034 , \21031 , \21033 );
xor \U$20052 ( \21035 , \20921 , \20925 );
xor \U$20053 ( \21036 , \21035 , \20930 );
and \U$20054 ( \21037 , \21033 , \21036 );
and \U$20055 ( \21038 , \21031 , \21036 );
or \U$20056 ( \21039 , \21034 , \21037 , \21038 );
and \U$20057 ( \21040 , \21029 , \21039 );
xor \U$20058 ( \21041 , \20939 , \20941 );
xor \U$20059 ( \21042 , \21041 , \20944 );
and \U$20060 ( \21043 , \21039 , \21042 );
and \U$20061 ( \21044 , \21029 , \21042 );
or \U$20062 ( \21045 , \21040 , \21043 , \21044 );
xor \U$20063 ( \21046 , \20888 , \20936 );
xor \U$20064 ( \21047 , \21046 , \20947 );
and \U$20065 ( \21048 , \21045 , \21047 );
xor \U$20066 ( \21049 , \20952 , \20954 );
xor \U$20067 ( \21050 , \21049 , \20956 );
and \U$20068 ( \21051 , \21047 , \21050 );
and \U$20069 ( \21052 , \21045 , \21050 );
or \U$20070 ( \21053 , \21048 , \21051 , \21052 );
xor \U$20071 ( \21054 , \20817 , \20827 );
xor \U$20072 ( \21055 , \21054 , \20833 );
and \U$20073 ( \21056 , \21053 , \21055 );
xor \U$20074 ( \21057 , \20950 , \20959 );
xor \U$20075 ( \21058 , \21057 , \20962 );
and \U$20076 ( \21059 , \21055 , \21058 );
and \U$20077 ( \21060 , \21053 , \21058 );
or \U$20078 ( \21061 , \21056 , \21059 , \21060 );
and \U$20079 ( \21062 , \20977 , \21061 );
xor \U$20080 ( \21063 , \20977 , \21061 );
xor \U$20081 ( \21064 , \21053 , \21055 );
xor \U$20082 ( \21065 , \21064 , \21058 );
and \U$20083 ( \21066 , \6816 , \11482 );
and \U$20084 ( \21067 , \6444 , \11479 );
nor \U$20085 ( \21068 , \21066 , \21067 );
xnor \U$20086 ( \21069 , \21068 , \10427 );
and \U$20087 ( \21070 , \7168 , \10669 );
and \U$20088 ( \21071 , \6825 , \10667 );
nor \U$20089 ( \21072 , \21070 , \21071 );
xnor \U$20090 ( \21073 , \21072 , \10430 );
and \U$20091 ( \21074 , \21069 , \21073 );
and \U$20092 ( \21075 , \21073 , \6073 );
and \U$20093 ( \21076 , \21069 , \6073 );
or \U$20094 ( \21077 , \21074 , \21075 , \21076 );
and \U$20095 ( \21078 , \9365 , \8435 );
and \U$20096 ( \21079 , \9046 , \8433 );
nor \U$20097 ( \21080 , \21078 , \21079 );
xnor \U$20098 ( \21081 , \21080 , \8186 );
and \U$20099 ( \21082 , \10218 , \7906 );
and \U$20100 ( \21083 , \9649 , \7904 );
nor \U$20101 ( \21084 , \21082 , \21083 );
xnor \U$20102 ( \21085 , \21084 , \7646 );
and \U$20103 ( \21086 , \21081 , \21085 );
and \U$20104 ( \21087 , \10829 , \7412 );
and \U$20105 ( \21088 , \10226 , \7410 );
nor \U$20106 ( \21089 , \21087 , \21088 );
xnor \U$20107 ( \21090 , \21089 , \7097 );
and \U$20108 ( \21091 , \21085 , \21090 );
and \U$20109 ( \21092 , \21081 , \21090 );
or \U$20110 ( \21093 , \21086 , \21091 , \21092 );
and \U$20111 ( \21094 , \21077 , \21093 );
and \U$20112 ( \21095 , \7673 , \10101 );
and \U$20113 ( \21096 , \7370 , \10099 );
nor \U$20114 ( \21097 , \21095 , \21096 );
xnor \U$20115 ( \21098 , \21097 , \9791 );
and \U$20116 ( \21099 , \8371 , \9564 );
and \U$20117 ( \21100 , \7845 , \9562 );
nor \U$20118 ( \21101 , \21099 , \21100 );
xnor \U$20119 ( \21102 , \21101 , \9193 );
and \U$20120 ( \21103 , \21098 , \21102 );
and \U$20121 ( \21104 , \9041 , \9002 );
and \U$20122 ( \21105 , \8795 , \9000 );
nor \U$20123 ( \21106 , \21104 , \21105 );
xnor \U$20124 ( \21107 , \21106 , \8684 );
and \U$20125 ( \21108 , \21102 , \21107 );
and \U$20126 ( \21109 , \21098 , \21107 );
or \U$20127 ( \21110 , \21103 , \21108 , \21109 );
and \U$20128 ( \21111 , \21093 , \21110 );
and \U$20129 ( \21112 , \21077 , \21110 );
or \U$20130 ( \21113 , \21094 , \21111 , \21112 );
and \U$20131 ( \21114 , \11635 , \6314 );
and \U$20132 ( \21115 , \11015 , \6312 );
nor \U$20133 ( \21116 , \21114 , \21115 );
xnor \U$20134 ( \21117 , \21116 , \6073 );
xor \U$20135 ( \21118 , \20981 , \20985 );
xor \U$20136 ( \21119 , \21118 , \20990 );
and \U$20137 ( \21120 , \21117 , \21119 );
xor \U$20138 ( \21121 , \21014 , \21018 );
xor \U$20139 ( \21122 , \21121 , \21023 );
and \U$20140 ( \21123 , \21119 , \21122 );
and \U$20141 ( \21124 , \21117 , \21122 );
or \U$20142 ( \21125 , \21120 , \21123 , \21124 );
and \U$20143 ( \21126 , \21113 , \21125 );
xor \U$20144 ( \21127 , \20892 , \20896 );
xor \U$20145 ( \21128 , \21127 , \5660 );
and \U$20146 ( \21129 , \21125 , \21128 );
and \U$20147 ( \21130 , \21113 , \21128 );
or \U$20148 ( \21131 , \21126 , \21129 , \21130 );
xor \U$20149 ( \21132 , \20993 , \21009 );
xor \U$20150 ( \21133 , \21132 , \21026 );
xor \U$20151 ( \21134 , \21031 , \21033 );
xor \U$20152 ( \21135 , \21134 , \21036 );
and \U$20153 ( \21136 , \21133 , \21135 );
and \U$20154 ( \21137 , \21131 , \21136 );
xor \U$20155 ( \21138 , \20876 , \20880 );
xor \U$20156 ( \21139 , \21138 , \20885 );
and \U$20157 ( \21140 , \21136 , \21139 );
and \U$20158 ( \21141 , \21131 , \21139 );
or \U$20159 ( \21142 , \21137 , \21140 , \21141 );
xor \U$20160 ( \21143 , \20900 , \20916 );
xor \U$20161 ( \21144 , \21143 , \20933 );
xor \U$20162 ( \21145 , \21029 , \21039 );
xor \U$20163 ( \21146 , \21145 , \21042 );
and \U$20164 ( \21147 , \21144 , \21146 );
and \U$20165 ( \21148 , \21142 , \21147 );
xor \U$20166 ( \21149 , \21045 , \21047 );
xor \U$20167 ( \21150 , \21149 , \21050 );
and \U$20168 ( \21151 , \21147 , \21150 );
and \U$20169 ( \21152 , \21142 , \21150 );
or \U$20170 ( \21153 , \21148 , \21151 , \21152 );
and \U$20171 ( \21154 , \21065 , \21153 );
xor \U$20172 ( \21155 , \21065 , \21153 );
xor \U$20173 ( \21156 , \21142 , \21147 );
xor \U$20174 ( \21157 , \21156 , \21150 );
and \U$20175 ( \21158 , \8795 , \9564 );
and \U$20176 ( \21159 , \8371 , \9562 );
nor \U$20177 ( \21160 , \21158 , \21159 );
xnor \U$20178 ( \21161 , \21160 , \9193 );
and \U$20179 ( \21162 , \9046 , \9002 );
and \U$20180 ( \21163 , \9041 , \9000 );
nor \U$20181 ( \21164 , \21162 , \21163 );
xnor \U$20182 ( \21165 , \21164 , \8684 );
and \U$20183 ( \21166 , \21161 , \21165 );
and \U$20184 ( \21167 , \9649 , \8435 );
and \U$20185 ( \21168 , \9365 , \8433 );
nor \U$20186 ( \21169 , \21167 , \21168 );
xnor \U$20187 ( \21170 , \21169 , \8186 );
and \U$20188 ( \21171 , \21165 , \21170 );
and \U$20189 ( \21172 , \21161 , \21170 );
or \U$20190 ( \21173 , \21166 , \21171 , \21172 );
and \U$20191 ( \21174 , \6825 , \11482 );
and \U$20192 ( \21175 , \6816 , \11479 );
nor \U$20193 ( \21176 , \21174 , \21175 );
xnor \U$20194 ( \21177 , \21176 , \10427 );
and \U$20195 ( \21178 , \7370 , \10669 );
and \U$20196 ( \21179 , \7168 , \10667 );
nor \U$20197 ( \21180 , \21178 , \21179 );
xnor \U$20198 ( \21181 , \21180 , \10430 );
and \U$20199 ( \21182 , \21177 , \21181 );
and \U$20200 ( \21183 , \7845 , \10101 );
and \U$20201 ( \21184 , \7673 , \10099 );
nor \U$20202 ( \21185 , \21183 , \21184 );
xnor \U$20203 ( \21186 , \21185 , \9791 );
and \U$20204 ( \21187 , \21181 , \21186 );
and \U$20205 ( \21188 , \21177 , \21186 );
or \U$20206 ( \21189 , \21182 , \21187 , \21188 );
and \U$20207 ( \21190 , \21173 , \21189 );
and \U$20208 ( \21191 , \10226 , \7906 );
and \U$20209 ( \21192 , \10218 , \7904 );
nor \U$20210 ( \21193 , \21191 , \21192 );
xnor \U$20211 ( \21194 , \21193 , \7646 );
and \U$20212 ( \21195 , \10834 , \7412 );
and \U$20213 ( \21196 , \10829 , \7410 );
nor \U$20214 ( \21197 , \21195 , \21196 );
xnor \U$20215 ( \21198 , \21197 , \7097 );
and \U$20216 ( \21199 , \21194 , \21198 );
and \U$20217 ( \21200 , \11635 , \6903 );
and \U$20218 ( \21201 , \11015 , \6901 );
nor \U$20219 ( \21202 , \21200 , \21201 );
xnor \U$20220 ( \21203 , \21202 , \6563 );
and \U$20221 ( \21204 , \21198 , \21203 );
and \U$20222 ( \21205 , \21194 , \21203 );
or \U$20223 ( \21206 , \21199 , \21204 , \21205 );
and \U$20224 ( \21207 , \21189 , \21206 );
and \U$20225 ( \21208 , \21173 , \21206 );
or \U$20226 ( \21209 , \21190 , \21207 , \21208 );
and \U$20227 ( \21210 , \11015 , \6903 );
and \U$20228 ( \21211 , \10834 , \6901 );
nor \U$20229 ( \21212 , \21210 , \21211 );
xnor \U$20230 ( \21213 , \21212 , \6563 );
nand \U$20231 ( \21214 , \11635 , \6312 );
xnor \U$20232 ( \21215 , \21214 , \6073 );
and \U$20233 ( \21216 , \21213 , \21215 );
xor \U$20234 ( \21217 , \21081 , \21085 );
xor \U$20235 ( \21218 , \21217 , \21090 );
and \U$20236 ( \21219 , \21215 , \21218 );
and \U$20237 ( \21220 , \21213 , \21218 );
or \U$20238 ( \21221 , \21216 , \21219 , \21220 );
and \U$20239 ( \21222 , \21209 , \21221 );
xor \U$20240 ( \21223 , \20997 , \21001 );
xor \U$20241 ( \21224 , \21223 , \21006 );
and \U$20242 ( \21225 , \21221 , \21224 );
and \U$20243 ( \21226 , \21209 , \21224 );
or \U$20244 ( \21227 , \21222 , \21225 , \21226 );
xor \U$20245 ( \21228 , \21113 , \21125 );
xor \U$20246 ( \21229 , \21228 , \21128 );
and \U$20247 ( \21230 , \21227 , \21229 );
xor \U$20248 ( \21231 , \21133 , \21135 );
and \U$20249 ( \21232 , \21229 , \21231 );
and \U$20250 ( \21233 , \21227 , \21231 );
or \U$20251 ( \21234 , \21230 , \21232 , \21233 );
xor \U$20252 ( \21235 , \21131 , \21136 );
xor \U$20253 ( \21236 , \21235 , \21139 );
and \U$20254 ( \21237 , \21234 , \21236 );
xor \U$20255 ( \21238 , \21144 , \21146 );
and \U$20256 ( \21239 , \21236 , \21238 );
and \U$20257 ( \21240 , \21234 , \21238 );
or \U$20258 ( \21241 , \21237 , \21239 , \21240 );
and \U$20259 ( \21242 , \21157 , \21241 );
xor \U$20260 ( \21243 , \21157 , \21241 );
xor \U$20261 ( \21244 , \21234 , \21236 );
xor \U$20262 ( \21245 , \21244 , \21238 );
and \U$20263 ( \21246 , \8371 , \10101 );
and \U$20264 ( \21247 , \7845 , \10099 );
nor \U$20265 ( \21248 , \21246 , \21247 );
xnor \U$20266 ( \21249 , \21248 , \9791 );
and \U$20267 ( \21250 , \9041 , \9564 );
and \U$20268 ( \21251 , \8795 , \9562 );
nor \U$20269 ( \21252 , \21250 , \21251 );
xnor \U$20270 ( \21253 , \21252 , \9193 );
and \U$20271 ( \21254 , \21249 , \21253 );
and \U$20272 ( \21255 , \9365 , \9002 );
and \U$20273 ( \21256 , \9046 , \9000 );
nor \U$20274 ( \21257 , \21255 , \21256 );
xnor \U$20275 ( \21258 , \21257 , \8684 );
and \U$20276 ( \21259 , \21253 , \21258 );
and \U$20277 ( \21260 , \21249 , \21258 );
or \U$20278 ( \21261 , \21254 , \21259 , \21260 );
and \U$20279 ( \21262 , \7168 , \11482 );
and \U$20280 ( \21263 , \6825 , \11479 );
nor \U$20281 ( \21264 , \21262 , \21263 );
xnor \U$20282 ( \21265 , \21264 , \10427 );
and \U$20283 ( \21266 , \7673 , \10669 );
and \U$20284 ( \21267 , \7370 , \10667 );
nor \U$20285 ( \21268 , \21266 , \21267 );
xnor \U$20286 ( \21269 , \21268 , \10430 );
and \U$20287 ( \21270 , \21265 , \21269 );
and \U$20288 ( \21271 , \21269 , \6563 );
and \U$20289 ( \21272 , \21265 , \6563 );
or \U$20290 ( \21273 , \21270 , \21271 , \21272 );
and \U$20291 ( \21274 , \21261 , \21273 );
and \U$20292 ( \21275 , \10218 , \8435 );
and \U$20293 ( \21276 , \9649 , \8433 );
nor \U$20294 ( \21277 , \21275 , \21276 );
xnor \U$20295 ( \21278 , \21277 , \8186 );
and \U$20296 ( \21279 , \10829 , \7906 );
and \U$20297 ( \21280 , \10226 , \7904 );
nor \U$20298 ( \21281 , \21279 , \21280 );
xnor \U$20299 ( \21282 , \21281 , \7646 );
and \U$20300 ( \21283 , \21278 , \21282 );
and \U$20301 ( \21284 , \11015 , \7412 );
and \U$20302 ( \21285 , \10834 , \7410 );
nor \U$20303 ( \21286 , \21284 , \21285 );
xnor \U$20304 ( \21287 , \21286 , \7097 );
and \U$20305 ( \21288 , \21282 , \21287 );
and \U$20306 ( \21289 , \21278 , \21287 );
or \U$20307 ( \21290 , \21283 , \21288 , \21289 );
and \U$20308 ( \21291 , \21273 , \21290 );
and \U$20309 ( \21292 , \21261 , \21290 );
or \U$20310 ( \21293 , \21274 , \21291 , \21292 );
xor \U$20311 ( \21294 , \21161 , \21165 );
xor \U$20312 ( \21295 , \21294 , \21170 );
xor \U$20313 ( \21296 , \21177 , \21181 );
xor \U$20314 ( \21297 , \21296 , \21186 );
and \U$20315 ( \21298 , \21295 , \21297 );
xor \U$20316 ( \21299 , \21194 , \21198 );
xor \U$20317 ( \21300 , \21299 , \21203 );
and \U$20318 ( \21301 , \21297 , \21300 );
and \U$20319 ( \21302 , \21295 , \21300 );
or \U$20320 ( \21303 , \21298 , \21301 , \21302 );
and \U$20321 ( \21304 , \21293 , \21303 );
xor \U$20322 ( \21305 , \21098 , \21102 );
xor \U$20323 ( \21306 , \21305 , \21107 );
and \U$20324 ( \21307 , \21303 , \21306 );
and \U$20325 ( \21308 , \21293 , \21306 );
or \U$20326 ( \21309 , \21304 , \21307 , \21308 );
xor \U$20327 ( \21310 , \21069 , \21073 );
xor \U$20328 ( \21311 , \21310 , \6073 );
xor \U$20329 ( \21312 , \21173 , \21189 );
xor \U$20330 ( \21313 , \21312 , \21206 );
and \U$20331 ( \21314 , \21311 , \21313 );
xor \U$20332 ( \21315 , \21213 , \21215 );
xor \U$20333 ( \21316 , \21315 , \21218 );
and \U$20334 ( \21317 , \21313 , \21316 );
and \U$20335 ( \21318 , \21311 , \21316 );
or \U$20336 ( \21319 , \21314 , \21317 , \21318 );
and \U$20337 ( \21320 , \21309 , \21319 );
xor \U$20338 ( \21321 , \21117 , \21119 );
xor \U$20339 ( \21322 , \21321 , \21122 );
and \U$20340 ( \21323 , \21319 , \21322 );
and \U$20341 ( \21324 , \21309 , \21322 );
or \U$20342 ( \21325 , \21320 , \21323 , \21324 );
xor \U$20343 ( \21326 , \21077 , \21093 );
xor \U$20344 ( \21327 , \21326 , \21110 );
xor \U$20345 ( \21328 , \21209 , \21221 );
xor \U$20346 ( \21329 , \21328 , \21224 );
and \U$20347 ( \21330 , \21327 , \21329 );
and \U$20348 ( \21331 , \21325 , \21330 );
xor \U$20349 ( \21332 , \21227 , \21229 );
xor \U$20350 ( \21333 , \21332 , \21231 );
and \U$20351 ( \21334 , \21330 , \21333 );
and \U$20352 ( \21335 , \21325 , \21333 );
or \U$20353 ( \21336 , \21331 , \21334 , \21335 );
and \U$20354 ( \21337 , \21245 , \21336 );
xor \U$20355 ( \21338 , \21245 , \21336 );
xor \U$20356 ( \21339 , \21325 , \21330 );
xor \U$20357 ( \21340 , \21339 , \21333 );
and \U$20358 ( \21341 , \7370 , \11482 );
and \U$20359 ( \21342 , \7168 , \11479 );
nor \U$20360 ( \21343 , \21341 , \21342 );
xnor \U$20361 ( \21344 , \21343 , \10427 );
and \U$20362 ( \21345 , \7845 , \10669 );
and \U$20363 ( \21346 , \7673 , \10667 );
nor \U$20364 ( \21347 , \21345 , \21346 );
xnor \U$20365 ( \21348 , \21347 , \10430 );
and \U$20366 ( \21349 , \21344 , \21348 );
and \U$20367 ( \21350 , \8795 , \10101 );
and \U$20368 ( \21351 , \8371 , \10099 );
nor \U$20369 ( \21352 , \21350 , \21351 );
xnor \U$20370 ( \21353 , \21352 , \9791 );
and \U$20371 ( \21354 , \21348 , \21353 );
and \U$20372 ( \21355 , \21344 , \21353 );
or \U$20373 ( \21356 , \21349 , \21354 , \21355 );
and \U$20374 ( \21357 , \9046 , \9564 );
and \U$20375 ( \21358 , \9041 , \9562 );
nor \U$20376 ( \21359 , \21357 , \21358 );
xnor \U$20377 ( \21360 , \21359 , \9193 );
and \U$20378 ( \21361 , \9649 , \9002 );
and \U$20379 ( \21362 , \9365 , \9000 );
nor \U$20380 ( \21363 , \21361 , \21362 );
xnor \U$20381 ( \21364 , \21363 , \8684 );
and \U$20382 ( \21365 , \21360 , \21364 );
and \U$20383 ( \21366 , \10226 , \8435 );
and \U$20384 ( \21367 , \10218 , \8433 );
nor \U$20385 ( \21368 , \21366 , \21367 );
xnor \U$20386 ( \21369 , \21368 , \8186 );
and \U$20387 ( \21370 , \21364 , \21369 );
and \U$20388 ( \21371 , \21360 , \21369 );
or \U$20389 ( \21372 , \21365 , \21370 , \21371 );
and \U$20390 ( \21373 , \21356 , \21372 );
and \U$20391 ( \21374 , \10834 , \7906 );
and \U$20392 ( \21375 , \10829 , \7904 );
nor \U$20393 ( \21376 , \21374 , \21375 );
xnor \U$20394 ( \21377 , \21376 , \7646 );
and \U$20395 ( \21378 , \11635 , \7412 );
and \U$20396 ( \21379 , \11015 , \7410 );
nor \U$20397 ( \21380 , \21378 , \21379 );
xnor \U$20398 ( \21381 , \21380 , \7097 );
and \U$20399 ( \21382 , \21377 , \21381 );
and \U$20400 ( \21383 , \21372 , \21382 );
and \U$20401 ( \21384 , \21356 , \21382 );
or \U$20402 ( \21385 , \21373 , \21383 , \21384 );
nand \U$20403 ( \21386 , \11635 , \6901 );
xnor \U$20404 ( \21387 , \21386 , \6563 );
xor \U$20405 ( \21388 , \21249 , \21253 );
xor \U$20406 ( \21389 , \21388 , \21258 );
and \U$20407 ( \21390 , \21387 , \21389 );
xor \U$20408 ( \21391 , \21278 , \21282 );
xor \U$20409 ( \21392 , \21391 , \21287 );
and \U$20410 ( \21393 , \21389 , \21392 );
and \U$20411 ( \21394 , \21387 , \21392 );
or \U$20412 ( \21395 , \21390 , \21393 , \21394 );
and \U$20413 ( \21396 , \21385 , \21395 );
xor \U$20414 ( \21397 , \21295 , \21297 );
xor \U$20415 ( \21398 , \21397 , \21300 );
and \U$20416 ( \21399 , \21395 , \21398 );
and \U$20417 ( \21400 , \21385 , \21398 );
or \U$20418 ( \21401 , \21396 , \21399 , \21400 );
xor \U$20419 ( \21402 , \21293 , \21303 );
xor \U$20420 ( \21403 , \21402 , \21306 );
and \U$20421 ( \21404 , \21401 , \21403 );
xor \U$20422 ( \21405 , \21311 , \21313 );
xor \U$20423 ( \21406 , \21405 , \21316 );
and \U$20424 ( \21407 , \21403 , \21406 );
and \U$20425 ( \21408 , \21401 , \21406 );
or \U$20426 ( \21409 , \21404 , \21407 , \21408 );
xor \U$20427 ( \21410 , \21309 , \21319 );
xor \U$20428 ( \21411 , \21410 , \21322 );
and \U$20429 ( \21412 , \21409 , \21411 );
xor \U$20430 ( \21413 , \21327 , \21329 );
and \U$20431 ( \21414 , \21411 , \21413 );
and \U$20432 ( \21415 , \21409 , \21413 );
or \U$20433 ( \21416 , \21412 , \21414 , \21415 );
and \U$20434 ( \21417 , \21340 , \21416 );
xor \U$20435 ( \21418 , \21340 , \21416 );
xor \U$20436 ( \21419 , \21409 , \21411 );
xor \U$20437 ( \21420 , \21419 , \21413 );
and \U$20438 ( \21421 , \10829 , \8435 );
and \U$20439 ( \21422 , \10226 , \8433 );
nor \U$20440 ( \21423 , \21421 , \21422 );
xnor \U$20441 ( \21424 , \21423 , \8186 );
and \U$20442 ( \21425 , \11015 , \7906 );
and \U$20443 ( \21426 , \10834 , \7904 );
nor \U$20444 ( \21427 , \21425 , \21426 );
xnor \U$20445 ( \21428 , \21427 , \7646 );
and \U$20446 ( \21429 , \21424 , \21428 );
nand \U$20447 ( \21430 , \11635 , \7410 );
xnor \U$20448 ( \21431 , \21430 , \7097 );
and \U$20449 ( \21432 , \21428 , \21431 );
and \U$20450 ( \21433 , \21424 , \21431 );
or \U$20451 ( \21434 , \21429 , \21432 , \21433 );
and \U$20452 ( \21435 , \7673 , \11482 );
and \U$20453 ( \21436 , \7370 , \11479 );
nor \U$20454 ( \21437 , \21435 , \21436 );
xnor \U$20455 ( \21438 , \21437 , \10427 );
and \U$20456 ( \21439 , \8371 , \10669 );
and \U$20457 ( \21440 , \7845 , \10667 );
nor \U$20458 ( \21441 , \21439 , \21440 );
xnor \U$20459 ( \21442 , \21441 , \10430 );
and \U$20460 ( \21443 , \21438 , \21442 );
and \U$20461 ( \21444 , \21442 , \7097 );
and \U$20462 ( \21445 , \21438 , \7097 );
or \U$20463 ( \21446 , \21443 , \21444 , \21445 );
and \U$20464 ( \21447 , \21434 , \21446 );
and \U$20465 ( \21448 , \9041 , \10101 );
and \U$20466 ( \21449 , \8795 , \10099 );
nor \U$20467 ( \21450 , \21448 , \21449 );
xnor \U$20468 ( \21451 , \21450 , \9791 );
and \U$20469 ( \21452 , \9365 , \9564 );
and \U$20470 ( \21453 , \9046 , \9562 );
nor \U$20471 ( \21454 , \21452 , \21453 );
xnor \U$20472 ( \21455 , \21454 , \9193 );
and \U$20473 ( \21456 , \21451 , \21455 );
and \U$20474 ( \21457 , \10218 , \9002 );
and \U$20475 ( \21458 , \9649 , \9000 );
nor \U$20476 ( \21459 , \21457 , \21458 );
xnor \U$20477 ( \21460 , \21459 , \8684 );
and \U$20478 ( \21461 , \21455 , \21460 );
and \U$20479 ( \21462 , \21451 , \21460 );
or \U$20480 ( \21463 , \21456 , \21461 , \21462 );
and \U$20481 ( \21464 , \21446 , \21463 );
and \U$20482 ( \21465 , \21434 , \21463 );
or \U$20483 ( \21466 , \21447 , \21464 , \21465 );
xor \U$20484 ( \21467 , \21344 , \21348 );
xor \U$20485 ( \21468 , \21467 , \21353 );
xor \U$20486 ( \21469 , \21360 , \21364 );
xor \U$20487 ( \21470 , \21469 , \21369 );
and \U$20488 ( \21471 , \21468 , \21470 );
xor \U$20489 ( \21472 , \21377 , \21381 );
and \U$20490 ( \21473 , \21470 , \21472 );
and \U$20491 ( \21474 , \21468 , \21472 );
or \U$20492 ( \21475 , \21471 , \21473 , \21474 );
and \U$20493 ( \21476 , \21466 , \21475 );
xor \U$20494 ( \21477 , \21265 , \21269 );
xor \U$20495 ( \21478 , \21477 , \6563 );
and \U$20496 ( \21479 , \21475 , \21478 );
and \U$20497 ( \21480 , \21466 , \21478 );
or \U$20498 ( \21481 , \21476 , \21479 , \21480 );
xor \U$20499 ( \21482 , \21356 , \21372 );
xor \U$20500 ( \21483 , \21482 , \21382 );
xor \U$20501 ( \21484 , \21387 , \21389 );
xor \U$20502 ( \21485 , \21484 , \21392 );
and \U$20503 ( \21486 , \21483 , \21485 );
and \U$20504 ( \21487 , \21481 , \21486 );
xor \U$20505 ( \21488 , \21261 , \21273 );
xor \U$20506 ( \21489 , \21488 , \21290 );
and \U$20507 ( \21490 , \21486 , \21489 );
and \U$20508 ( \21491 , \21481 , \21489 );
or \U$20509 ( \21492 , \21487 , \21490 , \21491 );
xor \U$20510 ( \21493 , \21401 , \21403 );
xor \U$20511 ( \21494 , \21493 , \21406 );
and \U$20512 ( \21495 , \21492 , \21494 );
and \U$20513 ( \21496 , \21420 , \21495 );
xor \U$20514 ( \21497 , \21420 , \21495 );
xor \U$20515 ( \21498 , \21492 , \21494 );
xor \U$20516 ( \21499 , \21481 , \21486 );
xor \U$20517 ( \21500 , \21499 , \21489 );
xor \U$20518 ( \21501 , \21385 , \21395 );
xor \U$20519 ( \21502 , \21501 , \21398 );
and \U$20520 ( \21503 , \21500 , \21502 );
and \U$20521 ( \21504 , \21498 , \21503 );
xor \U$20522 ( \21505 , \21498 , \21503 );
xor \U$20523 ( \21506 , \21500 , \21502 );
and \U$20524 ( \21507 , \7845 , \11482 );
and \U$20525 ( \21508 , \7673 , \11479 );
nor \U$20526 ( \21509 , \21507 , \21508 );
xnor \U$20527 ( \21510 , \21509 , \10427 );
and \U$20528 ( \21511 , \8795 , \10669 );
and \U$20529 ( \21512 , \8371 , \10667 );
nor \U$20530 ( \21513 , \21511 , \21512 );
xnor \U$20531 ( \21514 , \21513 , \10430 );
and \U$20532 ( \21515 , \21510 , \21514 );
and \U$20533 ( \21516 , \9046 , \10101 );
and \U$20534 ( \21517 , \9041 , \10099 );
nor \U$20535 ( \21518 , \21516 , \21517 );
xnor \U$20536 ( \21519 , \21518 , \9791 );
and \U$20537 ( \21520 , \21514 , \21519 );
and \U$20538 ( \21521 , \21510 , \21519 );
or \U$20539 ( \21522 , \21515 , \21520 , \21521 );
and \U$20540 ( \21523 , \9649 , \9564 );
and \U$20541 ( \21524 , \9365 , \9562 );
nor \U$20542 ( \21525 , \21523 , \21524 );
xnor \U$20543 ( \21526 , \21525 , \9193 );
and \U$20544 ( \21527 , \10226 , \9002 );
and \U$20545 ( \21528 , \10218 , \9000 );
nor \U$20546 ( \21529 , \21527 , \21528 );
xnor \U$20547 ( \21530 , \21529 , \8684 );
and \U$20548 ( \21531 , \21526 , \21530 );
and \U$20549 ( \21532 , \10834 , \8435 );
and \U$20550 ( \21533 , \10829 , \8433 );
nor \U$20551 ( \21534 , \21532 , \21533 );
xnor \U$20552 ( \21535 , \21534 , \8186 );
and \U$20553 ( \21536 , \21530 , \21535 );
and \U$20554 ( \21537 , \21526 , \21535 );
or \U$20555 ( \21538 , \21531 , \21536 , \21537 );
and \U$20556 ( \21539 , \21522 , \21538 );
xor \U$20557 ( \21540 , \21424 , \21428 );
xor \U$20558 ( \21541 , \21540 , \21431 );
and \U$20559 ( \21542 , \21538 , \21541 );
and \U$20560 ( \21543 , \21522 , \21541 );
or \U$20561 ( \21544 , \21539 , \21542 , \21543 );
xor \U$20562 ( \21545 , \21438 , \21442 );
xor \U$20563 ( \21546 , \21545 , \7097 );
xor \U$20564 ( \21547 , \21451 , \21455 );
xor \U$20565 ( \21548 , \21547 , \21460 );
and \U$20566 ( \21549 , \21546 , \21548 );
and \U$20567 ( \21550 , \21544 , \21549 );
xor \U$20568 ( \21551 , \21468 , \21470 );
xor \U$20569 ( \21552 , \21551 , \21472 );
and \U$20570 ( \21553 , \21549 , \21552 );
and \U$20571 ( \21554 , \21544 , \21552 );
or \U$20572 ( \21555 , \21550 , \21553 , \21554 );
xor \U$20573 ( \21556 , \21466 , \21475 );
xor \U$20574 ( \21557 , \21556 , \21478 );
and \U$20575 ( \21558 , \21555 , \21557 );
xor \U$20576 ( \21559 , \21483 , \21485 );
and \U$20577 ( \21560 , \21557 , \21559 );
and \U$20578 ( \21561 , \21555 , \21559 );
or \U$20579 ( \21562 , \21558 , \21560 , \21561 );
and \U$20580 ( \21563 , \21506 , \21562 );
xor \U$20581 ( \21564 , \21506 , \21562 );
xor \U$20582 ( \21565 , \21555 , \21557 );
xor \U$20583 ( \21566 , \21565 , \21559 );
and \U$20584 ( \21567 , \8371 , \11482 );
and \U$20585 ( \21568 , \7845 , \11479 );
nor \U$20586 ( \21569 , \21567 , \21568 );
xnor \U$20587 ( \21570 , \21569 , \10427 );
and \U$20588 ( \21571 , \9041 , \10669 );
and \U$20589 ( \21572 , \8795 , \10667 );
nor \U$20590 ( \21573 , \21571 , \21572 );
xnor \U$20591 ( \21574 , \21573 , \10430 );
and \U$20592 ( \21575 , \21570 , \21574 );
and \U$20593 ( \21576 , \21574 , \7646 );
and \U$20594 ( \21577 , \21570 , \7646 );
or \U$20595 ( \21578 , \21575 , \21576 , \21577 );
and \U$20596 ( \21579 , \9365 , \10101 );
and \U$20597 ( \21580 , \9046 , \10099 );
nor \U$20598 ( \21581 , \21579 , \21580 );
xnor \U$20599 ( \21582 , \21581 , \9791 );
and \U$20600 ( \21583 , \10218 , \9564 );
and \U$20601 ( \21584 , \9649 , \9562 );
nor \U$20602 ( \21585 , \21583 , \21584 );
xnor \U$20603 ( \21586 , \21585 , \9193 );
and \U$20604 ( \21587 , \21582 , \21586 );
and \U$20605 ( \21588 , \10829 , \9002 );
and \U$20606 ( \21589 , \10226 , \9000 );
nor \U$20607 ( \21590 , \21588 , \21589 );
xnor \U$20608 ( \21591 , \21590 , \8684 );
and \U$20609 ( \21592 , \21586 , \21591 );
and \U$20610 ( \21593 , \21582 , \21591 );
or \U$20611 ( \21594 , \21587 , \21592 , \21593 );
and \U$20612 ( \21595 , \21578 , \21594 );
and \U$20613 ( \21596 , \11635 , \7906 );
and \U$20614 ( \21597 , \11015 , \7904 );
nor \U$20615 ( \21598 , \21596 , \21597 );
xnor \U$20616 ( \21599 , \21598 , \7646 );
and \U$20617 ( \21600 , \21594 , \21599 );
and \U$20618 ( \21601 , \21578 , \21599 );
or \U$20619 ( \21602 , \21595 , \21600 , \21601 );
xor \U$20620 ( \21603 , \21522 , \21538 );
xor \U$20621 ( \21604 , \21603 , \21541 );
and \U$20622 ( \21605 , \21602 , \21604 );
xor \U$20623 ( \21606 , \21546 , \21548 );
and \U$20624 ( \21607 , \21604 , \21606 );
and \U$20625 ( \21608 , \21602 , \21606 );
or \U$20626 ( \21609 , \21605 , \21607 , \21608 );
xor \U$20627 ( \21610 , \21434 , \21446 );
xor \U$20628 ( \21611 , \21610 , \21463 );
and \U$20629 ( \21612 , \21609 , \21611 );
xor \U$20630 ( \21613 , \21544 , \21549 );
xor \U$20631 ( \21614 , \21613 , \21552 );
and \U$20632 ( \21615 , \21611 , \21614 );
and \U$20633 ( \21616 , \21609 , \21614 );
or \U$20634 ( \21617 , \21612 , \21615 , \21616 );
and \U$20635 ( \21618 , \21566 , \21617 );
xor \U$20636 ( \21619 , \21566 , \21617 );
xor \U$20637 ( \21620 , \21609 , \21611 );
xor \U$20638 ( \21621 , \21620 , \21614 );
and \U$20639 ( \21622 , \10226 , \9564 );
and \U$20640 ( \21623 , \10218 , \9562 );
nor \U$20641 ( \21624 , \21622 , \21623 );
xnor \U$20642 ( \21625 , \21624 , \9193 );
and \U$20643 ( \21626 , \10834 , \9002 );
and \U$20644 ( \21627 , \10829 , \9000 );
nor \U$20645 ( \21628 , \21626 , \21627 );
xnor \U$20646 ( \21629 , \21628 , \8684 );
and \U$20647 ( \21630 , \21625 , \21629 );
and \U$20648 ( \21631 , \11635 , \8435 );
and \U$20649 ( \21632 , \11015 , \8433 );
nor \U$20650 ( \21633 , \21631 , \21632 );
xnor \U$20651 ( \21634 , \21633 , \8186 );
and \U$20652 ( \21635 , \21629 , \21634 );
and \U$20653 ( \21636 , \21625 , \21634 );
or \U$20654 ( \21637 , \21630 , \21635 , \21636 );
and \U$20655 ( \21638 , \8795 , \11482 );
and \U$20656 ( \21639 , \8371 , \11479 );
nor \U$20657 ( \21640 , \21638 , \21639 );
xnor \U$20658 ( \21641 , \21640 , \10427 );
and \U$20659 ( \21642 , \9046 , \10669 );
and \U$20660 ( \21643 , \9041 , \10667 );
nor \U$20661 ( \21644 , \21642 , \21643 );
xnor \U$20662 ( \21645 , \21644 , \10430 );
and \U$20663 ( \21646 , \21641 , \21645 );
and \U$20664 ( \21647 , \9649 , \10101 );
and \U$20665 ( \21648 , \9365 , \10099 );
nor \U$20666 ( \21649 , \21647 , \21648 );
xnor \U$20667 ( \21650 , \21649 , \9791 );
and \U$20668 ( \21651 , \21645 , \21650 );
and \U$20669 ( \21652 , \21641 , \21650 );
or \U$20670 ( \21653 , \21646 , \21651 , \21652 );
and \U$20671 ( \21654 , \21637 , \21653 );
and \U$20672 ( \21655 , \11015 , \8435 );
and \U$20673 ( \21656 , \10834 , \8433 );
nor \U$20674 ( \21657 , \21655 , \21656 );
xnor \U$20675 ( \21658 , \21657 , \8186 );
and \U$20676 ( \21659 , \21653 , \21658 );
and \U$20677 ( \21660 , \21637 , \21658 );
or \U$20678 ( \21661 , \21654 , \21659 , \21660 );
nand \U$20679 ( \21662 , \11635 , \7904 );
xnor \U$20680 ( \21663 , \21662 , \7646 );
xor \U$20681 ( \21664 , \21570 , \21574 );
xor \U$20682 ( \21665 , \21664 , \7646 );
and \U$20683 ( \21666 , \21663 , \21665 );
xor \U$20684 ( \21667 , \21582 , \21586 );
xor \U$20685 ( \21668 , \21667 , \21591 );
and \U$20686 ( \21669 , \21665 , \21668 );
and \U$20687 ( \21670 , \21663 , \21668 );
or \U$20688 ( \21671 , \21666 , \21669 , \21670 );
and \U$20689 ( \21672 , \21661 , \21671 );
xor \U$20690 ( \21673 , \21526 , \21530 );
xor \U$20691 ( \21674 , \21673 , \21535 );
and \U$20692 ( \21675 , \21671 , \21674 );
and \U$20693 ( \21676 , \21661 , \21674 );
or \U$20694 ( \21677 , \21672 , \21675 , \21676 );
xor \U$20695 ( \21678 , \21510 , \21514 );
xor \U$20696 ( \21679 , \21678 , \21519 );
xor \U$20697 ( \21680 , \21578 , \21594 );
xor \U$20698 ( \21681 , \21680 , \21599 );
and \U$20699 ( \21682 , \21679 , \21681 );
and \U$20700 ( \21683 , \21677 , \21682 );
xor \U$20701 ( \21684 , \21602 , \21604 );
xor \U$20702 ( \21685 , \21684 , \21606 );
and \U$20703 ( \21686 , \21682 , \21685 );
and \U$20704 ( \21687 , \21677 , \21685 );
or \U$20705 ( \21688 , \21683 , \21686 , \21687 );
and \U$20706 ( \21689 , \21621 , \21688 );
xor \U$20707 ( \21690 , \21621 , \21688 );
xor \U$20708 ( \21691 , \21677 , \21682 );
xor \U$20709 ( \21692 , \21691 , \21685 );
and \U$20710 ( \21693 , \10218 , \10101 );
and \U$20711 ( \21694 , \9649 , \10099 );
nor \U$20712 ( \21695 , \21693 , \21694 );
xnor \U$20713 ( \21696 , \21695 , \9791 );
and \U$20714 ( \21697 , \10829 , \9564 );
and \U$20715 ( \21698 , \10226 , \9562 );
nor \U$20716 ( \21699 , \21697 , \21698 );
xnor \U$20717 ( \21700 , \21699 , \9193 );
and \U$20718 ( \21701 , \21696 , \21700 );
and \U$20719 ( \21702 , \11015 , \9002 );
and \U$20720 ( \21703 , \10834 , \9000 );
nor \U$20721 ( \21704 , \21702 , \21703 );
xnor \U$20722 ( \21705 , \21704 , \8684 );
and \U$20723 ( \21706 , \21700 , \21705 );
and \U$20724 ( \21707 , \21696 , \21705 );
or \U$20725 ( \21708 , \21701 , \21706 , \21707 );
and \U$20726 ( \21709 , \9041 , \11482 );
and \U$20727 ( \21710 , \8795 , \11479 );
nor \U$20728 ( \21711 , \21709 , \21710 );
xnor \U$20729 ( \21712 , \21711 , \10427 );
and \U$20730 ( \21713 , \9365 , \10669 );
and \U$20731 ( \21714 , \9046 , \10667 );
nor \U$20732 ( \21715 , \21713 , \21714 );
xnor \U$20733 ( \21716 , \21715 , \10430 );
and \U$20734 ( \21717 , \21712 , \21716 );
and \U$20735 ( \21718 , \21716 , \8186 );
and \U$20736 ( \21719 , \21712 , \8186 );
or \U$20737 ( \21720 , \21717 , \21718 , \21719 );
and \U$20738 ( \21721 , \21708 , \21720 );
xor \U$20739 ( \21722 , \21625 , \21629 );
xor \U$20740 ( \21723 , \21722 , \21634 );
and \U$20741 ( \21724 , \21720 , \21723 );
and \U$20742 ( \21725 , \21708 , \21723 );
or \U$20743 ( \21726 , \21721 , \21724 , \21725 );
xor \U$20744 ( \21727 , \21637 , \21653 );
xor \U$20745 ( \21728 , \21727 , \21658 );
and \U$20746 ( \21729 , \21726 , \21728 );
xor \U$20747 ( \21730 , \21663 , \21665 );
xor \U$20748 ( \21731 , \21730 , \21668 );
and \U$20749 ( \21732 , \21728 , \21731 );
and \U$20750 ( \21733 , \21726 , \21731 );
or \U$20751 ( \21734 , \21729 , \21732 , \21733 );
xor \U$20752 ( \21735 , \21661 , \21671 );
xor \U$20753 ( \21736 , \21735 , \21674 );
and \U$20754 ( \21737 , \21734 , \21736 );
xor \U$20755 ( \21738 , \21679 , \21681 );
and \U$20756 ( \21739 , \21736 , \21738 );
and \U$20757 ( \21740 , \21734 , \21738 );
or \U$20758 ( \21741 , \21737 , \21739 , \21740 );
and \U$20759 ( \21742 , \21692 , \21741 );
xor \U$20760 ( \21743 , \21692 , \21741 );
xor \U$20761 ( \21744 , \21734 , \21736 );
xor \U$20762 ( \21745 , \21744 , \21738 );
and \U$20763 ( \21746 , \9046 , \11482 );
and \U$20764 ( \21747 , \9041 , \11479 );
nor \U$20765 ( \21748 , \21746 , \21747 );
xnor \U$20766 ( \21749 , \21748 , \10427 );
and \U$20767 ( \21750 , \9649 , \10669 );
and \U$20768 ( \21751 , \9365 , \10667 );
nor \U$20769 ( \21752 , \21750 , \21751 );
xnor \U$20770 ( \21753 , \21752 , \10430 );
and \U$20771 ( \21754 , \21749 , \21753 );
and \U$20772 ( \21755 , \10226 , \10101 );
and \U$20773 ( \21756 , \10218 , \10099 );
nor \U$20774 ( \21757 , \21755 , \21756 );
xnor \U$20775 ( \21758 , \21757 , \9791 );
and \U$20776 ( \21759 , \21753 , \21758 );
and \U$20777 ( \21760 , \21749 , \21758 );
or \U$20778 ( \21761 , \21754 , \21759 , \21760 );
nand \U$20779 ( \21762 , \11635 , \8433 );
xnor \U$20780 ( \21763 , \21762 , \8186 );
and \U$20781 ( \21764 , \21761 , \21763 );
xor \U$20782 ( \21765 , \21696 , \21700 );
xor \U$20783 ( \21766 , \21765 , \21705 );
and \U$20784 ( \21767 , \21763 , \21766 );
and \U$20785 ( \21768 , \21761 , \21766 );
or \U$20786 ( \21769 , \21764 , \21767 , \21768 );
xor \U$20787 ( \21770 , \21641 , \21645 );
xor \U$20788 ( \21771 , \21770 , \21650 );
and \U$20789 ( \21772 , \21769 , \21771 );
xor \U$20790 ( \21773 , \21708 , \21720 );
xor \U$20791 ( \21774 , \21773 , \21723 );
and \U$20792 ( \21775 , \21771 , \21774 );
and \U$20793 ( \21776 , \21769 , \21774 );
or \U$20794 ( \21777 , \21772 , \21775 , \21776 );
xor \U$20795 ( \21778 , \21726 , \21728 );
xor \U$20796 ( \21779 , \21778 , \21731 );
and \U$20797 ( \21780 , \21777 , \21779 );
and \U$20798 ( \21781 , \21745 , \21780 );
xor \U$20799 ( \21782 , \21745 , \21780 );
xor \U$20800 ( \21783 , \21777 , \21779 );
and \U$20801 ( \21784 , \10829 , \10101 );
and \U$20802 ( \21785 , \10226 , \10099 );
nor \U$20803 ( \21786 , \21784 , \21785 );
xnor \U$20804 ( \21787 , \21786 , \9791 );
and \U$20805 ( \21788 , \11015 , \9564 );
and \U$20806 ( \21789 , \10834 , \9562 );
nor \U$20807 ( \21790 , \21788 , \21789 );
xnor \U$20808 ( \21791 , \21790 , \9193 );
and \U$20809 ( \21792 , \21787 , \21791 );
nand \U$20810 ( \21793 , \11635 , \9000 );
xnor \U$20811 ( \21794 , \21793 , \8684 );
and \U$20812 ( \21795 , \21791 , \21794 );
and \U$20813 ( \21796 , \21787 , \21794 );
or \U$20814 ( \21797 , \21792 , \21795 , \21796 );
and \U$20815 ( \21798 , \9365 , \11482 );
and \U$20816 ( \21799 , \9046 , \11479 );
nor \U$20817 ( \21800 , \21798 , \21799 );
xnor \U$20818 ( \21801 , \21800 , \10427 );
and \U$20819 ( \21802 , \10218 , \10669 );
and \U$20820 ( \21803 , \9649 , \10667 );
nor \U$20821 ( \21804 , \21802 , \21803 );
xnor \U$20822 ( \21805 , \21804 , \10430 );
and \U$20823 ( \21806 , \21801 , \21805 );
and \U$20824 ( \21807 , \21805 , \8684 );
and \U$20825 ( \21808 , \21801 , \8684 );
or \U$20826 ( \21809 , \21806 , \21807 , \21808 );
and \U$20827 ( \21810 , \21797 , \21809 );
and \U$20828 ( \21811 , \10834 , \9564 );
and \U$20829 ( \21812 , \10829 , \9562 );
nor \U$20830 ( \21813 , \21811 , \21812 );
xnor \U$20831 ( \21814 , \21813 , \9193 );
and \U$20832 ( \21815 , \21809 , \21814 );
and \U$20833 ( \21816 , \21797 , \21814 );
or \U$20834 ( \21817 , \21810 , \21815 , \21816 );
and \U$20835 ( \21818 , \11635 , \9002 );
and \U$20836 ( \21819 , \11015 , \9000 );
nor \U$20837 ( \21820 , \21818 , \21819 );
xnor \U$20838 ( \21821 , \21820 , \8684 );
xor \U$20839 ( \21822 , \21749 , \21753 );
xor \U$20840 ( \21823 , \21822 , \21758 );
and \U$20841 ( \21824 , \21821 , \21823 );
and \U$20842 ( \21825 , \21817 , \21824 );
xor \U$20843 ( \21826 , \21712 , \21716 );
xor \U$20844 ( \21827 , \21826 , \8186 );
and \U$20845 ( \21828 , \21824 , \21827 );
and \U$20846 ( \21829 , \21817 , \21827 );
or \U$20847 ( \21830 , \21825 , \21828 , \21829 );
xor \U$20848 ( \21831 , \21769 , \21771 );
xor \U$20849 ( \21832 , \21831 , \21774 );
and \U$20850 ( \21833 , \21830 , \21832 );
and \U$20851 ( \21834 , \21783 , \21833 );
xor \U$20852 ( \21835 , \21783 , \21833 );
xor \U$20853 ( \21836 , \21830 , \21832 );
xor \U$20854 ( \21837 , \21761 , \21763 );
xor \U$20855 ( \21838 , \21837 , \21766 );
xor \U$20856 ( \21839 , \21817 , \21824 );
xor \U$20857 ( \21840 , \21839 , \21827 );
and \U$20858 ( \21841 , \21838 , \21840 );
and \U$20859 ( \21842 , \21836 , \21841 );
xor \U$20860 ( \21843 , \21836 , \21841 );
xor \U$20861 ( \21844 , \21838 , \21840 );
and \U$20862 ( \21845 , \9649 , \11482 );
and \U$20863 ( \21846 , \9365 , \11479 );
nor \U$20864 ( \21847 , \21845 , \21846 );
xnor \U$20865 ( \21848 , \21847 , \10427 );
and \U$20866 ( \21849 , \10226 , \10669 );
and \U$20867 ( \21850 , \10218 , \10667 );
nor \U$20868 ( \21851 , \21849 , \21850 );
xnor \U$20869 ( \21852 , \21851 , \10430 );
and \U$20870 ( \21853 , \21848 , \21852 );
and \U$20871 ( \21854 , \10834 , \10101 );
and \U$20872 ( \21855 , \10829 , \10099 );
nor \U$20873 ( \21856 , \21854 , \21855 );
xnor \U$20874 ( \21857 , \21856 , \9791 );
and \U$20875 ( \21858 , \21852 , \21857 );
and \U$20876 ( \21859 , \21848 , \21857 );
or \U$20877 ( \21860 , \21853 , \21858 , \21859 );
xor \U$20878 ( \21861 , \21787 , \21791 );
xor \U$20879 ( \21862 , \21861 , \21794 );
and \U$20880 ( \21863 , \21860 , \21862 );
xor \U$20881 ( \21864 , \21801 , \21805 );
xor \U$20882 ( \21865 , \21864 , \8684 );
and \U$20883 ( \21866 , \21862 , \21865 );
and \U$20884 ( \21867 , \21860 , \21865 );
or \U$20885 ( \21868 , \21863 , \21866 , \21867 );
xor \U$20886 ( \21869 , \21797 , \21809 );
xor \U$20887 ( \21870 , \21869 , \21814 );
and \U$20888 ( \21871 , \21868 , \21870 );
xor \U$20889 ( \21872 , \21821 , \21823 );
and \U$20890 ( \21873 , \21870 , \21872 );
and \U$20891 ( \21874 , \21868 , \21872 );
or \U$20892 ( \21875 , \21871 , \21873 , \21874 );
and \U$20893 ( \21876 , \21844 , \21875 );
xor \U$20894 ( \21877 , \21844 , \21875 );
xor \U$20895 ( \21878 , \21868 , \21870 );
xor \U$20896 ( \21879 , \21878 , \21872 );
and \U$20897 ( \21880 , \10218 , \11482 );
and \U$20898 ( \21881 , \9649 , \11479 );
nor \U$20899 ( \21882 , \21880 , \21881 );
xnor \U$20900 ( \21883 , \21882 , \10427 );
and \U$20901 ( \21884 , \10829 , \10669 );
and \U$20902 ( \21885 , \10226 , \10667 );
nor \U$20903 ( \21886 , \21884 , \21885 );
xnor \U$20904 ( \21887 , \21886 , \10430 );
and \U$20905 ( \21888 , \21883 , \21887 );
and \U$20906 ( \21889 , \21887 , \9193 );
and \U$20907 ( \21890 , \21883 , \9193 );
or \U$20908 ( \21891 , \21888 , \21889 , \21890 );
and \U$20909 ( \21892 , \11015 , \10101 );
and \U$20910 ( \21893 , \10834 , \10099 );
nor \U$20911 ( \21894 , \21892 , \21893 );
xnor \U$20912 ( \21895 , \21894 , \9791 );
nand \U$20913 ( \21896 , \11635 , \9562 );
xnor \U$20914 ( \21897 , \21896 , \9193 );
and \U$20915 ( \21898 , \21895 , \21897 );
and \U$20916 ( \21899 , \21891 , \21898 );
and \U$20917 ( \21900 , \11635 , \9564 );
and \U$20918 ( \21901 , \11015 , \9562 );
nor \U$20919 ( \21902 , \21900 , \21901 );
xnor \U$20920 ( \21903 , \21902 , \9193 );
and \U$20921 ( \21904 , \21898 , \21903 );
and \U$20922 ( \21905 , \21891 , \21903 );
or \U$20923 ( \21906 , \21899 , \21904 , \21905 );
xor \U$20924 ( \21907 , \21860 , \21862 );
xor \U$20925 ( \21908 , \21907 , \21865 );
and \U$20926 ( \21909 , \21906 , \21908 );
and \U$20927 ( \21910 , \21879 , \21909 );
xor \U$20928 ( \21911 , \21879 , \21909 );
xor \U$20929 ( \21912 , \21906 , \21908 );
xor \U$20930 ( \21913 , \21848 , \21852 );
xor \U$20931 ( \21914 , \21913 , \21857 );
xor \U$20932 ( \21915 , \21891 , \21898 );
xor \U$20933 ( \21916 , \21915 , \21903 );
and \U$20934 ( \21917 , \21914 , \21916 );
and \U$20935 ( \21918 , \21912 , \21917 );
xor \U$20936 ( \21919 , \21912 , \21917 );
xor \U$20937 ( \21920 , \21914 , \21916 );
and \U$20938 ( \21921 , \10226 , \11482 );
and \U$20939 ( \21922 , \10218 , \11479 );
nor \U$20940 ( \21923 , \21921 , \21922 );
xnor \U$20941 ( \21924 , \21923 , \10427 );
and \U$20942 ( \21925 , \10834 , \10669 );
and \U$20943 ( \21926 , \10829 , \10667 );
nor \U$20944 ( \21927 , \21925 , \21926 );
xnor \U$20945 ( \21928 , \21927 , \10430 );
and \U$20946 ( \21929 , \21924 , \21928 );
and \U$20947 ( \21930 , \11635 , \10101 );
and \U$20948 ( \21931 , \11015 , \10099 );
nor \U$20949 ( \21932 , \21930 , \21931 );
xnor \U$20950 ( \21933 , \21932 , \9791 );
and \U$20951 ( \21934 , \21928 , \21933 );
and \U$20952 ( \21935 , \21924 , \21933 );
or \U$20953 ( \21936 , \21929 , \21934 , \21935 );
xor \U$20954 ( \21937 , \21883 , \21887 );
xor \U$20955 ( \21938 , \21937 , \9193 );
and \U$20956 ( \21939 , \21936 , \21938 );
xor \U$20957 ( \21940 , \21895 , \21897 );
and \U$20958 ( \21941 , \21938 , \21940 );
and \U$20959 ( \21942 , \21936 , \21940 );
or \U$20960 ( \21943 , \21939 , \21941 , \21942 );
and \U$20961 ( \21944 , \21920 , \21943 );
xor \U$20962 ( \21945 , \21920 , \21943 );
xor \U$20963 ( \21946 , \21936 , \21938 );
xor \U$20964 ( \21947 , \21946 , \21940 );
and \U$20965 ( \21948 , \10829 , \11482 );
and \U$20966 ( \21949 , \10226 , \11479 );
nor \U$20967 ( \21950 , \21948 , \21949 );
xnor \U$20968 ( \21951 , \21950 , \10427 );
and \U$20969 ( \21952 , \11015 , \10669 );
and \U$20970 ( \21953 , \10834 , \10667 );
nor \U$20971 ( \21954 , \21952 , \21953 );
xnor \U$20972 ( \21955 , \21954 , \10430 );
and \U$20973 ( \21956 , \21951 , \21955 );
and \U$20974 ( \21957 , \21955 , \9791 );
and \U$20975 ( \21958 , \21951 , \9791 );
or \U$20976 ( \21959 , \21956 , \21957 , \21958 );
xor \U$20977 ( \21960 , \21924 , \21928 );
xor \U$20978 ( \21961 , \21960 , \21933 );
and \U$20979 ( \21962 , \21959 , \21961 );
and \U$20980 ( \21963 , \21947 , \21962 );
xor \U$20981 ( \21964 , \21947 , \21962 );
xor \U$20982 ( \21965 , \21959 , \21961 );
nand \U$20983 ( \21966 , \11635 , \10099 );
xnor \U$20984 ( \21967 , \21966 , \9791 );
xor \U$20985 ( \21968 , \21951 , \21955 );
xor \U$20986 ( \21969 , \21968 , \9791 );
and \U$20987 ( \21970 , \21967 , \21969 );
and \U$20988 ( \21971 , \21965 , \21970 );
xor \U$20989 ( \21972 , \21965 , \21970 );
xor \U$20990 ( \21973 , \21967 , \21969 );
and \U$20991 ( \21974 , \10834 , \11482 );
and \U$20992 ( \21975 , \10829 , \11479 );
nor \U$20993 ( \21976 , \21974 , \21975 );
xnor \U$20994 ( \21977 , \21976 , \10427 );
and \U$20995 ( \21978 , \11635 , \10669 );
and \U$20996 ( \21979 , \11015 , \10667 );
nor \U$20997 ( \21980 , \21978 , \21979 );
xnor \U$20998 ( \21981 , \21980 , \10430 );
and \U$20999 ( \21982 , \21977 , \21981 );
and \U$21000 ( \21983 , \21973 , \21982 );
xor \U$21001 ( \21984 , \21973 , \21982 );
xor \U$21002 ( \21985 , \21977 , \21981 );
and \U$21003 ( \21986 , \11015 , \11482 );
and \U$21004 ( \21987 , \10834 , \11479 );
nor \U$21005 ( \21988 , \21986 , \21987 );
xnor \U$21006 ( \21989 , \21988 , \10427 );
and \U$21007 ( \21990 , \21989 , \10430 );
and \U$21008 ( \21991 , \21985 , \21990 );
xor \U$21009 ( \21992 , \21985 , \21990 );
nand \U$21010 ( \21993 , \11635 , \10667 );
xnor \U$21011 ( \21994 , \21993 , \10430 );
xor \U$21012 ( \21995 , \21989 , \10430 );
and \U$21013 ( \21996 , \21994 , \21995 );
xor \U$21014 ( \21997 , \21994 , \21995 );
and \U$21015 ( \21998 , \11635 , \11482 );
and \U$21016 ( \21999 , \11015 , \11479 );
nor \U$21017 ( \22000 , \21998 , \21999 );
xnor \U$21018 ( \22001 , \22000 , \10427 );
nand \U$21019 ( \22002 , \11635 , \11479 );
xnor \U$21020 ( \22003 , \22002 , \10427 );
and \U$21021 ( \22004 , \22003 , \10427 );
and \U$21022 ( \22005 , \22001 , \22004 );
and \U$21023 ( \22006 , \21997 , \22005 );
or \U$21024 ( \22007 , \21996 , \22006 );
and \U$21025 ( \22008 , \21992 , \22007 );
or \U$21026 ( \22009 , \21991 , \22008 );
and \U$21027 ( \22010 , \21984 , \22009 );
or \U$21028 ( \22011 , \21983 , \22010 );
and \U$21029 ( \22012 , \21972 , \22011 );
or \U$21030 ( \22013 , \21971 , \22012 );
and \U$21031 ( \22014 , \21964 , \22013 );
or \U$21032 ( \22015 , \21963 , \22014 );
and \U$21033 ( \22016 , \21945 , \22015 );
or \U$21034 ( \22017 , \21944 , \22016 );
and \U$21035 ( \22018 , \21919 , \22017 );
or \U$21036 ( \22019 , \21918 , \22018 );
and \U$21037 ( \22020 , \21911 , \22019 );
or \U$21038 ( \22021 , \21910 , \22020 );
and \U$21039 ( \22022 , \21877 , \22021 );
or \U$21040 ( \22023 , \21876 , \22022 );
and \U$21041 ( \22024 , \21843 , \22023 );
or \U$21042 ( \22025 , \21842 , \22024 );
and \U$21043 ( \22026 , \21835 , \22025 );
or \U$21044 ( \22027 , \21834 , \22026 );
and \U$21045 ( \22028 , \21782 , \22027 );
or \U$21046 ( \22029 , \21781 , \22028 );
and \U$21047 ( \22030 , \21743 , \22029 );
or \U$21048 ( \22031 , \21742 , \22030 );
and \U$21049 ( \22032 , \21690 , \22031 );
or \U$21050 ( \22033 , \21689 , \22032 );
and \U$21051 ( \22034 , \21619 , \22033 );
or \U$21052 ( \22035 , \21618 , \22034 );
and \U$21053 ( \22036 , \21564 , \22035 );
or \U$21054 ( \22037 , \21563 , \22036 );
and \U$21055 ( \22038 , \21505 , \22037 );
or \U$21056 ( \22039 , \21504 , \22038 );
and \U$21057 ( \22040 , \21497 , \22039 );
or \U$21058 ( \22041 , \21496 , \22040 );
and \U$21059 ( \22042 , \21418 , \22041 );
or \U$21060 ( \22043 , \21417 , \22042 );
and \U$21061 ( \22044 , \21338 , \22043 );
or \U$21062 ( \22045 , \21337 , \22044 );
and \U$21063 ( \22046 , \21243 , \22045 );
or \U$21064 ( \22047 , \21242 , \22046 );
and \U$21065 ( \22048 , \21155 , \22047 );
or \U$21066 ( \22049 , \21154 , \22048 );
and \U$21067 ( \22050 , \21063 , \22049 );
or \U$21068 ( \22051 , \21062 , \22050 );
and \U$21069 ( \22052 , \20975 , \22051 );
or \U$21070 ( \22053 , \20974 , \22052 );
and \U$21071 ( \22054 , \20860 , \22053 );
or \U$21072 ( \22055 , \20859 , \22054 );
and \U$21073 ( \22056 , \20764 , \22055 );
or \U$21074 ( \22057 , \20763 , \22056 );
and \U$21075 ( \22058 , \20756 , \22057 );
or \U$21076 ( \22059 , \20755 , \22058 );
and \U$21077 ( \22060 , \20641 , \22059 );
or \U$21078 ( \22061 , \20640 , \22060 );
and \U$21079 ( \22062 , \20517 , \22061 );
or \U$21080 ( \22063 , \20516 , \22062 );
and \U$21081 ( \22064 , \20377 , \22063 );
or \U$21082 ( \22065 , \20376 , \22064 );
and \U$21083 ( \22066 , \20253 , \22065 );
or \U$21084 ( \22067 , \20252 , \22066 );
and \U$21085 ( \22068 , \20109 , \22067 );
or \U$21086 ( \22069 , \20108 , \22068 );
and \U$21087 ( \22070 , \19984 , \22069 );
or \U$21088 ( \22071 , \19983 , \22070 );
and \U$21089 ( \22072 , \19845 , \22071 );
or \U$21090 ( \22073 , \19844 , \22072 );
and \U$21091 ( \22074 , \19681 , \22073 );
or \U$21092 ( \22075 , \19680 , \22074 );
and \U$21093 ( \22076 , \19529 , \22075 );
or \U$21094 ( \22077 , \19528 , \22076 );
and \U$21095 ( \22078 , \19389 , \22077 );
or \U$21096 ( \22079 , \19388 , \22078 );
and \U$21097 ( \22080 , \19221 , \22079 );
or \U$21098 ( \22081 , \19220 , \22080 );
and \U$21099 ( \22082 , \19213 , \22081 );
or \U$21100 ( \22083 , \19212 , \22082 );
and \U$21101 ( \22084 , \19042 , \22083 );
or \U$21102 ( \22085 , \19041 , \22084 );
and \U$21103 ( \22086 , \18866 , \22085 );
or \U$21104 ( \22087 , \18865 , \22086 );
and \U$21105 ( \22088 , \18676 , \22087 );
or \U$21106 ( \22089 , \18675 , \22088 );
and \U$21107 ( \22090 , \18489 , \22089 );
or \U$21108 ( \22091 , \18488 , \22090 );
and \U$21109 ( \22092 , \18304 , \22091 );
or \U$21110 ( \22093 , \18303 , \22092 );
and \U$21111 ( \22094 , \18096 , \22093 );
or \U$21112 ( \22095 , \18095 , \22094 );
and \U$21113 ( \22096 , \17900 , \22095 );
or \U$21114 ( \22097 , \17899 , \22096 );
and \U$21115 ( \22098 , \17703 , \22097 );
or \U$21116 ( \22099 , \17702 , \22098 );
and \U$21117 ( \22100 , \17490 , \22099 );
or \U$21118 ( \22101 , \17489 , \22100 );
and \U$21119 ( \22102 , \17279 , \22101 );
or \U$21120 ( \22103 , \17278 , \22102 );
and \U$21121 ( \22104 , \17048 , \22103 );
or \U$21122 ( \22105 , \17047 , \22104 );
and \U$21123 ( \22106 , \16818 , \22105 );
or \U$21124 ( \22107 , \16817 , \22106 );
and \U$21125 ( \22108 , \16599 , \22107 );
or \U$21126 ( \22109 , \16598 , \22108 );
and \U$21127 ( \22110 , \16374 , \22109 );
or \U$21128 ( \22111 , \16373 , \22110 );
and \U$21129 ( \22112 , \16124 , \22111 );
or \U$21130 ( \22113 , \16123 , \22112 );
and \U$21131 ( \22114 , \15894 , \22113 );
or \U$21132 ( \22115 , \15893 , \22114 );
and \U$21133 ( \22116 , \15648 , \22115 );
or \U$21134 ( \22117 , \15647 , \22116 );
and \U$21135 ( \22118 , \15640 , \22117 );
or \U$21136 ( \22119 , \15639 , \22118 );
and \U$21137 ( \22120 , \15379 , \22119 );
or \U$21138 ( \22121 , \15378 , \22120 );
and \U$21139 ( \22122 , \15117 , \22121 );
or \U$21140 ( \22123 , \15116 , \22122 );
and \U$21141 ( \22124 , \14847 , \22123 );
or \U$21142 ( \22125 , \14846 , \22124 );
and \U$21143 ( \22126 , \14570 , \22125 );
or \U$21144 ( \22127 , \14569 , \22126 );
and \U$21145 ( \22128 , \14294 , \22127 );
or \U$21146 ( \22129 , \14293 , \22128 );
and \U$21147 ( \22130 , \14023 , \22129 );
or \U$21148 ( \22131 , \14022 , \22130 );
and \U$21149 ( \22132 , \13720 , \22131 );
or \U$21150 ( \22133 , \13719 , \22132 );
and \U$21151 ( \22134 , \13441 , \22133 );
or \U$21152 ( \22135 , \13440 , \22134 );
and \U$21153 ( \22136 , \13156 , \22135 );
or \U$21154 ( \22137 , \13155 , \22136 );
and \U$21155 ( \22138 , \12840 , \22137 );
or \U$21156 ( \22139 , \12839 , \22138 );
and \U$21157 ( \22140 , \12540 , \22139 );
or \U$21158 ( \22141 , \12539 , \22140 );
and \U$21159 ( \22142 , \12224 , \22141 );
or \U$21160 ( \22143 , \12223 , \22142 );
and \U$21161 ( \22144 , \11906 , \22143 );
or \U$21162 ( \22145 , \11905 , \22144 );
and \U$21163 ( \22146 , \11595 , \22145 );
or \U$21164 ( \22147 , \11594 , \22146 );
and \U$21165 ( \22148 , \11282 , \22147 );
or \U$21166 ( \22149 , \11281 , \22148 );
and \U$21167 ( \22150 , \10966 , \22149 );
or \U$21168 ( \22151 , \10965 , \22150 );
and \U$21169 ( \22152 , \10648 , \22151 );
or \U$21170 ( \22153 , \10647 , \22152 );
and \U$21171 ( \22154 , \10339 , \22153 );
or \U$21172 ( \22155 , \10338 , \22154 );
and \U$21173 ( \22156 , \10043 , \22155 );
or \U$21174 ( \22157 , \10042 , \22156 );
and \U$21175 ( \22158 , \9742 , \22157 );
or \U$21176 ( \22159 , \9741 , \22158 );
and \U$21177 ( \22160 , \9454 , \22159 );
or \U$21178 ( \22161 , \9453 , \22160 );
and \U$21179 ( \22162 , \9171 , \22161 );
or \U$21180 ( \22163 , \9170 , \22162 );
and \U$21181 ( \22164 , \8876 , \22163 );
or \U$21182 ( \22165 , \8875 , \22164 );
and \U$21183 ( \22166 , \8610 , \22165 );
or \U$21184 ( \22167 , \8609 , \22166 );
and \U$21185 ( \22168 , \8344 , \22167 );
or \U$21186 ( \22169 , \8343 , \22168 );
and \U$21187 ( \22170 , \8083 , \22169 );
or \U$21188 ( \22171 , \8082 , \22170 );
and \U$21189 ( \22172 , \7818 , \22171 );
or \U$21190 ( \22173 , \7817 , \22172 );
and \U$21191 ( \22174 , \7555 , \22173 );
or \U$21192 ( \22175 , \7554 , \22174 );
and \U$21193 ( \22176 , \7298 , \22175 );
or \U$21194 ( \22177 , \7297 , \22176 );
and \U$21195 ( \22178 , \7042 , \22177 );
or \U$21196 ( \22179 , \7041 , \22178 );
and \U$21197 ( \22180 , \6789 , \22179 );
or \U$21198 ( \22181 , \6788 , \22180 );
and \U$21199 ( \22182 , \6541 , \22181 );
or \U$21200 ( \22183 , \6540 , \22182 );
and \U$21201 ( \22184 , \6309 , \22183 );
or \U$21202 ( \22185 , \6308 , \22184 );
and \U$21203 ( \22186 , \6066 , \22185 );
or \U$21204 ( \22187 , \6065 , \22186 );
and \U$21205 ( \22188 , \5637 , \22187 );
or \U$21206 ( \22189 , \5636 , \22188 );
and \U$21207 ( \22190 , \5427 , \22189 );
or \U$21208 ( \22191 , \5426 , \22190 );
and \U$21209 ( \22192 , \5220 , \22191 );
or \U$21210 ( \22193 , \5219 , \22192 );
and \U$21211 ( \22194 , \5018 , \22193 );
or \U$21212 ( \22195 , \5017 , \22194 );
and \U$21213 ( \22196 , \4822 , \22195 );
or \U$21214 ( \22197 , \4821 , \22196 );
and \U$21215 ( \22198 , \4625 , \22197 );
or \U$21216 ( \22199 , \4624 , \22198 );
and \U$21217 ( \22200 , \4448 , \22199 );
or \U$21218 ( \22201 , \4447 , \22200 );
and \U$21219 ( \22202 , \4267 , \22201 );
or \U$21220 ( \22203 , \4266 , \22202 );
and \U$21221 ( \22204 , \4096 , \22203 );
or \U$21222 ( \22205 , \4095 , \22204 );
and \U$21223 ( \22206 , \3921 , \22205 );
or \U$21224 ( \22207 , \3920 , \22206 );
and \U$21225 ( \22208 , \3748 , \22207 );
or \U$21226 ( \22209 , \3747 , \22208 );
and \U$21227 ( \22210 , \3581 , \22209 );
or \U$21228 ( \22211 , \3580 , \22210 );
and \U$21229 ( \22212 , \3415 , \22211 );
or \U$21230 ( \22213 , \3414 , \22212 );
and \U$21231 ( \22214 , \3242 , \22213 );
or \U$21232 ( \22215 , \3241 , \22214 );
and \U$21233 ( \22216 , \2962 , \22215 );
or \U$21234 ( \22217 , \2961 , \22216 );
and \U$21235 ( \22218 , \2825 , \22217 );
or \U$21236 ( \22219 , \2824 , \22218 );
and \U$21237 ( \22220 , \2692 , \22219 );
or \U$21238 ( \22221 , \2691 , \22220 );
and \U$21239 ( \22222 , \2571 , \22221 );
or \U$21240 ( \22223 , \2570 , \22222 );
and \U$21241 ( \22224 , \2448 , \22223 );
or \U$21242 ( \22225 , \2447 , \22224 );
and \U$21243 ( \22226 , \2332 , \22225 );
or \U$21244 ( \22227 , \2331 , \22226 );
and \U$21245 ( \22228 , \2217 , \22227 );
or \U$21246 ( \22229 , \2216 , \22228 );
and \U$21247 ( \22230 , \2103 , \22229 );
or \U$21248 ( \22231 , \2102 , \22230 );
and \U$21249 ( \22232 , \1989 , \22231 );
or \U$21250 ( \22233 , \1988 , \22232 );
and \U$21251 ( \22234 , \1807 , \22233 );
or \U$21252 ( \22235 , \1806 , \22234 );
and \U$21253 ( \22236 , \1728 , \22235 );
or \U$21254 ( \22237 , \1727 , \22236 );
and \U$21255 ( \22238 , \1645 , \22237 );
or \U$21256 ( \22239 , \1644 , \22238 );
and \U$21257 ( \22240 , \1564 , \22239 );
or \U$21258 ( \22241 , \1563 , \22240 );
and \U$21259 ( \22242 , \1489 , \22241 );
or \U$21260 ( \22243 , \1488 , \22242 );
and \U$21261 ( \22244 , \1415 , \22243 );
or \U$21262 ( \22245 , \1414 , \22244 );
and \U$21263 ( \22246 , \1295 , \22245 );
or \U$21264 ( \22247 , \1294 , \22246 );
and \U$21265 ( \22248 , \1242 , \22247 );
or \U$21266 ( \22249 , \1241 , \22248 );
and \U$21267 ( \22250 , \1192 , \22249 );
or \U$21268 ( \22251 , \1191 , \22250 );
and \U$21269 ( \22252 , \1140 , \22251 );
or \U$21270 ( \22253 , \1139 , \22252 );
and \U$21271 ( \22254 , \1070 , \22253 );
or \U$21272 ( \22255 , \1069 , \22254 );
xor \U$21273 ( \22256 , \1023 , \22255 );
buf g5617_GF_PartitionCandidate( \22257_nG5617 , \22256 );
buf \U$21274 ( \22258 , \22257_nG5617 );
xor \U$21276 ( \22259 , \22258 , 1'b0 );
xor \U$21279 ( \22260 , \1070 , \22253 );
buf g561a_GF_PartitionCandidate( \22261_nG561a , \22260 );
buf \U$21280 ( \22262 , \22261_nG561a );
xor \U$21283 ( \22263 , \1140 , \22251 );
buf g561d_GF_PartitionCandidate( \22264_nG561d , \22263 );
buf \U$21284 ( \22265 , \22264_nG561d );
xor \U$21287 ( \22266 , \1192 , \22249 );
buf g5620_GF_PartitionCandidate( \22267_nG5620 , \22266 );
buf \U$21288 ( \22268 , \22267_nG5620 );
xor \U$21291 ( \22269 , \1242 , \22247 );
buf g5623_GF_PartitionCandidate( \22270_nG5623 , \22269 );
buf \U$21292 ( \22271 , \22270_nG5623 );
xor \U$21295 ( \22272 , \1295 , \22245 );
buf g5626_GF_PartitionCandidate( \22273_nG5626 , \22272 );
buf \U$21296 ( \22274 , \22273_nG5626 );
xor \U$21299 ( \22275 , \1415 , \22243 );
buf g5629_GF_PartitionCandidate( \22276_nG5629 , \22275 );
buf \U$21300 ( \22277 , \22276_nG5629 );
xor \U$21303 ( \22278 , \1489 , \22241 );
buf g562c_GF_PartitionCandidate( \22279_nG562c , \22278 );
buf \U$21304 ( \22280 , \22279_nG562c );
xor \U$21307 ( \22281 , \1564 , \22239 );
buf g562f_GF_PartitionCandidate( \22282_nG562f , \22281 );
buf \U$21308 ( \22283 , \22282_nG562f );
xor \U$21311 ( \22284 , \1645 , \22237 );
buf g5632_GF_PartitionCandidate( \22285_nG5632 , \22284 );
buf \U$21312 ( \22286 , \22285_nG5632 );
xor \U$21315 ( \22287 , \1728 , \22235 );
buf g5635_GF_PartitionCandidate( \22288_nG5635 , \22287 );
buf \U$21316 ( \22289 , \22288_nG5635 );
xor \U$21319 ( \22290 , \1807 , \22233 );
buf g5638_GF_PartitionCandidate( \22291_nG5638 , \22290 );
buf \U$21320 ( \22292 , \22291_nG5638 );
xor \U$21323 ( \22293 , \1989 , \22231 );
buf g563b_GF_PartitionCandidate( \22294_nG563b , \22293 );
buf \U$21324 ( \22295 , \22294_nG563b );
xor \U$21327 ( \22296 , \2103 , \22229 );
buf g563e_GF_PartitionCandidate( \22297_nG563e , \22296 );
buf \U$21328 ( \22298 , \22297_nG563e );
xor \U$21331 ( \22299 , \2217 , \22227 );
buf g5641_GF_PartitionCandidate( \22300_nG5641 , \22299 );
buf \U$21332 ( \22301 , \22300_nG5641 );
xor \U$21335 ( \22302 , \2332 , \22225 );
buf g5644_GF_PartitionCandidate( \22303_nG5644 , \22302 );
buf \U$21336 ( \22304 , \22303_nG5644 );
xor \U$21339 ( \22305 , \2448 , \22223 );
buf g5647_GF_PartitionCandidate( \22306_nG5647 , \22305 );
buf \U$21340 ( \22307 , \22306_nG5647 );
xor \U$21343 ( \22308 , \2571 , \22221 );
buf g564a_GF_PartitionCandidate( \22309_nG564a , \22308 );
buf \U$21344 ( \22310 , \22309_nG564a );
xor \U$21347 ( \22311 , \2692 , \22219 );
buf g564d_GF_PartitionCandidate( \22312_nG564d , \22311 );
buf \U$21348 ( \22313 , \22312_nG564d );
xor \U$21351 ( \22314 , \2825 , \22217 );
buf g5650_GF_PartitionCandidate( \22315_nG5650 , \22314 );
buf \U$21352 ( \22316 , \22315_nG5650 );
xor \U$21355 ( \22317 , \2962 , \22215 );
buf g5653_GF_PartitionCandidate( \22318_nG5653 , \22317 );
buf \U$21356 ( \22319 , \22318_nG5653 );
xor \U$21359 ( \22320 , \3242 , \22213 );
buf g5656_GF_PartitionCandidate( \22321_nG5656 , \22320 );
buf \U$21360 ( \22322 , \22321_nG5656 );
xor \U$21363 ( \22323 , \3415 , \22211 );
buf g5659_GF_PartitionCandidate( \22324_nG5659 , \22323 );
buf \U$21364 ( \22325 , \22324_nG5659 );
xor \U$21367 ( \22326 , \3581 , \22209 );
buf g565c_GF_PartitionCandidate( \22327_nG565c , \22326 );
buf \U$21368 ( \22328 , \22327_nG565c );
xor \U$21371 ( \22329 , \3748 , \22207 );
buf g565f_GF_PartitionCandidate( \22330_nG565f , \22329 );
buf \U$21372 ( \22331 , \22330_nG565f );
xor \U$21375 ( \22332 , \3921 , \22205 );
buf g5662_GF_PartitionCandidate( \22333_nG5662 , \22332 );
buf \U$21376 ( \22334 , \22333_nG5662 );
xor \U$21379 ( \22335 , \4096 , \22203 );
buf g5665_GF_PartitionCandidate( \22336_nG5665 , \22335 );
buf \U$21380 ( \22337 , \22336_nG5665 );
xor \U$21383 ( \22338 , \4267 , \22201 );
buf g5668_GF_PartitionCandidate( \22339_nG5668 , \22338 );
buf \U$21384 ( \22340 , \22339_nG5668 );
xor \U$21387 ( \22341 , \4448 , \22199 );
buf g566b_GF_PartitionCandidate( \22342_nG566b , \22341 );
buf \U$21388 ( \22343 , \22342_nG566b );
xor \U$21391 ( \22344 , \4625 , \22197 );
buf g566e_GF_PartitionCandidate( \22345_nG566e , \22344 );
buf \U$21392 ( \22346 , \22345_nG566e );
xor \U$21395 ( \22347 , \4822 , \22195 );
buf g5671_GF_PartitionCandidate( \22348_nG5671 , \22347 );
buf \U$21396 ( \22349 , \22348_nG5671 );
xor \U$21399 ( \22350 , \5018 , \22193 );
buf g5674_GF_PartitionCandidate( \22351_nG5674 , \22350 );
buf \U$21400 ( \22352 , \22351_nG5674 );
xor \U$21403 ( \22353 , \5220 , \22191 );
buf g5677_GF_PartitionCandidate( \22354_nG5677 , \22353 );
buf \U$21404 ( \22355 , \22354_nG5677 );
xor \U$21407 ( \22356 , \5427 , \22189 );
buf g567a_GF_PartitionCandidate( \22357_nG567a , \22356 );
buf \U$21408 ( \22358 , \22357_nG567a );
xor \U$21411 ( \22359 , \5637 , \22187 );
buf g567d_GF_PartitionCandidate( \22360_nG567d , \22359 );
buf \U$21412 ( \22361 , \22360_nG567d );
xor \U$21415 ( \22362 , \6066 , \22185 );
buf g5680_GF_PartitionCandidate( \22363_nG5680 , \22362 );
buf \U$21416 ( \22364 , \22363_nG5680 );
xor \U$21419 ( \22365 , \6309 , \22183 );
buf g5683_GF_PartitionCandidate( \22366_nG5683 , \22365 );
buf \U$21420 ( \22367 , \22366_nG5683 );
xor \U$21423 ( \22368 , \6541 , \22181 );
buf g5686_GF_PartitionCandidate( \22369_nG5686 , \22368 );
buf \U$21424 ( \22370 , \22369_nG5686 );
xor \U$21427 ( \22371 , \6789 , \22179 );
buf g5689_GF_PartitionCandidate( \22372_nG5689 , \22371 );
buf \U$21428 ( \22373 , \22372_nG5689 );
xor \U$21431 ( \22374 , \7042 , \22177 );
buf g568c_GF_PartitionCandidate( \22375_nG568c , \22374 );
buf \U$21432 ( \22376 , \22375_nG568c );
xor \U$21435 ( \22377 , \7298 , \22175 );
buf g568f_GF_PartitionCandidate( \22378_nG568f , \22377 );
buf \U$21436 ( \22379 , \22378_nG568f );
xor \U$21439 ( \22380 , \7555 , \22173 );
buf g5692_GF_PartitionCandidate( \22381_nG5692 , \22380 );
buf \U$21440 ( \22382 , \22381_nG5692 );
xor \U$21443 ( \22383 , \7818 , \22171 );
buf g5695_GF_PartitionCandidate( \22384_nG5695 , \22383 );
buf \U$21444 ( \22385 , \22384_nG5695 );
xor \U$21447 ( \22386 , \8083 , \22169 );
buf g5698_GF_PartitionCandidate( \22387_nG5698 , \22386 );
buf \U$21448 ( \22388 , \22387_nG5698 );
xor \U$21451 ( \22389 , \8344 , \22167 );
buf g569b_GF_PartitionCandidate( \22390_nG569b , \22389 );
buf \U$21452 ( \22391 , \22390_nG569b );
xor \U$21455 ( \22392 , \8610 , \22165 );
buf g569e_GF_PartitionCandidate( \22393_nG569e , \22392 );
buf \U$21456 ( \22394 , \22393_nG569e );
xor \U$21459 ( \22395 , \8876 , \22163 );
buf g56a1_GF_PartitionCandidate( \22396_nG56a1 , \22395 );
buf \U$21460 ( \22397 , \22396_nG56a1 );
xor \U$21463 ( \22398 , \9171 , \22161 );
buf g56a4_GF_PartitionCandidate( \22399_nG56a4 , \22398 );
buf \U$21464 ( \22400 , \22399_nG56a4 );
xor \U$21467 ( \22401 , \9454 , \22159 );
buf g56a7_GF_PartitionCandidate( \22402_nG56a7 , \22401 );
buf \U$21468 ( \22403 , \22402_nG56a7 );
xor \U$21471 ( \22404 , \9742 , \22157 );
buf g56aa_GF_PartitionCandidate( \22405_nG56aa , \22404 );
buf \U$21472 ( \22406 , \22405_nG56aa );
xor \U$21475 ( \22407 , \10043 , \22155 );
buf g56ad_GF_PartitionCandidate( \22408_nG56ad , \22407 );
buf \U$21476 ( \22409 , \22408_nG56ad );
xor \U$21479 ( \22410 , \10339 , \22153 );
buf g56b0_GF_PartitionCandidate( \22411_nG56b0 , \22410 );
buf \U$21480 ( \22412 , \22411_nG56b0 );
xor \U$21483 ( \22413 , \10648 , \22151 );
buf g56b3_GF_PartitionCandidate( \22414_nG56b3 , \22413 );
buf \U$21484 ( \22415 , \22414_nG56b3 );
xor \U$21487 ( \22416 , \10966 , \22149 );
buf g56b6_GF_PartitionCandidate( \22417_nG56b6 , \22416 );
buf \U$21488 ( \22418 , \22417_nG56b6 );
xor \U$21491 ( \22419 , \11282 , \22147 );
buf g56b9_GF_PartitionCandidate( \22420_nG56b9 , \22419 );
buf \U$21492 ( \22421 , \22420_nG56b9 );
xor \U$21495 ( \22422 , \11595 , \22145 );
buf g56bc_GF_PartitionCandidate( \22423_nG56bc , \22422 );
buf \U$21496 ( \22424 , \22423_nG56bc );
xor \U$21499 ( \22425 , \11906 , \22143 );
buf g56bf_GF_PartitionCandidate( \22426_nG56bf , \22425 );
buf \U$21500 ( \22427 , \22426_nG56bf );
xor \U$21503 ( \22428 , \12224 , \22141 );
buf g56c2_GF_PartitionCandidate( \22429_nG56c2 , \22428 );
buf \U$21504 ( \22430 , \22429_nG56c2 );
xor \U$21507 ( \22431 , \12540 , \22139 );
buf g56c5_GF_PartitionCandidate( \22432_nG56c5 , \22431 );
buf \U$21508 ( \22433 , \22432_nG56c5 );
xor \U$21511 ( \22434 , \12840 , \22137 );
buf g56c8_GF_PartitionCandidate( \22435_nG56c8 , \22434 );
buf \U$21512 ( \22436 , \22435_nG56c8 );
xor \U$21515 ( \22437 , \13156 , \22135 );
buf g56cb_GF_PartitionCandidate( \22438_nG56cb , \22437 );
buf \U$21516 ( \22439 , \22438_nG56cb );
xor \U$21519 ( \22440 , \13441 , \22133 );
buf g56ce_GF_PartitionCandidate( \22441_nG56ce , \22440 );
buf \U$21520 ( \22442 , \22441_nG56ce );
xor \U$21523 ( \22443 , \13720 , \22131 );
buf g56d1_GF_PartitionCandidate( \22444_nG56d1 , \22443 );
buf \U$21524 ( \22445 , \22444_nG56d1 );
xor \U$21527 ( \22446 , \14023 , \22129 );
buf g56d4_GF_PartitionCandidate( \22447_nG56d4 , \22446 );
buf \U$21528 ( \22448 , \22447_nG56d4 );
xor \U$21531 ( \22449 , \14294 , \22127 );
buf g56d7_GF_PartitionCandidate( \22450_nG56d7 , \22449 );
buf \U$21532 ( \22451 , \22450_nG56d7 );
xor \U$21535 ( \22452 , \14570 , \22125 );
buf g56da_GF_PartitionCandidate( \22453_nG56da , \22452 );
buf \U$21536 ( \22454 , \22453_nG56da );
xor \U$21539 ( \22455 , \14847 , \22123 );
buf g56dd_GF_PartitionCandidate( \22456_nG56dd , \22455 );
buf \U$21540 ( \22457 , \22456_nG56dd );
xor \U$21543 ( \22458 , \15117 , \22121 );
buf g56e0_GF_PartitionCandidate( \22459_nG56e0 , \22458 );
buf \U$21544 ( \22460 , \22459_nG56e0 );
xor \U$21547 ( \22461 , \15379 , \22119 );
buf g56e3_GF_PartitionCandidate( \22462_nG56e3 , \22461 );
buf \U$21548 ( \22463 , \22462_nG56e3 );
xor \U$21551 ( \22464 , \15640 , \22117 );
buf g56e6_GF_PartitionCandidate( \22465_nG56e6 , \22464 );
buf \U$21552 ( \22466 , \22465_nG56e6 );
xor \U$21555 ( \22467 , \15648 , \22115 );
buf g56e9_GF_PartitionCandidate( \22468_nG56e9 , \22467 );
buf \U$21556 ( \22469 , \22468_nG56e9 );
xor \U$21559 ( \22470 , \15894 , \22113 );
buf g56ec_GF_PartitionCandidate( \22471_nG56ec , \22470 );
buf \U$21560 ( \22472 , \22471_nG56ec );
xor \U$21563 ( \22473 , \16124 , \22111 );
buf g56ef_GF_PartitionCandidate( \22474_nG56ef , \22473 );
buf \U$21564 ( \22475 , \22474_nG56ef );
xor \U$21567 ( \22476 , \16374 , \22109 );
buf g56f2_GF_PartitionCandidate( \22477_nG56f2 , \22476 );
buf \U$21568 ( \22478 , \22477_nG56f2 );
xor \U$21571 ( \22479 , \16599 , \22107 );
buf g56f5_GF_PartitionCandidate( \22480_nG56f5 , \22479 );
buf \U$21572 ( \22481 , \22480_nG56f5 );
xor \U$21575 ( \22482 , \16818 , \22105 );
buf g56f8_GF_PartitionCandidate( \22483_nG56f8 , \22482 );
buf \U$21576 ( \22484 , \22483_nG56f8 );
xor \U$21579 ( \22485 , \17048 , \22103 );
buf g56fb_GF_PartitionCandidate( \22486_nG56fb , \22485 );
buf \U$21580 ( \22487 , \22486_nG56fb );
xor \U$21583 ( \22488 , \17279 , \22101 );
buf g56fe_GF_PartitionCandidate( \22489_nG56fe , \22488 );
buf \U$21584 ( \22490 , \22489_nG56fe );
xor \U$21587 ( \22491 , \17490 , \22099 );
buf g5701_GF_PartitionCandidate( \22492_nG5701 , \22491 );
buf \U$21588 ( \22493 , \22492_nG5701 );
xor \U$21591 ( \22494 , \17703 , \22097 );
buf g5704_GF_PartitionCandidate( \22495_nG5704 , \22494 );
buf \U$21592 ( \22496 , \22495_nG5704 );
xor \U$21595 ( \22497 , \17900 , \22095 );
buf g5707_GF_PartitionCandidate( \22498_nG5707 , \22497 );
buf \U$21596 ( \22499 , \22498_nG5707 );
xor \U$21599 ( \22500 , \18096 , \22093 );
buf g570a_GF_PartitionCandidate( \22501_nG570a , \22500 );
buf \U$21600 ( \22502 , \22501_nG570a );
xor \U$21603 ( \22503 , \18304 , \22091 );
buf g570d_GF_PartitionCandidate( \22504_nG570d , \22503 );
buf \U$21604 ( \22505 , \22504_nG570d );
xor \U$21607 ( \22506 , \18489 , \22089 );
buf g5710_GF_PartitionCandidate( \22507_nG5710 , \22506 );
buf \U$21608 ( \22508 , \22507_nG5710 );
xor \U$21611 ( \22509 , \18676 , \22087 );
buf g5713_GF_PartitionCandidate( \22510_nG5713 , \22509 );
buf \U$21612 ( \22511 , \22510_nG5713 );
xor \U$21615 ( \22512 , \18866 , \22085 );
buf g5716_GF_PartitionCandidate( \22513_nG5716 , \22512 );
buf \U$21616 ( \22514 , \22513_nG5716 );
xor \U$21619 ( \22515 , \19042 , \22083 );
buf g5719_GF_PartitionCandidate( \22516_nG5719 , \22515 );
buf \U$21620 ( \22517 , \22516_nG5719 );
xor \U$21623 ( \22518 , \19213 , \22081 );
buf g571c_GF_PartitionCandidate( \22519_nG571c , \22518 );
buf \U$21624 ( \22520 , \22519_nG571c );
xor \U$21627 ( \22521 , \19221 , \22079 );
buf g571f_GF_PartitionCandidate( \22522_nG571f , \22521 );
buf \U$21628 ( \22523 , \22522_nG571f );
xor \U$21631 ( \22524 , \19389 , \22077 );
buf g5722_GF_PartitionCandidate( \22525_nG5722 , \22524 );
buf \U$21632 ( \22526 , \22525_nG5722 );
xor \U$21635 ( \22527 , \19529 , \22075 );
buf g5725_GF_PartitionCandidate( \22528_nG5725 , \22527 );
buf \U$21636 ( \22529 , \22528_nG5725 );
xor \U$21639 ( \22530 , \19681 , \22073 );
buf g5728_GF_PartitionCandidate( \22531_nG5728 , \22530 );
buf \U$21640 ( \22532 , \22531_nG5728 );
xor \U$21643 ( \22533 , \19845 , \22071 );
buf g572b_GF_PartitionCandidate( \22534_nG572b , \22533 );
buf \U$21644 ( \22535 , \22534_nG572b );
xor \U$21647 ( \22536 , \19984 , \22069 );
buf g572e_GF_PartitionCandidate( \22537_nG572e , \22536 );
buf \U$21648 ( \22538 , \22537_nG572e );
xor \U$21651 ( \22539 , \20109 , \22067 );
buf g5731_GF_PartitionCandidate( \22540_nG5731 , \22539 );
buf \U$21652 ( \22541 , \22540_nG5731 );
xor \U$21655 ( \22542 , \20253 , \22065 );
buf g5734_GF_PartitionCandidate( \22543_nG5734 , \22542 );
buf \U$21656 ( \22544 , \22543_nG5734 );
xor \U$21659 ( \22545 , \20377 , \22063 );
buf g5737_GF_PartitionCandidate( \22546_nG5737 , \22545 );
buf \U$21660 ( \22547 , \22546_nG5737 );
xor \U$21663 ( \22548 , \20517 , \22061 );
buf g573a_GF_PartitionCandidate( \22549_nG573a , \22548 );
buf \U$21664 ( \22550 , \22549_nG573a );
xor \U$21667 ( \22551 , \20641 , \22059 );
buf g573d_GF_PartitionCandidate( \22552_nG573d , \22551 );
buf \U$21668 ( \22553 , \22552_nG573d );
xor \U$21671 ( \22554 , \20756 , \22057 );
buf g5740_GF_PartitionCandidate( \22555_nG5740 , \22554 );
buf \U$21672 ( \22556 , \22555_nG5740 );
xor \U$21675 ( \22557 , \20764 , \22055 );
buf g5743_GF_PartitionCandidate( \22558_nG5743 , \22557 );
buf \U$21676 ( \22559 , \22558_nG5743 );
xor \U$21679 ( \22560 , \20860 , \22053 );
buf g5746_GF_PartitionCandidate( \22561_nG5746 , \22560 );
buf \U$21680 ( \22562 , \22561_nG5746 );
xor \U$21683 ( \22563 , \20975 , \22051 );
buf g5749_GF_PartitionCandidate( \22564_nG5749 , \22563 );
buf \U$21684 ( \22565 , \22564_nG5749 );
xor \U$21687 ( \22566 , \21063 , \22049 );
buf g574c_GF_PartitionCandidate( \22567_nG574c , \22566 );
buf \U$21688 ( \22568 , \22567_nG574c );
xor \U$21691 ( \22569 , \21155 , \22047 );
buf g574f_GF_PartitionCandidate( \22570_nG574f , \22569 );
buf \U$21692 ( \22571 , \22570_nG574f );
xor \U$21695 ( \22572 , \21243 , \22045 );
buf g5752_GF_PartitionCandidate( \22573_nG5752 , \22572 );
buf \U$21696 ( \22574 , \22573_nG5752 );
xor \U$21699 ( \22575 , \21338 , \22043 );
buf g5755_GF_PartitionCandidate( \22576_nG5755 , \22575 );
buf \U$21700 ( \22577 , \22576_nG5755 );
xor \U$21703 ( \22578 , \21418 , \22041 );
buf g5758_GF_PartitionCandidate( \22579_nG5758 , \22578 );
buf \U$21704 ( \22580 , \22579_nG5758 );
xor \U$21707 ( \22581 , \21497 , \22039 );
buf g575b_GF_PartitionCandidate( \22582_nG575b , \22581 );
buf \U$21708 ( \22583 , \22582_nG575b );
xor \U$21711 ( \22584 , \21505 , \22037 );
buf g575e_GF_PartitionCandidate( \22585_nG575e , \22584 );
buf \U$21712 ( \22586 , \22585_nG575e );
xor \U$21715 ( \22587 , \21564 , \22035 );
buf g5761_GF_PartitionCandidate( \22588_nG5761 , \22587 );
buf \U$21716 ( \22589 , \22588_nG5761 );
xor \U$21719 ( \22590 , \21619 , \22033 );
buf g5764_GF_PartitionCandidate( \22591_nG5764 , \22590 );
buf \U$21720 ( \22592 , \22591_nG5764 );
xor \U$21723 ( \22593 , \21690 , \22031 );
buf g5767_GF_PartitionCandidate( \22594_nG5767 , \22593 );
buf \U$21724 ( \22595 , \22594_nG5767 );
xor \U$21727 ( \22596 , \21743 , \22029 );
buf g576a_GF_PartitionCandidate( \22597_nG576a , \22596 );
buf \U$21728 ( \22598 , \22597_nG576a );
xor \U$21731 ( \22599 , \21782 , \22027 );
buf g576d_GF_PartitionCandidate( \22600_nG576d , \22599 );
buf \U$21732 ( \22601 , \22600_nG576d );
xor \U$21735 ( \22602 , \21835 , \22025 );
buf g5770_GF_PartitionCandidate( \22603_nG5770 , \22602 );
buf \U$21736 ( \22604 , \22603_nG5770 );
xor \U$21739 ( \22605 , \21843 , \22023 );
buf g5773_GF_PartitionCandidate( \22606_nG5773 , \22605 );
buf \U$21740 ( \22607 , \22606_nG5773 );
xor \U$21743 ( \22608 , \21877 , \22021 );
buf g5776_GF_PartitionCandidate( \22609_nG5776 , \22608 );
buf \U$21744 ( \22610 , \22609_nG5776 );
xor \U$21747 ( \22611 , \21911 , \22019 );
buf g5779_GF_PartitionCandidate( \22612_nG5779 , \22611 );
buf \U$21748 ( \22613 , \22612_nG5779 );
xor \U$21751 ( \22614 , \21919 , \22017 );
buf g577c_GF_PartitionCandidate( \22615_nG577c , \22614 );
buf \U$21752 ( \22616 , \22615_nG577c );
xor \U$21755 ( \22617 , \21945 , \22015 );
buf g577f_GF_PartitionCandidate( \22618_nG577f , \22617 );
buf \U$21756 ( \22619 , \22618_nG577f );
xor \U$21759 ( \22620 , \21964 , \22013 );
buf g5782_GF_PartitionCandidate( \22621_nG5782 , \22620 );
buf \U$21760 ( \22622 , \22621_nG5782 );
xor \U$21763 ( \22623 , \21972 , \22011 );
buf g5785_GF_PartitionCandidate( \22624_nG5785 , \22623 );
buf \U$21764 ( \22625 , \22624_nG5785 );
xor \U$21767 ( \22626 , \21984 , \22009 );
buf g5788_GF_PartitionCandidate( \22627_nG5788 , \22626 );
buf \U$21768 ( \22628 , \22627_nG5788 );
xor \U$21771 ( \22629 , \21992 , \22007 );
buf g578b_GF_PartitionCandidate( \22630_nG578b , \22629 );
buf \U$21772 ( \22631 , \22630_nG578b );
xor \U$21775 ( \22632 , \21997 , \22005 );
buf g578e_GF_PartitionCandidate( \22633_nG578e , \22632 );
buf \U$21776 ( \22634 , \22633_nG578e );
xor \U$21779 ( \22635 , \22001 , \22004 );
buf g5791_GF_PartitionCandidate( \22636_nG5791 , \22635 );
buf \U$21780 ( \22637 , \22636_nG5791 );
xor \U$21781 ( \22638 , \22003 , \10427 );
buf g5794_GF_PartitionCandidate( \22639_nG5794 , \22638 );
buf \U$21782 ( \22640 , \22639_nG5794 );
_DC g2fd ( \22641_nG2fd , 1'b0 , 1'b1 );
_DC g5796 ( \22642_nG5796 , 1'b0 , 1'b1 );
and g5797_GF_PartitionCandidate( \22643_nG5797 , \22641_nG2fd , \22642_nG5796 );
buf \U$21785 ( \22644 , \22643_nG5797 );
and \U$21786 ( \22645 , \22640 , \22644 );
and \U$21787 ( \22646 , \22637 , \22645 );
or \U$21788 ( \22647 , 1'b0 , 1'b0 , \22646 );
and \U$21789 ( \22648 , \22634 , \22647 );
or \U$21790 ( \22649 , 1'b0 , 1'b0 , \22648 );
and \U$21791 ( \22650 , \22631 , \22649 );
or \U$21792 ( \22651 , 1'b0 , 1'b0 , \22650 );
and \U$21793 ( \22652 , \22628 , \22651 );
or \U$21794 ( \22653 , 1'b0 , 1'b0 , \22652 );
and \U$21795 ( \22654 , \22625 , \22653 );
or \U$21796 ( \22655 , 1'b0 , 1'b0 , \22654 );
and \U$21797 ( \22656 , \22622 , \22655 );
or \U$21798 ( \22657 , 1'b0 , 1'b0 , \22656 );
and \U$21799 ( \22658 , \22619 , \22657 );
or \U$21800 ( \22659 , 1'b0 , 1'b0 , \22658 );
and \U$21801 ( \22660 , \22616 , \22659 );
or \U$21802 ( \22661 , 1'b0 , 1'b0 , \22660 );
and \U$21803 ( \22662 , \22613 , \22661 );
or \U$21804 ( \22663 , 1'b0 , 1'b0 , \22662 );
and \U$21805 ( \22664 , \22610 , \22663 );
or \U$21806 ( \22665 , 1'b0 , 1'b0 , \22664 );
and \U$21807 ( \22666 , \22607 , \22665 );
or \U$21808 ( \22667 , 1'b0 , 1'b0 , \22666 );
and \U$21809 ( \22668 , \22604 , \22667 );
or \U$21810 ( \22669 , 1'b0 , 1'b0 , \22668 );
and \U$21811 ( \22670 , \22601 , \22669 );
or \U$21812 ( \22671 , 1'b0 , 1'b0 , \22670 );
and \U$21813 ( \22672 , \22598 , \22671 );
or \U$21814 ( \22673 , 1'b0 , 1'b0 , \22672 );
and \U$21815 ( \22674 , \22595 , \22673 );
or \U$21816 ( \22675 , 1'b0 , 1'b0 , \22674 );
and \U$21817 ( \22676 , \22592 , \22675 );
or \U$21818 ( \22677 , 1'b0 , 1'b0 , \22676 );
and \U$21819 ( \22678 , \22589 , \22677 );
or \U$21820 ( \22679 , 1'b0 , 1'b0 , \22678 );
and \U$21821 ( \22680 , \22586 , \22679 );
or \U$21822 ( \22681 , 1'b0 , 1'b0 , \22680 );
and \U$21823 ( \22682 , \22583 , \22681 );
or \U$21824 ( \22683 , 1'b0 , 1'b0 , \22682 );
and \U$21825 ( \22684 , \22580 , \22683 );
or \U$21826 ( \22685 , 1'b0 , 1'b0 , \22684 );
and \U$21827 ( \22686 , \22577 , \22685 );
or \U$21828 ( \22687 , 1'b0 , 1'b0 , \22686 );
and \U$21829 ( \22688 , \22574 , \22687 );
or \U$21830 ( \22689 , 1'b0 , 1'b0 , \22688 );
and \U$21831 ( \22690 , \22571 , \22689 );
or \U$21832 ( \22691 , 1'b0 , 1'b0 , \22690 );
and \U$21833 ( \22692 , \22568 , \22691 );
or \U$21834 ( \22693 , 1'b0 , 1'b0 , \22692 );
and \U$21835 ( \22694 , \22565 , \22693 );
or \U$21836 ( \22695 , 1'b0 , 1'b0 , \22694 );
and \U$21837 ( \22696 , \22562 , \22695 );
or \U$21838 ( \22697 , 1'b0 , 1'b0 , \22696 );
and \U$21839 ( \22698 , \22559 , \22697 );
or \U$21840 ( \22699 , 1'b0 , 1'b0 , \22698 );
and \U$21841 ( \22700 , \22556 , \22699 );
or \U$21842 ( \22701 , 1'b0 , 1'b0 , \22700 );
and \U$21843 ( \22702 , \22553 , \22701 );
or \U$21844 ( \22703 , 1'b0 , 1'b0 , \22702 );
and \U$21845 ( \22704 , \22550 , \22703 );
or \U$21846 ( \22705 , 1'b0 , 1'b0 , \22704 );
and \U$21847 ( \22706 , \22547 , \22705 );
or \U$21848 ( \22707 , 1'b0 , 1'b0 , \22706 );
and \U$21849 ( \22708 , \22544 , \22707 );
or \U$21850 ( \22709 , 1'b0 , 1'b0 , \22708 );
and \U$21851 ( \22710 , \22541 , \22709 );
or \U$21852 ( \22711 , 1'b0 , 1'b0 , \22710 );
and \U$21853 ( \22712 , \22538 , \22711 );
or \U$21854 ( \22713 , 1'b0 , 1'b0 , \22712 );
and \U$21855 ( \22714 , \22535 , \22713 );
or \U$21856 ( \22715 , 1'b0 , 1'b0 , \22714 );
and \U$21857 ( \22716 , \22532 , \22715 );
or \U$21858 ( \22717 , 1'b0 , 1'b0 , \22716 );
and \U$21859 ( \22718 , \22529 , \22717 );
or \U$21860 ( \22719 , 1'b0 , 1'b0 , \22718 );
and \U$21861 ( \22720 , \22526 , \22719 );
or \U$21862 ( \22721 , 1'b0 , 1'b0 , \22720 );
and \U$21863 ( \22722 , \22523 , \22721 );
or \U$21864 ( \22723 , 1'b0 , 1'b0 , \22722 );
and \U$21865 ( \22724 , \22520 , \22723 );
or \U$21866 ( \22725 , 1'b0 , 1'b0 , \22724 );
and \U$21867 ( \22726 , \22517 , \22725 );
or \U$21868 ( \22727 , 1'b0 , 1'b0 , \22726 );
and \U$21869 ( \22728 , \22514 , \22727 );
or \U$21870 ( \22729 , 1'b0 , 1'b0 , \22728 );
and \U$21871 ( \22730 , \22511 , \22729 );
or \U$21872 ( \22731 , 1'b0 , 1'b0 , \22730 );
and \U$21873 ( \22732 , \22508 , \22731 );
or \U$21874 ( \22733 , 1'b0 , 1'b0 , \22732 );
and \U$21875 ( \22734 , \22505 , \22733 );
or \U$21876 ( \22735 , 1'b0 , 1'b0 , \22734 );
and \U$21877 ( \22736 , \22502 , \22735 );
or \U$21878 ( \22737 , 1'b0 , 1'b0 , \22736 );
and \U$21879 ( \22738 , \22499 , \22737 );
or \U$21880 ( \22739 , 1'b0 , 1'b0 , \22738 );
and \U$21881 ( \22740 , \22496 , \22739 );
or \U$21882 ( \22741 , 1'b0 , 1'b0 , \22740 );
and \U$21883 ( \22742 , \22493 , \22741 );
or \U$21884 ( \22743 , 1'b0 , 1'b0 , \22742 );
and \U$21885 ( \22744 , \22490 , \22743 );
or \U$21886 ( \22745 , 1'b0 , 1'b0 , \22744 );
and \U$21887 ( \22746 , \22487 , \22745 );
or \U$21888 ( \22747 , 1'b0 , 1'b0 , \22746 );
and \U$21889 ( \22748 , \22484 , \22747 );
or \U$21890 ( \22749 , 1'b0 , 1'b0 , \22748 );
and \U$21891 ( \22750 , \22481 , \22749 );
or \U$21892 ( \22751 , 1'b0 , 1'b0 , \22750 );
and \U$21893 ( \22752 , \22478 , \22751 );
or \U$21894 ( \22753 , 1'b0 , 1'b0 , \22752 );
and \U$21895 ( \22754 , \22475 , \22753 );
or \U$21896 ( \22755 , 1'b0 , 1'b0 , \22754 );
and \U$21897 ( \22756 , \22472 , \22755 );
or \U$21898 ( \22757 , 1'b0 , 1'b0 , \22756 );
and \U$21899 ( \22758 , \22469 , \22757 );
or \U$21900 ( \22759 , 1'b0 , 1'b0 , \22758 );
and \U$21901 ( \22760 , \22466 , \22759 );
or \U$21902 ( \22761 , 1'b0 , 1'b0 , \22760 );
and \U$21903 ( \22762 , \22463 , \22761 );
or \U$21904 ( \22763 , 1'b0 , 1'b0 , \22762 );
and \U$21905 ( \22764 , \22460 , \22763 );
or \U$21906 ( \22765 , 1'b0 , 1'b0 , \22764 );
and \U$21907 ( \22766 , \22457 , \22765 );
or \U$21908 ( \22767 , 1'b0 , 1'b0 , \22766 );
and \U$21909 ( \22768 , \22454 , \22767 );
or \U$21910 ( \22769 , 1'b0 , 1'b0 , \22768 );
and \U$21911 ( \22770 , \22451 , \22769 );
or \U$21912 ( \22771 , 1'b0 , 1'b0 , \22770 );
and \U$21913 ( \22772 , \22448 , \22771 );
or \U$21914 ( \22773 , 1'b0 , 1'b0 , \22772 );
and \U$21915 ( \22774 , \22445 , \22773 );
or \U$21916 ( \22775 , 1'b0 , 1'b0 , \22774 );
and \U$21917 ( \22776 , \22442 , \22775 );
or \U$21918 ( \22777 , 1'b0 , 1'b0 , \22776 );
and \U$21919 ( \22778 , \22439 , \22777 );
or \U$21920 ( \22779 , 1'b0 , 1'b0 , \22778 );
and \U$21921 ( \22780 , \22436 , \22779 );
or \U$21922 ( \22781 , 1'b0 , 1'b0 , \22780 );
and \U$21923 ( \22782 , \22433 , \22781 );
or \U$21924 ( \22783 , 1'b0 , 1'b0 , \22782 );
and \U$21925 ( \22784 , \22430 , \22783 );
or \U$21926 ( \22785 , 1'b0 , 1'b0 , \22784 );
and \U$21927 ( \22786 , \22427 , \22785 );
or \U$21928 ( \22787 , 1'b0 , 1'b0 , \22786 );
and \U$21929 ( \22788 , \22424 , \22787 );
or \U$21930 ( \22789 , 1'b0 , 1'b0 , \22788 );
and \U$21931 ( \22790 , \22421 , \22789 );
or \U$21932 ( \22791 , 1'b0 , 1'b0 , \22790 );
and \U$21933 ( \22792 , \22418 , \22791 );
or \U$21934 ( \22793 , 1'b0 , 1'b0 , \22792 );
and \U$21935 ( \22794 , \22415 , \22793 );
or \U$21936 ( \22795 , 1'b0 , 1'b0 , \22794 );
and \U$21937 ( \22796 , \22412 , \22795 );
or \U$21938 ( \22797 , 1'b0 , 1'b0 , \22796 );
and \U$21939 ( \22798 , \22409 , \22797 );
or \U$21940 ( \22799 , 1'b0 , 1'b0 , \22798 );
and \U$21941 ( \22800 , \22406 , \22799 );
or \U$21942 ( \22801 , 1'b0 , 1'b0 , \22800 );
and \U$21943 ( \22802 , \22403 , \22801 );
or \U$21944 ( \22803 , 1'b0 , 1'b0 , \22802 );
and \U$21945 ( \22804 , \22400 , \22803 );
or \U$21946 ( \22805 , 1'b0 , 1'b0 , \22804 );
and \U$21947 ( \22806 , \22397 , \22805 );
or \U$21948 ( \22807 , 1'b0 , 1'b0 , \22806 );
and \U$21949 ( \22808 , \22394 , \22807 );
or \U$21950 ( \22809 , 1'b0 , 1'b0 , \22808 );
and \U$21951 ( \22810 , \22391 , \22809 );
or \U$21952 ( \22811 , 1'b0 , 1'b0 , \22810 );
and \U$21953 ( \22812 , \22388 , \22811 );
or \U$21954 ( \22813 , 1'b0 , 1'b0 , \22812 );
and \U$21955 ( \22814 , \22385 , \22813 );
or \U$21956 ( \22815 , 1'b0 , 1'b0 , \22814 );
and \U$21957 ( \22816 , \22382 , \22815 );
or \U$21958 ( \22817 , 1'b0 , 1'b0 , \22816 );
and \U$21959 ( \22818 , \22379 , \22817 );
or \U$21960 ( \22819 , 1'b0 , 1'b0 , \22818 );
and \U$21961 ( \22820 , \22376 , \22819 );
or \U$21962 ( \22821 , 1'b0 , 1'b0 , \22820 );
and \U$21963 ( \22822 , \22373 , \22821 );
or \U$21964 ( \22823 , 1'b0 , 1'b0 , \22822 );
and \U$21965 ( \22824 , \22370 , \22823 );
or \U$21966 ( \22825 , 1'b0 , 1'b0 , \22824 );
and \U$21967 ( \22826 , \22367 , \22825 );
or \U$21968 ( \22827 , 1'b0 , 1'b0 , \22826 );
and \U$21969 ( \22828 , \22364 , \22827 );
or \U$21970 ( \22829 , 1'b0 , 1'b0 , \22828 );
and \U$21971 ( \22830 , \22361 , \22829 );
or \U$21972 ( \22831 , 1'b0 , 1'b0 , \22830 );
and \U$21973 ( \22832 , \22358 , \22831 );
or \U$21974 ( \22833 , 1'b0 , 1'b0 , \22832 );
and \U$21975 ( \22834 , \22355 , \22833 );
or \U$21976 ( \22835 , 1'b0 , 1'b0 , \22834 );
and \U$21977 ( \22836 , \22352 , \22835 );
or \U$21978 ( \22837 , 1'b0 , 1'b0 , \22836 );
and \U$21979 ( \22838 , \22349 , \22837 );
or \U$21980 ( \22839 , 1'b0 , 1'b0 , \22838 );
and \U$21981 ( \22840 , \22346 , \22839 );
or \U$21982 ( \22841 , 1'b0 , 1'b0 , \22840 );
and \U$21983 ( \22842 , \22343 , \22841 );
or \U$21984 ( \22843 , 1'b0 , 1'b0 , \22842 );
and \U$21985 ( \22844 , \22340 , \22843 );
or \U$21986 ( \22845 , 1'b0 , 1'b0 , \22844 );
and \U$21987 ( \22846 , \22337 , \22845 );
or \U$21988 ( \22847 , 1'b0 , 1'b0 , \22846 );
and \U$21989 ( \22848 , \22334 , \22847 );
or \U$21990 ( \22849 , 1'b0 , 1'b0 , \22848 );
and \U$21991 ( \22850 , \22331 , \22849 );
or \U$21992 ( \22851 , 1'b0 , 1'b0 , \22850 );
and \U$21993 ( \22852 , \22328 , \22851 );
or \U$21994 ( \22853 , 1'b0 , 1'b0 , \22852 );
and \U$21995 ( \22854 , \22325 , \22853 );
or \U$21996 ( \22855 , 1'b0 , 1'b0 , \22854 );
and \U$21997 ( \22856 , \22322 , \22855 );
or \U$21998 ( \22857 , 1'b0 , 1'b0 , \22856 );
and \U$21999 ( \22858 , \22319 , \22857 );
or \U$22000 ( \22859 , 1'b0 , 1'b0 , \22858 );
and \U$22001 ( \22860 , \22316 , \22859 );
or \U$22002 ( \22861 , 1'b0 , 1'b0 , \22860 );
and \U$22003 ( \22862 , \22313 , \22861 );
or \U$22004 ( \22863 , 1'b0 , 1'b0 , \22862 );
and \U$22005 ( \22864 , \22310 , \22863 );
or \U$22006 ( \22865 , 1'b0 , 1'b0 , \22864 );
and \U$22007 ( \22866 , \22307 , \22865 );
or \U$22008 ( \22867 , 1'b0 , 1'b0 , \22866 );
and \U$22009 ( \22868 , \22304 , \22867 );
or \U$22010 ( \22869 , 1'b0 , 1'b0 , \22868 );
and \U$22011 ( \22870 , \22301 , \22869 );
or \U$22012 ( \22871 , 1'b0 , 1'b0 , \22870 );
and \U$22013 ( \22872 , \22298 , \22871 );
or \U$22014 ( \22873 , 1'b0 , 1'b0 , \22872 );
and \U$22015 ( \22874 , \22295 , \22873 );
or \U$22016 ( \22875 , 1'b0 , 1'b0 , \22874 );
and \U$22017 ( \22876 , \22292 , \22875 );
or \U$22018 ( \22877 , 1'b0 , 1'b0 , \22876 );
and \U$22019 ( \22878 , \22289 , \22877 );
or \U$22020 ( \22879 , 1'b0 , 1'b0 , \22878 );
and \U$22021 ( \22880 , \22286 , \22879 );
or \U$22022 ( \22881 , 1'b0 , 1'b0 , \22880 );
and \U$22023 ( \22882 , \22283 , \22881 );
or \U$22024 ( \22883 , 1'b0 , 1'b0 , \22882 );
and \U$22025 ( \22884 , \22280 , \22883 );
or \U$22026 ( \22885 , 1'b0 , 1'b0 , \22884 );
and \U$22027 ( \22886 , \22277 , \22885 );
or \U$22028 ( \22887 , 1'b0 , 1'b0 , \22886 );
and \U$22029 ( \22888 , \22274 , \22887 );
or \U$22030 ( \22889 , 1'b0 , 1'b0 , \22888 );
and \U$22031 ( \22890 , \22271 , \22889 );
or \U$22032 ( \22891 , 1'b0 , 1'b0 , \22890 );
and \U$22033 ( \22892 , \22268 , \22891 );
or \U$22034 ( \22893 , 1'b0 , 1'b0 , \22892 );
and \U$22035 ( \22894 , \22265 , \22893 );
or \U$22036 ( \22895 , 1'b0 , 1'b0 , \22894 );
and \U$22037 ( \22896 , \22262 , \22895 );
or \U$22038 ( \22897 , 1'b0 , 1'b0 , \22896 );
xor \U$22039 ( \22898 , \22259 , \22897 );
buf g5898_GF_PartitionCandidate( \22899_nG5898 , \22898 );
buf \U$22040 ( \22900 , \22899_nG5898 );
xor \U$22042 ( \22901 , \22262 , 1'b0 );
xor \U$22043 ( \22902 , \22901 , \22895 );
buf g589b_GF_PartitionCandidate( \22903_nG589b , \22902 );
buf \U$22044 ( \22904 , \22903_nG589b );
xor \U$22046 ( \22905 , \22265 , 1'b0 );
xor \U$22047 ( \22906 , \22905 , \22893 );
buf g589e_GF_PartitionCandidate( \22907_nG589e , \22906 );
buf \U$22048 ( \22908 , \22907_nG589e );
xor \U$22050 ( \22909 , \22268 , 1'b0 );
xor \U$22051 ( \22910 , \22909 , \22891 );
buf g58a1_GF_PartitionCandidate( \22911_nG58a1 , \22910 );
buf \U$22052 ( \22912 , \22911_nG58a1 );
xor \U$22054 ( \22913 , \22271 , 1'b0 );
xor \U$22055 ( \22914 , \22913 , \22889 );
buf g58a4_GF_PartitionCandidate( \22915_nG58a4 , \22914 );
buf \U$22056 ( \22916 , \22915_nG58a4 );
xor \U$22058 ( \22917 , \22274 , 1'b0 );
xor \U$22059 ( \22918 , \22917 , \22887 );
buf g58a7_GF_PartitionCandidate( \22919_nG58a7 , \22918 );
buf \U$22060 ( \22920 , \22919_nG58a7 );
xor \U$22062 ( \22921 , \22277 , 1'b0 );
xor \U$22063 ( \22922 , \22921 , \22885 );
buf g58aa_GF_PartitionCandidate( \22923_nG58aa , \22922 );
buf \U$22064 ( \22924 , \22923_nG58aa );
xor \U$22066 ( \22925 , \22280 , 1'b0 );
xor \U$22067 ( \22926 , \22925 , \22883 );
buf g58ad_GF_PartitionCandidate( \22927_nG58ad , \22926 );
buf \U$22068 ( \22928 , \22927_nG58ad );
xor \U$22070 ( \22929 , \22283 , 1'b0 );
xor \U$22071 ( \22930 , \22929 , \22881 );
buf g58b0_GF_PartitionCandidate( \22931_nG58b0 , \22930 );
buf \U$22072 ( \22932 , \22931_nG58b0 );
xor \U$22074 ( \22933 , \22286 , 1'b0 );
xor \U$22075 ( \22934 , \22933 , \22879 );
buf g58b3_GF_PartitionCandidate( \22935_nG58b3 , \22934 );
buf \U$22076 ( \22936 , \22935_nG58b3 );
xor \U$22078 ( \22937 , \22289 , 1'b0 );
xor \U$22079 ( \22938 , \22937 , \22877 );
buf g58b6_GF_PartitionCandidate( \22939_nG58b6 , \22938 );
buf \U$22080 ( \22940 , \22939_nG58b6 );
xor \U$22082 ( \22941 , \22292 , 1'b0 );
xor \U$22083 ( \22942 , \22941 , \22875 );
buf g58b9_GF_PartitionCandidate( \22943_nG58b9 , \22942 );
buf \U$22084 ( \22944 , \22943_nG58b9 );
xor \U$22086 ( \22945 , \22295 , 1'b0 );
xor \U$22087 ( \22946 , \22945 , \22873 );
buf g58bc_GF_PartitionCandidate( \22947_nG58bc , \22946 );
buf \U$22088 ( \22948 , \22947_nG58bc );
xor \U$22090 ( \22949 , \22298 , 1'b0 );
xor \U$22091 ( \22950 , \22949 , \22871 );
buf g58bf_GF_PartitionCandidate( \22951_nG58bf , \22950 );
buf \U$22092 ( \22952 , \22951_nG58bf );
xor \U$22094 ( \22953 , \22301 , 1'b0 );
xor \U$22095 ( \22954 , \22953 , \22869 );
buf g58c2_GF_PartitionCandidate( \22955_nG58c2 , \22954 );
buf \U$22096 ( \22956 , \22955_nG58c2 );
xor \U$22098 ( \22957 , \22304 , 1'b0 );
xor \U$22099 ( \22958 , \22957 , \22867 );
buf g58c5_GF_PartitionCandidate( \22959_nG58c5 , \22958 );
buf \U$22100 ( \22960 , \22959_nG58c5 );
xor \U$22102 ( \22961 , \22307 , 1'b0 );
xor \U$22103 ( \22962 , \22961 , \22865 );
buf g58c8_GF_PartitionCandidate( \22963_nG58c8 , \22962 );
buf \U$22104 ( \22964 , \22963_nG58c8 );
xor \U$22106 ( \22965 , \22310 , 1'b0 );
xor \U$22107 ( \22966 , \22965 , \22863 );
buf g58cb_GF_PartitionCandidate( \22967_nG58cb , \22966 );
buf \U$22108 ( \22968 , \22967_nG58cb );
xor \U$22110 ( \22969 , \22313 , 1'b0 );
xor \U$22111 ( \22970 , \22969 , \22861 );
buf g58ce_GF_PartitionCandidate( \22971_nG58ce , \22970 );
buf \U$22112 ( \22972 , \22971_nG58ce );
xor \U$22114 ( \22973 , \22316 , 1'b0 );
xor \U$22115 ( \22974 , \22973 , \22859 );
buf g58d1_GF_PartitionCandidate( \22975_nG58d1 , \22974 );
buf \U$22116 ( \22976 , \22975_nG58d1 );
xor \U$22118 ( \22977 , \22319 , 1'b0 );
xor \U$22119 ( \22978 , \22977 , \22857 );
buf g58d4_GF_PartitionCandidate( \22979_nG58d4 , \22978 );
buf \U$22120 ( \22980 , \22979_nG58d4 );
xor \U$22122 ( \22981 , \22322 , 1'b0 );
xor \U$22123 ( \22982 , \22981 , \22855 );
buf g58d7_GF_PartitionCandidate( \22983_nG58d7 , \22982 );
buf \U$22124 ( \22984 , \22983_nG58d7 );
xor \U$22126 ( \22985 , \22325 , 1'b0 );
xor \U$22127 ( \22986 , \22985 , \22853 );
buf g58da_GF_PartitionCandidate( \22987_nG58da , \22986 );
buf \U$22128 ( \22988 , \22987_nG58da );
xor \U$22130 ( \22989 , \22328 , 1'b0 );
xor \U$22131 ( \22990 , \22989 , \22851 );
buf g58dd_GF_PartitionCandidate( \22991_nG58dd , \22990 );
buf \U$22132 ( \22992 , \22991_nG58dd );
xor \U$22134 ( \22993 , \22331 , 1'b0 );
xor \U$22135 ( \22994 , \22993 , \22849 );
buf g58e0_GF_PartitionCandidate( \22995_nG58e0 , \22994 );
buf \U$22136 ( \22996 , \22995_nG58e0 );
xor \U$22138 ( \22997 , \22334 , 1'b0 );
xor \U$22139 ( \22998 , \22997 , \22847 );
buf g58e3_GF_PartitionCandidate( \22999_nG58e3 , \22998 );
buf \U$22140 ( \23000 , \22999_nG58e3 );
xor \U$22142 ( \23001 , \22337 , 1'b0 );
xor \U$22143 ( \23002 , \23001 , \22845 );
buf g58e6_GF_PartitionCandidate( \23003_nG58e6 , \23002 );
buf \U$22144 ( \23004 , \23003_nG58e6 );
xor \U$22146 ( \23005 , \22340 , 1'b0 );
xor \U$22147 ( \23006 , \23005 , \22843 );
buf g58e9_GF_PartitionCandidate( \23007_nG58e9 , \23006 );
buf \U$22148 ( \23008 , \23007_nG58e9 );
xor \U$22150 ( \23009 , \22343 , 1'b0 );
xor \U$22151 ( \23010 , \23009 , \22841 );
buf g58ec_GF_PartitionCandidate( \23011_nG58ec , \23010 );
buf \U$22152 ( \23012 , \23011_nG58ec );
xor \U$22154 ( \23013 , \22346 , 1'b0 );
xor \U$22155 ( \23014 , \23013 , \22839 );
buf g58ef_GF_PartitionCandidate( \23015_nG58ef , \23014 );
buf \U$22156 ( \23016 , \23015_nG58ef );
xor \U$22158 ( \23017 , \22349 , 1'b0 );
xor \U$22159 ( \23018 , \23017 , \22837 );
buf g58f2_GF_PartitionCandidate( \23019_nG58f2 , \23018 );
buf \U$22160 ( \23020 , \23019_nG58f2 );
xor \U$22162 ( \23021 , \22352 , 1'b0 );
xor \U$22163 ( \23022 , \23021 , \22835 );
buf g58f5_GF_PartitionCandidate( \23023_nG58f5 , \23022 );
buf \U$22164 ( \23024 , \23023_nG58f5 );
xor \U$22166 ( \23025 , \22355 , 1'b0 );
xor \U$22167 ( \23026 , \23025 , \22833 );
buf g58f8_GF_PartitionCandidate( \23027_nG58f8 , \23026 );
buf \U$22168 ( \23028 , \23027_nG58f8 );
xor \U$22170 ( \23029 , \22358 , 1'b0 );
xor \U$22171 ( \23030 , \23029 , \22831 );
buf g58fb_GF_PartitionCandidate( \23031_nG58fb , \23030 );
buf \U$22172 ( \23032 , \23031_nG58fb );
xor \U$22174 ( \23033 , \22361 , 1'b0 );
xor \U$22175 ( \23034 , \23033 , \22829 );
buf g58fe_GF_PartitionCandidate( \23035_nG58fe , \23034 );
buf \U$22176 ( \23036 , \23035_nG58fe );
xor \U$22178 ( \23037 , \22364 , 1'b0 );
xor \U$22179 ( \23038 , \23037 , \22827 );
buf g5901_GF_PartitionCandidate( \23039_nG5901 , \23038 );
buf \U$22180 ( \23040 , \23039_nG5901 );
xor \U$22182 ( \23041 , \22367 , 1'b0 );
xor \U$22183 ( \23042 , \23041 , \22825 );
buf g5904_GF_PartitionCandidate( \23043_nG5904 , \23042 );
buf \U$22184 ( \23044 , \23043_nG5904 );
xor \U$22186 ( \23045 , \22370 , 1'b0 );
xor \U$22187 ( \23046 , \23045 , \22823 );
buf g5907_GF_PartitionCandidate( \23047_nG5907 , \23046 );
buf \U$22188 ( \23048 , \23047_nG5907 );
xor \U$22190 ( \23049 , \22373 , 1'b0 );
xor \U$22191 ( \23050 , \23049 , \22821 );
buf g590a_GF_PartitionCandidate( \23051_nG590a , \23050 );
buf \U$22192 ( \23052 , \23051_nG590a );
xor \U$22194 ( \23053 , \22376 , 1'b0 );
xor \U$22195 ( \23054 , \23053 , \22819 );
buf g590d_GF_PartitionCandidate( \23055_nG590d , \23054 );
buf \U$22196 ( \23056 , \23055_nG590d );
xor \U$22198 ( \23057 , \22379 , 1'b0 );
xor \U$22199 ( \23058 , \23057 , \22817 );
buf g5910_GF_PartitionCandidate( \23059_nG5910 , \23058 );
buf \U$22200 ( \23060 , \23059_nG5910 );
xor \U$22202 ( \23061 , \22382 , 1'b0 );
xor \U$22203 ( \23062 , \23061 , \22815 );
buf g5913_GF_PartitionCandidate( \23063_nG5913 , \23062 );
buf \U$22204 ( \23064 , \23063_nG5913 );
xor \U$22206 ( \23065 , \22385 , 1'b0 );
xor \U$22207 ( \23066 , \23065 , \22813 );
buf g5916_GF_PartitionCandidate( \23067_nG5916 , \23066 );
buf \U$22208 ( \23068 , \23067_nG5916 );
xor \U$22210 ( \23069 , \22388 , 1'b0 );
xor \U$22211 ( \23070 , \23069 , \22811 );
buf g5919_GF_PartitionCandidate( \23071_nG5919 , \23070 );
buf \U$22212 ( \23072 , \23071_nG5919 );
xor \U$22214 ( \23073 , \22391 , 1'b0 );
xor \U$22215 ( \23074 , \23073 , \22809 );
buf g591c_GF_PartitionCandidate( \23075_nG591c , \23074 );
buf \U$22216 ( \23076 , \23075_nG591c );
xor \U$22218 ( \23077 , \22394 , 1'b0 );
xor \U$22219 ( \23078 , \23077 , \22807 );
buf g591f_GF_PartitionCandidate( \23079_nG591f , \23078 );
buf \U$22220 ( \23080 , \23079_nG591f );
xor \U$22222 ( \23081 , \22397 , 1'b0 );
xor \U$22223 ( \23082 , \23081 , \22805 );
buf g5922_GF_PartitionCandidate( \23083_nG5922 , \23082 );
buf \U$22224 ( \23084 , \23083_nG5922 );
xor \U$22226 ( \23085 , \22400 , 1'b0 );
xor \U$22227 ( \23086 , \23085 , \22803 );
buf g5925_GF_PartitionCandidate( \23087_nG5925 , \23086 );
buf \U$22228 ( \23088 , \23087_nG5925 );
xor \U$22230 ( \23089 , \22403 , 1'b0 );
xor \U$22231 ( \23090 , \23089 , \22801 );
buf g5928_GF_PartitionCandidate( \23091_nG5928 , \23090 );
buf \U$22232 ( \23092 , \23091_nG5928 );
xor \U$22234 ( \23093 , \22406 , 1'b0 );
xor \U$22235 ( \23094 , \23093 , \22799 );
buf g592b_GF_PartitionCandidate( \23095_nG592b , \23094 );
buf \U$22236 ( \23096 , \23095_nG592b );
xor \U$22238 ( \23097 , \22409 , 1'b0 );
xor \U$22239 ( \23098 , \23097 , \22797 );
buf g592e_GF_PartitionCandidate( \23099_nG592e , \23098 );
buf \U$22240 ( \23100 , \23099_nG592e );
xor \U$22242 ( \23101 , \22412 , 1'b0 );
xor \U$22243 ( \23102 , \23101 , \22795 );
buf g5931_GF_PartitionCandidate( \23103_nG5931 , \23102 );
buf \U$22244 ( \23104 , \23103_nG5931 );
xor \U$22246 ( \23105 , \22415 , 1'b0 );
xor \U$22247 ( \23106 , \23105 , \22793 );
buf g5934_GF_PartitionCandidate( \23107_nG5934 , \23106 );
buf \U$22248 ( \23108 , \23107_nG5934 );
xor \U$22250 ( \23109 , \22418 , 1'b0 );
xor \U$22251 ( \23110 , \23109 , \22791 );
buf g5937_GF_PartitionCandidate( \23111_nG5937 , \23110 );
buf \U$22252 ( \23112 , \23111_nG5937 );
xor \U$22254 ( \23113 , \22421 , 1'b0 );
xor \U$22255 ( \23114 , \23113 , \22789 );
buf g593a_GF_PartitionCandidate( \23115_nG593a , \23114 );
buf \U$22256 ( \23116 , \23115_nG593a );
xor \U$22258 ( \23117 , \22424 , 1'b0 );
xor \U$22259 ( \23118 , \23117 , \22787 );
buf g593d_GF_PartitionCandidate( \23119_nG593d , \23118 );
buf \U$22260 ( \23120 , \23119_nG593d );
xor \U$22262 ( \23121 , \22427 , 1'b0 );
xor \U$22263 ( \23122 , \23121 , \22785 );
buf g5940_GF_PartitionCandidate( \23123_nG5940 , \23122 );
buf \U$22264 ( \23124 , \23123_nG5940 );
xor \U$22266 ( \23125 , \22430 , 1'b0 );
xor \U$22267 ( \23126 , \23125 , \22783 );
buf g5943_GF_PartitionCandidate( \23127_nG5943 , \23126 );
buf \U$22268 ( \23128 , \23127_nG5943 );
xor \U$22270 ( \23129 , \22433 , 1'b0 );
xor \U$22271 ( \23130 , \23129 , \22781 );
buf g5946_GF_PartitionCandidate( \23131_nG5946 , \23130 );
buf \U$22272 ( \23132 , \23131_nG5946 );
xor \U$22274 ( \23133 , \22436 , 1'b0 );
xor \U$22275 ( \23134 , \23133 , \22779 );
buf g5949_GF_PartitionCandidate( \23135_nG5949 , \23134 );
buf \U$22276 ( \23136 , \23135_nG5949 );
xor \U$22278 ( \23137 , \22439 , 1'b0 );
xor \U$22279 ( \23138 , \23137 , \22777 );
buf g594c_GF_PartitionCandidate( \23139_nG594c , \23138 );
buf \U$22280 ( \23140 , \23139_nG594c );
xor \U$22282 ( \23141 , \22442 , 1'b0 );
xor \U$22283 ( \23142 , \23141 , \22775 );
buf g594f_GF_PartitionCandidate( \23143_nG594f , \23142 );
buf \U$22284 ( \23144 , \23143_nG594f );
xor \U$22286 ( \23145 , \22445 , 1'b0 );
xor \U$22287 ( \23146 , \23145 , \22773 );
buf g5952_GF_PartitionCandidate( \23147_nG5952 , \23146 );
buf \U$22288 ( \23148 , \23147_nG5952 );
xor \U$22290 ( \23149 , \22448 , 1'b0 );
xor \U$22291 ( \23150 , \23149 , \22771 );
buf g5955_GF_PartitionCandidate( \23151_nG5955 , \23150 );
buf \U$22292 ( \23152 , \23151_nG5955 );
xor \U$22294 ( \23153 , \22451 , 1'b0 );
xor \U$22295 ( \23154 , \23153 , \22769 );
buf g5958_GF_PartitionCandidate( \23155_nG5958 , \23154 );
buf \U$22296 ( \23156 , \23155_nG5958 );
xor \U$22298 ( \23157 , \22454 , 1'b0 );
xor \U$22299 ( \23158 , \23157 , \22767 );
buf g595b_GF_PartitionCandidate( \23159_nG595b , \23158 );
buf \U$22300 ( \23160 , \23159_nG595b );
xor \U$22302 ( \23161 , \22457 , 1'b0 );
xor \U$22303 ( \23162 , \23161 , \22765 );
buf g595e_GF_PartitionCandidate( \23163_nG595e , \23162 );
buf \U$22304 ( \23164 , \23163_nG595e );
xor \U$22306 ( \23165 , \22460 , 1'b0 );
xor \U$22307 ( \23166 , \23165 , \22763 );
buf g5961_GF_PartitionCandidate( \23167_nG5961 , \23166 );
buf \U$22308 ( \23168 , \23167_nG5961 );
xor \U$22310 ( \23169 , \22463 , 1'b0 );
xor \U$22311 ( \23170 , \23169 , \22761 );
buf g5964_GF_PartitionCandidate( \23171_nG5964 , \23170 );
buf \U$22312 ( \23172 , \23171_nG5964 );
xor \U$22314 ( \23173 , \22466 , 1'b0 );
xor \U$22315 ( \23174 , \23173 , \22759 );
buf g5967_GF_PartitionCandidate( \23175_nG5967 , \23174 );
buf \U$22316 ( \23176 , \23175_nG5967 );
xor \U$22318 ( \23177 , \22469 , 1'b0 );
xor \U$22319 ( \23178 , \23177 , \22757 );
buf g596a_GF_PartitionCandidate( \23179_nG596a , \23178 );
buf \U$22320 ( \23180 , \23179_nG596a );
xor \U$22322 ( \23181 , \22472 , 1'b0 );
xor \U$22323 ( \23182 , \23181 , \22755 );
buf g596d_GF_PartitionCandidate( \23183_nG596d , \23182 );
buf \U$22324 ( \23184 , \23183_nG596d );
xor \U$22326 ( \23185 , \22475 , 1'b0 );
xor \U$22327 ( \23186 , \23185 , \22753 );
buf g5970_GF_PartitionCandidate( \23187_nG5970 , \23186 );
buf \U$22328 ( \23188 , \23187_nG5970 );
xor \U$22330 ( \23189 , \22478 , 1'b0 );
xor \U$22331 ( \23190 , \23189 , \22751 );
buf g5973_GF_PartitionCandidate( \23191_nG5973 , \23190 );
buf \U$22332 ( \23192 , \23191_nG5973 );
xor \U$22334 ( \23193 , \22481 , 1'b0 );
xor \U$22335 ( \23194 , \23193 , \22749 );
buf g5976_GF_PartitionCandidate( \23195_nG5976 , \23194 );
buf \U$22336 ( \23196 , \23195_nG5976 );
xor \U$22338 ( \23197 , \22484 , 1'b0 );
xor \U$22339 ( \23198 , \23197 , \22747 );
buf g5979_GF_PartitionCandidate( \23199_nG5979 , \23198 );
buf \U$22340 ( \23200 , \23199_nG5979 );
xor \U$22342 ( \23201 , \22487 , 1'b0 );
xor \U$22343 ( \23202 , \23201 , \22745 );
buf g597c_GF_PartitionCandidate( \23203_nG597c , \23202 );
buf \U$22344 ( \23204 , \23203_nG597c );
xor \U$22346 ( \23205 , \22490 , 1'b0 );
xor \U$22347 ( \23206 , \23205 , \22743 );
buf g597f_GF_PartitionCandidate( \23207_nG597f , \23206 );
buf \U$22348 ( \23208 , \23207_nG597f );
xor \U$22350 ( \23209 , \22493 , 1'b0 );
xor \U$22351 ( \23210 , \23209 , \22741 );
buf g5982_GF_PartitionCandidate( \23211_nG5982 , \23210 );
buf \U$22352 ( \23212 , \23211_nG5982 );
xor \U$22354 ( \23213 , \22496 , 1'b0 );
xor \U$22355 ( \23214 , \23213 , \22739 );
buf g5985_GF_PartitionCandidate( \23215_nG5985 , \23214 );
buf \U$22356 ( \23216 , \23215_nG5985 );
xor \U$22358 ( \23217 , \22499 , 1'b0 );
xor \U$22359 ( \23218 , \23217 , \22737 );
buf g5988_GF_PartitionCandidate( \23219_nG5988 , \23218 );
buf \U$22360 ( \23220 , \23219_nG5988 );
xor \U$22362 ( \23221 , \22502 , 1'b0 );
xor \U$22363 ( \23222 , \23221 , \22735 );
buf g598b_GF_PartitionCandidate( \23223_nG598b , \23222 );
buf \U$22364 ( \23224 , \23223_nG598b );
xor \U$22366 ( \23225 , \22505 , 1'b0 );
xor \U$22367 ( \23226 , \23225 , \22733 );
buf g598e_GF_PartitionCandidate( \23227_nG598e , \23226 );
buf \U$22368 ( \23228 , \23227_nG598e );
xor \U$22370 ( \23229 , \22508 , 1'b0 );
xor \U$22371 ( \23230 , \23229 , \22731 );
buf g5991_GF_PartitionCandidate( \23231_nG5991 , \23230 );
buf \U$22372 ( \23232 , \23231_nG5991 );
xor \U$22374 ( \23233 , \22511 , 1'b0 );
xor \U$22375 ( \23234 , \23233 , \22729 );
buf g5994_GF_PartitionCandidate( \23235_nG5994 , \23234 );
buf \U$22376 ( \23236 , \23235_nG5994 );
xor \U$22378 ( \23237 , \22514 , 1'b0 );
xor \U$22379 ( \23238 , \23237 , \22727 );
buf g5997_GF_PartitionCandidate( \23239_nG5997 , \23238 );
buf \U$22380 ( \23240 , \23239_nG5997 );
xor \U$22382 ( \23241 , \22517 , 1'b0 );
xor \U$22383 ( \23242 , \23241 , \22725 );
buf g599a_GF_PartitionCandidate( \23243_nG599a , \23242 );
buf \U$22384 ( \23244 , \23243_nG599a );
xor \U$22386 ( \23245 , \22520 , 1'b0 );
xor \U$22387 ( \23246 , \23245 , \22723 );
buf g599d_GF_PartitionCandidate( \23247_nG599d , \23246 );
buf \U$22388 ( \23248 , \23247_nG599d );
xor \U$22390 ( \23249 , \22523 , 1'b0 );
xor \U$22391 ( \23250 , \23249 , \22721 );
buf g59a0_GF_PartitionCandidate( \23251_nG59a0 , \23250 );
buf \U$22392 ( \23252 , \23251_nG59a0 );
xor \U$22394 ( \23253 , \22526 , 1'b0 );
xor \U$22395 ( \23254 , \23253 , \22719 );
buf g59a3_GF_PartitionCandidate( \23255_nG59a3 , \23254 );
buf \U$22396 ( \23256 , \23255_nG59a3 );
xor \U$22398 ( \23257 , \22529 , 1'b0 );
xor \U$22399 ( \23258 , \23257 , \22717 );
buf g59a6_GF_PartitionCandidate( \23259_nG59a6 , \23258 );
buf \U$22400 ( \23260 , \23259_nG59a6 );
xor \U$22402 ( \23261 , \22532 , 1'b0 );
xor \U$22403 ( \23262 , \23261 , \22715 );
buf g59a9_GF_PartitionCandidate( \23263_nG59a9 , \23262 );
buf \U$22404 ( \23264 , \23263_nG59a9 );
xor \U$22406 ( \23265 , \22535 , 1'b0 );
xor \U$22407 ( \23266 , \23265 , \22713 );
buf g59ac_GF_PartitionCandidate( \23267_nG59ac , \23266 );
buf \U$22408 ( \23268 , \23267_nG59ac );
xor \U$22410 ( \23269 , \22538 , 1'b0 );
xor \U$22411 ( \23270 , \23269 , \22711 );
buf g59af_GF_PartitionCandidate( \23271_nG59af , \23270 );
buf \U$22412 ( \23272 , \23271_nG59af );
xor \U$22414 ( \23273 , \22541 , 1'b0 );
xor \U$22415 ( \23274 , \23273 , \22709 );
buf g59b2_GF_PartitionCandidate( \23275_nG59b2 , \23274 );
buf \U$22416 ( \23276 , \23275_nG59b2 );
xor \U$22418 ( \23277 , \22544 , 1'b0 );
xor \U$22419 ( \23278 , \23277 , \22707 );
buf g59b5_GF_PartitionCandidate( \23279_nG59b5 , \23278 );
buf \U$22420 ( \23280 , \23279_nG59b5 );
xor \U$22422 ( \23281 , \22547 , 1'b0 );
xor \U$22423 ( \23282 , \23281 , \22705 );
buf g59b8_GF_PartitionCandidate( \23283_nG59b8 , \23282 );
buf \U$22424 ( \23284 , \23283_nG59b8 );
xor \U$22426 ( \23285 , \22550 , 1'b0 );
xor \U$22427 ( \23286 , \23285 , \22703 );
buf g59bb_GF_PartitionCandidate( \23287_nG59bb , \23286 );
buf \U$22428 ( \23288 , \23287_nG59bb );
xor \U$22430 ( \23289 , \22553 , 1'b0 );
xor \U$22431 ( \23290 , \23289 , \22701 );
buf g59be_GF_PartitionCandidate( \23291_nG59be , \23290 );
buf \U$22432 ( \23292 , \23291_nG59be );
xor \U$22434 ( \23293 , \22556 , 1'b0 );
xor \U$22435 ( \23294 , \23293 , \22699 );
buf g59c1_GF_PartitionCandidate( \23295_nG59c1 , \23294 );
buf \U$22436 ( \23296 , \23295_nG59c1 );
xor \U$22438 ( \23297 , \22559 , 1'b0 );
xor \U$22439 ( \23298 , \23297 , \22697 );
buf g59c4_GF_PartitionCandidate( \23299_nG59c4 , \23298 );
buf \U$22440 ( \23300 , \23299_nG59c4 );
xor \U$22442 ( \23301 , \22562 , 1'b0 );
xor \U$22443 ( \23302 , \23301 , \22695 );
buf g59c7_GF_PartitionCandidate( \23303_nG59c7 , \23302 );
buf \U$22444 ( \23304 , \23303_nG59c7 );
xor \U$22446 ( \23305 , \22565 , 1'b0 );
xor \U$22447 ( \23306 , \23305 , \22693 );
buf g59ca_GF_PartitionCandidate( \23307_nG59ca , \23306 );
buf \U$22448 ( \23308 , \23307_nG59ca );
xor \U$22450 ( \23309 , \22568 , 1'b0 );
xor \U$22451 ( \23310 , \23309 , \22691 );
buf g59cd_GF_PartitionCandidate( \23311_nG59cd , \23310 );
buf \U$22452 ( \23312 , \23311_nG59cd );
xor \U$22454 ( \23313 , \22571 , 1'b0 );
xor \U$22455 ( \23314 , \23313 , \22689 );
buf g59d0_GF_PartitionCandidate( \23315_nG59d0 , \23314 );
buf \U$22456 ( \23316 , \23315_nG59d0 );
xor \U$22458 ( \23317 , \22574 , 1'b0 );
xor \U$22459 ( \23318 , \23317 , \22687 );
buf g59d3_GF_PartitionCandidate( \23319_nG59d3 , \23318 );
buf \U$22460 ( \23320 , \23319_nG59d3 );
xor \U$22462 ( \23321 , \22577 , 1'b0 );
xor \U$22463 ( \23322 , \23321 , \22685 );
buf g59d6_GF_PartitionCandidate( \23323_nG59d6 , \23322 );
buf \U$22464 ( \23324 , \23323_nG59d6 );
xor \U$22466 ( \23325 , \22580 , 1'b0 );
xor \U$22467 ( \23326 , \23325 , \22683 );
buf g59d9_GF_PartitionCandidate( \23327_nG59d9 , \23326 );
buf \U$22468 ( \23328 , \23327_nG59d9 );
xor \U$22470 ( \23329 , \22583 , 1'b0 );
xor \U$22471 ( \23330 , \23329 , \22681 );
buf g59dc_GF_PartitionCandidate( \23331_nG59dc , \23330 );
buf \U$22472 ( \23332 , \23331_nG59dc );
xor \U$22474 ( \23333 , \22586 , 1'b0 );
xor \U$22475 ( \23334 , \23333 , \22679 );
buf g59df_GF_PartitionCandidate( \23335_nG59df , \23334 );
buf \U$22476 ( \23336 , \23335_nG59df );
xor \U$22478 ( \23337 , \22589 , 1'b0 );
xor \U$22479 ( \23338 , \23337 , \22677 );
buf g59e2_GF_PartitionCandidate( \23339_nG59e2 , \23338 );
buf \U$22480 ( \23340 , \23339_nG59e2 );
xor \U$22482 ( \23341 , \22592 , 1'b0 );
xor \U$22483 ( \23342 , \23341 , \22675 );
buf g59e5_GF_PartitionCandidate( \23343_nG59e5 , \23342 );
buf \U$22484 ( \23344 , \23343_nG59e5 );
xor \U$22486 ( \23345 , \22595 , 1'b0 );
xor \U$22487 ( \23346 , \23345 , \22673 );
buf g59e8_GF_PartitionCandidate( \23347_nG59e8 , \23346 );
buf \U$22488 ( \23348 , \23347_nG59e8 );
xor \U$22490 ( \23349 , \22598 , 1'b0 );
xor \U$22491 ( \23350 , \23349 , \22671 );
buf g59eb_GF_PartitionCandidate( \23351_nG59eb , \23350 );
buf \U$22492 ( \23352 , \23351_nG59eb );
xor \U$22494 ( \23353 , \22601 , 1'b0 );
xor \U$22495 ( \23354 , \23353 , \22669 );
buf g59ee_GF_PartitionCandidate( \23355_nG59ee , \23354 );
buf \U$22496 ( \23356 , \23355_nG59ee );
endmodule

