//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RIc224f40_83,RIc229e00_147,RIc224ec8_84,RIc229e78_148,RIc224fb8_82,RIc229d88_146,RIc225030_81,RIc229d10_145,RIc224d60_87,
        RIc229fe0_151,RIc224ce8_88,RIc22a058_152,RIc224e50_85,RIc229ef0_149,RIc224dd8_86,RIc229f68_150,RIc224a90_93,RIc22a2b0_157,RIc224a18_94,
        RIc22a328_158,RIc2249a0_95,RIc22a3a0_159,RIc224928_96,RIc22a418_160,RIc224bf8_90,RIc22a148_154,RIc224c70_89,RIc22a0d0_153,RIc224b80_91,
        RIc22a1c0_155,RIc224b08_92,RIc22a238_156,RIc225300_75,RIc229a40_139,RIc225288_76,RIc229ab8_140,RIc2253f0_73,RIc229950_137,RIc225378_74,
        RIc2299c8_138,RIc2250a8_80,RIc229c98_144,RIc225120_79,RIc229c20_143,RIc225210_77,RIc229b30_141,RIc225198_78,RIc229ba8_142,RIc225558_70,
        RIc2297e8_134,RIc2255d0_69,RIc229770_133,RIc2254e0_71,RIc229860_135,RIc225468_72,RIc2298d8_136,RIc225648_68,RIc2296f8_132,RIc223f50_117,
        RIc22adf0_181,RIc223ed8_118,RIc22ae68_182,RIc223e60_119,RIc22aee0_183,RIc223de8_120,RIc22af58_184,RIc224040_115,RIc22ad00_179,RIc22ad78_180,
        RIc223fc8_116,RIc2240b8_114,RIc22ac88_178,RIc224130_113,RIc22ac10_177,RIc223b90_125,RIc22b1b0_189,RIc2294a0_127,RIc22b2a0_191,RIc229518_128,
        RIc22b318_192,RIc22b228_190,RIc223b18_126,RIc223cf8_122,RIc22b048_186,RIc223d70_121,RIc22afd0_185,RIc223c80_123,RIc22b0c0_187,RIc223c08_124,
        RIc22b138_188,RIc2245e0_103,RIc22a760_167,RIc224568_104,RIc22a7d8_168,RIc224658_102,RIc22a6e8_166,RIc2246d0_101,RIc22a670_165,RIc224298_110,
        RIc22aaa8_174,RIc224310_109,RIc22aa30_173,RIc224220_111,RIc22ab20_175,RIc224388_108,RIc22a9b8_172,RIc2241a8_112,RIc22ab98_176,RIc224478_106,
        RIc22a8c8_170,RIc22a850_169,RIc2244f0_105,RIc224400_107,RIc22a940_171,RIc2248b0_97,RIc22a490_161,RIc224838_98,RIc22a508_162,RIc2247c0_99,
        RIc22a580_163,RIc224748_100,RIc22a5f8_164,RIc2256c0_67,RIc229680_131,RIc2275b0_1,RIc2274c0_3,RIc227538_2,RIc225738_66,RIc229608_130,
        RIc2257b0_65,RIc229590_129,RIc2273d0_5,RIc227358_6,RIc2272e0_7,RIc227448_4,RIc2271f0_9,RIc227268_8,RIc227100_11,RIc227088_12,
        RIc227010_13,RIc227178_10,RIc226f98_14,RIc226f20_15,RIc226ae8_24,RIc226a70_25,RIc226b60_23,RIc226db8_18,RIc226e30_17,RIc226d40_19,
        RIc226818_30,RIc2267a0_31,RIc226890_29,RIc226908_28,RIc226980_27,RIc2269f8_26,RIc226ea8_16,RIc226bd8_22,RIc226c50_21,RIc226cc8_20,
        RIc226728_32,RIc2266b0_33,RIc2265c0_35,RIc226638_34,RIc2264d0_37,RIc226548_36,RIc226458_38,RIc2263e0_39,RIc226368_40,RIc2262f0_41,
        RIc225c60_55,RIc225cd8_54,RIc225d50_53,RIc226188_44,RIc226110_45,RIc226200_43,RIc226098_46,RIc226020_47,RIc225dc8_52,RIc225e40_51,
        RIc225f30_49,RIc225eb8_50,RIc225fa8_48,RIc226278_42,RIc225a80_59,RIc225af8_58,RIc225b70_57,RIc225a08_60,RIc225990_61,RIc225be8_56,
        RIc225918_62,RIc2258a0_63,RIc225828_64,RIc22c560_231,RIc22cb78_244,RIc22c218_224,RIc22b660_199,RIc22b840_203,RIc22cd58_248,RIc22b9a8_206,
        RIc22c038_220,RIc22c0b0_221,RIc22b930_205,RIc22c740_235,RIc22cc68_246,RIc22bc00_211,RIc22cce0_247,RIc22bed0_217,RIc22bcf0_213,RIc22c8a8_238,
        RIc22ba20_207,RIc22c4e8_230,RIc22ce48_250,RIc22b480_195,RIc22cfb0_253,RIc22c998_240,RIc22b6d8_200,RIc22b8b8_204,RIc22c920_239,RIc22b7c8_202,
        RIc22c128_222,RIc22c6c8_234,RIc22d028_254,RIc22c650_233,RIc22c5d8_232,RIc22bde0_215,RIc22bd68_214,RIc22be58_216,RIc22c7b8_236,RIc22b408_194,
        RIc22d0a0_255,RIc22b750_201,RIc22c1a0_223,RIc22bb88_210,RIc22cf38_252,RIc22bc78_212,RIc22c830_237,RIc22c290_225,RIc22b5e8_198,RIc22cbf0_245,
        RIc22cec0_251,RIc22bf48_218,RIc22bb10_209,RIc22c3f8_228,RIc22ca88_242,RIc22b4f8_196,RIc22cdd0_249,RIc22ba98_208,RIc22bfc0_219,RIc22ca10_241,
        RIc22b570_197,RIc22c470_229,RIc22cb00_243,RIc22b390_193,RIc22d118_256,RIc22c380_227,RIc22c308_226,R_101_9cd3d68,R_102_9cd3e10,R_103_9cd3eb8,
        R_104_9cd3f60,R_105_9cd4008,R_106_9cd40b0,R_107_9cd4158,R_108_9cd4200,R_109_9cd42a8,R_10a_9cd4350,R_10b_9cd43f8,R_10c_9cd44a0,R_10d_9cd4548,
        R_10e_9cd45f0,R_10f_9cd4698,R_110_9cd4740,R_111_9cd47e8,R_112_9cd4890,R_113_9cd4938,R_114_9cd49e0,R_115_9cd4a88,R_116_9cd4b30,R_117_9cd4bd8,
        R_118_9cd4c80,R_119_9cd4d28,R_11a_9cd4dd0,R_11b_9cd4e78,R_11c_9cd4f20,R_11d_9cd4fc8,R_11e_9cd5070,R_11f_9cd5118,R_120_9cd51c0,R_121_9cd5268,
        R_122_9cd5310,R_123_9cd53b8,R_124_9cd5460,R_125_9cd5508,R_126_9cd55b0,R_127_9cd5658,R_128_9cd5700,R_129_9cd57a8,R_12a_9cd5850,R_12b_9cd58f8,
        R_12c_9cd59a0,R_12d_9cd5a48,R_12e_9cd5af0,R_12f_9cd5b98,R_130_9cd5c40,R_131_9cd5ce8,R_132_9cd5d90,R_133_9cd5e38,R_134_9cd5ee0,R_135_9cd5f88,
        R_136_9cd6030,R_137_9cd60d8,R_138_9cd6180,R_139_9cd6228,R_13a_9cd62d0,R_13b_9cd6378,R_13c_9cd6420,R_13d_9cd64c8,R_13e_9cd6570,R_13f_9cd6618,
        R_140_9cd66c0,R_141_9cd6768,R_142_9cd6810,R_143_9cd68b8,R_144_9cd6960,R_145_9cd6a08,R_146_9cd6ab0,R_147_9cd6b58,R_148_9cd6c00,R_149_9cd6ca8,
        R_14a_9cd6d50,R_14b_9cd6df8,R_14c_9cd6ea0,R_14d_9cd6f48,R_14e_9cd6ff0,R_14f_9cd7098,R_150_9cd7140,R_151_9cd71e8,R_152_9cd7290,R_153_9cd7338,
        R_154_9cd73e0,R_155_9cd7488,R_156_9cd7530,R_157_9cd75d8,R_158_9cd7680,R_159_9cd7728,R_15a_9cd77d0,R_15b_9cd7878,R_15c_9cd7920,R_15d_9cd79c8,
        R_15e_9cd7a70,R_15f_9cd7b18,R_160_9cd7bc0,R_161_9cd7c68,R_162_9cd7d10,R_163_9cd7db8,R_164_9cd7e60,R_165_9cd7f08,R_166_9cd7fb0,R_167_9cd8058,
        R_168_9cd8100,R_169_9cd81a8,R_16a_9cd8250,R_16b_9cd82f8,R_16c_9cd83a0,R_16d_9cd8448,R_16e_9cd84f0,R_16f_9cd8598,R_170_9cd8640,R_171_9cd86e8,
        R_172_9cd8790,R_173_9cd8838,R_174_9cd88e0,R_175_9cd8988,R_176_9cd8a30,R_177_9cd8ad8);
input RIc224f40_83,RIc229e00_147,RIc224ec8_84,RIc229e78_148,RIc224fb8_82,RIc229d88_146,RIc225030_81,RIc229d10_145,RIc224d60_87,
        RIc229fe0_151,RIc224ce8_88,RIc22a058_152,RIc224e50_85,RIc229ef0_149,RIc224dd8_86,RIc229f68_150,RIc224a90_93,RIc22a2b0_157,RIc224a18_94,
        RIc22a328_158,RIc2249a0_95,RIc22a3a0_159,RIc224928_96,RIc22a418_160,RIc224bf8_90,RIc22a148_154,RIc224c70_89,RIc22a0d0_153,RIc224b80_91,
        RIc22a1c0_155,RIc224b08_92,RIc22a238_156,RIc225300_75,RIc229a40_139,RIc225288_76,RIc229ab8_140,RIc2253f0_73,RIc229950_137,RIc225378_74,
        RIc2299c8_138,RIc2250a8_80,RIc229c98_144,RIc225120_79,RIc229c20_143,RIc225210_77,RIc229b30_141,RIc225198_78,RIc229ba8_142,RIc225558_70,
        RIc2297e8_134,RIc2255d0_69,RIc229770_133,RIc2254e0_71,RIc229860_135,RIc225468_72,RIc2298d8_136,RIc225648_68,RIc2296f8_132,RIc223f50_117,
        RIc22adf0_181,RIc223ed8_118,RIc22ae68_182,RIc223e60_119,RIc22aee0_183,RIc223de8_120,RIc22af58_184,RIc224040_115,RIc22ad00_179,RIc22ad78_180,
        RIc223fc8_116,RIc2240b8_114,RIc22ac88_178,RIc224130_113,RIc22ac10_177,RIc223b90_125,RIc22b1b0_189,RIc2294a0_127,RIc22b2a0_191,RIc229518_128,
        RIc22b318_192,RIc22b228_190,RIc223b18_126,RIc223cf8_122,RIc22b048_186,RIc223d70_121,RIc22afd0_185,RIc223c80_123,RIc22b0c0_187,RIc223c08_124,
        RIc22b138_188,RIc2245e0_103,RIc22a760_167,RIc224568_104,RIc22a7d8_168,RIc224658_102,RIc22a6e8_166,RIc2246d0_101,RIc22a670_165,RIc224298_110,
        RIc22aaa8_174,RIc224310_109,RIc22aa30_173,RIc224220_111,RIc22ab20_175,RIc224388_108,RIc22a9b8_172,RIc2241a8_112,RIc22ab98_176,RIc224478_106,
        RIc22a8c8_170,RIc22a850_169,RIc2244f0_105,RIc224400_107,RIc22a940_171,RIc2248b0_97,RIc22a490_161,RIc224838_98,RIc22a508_162,RIc2247c0_99,
        RIc22a580_163,RIc224748_100,RIc22a5f8_164,RIc2256c0_67,RIc229680_131,RIc2275b0_1,RIc2274c0_3,RIc227538_2,RIc225738_66,RIc229608_130,
        RIc2257b0_65,RIc229590_129,RIc2273d0_5,RIc227358_6,RIc2272e0_7,RIc227448_4,RIc2271f0_9,RIc227268_8,RIc227100_11,RIc227088_12,
        RIc227010_13,RIc227178_10,RIc226f98_14,RIc226f20_15,RIc226ae8_24,RIc226a70_25,RIc226b60_23,RIc226db8_18,RIc226e30_17,RIc226d40_19,
        RIc226818_30,RIc2267a0_31,RIc226890_29,RIc226908_28,RIc226980_27,RIc2269f8_26,RIc226ea8_16,RIc226bd8_22,RIc226c50_21,RIc226cc8_20,
        RIc226728_32,RIc2266b0_33,RIc2265c0_35,RIc226638_34,RIc2264d0_37,RIc226548_36,RIc226458_38,RIc2263e0_39,RIc226368_40,RIc2262f0_41,
        RIc225c60_55,RIc225cd8_54,RIc225d50_53,RIc226188_44,RIc226110_45,RIc226200_43,RIc226098_46,RIc226020_47,RIc225dc8_52,RIc225e40_51,
        RIc225f30_49,RIc225eb8_50,RIc225fa8_48,RIc226278_42,RIc225a80_59,RIc225af8_58,RIc225b70_57,RIc225a08_60,RIc225990_61,RIc225be8_56,
        RIc225918_62,RIc2258a0_63,RIc225828_64,RIc22c560_231,RIc22cb78_244,RIc22c218_224,RIc22b660_199,RIc22b840_203,RIc22cd58_248,RIc22b9a8_206,
        RIc22c038_220,RIc22c0b0_221,RIc22b930_205,RIc22c740_235,RIc22cc68_246,RIc22bc00_211,RIc22cce0_247,RIc22bed0_217,RIc22bcf0_213,RIc22c8a8_238,
        RIc22ba20_207,RIc22c4e8_230,RIc22ce48_250,RIc22b480_195,RIc22cfb0_253,RIc22c998_240,RIc22b6d8_200,RIc22b8b8_204,RIc22c920_239,RIc22b7c8_202,
        RIc22c128_222,RIc22c6c8_234,RIc22d028_254,RIc22c650_233,RIc22c5d8_232,RIc22bde0_215,RIc22bd68_214,RIc22be58_216,RIc22c7b8_236,RIc22b408_194,
        RIc22d0a0_255,RIc22b750_201,RIc22c1a0_223,RIc22bb88_210,RIc22cf38_252,RIc22bc78_212,RIc22c830_237,RIc22c290_225,RIc22b5e8_198,RIc22cbf0_245,
        RIc22cec0_251,RIc22bf48_218,RIc22bb10_209,RIc22c3f8_228,RIc22ca88_242,RIc22b4f8_196,RIc22cdd0_249,RIc22ba98_208,RIc22bfc0_219,RIc22ca10_241,
        RIc22b570_197,RIc22c470_229,RIc22cb00_243,RIc22b390_193,RIc22d118_256,RIc22c380_227,RIc22c308_226;
output R_101_9cd3d68,R_102_9cd3e10,R_103_9cd3eb8,R_104_9cd3f60,R_105_9cd4008,R_106_9cd40b0,R_107_9cd4158,R_108_9cd4200,R_109_9cd42a8,
        R_10a_9cd4350,R_10b_9cd43f8,R_10c_9cd44a0,R_10d_9cd4548,R_10e_9cd45f0,R_10f_9cd4698,R_110_9cd4740,R_111_9cd47e8,R_112_9cd4890,R_113_9cd4938,
        R_114_9cd49e0,R_115_9cd4a88,R_116_9cd4b30,R_117_9cd4bd8,R_118_9cd4c80,R_119_9cd4d28,R_11a_9cd4dd0,R_11b_9cd4e78,R_11c_9cd4f20,R_11d_9cd4fc8,
        R_11e_9cd5070,R_11f_9cd5118,R_120_9cd51c0,R_121_9cd5268,R_122_9cd5310,R_123_9cd53b8,R_124_9cd5460,R_125_9cd5508,R_126_9cd55b0,R_127_9cd5658,
        R_128_9cd5700,R_129_9cd57a8,R_12a_9cd5850,R_12b_9cd58f8,R_12c_9cd59a0,R_12d_9cd5a48,R_12e_9cd5af0,R_12f_9cd5b98,R_130_9cd5c40,R_131_9cd5ce8,
        R_132_9cd5d90,R_133_9cd5e38,R_134_9cd5ee0,R_135_9cd5f88,R_136_9cd6030,R_137_9cd60d8,R_138_9cd6180,R_139_9cd6228,R_13a_9cd62d0,R_13b_9cd6378,
        R_13c_9cd6420,R_13d_9cd64c8,R_13e_9cd6570,R_13f_9cd6618,R_140_9cd66c0,R_141_9cd6768,R_142_9cd6810,R_143_9cd68b8,R_144_9cd6960,R_145_9cd6a08,
        R_146_9cd6ab0,R_147_9cd6b58,R_148_9cd6c00,R_149_9cd6ca8,R_14a_9cd6d50,R_14b_9cd6df8,R_14c_9cd6ea0,R_14d_9cd6f48,R_14e_9cd6ff0,R_14f_9cd7098,
        R_150_9cd7140,R_151_9cd71e8,R_152_9cd7290,R_153_9cd7338,R_154_9cd73e0,R_155_9cd7488,R_156_9cd7530,R_157_9cd75d8,R_158_9cd7680,R_159_9cd7728,
        R_15a_9cd77d0,R_15b_9cd7878,R_15c_9cd7920,R_15d_9cd79c8,R_15e_9cd7a70,R_15f_9cd7b18,R_160_9cd7bc0,R_161_9cd7c68,R_162_9cd7d10,R_163_9cd7db8,
        R_164_9cd7e60,R_165_9cd7f08,R_166_9cd7fb0,R_167_9cd8058,R_168_9cd8100,R_169_9cd81a8,R_16a_9cd8250,R_16b_9cd82f8,R_16c_9cd83a0,R_16d_9cd8448,
        R_16e_9cd84f0,R_16f_9cd8598,R_170_9cd8640,R_171_9cd86e8,R_172_9cd8790,R_173_9cd8838,R_174_9cd88e0,R_175_9cd8988,R_176_9cd8a30,R_177_9cd8ad8;

wire \376_ZERO , \377_ONE , \378 , \379 , \380 , \381 , \382 , \383 , \384 ,
         \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 , \394 ,
         \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 , \404 ,
         \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 , \414 ,
         \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 , \424 ,
         \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 , \434 ,
         \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 , \444 ,
         \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 , \454 ,
         \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 ,
         \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 , \474 ,
         \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 , \484 ,
         \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 , \494 ,
         \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 ,
         \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 ,
         \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 , \524 ,
         \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 , \534 ,
         \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 , \544 ,
         \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 , \554 ,
         \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 , \564 ,
         \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 , \574 ,
         \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 , \584 ,
         \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 , \594 ,
         \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 , \604 ,
         \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 , \614 ,
         \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 , \624 ,
         \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 , \634 ,
         \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 ,
         \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 ,
         \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 , \664 ,
         \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 , \674 ,
         \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 , \684 ,
         \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 , \694 ,
         \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 ,
         \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 , \714 ,
         \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 , \724 ,
         \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 ,
         \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 , \744 ,
         \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 , \754 ,
         \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 , \764 ,
         \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 , \774 ,
         \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 , \784 ,
         \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794 ,
         \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 , \804 ,
         \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 ,
         \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 , \824 ,
         \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 , \834 ,
         \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 , \844 ,
         \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 , \854 ,
         \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 , \864 ,
         \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 ,
         \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 , \884 ,
         \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 , \894 ,
         \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 , \904 ,
         \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 , \914 ,
         \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 , \924 ,
         \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 , \934 ,
         \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 , \944 ,
         \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 ,
         \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 , \964 ,
         \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 , \974 ,
         \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 , \984 ,
         \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 , \994 ,
         \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 ,
         \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 ,
         \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 ,
         \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 ,
         \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 ,
         \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 ,
         \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 ,
         \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 ,
         \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 ,
         \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 ,
         \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 ,
         \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 ,
         \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 ,
         \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 ,
         \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 ,
         \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 ,
         \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 ,
         \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 ,
         \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 ,
         \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 ,
         \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 ,
         \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 ,
         \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 ,
         \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 ,
         \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 ,
         \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 ,
         \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 ,
         \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 ,
         \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 ,
         \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 ,
         \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 ,
         \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 ,
         \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 ,
         \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 ,
         \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 ,
         \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 ,
         \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 ,
         \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 ,
         \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 ,
         \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 ,
         \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 ,
         \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 ,
         \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 ,
         \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 ,
         \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 ,
         \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 ,
         \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 ,
         \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 ,
         \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 ,
         \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 ,
         \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 ,
         \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 ,
         \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 ,
         \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 ,
         \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 ,
         \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 ,
         \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 ,
         \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 ,
         \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 ,
         \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 ,
         \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 ,
         \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 ,
         \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 ,
         \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 ,
         \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 ,
         \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 ,
         \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 ,
         \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 ,
         \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 ,
         \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 ,
         \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 ,
         \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 ,
         \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 ,
         \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 ,
         \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 ,
         \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 ,
         \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 ,
         \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 ,
         \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 ,
         \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 ,
         \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 ,
         \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 ,
         \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 ,
         \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 ,
         \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 ,
         \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 ,
         \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 ,
         \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 ,
         \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 ,
         \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 ,
         \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 ,
         \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 ,
         \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 ,
         \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 ,
         \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 ,
         \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 ,
         \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 ,
         \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 ,
         \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 ,
         \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 ,
         \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 ,
         \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 ,
         \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 ,
         \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 ,
         \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 ,
         \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 ,
         \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 ,
         \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 ,
         \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 ,
         \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 ,
         \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 ,
         \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 ,
         \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 ,
         \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 ,
         \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 ,
         \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 ,
         \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 ,
         \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 ,
         \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 ,
         \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 ,
         \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 ,
         \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 ,
         \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 ,
         \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 ,
         \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 ,
         \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 ,
         \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 ,
         \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 ,
         \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 ,
         \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 ,
         \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 ,
         \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 ,
         \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 ,
         \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 ,
         \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 ,
         \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 ,
         \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 ,
         \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 ,
         \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 ,
         \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 ,
         \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 ,
         \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 ,
         \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 ,
         \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 ,
         \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 ,
         \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 ,
         \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 ,
         \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 ,
         \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 ,
         \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 ,
         \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 ,
         \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 ,
         \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 ,
         \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 ,
         \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 ,
         \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 ,
         \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 ,
         \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 ,
         \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 ,
         \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 ,
         \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 ,
         \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 ,
         \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 ,
         \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 ,
         \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 ,
         \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 ,
         \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 ,
         \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 ,
         \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 ,
         \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 ,
         \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 ,
         \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 ,
         \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 ,
         \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 ,
         \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 ,
         \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 ,
         \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 ,
         \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 ,
         \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 ,
         \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 ,
         \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 ,
         \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 ,
         \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 ,
         \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 ,
         \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 ,
         \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 ,
         \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 ,
         \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 ,
         \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 ,
         \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 ,
         \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 ,
         \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 ,
         \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 ,
         \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 ,
         \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 ,
         \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 ,
         \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 ,
         \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 ,
         \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 ,
         \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 ,
         \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 ,
         \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 ,
         \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 ,
         \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 ,
         \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 ,
         \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 ,
         \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 ,
         \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 ,
         \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 ,
         \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 ,
         \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 ,
         \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 ,
         \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 ,
         \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 ,
         \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 ,
         \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 ,
         \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 ,
         \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 ,
         \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 ,
         \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 ,
         \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 ,
         \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 ,
         \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 ,
         \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 ,
         \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 ,
         \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 ,
         \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 ,
         \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 ,
         \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 ,
         \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 ,
         \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 ,
         \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 ,
         \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 ,
         \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 ,
         \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 ,
         \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 ,
         \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 ,
         \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 ,
         \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 ,
         \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 ,
         \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 ,
         \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 ,
         \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 ,
         \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 ,
         \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 ,
         \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 ,
         \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 ,
         \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 ,
         \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 ,
         \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 ,
         \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 ,
         \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 ,
         \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 ,
         \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 ,
         \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 ,
         \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 ,
         \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 ,
         \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 ,
         \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 ,
         \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 ,
         \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 ,
         \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 ,
         \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 ,
         \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 ,
         \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 ,
         \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 ,
         \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 ,
         \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 ,
         \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 ,
         \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 ,
         \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 ,
         \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 ,
         \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 ,
         \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 ,
         \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 ,
         \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 ,
         \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 ,
         \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 ,
         \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 ,
         \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 ,
         \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 ,
         \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 ,
         \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 ,
         \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 ,
         \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 ,
         \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 ,
         \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 ,
         \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 ,
         \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 ,
         \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 ,
         \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 ,
         \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 ,
         \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 ,
         \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 ,
         \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 ,
         \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 ,
         \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 ,
         \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 ,
         \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 ,
         \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 ,
         \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 ,
         \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 ,
         \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 ,
         \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 ,
         \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 ,
         \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 ,
         \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 ,
         \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 ,
         \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 ,
         \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 ,
         \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 ,
         \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 ,
         \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 ,
         \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 ,
         \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 ,
         \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 ,
         \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 ,
         \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 ,
         \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 ,
         \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 ,
         \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 ,
         \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 ,
         \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 ,
         \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 ,
         \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 ,
         \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 ,
         \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 ,
         \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 ,
         \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 ,
         \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 ,
         \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 ,
         \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 ,
         \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 ,
         \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 ,
         \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 ,
         \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 ,
         \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 ,
         \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 ,
         \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 ,
         \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 ,
         \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 ,
         \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 ,
         \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 ,
         \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 ,
         \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 ,
         \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 ,
         \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 ,
         \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 ,
         \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 ,
         \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 ,
         \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 ,
         \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 ,
         \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 ,
         \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 ,
         \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 ,
         \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 ,
         \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 ,
         \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 ,
         \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 ,
         \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 ,
         \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 ,
         \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 ,
         \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 ,
         \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 ,
         \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 ,
         \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 ,
         \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 ,
         \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 ,
         \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 ,
         \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 ,
         \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 ,
         \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 ,
         \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 ,
         \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 ,
         \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 ,
         \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 ,
         \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 ,
         \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 ,
         \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 ,
         \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 ,
         \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 ,
         \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 ,
         \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 ,
         \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 ,
         \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 ,
         \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 ,
         \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 ,
         \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 ,
         \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 ,
         \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 ,
         \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 ,
         \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 ,
         \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 ,
         \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 ,
         \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 ,
         \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 ,
         \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 ,
         \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 ,
         \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 ,
         \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 ,
         \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 ,
         \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 ,
         \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 ,
         \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 ,
         \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 ,
         \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 ,
         \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 ,
         \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 ,
         \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 ,
         \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 ,
         \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 ,
         \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 ,
         \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 ,
         \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 ,
         \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 ,
         \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 ,
         \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 ,
         \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 ,
         \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 ,
         \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 ,
         \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 ,
         \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 ,
         \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 ,
         \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 ,
         \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 ,
         \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 ,
         \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 ,
         \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 ,
         \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 ,
         \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 ,
         \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 ,
         \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 ,
         \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 ,
         \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 ,
         \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 ,
         \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 ,
         \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 ,
         \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 ,
         \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 ,
         \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 ,
         \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 ,
         \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 ,
         \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 ,
         \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 ,
         \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 ,
         \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 ,
         \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 ,
         \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 ,
         \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 ,
         \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 ,
         \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 ,
         \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 ,
         \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 ,
         \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 ,
         \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 ,
         \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 ,
         \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 ,
         \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 ,
         \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 ,
         \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 ,
         \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 ,
         \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 ,
         \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 ,
         \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 ,
         \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 ,
         \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 ,
         \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 ,
         \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 ,
         \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 ,
         \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 ,
         \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 ,
         \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 ,
         \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 ,
         \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 ,
         \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 ,
         \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 ,
         \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 ,
         \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 ,
         \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 ,
         \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 ,
         \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 ,
         \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 ,
         \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 ,
         \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 ,
         \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 ,
         \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 ,
         \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 ,
         \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 ,
         \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 ,
         \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 ,
         \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 ,
         \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 ,
         \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 ,
         \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 ,
         \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 ,
         \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 ,
         \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 ,
         \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 ,
         \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 ,
         \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 ,
         \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 ,
         \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 ,
         \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 ,
         \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 ,
         \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 ,
         \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 ,
         \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 ,
         \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 ,
         \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 ,
         \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 ,
         \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 ,
         \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 ,
         \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 ,
         \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 ,
         \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 ,
         \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 ,
         \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 ,
         \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 ,
         \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 ,
         \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 ,
         \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 ,
         \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 ,
         \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 ,
         \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 ,
         \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 ,
         \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 ,
         \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 ,
         \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 ,
         \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 ,
         \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 ,
         \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 ,
         \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 ,
         \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 ,
         \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 ,
         \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 ,
         \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 ,
         \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 ,
         \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 ,
         \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 ,
         \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 ,
         \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 ,
         \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 ,
         \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 ,
         \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 ,
         \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 ,
         \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 ,
         \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 ,
         \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 ,
         \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 ,
         \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 ,
         \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 ,
         \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 ,
         \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 ,
         \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 ,
         \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 ,
         \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 ,
         \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 ,
         \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 ,
         \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 ,
         \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 ,
         \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 ,
         \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 ,
         \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 ,
         \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 ,
         \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 ,
         \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 ,
         \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 ,
         \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 ,
         \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 ,
         \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 ,
         \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 ,
         \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 ,
         \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 ,
         \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 ,
         \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 ,
         \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 ,
         \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 ,
         \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 ,
         \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 ,
         \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 ,
         \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 ,
         \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 ,
         \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 ,
         \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 ,
         \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 ,
         \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 ,
         \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 ,
         \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 ,
         \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 ,
         \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 ,
         \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 ,
         \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 ,
         \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 ,
         \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 ,
         \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 ,
         \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 ,
         \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 ,
         \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 ,
         \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 ,
         \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 ,
         \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 ,
         \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 ,
         \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 ,
         \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 ,
         \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 ,
         \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 ,
         \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 ,
         \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 ,
         \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 ,
         \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 ,
         \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 ,
         \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 ,
         \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 ,
         \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 ,
         \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 ,
         \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 ,
         \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 ,
         \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 ,
         \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 ,
         \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 ,
         \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 ,
         \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 ,
         \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 ,
         \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 ,
         \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 ,
         \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 ,
         \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 ,
         \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 ,
         \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 ,
         \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 ,
         \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 ,
         \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 ,
         \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 ,
         \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 ,
         \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 ,
         \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 ,
         \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 ,
         \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 ,
         \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 ,
         \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 ,
         \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 ,
         \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 ,
         \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 ,
         \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 ,
         \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 ,
         \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 ,
         \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 ,
         \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 ,
         \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 ,
         \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 ,
         \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 ,
         \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 ,
         \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 ,
         \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 ,
         \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 ,
         \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 ,
         \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 ,
         \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 ,
         \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 ,
         \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 ,
         \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 ,
         \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 ,
         \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 ,
         \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 ,
         \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 ,
         \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 ,
         \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 ,
         \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 ,
         \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 ,
         \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 ,
         \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 ,
         \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 ,
         \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 ,
         \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 ,
         \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 ,
         \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 ,
         \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 ,
         \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 , \7773 , \7774 ,
         \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 ,
         \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 ,
         \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 ,
         \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 ,
         \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 ,
         \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 ,
         \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 ,
         \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 ,
         \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 ,
         \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 ,
         \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 ,
         \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 ,
         \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 ,
         \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 ,
         \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 ,
         \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 ,
         \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 ,
         \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 ,
         \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 ,
         \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 ,
         \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 ,
         \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 ,
         \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 ,
         \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 ,
         \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 ,
         \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 ,
         \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 ,
         \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 ,
         \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 ,
         \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 ,
         \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 ,
         \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 ,
         \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 ,
         \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 ,
         \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 ,
         \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 ,
         \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 ,
         \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 ,
         \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 ,
         \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 ,
         \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 ,
         \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 ,
         \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 ,
         \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 ,
         \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 ,
         \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 ,
         \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 ,
         \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 ,
         \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 ,
         \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 ,
         \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 ,
         \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 ,
         \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 ,
         \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 ,
         \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 ,
         \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 ,
         \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 ,
         \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 ,
         \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 ,
         \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 ,
         \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 ,
         \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 ,
         \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 ,
         \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 ,
         \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 ,
         \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 ,
         \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 ,
         \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 ,
         \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 ,
         \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 ,
         \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 ,
         \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 ,
         \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 ,
         \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 ,
         \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 ,
         \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 ,
         \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 ,
         \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 ,
         \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 ,
         \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 ,
         \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 ,
         \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 ,
         \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 ,
         \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 ,
         \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 ,
         \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 ,
         \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 ,
         \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 ,
         \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 ,
         \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 ,
         \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 ,
         \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 ,
         \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 ,
         \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 ,
         \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 ,
         \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 ,
         \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 ,
         \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 ,
         \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 ,
         \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 ,
         \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 ,
         \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 ,
         \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 ,
         \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 ,
         \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 ,
         \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 ,
         \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 ,
         \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 ,
         \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 ,
         \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 ,
         \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 ,
         \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 ,
         \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 ,
         \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 ,
         \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 ,
         \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 ,
         \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 ,
         \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 ,
         \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 ,
         \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 ,
         \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 ,
         \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 ,
         \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 ,
         \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 ,
         \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 ,
         \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 ,
         \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 ,
         \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 ,
         \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 ,
         \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 ,
         \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 ,
         \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 ,
         \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 ,
         \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 ,
         \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 ,
         \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 ,
         \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 ,
         \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 ,
         \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 ,
         \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 ,
         \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 ,
         \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 ,
         \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 ,
         \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 ,
         \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 ,
         \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 ,
         \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 ,
         \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 ,
         \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 ,
         \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 ,
         \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 ,
         \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 ,
         \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 ,
         \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 ,
         \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 ,
         \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 ,
         \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 ,
         \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 ,
         \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 ,
         \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 ,
         \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 ,
         \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 ,
         \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 ,
         \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 ,
         \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 ,
         \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 ,
         \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 ,
         \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 ,
         \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 ,
         \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 ,
         \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 ,
         \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 ,
         \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 ,
         \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 ,
         \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 ,
         \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 ,
         \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 ,
         \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 ,
         \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 ,
         \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 ,
         \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 ,
         \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 ,
         \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 ,
         \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 ,
         \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 ,
         \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 ,
         \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 ,
         \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 ,
         \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 ,
         \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 ,
         \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 ,
         \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 ,
         \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 ,
         \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 ,
         \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 ,
         \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 ,
         \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 ,
         \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 ,
         \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 ,
         \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 ,
         \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 ,
         \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 ,
         \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 ,
         \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 ,
         \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 ,
         \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 ,
         \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 ,
         \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 ,
         \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 ,
         \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 ,
         \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 ,
         \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 ,
         \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 ,
         \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 ,
         \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 ,
         \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 ,
         \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 ,
         \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 ,
         \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 ,
         \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 ,
         \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 ,
         \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 ,
         \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 ,
         \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 ,
         \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 ,
         \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 ,
         \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 ,
         \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 ,
         \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 ,
         \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 ,
         \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 ,
         \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 ,
         \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 ,
         \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 ,
         \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 ,
         \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 ,
         \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 ,
         \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 ,
         \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 ,
         \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 ,
         \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 ,
         \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 ,
         \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 ,
         \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 ,
         \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 ,
         \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 ,
         \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 ,
         \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 ,
         \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 ,
         \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 ,
         \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 ,
         \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 ,
         \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 ,
         \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 ,
         \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 ,
         \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 ,
         \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 ,
         \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 ,
         \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 ,
         \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 ,
         \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 ,
         \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 ,
         \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 ,
         \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 ,
         \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 ,
         \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 ,
         \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 ,
         \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 ,
         \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 ,
         \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 ,
         \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 ,
         \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 ,
         \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 ,
         \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 ,
         \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 ,
         \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 ,
         \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 ,
         \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 ,
         \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 ,
         \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 ,
         \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 ,
         \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 ,
         \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 ,
         \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 ,
         \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 ,
         \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 ,
         \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 ,
         \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 ,
         \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 ,
         \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 ,
         \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 ,
         \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 ,
         \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 ,
         \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 ,
         \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 ,
         \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 ,
         \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 ,
         \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 ,
         \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 ,
         \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 ,
         \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 ,
         \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 ,
         \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 ,
         \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 ,
         \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 ,
         \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 ,
         \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 ,
         \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 ,
         \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 ,
         \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 ,
         \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 ,
         \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 ,
         \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 ,
         \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 ,
         \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 ,
         \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 ,
         \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 ,
         \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 ,
         \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 ,
         \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 ,
         \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 ,
         \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 ,
         \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 ,
         \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 ,
         \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 ,
         \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 ,
         \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 ,
         \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 ,
         \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 ,
         \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 ,
         \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 ,
         \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 ,
         \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 ,
         \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 ,
         \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 ,
         \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 ,
         \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 ,
         \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 ,
         \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 ,
         \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 ,
         \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 ,
         \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 ,
         \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 ,
         \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 ,
         \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 ,
         \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 ,
         \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 ,
         \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 ,
         \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 ,
         \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 ,
         \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 ,
         \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 ,
         \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 ,
         \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 ,
         \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 ,
         \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 ,
         \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 ,
         \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 ,
         \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 ,
         \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 ,
         \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 ,
         \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 ,
         \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 ,
         \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 ,
         \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 ,
         \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 ,
         \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 ,
         \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 ,
         \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 ,
         \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 ,
         \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 ,
         \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 ,
         \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 ,
         \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 ,
         \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 ,
         \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 ,
         \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 ,
         \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 ,
         \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 ,
         \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 ,
         \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 ,
         \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 ,
         \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 ,
         \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 ,
         \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 ,
         \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 ,
         \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 ,
         \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 ,
         \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 ,
         \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 ,
         \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 ,
         \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 ,
         \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 ,
         \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 ,
         \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 ,
         \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 ,
         \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 ,
         \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 ,
         \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 ,
         \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 ,
         \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 ,
         \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 ,
         \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 ,
         \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 ,
         \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 ,
         \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 ,
         \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 ,
         \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 ,
         \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 ,
         \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 ,
         \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 ,
         \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 ,
         \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 ,
         \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 ,
         \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 ,
         \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 ,
         \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 ,
         \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 ,
         \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 ,
         \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 ,
         \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 ,
         \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 ,
         \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 ,
         \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 ,
         \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 ,
         \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 ,
         \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 ,
         \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 ,
         \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 ,
         \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 ,
         \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 ,
         \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 ,
         \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 ,
         \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 ,
         \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 ,
         \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 ,
         \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 ,
         \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 ,
         \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 ,
         \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 ,
         \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 ,
         \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 ,
         \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 ,
         \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 ,
         \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 ,
         \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 ,
         \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 ,
         \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 ,
         \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 ,
         \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 ,
         \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 ,
         \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 ,
         \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 ,
         \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 ,
         \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 ,
         \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 ,
         \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 ,
         \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 ,
         \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 ,
         \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 ,
         \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 ,
         \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 ,
         \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 ,
         \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 ,
         \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 ,
         \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 ,
         \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 ,
         \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 ,
         \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 ,
         \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 ,
         \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 ,
         \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 ,
         \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 ,
         \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 ,
         \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 ,
         \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 ,
         \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 ,
         \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 ,
         \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 ,
         \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 ,
         \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 ,
         \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 ,
         \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 ,
         \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 ,
         \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 ,
         \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 ,
         \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 ,
         \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 ,
         \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 ,
         \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 ,
         \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 ,
         \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 ,
         \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 ,
         \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 ,
         \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 ,
         \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 ,
         \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 ,
         \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 ,
         \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 ,
         \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 ,
         \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 ,
         \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 ,
         \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 ,
         \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 ,
         \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 ,
         \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 ,
         \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 ,
         \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 ,
         \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 ,
         \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 ,
         \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 ,
         \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 ,
         \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 ,
         \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 ,
         \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 ,
         \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 ,
         \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 ,
         \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 ,
         \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 ,
         \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 ,
         \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 ,
         \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 ,
         \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 ,
         \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 ,
         \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 ,
         \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 ,
         \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 ,
         \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 ,
         \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 ,
         \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 ,
         \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 ,
         \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 ,
         \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 ,
         \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 ,
         \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 ,
         \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 ,
         \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 ,
         \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 ,
         \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 ,
         \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 ,
         \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 ,
         \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 ,
         \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 ,
         \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 ,
         \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 ,
         \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 ,
         \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 ,
         \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 ,
         \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 ,
         \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 ,
         \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 ,
         \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 ,
         \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 ,
         \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 ,
         \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 ,
         \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 ,
         \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 ,
         \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 ,
         \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 ,
         \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 ,
         \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 ,
         \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 ,
         \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 ,
         \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 ,
         \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 ,
         \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 ,
         \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 ,
         \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 ,
         \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 ,
         \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 ,
         \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 ,
         \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 ,
         \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 ,
         \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 ,
         \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 ,
         \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 ,
         \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 ,
         \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 ,
         \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 ,
         \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 ,
         \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 ,
         \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 ,
         \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 ,
         \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 ,
         \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 ,
         \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 ,
         \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 ,
         \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 ,
         \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 ,
         \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 ,
         \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 ,
         \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 ,
         \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 ,
         \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 ,
         \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 ,
         \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 ,
         \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 ,
         \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 ,
         \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 ,
         \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 ,
         \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 ,
         \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 ,
         \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 ,
         \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 ,
         \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 ,
         \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 ,
         \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 ,
         \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 ,
         \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 ,
         \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 ,
         \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 ,
         \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 ,
         \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 ,
         \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 ,
         \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 ,
         \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 ,
         \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 ,
         \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 ,
         \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 ,
         \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 ,
         \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 ,
         \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 ,
         \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 ,
         \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 ,
         \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 ,
         \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 ,
         \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 ,
         \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 ,
         \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 ,
         \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 ,
         \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 ,
         \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 ,
         \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 ,
         \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 ,
         \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 ,
         \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 ,
         \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 ,
         \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 ,
         \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 ,
         \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 ,
         \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 ,
         \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 ,
         \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 ,
         \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 ,
         \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 ,
         \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 ,
         \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 ,
         \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 ,
         \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 ,
         \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 ,
         \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 ,
         \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 ,
         \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 ,
         \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 ,
         \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 ,
         \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 ,
         \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 ,
         \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 ,
         \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 ,
         \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 ,
         \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 ,
         \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 ,
         \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 ,
         \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 ,
         \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 ,
         \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 ,
         \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 ,
         \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 ,
         \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 ,
         \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 ,
         \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 ,
         \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 ,
         \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 ,
         \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 ,
         \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 ,
         \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 ,
         \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 ,
         \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 ,
         \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 ,
         \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 ,
         \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 ,
         \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 ,
         \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 ,
         \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 ,
         \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 ,
         \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 ,
         \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 ,
         \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 ,
         \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 ,
         \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 ,
         \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 ,
         \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 ,
         \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 ,
         \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 ,
         \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 ,
         \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 ,
         \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 ,
         \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 ,
         \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 ,
         \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 ,
         \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 ,
         \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 ,
         \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 ,
         \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 ,
         \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 ,
         \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 ,
         \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 ,
         \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 ,
         \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 ,
         \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 ,
         \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 ,
         \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 ,
         \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 ,
         \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 ,
         \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 ,
         \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 ,
         \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 ,
         \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 ,
         \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 ,
         \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 ,
         \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 ,
         \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 ,
         \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 ,
         \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 ,
         \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 ,
         \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 ,
         \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 ,
         \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 ,
         \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 ,
         \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 ,
         \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 ,
         \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 ,
         \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 ,
         \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 ,
         \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 ,
         \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 ,
         \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 ,
         \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 ,
         \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 ,
         \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 ,
         \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 ,
         \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 ,
         \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 ,
         \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 ,
         \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 ,
         \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 ,
         \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 ,
         \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 ,
         \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 ,
         \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 ,
         \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 ,
         \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 ,
         \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 ,
         \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 ,
         \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 ,
         \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 ,
         \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 ,
         \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 ,
         \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 ,
         \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 ,
         \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 ,
         \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 ,
         \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 ,
         \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 ,
         \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 ,
         \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 ,
         \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 ,
         \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 ,
         \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 ,
         \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 ,
         \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 ,
         \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 ,
         \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 ,
         \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 ,
         \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 ,
         \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 ,
         \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 ,
         \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 ,
         \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 ,
         \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 ,
         \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 ,
         \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 ,
         \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 ,
         \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 ,
         \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 ,
         \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 ,
         \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 ,
         \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 ,
         \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 ,
         \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 ,
         \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 ,
         \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 ,
         \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 ,
         \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 ,
         \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 ,
         \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 ,
         \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 ,
         \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 ,
         \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 ,
         \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 ,
         \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 ,
         \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 ,
         \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 ,
         \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 ,
         \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 ,
         \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 ,
         \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 ,
         \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 ,
         \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 ,
         \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 ,
         \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 ,
         \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 ,
         \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 ,
         \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 ,
         \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 ,
         \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 ,
         \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 ,
         \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 ,
         \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 ,
         \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 ,
         \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 ,
         \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 ,
         \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 ,
         \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 ,
         \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 ,
         \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 ,
         \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 ,
         \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 ,
         \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 ,
         \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 ,
         \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 ,
         \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 ,
         \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 ,
         \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 ,
         \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 ,
         \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 ,
         \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 ,
         \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 ,
         \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 ,
         \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 ,
         \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 ,
         \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 ,
         \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 ,
         \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 ,
         \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 ,
         \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 ,
         \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 ,
         \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 ,
         \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 ,
         \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 ,
         \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 ,
         \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 ,
         \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 ,
         \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 ,
         \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 ,
         \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 ,
         \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 ,
         \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 ,
         \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 ,
         \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 ,
         \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 ,
         \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 ,
         \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 ,
         \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 ,
         \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 ,
         \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 ,
         \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 ,
         \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 ,
         \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 ,
         \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 ,
         \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 ,
         \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 ,
         \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 ,
         \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 ,
         \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 ,
         \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 ,
         \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 ,
         \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 ,
         \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 ,
         \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 ,
         \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 ,
         \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 ,
         \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 ,
         \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 ,
         \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 ,
         \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 ,
         \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 ,
         \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 ,
         \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 ,
         \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 ,
         \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 ,
         \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 ,
         \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 ,
         \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 ,
         \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 ,
         \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 ,
         \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 ,
         \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 ,
         \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 ,
         \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 ,
         \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 ,
         \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 ,
         \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 ,
         \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 ,
         \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 ,
         \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 ,
         \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 ,
         \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 ,
         \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 ,
         \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 ,
         \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 ,
         \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 ,
         \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 ,
         \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 ,
         \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 ,
         \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 ,
         \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 ,
         \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 ,
         \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 ,
         \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 ,
         \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 ,
         \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 ,
         \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 ,
         \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 ,
         \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 ,
         \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 ,
         \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 ,
         \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 ,
         \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 ,
         \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 ,
         \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 ,
         \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 ,
         \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 ,
         \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 ,
         \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 ,
         \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 ,
         \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 ,
         \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 ,
         \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 ,
         \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 ,
         \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 ,
         \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 ,
         \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 ,
         \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 ,
         \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 ,
         \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 ,
         \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 ,
         \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 ,
         \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 ,
         \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 ,
         \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 ,
         \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 ,
         \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 ,
         \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 ,
         \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 ,
         \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 ,
         \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 ,
         \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 ,
         \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 ,
         \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 ,
         \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 ,
         \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 ,
         \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 ,
         \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 ,
         \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 ,
         \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 ,
         \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 ,
         \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 ,
         \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 ,
         \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 ,
         \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 ,
         \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 ,
         \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 ,
         \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 ,
         \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 ,
         \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 ,
         \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 ,
         \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 ,
         \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 ,
         \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 ,
         \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 ,
         \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 ,
         \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 ,
         \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 ,
         \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 ,
         \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 ,
         \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 ,
         \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 ,
         \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 ,
         \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 ,
         \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 ,
         \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 ,
         \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 ,
         \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 ,
         \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 ,
         \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 ,
         \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 ,
         \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 ,
         \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 ,
         \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 ,
         \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 ,
         \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 ,
         \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 ,
         \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 ,
         \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 ,
         \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 ,
         \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 ,
         \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 ,
         \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 ,
         \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 ,
         \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 ,
         \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 ,
         \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 ,
         \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 ,
         \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 ,
         \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 ,
         \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 ,
         \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 ,
         \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 ,
         \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 ,
         \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 ,
         \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 ,
         \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 ,
         \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 ,
         \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 ,
         \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 , \18033 , \18034 ,
         \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 ,
         \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 ,
         \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 ,
         \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 ,
         \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 ,
         \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 ,
         \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 ,
         \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 ,
         \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 ,
         \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 ,
         \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 ,
         \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 ,
         \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 ,
         \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 ,
         \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 ,
         \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 ,
         \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 ,
         \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 ,
         \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 ,
         \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 ,
         \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 ,
         \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 ,
         \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 ,
         \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 ,
         \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 ,
         \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 ,
         \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 ,
         \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 ,
         \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 ,
         \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 ,
         \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 ,
         \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 ,
         \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 ,
         \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 ,
         \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 ,
         \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 ,
         \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 ,
         \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 ,
         \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 ,
         \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 ,
         \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 ,
         \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 ,
         \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 ,
         \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 ,
         \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 ,
         \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 ,
         \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 ,
         \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 ,
         \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 ,
         \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 ,
         \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 ,
         \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 ,
         \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 ,
         \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 ,
         \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 ,
         \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 ,
         \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 ,
         \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 ,
         \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 ,
         \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 ,
         \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 ,
         \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 ,
         \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 ,
         \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 ,
         \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 ,
         \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 ,
         \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 ,
         \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 ,
         \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 ,
         \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 ,
         \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 ,
         \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 ,
         \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 ,
         \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 ,
         \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 ,
         \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 ,
         \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 ,
         \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 ,
         \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 ,
         \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 ,
         \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 ,
         \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 ,
         \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 ,
         \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 ,
         \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 ,
         \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 ,
         \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 ,
         \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 ,
         \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 ,
         \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 ,
         \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 ,
         \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 ,
         \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 ,
         \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 ,
         \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 ,
         \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 ,
         \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 ,
         \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 ,
         \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 ,
         \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 ,
         \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 ,
         \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 ,
         \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 ,
         \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 ,
         \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 ,
         \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 , \19093 , \19094 ,
         \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 ,
         \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 ,
         \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 ,
         \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 ,
         \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 ,
         \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 ,
         \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 ,
         \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 ,
         \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 ,
         \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 ,
         \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 ,
         \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 ,
         \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 ,
         \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 ,
         \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 ,
         \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 ,
         \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 ,
         \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 ,
         \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 ,
         \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 ,
         \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 ,
         \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 ,
         \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 ,
         \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 ,
         \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 ,
         \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 ,
         \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 ,
         \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 ,
         \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 ,
         \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 ,
         \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 ,
         \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 ,
         \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 ,
         \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 ,
         \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 ,
         \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 ,
         \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 ,
         \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 ,
         \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 ,
         \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 ,
         \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 ,
         \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 ,
         \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 ,
         \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 ,
         \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 ,
         \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 ,
         \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 ,
         \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 ,
         \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 ,
         \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 ,
         \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 ,
         \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 ,
         \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 ,
         \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 ,
         \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 ,
         \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 ,
         \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 ,
         \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 ,
         \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 ,
         \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 ,
         \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 ,
         \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 ,
         \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 ,
         \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 ,
         \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 ,
         \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 ,
         \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 ,
         \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 ,
         \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 ,
         \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 ,
         \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 ,
         \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 ,
         \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 ,
         \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 ,
         \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 ,
         \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 ,
         \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 ,
         \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 ,
         \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 ,
         \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 ,
         \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 ,
         \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 ,
         \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 ,
         \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 ,
         \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 ,
         \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 ,
         \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 ,
         \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 ,
         \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 ,
         \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 ,
         \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 , \20003 , \20004 ,
         \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 ,
         \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 ,
         \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 ,
         \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 ,
         \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 ,
         \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 ,
         \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 ,
         \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 ,
         \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 ,
         \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 ,
         \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 ,
         \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 ,
         \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 ,
         \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 ,
         \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 ,
         \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 ,
         \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 ,
         \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 ,
         \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 ,
         \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 ,
         \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 ,
         \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 ,
         \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 ,
         \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 ,
         \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 ,
         \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 ,
         \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 ,
         \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 ,
         \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 ,
         \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 ,
         \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 ,
         \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 ,
         \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 ,
         \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 ,
         \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 ,
         \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 ,
         \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 ,
         \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 ,
         \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 ,
         \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 ,
         \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 ,
         \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 ,
         \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 ,
         \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 ,
         \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 ,
         \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 ,
         \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 ,
         \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 ,
         \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 ,
         \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 ,
         \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 ,
         \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 ,
         \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 ,
         \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 ,
         \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 ,
         \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 ,
         \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 ,
         \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 ,
         \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 ,
         \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 ,
         \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 ,
         \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 ,
         \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 ,
         \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 ,
         \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 ,
         \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 ,
         \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 ,
         \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 ,
         \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 ,
         \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 ,
         \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 ,
         \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 , \20723 , \20724 ,
         \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 ,
         \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 ,
         \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 ,
         \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 ,
         \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 ,
         \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 ,
         \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 ,
         \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 ,
         \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 ,
         \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 ,
         \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 ,
         \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 ,
         \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 ,
         \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 ,
         \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 ,
         \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 ,
         \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 ,
         \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 ,
         \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 ,
         \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 ,
         \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 ,
         \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 ,
         \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 ,
         \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 ,
         \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 ,
         \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 ,
         \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 ,
         \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 ,
         \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 ,
         \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 ,
         \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 ,
         \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 ,
         \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 ,
         \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 ,
         \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 ,
         \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 ,
         \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 ,
         \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 ,
         \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 ,
         \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 ,
         \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 ,
         \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 ,
         \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 ,
         \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 ,
         \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 ,
         \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 ,
         \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 ,
         \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 ,
         \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 ,
         \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 ,
         \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 ,
         \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 ,
         \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 ,
         \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 ,
         \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 ,
         \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 ,
         \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 ,
         \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 ,
         \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 ,
         \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 ,
         \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 ,
         \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 ,
         \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 ,
         \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 ,
         \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 ,
         \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 ,
         \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 ,
         \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 ,
         \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 ,
         \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 ,
         \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 ,
         \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 ,
         \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 ,
         \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 ,
         \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 ,
         \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 ,
         \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 ,
         \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 ,
         \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 ,
         \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 ,
         \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 ,
         \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 ,
         \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 ,
         \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 ,
         \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 ,
         \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 ,
         \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 ,
         \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 ,
         \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 ,
         \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 ,
         \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 ,
         \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 ,
         \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 , \21653 , \21654 ,
         \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 ,
         \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 ,
         \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 ,
         \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 ,
         \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 ,
         \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 ,
         \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 ,
         \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 ,
         \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 ,
         \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 ,
         \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 ,
         \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 ,
         \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 ,
         \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 ,
         \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 ,
         \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 ,
         \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 ,
         \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 ,
         \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 ,
         \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 ,
         \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 ,
         \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 ,
         \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 ,
         \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 ,
         \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 ,
         \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 ,
         \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 ,
         \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 ,
         \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 ,
         \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 ,
         \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 ,
         \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 ,
         \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 ,
         \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 ,
         \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 ,
         \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 ,
         \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 ,
         \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 ,
         \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 ,
         \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 ,
         \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 ,
         \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 , \22073 , \22074 ,
         \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 ,
         \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 , \22093 , \22094 ,
         \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 , \22103 , \22104 ,
         \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 , \22113 , \22114 ,
         \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 , \22123 , \22124 ,
         \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 , \22133 , \22134 ,
         \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 ,
         \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 , \22153 , \22154 ,
         \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , \22163 , \22164 ,
         \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 , \22173 , \22174 ,
         \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 , \22183 , \22184 ,
         \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , \22193 , \22194 ,
         \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 ,
         \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 , \22213 , \22214 ,
         \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , \22223 , \22224 ,
         \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 ,
         \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 , \22243 , \22244 ,
         \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 ,
         \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 , \22263 , \22264 ,
         \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 , \22273 , \22274 ,
         \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 ,
         \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 ,
         \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 , \22303 , \22304 ,
         \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 ,
         \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 ,
         \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 , \22333 , \22334 ,
         \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 ,
         \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 , \22353 , \22354 ,
         \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 , \22363 , \22364 ,
         \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 , \22373 , \22374 ,
         \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 ,
         \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 ,
         \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 ,
         \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 , \22413 , \22414 ,
         \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 ,
         \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 ,
         \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 ,
         \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 ,
         \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 ,
         \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 , \22473 , \22474 ,
         \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 ,
         \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 , \22493 , \22494 ,
         \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 ,
         \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 ,
         \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 ,
         \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 ,
         \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 ,
         \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 , \22553 , \22554 ,
         \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 ,
         \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 , \22573 , \22574 ,
         \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 ,
         \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 , \22593 , \22594 ,
         \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 , \22603 , \22604 ,
         \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 , \22613 , \22614 ,
         \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 ,
         \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 , \22633 , \22634 ,
         \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 ,
         \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653 , \22654 ,
         \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 ,
         \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 ,
         \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 ,
         \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 ,
         \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 ,
         \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 , \22714 ,
         \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 ,
         \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 ,
         \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 ,
         \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 ,
         \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 ,
         \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 ,
         \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 , \22783 , \22784 ,
         \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 ,
         \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 ,
         \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 ,
         \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 ,
         \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 ,
         \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 ,
         \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 ,
         \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 ,
         \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 ,
         \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 ,
         \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 ,
         \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 ,
         \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914 ,
         \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 ,
         \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 ,
         \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 ,
         \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 ,
         \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 ,
         \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 ,
         \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 ,
         \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 ,
         \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 ,
         \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 ,
         \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 ,
         \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 ,
         \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 ,
         \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 ,
         \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 ,
         \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 ,
         \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 ,
         \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 ,
         \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 ,
         \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 , \23114 ,
         \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 ,
         \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 ,
         \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 ,
         \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 ,
         \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 ,
         \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 ,
         \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 , \23183 , \23184 ,
         \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 , \23193 , \23194 ,
         \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 ,
         \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 ,
         \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 , \23223 , \23224 ,
         \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 ,
         \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 ,
         \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 ,
         \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 ,
         \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 , \23274 ,
         \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 ,
         \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 ,
         \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 , \23303 , \23304 ,
         \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 ,
         \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 ,
         \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 , \23333 , \23334 ,
         \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 ,
         \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 ,
         \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 ,
         \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 ,
         \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 ,
         \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 ,
         \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 ,
         \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 ,
         \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 ,
         \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 ,
         \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 ,
         \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 , \23453 , \23454 ,
         \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 ,
         \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 , \23473 , \23474 ,
         \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483 , \23484 ,
         \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 , \23493 , \23494 ,
         \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 ,
         \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 , \23514 ,
         \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 ,
         \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 ,
         \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 ,
         \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 ,
         \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 , \23563 , \23564 ,
         \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 ,
         \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 ,
         \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 ,
         \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 ,
         \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 ,
         \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 , \23623 , \23624 ,
         \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 ,
         \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643 , \23644 ,
         \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 ,
         \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 , \23663 , \23664 ,
         \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 , \23673 , \23674 ,
         \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 , \23683 , \23684 ,
         \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 ,
         \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 , \23703 , \23704 ,
         \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 ,
         \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 ,
         \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 ,
         \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 ,
         \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753 , \23754 ,
         \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 ,
         \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 , \23773 , \23774 ,
         \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 , \23783 , \23784 ,
         \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 , \23793 , \23794 ,
         \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 ,
         \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 , \23813 , \23814 ,
         \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 ,
         \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 ,
         \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844 ,
         \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 ,
         \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 , \23863 , \23864 ,
         \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 ,
         \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 ,
         \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 ,
         \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 ,
         \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 ,
         \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 ,
         \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934 ,
         \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 ,
         \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 ,
         \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 ,
         \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 , \23973 , \23974 ,
         \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 ,
         \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 ,
         \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 , \24003 , \24004 ,
         \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 ,
         \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 ,
         \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 ,
         \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 ,
         \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 ,
         \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24064 ,
         \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 ,
         \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 ,
         \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 ,
         \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 ,
         \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 ,
         \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 ,
         \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133 , \24134 ,
         \24135 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 , \24143 , \24144 ,
         \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153 , \24154 ,
         \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 , \24163 , \24164 ,
         \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173 , \24174 ,
         \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 , \24183 , \24184 ,
         \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 , \24193 , \24194 ,
         \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 ,
         \24205 , \24206 , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 , \24213 , \24214 ,
         \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 ,
         \24225 , \24226 , \24227 , \24228 , \24229 , \24230 , \24231 , \24232 , \24233 , \24234 ,
         \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 , \24243 , \24244 ,
         \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 ,
         \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263 , \24264 ,
         \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 ,
         \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 , \24283 , \24284 ,
         \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 ,
         \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 , \24303 , \24304 ,
         \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 ,
         \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 ,
         \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333 , \24334 ,
         \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 ,
         \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 , \24353 , \24354 ,
         \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 ,
         \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 , \24373 , \24374 ,
         \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 , \24383 , \24384 ,
         \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 ,
         \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 ,
         \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413 , \24414 ,
         \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 ,
         \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 , \24433 , \24434 ,
         \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 ,
         \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 ,
         \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 , \24463 , \24464 ,
         \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 ,
         \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 , \24483 , \24484 ,
         \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494 ,
         \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 ,
         \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 , \24513 , \24514 ,
         \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 ,
         \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534 ,
         \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 , \24543 , \24544 ,
         \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 ,
         \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 ,
         \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 , \24573 , \24574 ,
         \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 ,
         \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 ,
         \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 ,
         \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 ,
         \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 ,
         \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 ,
         \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 , \24643 , \24644 ,
         \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 ,
         \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 ,
         \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 ,
         \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 ,
         \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 , \24693 , \24694 ,
         \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 ,
         \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 ,
         \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 ,
         \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 ,
         \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 ,
         \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 ,
         \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 ,
         \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 , \24773 , \24774 ,
         \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 , \24783 , \24784 ,
         \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 ,
         \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 , \24803 , \24804 ,
         \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 ,
         \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 ,
         \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834 ,
         \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 ,
         \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 , \24853 , \24854 ,
         \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 ,
         \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 ,
         \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 , \24883 , \24884 ,
         \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 ,
         \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 , \24903 , \24904 ,
         \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 ,
         \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 , \24923 , \24924 ,
         \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 , \24934 ,
         \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 ,
         \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954 ,
         \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 , \24963 , \24964 ,
         \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 , \24973 , \24974 ,
         \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 ,
         \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 , \24993 , \24994 ,
         \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 ,
         \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 ,
         \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 , \25023 , \25024 ,
         \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 ,
         \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 ,
         \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 ,
         \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 ,
         \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 ,
         \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 ,
         \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 , \25093 , \25094 ,
         \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 ,
         \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 ,
         \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124 ,
         \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 , \25133 , \25134 ,
         \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 ,
         \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 ,
         \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 ,
         \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 ,
         \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 ,
         \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 , \25194 ,
         \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 ,
         \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 ,
         \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 ,
         \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 ,
         \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 ,
         \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 ,
         \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 , \25263 , \25264 ,
         \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 , \25273 , \25274 ,
         \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 , \25283 , \25284 ,
         \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294 ,
         \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 ,
         \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 , \25313 , \25314 ,
         \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 ,
         \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 ,
         \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 ,
         \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 ,
         \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 , \25363 , \25364 ,
         \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 ,
         \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 , \25383 , \25384 ,
         \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 , \25393 , \25394 ,
         \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 ,
         \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413 , \25414 ,
         \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 , \25423 , \25424 ,
         \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 , \25433 , \25434 ,
         \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 ,
         \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 ,
         \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 ,
         \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 , \25473 , \25474 ,
         \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 , \25483 , \25484 ,
         \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 ,
         \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 , \25503 , \25504 ,
         \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 ,
         \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 ,
         \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533 , \25534 ,
         \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 ,
         \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 ,
         \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 ,
         \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 ,
         \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 ,
         \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 ,
         \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 , \25603 , \25604 ,
         \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 ,
         \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 ,
         \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 , \25634 ,
         \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 ,
         \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653 , \25654 ,
         \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 ,
         \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 , \25673 , \25674 ,
         \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 ,
         \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 , \25693 , \25694 ,
         \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704 ,
         \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713 , \25714 ,
         \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 ,
         \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 ,
         \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 ,
         \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 ,
         \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 ,
         \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 , \25773 , \25774 ,
         \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 , \25783 , \25784 ,
         \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 , \25793 , \25794 ,
         \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 ,
         \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 , \25813 , \25814 ,
         \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 ,
         \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 ,
         \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843 , \25844 ,
         \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 ,
         \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 , \25863 , \25864 ,
         \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 , \25873 , \25874 ,
         \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 ,
         \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 ,
         \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 , \25903 , \25904 ,
         \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 ,
         \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 ,
         \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 ,
         \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 , \25944 ,
         \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 ,
         \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 ,
         \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 ,
         \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984 ,
         \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 ,
         \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 ,
         \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 , \26013 , \26014 ,
         \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 ,
         \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 ,
         \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 ,
         \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 ,
         \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 ,
         \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 ,
         \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 ,
         \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 ,
         \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 ,
         \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 , \26114 ,
         \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 ,
         \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 ,
         \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 , \26143 , \26144 ,
         \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 ,
         \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 ,
         \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 ,
         \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 ,
         \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 ,
         \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 ,
         \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 , \26213 , \26214 ,
         \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 ,
         \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 ,
         \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 ,
         \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 ,
         \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 ,
         \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273 , \26274 ,
         \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 , \26283 , \26284 ,
         \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294 ,
         \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 ,
         \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 ,
         \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 , \26323 , \26324 ,
         \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 ,
         \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 , \26343 , \26344 ,
         \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 ,
         \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 , \26363 , \26364 ,
         \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 ,
         \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 , \26383 , \26384 ,
         \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 ,
         \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404 ,
         \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 , \26413 , \26414 ,
         \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 , \26423 , \26424 ,
         \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 , \26433 , \26434 ,
         \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 , \26443 , \26444 ,
         \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 , \26453 , \26454 ,
         \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 , \26463 , \26464 ,
         \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 , \26473 , \26474 ,
         \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 , \26483 , \26484 ,
         \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 , \26493 , \26494 ,
         \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 , \26503 , \26504 ,
         \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 ,
         \26515 , \26516 , \26517 , \26518 , \26519 , \26520 , \26521 , \26522 , \26523 , \26524 ,
         \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 , \26533 , \26534 ,
         \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 ,
         \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 , \26553 , \26554 ,
         \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 ,
         \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574 ,
         \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584 ,
         \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 ,
         \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 , \26603 , \26604 ,
         \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 ,
         \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 ,
         \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , \26634 ,
         \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644 ,
         \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654 ,
         \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 ,
         \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 , \26673 , \26674 ,
         \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 ,
         \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 ,
         \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704 ,
         \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 ,
         \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 , \26723 , \26724 ,
         \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 ,
         \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 ,
         \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 ,
         \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763 , \26764 ,
         \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 , \26773 , \26774 ,
         \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 , \26783 , \26784 ,
         \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 ,
         \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804 ,
         \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 , \26813 , \26814 ,
         \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 , \26823 , \26824 ,
         \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 ,
         \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 , \26843 , \26844 ,
         \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 , \26853 , \26854 ,
         \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 ,
         \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 , \26873 , \26874 ,
         \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 , \26883 , \26884 ,
         \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 ,
         \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 , \26903 , \26904 ,
         \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 ,
         \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 ,
         \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 , \26933 , \26934 ,
         \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 ,
         \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 ,
         \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 , \26963 , \26964 ,
         \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 ,
         \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 ,
         \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 , \26993 , \26994 ,
         \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 ,
         \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 , \27013 , \27014 ,
         \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 , \27023 , \27024 ,
         \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 ,
         \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 ,
         \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 ,
         \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 ,
         \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 ,
         \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 ,
         \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 , \27094 ,
         \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 ,
         \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 ,
         \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 ,
         \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 ,
         \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 ,
         \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 ,
         \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 ,
         \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 ,
         \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 ,
         \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 ,
         \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 ,
         \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 ,
         \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 ,
         \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 ,
         \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 ,
         \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 ,
         \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 ,
         \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 ,
         \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 ,
         \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 , \27293 , \27294 ,
         \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 , \27303 , \27304 ,
         \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 , \27313 , \27314 ,
         \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 ,
         \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 ,
         \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344 ,
         \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 ,
         \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 , \27363 , \27364 ,
         \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 ,
         \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 ,
         \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 , \27393 , \27394 ,
         \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 ,
         \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 , \27413 , \27414 ,
         \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 ,
         \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 ,
         \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 , \27443 , \27444 ,
         \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 ,
         \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 ,
         \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 , \27473 , \27474 ,
         \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 ,
         \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 ,
         \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 ,
         \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 ,
         \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 , \27523 , \27524 ,
         \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 ,
         \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 ,
         \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 , \27553 , \27554 ,
         \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 ,
         \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 ,
         \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 ,
         \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 ,
         \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 ,
         \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 ,
         \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 ,
         \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 , \27633 , \27634 ,
         \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 ,
         \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 ,
         \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 ,
         \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 ,
         \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 ,
         \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 ,
         \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 ,
         \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714 ,
         \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 ,
         \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 ,
         \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 ,
         \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 ,
         \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 ,
         \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 ,
         \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 ,
         \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 ,
         \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 ,
         \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 , \27813 , \27814 ,
         \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 ,
         \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 , \27833 , \27834 ,
         \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 , \27843 , \27844 ,
         \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 ,
         \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 , \27863 , \27864 ,
         \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 ,
         \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883 , \27884 ,
         \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 ,
         \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 , \27903 , \27904 ,
         \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 ,
         \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 ,
         \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 ,
         \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 ,
         \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 , \27953 , \27954 ,
         \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 , \27963 , \27964 ,
         \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 , \27973 , \27974 ,
         \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 ,
         \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 ,
         \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 ,
         \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 ,
         \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 ,
         \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 , \28033 , \28034 ,
         \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 ,
         \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 ,
         \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 ,
         \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 ,
         \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 ,
         \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 ,
         \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 ,
         \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 , \28113 , \28114 ,
         \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 ,
         \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133 , \28134 ,
         \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 , \28143 , \28144 ,
         \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 , \28153 , \28154 ,
         \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 ,
         \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 , \28173 , \28174 ,
         \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 ,
         \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 , \28193 , \28194 ,
         \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 ,
         \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 , \28213 , \28214 ,
         \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 , \28223 , \28224 ,
         \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 ,
         \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 ,
         \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 ,
         \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 ,
         \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 ,
         \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 ,
         \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 ,
         \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 ,
         \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 ,
         \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324 ,
         \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 ,
         \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 ,
         \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 ,
         \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 ,
         \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 ,
         \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 , \28383 , \28384 ,
         \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 , \28393 , \28394 ,
         \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 ,
         \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 ,
         \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 ,
         \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 ,
         \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 ,
         \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 ,
         \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 ,
         \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 ,
         \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 , \28483 , \28484 ,
         \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 ,
         \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 ,
         \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 ,
         \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 , \28523 , \28524 ,
         \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 , \28533 , \28534 ,
         \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 , \28543 , \28544 ,
         \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 , \28553 , \28554 ,
         \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 , \28563 , \28564 ,
         \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 , \28573 , \28574 ,
         \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 , \28583 , \28584 ,
         \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 ,
         \28595 , \28596 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 , \28603 , \28604 ,
         \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 ,
         \28615 , \28616 , \28617 , \28618 , \28619 , \28620 , \28621 , \28622 , \28623 , \28624 ,
         \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 ,
         \28635 , \28636 , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 , \28643 , \28644 ,
         \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 , \28653 , \28654 ,
         \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 , \28663 , \28664 ,
         \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 , \28673 , \28674 ,
         \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 , \28683 , \28684 ,
         \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 , \28693 , \28694 ,
         \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 , \28703 , \28704 ,
         \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 , \28713 , \28714 ,
         \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 , \28723 , \28724 ,
         \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 ,
         \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 , \28743 , \28744 ,
         \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 , \28753 , \28754 ,
         \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 ,
         \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771 , \28772 , \28773 , \28774 ,
         \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 ,
         \28785 , \28786 , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 , \28793 , \28794 ,
         \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804 ,
         \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 ,
         \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , \28824 ,
         \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 ,
         \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 , \28843 , \28844 ,
         \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 ,
         \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 , \28863 , \28864 ,
         \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 ,
         \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 , \28883 , \28884 ,
         \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 ,
         \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904 ,
         \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 ,
         \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 , \28923 , \28924 ,
         \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , \28933 , \28934 ,
         \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 ,
         \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 , \28953 , \28954 ,
         \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 ,
         \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 , \28973 , \28974 ,
         \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 ,
         \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 ,
         \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 ,
         \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014 ,
         \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 , \29023 , \29024 ,
         \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 ,
         \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 ,
         \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 ,
         \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 , \29063 , \29064 ,
         \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 ,
         \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 , \29083 , \29084 ,
         \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094 ,
         \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 ,
         \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 , \29113 , \29114 ,
         \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 ,
         \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 , \29133 , \29134 ,
         \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 , \29143 , \29144 ,
         \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 ,
         \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 ,
         \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 ,
         \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 , \29183 , \29184 ,
         \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 , \29193 , \29194 ,
         \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 , \29203 , \29204 ,
         \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 ,
         \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 , \29223 , \29224 ,
         \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 ,
         \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 ,
         \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 ,
         \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 ,
         \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 , \29274 ,
         \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 ,
         \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 , \29293 , \29294 ,
         \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 , \29303 , \29304 ,
         \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 ,
         \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 ,
         \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 ,
         \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 ,
         \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 ,
         \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 ,
         \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 ,
         \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 ,
         \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 ,
         \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 ,
         \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 , \29413 , \29414 ,
         \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 ,
         \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433 , \29434 ,
         \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 ,
         \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 ,
         \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 , \29463 , \29464 ,
         \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 ,
         \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 ,
         \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 ,
         \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 , \29503 , \29504 ,
         \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 ,
         \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 ,
         \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533 , \29534 ,
         \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 , \29543 , \29544 ,
         \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 ,
         \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 ,
         \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 , \29573 , \29574 ,
         \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 ,
         \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 ,
         \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 ,
         \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 ,
         \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624 ,
         \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 ,
         \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 ,
         \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 ,
         \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 ,
         \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 ,
         \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 ,
         \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 ,
         \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 , \29703 , \29704 ,
         \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 ,
         \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 ,
         \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 , \29733 , \29734 ,
         \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 ,
         \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 ,
         \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 ,
         \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 ,
         \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 ,
         \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 ,
         \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 ,
         \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 ,
         \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 ,
         \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833 , \29834 ,
         \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 , \29843 , \29844 ,
         \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 ,
         \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 ,
         \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873 , \29874 ,
         \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 ,
         \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 , \29893 , \29894 ,
         \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 ,
         \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 , \29913 , \29914 ,
         \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 , \29923 , \29924 ,
         \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 ,
         \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 ,
         \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 ,
         \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 , \29963 , \29964 ,
         \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 , \29974 ,
         \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 , \29983 , \29984 ,
         \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 ,
         \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 ,
         \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 ,
         \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 ,
         \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 ,
         \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 , \30044 ,
         \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 , \30053 , \30054 ,
         \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 ,
         \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073 , \30074 ,
         \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 ,
         \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 ,
         \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 ,
         \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 , \30113 , \30114 ,
         \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 ,
         \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 ,
         \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 , \30143 , \30144 ,
         \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 ,
         \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 , \30163 , \30164 ,
         \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 ,
         \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 , \30183 , \30184 ,
         \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 ,
         \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 ,
         \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 , \30213 , \30214 ,
         \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 ,
         \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 ,
         \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 , \30243 , \30244 ,
         \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 ,
         \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263 , \30264 ,
         \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 ,
         \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 , \30283 , \30284 ,
         \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 , \30293 , \30294 ,
         \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 ,
         \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314 ,
         \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 , \30323 , \30324 ,
         \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 , \30333 , \30334 ,
         \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 ,
         \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 ,
         \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 ,
         \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 , \30373 , \30374 ,
         \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 , \30383 , \30384 ,
         \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 ,
         \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 , \30403 , \30404 ,
         \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 ,
         \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 ,
         \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 , \30433 , \30434 ,
         \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 ,
         \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 , \30454 ,
         \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463 , \30464 ,
         \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 ,
         \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 , \30483 , \30484 ,
         \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 ,
         \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 ,
         \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 , \30513 , \30514 ,
         \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 ,
         \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 , \30533 , \30534 ,
         \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 ,
         \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 ,
         \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564 ,
         \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 ,
         \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 ,
         \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 ,
         \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 , \30603 , \30604 ,
         \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 ,
         \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 ,
         \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 ,
         \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 ,
         \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 ,
         \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 ,
         \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 ,
         \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 ,
         \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 ,
         \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 ,
         \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 ,
         \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 , \30723 , \30724 ,
         \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 ,
         \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 , \30743 , \30744 ,
         \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 ,
         \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764 ,
         \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 ,
         \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 ,
         \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 ,
         \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 , \30803 , \30804 ,
         \30805 , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 , \30813 , \30814 ,
         \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 , \30823 , \30824 ,
         \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 , \30833 , \30834 ,
         \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 , \30843 , \30844 ,
         \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 , \30853 , \30854 ,
         \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 ,
         \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 , \30873 , \30874 ,
         \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 , \30883 , \30884 ,
         \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892 , \30893 , \30894 ,
         \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 , \30903 , \30904 ,
         \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 , \30913 , \30914 ,
         \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 , \30923 , \30924 ,
         \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 , \30933 , \30934 ,
         \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 , \30943 , \30944 ,
         \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952 , \30953 , \30954 ,
         \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 ,
         \30965 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 , \30973 , \30974 ,
         \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 , \30983 , \30984 ,
         \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 , \30993 , \30994 ,
         \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 ,
         \31005 , \31006 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 , \31013 , \31014 ,
         \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023 , \31024 ,
         \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 , \31033 , \31034 ,
         \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 , \31043 , \31044 ,
         \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 , \31053 , \31054 ,
         \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 , \31063 , \31064 ,
         \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 ,
         \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082 , \31083 , \31084 ,
         \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 ,
         \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 , \31103 , \31104 ,
         \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 ,
         \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 , \31123 , \31124 ,
         \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 ,
         \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 , \31143 , \31144 ,
         \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 , \31153 , \31154 ,
         \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 , \31163 , \31164 ,
         \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 ,
         \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 ,
         \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 ,
         \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 ,
         \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 ,
         \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 , \31223 , \31224 ,
         \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 ,
         \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 ,
         \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , \31253 , \31254 ,
         \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 , \31263 , \31264 ,
         \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 ,
         \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 ,
         \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 ,
         \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 ,
         \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 ,
         \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 ,
         \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333 , \31334 ,
         \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 ,
         \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 , \31353 , \31354 ,
         \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 , \31363 , \31364 ,
         \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 ,
         \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 ,
         \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 ,
         \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 ,
         \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 ,
         \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 ,
         \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 ,
         \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 ,
         \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 ,
         \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 ,
         \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474 ,
         \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483 , \31484 ,
         \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 ,
         \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 ,
         \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 ,
         \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 ,
         \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 ,
         \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 ,
         \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 , \31553 , \31554 ,
         \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 ,
         \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 ,
         \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 ,
         \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 ,
         \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 , \31603 , \31604 ,
         \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614 ,
         \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 ,
         \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 , \31633 , \31634 ,
         \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 , \31643 , \31644 ,
         \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 ,
         \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 ,
         \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 , \31673 , \31674 ,
         \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 , \31684 ,
         \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 ,
         \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 ,
         \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 , \31713 , \31714 ,
         \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 ,
         \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 ,
         \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 , \31743 , \31744 ,
         \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 , \31753 , \31754 ,
         \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 ,
         \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 ,
         \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 , \31783 , \31784 ,
         \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 , \31793 , \31794 ,
         \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 ,
         \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 ,
         \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 ,
         \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 ,
         \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 ,
         \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 ,
         \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 ,
         \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 ,
         \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 ,
         \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 ,
         \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 ,
         \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 ,
         \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 , \31923 , \31924 ,
         \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 ,
         \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 ,
         \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 ,
         \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 ,
         \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 ,
         \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 ,
         \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 ,
         \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 ,
         \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 ,
         \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 ,
         \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 , \32033 , \32034 ,
         \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 ,
         \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 , \32053 , \32054 ,
         \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 , \32063 , \32064 ,
         \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 ,
         \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 ,
         \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 , \32093 , \32094 ,
         \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 ,
         \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 , \32114 ,
         \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 , \32123 , \32124 ,
         \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 ,
         \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 , \32143 , \32144 ,
         \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 , \32153 , \32154 ,
         \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 ,
         \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 , \32173 , \32174 ,
         \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 , \32183 , \32184 ,
         \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 ,
         \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 ,
         \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 , \32213 , \32214 ,
         \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 , \32223 , \32224 ,
         \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 ,
         \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 , \32243 , \32244 ,
         \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 ,
         \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 , \32263 , \32264 ,
         \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 , \32273 , \32274 ,
         \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 ,
         \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 , \32293 , \32294 ,
         \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302 , \32303 , \32304 ,
         \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314 ,
         \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 , \32323 , \32324 ,
         \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 ,
         \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 , \32343 , \32344 ,
         \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 ,
         \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 , \32364 ,
         \32365 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 , \32373 , \32374 ,
         \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 ,
         \32385 , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 , \32393 , \32394 ,
         \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 ,
         \32405 , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 , \32413 , \32414 ,
         \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 ,
         \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 , \32433 , \32434 ,
         \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 ,
         \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 , \32453 , \32454 ,
         \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 , \32463 , \32464 ,
         \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 ,
         \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 ,
         \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 ,
         \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 ,
         \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 , \32513 , \32514 ,
         \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 ,
         \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 ,
         \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 ,
         \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 ,
         \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 ,
         \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 ,
         \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 ,
         \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 , \32594 ,
         \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 ,
         \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 ,
         \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 ,
         \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 ,
         \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 ,
         \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 ,
         \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 , \32663 , \32664 ,
         \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 ,
         \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 ,
         \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 ,
         \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704 ,
         \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 ,
         \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 ,
         \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733 , \32734 ,
         \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 ,
         \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 ,
         \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 ,
         \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 ,
         \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 ,
         \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 , \32793 , \32794 ,
         \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 , \32803 , \32804 ,
         \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 , \32813 , \32814 ,
         \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 , \32823 , \32824 ,
         \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 ,
         \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 , \32843 , \32844 ,
         \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 ,
         \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 , \32863 , \32864 ,
         \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 ,
         \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884 ,
         \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 , \32893 , \32894 ,
         \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 ,
         \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 ,
         \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924 ,
         \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 , \32933 , \32934 ,
         \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944 ,
         \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 ,
         \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 , \32963 , \32964 ,
         \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 , \32973 , \32974 ,
         \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984 ,
         \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 , \32993 , \32994 ,
         \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004 ,
         \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 , \33013 , \33014 ,
         \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024 ,
         \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 , \33033 , \33034 ,
         \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 , \33043 , \33044 ,
         \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 ,
         \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 , \33063 , \33064 ,
         \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 ,
         \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081 , \33082 , \33083 , \33084 ,
         \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 ,
         \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101 , \33102 , \33103 , \33104 ,
         \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 ,
         \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122 , \33123 , \33124 ,
         \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 , \33133 , \33134 ,
         \33135 , \33136 , \33137 , \33138 , \33139 , \33140 , \33141 , \33142 , \33143 , \33144 ,
         \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 , \33153 , \33154 ,
         \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 , \33163 , \33164 ,
         \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 , \33173 , \33174 ,
         \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 , \33183 , \33184 ,
         \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 , \33193 , \33194 ,
         \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 , \33203 , \33204 ,
         \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 ,
         \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , \33223 , \33224 ,
         \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 ,
         \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 , \33243 , \33244 ,
         \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 ,
         \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 , \33263 , \33264 ,
         \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 ,
         \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 , \33283 , \33284 ,
         \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294 ,
         \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 , \33303 , \33304 ,
         \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 ,
         \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 , \33323 , \33324 ,
         \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334 ,
         \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 , \33343 , \33344 ,
         \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354 ,
         \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 , \33363 , \33364 ,
         \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 , \33373 , \33374 ,
         \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , \33384 ,
         \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 , \33393 , \33394 ,
         \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , \33403 , \33404 ,
         \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 , \33413 , \33414 ,
         \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , \33423 , \33424 ,
         \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 , \33433 , \33434 ,
         \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , \33443 , \33444 ,
         \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 , \33453 , \33454 ,
         \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , \33463 , \33464 ,
         \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 , \33473 , \33474 ,
         \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , \33483 , \33484 ,
         \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 ,
         \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , \33503 , \33504 ,
         \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 ,
         \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , \33523 , \33524 ,
         \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532 , \33533 , \33534 ,
         \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 , \33543 , \33544 ,
         \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 ,
         \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 ,
         \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 , \33573 , \33574 ,
         \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 ,
         \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 ,
         \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 , \33603 , \33604 ,
         \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613 , \33614 ,
         \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 , \33623 , \33624 ,
         \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 , \33633 , \33634 ,
         \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 , \33643 , \33644 ,
         \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 ,
         \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 , \33663 , \33664 ,
         \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 ,
         \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 , \33683 , \33684 ,
         \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 ,
         \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 , \33703 , \33704 ,
         \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 , \33713 , \33714 ,
         \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 , \33723 , \33724 ,
         \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 ,
         \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 , \33743 , \33744 ,
         \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 ,
         \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 ,
         \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 ,
         \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 ,
         \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 , \33793 , \33794 ,
         \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 ,
         \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 ,
         \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 , \33823 , \33824 ,
         \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834 ,
         \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 ,
         \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853 , \33854 ,
         \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 ,
         \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 , \33873 , \33874 ,
         \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 ,
         \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 , \33893 , \33894 ,
         \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 , \33903 , \33904 ,
         \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 , \33913 , \33914 ,
         \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 ,
         \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 , \33933 , \33934 ,
         \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 ,
         \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 , \33953 , \33954 ,
         \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 ,
         \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 ,
         \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 , \33983 , \33984 ,
         \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 ,
         \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004 ,
         \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 ,
         \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 , \34023 , \34024 ,
         \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 ,
         \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 , \34043 , \34044 ,
         \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 , \34053 , \34054 ,
         \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061 , \34062 , \34063 , \34064 ,
         \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 ,
         \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 , \34083 , \34084 ,
         \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 ,
         \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 , \34103 , \34104 ,
         \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 , \34114 ,
         \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 ,
         \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 ,
         \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 , \34143 , \34144 ,
         \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153 , \34154 ,
         \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 ,
         \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 , \34173 , \34174 ,
         \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 ,
         \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 , \34193 , \34194 ,
         \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 ,
         \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 ,
         \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 , \34223 , \34224 ,
         \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 ,
         \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243 , \34244 ,
         \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 , \34253 , \34254 ,
         \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 , \34263 , \34264 ,
         \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 ,
         \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 , \34283 , \34284 ,
         \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294 ,
         \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 , \34303 , \34304 ,
         \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 ,
         \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 ,
         \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 , \34333 , \34334 ,
         \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 ,
         \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353 , \34354 ,
         \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 ,
         \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 , \34373 , \34374 ,
         \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 , \34384 ,
         \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 , \34393 , \34394 ,
         \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 ,
         \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 , \34413 , \34414 ,
         \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 ,
         \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 ,
         \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 , \34443 , \34444 ,
         \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 ,
         \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 , \34463 , \34464 ,
         \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 ,
         \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 , \34483 , \34484 ,
         \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 , \34493 , \34494 ,
         \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 ,
         \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 ,
         \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 ,
         \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 , \34533 , \34534 ,
         \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 ,
         \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 , \34553 , \34554 ,
         \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 , \34563 , \34564 ,
         \34565 , \34566 , \34567 , \34568 , \34569 , \34570 , \34571 , \34572 , \34573 , \34574 ,
         \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 ,
         \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591 , \34592 , \34593 , \34594 ,
         \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 ,
         \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 , \34613 , \34614 ,
         \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623 , \34624 ,
         \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 , \34634 ,
         \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 , \34643 , \34644 ,
         \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 ,
         \34655 , \34656 , \34657 , \34658 , \34659 , \34660 , \34661 , \34662 , \34663 , \34664 ,
         \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 ,
         \34675 , \34676 , \34677 , \34678 , \34679 , \34680 , \34681 , \34682 , \34683 , \34684 ,
         \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 ,
         \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 , \34703 , \34704 ,
         \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 ,
         \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 , \34723 , \34724 ,
         \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 , \34733 , \34734 ,
         \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 ,
         \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 , \34753 , \34754 ,
         \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 ,
         \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 , \34773 , \34774 ,
         \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 , \34783 , \34784 ,
         \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 ,
         \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 ,
         \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 , \34813 , \34814 ,
         \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823 , \34824 ,
         \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 ,
         \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 , \34843 , \34844 ,
         \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 ,
         \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 , \34863 , \34864 ,
         \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 ,
         \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 ,
         \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 , \34893 , \34894 ,
         \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 ,
         \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913 , \34914 ,
         \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 , \34923 , \34924 ,
         \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933 , \34934 ,
         \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 ,
         \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 , \34953 , \34954 ,
         \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 ,
         \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 , \34973 , \34974 ,
         \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 ,
         \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 ,
         \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 , \35003 , \35004 ,
         \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 ,
         \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023 , \35024 ,
         \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 ,
         \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 , \35043 , \35044 ,
         \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 , \35053 , \35054 ,
         \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 , \35063 , \35064 ,
         \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 ,
         \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 , \35083 , \35084 ,
         \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094 ,
         \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 ,
         \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 , \35113 , \35114 ,
         \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 ,
         \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 , \35133 , \35134 ,
         \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 ,
         \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 ,
         \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 , \35163 , \35164 ,
         \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 ,
         \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 , \35183 , \35184 ,
         \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 ,
         \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 , \35203 , \35204 ,
         \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 ,
         \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 ,
         \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 , \35233 , \35234 ,
         \35235 , \35236 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 , \35243 , \35244 ,
         \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 ,
         \35255 , \35256 , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 , \35263 , \35264 ,
         \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 , \35273 , \35274 ,
         \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 , \35283 , \35284 ,
         \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 , \35293 , \35294 ,
         \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 , \35303 , \35304 ,
         \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 ,
         \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 ,
         \35325 , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 , \35333 , \35334 ,
         \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 , \35343 , \35344 ,
         \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 , \35353 , \35354 ,
         \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 , \35363 , \35364 ,
         \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 , \35373 , \35374 ,
         \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 ,
         \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 , \35393 , \35394 ,
         \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 , \35403 , \35404 ,
         \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411 , \35412 , \35413 , \35414 ,
         \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 , \35423 , \35424 ,
         \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 , \35433 , \35434 ,
         \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 , \35443 , \35444 ,
         \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 , \35453 , \35454 ,
         \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 , \35463 , \35464 ,
         \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 , \35473 , \35474 ,
         \35475 , \35476 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 , \35483 , \35484 ,
         \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , \35494 ,
         \35495 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 ,
         \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513 , \35514 ,
         \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 , \35523 , \35524 ,
         \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 , \35533 , \35534 ,
         \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 , \35543 , \35544 ,
         \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 ,
         \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 , \35563 , \35564 ,
         \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 , \35573 , \35574 ,
         \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582 , \35583 , \35584 ,
         \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 ,
         \35595 , \35596 , \35597 , \35598 , \35599 , \35600 , \35601 , \35602 , \35603 , \35604 ,
         \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 ,
         \35615 , \35616 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 , \35623 , \35624 ,
         \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633 , \35634 ,
         \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 , \35643 , \35644 ,
         \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 , \35653 , \35654 ,
         \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , \35663 , \35664 ,
         \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 ,
         \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , \35683 , \35684 ,
         \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 ,
         \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 , \35703 , \35704 ,
         \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 , \35713 , \35714 ,
         \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 ,
         \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 , \35733 , \35734 ,
         \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 ,
         \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752 , \35753 , \35754 ,
         \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 ,
         \35765 , \35766 , \35767 , \35768 , \35769 , \35770 , \35771 , \35772 , \35773 , \35774 ,
         \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 ,
         \35785 , \35786 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 , \35793 , \35794 ,
         \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 , \35803 , \35804 ,
         \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 , \35813 , \35814 ,
         \35815 , \35816 , \35817 , \35818 , \35819 , \35820 , \35821 , \35822 , \35823 , \35824 ,
         \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 , \35833 , \35834 ,
         \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 ,
         \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854 ,
         \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 , \35863 , \35864 ,
         \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 , \35873 , \35874 ,
         \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 ,
         \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 , \35893 , \35894 ,
         \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 ,
         \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 ,
         \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 , \35923 , \35924 ,
         \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 ,
         \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 , \35943 , \35944 ,
         \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 ,
         \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 ,
         \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 , \35973 , \35974 ,
         \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 ,
         \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 , \35993 , \35994 ,
         \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 ,
         \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 ,
         \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 , \36024 ,
         \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 ,
         \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 , \36043 , \36044 ,
         \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 , \36053 , \36054 ,
         \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 ,
         \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 ,
         \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 , \36083 , \36084 ,
         \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 , \36093 , \36094 ,
         \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 ,
         \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 , \36113 , \36114 ,
         \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 ,
         \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 , \36133 , \36134 ,
         \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143 , \36144 ,
         \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 ,
         \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 , \36163 , \36164 ,
         \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 , \36173 , \36174 ,
         \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 ,
         \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 ,
         \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 ,
         \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 , \36213 , \36214 ,
         \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 ,
         \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 , \36233 , \36234 ,
         \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 , \36243 , \36244 ,
         \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 ,
         \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 ,
         \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 , \36273 , \36274 ,
         \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 ,
         \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 , \36293 , \36294 ,
         \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 , \36303 , \36304 ,
         \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 ,
         \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 , \36323 , \36324 ,
         \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36334 ,
         \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 , \36343 , \36344 ,
         \36345 , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 , \36353 , \36354 ,
         \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364 ,
         \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 , \36373 , \36374 ,
         \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 , \36383 , \36384 ,
         \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393 , \36394 ,
         \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 , \36403 , \36404 ,
         \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 ,
         \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 , \36423 , \36424 ,
         \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 ,
         \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 ,
         \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 , \36453 , \36454 ,
         \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464 ,
         \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 ,
         \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 , \36483 , \36484 ,
         \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 , \36493 , \36494 ,
         \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 ,
         \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 , \36513 , \36514 ,
         \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 , \36523 , \36524 ,
         \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534 ,
         \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 ,
         \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 , \36553 , \36554 ,
         \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 , \36563 , \36564 ,
         \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 ,
         \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 ,
         \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 , \36593 , \36594 ,
         \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 ,
         \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 ,
         \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 , \36623 , \36624 ,
         \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633 , \36634 ,
         \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 , \36643 , \36644 ,
         \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 ,
         \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 , \36663 , \36664 ,
         \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 , \36673 , \36674 ,
         \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 ,
         \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 , \36693 , \36694 ,
         \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704 ,
         \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 ,
         \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 , \36723 , \36724 ,
         \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 , \36733 , \36734 ,
         \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 ,
         \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 , \36753 , \36754 ,
         \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 , \36763 , \36764 ,
         \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774 ,
         \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 , \36783 , \36784 ,
         \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 ,
         \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 , \36803 , \36804 ,
         \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 , \36814 ,
         \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 ,
         \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 , \36833 , \36834 ,
         \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844 ,
         \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 , \36853 , \36854 ,
         \36855 , \36856 , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 , \36863 , \36864 ,
         \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 , \36873 , \36874 ,
         \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 , \36883 , \36884 ,
         \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 ,
         \36895 , \36896 , \36897 , \36898 , \36899 , \36900 , \36901 , \36902 , \36903 , \36904 ,
         \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914 ,
         \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 , \36923 , \36924 ,
         \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 ,
         \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 , \36943 , \36944 ,
         \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 ,
         \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 , \36964 ,
         \36965 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 , \36973 , \36974 ,
         \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984 ,
         \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 , \36993 , \36994 ,
         \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 ,
         \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012 , \37013 , \37014 ,
         \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 ,
         \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 ,
         \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 , \37043 , \37044 ,
         \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054 ,
         \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 ,
         \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 , \37073 , \37074 ,
         \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 , \37083 , \37084 ,
         \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 ,
         \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 ,
         \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 , \37113 , \37114 ,
         \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 , \37123 , \37124 ,
         \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 ,
         \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 ,
         \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 , \37153 , \37154 ,
         \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 ,
         \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 ,
         \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 ,
         \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 ,
         \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203 , \37204 ,
         \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 ,
         \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 , \37223 , \37224 ,
         \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 , \37233 , \37234 ,
         \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 ,
         \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 , \37253 , \37254 ,
         \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 , \37263 , \37264 ,
         \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 , \37273 , \37274 ,
         \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 ,
         \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 ,
         \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304 ,
         \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 , \37313 , \37314 ,
         \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 , \37323 , \37324 ,
         \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334 ,
         \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 , \37343 , \37344 ,
         \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 , \37353 , \37354 ,
         \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364 ,
         \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 ,
         \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 , \37383 , \37384 ,
         \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 , \37393 , \37394 ,
         \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 ,
         \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 , \37413 , \37414 ,
         \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 , \37423 , \37424 ,
         \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 ,
         \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 , \37443 , \37444 ,
         \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 , \37453 , \37454 ,
         \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 ,
         \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 , \37473 , \37474 ,
         \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 , \37483 , \37484 ,
         \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 ,
         \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 , \37503 , \37504 ,
         \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37514 ,
         \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 , \37523 , \37524 ,
         \37525 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 , \37533 , \37534 ,
         \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544 ,
         \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 , \37553 , \37554 ,
         \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 , \37563 , \37564 ,
         \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 , \37573 , \37574 ,
         \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 ,
         \37585 , \37586 , \37587 , \37588 , \37589 , \37590 , \37591 , \37592 , \37593 , \37594 ,
         \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604 ,
         \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 , \37613 , \37614 ,
         \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 , \37623 , \37624 ,
         \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 , \37633 , \37634 ,
         \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 ,
         \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 , \37653 , \37654 ,
         \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 , \37663 , \37664 ,
         \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 ,
         \37675 , \37676 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 , \37683 , \37684 ,
         \37685 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 , \37693 , \37694 ,
         \37695 , \37696 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 , \37703 , \37704 ,
         \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 , \37713 , \37714 ,
         \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 , \37723 , \37724 ,
         \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 , \37733 , \37734 ,
         \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 , \37743 , \37744 ,
         \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 , \37753 , \37754 ,
         \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 , \37763 , \37764 ,
         \37765 , \37766 , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 ,
         \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 ,
         \37785 , \37786 , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 , \37793 , \37794 ,
         \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 ,
         \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 , \37813 , \37814 ,
         \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 ,
         \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 , \37833 , \37834 ,
         \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 ,
         \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 , \37853 , \37854 ,
         \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 ,
         \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 , \37873 , \37874 ,
         \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 ,
         \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 , \37894 ,
         \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 , \37903 , \37904 ,
         \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 ,
         \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 , \37923 , \37924 ,
         \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 ,
         \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 , \37943 , \37944 ,
         \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 ,
         \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 , \37963 , \37964 ,
         \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974 ,
         \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 , \37983 , \37984 ,
         \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 ,
         \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 , \38003 , \38004 ,
         \38005 , \38006 , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 , \38013 , \38014 ,
         \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 ,
         \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 , \38033 , \38034 ,
         \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 ,
         \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 , \38053 , \38054 ,
         \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 ,
         \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072 , \38073 , \38074 ,
         \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 ,
         \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 , \38093 , \38094 ,
         \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 ,
         \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 ,
         \38115 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 , \38123 , \38124 ,
         \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 , \38133 , \38134 ,
         \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 ,
         \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 ,
         \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 , \38164 ,
         \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 , \38173 , \38174 ,
         \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 , \38183 , \38184 ,
         \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 ,
         \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 , \38203 , \38204 ,
         \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 ,
         \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 , \38223 , \38224 ,
         \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 ,
         \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 , \38243 , \38244 ,
         \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 , \38253 , \38254 ,
         \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 , \38263 , \38264 ,
         \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 ,
         \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 , \38283 , \38284 ,
         \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 ,
         \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 , \38303 , \38304 ,
         \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 ,
         \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 , \38323 , \38324 ,
         \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 , \38333 , \38334 ,
         \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 , \38343 , \38344 ,
         \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 ,
         \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 , \38363 , \38364 ,
         \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 ,
         \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 , \38383 , \38384 ,
         \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 ,
         \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 ,
         \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 , \38413 , \38414 ,
         \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 ,
         \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 ,
         \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 , \38443 , \38444 ,
         \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453 , \38454 ,
         \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 ,
         \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 , \38473 , \38474 ,
         \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 ,
         \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 , \38493 , \38494 ,
         \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 ,
         \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 , \38513 , \38514 ,
         \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 , \38523 , \38524 ,
         \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 ,
         \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 ,
         \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 ,
         \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 ,
         \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 , \38573 , \38574 ,
         \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583 , \38584 ,
         \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 ,
         \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 , \38603 , \38604 ,
         \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 , \38613 , \38614 ,
         \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 , \38623 , \38624 ,
         \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 ,
         \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 , \38643 , \38644 ,
         \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 , \38653 , \38654 ,
         \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663 , \38664 ,
         \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 ,
         \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 , \38683 , \38684 ,
         \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 ,
         \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703 , \38704 ,
         \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 ,
         \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723 , \38724 ,
         \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 , \38733 , \38734 ,
         \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744 ,
         \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 ,
         \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 , \38763 , \38764 ,
         \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 ,
         \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783 , \38784 ,
         \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 ,
         \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 , \38803 , \38804 ,
         \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 , \38814 ,
         \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 , \38823 , \38824 ,
         \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 ,
         \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 , \38843 , \38844 ,
         \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 ,
         \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 ,
         \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 , \38873 , \38874 ,
         \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 ,
         \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893 , \38894 ,
         \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 ,
         \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 , \38913 , \38914 ,
         \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 , \38923 , \38924 ,
         \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 , \38933 , \38934 ,
         \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 ,
         \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 , \38953 , \38954 ,
         \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 ,
         \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 ,
         \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 ,
         \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 ,
         \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 , \39003 , \39004 ,
         \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 ,
         \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024 ,
         \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 , \39033 , \39034 ,
         \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043 , \39044 ,
         \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 ,
         \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064 ,
         \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 ,
         \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 , \39084 ,
         \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 ,
         \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103 , \39104 ,
         \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 ,
         \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 , \39123 , \39124 ,
         \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 ,
         \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 , \39143 , \39144 ,
         \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 , \39153 , \39154 ,
         \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162 , \39163 , \39164 ,
         \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 ,
         \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 , \39183 , \39184 ,
         \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 ,
         \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 , \39203 , \39204 ,
         \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 , \39213 , \39214 ,
         \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 , \39223 , \39224 ,
         \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 , \39233 , \39234 ,
         \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 , \39243 , \39244 ,
         \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 , \39253 , \39254 ,
         \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 , \39263 , \39264 ,
         \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 , \39273 , \39274 ,
         \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 , \39283 , \39284 ,
         \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 , \39293 , \39294 ,
         \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 ,
         \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 , \39314 ,
         \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 , \39323 , \39324 ,
         \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 , \39333 , \39334 ,
         \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 ,
         \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 , \39353 , \39354 ,
         \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 ,
         \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 , \39373 , \39374 ,
         \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 ,
         \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 , \39393 , \39394 ,
         \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 , \39403 , \39404 ,
         \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 , \39413 , \39414 ,
         \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 ,
         \39425 , \39426 , \39427 , \39428 , \39429 , \39430 , \39431 , \39432 , \39433 , \39434 ,
         \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 ,
         \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 ,
         \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 ,
         \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 ,
         \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 , \39483 , \39484 ,
         \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 ,
         \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 , \39503 , \39504 ,
         \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 , \39513 , \39514 ,
         \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 , \39523 , \39524 ,
         \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 ,
         \39535 , \39536 , \39537 , \39538 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 ,
         \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 ,
         \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 , \39564 ,
         \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574 ,
         \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 ,
         \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592 , \39593 , \39594 ,
         \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 ,
         \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 , \39613 , \39614 ,
         \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 , \39623 , \39624 ,
         \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 ,
         \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 ,
         \39645 , \39646 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 ,
         \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664 ,
         \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 , \39673 , \39674 ,
         \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 , \39683 , \39684 ,
         \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 ,
         \39695 , \39696 , \39697 , \39698 , \39699 , \39700 , \39701 , \39702 , \39703 , \39704 ,
         \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 ,
         \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 ,
         \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 ,
         \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 ,
         \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 , \39753 , \39754 ,
         \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 ,
         \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 , \39773 , \39774 ,
         \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 ,
         \39785 , \39786 , \39787 , \39788 , \39789 , \39790 , \39791 , \39792 , \39793 , \39794 ,
         \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 ,
         \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 ,
         \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 , \39823 , \39824 ,
         \39825 , \39826 , \39827 , \39828 , \39829 , \39830 , \39831 , \39832 , \39833 , \39834 ,
         \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844 ,
         \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852 , \39853 , \39854 ,
         \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 , \39863 , \39864 ,
         \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 , \39873 , \39874 ,
         \39875 , \39876 , \39877 , \39878 , \39879 , \39880 , \39881 , \39882 , \39883 , \39884 ,
         \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 ,
         \39895 , \39896 , \39897 , \39898 , \39899 , \39900 , \39901 , \39902 , \39903 , \39904 ,
         \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 ,
         \39915 , \39916 , \39917 , \39918 , \39919 , \39920 , \39921 , \39922 , \39923 , \39924 ,
         \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934 ,
         \39935 , \39936 , \39937 , \39938 , \39939 , \39940 , \39941 , \39942 , \39943 , \39944 ,
         \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 , \39953 , \39954 ,
         \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962 , \39963 , \39964 ,
         \39965 , \39966 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 , \39973 , \39974 ,
         \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 , \39983 , \39984 ,
         \39985 , \39986 , \39987 , \39988 , \39989 , \39990 , \39991 , \39992 , \39993 , \39994 ,
         \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002 , \40003 , \40004 ,
         \40005 , \40006 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 , \40013 , \40014 ,
         \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 , \40023 , \40024 ,
         \40025 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 , \40033 , \40034 ,
         \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 , \40043 , \40044 ,
         \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 , \40053 , \40054 ,
         \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 , \40063 , \40064 ,
         \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 , \40073 , \40074 ,
         \40075 , \40076 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 , \40083 , \40084 ,
         \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 , \40093 , \40094 ,
         \40095 , \40096 , \40097 , \40098 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 ,
         \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 ,
         \40115 , \40116 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 , \40123 , \40124 ,
         \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133 , \40134 ,
         \40135 , \40136 , \40137 , \40138 , \40139 , \40140 , \40141 , \40142 , \40143 , \40144 ,
         \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 , \40153 , \40154 ,
         \40155 , \40156 , \40157 , \40158 , \40159 , \40160 , \40161 , \40162 , \40163 , \40164 ,
         \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 , \40173 , \40174 ,
         \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182 , \40183 , \40184 ,
         \40185 , \40186 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 ,
         \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 , \40203 , \40204 ,
         \40205 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 ,
         \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223 , \40224 ,
         \40225 , \40226 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 , \40233 , \40234 ,
         \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 , \40243 , \40244 ,
         \40245 , \40246 , \40247 , \40248 , \40249 , \40250 , \40251 , \40252 , \40253 , \40254 ,
         \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 , \40263 , \40264 ,
         \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271 , \40272 , \40273 , \40274 ,
         \40275 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 ,
         \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 , \40293 , \40294 ,
         \40295 , \40296 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 ,
         \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 , \40314 ,
         \40315 , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 , \40323 , \40324 ,
         \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 , \40333 , \40334 ,
         \40335 , \40336 , \40337 , \40338 , \40339 , \40340 , \40341 , \40342 , \40343 , \40344 ,
         \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 , \40353 , \40354 ,
         \40355 , \40356 , \40357 , \40358 , \40359 , \40360 , \40361 , \40362 , \40363 , \40364 ,
         \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 ,
         \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381 , \40382 , \40383 , \40384 ,
         \40385 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 ,
         \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 , \40403 , \40404 ,
         \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411 , \40412 , \40413 , \40414 ,
         \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422 , \40423 , \40424 ,
         \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 ,
         \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 , \40443 , \40444 ,
         \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 , \40453 , \40454 ,
         \40455 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 ,
         \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 ,
         \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 , \40483 , \40484 ,
         \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 ,
         \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 ,
         \40505 , \40506 , \40507 , \40508 , \40509 , \40510 , \40511 , \40512 , \40513 , \40514 ,
         \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 ,
         \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 ,
         \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 , \40543 , \40544 ,
         \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 ,
         \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563 , \40564 ,
         \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 ,
         \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 , \40583 , \40584 ,
         \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 , \40594 ,
         \40595 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 , \40603 , \40604 ,
         \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 ,
         \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 , \40623 , \40624 ,
         \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633 , \40634 ,
         \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 ,
         \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651 , \40652 , \40653 , \40654 ,
         \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 ,
         \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 , \40673 , \40674 ,
         \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 , \40683 , \40684 ,
         \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 ,
         \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 ,
         \40705 , \40706 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 ,
         \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724 ,
         \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 , \40734 ,
         \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 , \40743 , \40744 ,
         \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 ,
         \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 , \40762 , \40763 , \40764 ,
         \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 ,
         \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 ,
         \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792 , \40793 , \40794 ,
         \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 ,
         \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 , \40813 , \40814 ,
         \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 , \40823 , \40824 ,
         \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 ,
         \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843 , \40844 ,
         \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 , \40853 , \40854 ,
         \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 , \40863 , \40864 ,
         \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 ,
         \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 , \40882 , \40883 , \40884 ,
         \40885 , \40886 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 ,
         \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 ,
         \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 , \40913 , \40914 ,
         \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 ,
         \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 , \40933 , \40934 ,
         \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 , \40943 , \40944 ,
         \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 ,
         \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963 , \40964 ,
         \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 , \40973 , \40974 ,
         \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 , \40983 , \40984 ,
         \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 ,
         \40995 , \40996 , \40997 , \40998 , \40999 , \41000 , \41001 , \41002 , \41003 , \41004 ,
         \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014 ,
         \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 ,
         \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031 , \41032 , \41033 , \41034 ,
         \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 , \41043 , \41044 ,
         \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 ,
         \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 ,
         \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 ,
         \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 , \41083 , \41084 ,
         \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 ,
         \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 , \41103 , \41104 ,
         \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 , \41113 , \41114 ,
         \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 ,
         \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133 , \41134 ,
         \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 , \41143 , \41144 ,
         \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 , \41153 , \41154 ,
         \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 ,
         \41165 , \41166 , \41167 , \41168 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 ,
         \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184 ,
         \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 ,
         \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 , \41203 , \41204 ,
         \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 ,
         \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 , \41223 , \41224 ,
         \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 ,
         \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 ,
         \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252 , \41253 , \41254 ,
         \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 ,
         \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 , \41273 , \41274 ,
         \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 , \41283 , \41284 ,
         \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 ,
         \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304 ,
         \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 , \41313 , \41314 ,
         \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 , \41323 , \41324 ,
         \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 ,
         \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 , \41343 , \41344 ,
         \41345 , \41346 , \41347 , \41348 , \41349 , \41350 , \41351 , \41352 , \41353 , \41354 ,
         \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 ,
         \41365 , \41366 , \41367 , \41368 , \41369 , \41370 , \41371 , \41372 , \41373 , \41374 ,
         \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 , \41383 , \41384 ,
         \41385 , \41386 , \41387 , \41388 , \41389 , \41390 , \41391 , \41392 , \41393 , \41394 ,
         \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 ,
         \41405 , \41406 , \41407 , \41408 , \41409 , \41410 , \41411 , \41412 , \41413 , \41414 ,
         \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424 ,
         \41425 , \41426 , \41427 , \41428 , \41429 , \41430 , \41431 , \41432 , \41433 , \41434 ,
         \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 , \41443 , \41444 ,
         \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451 , \41452 , \41453 , \41454 ,
         \41455 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 ,
         \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472 , \41473 , \41474 ,
         \41475 , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 ,
         \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492 , \41493 , \41494 ,
         \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 , \41503 , \41504 ,
         \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 , \41513 , \41514 ,
         \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 ,
         \41525 , \41526 , \41527 , \41528 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 ,
         \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544 ,
         \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 ,
         \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 , \41563 , \41564 ,
         \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 ,
         \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 , \41583 , \41584 ,
         \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 ,
         \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 ,
         \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 , \41613 , \41614 ,
         \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 , \41623 , \41624 ,
         \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 ,
         \41635 , \41636 , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 , \41643 , \41644 ,
         \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653 , \41654 ,
         \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 ,
         \41665 , \41666 , \41667 , \41668 , \41669 , \41670 , \41671 , \41672 , \41673 , \41674 ,
         \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683 , \41684 ,
         \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 ,
         \41695 , \41696 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 ,
         \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 , \41713 , \41714 ,
         \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 , \41723 , \41724 ,
         \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 ,
         \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 , \41743 , \41744 ,
         \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 , \41753 , \41754 ,
         \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 ,
         \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 , \41773 , \41774 ,
         \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 , \41783 , \41784 ,
         \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 ,
         \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 ,
         \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811 , \41812 , \41813 , \41814 ,
         \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 ,
         \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 ,
         \41835 , \41836 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 , \41843 , \41844 ,
         \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854 ,
         \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 , \41863 , \41864 ,
         \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 ,
         \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 , \41883 , \41884 ,
         \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 , \41893 , \41894 ,
         \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 ,
         \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 , \41913 , \41914 ,
         \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 , \41923 , \41924 ,
         \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 ,
         \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 ,
         \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 , \41953 , \41954 ,
         \41955 , \41956 , \41957 , \41958 , \41959 , \41960 , \41961 , \41962 , \41963 , \41964 ,
         \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 ,
         \41975 , \41976 , \41977 , \41978 , \41979 , \41980 , \41981 , \41982 , \41983 , \41984 ,
         \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994 ,
         \41995 , \41996 , \41997 , \41998 , \41999 , \42000 , \42001 , \42002 , \42003 , \42004 ,
         \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 ,
         \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021 , \42022 , \42023 , \42024 ,
         \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 ,
         \42035 , \42036 , \42037 , \42038 , \42039 , \42040 , \42041 , \42042 , \42043 , \42044 ,
         \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 , \42053 , \42054 ,
         \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 , \42063 , \42064 ,
         \42065 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 ,
         \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 , \42083 , \42084 ,
         \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 , \42093 , \42094 ,
         \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 , \42104 ,
         \42105 , \42106 , \42107 , \42108 , \42109 , \42110 , \42111 , \42112 , \42113 , \42114 ,
         \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121 , \42122 , \42123 , \42124 ,
         \42125 , \42126 , \42127 , \42128 , \42129 , \42130 , \42131 , \42132 , \42133 , \42134 ,
         \42135 , \42136 , \42137 , \42138 , \42139 , \42140 , \42141 , \42142 , \42143 , \42144 ,
         \42145 , \42146 , \42147 , \42148 , \42149 , \42150 , \42151 , \42152 , \42153 , \42154 ,
         \42155 , \42156 , \42157 , \42158 , \42159 , \42160 , \42161 , \42162 , \42163 , \42164 ,
         \42165 , \42166 , \42167 , \42168 , \42169 , \42170 , \42171 , \42172 , \42173 , \42174 ,
         \42175 , \42176 , \42177 , \42178 , \42179 , \42180 , \42181 , \42182 , \42183 , \42184 ,
         \42185 , \42186 , \42187 , \42188 , \42189 , \42190 , \42191 , \42192 , \42193 , \42194 ,
         \42195 , \42196 , \42197 , \42198 , \42199 , \42200 , \42201 , \42202 , \42203 , \42204 ,
         \42205 , \42206 , \42207 , \42208 , \42209 , \42210 , \42211 , \42212 , \42213 , \42214 ,
         \42215 , \42216 , \42217 , \42218 , \42219 , \42220 , \42221 , \42222 , \42223 , \42224 ,
         \42225 , \42226 , \42227 , \42228 , \42229 , \42230 , \42231 , \42232 , \42233 , \42234 ,
         \42235 , \42236 , \42237 , \42238 , \42239 , \42240 , \42241 , \42242 , \42243 , \42244 ,
         \42245 , \42246 , \42247 , \42248 , \42249 , \42250 , \42251 , \42252 , \42253 , \42254 ,
         \42255 , \42256 , \42257 , \42258 , \42259 , \42260 , \42261 , \42262 , \42263 , \42264 ,
         \42265 , \42266 , \42267 , \42268 , \42269 , \42270 , \42271 , \42272 , \42273 , \42274 ,
         \42275 , \42276 , \42277 , \42278 , \42279 , \42280 , \42281 , \42282 , \42283 , \42284 ,
         \42285 , \42286 , \42287 , \42288 , \42289 , \42290 , \42291 , \42292 , \42293 , \42294 ,
         \42295 , \42296 , \42297 , \42298 , \42299 , \42300 , \42301 , \42302 , \42303 , \42304 ,
         \42305 , \42306 , \42307 , \42308 , \42309 , \42310 , \42311 , \42312 , \42313 , \42314 ,
         \42315 , \42316 , \42317 , \42318 , \42319 , \42320 , \42321 , \42322 , \42323 , \42324 ,
         \42325 , \42326 , \42327 , \42328 , \42329 , \42330 , \42331 , \42332 , \42333 , \42334 ,
         \42335 , \42336 , \42337 , \42338 , \42339 , \42340 , \42341 , \42342 , \42343 , \42344 ,
         \42345 , \42346 , \42347 , \42348 , \42349 , \42350 , \42351 , \42352 , \42353 , \42354 ,
         \42355 , \42356 , \42357 , \42358 , \42359 , \42360 , \42361 , \42362 , \42363 , \42364 ,
         \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 , \42373 , \42374 ,
         \42375 , \42376 , \42377 , \42378 , \42379 , \42380 , \42381 , \42382 , \42383 , \42384 ,
         \42385 , \42386 , \42387 , \42388 , \42389 , \42390 , \42391 , \42392 , \42393 , \42394 ,
         \42395 , \42396 , \42397 , \42398 , \42399 , \42400 , \42401 , \42402 , \42403 , \42404 ,
         \42405 , \42406 , \42407 , \42408 , \42409 , \42410 , \42411 , \42412 , \42413 , \42414 ,
         \42415 , \42416 , \42417 , \42418 , \42419 , \42420 , \42421 , \42422 , \42423 , \42424 ,
         \42425 , \42426 , \42427 , \42428 , \42429 , \42430 , \42431 , \42432 , \42433 , \42434 ,
         \42435 , \42436 , \42437 , \42438 , \42439 , \42440 , \42441 , \42442 , \42443 , \42444 ,
         \42445 , \42446 , \42447 , \42448 , \42449 , \42450 , \42451 , \42452 , \42453 , \42454 ,
         \42455 , \42456 , \42457 , \42458 , \42459 , \42460 , \42461 , \42462 , \42463 , \42464 ,
         \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471 , \42472 , \42473 , \42474 ,
         \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 , \42483 , \42484 ,
         \42485 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 , \42493 , \42494 ,
         \42495 , \42496 , \42497 , \42498 , \42499 , \42500 , \42501 , \42502 , \42503 , \42504 ,
         \42505 , \42506 , \42507 , \42508 , \42509 , \42510 , \42511 , \42512 , \42513 , \42514 ,
         \42515 , \42516 , \42517 , \42518 , \42519 , \42520 , \42521 , \42522 , \42523 , \42524 ,
         \42525 , \42526 , \42527 , \42528 , \42529 , \42530 , \42531 , \42532 , \42533 , \42534 ,
         \42535 , \42536 , \42537 , \42538 , \42539 , \42540 , \42541 , \42542 , \42543 , \42544 ,
         \42545 , \42546 , \42547 , \42548 , \42549 , \42550 , \42551 , \42552 , \42553 , \42554 ,
         \42555 , \42556 , \42557 , \42558 , \42559 , \42560 , \42561 , \42562 , \42563 , \42564 ,
         \42565 , \42566 , \42567 , \42568 , \42569 , \42570 , \42571 , \42572 , \42573 , \42574 ,
         \42575 , \42576 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582 , \42583 , \42584 ,
         \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591 , \42592 , \42593 , \42594 ,
         \42595 , \42596 , \42597 , \42598 , \42599 , \42600 , \42601 , \42602 , \42603 , \42604 ,
         \42605 , \42606 , \42607 , \42608 , \42609 , \42610 , \42611 , \42612 , \42613 , \42614 ,
         \42615 , \42616 , \42617 , \42618 , \42619 , \42620 , \42621 , \42622 , \42623 , \42624 ,
         \42625 , \42626 , \42627 , \42628 , \42629 , \42630 , \42631 , \42632 , \42633 , \42634 ,
         \42635 , \42636 , \42637 , \42638 , \42639 , \42640 , \42641 , \42642 , \42643 , \42644 ,
         \42645 , \42646 , \42647 , \42648 , \42649 , \42650 , \42651 , \42652 , \42653 , \42654 ,
         \42655 , \42656 , \42657 , \42658 , \42659 , \42660 , \42661 , \42662 , \42663 , \42664 ,
         \42665 , \42666 , \42667 , \42668 , \42669 , \42670 , \42671 , \42672 , \42673 , \42674 ,
         \42675 , \42676 , \42677 , \42678 , \42679 , \42680 , \42681 , \42682 , \42683 , \42684 ,
         \42685 , \42686 , \42687 , \42688 , \42689 , \42690 , \42691 , \42692 , \42693 , \42694 ,
         \42695 , \42696 , \42697 , \42698 , \42699 , \42700 , \42701 , \42702 , \42703 , \42704 ,
         \42705 , \42706 , \42707 , \42708 , \42709 , \42710 , \42711 , \42712 , \42713 , \42714 ,
         \42715 , \42716 , \42717 , \42718 , \42719 , \42720 , \42721 , \42722 , \42723 , \42724 ,
         \42725 , \42726 , \42727 , \42728 , \42729 , \42730 , \42731 , \42732 , \42733 , \42734 ,
         \42735 , \42736 , \42737 , \42738 , \42739 , \42740 , \42741 , \42742 , \42743 , \42744 ,
         \42745 , \42746 , \42747 , \42748 , \42749 , \42750 , \42751 , \42752 , \42753 , \42754 ,
         \42755 , \42756 , \42757 , \42758 , \42759 , \42760 , \42761 , \42762 , \42763 , \42764 ,
         \42765 , \42766 , \42767 , \42768 , \42769 , \42770 , \42771 , \42772 , \42773 , \42774 ,
         \42775 , \42776 , \42777 , \42778 , \42779 , \42780 , \42781 , \42782 , \42783 , \42784 ,
         \42785 , \42786 , \42787 , \42788 , \42789 , \42790 , \42791 , \42792 , \42793 , \42794 ,
         \42795 , \42796 , \42797 , \42798 , \42799 , \42800 , \42801 , \42802 , \42803 , \42804 ,
         \42805 , \42806 , \42807 , \42808 , \42809 , \42810 , \42811 , \42812 , \42813 , \42814 ,
         \42815 , \42816 , \42817 , \42818 , \42819 , \42820 , \42821 , \42822 , \42823 , \42824 ,
         \42825 , \42826 , \42827 , \42828 , \42829 , \42830 , \42831 , \42832 , \42833 , \42834 ,
         \42835 , \42836 , \42837 , \42838 , \42839 , \42840 , \42841 , \42842 , \42843 , \42844 ,
         \42845 , \42846 , \42847 , \42848 , \42849 , \42850 , \42851 , \42852 , \42853 , \42854 ,
         \42855 , \42856 , \42857 , \42858 , \42859 , \42860 , \42861 , \42862 , \42863 , \42864 ,
         \42865 , \42866 , \42867 , \42868 , \42869 , \42870 , \42871 , \42872 , \42873 , \42874 ,
         \42875 , \42876 , \42877 , \42878 , \42879 , \42880 , \42881 , \42882 , \42883 , \42884 ,
         \42885 , \42886 , \42887 , \42888 , \42889 , \42890 , \42891 , \42892 , \42893 , \42894 ,
         \42895 , \42896 , \42897 , \42898 , \42899 , \42900 , \42901 , \42902 , \42903 , \42904 ,
         \42905 , \42906 , \42907 , \42908 , \42909 , \42910 , \42911 , \42912 , \42913 , \42914 ,
         \42915 , \42916 , \42917 , \42918 , \42919 , \42920 , \42921 , \42922 , \42923 , \42924 ,
         \42925 , \42926 , \42927 , \42928 , \42929 , \42930 , \42931 , \42932 , \42933 , \42934 ,
         \42935 , \42936 , \42937 , \42938 , \42939 , \42940 , \42941 , \42942 , \42943 , \42944 ,
         \42945 , \42946 , \42947 , \42948 , \42949 , \42950 , \42951 , \42952 , \42953 , \42954 ,
         \42955 , \42956 , \42957 , \42958 , \42959 , \42960 , \42961 , \42962 , \42963 , \42964 ,
         \42965 , \42966 , \42967 , \42968 , \42969 , \42970 , \42971 , \42972 , \42973 , \42974 ,
         \42975 , \42976 , \42977 , \42978 , \42979 , \42980 , \42981 , \42982 , \42983 , \42984 ,
         \42985 , \42986 , \42987 , \42988 , \42989 , \42990 , \42991 , \42992 , \42993 , \42994 ,
         \42995 , \42996 , \42997 , \42998 , \42999 , \43000 , \43001 , \43002 , \43003 , \43004 ,
         \43005 , \43006 , \43007 , \43008 , \43009 , \43010 , \43011 , \43012 , \43013 , \43014 ,
         \43015 , \43016 , \43017 , \43018 , \43019 , \43020 , \43021 , \43022 , \43023 , \43024 ,
         \43025 , \43026 , \43027 , \43028 , \43029 , \43030 , \43031 , \43032 , \43033 , \43034 ,
         \43035 , \43036 , \43037 , \43038 , \43039 , \43040 , \43041 , \43042 , \43043 , \43044 ,
         \43045 , \43046 , \43047 , \43048 , \43049 , \43050 , \43051 , \43052 , \43053 , \43054 ,
         \43055 , \43056 , \43057 , \43058 , \43059 , \43060 , \43061 , \43062 , \43063 , \43064 ,
         \43065 , \43066 , \43067 , \43068 , \43069 , \43070 , \43071 , \43072 , \43073 , \43074 ,
         \43075 , \43076 , \43077 , \43078 , \43079 , \43080 , \43081 , \43082 , \43083 , \43084 ,
         \43085 , \43086 , \43087 , \43088 , \43089 , \43090 , \43091 , \43092 , \43093 , \43094 ,
         \43095 , \43096 , \43097 , \43098 , \43099 , \43100 , \43101 , \43102 , \43103 , \43104 ,
         \43105 , \43106 , \43107 , \43108 , \43109 , \43110 , \43111 , \43112 , \43113 , \43114 ,
         \43115 , \43116 , \43117 , \43118 , \43119 , \43120 , \43121 , \43122 , \43123 , \43124 ,
         \43125 , \43126 , \43127 , \43128 , \43129 , \43130 , \43131 , \43132 , \43133 , \43134 ,
         \43135 , \43136 , \43137 , \43138 , \43139 , \43140 , \43141 , \43142 , \43143 , \43144 ,
         \43145 , \43146 , \43147 , \43148 , \43149 , \43150 , \43151 , \43152 , \43153 , \43154 ,
         \43155 , \43156 , \43157 , \43158 , \43159 , \43160 , \43161 , \43162 , \43163 , \43164 ,
         \43165 , \43166 , \43167 , \43168 , \43169 , \43170 , \43171 , \43172 , \43173 , \43174 ,
         \43175 , \43176 , \43177 , \43178 , \43179 , \43180 , \43181 , \43182 , \43183 , \43184 ,
         \43185 , \43186 , \43187 , \43188 , \43189 , \43190 , \43191 , \43192 , \43193 , \43194 ,
         \43195 , \43196 , \43197 , \43198 , \43199 , \43200 , \43201 , \43202 , \43203 , \43204 ,
         \43205 , \43206 , \43207 , \43208 , \43209 , \43210 , \43211 , \43212 , \43213 , \43214 ,
         \43215 , \43216 , \43217 , \43218 , \43219 , \43220 , \43221 , \43222 , \43223 , \43224 ,
         \43225 , \43226 , \43227 , \43228 , \43229 , \43230 , \43231 , \43232 , \43233 , \43234 ,
         \43235 , \43236 , \43237 , \43238 , \43239 , \43240 , \43241 , \43242 , \43243 , \43244 ,
         \43245 , \43246 , \43247 , \43248 , \43249 , \43250 , \43251 , \43252 , \43253 , \43254 ,
         \43255 , \43256 , \43257 , \43258 , \43259 , \43260 , \43261 , \43262 , \43263 , \43264 ,
         \43265 , \43266 , \43267 , \43268 , \43269 , \43270 , \43271 , \43272 , \43273 , \43274 ,
         \43275 , \43276 , \43277 , \43278 , \43279 , \43280 , \43281 , \43282 , \43283 , \43284 ,
         \43285 , \43286 , \43287 , \43288 , \43289 , \43290 , \43291 , \43292 , \43293 , \43294 ,
         \43295 , \43296 , \43297 , \43298 , \43299 , \43300 , \43301 , \43302 , \43303 , \43304 ,
         \43305 , \43306 , \43307 , \43308 , \43309 , \43310 , \43311 , \43312 , \43313 , \43314 ,
         \43315 , \43316 , \43317 , \43318 , \43319 , \43320 , \43321 , \43322 , \43323 , \43324 ,
         \43325 , \43326 , \43327 , \43328 , \43329 , \43330 , \43331 , \43332 , \43333 , \43334 ,
         \43335 , \43336 , \43337 , \43338 , \43339 , \43340 , \43341 , \43342 , \43343 , \43344 ,
         \43345 , \43346 , \43347 , \43348 , \43349 , \43350 , \43351 , \43352 , \43353 , \43354 ,
         \43355 , \43356 , \43357 , \43358 , \43359 , \43360 , \43361 , \43362 , \43363 , \43364 ,
         \43365 , \43366 , \43367 , \43368 , \43369 , \43370 , \43371 , \43372 , \43373 , \43374 ,
         \43375 , \43376 , \43377 , \43378 , \43379 , \43380 , \43381 , \43382 , \43383 , \43384 ,
         \43385 , \43386 , \43387 , \43388 , \43389 , \43390 , \43391 , \43392 , \43393 , \43394 ,
         \43395 , \43396 , \43397 , \43398 , \43399 , \43400 , \43401 , \43402 , \43403 , \43404 ,
         \43405 , \43406 , \43407 , \43408 , \43409 , \43410 , \43411 , \43412 , \43413 , \43414 ,
         \43415 , \43416 , \43417 , \43418 , \43419 , \43420 , \43421 , \43422 , \43423 , \43424 ,
         \43425 , \43426 , \43427 , \43428 , \43429 , \43430 , \43431 , \43432 , \43433 , \43434 ,
         \43435 , \43436 , \43437 , \43438 , \43439 , \43440 , \43441 , \43442 , \43443 , \43444 ,
         \43445 , \43446 , \43447 , \43448 , \43449 , \43450 , \43451 , \43452 , \43453 , \43454 ,
         \43455 , \43456 , \43457 , \43458 , \43459 , \43460 , \43461 , \43462 , \43463 , \43464 ,
         \43465 , \43466 , \43467 , \43468 , \43469 , \43470 , \43471 , \43472 , \43473 , \43474 ,
         \43475 , \43476 , \43477 , \43478 , \43479 , \43480 , \43481 , \43482 , \43483 , \43484 ,
         \43485 , \43486 , \43487 , \43488 , \43489 ;
buf \U$labaj4393 ( R_101_9cd3d68, \41984 );
buf \U$labaj4394 ( R_102_9cd3e10, \42007 );
buf \U$labaj4395 ( R_103_9cd3eb8, \42020 );
buf \U$labaj4396 ( R_104_9cd3f60, \42028 );
buf \U$labaj4397 ( R_105_9cd4008, \42040 );
buf \U$labaj4398 ( R_106_9cd40b0, \42049 );
buf \U$labaj4399 ( R_107_9cd4158, \42058 );
buf \U$labaj4400 ( R_108_9cd4200, \42063 );
buf \U$labaj4401 ( R_109_9cd42a8, \42073 );
buf \U$labaj4402 ( R_10a_9cd4350, \42091 );
buf \U$labaj4403 ( R_10b_9cd43f8, \42101 );
buf \U$labaj4404 ( R_10c_9cd44a0, \42109 );
buf \U$labaj4405 ( R_10d_9cd4548, \42123 );
buf \U$labaj4406 ( R_10e_9cd45f0, \42127 );
buf \U$labaj4407 ( R_10f_9cd4698, \42137 );
buf \U$labaj4408 ( R_110_9cd4740, \42141 );
buf \U$labaj4409 ( R_111_9cd47e8, \42159 );
buf \U$labaj4410 ( R_112_9cd4890, \42175 );
buf \U$labaj4411 ( R_113_9cd4938, \42183 );
buf \U$labaj4412 ( R_114_9cd49e0, \42188 );
buf \U$labaj4413 ( R_115_9cd4a88, \42204 );
buf \U$labaj4414 ( R_116_9cd4b30, \42208 );
buf \U$labaj4415 ( R_117_9cd4bd8, \42217 );
buf \U$labaj4416 ( R_118_9cd4c80, \42221 );
buf \U$labaj4417 ( R_119_9cd4d28, \42236 );
buf \U$labaj4418 ( R_11a_9cd4dd0, \42246 );
buf \U$labaj4419 ( R_11b_9cd4e78, \42261 );
buf \U$labaj4420 ( R_11c_9cd4f20, \42265 );
buf \U$labaj4421 ( R_11d_9cd4fc8, \42274 );
buf \U$labaj4422 ( R_11e_9cd5070, \42284 );
buf \U$labaj4423 ( R_11f_9cd5118, \42293 );
buf \U$labaj4424 ( R_120_9cd51c0, \42298 );
buf \U$labaj4425 ( R_121_9cd5268, \42328 );
buf \U$labaj4426 ( R_122_9cd5310, \42345 );
buf \U$labaj4427 ( R_123_9cd53b8, \42353 );
buf \U$labaj4428 ( R_124_9cd5460, \42357 );
buf \U$labaj4429 ( R_125_9cd5508, \42382 );
buf \U$labaj4430 ( R_126_9cd55b0, \42390 );
buf \U$labaj4431 ( R_127_9cd5658, \42400 );
buf \U$labaj4432 ( R_128_9cd5700, \42408 );
buf \U$labaj4433 ( R_129_9cd57a8, \42431 );
buf \U$labaj4434 ( R_12a_9cd5850, \42444 );
buf \U$labaj4435 ( R_12b_9cd58f8, \42454 );
buf \U$labaj4436 ( R_12c_9cd59a0, \42462 );
buf \U$labaj4437 ( R_12d_9cd5a48, \42472 );
buf \U$labaj4438 ( R_12e_9cd5af0, \42478 );
buf \U$labaj4439 ( R_12f_9cd5b98, \42487 );
buf \U$labaj4440 ( R_130_9cd5c40, \42495 );
buf \U$labaj4441 ( R_131_9cd5ce8, \42522 );
buf \U$labaj4442 ( R_132_9cd5d90, \42526 );
buf \U$labaj4443 ( R_133_9cd5e38, \42540 );
buf \U$labaj4444 ( R_134_9cd5ee0, \42544 );
buf \U$labaj4445 ( R_135_9cd5f88, \42556 );
buf \U$labaj4446 ( R_136_9cd6030, \42567 );
buf \U$labaj4447 ( R_137_9cd60d8, \42579 );
buf \U$labaj4448 ( R_138_9cd6180, \42587 );
buf \U$labaj4449 ( R_139_9cd6228, \42603 );
buf \U$labaj4450 ( R_13a_9cd62d0, \42612 );
buf \U$labaj4451 ( R_13b_9cd6378, \42621 );
buf \U$labaj4452 ( R_13c_9cd6420, \42629 );
buf \U$labaj4453 ( R_13d_9cd64c8, \42646 );
buf \U$labaj4454 ( R_13e_9cd6570, \42651 );
buf \U$labaj4455 ( R_13f_9cd6618, \42664 );
buf \U$labaj4456 ( R_140_9cd66c0, \42672 );
buf \U$labaj4457 ( R_141_9cd6768, \42705 );
buf \U$labaj4458 ( R_142_9cd6810, \42717 );
buf \U$labaj4459 ( R_143_9cd68b8, \42734 );
buf \U$labaj4460 ( R_144_9cd6960, \42746 );
buf \U$labaj4461 ( R_145_9cd6a08, \42769 );
buf \U$labaj4462 ( R_146_9cd6ab0, \42782 );
buf \U$labaj4463 ( R_147_9cd6b58, \42801 );
buf \U$labaj4464 ( R_148_9cd6c00, \42809 );
buf \U$labaj4465 ( R_149_9cd6ca8, \42839 );
buf \U$labaj4466 ( R_14a_9cd6d50, \42851 );
buf \U$labaj4467 ( R_14b_9cd6df8, \42868 );
buf \U$labaj4468 ( R_14c_9cd6ea0, \42880 );
buf \U$labaj4469 ( R_14d_9cd6f48, \42902 );
buf \U$labaj4470 ( R_14e_9cd6ff0, \42914 );
buf \U$labaj4471 ( R_14f_9cd7098, \42934 );
buf \U$labaj4472 ( R_150_9cd7140, \42941 );
buf \U$labaj4473 ( R_151_9cd71e8, \42974 );
buf \U$labaj4474 ( R_152_9cd7290, \42985 );
buf \U$labaj4475 ( R_153_9cd7338, \43002 );
buf \U$labaj4476 ( R_154_9cd73e0, \43009 );
buf \U$labaj4477 ( R_155_9cd7488, \43031 );
buf \U$labaj4478 ( R_156_9cd7530, \43042 );
buf \U$labaj4479 ( R_157_9cd75d8, \43058 );
buf \U$labaj4480 ( R_158_9cd7680, \43065 );
buf \U$labaj4481 ( R_159_9cd7728, \43090 );
buf \U$labaj4482 ( R_15a_9cd77d0, \43101 );
buf \U$labaj4483 ( R_15b_9cd7878, \43117 );
buf \U$labaj4484 ( R_15c_9cd7920, \43129 );
buf \U$labaj4485 ( R_15d_9cd79c8, \43150 );
buf \U$labaj4486 ( R_15e_9cd7a70, \43162 );
buf \U$labaj4487 ( R_15f_9cd7b18, \43179 );
buf \U$labaj4488 ( R_160_9cd7bc0, \43186 );
buf \U$labaj4489 ( R_161_9cd7c68, \43217 );
buf \U$labaj4490 ( R_162_9cd7d10, \43229 );
buf \U$labaj4491 ( R_163_9cd7db8, \43241 );
buf \U$labaj4492 ( R_164_9cd7e60, \43252 );
buf \U$labaj4493 ( R_165_9cd7f08, \43273 );
buf \U$labaj4494 ( R_166_9cd7fb0, \43280 );
buf \U$labaj4495 ( R_167_9cd8058, \43296 );
buf \U$labaj4496 ( R_168_9cd8100, \43303 );
buf \U$labaj4497 ( R_169_9cd81a8, \43324 );
buf \U$labaj4498 ( R_16a_9cd8250, \43332 );
buf \U$labaj4499 ( R_16b_9cd82f8, \43347 );
buf \U$labaj4500 ( R_16c_9cd83a0, \43354 );
buf \U$labaj4501 ( R_16d_9cd8448, \43375 );
buf \U$labaj4502 ( R_16e_9cd84f0, \43388 );
buf \U$labaj4503 ( R_16f_9cd8598, \43404 );
buf \U$labaj4504 ( R_170_9cd8640, \43411 );
buf \U$labaj4505 ( R_171_9cd86e8, \43431 );
buf \U$labaj4506 ( R_172_9cd8790, \43438 );
buf \U$labaj4507 ( R_173_9cd8838, \43451 );
buf \U$labaj4508 ( R_174_9cd88e0, \43463 );
buf \U$labaj4509 ( R_175_9cd8988, \43471 );
buf \U$labaj4510 ( R_176_9cd8a30, \43479 );
buf \U$labaj4511 ( R_177_9cd8ad8, \43489 );
not \U$1 ( \378 , RIc224f40_83);
not \U$2 ( \379 , RIc229e00_147);
and \U$3 ( \380 , \378 , \379 );
nor \U$4 ( \381 , RIc224ec8_84, RIc229e78_148);
nor \U$5 ( \382 , \380 , \381 );
nor \U$6 ( \383 , RIc224fb8_82, RIc229d88_146);
nor \U$7 ( \384 , RIc225030_81, RIc229d10_145);
nor \U$8 ( \385 , \383 , \384 );
nand \U$9 ( \386 , \382 , \385 );
not \U$10 ( \387 , \386 );
nor \U$11 ( \388 , RIc224d60_87, RIc229fe0_151);
nor \U$12 ( \389 , RIc224ce8_88, RIc22a058_152);
nor \U$13 ( \390 , \388 , \389 );
or \U$14 ( \391 , RIc224e50_85, RIc229ef0_149);
nor \U$15 ( \392 , RIc224dd8_86, RIc229f68_150);
not \U$16 ( \393 , \392 );
nand \U$17 ( \394 , \390 , \391 , \393 );
not \U$18 ( \395 , \394 );
not \U$19 ( \396 , RIc224a90_93);
not \U$20 ( \397 , RIc22a2b0_157);
and \U$21 ( \398 , \396 , \397 );
nor \U$22 ( \399 , RIc224a18_94, RIc22a328_158);
nor \U$23 ( \400 , \398 , \399 );
nor \U$24 ( \401 , RIc2249a0_95, RIc22a3a0_159);
nor \U$25 ( \402 , RIc224928_96, RIc22a418_160);
nor \U$26 ( \403 , \401 , \402 );
nand \U$27 ( \404 , \400 , \403 );
not \U$28 ( \405 , RIc224bf8_90);
not \U$29 ( \406 , RIc22a148_154);
and \U$30 ( \407 , \405 , \406 );
nor \U$31 ( \408 , RIc224c70_89, RIc22a0d0_153);
nor \U$32 ( \409 , \407 , \408 );
nor \U$33 ( \410 , RIc224b80_91, RIc22a1c0_155);
nor \U$34 ( \411 , RIc224b08_92, RIc22a238_156);
nor \U$35 ( \412 , \410 , \411 );
nand \U$36 ( \413 , \409 , \412 );
nor \U$37 ( \414 , \404 , \413 );
and \U$38 ( \415 , \387 , \395 , \414 );
buf \U$39 ( \416 , \415 );
nor \U$40 ( \417 , RIc225300_75, RIc229a40_139);
nor \U$41 ( \418 , RIc225288_76, RIc229ab8_140);
nor \U$42 ( \419 , \417 , \418 );
not \U$43 ( \420 , \419 );
nor \U$44 ( \421 , RIc2253f0_73, RIc229950_137);
not \U$45 ( \422 , \421 );
or \U$46 ( \423 , RIc225378_74, RIc2299c8_138);
nand \U$47 ( \424 , \422 , \423 );
nor \U$48 ( \425 , \420 , \424 );
nor \U$49 ( \426 , RIc2250a8_80, RIc229c98_144);
nor \U$50 ( \427 , RIc225120_79, RIc229c20_143);
nor \U$51 ( \428 , \426 , \427 );
or \U$52 ( \429 , RIc225210_77, RIc229b30_141);
or \U$53 ( \430 , RIc225198_78, RIc229ba8_142);
and \U$54 ( \431 , \428 , \429 , \430 );
and \U$55 ( \432 , \425 , \431 );
not \U$56 ( \433 , \432 );
nor \U$57 ( \434 , RIc225558_70, RIc2297e8_134);
nor \U$58 ( \435 , RIc2255d0_69, RIc229770_133);
nor \U$59 ( \436 , \434 , \435 );
nor \U$60 ( \437 , RIc2254e0_71, RIc229860_135);
nor \U$61 ( \438 , RIc225468_72, RIc2298d8_136);
nor \U$62 ( \439 , \437 , \438 );
and \U$63 ( \440 , \436 , \439 );
nor \U$64 ( \441 , RIc225648_68, RIc2296f8_132);
not \U$65 ( \442 , \441 );
nand \U$66 ( \443 , \440 , \442 );
nor \U$67 ( \444 , \433 , \443 );
and \U$68 ( \445 , \416 , \444 );
not \U$69 ( \446 , \445 );
nand \U$70 ( \447 , RIc223f50_117, RIc22adf0_181);
nand \U$71 ( \448 , RIc223ed8_118, RIc22ae68_182);
and \U$72 ( \449 , \447 , \448 );
not \U$73 ( \450 , \449 );
nor \U$74 ( \451 , RIc223e60_119, RIc22aee0_183);
nand \U$75 ( \452 , RIc223de8_120, RIc22af58_184);
or \U$76 ( \453 , \451 , \452 );
nand \U$77 ( \454 , RIc223e60_119, RIc22aee0_183);
nand \U$78 ( \455 , \453 , \454 );
nor \U$79 ( \456 , RIc223ed8_118, RIc22ae68_182);
not \U$80 ( \457 , \456 );
nand \U$81 ( \458 , \455 , \457 );
not \U$82 ( \459 , \458 );
or \U$83 ( \460 , \450 , \459 );
nor \U$84 ( \461 , RIc224040_115, RIc22ad00_179);
not \U$85 ( \462 , \461 );
not \U$86 ( \463 , RIc22ad78_180);
not \U$87 ( \464 , RIc223fc8_116);
nand \U$88 ( \465 , \463 , \464 );
nand \U$89 ( \466 , \462 , \465 );
not \U$90 ( \467 , \466 );
not \U$91 ( \468 , RIc2240b8_114);
not \U$92 ( \469 , RIc22ac88_178);
and \U$93 ( \470 , \468 , \469 );
nor \U$94 ( \471 , RIc224130_113, RIc22ac10_177);
nor \U$95 ( \472 , \470 , \471 );
nand \U$96 ( \473 , \467 , \472 );
nor \U$97 ( \474 , RIc223f50_117, RIc22adf0_181);
buf \U$98 ( \475 , \474 );
nor \U$99 ( \476 , \473 , \475 );
nand \U$100 ( \477 , \460 , \476 );
not \U$101 ( \478 , \477 );
not \U$102 ( \479 , RIc223b90_125);
not \U$103 ( \480 , RIc22b1b0_189);
and \U$104 ( \481 , \479 , \480 );
nor \U$105 ( \482 , RIc2294a0_127, RIc22b2a0_191);
nor \U$106 ( \483 , \481 , \482 );
not \U$107 ( \484 , RIc2294a0_127);
not \U$108 ( \485 , RIc22b2a0_191);
or \U$109 ( \486 , \484 , \485 );
nand \U$110 ( \487 , RIc229518_128, RIc22b318_192);
nand \U$111 ( \488 , \486 , \487 );
not \U$112 ( \489 , RIc22b228_190);
not \U$113 ( \490 , RIc223b18_126);
nand \U$114 ( \491 , \489 , \490 );
nand \U$115 ( \492 , \483 , \488 , \491 );
nand \U$116 ( \493 , RIc223b18_126, RIc22b228_190);
not \U$117 ( \494 , \493 );
not \U$118 ( \495 , RIc223b90_125);
not \U$119 ( \496 , RIc22b1b0_189);
nand \U$120 ( \497 , \495 , \496 );
and \U$121 ( \498 , \494 , \497 );
nand \U$122 ( \499 , RIc223b90_125, RIc22b1b0_189);
not \U$123 ( \500 , \499 );
nor \U$124 ( \501 , \498 , \500 );
nand \U$125 ( \502 , \492 , \501 );
or \U$126 ( \503 , RIc223cf8_122, RIc22b048_186);
or \U$127 ( \504 , RIc2240b8_114, RIc22ac88_178);
or \U$128 ( \505 , RIc223fc8_116, RIc22ad78_180);
nand \U$129 ( \506 , \503 , \504 , \505 , \457 );
nor \U$130 ( \507 , RIc223d70_121, RIc22afd0_185);
not \U$131 ( \508 , \507 );
not \U$132 ( \509 , \474 );
not \U$133 ( \510 , \471 );
nand \U$134 ( \511 , \508 , \509 , \462 , \510 );
nor \U$135 ( \512 , RIc223de8_120, RIc22af58_184);
nor \U$136 ( \513 , \451 , \512 );
not \U$137 ( \514 , RIc223c80_123);
not \U$138 ( \515 , RIc22b0c0_187);
and \U$139 ( \516 , \514 , \515 );
nor \U$140 ( \517 , RIc223c08_124, RIc22b138_188);
nor \U$141 ( \518 , \516 , \517 );
nand \U$142 ( \519 , \513 , \518 );
nor \U$143 ( \520 , \506 , \511 , \519 );
nand \U$144 ( \521 , \502 , \520 );
not \U$145 ( \522 , \521 );
or \U$146 ( \523 , \478 , \522 );
not \U$147 ( \524 , RIc2245e0_103);
not \U$148 ( \525 , RIc22a760_167);
and \U$149 ( \526 , \524 , \525 );
nor \U$150 ( \527 , RIc224568_104, RIc22a7d8_168);
nor \U$151 ( \528 , \526 , \527 );
nor \U$152 ( \529 , RIc224658_102, RIc22a6e8_166);
nor \U$153 ( \530 , RIc2246d0_101, RIc22a670_165);
nor \U$154 ( \531 , \529 , \530 );
and \U$155 ( \532 , \528 , \531 );
nor \U$156 ( \533 , RIc224298_110, RIc22aaa8_174);
not \U$157 ( \534 , \533 );
not \U$158 ( \535 , RIc224310_109);
not \U$159 ( \536 , RIc22aa30_173);
and \U$160 ( \537 , \535 , \536 );
nor \U$161 ( \538 , RIc224220_111, RIc22ab20_175);
nor \U$162 ( \539 , \537 , \538 );
nor \U$163 ( \540 , RIc224388_108, RIc22a9b8_172);
not \U$164 ( \541 , \540 );
nand \U$165 ( \542 , \534 , \539 , \541 );
nor \U$166 ( \543 , RIc2241a8_112, RIc22ab98_176);
not \U$167 ( \544 , \543 );
or \U$168 ( \545 , RIc224478_106, RIc22a8c8_170);
or \U$169 ( \546 , RIc22a850_169, RIc2244f0_105);
or \U$170 ( \547 , RIc224400_107, RIc22a940_171);
nand \U$171 ( \548 , \544 , \545 , \546 , \547 );
nor \U$172 ( \549 , \542 , \548 );
nor \U$173 ( \550 , RIc2248b0_97, RIc22a490_161);
nor \U$174 ( \551 , RIc224838_98, RIc22a508_162);
nor \U$175 ( \552 , \550 , \551 );
nor \U$176 ( \553 , RIc2247c0_99, RIc22a580_163);
nor \U$177 ( \554 , RIc224748_100, RIc22a5f8_164);
nor \U$178 ( \555 , \553 , \554 );
nand \U$179 ( \556 , \552 , \555 );
not \U$180 ( \557 , \556 );
and \U$181 ( \558 , \532 , \549 , \557 );
nand \U$182 ( \559 , \523 , \558 );
nor \U$183 ( \560 , \451 , \512 );
nor \U$184 ( \561 , \474 , \456 );
nand \U$185 ( \562 , \560 , \561 );
nor \U$186 ( \563 , \473 , \562 );
nor \U$187 ( \564 , RIc223c80_123, RIc22b0c0_187);
nand \U$188 ( \565 , RIc223c08_124, RIc22b138_188);
or \U$189 ( \566 , \564 , \565 );
nand \U$190 ( \567 , RIc223c80_123, RIc22b0c0_187);
nand \U$191 ( \568 , \566 , \567 );
not \U$192 ( \569 , \568 );
not \U$193 ( \570 , RIc223cf8_122);
not \U$194 ( \571 , RIc22b048_186);
and \U$195 ( \572 , \570 , \571 );
nor \U$196 ( \573 , \572 , \507 );
not \U$197 ( \574 , \573 );
or \U$198 ( \575 , \569 , \574 );
not \U$199 ( \576 , \507 );
nand \U$200 ( \577 , RIc223cf8_122, RIc22b048_186);
not \U$201 ( \578 , \577 );
and \U$202 ( \579 , \576 , \578 );
nand \U$203 ( \580 , RIc223d70_121, RIc22afd0_185);
not \U$204 ( \581 , \580 );
nor \U$205 ( \582 , \579 , \581 );
nand \U$206 ( \583 , \575 , \582 );
nand \U$207 ( \584 , \563 , \583 );
not \U$208 ( \585 , \584 );
and \U$209 ( \586 , RIc223fc8_116, RIc22ad78_180);
not \U$210 ( \587 , \586 );
not \U$211 ( \588 , \462 );
or \U$212 ( \589 , \587 , \588 );
nand \U$213 ( \590 , RIc224040_115, RIc22ad00_179);
nand \U$214 ( \591 , \589 , \590 );
nand \U$215 ( \592 , \591 , \472 );
or \U$216 ( \593 , RIc224130_113, RIc22ac10_177);
nand \U$217 ( \594 , \593 , RIc2240b8_114, RIc22ac88_178);
nand \U$218 ( \595 , RIc224310_109, RIc22aa30_173);
nand \U$219 ( \596 , RIc224130_113, RIc22ac10_177);
and \U$220 ( \597 , \594 , \595 , \596 );
nand \U$221 ( \598 , \592 , \597 );
nor \U$222 ( \599 , RIc224220_111, RIc22ab20_175);
nand \U$223 ( \600 , RIc2241a8_112, RIc22ab98_176);
nor \U$224 ( \601 , \599 , \600 );
not \U$225 ( \602 , \601 );
nor \U$226 ( \603 , RIc224310_109, RIc22aa30_173);
nor \U$227 ( \604 , \603 , \533 );
not \U$228 ( \605 , \604 );
or \U$229 ( \606 , \602 , \605 );
nand \U$230 ( \607 , RIc224220_111, RIc22ab20_175);
nand \U$231 ( \608 , RIc224298_110, RIc22aaa8_174);
nand \U$232 ( \609 , \607 , \608 );
nand \U$233 ( \610 , \604 , \609 );
nand \U$234 ( \611 , \606 , \610 );
nor \U$235 ( \612 , \598 , \611 );
not \U$236 ( \613 , \612 );
or \U$237 ( \614 , \585 , \613 );
and \U$238 ( \615 , \595 , \607 , \608 );
not \U$239 ( \616 , \615 );
nor \U$240 ( \617 , \543 , \533 );
nand \U$241 ( \618 , \617 , \539 );
not \U$242 ( \619 , \618 );
or \U$243 ( \620 , \616 , \619 );
not \U$244 ( \621 , \603 );
not \U$245 ( \622 , \621 );
not \U$246 ( \623 , \534 );
or \U$247 ( \624 , \622 , \623 );
nand \U$248 ( \625 , \624 , \595 );
nand \U$249 ( \626 , \620 , \625 );
not \U$250 ( \627 , RIc224400_107);
not \U$251 ( \628 , RIc22a940_171);
and \U$252 ( \629 , \627 , \628 );
nor \U$253 ( \630 , \629 , \540 );
not \U$254 ( \631 , RIc224478_106);
not \U$255 ( \632 , RIc22a8c8_170);
and \U$256 ( \633 , \631 , \632 );
nor \U$257 ( \634 , RIc2244f0_105, RIc22a850_169);
nor \U$258 ( \635 , \633 , \634 );
and \U$259 ( \636 , \630 , \635 );
nand \U$260 ( \637 , \532 , \636 , \557 );
nor \U$261 ( \638 , \626 , \637 );
nand \U$262 ( \639 , \614 , \638 );
nor \U$263 ( \640 , \556 , \530 );
not \U$264 ( \641 , \640 );
and \U$265 ( \642 , RIc224568_104, RIc22a7d8_168);
not \U$266 ( \643 , \642 );
or \U$267 ( \644 , RIc22a760_167, RIc2245e0_103);
not \U$268 ( \645 , \644 );
or \U$269 ( \646 , \643 , \645 );
nand \U$270 ( \647 , RIc2245e0_103, RIc22a760_167);
nand \U$271 ( \648 , \646 , \647 );
not \U$272 ( \649 , \529 );
nand \U$273 ( \650 , \648 , \649 );
nand \U$274 ( \651 , RIc2246d0_101, RIc22a670_165);
nand \U$275 ( \652 , RIc224658_102, RIc22a6e8_166);
and \U$276 ( \653 , \651 , \652 );
nand \U$277 ( \654 , \650 , \653 );
not \U$278 ( \655 , \654 );
or \U$279 ( \656 , \641 , \655 );
nand \U$280 ( \657 , RIc224748_100, RIc22a5f8_164);
or \U$281 ( \658 , \553 , \657 );
nand \U$282 ( \659 , RIc2247c0_99, RIc22a580_163);
nand \U$283 ( \660 , \658 , \659 );
and \U$284 ( \661 , \660 , \552 );
nand \U$285 ( \662 , RIc224838_98, RIc22a508_162);
or \U$286 ( \663 , \550 , \662 );
nand \U$287 ( \664 , RIc2248b0_97, RIc22a490_161);
nand \U$288 ( \665 , \663 , \664 );
nor \U$289 ( \666 , \661 , \665 );
nand \U$290 ( \667 , \656 , \666 );
not \U$291 ( \668 , \667 );
not \U$292 ( \669 , \635 );
and \U$293 ( \670 , RIc224388_108, RIc22a9b8_172);
not \U$294 ( \671 , \670 );
not \U$295 ( \672 , \547 );
or \U$296 ( \673 , \671 , \672 );
nand \U$297 ( \674 , RIc224400_107, RIc22a940_171);
nand \U$298 ( \675 , \673 , \674 );
not \U$299 ( \676 , \675 );
or \U$300 ( \677 , \669 , \676 );
not \U$301 ( \678 , \634 );
nand \U$302 ( \679 , RIc224478_106, RIc22a8c8_170);
not \U$303 ( \680 , \679 );
and \U$304 ( \681 , \678 , \680 );
and \U$305 ( \682 , RIc2244f0_105, RIc22a850_169);
nor \U$306 ( \683 , \681 , \682 );
nand \U$307 ( \684 , \677 , \683 );
buf \U$308 ( \685 , \532 );
nand \U$309 ( \686 , \684 , \685 , \557 );
nand \U$310 ( \687 , \559 , \639 , \668 , \686 );
buf \U$311 ( \688 , \687 );
not \U$312 ( \689 , \688 );
or \U$313 ( \690 , \446 , \689 );
nand \U$314 ( \691 , RIc224b08_92, RIc22a238_156);
or \U$315 ( \692 , \410 , \691 );
nand \U$316 ( \693 , RIc224b80_91, RIc22a1c0_155);
nand \U$317 ( \694 , \692 , \693 );
and \U$318 ( \695 , \694 , \409 );
nand \U$319 ( \696 , RIc224bf8_90, RIc22a148_154);
or \U$320 ( \697 , \408 , \696 );
nand \U$321 ( \698 , RIc224c70_89, RIc22a0d0_153);
nand \U$322 ( \699 , \697 , \698 );
nor \U$323 ( \700 , \695 , \699 );
nand \U$324 ( \701 , RIc224a18_94, RIc22a328_158);
nand \U$325 ( \702 , RIc224a90_93, RIc22a2b0_157);
nand \U$326 ( \703 , RIc2249a0_95, RIc22a3a0_159);
nand \U$327 ( \704 , \701 , \702 , \703 );
not \U$328 ( \705 , \704 );
nand \U$329 ( \706 , RIc224928_96, RIc22a418_160);
or \U$330 ( \707 , \401 , \706 );
nand \U$331 ( \708 , \705 , \707 );
or \U$332 ( \709 , RIc224a90_93, RIc22a2b0_157);
not \U$333 ( \710 , \709 );
or \U$334 ( \711 , RIc224a18_94, RIc22a328_158);
not \U$335 ( \712 , \711 );
or \U$336 ( \713 , \710 , \712 );
nand \U$337 ( \714 , \713 , \702 );
or \U$338 ( \715 , \408 , \410 );
or \U$339 ( \716 , RIc224bf8_90, RIc22a148_154);
or \U$340 ( \717 , RIc224b08_92, RIc22a238_156);
nand \U$341 ( \718 , \716 , \717 );
nor \U$342 ( \719 , \715 , \718 );
nand \U$343 ( \720 , \708 , \714 , \719 );
nand \U$344 ( \721 , \700 , \720 );
not \U$345 ( \722 , \721 );
nor \U$346 ( \723 , \386 , \394 );
not \U$347 ( \724 , \723 );
or \U$348 ( \725 , \722 , \724 );
nor \U$349 ( \726 , RIc224e50_85, RIc229ef0_149);
nor \U$350 ( \727 , \726 , \392 );
not \U$351 ( \728 , \727 );
nand \U$352 ( \729 , RIc224ce8_88, RIc22a058_152);
or \U$353 ( \730 , \388 , \729 );
nand \U$354 ( \731 , RIc224d60_87, RIc229fe0_151);
nand \U$355 ( \732 , \730 , \731 );
not \U$356 ( \733 , \732 );
or \U$357 ( \734 , \728 , \733 );
nand \U$358 ( \735 , RIc224dd8_86, RIc229f68_150);
not \U$359 ( \736 , \735 );
and \U$360 ( \737 , \391 , \736 );
and \U$361 ( \738 , RIc224e50_85, RIc229ef0_149);
nor \U$362 ( \739 , \737 , \738 );
nand \U$363 ( \740 , \734 , \739 );
and \U$364 ( \741 , \740 , \387 );
not \U$365 ( \742 , \385 );
not \U$366 ( \743 , RIc224ec8_84);
not \U$367 ( \744 , RIc229e78_148);
nor \U$368 ( \745 , \743 , \744 );
not \U$369 ( \746 , \745 );
or \U$370 ( \747 , RIc224f40_83, RIc229e00_147);
not \U$371 ( \748 , \747 );
or \U$372 ( \749 , \746 , \748 );
nand \U$373 ( \750 , RIc224f40_83, RIc229e00_147);
nand \U$374 ( \751 , \749 , \750 );
not \U$375 ( \752 , \751 );
or \U$376 ( \753 , \742 , \752 );
nand \U$377 ( \754 , RIc224fb8_82, RIc229d88_146);
not \U$378 ( \755 , \754 );
not \U$379 ( \756 , \384 );
and \U$380 ( \757 , \755 , \756 );
and \U$381 ( \758 , RIc225030_81, RIc229d10_145);
nor \U$382 ( \759 , \757 , \758 );
nand \U$383 ( \760 , \753 , \759 );
nor \U$384 ( \761 , \741 , \760 );
nand \U$385 ( \762 , \725 , \761 );
buf \U$386 ( \763 , \762 );
nor \U$387 ( \764 , \433 , \443 );
and \U$388 ( \765 , \763 , \764 );
not \U$389 ( \766 , \443 );
not \U$390 ( \767 , \766 );
not \U$391 ( \768 , \425 );
not \U$392 ( \769 , \429 );
not \U$393 ( \770 , \430 );
nor \U$394 ( \771 , \769 , \770 );
not \U$395 ( \772 , \771 );
nand \U$396 ( \773 , RIc2250a8_80, RIc229c98_144);
or \U$397 ( \774 , \427 , \773 );
nand \U$398 ( \775 , RIc225120_79, RIc229c20_143);
nand \U$399 ( \776 , \774 , \775 );
not \U$400 ( \777 , \776 );
or \U$401 ( \778 , \772 , \777 );
nand \U$402 ( \779 , RIc225198_78, RIc229ba8_142);
not \U$403 ( \780 , \779 );
and \U$404 ( \781 , \429 , \780 );
nand \U$405 ( \782 , RIc225210_77, RIc229b30_141);
not \U$406 ( \783 , \782 );
nor \U$407 ( \784 , \781 , \783 );
nand \U$408 ( \785 , \778 , \784 );
not \U$409 ( \786 , \785 );
or \U$410 ( \787 , \768 , \786 );
not \U$411 ( \788 , \424 );
not \U$412 ( \789 , \788 );
nand \U$413 ( \790 , RIc225288_76, RIc229ab8_140);
not \U$414 ( \791 , \790 );
not \U$415 ( \792 , \791 );
not \U$416 ( \793 , \417 );
not \U$417 ( \794 , \793 );
or \U$418 ( \795 , \792 , \794 );
nand \U$419 ( \796 , RIc225300_75, RIc229a40_139);
nand \U$420 ( \797 , \795 , \796 );
not \U$421 ( \798 , \797 );
or \U$422 ( \799 , \789 , \798 );
not \U$423 ( \800 , \421 );
nand \U$424 ( \801 , RIc225378_74, RIc2299c8_138);
not \U$425 ( \802 , \801 );
and \U$426 ( \803 , \800 , \802 );
and \U$427 ( \804 , RIc2253f0_73, RIc229950_137);
nor \U$428 ( \805 , \803 , \804 );
nand \U$429 ( \806 , \799 , \805 );
not \U$430 ( \807 , \806 );
nand \U$431 ( \808 , \787 , \807 );
not \U$432 ( \809 , \808 );
or \U$433 ( \810 , \767 , \809 );
not \U$434 ( \811 , \436 );
nand \U$435 ( \812 , RIc225468_72, RIc2298d8_136);
or \U$436 ( \813 , \437 , \812 );
nand \U$437 ( \814 , RIc2254e0_71, RIc229860_135);
nand \U$438 ( \815 , \813 , \814 );
not \U$439 ( \816 , \815 );
or \U$440 ( \817 , \811 , \816 );
not \U$441 ( \818 , \435 );
nand \U$442 ( \819 , RIc225558_70, RIc2297e8_134);
not \U$443 ( \820 , \819 );
and \U$444 ( \821 , \818 , \820 );
and \U$445 ( \822 , RIc2255d0_69, RIc229770_133);
nor \U$446 ( \823 , \821 , \822 );
nand \U$447 ( \824 , \817 , \823 );
and \U$448 ( \825 , \824 , \442 );
and \U$449 ( \826 , RIc225648_68, RIc2296f8_132);
nor \U$450 ( \827 , \825 , \826 );
nand \U$451 ( \828 , \810 , \827 );
nor \U$452 ( \829 , \765 , \828 );
nand \U$453 ( \830 , \690 , \829 );
nor \U$454 ( \831 , RIc2256c0_67, RIc229680_131);
not \U$455 ( \832 , \831 );
nand \U$456 ( \833 , RIc2256c0_67, RIc229680_131);
nand \U$457 ( \834 , \832 , \833 );
not \U$458 ( \835 , \834 );
and \U$459 ( \836 , \830 , \835 );
not \U$460 ( \837 , \830 );
and \U$461 ( \838 , \837 , \834 );
nor \U$462 ( \839 , \836 , \838 );
buf \U$463 ( \840 , \839 );
buf \U$464 ( \841 , \840 );
not \U$465 ( \842 , \841 );
xor \U$466 ( \843 , \842 , RIc2275b0_1);
not \U$467 ( \844 , RIc227538_2);
and \U$468 ( \845 , RIc2274c0_3, \844 );
not \U$469 ( \846 , RIc2274c0_3);
and \U$470 ( \847 , \846 , RIc227538_2);
nor \U$471 ( \848 , \845 , \847 );
and \U$472 ( \849 , RIc2275b0_1, RIc227538_2);
not \U$473 ( \850 , RIc2275b0_1);
and \U$474 ( \851 , \850 , \844 );
nor \U$475 ( \852 , \849 , \851 );
and \U$476 ( \853 , \848 , \852 );
buf \U$477 ( \854 , \853 );
not \U$478 ( \855 , \854 );
or \U$479 ( \856 , \843 , \855 );
nor \U$480 ( \857 , \831 , \441 );
nand \U$481 ( \858 , \440 , \857 );
nor \U$482 ( \859 , \433 , \858 );
and \U$483 ( \860 , \416 , \859 );
not \U$484 ( \861 , \860 );
not \U$485 ( \862 , \688 );
or \U$486 ( \863 , \861 , \862 );
nor \U$487 ( \864 , \433 , \858 );
and \U$488 ( \865 , \763 , \864 );
not \U$489 ( \866 , \858 );
not \U$490 ( \867 , \866 );
not \U$491 ( \868 , \808 );
or \U$492 ( \869 , \867 , \868 );
and \U$493 ( \870 , \824 , \857 );
not \U$494 ( \871 , \826 );
not \U$495 ( \872 , \832 );
or \U$496 ( \873 , \871 , \872 );
nand \U$497 ( \874 , \873 , \833 );
nor \U$498 ( \875 , \870 , \874 );
nand \U$499 ( \876 , \869 , \875 );
nor \U$500 ( \877 , \865 , \876 );
nand \U$501 ( \878 , \863 , \877 );
nor \U$502 ( \879 , RIc225738_66, RIc229608_130);
not \U$503 ( \880 , \879 );
nand \U$504 ( \881 , RIc225738_66, RIc229608_130);
nand \U$505 ( \882 , \880 , \881 );
not \U$506 ( \883 , \882 );
and \U$507 ( \884 , \878 , \883 );
not \U$508 ( \885 , \878 );
and \U$509 ( \886 , \885 , \882 );
nor \U$510 ( \887 , \884 , \886 );
buf \U$511 ( \888 , \887 );
buf \U$512 ( \889 , \888 );
not \U$513 ( \890 , \889 );
not \U$514 ( \891 , \890 );
buf \U$515 ( \892 , \891 );
not \U$516 ( \893 , \892 );
and \U$517 ( \894 , RIc2275b0_1, \893 );
not \U$518 ( \895 , RIc2275b0_1);
and \U$519 ( \896 , \895 , \892 );
nor \U$520 ( \897 , \894 , \896 );
not \U$521 ( \898 , \848 );
not \U$522 ( \899 , \898 );
or \U$523 ( \900 , \897 , \899 );
nand \U$524 ( \901 , \856 , \900 );
not \U$525 ( \902 , \416 );
nor \U$526 ( \903 , RIc2257b0_65, RIc229590_129);
nor \U$527 ( \904 , \879 , \903 );
and \U$528 ( \905 , \857 , \904 );
and \U$529 ( \906 , \440 , \905 );
nand \U$530 ( \907 , \432 , \906 );
nor \U$531 ( \908 , \902 , \907 );
not \U$532 ( \909 , \908 );
not \U$533 ( \910 , \688 );
or \U$534 ( \911 , \909 , \910 );
not \U$535 ( \912 , \907 );
not \U$536 ( \913 , \912 );
not \U$537 ( \914 , \763 );
or \U$538 ( \915 , \913 , \914 );
and \U$539 ( \916 , \808 , \906 );
not \U$540 ( \917 , \905 );
not \U$541 ( \918 , \824 );
or \U$542 ( \919 , \917 , \918 );
and \U$543 ( \920 , \874 , \904 );
or \U$544 ( \921 , \903 , \881 );
nand \U$545 ( \922 , RIc2257b0_65, RIc229590_129);
nand \U$546 ( \923 , \921 , \922 );
nor \U$547 ( \924 , \920 , \923 );
nand \U$548 ( \925 , \919 , \924 );
nor \U$549 ( \926 , \916 , \925 );
nand \U$550 ( \927 , \915 , \926 );
not \U$551 ( \928 , \927 );
nand \U$552 ( \929 , \911 , \928 );
buf \U$553 ( \930 , \929 );
buf \U$554 ( \931 , \930 );
not \U$555 ( \932 , \931 );
and \U$556 ( \933 , \932 , RIc2273d0_5);
not \U$557 ( \934 , \932 );
not \U$558 ( \935 , RIc2273d0_5);
and \U$559 ( \936 , \934 , \935 );
nor \U$560 ( \937 , \933 , \936 );
and \U$561 ( \938 , RIc227358_6, RIc2272e0_7);
not \U$562 ( \939 , RIc227358_6);
not \U$563 ( \940 , RIc2272e0_7);
and \U$564 ( \941 , \939 , \940 );
nor \U$565 ( \942 , \938 , \941 );
not \U$566 ( \943 , \942 );
and \U$567 ( \944 , RIc227358_6, RIc2273d0_5);
not \U$568 ( \945 , RIc227358_6);
not \U$569 ( \946 , RIc2273d0_5);
and \U$570 ( \947 , \945 , \946 );
nor \U$571 ( \948 , \944 , \947 );
nand \U$572 ( \949 , \943 , \948 );
not \U$573 ( \950 , \949 );
buf \U$574 ( \951 , \950 );
not \U$575 ( \952 , \951 );
or \U$576 ( \953 , \937 , \952 );
buf \U$577 ( \954 , \942 );
not \U$578 ( \955 , \954 );
not \U$579 ( \956 , RIc2273d0_5);
or \U$580 ( \957 , \955 , \956 );
nand \U$581 ( \958 , \953 , \957 );
xor \U$582 ( \959 , \901 , \958 );
not \U$583 ( \960 , \440 );
nor \U$584 ( \961 , \433 , \960 );
and \U$585 ( \962 , \416 , \961 );
not \U$586 ( \963 , \962 );
not \U$587 ( \964 , \688 );
or \U$588 ( \965 , \963 , \964 );
nor \U$589 ( \966 , \433 , \960 );
and \U$590 ( \967 , \763 , \966 );
not \U$591 ( \968 , \440 );
not \U$592 ( \969 , \808 );
or \U$593 ( \970 , \968 , \969 );
not \U$594 ( \971 , \824 );
nand \U$595 ( \972 , \970 , \971 );
nor \U$596 ( \973 , \967 , \972 );
nand \U$597 ( \974 , \965 , \973 );
nor \U$598 ( \975 , \826 , \441 );
and \U$599 ( \976 , \974 , \975 );
not \U$600 ( \977 , \974 );
not \U$601 ( \978 , \975 );
and \U$602 ( \979 , \977 , \978 );
nor \U$603 ( \980 , \976 , \979 );
buf \U$604 ( \981 , \980 );
not \U$605 ( \982 , \981 );
buf \U$606 ( \983 , \982 );
not \U$607 ( \984 , \983 );
buf \U$608 ( \985 , \984 );
not \U$609 ( \986 , \985 );
and \U$610 ( \987 , RIc2275b0_1, \986 );
not \U$611 ( \988 , RIc2275b0_1);
and \U$612 ( \989 , \988 , \985 );
nor \U$613 ( \990 , \987 , \989 );
or \U$614 ( \991 , \990 , \855 );
or \U$615 ( \992 , \843 , \899 );
nand \U$616 ( \993 , \991 , \992 );
not \U$617 ( \994 , RIc2275b0_1);
not \U$618 ( \995 , \434 );
nand \U$619 ( \996 , \439 , \995 );
nor \U$620 ( \997 , \433 , \996 );
and \U$621 ( \998 , \416 , \997 );
not \U$622 ( \999 , \998 );
not \U$623 ( \1000 , \688 );
or \U$624 ( \1001 , \999 , \1000 );
nor \U$625 ( \1002 , \433 , \996 );
and \U$626 ( \1003 , \763 , \1002 );
not \U$627 ( \1004 , \996 );
not \U$628 ( \1005 , \1004 );
not \U$629 ( \1006 , \808 );
or \U$630 ( \1007 , \1005 , \1006 );
and \U$631 ( \1008 , \815 , \995 );
not \U$632 ( \1009 , \819 );
nor \U$633 ( \1010 , \1008 , \1009 );
nand \U$634 ( \1011 , \1007 , \1010 );
nor \U$635 ( \1012 , \1003 , \1011 );
nand \U$636 ( \1013 , \1001 , \1012 );
nor \U$637 ( \1014 , \435 , \822 );
and \U$638 ( \1015 , \1013 , \1014 );
not \U$639 ( \1016 , \1013 );
not \U$640 ( \1017 , \1014 );
and \U$641 ( \1018 , \1016 , \1017 );
nor \U$642 ( \1019 , \1015 , \1018 );
buf \U$643 ( \1020 , \1019 );
not \U$644 ( \1021 , \1020 );
buf \U$645 ( \1022 , \1021 );
nor \U$646 ( \1023 , \994 , \1022 );
xor \U$647 ( \1024 , \993 , \1023 );
and \U$648 ( \1025 , \893 , RIc2274c0_3);
not \U$649 ( \1026 , \893 );
not \U$650 ( \1027 , RIc2274c0_3);
and \U$651 ( \1028 , \1026 , \1027 );
nor \U$652 ( \1029 , \1025 , \1028 );
and \U$653 ( \1030 , RIc227448_4, RIc2274c0_3);
not \U$654 ( \1031 , RIc227448_4);
not \U$655 ( \1032 , RIc2274c0_3);
and \U$656 ( \1033 , \1031 , \1032 );
nor \U$657 ( \1034 , \1030 , \1033 );
and \U$658 ( \1035 , RIc227448_4, \946 );
not \U$659 ( \1036 , RIc227448_4);
and \U$660 ( \1037 , \1036 , RIc2273d0_5);
nor \U$661 ( \1038 , \1035 , \1037 );
and \U$662 ( \1039 , \1034 , \1038 );
buf \U$663 ( \1040 , \1039 );
not \U$664 ( \1041 , \1040 );
or \U$665 ( \1042 , \1029 , \1041 );
not \U$666 ( \1043 , \857 );
nor \U$667 ( \1044 , \1043 , \879 );
and \U$668 ( \1045 , \440 , \1044 );
nand \U$669 ( \1046 , \432 , \1045 );
nor \U$670 ( \1047 , \902 , \1046 );
not \U$671 ( \1048 , \1047 );
not \U$672 ( \1049 , \688 );
or \U$673 ( \1050 , \1048 , \1049 );
not \U$674 ( \1051 , \1046 );
and \U$675 ( \1052 , \763 , \1051 );
not \U$676 ( \1053 , \1045 );
not \U$677 ( \1054 , \808 );
or \U$678 ( \1055 , \1053 , \1054 );
and \U$679 ( \1056 , \824 , \1044 );
not \U$680 ( \1057 , \880 );
not \U$681 ( \1058 , \874 );
or \U$682 ( \1059 , \1057 , \1058 );
nand \U$683 ( \1060 , \1059 , \881 );
nor \U$684 ( \1061 , \1056 , \1060 );
nand \U$685 ( \1062 , \1055 , \1061 );
nor \U$686 ( \1063 , \1052 , \1062 );
nand \U$687 ( \1064 , \1050 , \1063 );
not \U$688 ( \1065 , \903 );
nand \U$689 ( \1066 , \1065 , \922 );
not \U$690 ( \1067 , \1066 );
and \U$691 ( \1068 , \1064 , \1067 );
not \U$692 ( \1069 , \1064 );
and \U$693 ( \1070 , \1069 , \1066 );
nor \U$694 ( \1071 , \1068 , \1070 );
buf \U$695 ( \1072 , \1071 );
buf \U$696 ( \1073 , \1072 );
not \U$697 ( \1074 , \1073 );
buf \U$698 ( \1075 , \1074 );
and \U$699 ( \1076 , \1075 , RIc2274c0_3);
not \U$700 ( \1077 , \1075 );
not \U$701 ( \1078 , RIc2274c0_3);
and \U$702 ( \1079 , \1077 , \1078 );
nor \U$703 ( \1080 , \1076 , \1079 );
not \U$704 ( \1081 , \1038 );
buf \U$705 ( \1082 , \1081 );
not \U$706 ( \1083 , \1082 );
or \U$707 ( \1084 , \1080 , \1083 );
nand \U$708 ( \1085 , \1042 , \1084 );
and \U$709 ( \1086 , \1024 , \1085 );
and \U$710 ( \1087 , \993 , \1023 );
or \U$711 ( \1088 , \1086 , \1087 );
xor \U$712 ( \1089 , \959 , \1088 );
not \U$713 ( \1090 , RIc2275b0_1);
nor \U$714 ( \1091 , \1090 , \986 );
or \U$715 ( \1092 , \951 , \954 );
nand \U$716 ( \1093 , \1092 , RIc2273d0_5);
xor \U$717 ( \1094 , \1091 , \1093 );
or \U$718 ( \1095 , \1080 , \1041 );
and \U$719 ( \1096 , \932 , RIc2274c0_3);
not \U$720 ( \1097 , \932 );
and \U$721 ( \1098 , \1097 , \1032 );
nor \U$722 ( \1099 , \1096 , \1098 );
or \U$723 ( \1100 , \1099 , \1083 );
nand \U$724 ( \1101 , \1095 , \1100 );
xor \U$725 ( \1102 , \1094 , \1101 );
and \U$726 ( \1103 , \1074 , RIc2273d0_5);
and \U$727 ( \1104 , \1073 , \946 );
nor \U$728 ( \1105 , \1103 , \1104 );
or \U$729 ( \1106 , \1105 , \952 );
or \U$730 ( \1107 , \937 , \955 );
nand \U$731 ( \1108 , \1106 , \1107 );
not \U$732 ( \1109 , RIc227268_8);
and \U$733 ( \1110 , RIc2271f0_9, \1109 );
not \U$734 ( \1111 , RIc2271f0_9);
and \U$735 ( \1112 , \1111 , RIc227268_8);
nor \U$736 ( \1113 , \1110 , \1112 );
and \U$737 ( \1114 , \940 , \1109 );
and \U$738 ( \1115 , RIc2272e0_7, RIc227268_8);
nor \U$739 ( \1116 , \1114 , \1115 );
nand \U$740 ( \1117 , \1113 , \1116 );
not \U$741 ( \1118 , \1117 );
buf \U$742 ( \1119 , \1113 );
not \U$743 ( \1120 , \1119 );
buf \U$744 ( \1121 , \1120 );
or \U$745 ( \1122 , \1118 , \1121 );
nand \U$746 ( \1123 , \1122 , RIc2272e0_7);
xor \U$747 ( \1124 , \1108 , \1123 );
and \U$748 ( \1125 , RIc2275b0_1, \1022 );
not \U$749 ( \1126 , RIc2275b0_1);
not \U$750 ( \1127 , \1022 );
and \U$751 ( \1128 , \1126 , \1127 );
nor \U$752 ( \1129 , \1125 , \1128 );
or \U$753 ( \1130 , \1129 , \855 );
or \U$754 ( \1131 , \990 , \899 );
nand \U$755 ( \1132 , \1130 , \1131 );
and \U$756 ( \1133 , \1124 , \1132 );
and \U$757 ( \1134 , \1108 , \1123 );
or \U$758 ( \1135 , \1133 , \1134 );
not \U$759 ( \1136 , \958 );
xor \U$760 ( \1137 , \1135 , \1136 );
and \U$761 ( \1138 , \932 , RIc2272e0_7);
not \U$762 ( \1139 , RIc2272e0_7);
and \U$763 ( \1140 , \931 , \1139 );
nor \U$764 ( \1141 , \1138 , \1140 );
not \U$765 ( \1142 , \1141 );
and \U$766 ( \1143 , \1142 , \1118 );
and \U$767 ( \1144 , \1121 , RIc2272e0_7);
nor \U$768 ( \1145 , \1143 , \1144 );
not \U$769 ( \1146 , \1145 );
not \U$770 ( \1147 , RIc2275b0_1);
not \U$771 ( \1148 , \439 );
nor \U$772 ( \1149 , \433 , \1148 );
and \U$773 ( \1150 , \416 , \1149 );
not \U$774 ( \1151 , \1150 );
not \U$775 ( \1152 , \688 );
or \U$776 ( \1153 , \1151 , \1152 );
nor \U$777 ( \1154 , \433 , \1148 );
and \U$778 ( \1155 , \763 , \1154 );
not \U$779 ( \1156 , \439 );
not \U$780 ( \1157 , \808 );
or \U$781 ( \1158 , \1156 , \1157 );
not \U$782 ( \1159 , \815 );
nand \U$783 ( \1160 , \1158 , \1159 );
nor \U$784 ( \1161 , \1155 , \1160 );
nand \U$785 ( \1162 , \1153 , \1161 );
nand \U$786 ( \1163 , \995 , \819 );
not \U$787 ( \1164 , \1163 );
and \U$788 ( \1165 , \1162 , \1164 );
not \U$789 ( \1166 , \1162 );
and \U$790 ( \1167 , \1166 , \1163 );
nor \U$791 ( \1168 , \1165 , \1167 );
buf \U$792 ( \1169 , \1168 );
not \U$793 ( \1170 , \1169 );
buf \U$794 ( \1171 , \1170 );
nor \U$795 ( \1172 , \1147 , \1171 );
xor \U$796 ( \1173 , \1146 , \1172 );
and \U$797 ( \1174 , \842 , RIc2274c0_3);
not \U$798 ( \1175 , \842 );
and \U$799 ( \1176 , \1175 , \1032 );
nor \U$800 ( \1177 , \1174 , \1176 );
or \U$801 ( \1178 , \1177 , \1041 );
or \U$802 ( \1179 , \1029 , \1083 );
nand \U$803 ( \1180 , \1178 , \1179 );
and \U$804 ( \1181 , \1173 , \1180 );
and \U$805 ( \1182 , \1146 , \1172 );
or \U$806 ( \1183 , \1181 , \1182 );
and \U$807 ( \1184 , \1137 , \1183 );
and \U$808 ( \1185 , \1135 , \1136 );
or \U$809 ( \1186 , \1184 , \1185 );
xor \U$810 ( \1187 , \1102 , \1186 );
xor \U$811 ( \1188 , \1089 , \1187 );
xor \U$812 ( \1189 , \993 , \1023 );
xor \U$813 ( \1190 , \1189 , \1085 );
xor \U$814 ( \1191 , \1135 , \1136 );
xor \U$815 ( \1192 , \1191 , \1183 );
and \U$816 ( \1193 , \1190 , \1192 );
and \U$817 ( \1194 , \893 , RIc2273d0_5);
and \U$818 ( \1195 , \889 , \946 );
nor \U$819 ( \1196 , \1194 , \1195 );
or \U$820 ( \1197 , \1196 , \952 );
or \U$821 ( \1198 , \1105 , \955 );
nand \U$822 ( \1199 , \1197 , \1198 );
not \U$823 ( \1200 , \438 );
nand \U$824 ( \1201 , \432 , \1200 );
nor \U$825 ( \1202 , \902 , \1201 );
not \U$826 ( \1203 , \1202 );
not \U$827 ( \1204 , \688 );
or \U$828 ( \1205 , \1203 , \1204 );
not \U$829 ( \1206 , \1201 );
and \U$830 ( \1207 , \763 , \1206 );
not \U$831 ( \1208 , \1200 );
not \U$832 ( \1209 , \808 );
or \U$833 ( \1210 , \1208 , \1209 );
nand \U$834 ( \1211 , \1210 , \812 );
nor \U$835 ( \1212 , \1207 , \1211 );
nand \U$836 ( \1213 , \1205 , \1212 );
not \U$837 ( \1214 , \814 );
nor \U$838 ( \1215 , \1214 , \437 );
and \U$839 ( \1216 , \1213 , \1215 );
not \U$840 ( \1217 , \1213 );
not \U$841 ( \1218 , \1215 );
and \U$842 ( \1219 , \1217 , \1218 );
nor \U$843 ( \1220 , \1216 , \1219 );
not \U$844 ( \1221 , \1220 );
buf \U$845 ( \1222 , \1221 );
not \U$846 ( \1223 , \1222 );
and \U$847 ( \1224 , \1223 , RIc2275b0_1);
xor \U$848 ( \1225 , \1199 , \1224 );
and \U$849 ( \1226 , RIc2275b0_1, \1171 );
not \U$850 ( \1227 , RIc2275b0_1);
not \U$851 ( \1228 , \1171 );
and \U$852 ( \1229 , \1227 , \1228 );
nor \U$853 ( \1230 , \1226 , \1229 );
or \U$854 ( \1231 , \1230 , \855 );
or \U$855 ( \1232 , \1129 , \899 );
nand \U$856 ( \1233 , \1231 , \1232 );
and \U$857 ( \1234 , \1225 , \1233 );
and \U$858 ( \1235 , \1199 , \1224 );
or \U$859 ( \1236 , \1234 , \1235 );
xor \U$860 ( \1237 , \1146 , \1172 );
xor \U$861 ( \1238 , \1237 , \1180 );
xor \U$862 ( \1239 , \1236 , \1238 );
xor \U$863 ( \1240 , \1108 , \1123 );
xor \U$864 ( \1241 , \1240 , \1132 );
and \U$865 ( \1242 , \1239 , \1241 );
and \U$866 ( \1243 , \1236 , \1238 );
or \U$867 ( \1244 , \1242 , \1243 );
xor \U$868 ( \1245 , \1135 , \1136 );
xor \U$869 ( \1246 , \1245 , \1183 );
and \U$870 ( \1247 , \1244 , \1246 );
and \U$871 ( \1248 , \1190 , \1244 );
or \U$872 ( \1249 , \1193 , \1247 , \1248 );
or \U$873 ( \1250 , \1188 , \1249 );
not \U$874 ( \1251 , \1250 );
xor \U$875 ( \1252 , \901 , \958 );
xor \U$876 ( \1253 , \1252 , \1088 );
and \U$877 ( \1254 , \1102 , \1253 );
xor \U$878 ( \1255 , \901 , \958 );
xor \U$879 ( \1256 , \1255 , \1088 );
and \U$880 ( \1257 , \1186 , \1256 );
and \U$881 ( \1258 , \1102 , \1186 );
or \U$882 ( \1259 , \1254 , \1257 , \1258 );
not \U$883 ( \1260 , \1099 );
not \U$884 ( \1261 , \1041 );
and \U$885 ( \1262 , \1260 , \1261 );
and \U$886 ( \1263 , \1082 , RIc2274c0_3);
nor \U$887 ( \1264 , \1262 , \1263 );
not \U$888 ( \1265 , RIc2275b0_1);
nor \U$889 ( \1266 , \1265 , \842 );
xor \U$890 ( \1267 , \1264 , \1266 );
or \U$891 ( \1268 , \897 , \855 );
and \U$892 ( \1269 , RIc2275b0_1, \1075 );
not \U$893 ( \1270 , RIc2275b0_1);
not \U$894 ( \1271 , \1075 );
and \U$895 ( \1272 , \1270 , \1271 );
nor \U$896 ( \1273 , \1269 , \1272 );
or \U$897 ( \1274 , \1273 , \899 );
nand \U$898 ( \1275 , \1268 , \1274 );
xor \U$899 ( \1276 , \1267 , \1275 );
xor \U$900 ( \1277 , \1091 , \1093 );
and \U$901 ( \1278 , \1277 , \1101 );
and \U$902 ( \1279 , \1091 , \1093 );
or \U$903 ( \1280 , \1278 , \1279 );
xor \U$904 ( \1281 , \901 , \958 );
and \U$905 ( \1282 , \1281 , \1088 );
and \U$906 ( \1283 , \901 , \958 );
or \U$907 ( \1284 , \1282 , \1283 );
xor \U$908 ( \1285 , \1280 , \1284 );
xor \U$909 ( \1286 , \1276 , \1285 );
nor \U$910 ( \1287 , \1259 , \1286 );
nor \U$911 ( \1288 , \1251 , \1287 );
not \U$912 ( \1289 , \1288 );
and \U$913 ( \1290 , \932 , RIc227100_11);
not \U$914 ( \1291 , RIc227100_11);
and \U$915 ( \1292 , \931 , \1291 );
nor \U$916 ( \1293 , \1290 , \1292 );
and \U$917 ( \1294 , RIc227088_12, RIc227010_13);
not \U$918 ( \1295 , RIc227088_12);
not \U$919 ( \1296 , RIc227010_13);
and \U$920 ( \1297 , \1295 , \1296 );
nor \U$921 ( \1298 , \1294 , \1297 );
not \U$922 ( \1299 , \1298 );
and \U$923 ( \1300 , RIc227088_12, RIc227100_11);
not \U$924 ( \1301 , RIc227088_12);
not \U$925 ( \1302 , RIc227100_11);
and \U$926 ( \1303 , \1301 , \1302 );
nor \U$927 ( \1304 , \1300 , \1303 );
nand \U$928 ( \1305 , \1299 , \1304 );
not \U$929 ( \1306 , \1305 );
buf \U$930 ( \1307 , \1306 );
not \U$931 ( \1308 , \1307 );
or \U$932 ( \1309 , \1293 , \1308 );
buf \U$933 ( \1310 , \1298 );
buf \U$934 ( \1311 , \1310 );
not \U$935 ( \1312 , \1311 );
or \U$936 ( \1313 , \1312 , \1302 );
nand \U$937 ( \1314 , \1309 , \1313 );
nand \U$938 ( \1315 , \431 , \419 );
nor \U$939 ( \1316 , \902 , \1315 );
not \U$940 ( \1317 , \1316 );
not \U$941 ( \1318 , \688 );
or \U$942 ( \1319 , \1317 , \1318 );
not \U$943 ( \1320 , \1315 );
and \U$944 ( \1321 , \763 , \1320 );
not \U$945 ( \1322 , \419 );
not \U$946 ( \1323 , \785 );
or \U$947 ( \1324 , \1322 , \1323 );
not \U$948 ( \1325 , \797 );
nand \U$949 ( \1326 , \1324 , \1325 );
nor \U$950 ( \1327 , \1321 , \1326 );
nand \U$951 ( \1328 , \1319 , \1327 );
nand \U$952 ( \1329 , \423 , \801 );
xnor \U$953 ( \1330 , \1328 , \1329 );
buf \U$954 ( \1331 , \1330 );
buf \U$955 ( \1332 , \1331 );
not \U$956 ( \1333 , \1332 );
buf \U$957 ( \1334 , \1333 );
not \U$958 ( \1335 , \1334 );
and \U$959 ( \1336 , \1335 , RIc2275b0_1);
xor \U$960 ( \1337 , \1314 , \1336 );
xor \U$961 ( \1338 , RIc227100_11, RIc227178_10);
buf \U$962 ( \1339 , \1338 );
buf \U$963 ( \1340 , \1339 );
not \U$964 ( \1341 , \1340 );
not \U$965 ( \1342 , RIc2271f0_9);
and \U$966 ( \1343 , \1342 , \1074 );
not \U$967 ( \1344 , \1342 );
and \U$968 ( \1345 , \1344 , \1073 );
nor \U$969 ( \1346 , \1343 , \1345 );
not \U$970 ( \1347 , \1346 );
or \U$971 ( \1348 , \1341 , \1347 );
not \U$972 ( \1349 , \889 );
and \U$973 ( \1350 , \1349 , RIc2271f0_9);
not \U$974 ( \1351 , RIc2271f0_9);
and \U$975 ( \1352 , \889 , \1351 );
nor \U$976 ( \1353 , \1350 , \1352 );
not \U$977 ( \1354 , RIc227178_10);
and \U$978 ( \1355 , RIc227100_11, \1354 );
not \U$979 ( \1356 , RIc227100_11);
and \U$980 ( \1357 , \1356 , RIc227178_10);
nor \U$981 ( \1358 , \1355 , \1357 );
and \U$982 ( \1359 , \1342 , \1354 );
and \U$983 ( \1360 , RIc2271f0_9, RIc227178_10);
nor \U$984 ( \1361 , \1359 , \1360 );
and \U$985 ( \1362 , \1358 , \1361 );
buf \U$986 ( \1363 , \1362 );
not \U$987 ( \1364 , \1363 );
or \U$988 ( \1365 , \1353 , \1364 );
nand \U$989 ( \1366 , \1348 , \1365 );
not \U$990 ( \1367 , \1082 );
and \U$991 ( \1368 , RIc2274c0_3, \1223 );
not \U$992 ( \1369 , RIc2274c0_3);
buf \U$993 ( \1370 , \1220 );
buf \U$994 ( \1371 , \1370 );
not \U$995 ( \1372 , \1371 );
and \U$996 ( \1373 , \1369 , \1372 );
nor \U$997 ( \1374 , \1368 , \1373 );
not \U$998 ( \1375 , \1374 );
or \U$999 ( \1376 , \1367 , \1375 );
nor \U$1000 ( \1377 , \902 , \433 );
not \U$1001 ( \1378 , \1377 );
not \U$1002 ( \1379 , \688 );
or \U$1003 ( \1380 , \1378 , \1379 );
not \U$1004 ( \1381 , \433 );
and \U$1005 ( \1382 , \763 , \1381 );
nor \U$1006 ( \1383 , \1382 , \808 );
nand \U$1007 ( \1384 , \1380 , \1383 );
nand \U$1008 ( \1385 , \1200 , \812 );
not \U$1009 ( \1386 , \1385 );
and \U$1010 ( \1387 , \1384 , \1386 );
not \U$1011 ( \1388 , \1384 );
and \U$1012 ( \1389 , \1388 , \1385 );
nor \U$1013 ( \1390 , \1387 , \1389 );
buf \U$1014 ( \1391 , \1390 );
not \U$1015 ( \1392 , \1391 );
buf \U$1016 ( \1393 , \1392 );
and \U$1017 ( \1394 , RIc2274c0_3, \1393 );
not \U$1018 ( \1395 , RIc2274c0_3);
not \U$1019 ( \1396 , \1393 );
and \U$1020 ( \1397 , \1395 , \1396 );
nor \U$1021 ( \1398 , \1394 , \1397 );
or \U$1022 ( \1399 , \1398 , \1041 );
nand \U$1023 ( \1400 , \1376 , \1399 );
xor \U$1024 ( \1401 , \1366 , \1400 );
not \U$1025 ( \1402 , \1169 );
not \U$1026 ( \1403 , \1402 );
not \U$1027 ( \1404 , \1403 );
and \U$1028 ( \1405 , \1404 , RIc2273d0_5);
and \U$1029 ( \1406 , \1228 , \946 );
nor \U$1030 ( \1407 , \1405 , \1406 );
or \U$1031 ( \1408 , \1407 , \952 );
and \U$1032 ( \1409 , \1022 , RIc2273d0_5);
and \U$1033 ( \1410 , \1127 , \946 );
nor \U$1034 ( \1411 , \1409 , \1410 );
or \U$1035 ( \1412 , \1411 , \955 );
nand \U$1036 ( \1413 , \1408 , \1412 );
and \U$1037 ( \1414 , \1401 , \1413 );
and \U$1038 ( \1415 , \1366 , \1400 );
or \U$1039 ( \1416 , \1414 , \1415 );
and \U$1040 ( \1417 , \1337 , \1416 );
and \U$1041 ( \1418 , \1314 , \1336 );
or \U$1042 ( \1419 , \1417 , \1418 );
not \U$1043 ( \1420 , \1118 );
and \U$1044 ( \1421 , \892 , RIc2272e0_7);
not \U$1045 ( \1422 , \892 );
not \U$1046 ( \1423 , RIc2272e0_7);
and \U$1047 ( \1424 , \1422 , \1423 );
nor \U$1048 ( \1425 , \1421 , \1424 );
not \U$1049 ( \1426 , \1425 );
or \U$1050 ( \1427 , \1420 , \1426 );
and \U$1051 ( \1428 , \1075 , RIc2272e0_7);
and \U$1052 ( \1429 , \1073 , \1139 );
nor \U$1053 ( \1430 , \1428 , \1429 );
not \U$1054 ( \1431 , \1121 );
or \U$1055 ( \1432 , \1430 , \1431 );
nand \U$1056 ( \1433 , \1427 , \1432 );
not \U$1057 ( \1434 , \854 );
xor \U$1058 ( \1435 , RIc2275b0_1, \1396 );
not \U$1059 ( \1436 , \1435 );
or \U$1060 ( \1437 , \1434 , \1436 );
not \U$1061 ( \1438 , \1370 );
not \U$1062 ( \1439 , \1438 );
not \U$1063 ( \1440 , \1439 );
buf \U$1064 ( \1441 , \1440 );
buf \U$1065 ( \1442 , \1441 );
and \U$1066 ( \1443 , RIc2275b0_1, \1442 );
not \U$1067 ( \1444 , RIc2275b0_1);
and \U$1068 ( \1445 , \1444 , \1223 );
nor \U$1069 ( \1446 , \1443 , \1445 );
or \U$1070 ( \1447 , \1446 , \899 );
nand \U$1071 ( \1448 , \1437 , \1447 );
xor \U$1072 ( \1449 , \1433 , \1448 );
and \U$1073 ( \1450 , \1404 , RIc2274c0_3);
and \U$1074 ( \1451 , \1403 , \1032 );
nor \U$1075 ( \1452 , \1450 , \1451 );
or \U$1076 ( \1453 , \1452 , \1041 );
buf \U$1077 ( \1454 , \1020 );
buf \U$1078 ( \1455 , \1454 );
not \U$1079 ( \1456 , \1455 );
and \U$1080 ( \1457 , \1456 , RIc2274c0_3);
and \U$1081 ( \1458 , \1127 , \1027 );
nor \U$1082 ( \1459 , \1457 , \1458 );
or \U$1083 ( \1460 , \1459 , \1083 );
nand \U$1084 ( \1461 , \1453 , \1460 );
xor \U$1085 ( \1462 , \1449 , \1461 );
xor \U$1086 ( \1463 , \1419 , \1462 );
not \U$1087 ( \1464 , RIc2275b0_1);
not \U$1088 ( \1465 , \431 );
nor \U$1089 ( \1466 , \1465 , \418 );
and \U$1090 ( \1467 , \416 , \1466 );
not \U$1091 ( \1468 , \1467 );
not \U$1092 ( \1469 , \688 );
or \U$1093 ( \1470 , \1468 , \1469 );
and \U$1094 ( \1471 , \763 , \1466 );
not \U$1095 ( \1472 , \418 );
not \U$1096 ( \1473 , \1472 );
not \U$1097 ( \1474 , \785 );
or \U$1098 ( \1475 , \1473 , \1474 );
nand \U$1099 ( \1476 , \1475 , \790 );
nor \U$1100 ( \1477 , \1471 , \1476 );
nand \U$1101 ( \1478 , \1470 , \1477 );
nand \U$1102 ( \1479 , \793 , \796 );
not \U$1103 ( \1480 , \1479 );
and \U$1104 ( \1481 , \1478 , \1480 );
not \U$1105 ( \1482 , \1478 );
and \U$1106 ( \1483 , \1482 , \1479 );
nor \U$1107 ( \1484 , \1481 , \1483 );
buf \U$1108 ( \1485 , \1484 );
buf \U$1109 ( \1486 , \1485 );
not \U$1110 ( \1487 , \1486 );
buf \U$1111 ( \1488 , \1487 );
nor \U$1112 ( \1489 , \1464 , \1488 );
buf \U$1113 ( \1490 , \983 );
and \U$1114 ( \1491 , \1490 , RIc2272e0_7);
and \U$1115 ( \1492 , \985 , \1139 );
nor \U$1116 ( \1493 , \1491 , \1492 );
or \U$1117 ( \1494 , \1493 , \1117 );
and \U$1118 ( \1495 , \842 , RIc2272e0_7);
and \U$1119 ( \1496 , \841 , \1423 );
nor \U$1120 ( \1497 , \1495 , \1496 );
or \U$1121 ( \1498 , \1497 , \1431 );
nand \U$1122 ( \1499 , \1494 , \1498 );
xor \U$1123 ( \1500 , \1489 , \1499 );
and \U$1124 ( \1501 , RIc2275b0_1, \1334 );
not \U$1125 ( \1502 , RIc2275b0_1);
and \U$1126 ( \1503 , \1502 , \1335 );
nor \U$1127 ( \1504 , \1501 , \1503 );
or \U$1128 ( \1505 , \1504 , \855 );
nand \U$1129 ( \1506 , \423 , \419 );
nor \U$1130 ( \1507 , \1506 , \1465 );
and \U$1131 ( \1508 , \416 , \1507 );
not \U$1132 ( \1509 , \1508 );
not \U$1133 ( \1510 , \688 );
or \U$1134 ( \1511 , \1509 , \1510 );
and \U$1135 ( \1512 , \763 , \1507 );
not \U$1136 ( \1513 , \1506 );
not \U$1137 ( \1514 , \1513 );
not \U$1138 ( \1515 , \785 );
or \U$1139 ( \1516 , \1514 , \1515 );
and \U$1140 ( \1517 , \797 , \423 );
not \U$1141 ( \1518 , \801 );
nor \U$1142 ( \1519 , \1517 , \1518 );
nand \U$1143 ( \1520 , \1516 , \1519 );
nor \U$1144 ( \1521 , \1512 , \1520 );
nand \U$1145 ( \1522 , \1511 , \1521 );
nor \U$1146 ( \1523 , \804 , \421 );
and \U$1147 ( \1524 , \1522 , \1523 );
not \U$1148 ( \1525 , \1522 );
not \U$1149 ( \1526 , \1523 );
and \U$1150 ( \1527 , \1525 , \1526 );
nor \U$1151 ( \1528 , \1524 , \1527 );
buf \U$1152 ( \1529 , \1528 );
not \U$1153 ( \1530 , \1529 );
buf \U$1154 ( \1531 , \1530 );
not \U$1155 ( \1532 , \1531 );
buf \U$1156 ( \1533 , \1532 );
not \U$1157 ( \1534 , \1533 );
and \U$1158 ( \1535 , RIc2275b0_1, \1534 );
not \U$1159 ( \1536 , RIc2275b0_1);
and \U$1160 ( \1537 , \1536 , \1533 );
nor \U$1161 ( \1538 , \1535 , \1537 );
or \U$1162 ( \1539 , \1538 , \899 );
nand \U$1163 ( \1540 , \1505 , \1539 );
and \U$1164 ( \1541 , \1500 , \1540 );
and \U$1165 ( \1542 , \1489 , \1499 );
or \U$1166 ( \1543 , \1541 , \1542 );
or \U$1167 ( \1544 , \1307 , \1311 );
nand \U$1168 ( \1545 , \1544 , RIc227100_11);
not \U$1169 ( \1546 , \1363 );
not \U$1170 ( \1547 , \1346 );
or \U$1171 ( \1548 , \1546 , \1547 );
and \U$1172 ( \1549 , \932 , RIc2271f0_9);
and \U$1173 ( \1550 , \931 , \1342 );
nor \U$1174 ( \1551 , \1549 , \1550 );
not \U$1175 ( \1552 , \1340 );
or \U$1176 ( \1553 , \1551 , \1552 );
nand \U$1177 ( \1554 , \1548 , \1553 );
xor \U$1178 ( \1555 , \1545 , \1554 );
or \U$1179 ( \1556 , \1411 , \952 );
not \U$1180 ( \1557 , \980 );
buf \U$1181 ( \1558 , \1557 );
buf \U$1182 ( \1559 , \1558 );
and \U$1183 ( \1560 , \1559 , RIc2273d0_5);
not \U$1184 ( \1561 , \1490 );
and \U$1185 ( \1562 , \1561 , \946 );
nor \U$1186 ( \1563 , \1560 , \1562 );
or \U$1187 ( \1564 , \1563 , \955 );
nand \U$1188 ( \1565 , \1556 , \1564 );
xor \U$1189 ( \1566 , \1555 , \1565 );
xor \U$1190 ( \1567 , \1543 , \1566 );
not \U$1191 ( \1568 , \1040 );
not \U$1192 ( \1569 , \1374 );
or \U$1193 ( \1570 , \1568 , \1569 );
or \U$1194 ( \1571 , \1452 , \1083 );
nand \U$1195 ( \1572 , \1570 , \1571 );
not \U$1196 ( \1573 , \1121 );
not \U$1197 ( \1574 , \1425 );
or \U$1198 ( \1575 , \1573 , \1574 );
or \U$1199 ( \1576 , \1497 , \1117 );
nand \U$1200 ( \1577 , \1575 , \1576 );
xor \U$1201 ( \1578 , \1572 , \1577 );
not \U$1202 ( \1579 , \899 );
not \U$1203 ( \1580 , \1579 );
not \U$1204 ( \1581 , \1435 );
or \U$1205 ( \1582 , \1580 , \1581 );
or \U$1206 ( \1583 , \1538 , \855 );
nand \U$1207 ( \1584 , \1582 , \1583 );
xor \U$1208 ( \1585 , \1578 , \1584 );
and \U$1209 ( \1586 , \1567 , \1585 );
and \U$1210 ( \1587 , \1543 , \1566 );
or \U$1211 ( \1588 , \1586 , \1587 );
and \U$1212 ( \1589 , \1463 , \1588 );
and \U$1213 ( \1590 , \1419 , \1462 );
or \U$1214 ( \1591 , \1589 , \1590 );
xor \U$1215 ( \1592 , \1545 , \1554 );
and \U$1216 ( \1593 , \1592 , \1565 );
and \U$1217 ( \1594 , \1545 , \1554 );
or \U$1218 ( \1595 , \1593 , \1594 );
not \U$1219 ( \1596 , \1551 );
not \U$1220 ( \1597 , \1364 );
and \U$1221 ( \1598 , \1596 , \1597 );
and \U$1222 ( \1599 , \1340 , RIc2271f0_9);
nor \U$1223 ( \1600 , \1598 , \1599 );
not \U$1224 ( \1601 , RIc2275b0_1);
not \U$1225 ( \1602 , \1533 );
nor \U$1226 ( \1603 , \1601 , \1602 );
xor \U$1227 ( \1604 , \1600 , \1603 );
not \U$1228 ( \1605 , \954 );
and \U$1229 ( \1606 , \841 , RIc2273d0_5);
not \U$1230 ( \1607 , \841 );
and \U$1231 ( \1608 , \1607 , \946 );
nor \U$1232 ( \1609 , \1606 , \1608 );
not \U$1233 ( \1610 , \1609 );
or \U$1234 ( \1611 , \1605 , \1610 );
or \U$1235 ( \1612 , \1563 , \952 );
nand \U$1236 ( \1613 , \1611 , \1612 );
xor \U$1237 ( \1614 , \1604 , \1613 );
xor \U$1238 ( \1615 , \1595 , \1614 );
xor \U$1239 ( \1616 , \1572 , \1577 );
and \U$1240 ( \1617 , \1616 , \1584 );
and \U$1241 ( \1618 , \1572 , \1577 );
or \U$1242 ( \1619 , \1617 , \1618 );
and \U$1243 ( \1620 , \1615 , \1619 );
and \U$1244 ( \1621 , \1595 , \1614 );
or \U$1245 ( \1622 , \1620 , \1621 );
xor \U$1246 ( \1623 , \1591 , \1622 );
or \U$1247 ( \1624 , \1459 , \1041 );
and \U$1248 ( \1625 , \986 , RIc2274c0_3);
and \U$1249 ( \1626 , \1561 , \1032 );
nor \U$1250 ( \1627 , \1625 , \1626 );
or \U$1251 ( \1628 , \1627 , \1083 );
nand \U$1252 ( \1629 , \1624 , \1628 );
or \U$1253 ( \1630 , \1597 , \1340 );
nand \U$1254 ( \1631 , \1630 , RIc2271f0_9);
xor \U$1255 ( \1632 , \1629 , \1631 );
not \U$1256 ( \1633 , \1118 );
not \U$1257 ( \1634 , \1430 );
not \U$1258 ( \1635 , \1634 );
or \U$1259 ( \1636 , \1633 , \1635 );
or \U$1260 ( \1637 , \1141 , \1431 );
nand \U$1261 ( \1638 , \1636 , \1637 );
xor \U$1262 ( \1639 , \1632 , \1638 );
xor \U$1263 ( \1640 , \1600 , \1603 );
and \U$1264 ( \1641 , \1640 , \1613 );
and \U$1265 ( \1642 , \1600 , \1603 );
or \U$1266 ( \1643 , \1641 , \1642 );
xor \U$1267 ( \1644 , \1433 , \1448 );
and \U$1268 ( \1645 , \1644 , \1461 );
and \U$1269 ( \1646 , \1433 , \1448 );
or \U$1270 ( \1647 , \1645 , \1646 );
not \U$1271 ( \1648 , \1600 );
xor \U$1272 ( \1649 , \1647 , \1648 );
and \U$1273 ( \1650 , RIc2275b0_1, \1396 );
not \U$1274 ( \1651 , \951 );
not \U$1275 ( \1652 , \1609 );
or \U$1276 ( \1653 , \1651 , \1652 );
or \U$1277 ( \1654 , \1196 , \955 );
nand \U$1278 ( \1655 , \1653 , \1654 );
xor \U$1279 ( \1656 , \1650 , \1655 );
or \U$1280 ( \1657 , \1446 , \855 );
or \U$1281 ( \1658 , \1230 , \899 );
nand \U$1282 ( \1659 , \1657 , \1658 );
xor \U$1283 ( \1660 , \1656 , \1659 );
xor \U$1284 ( \1661 , \1649 , \1660 );
xor \U$1285 ( \1662 , \1643 , \1661 );
xor \U$1286 ( \1663 , \1639 , \1662 );
xor \U$1287 ( \1664 , \1623 , \1663 );
xor \U$1288 ( \1665 , \1595 , \1614 );
xor \U$1289 ( \1666 , \1665 , \1619 );
xor \U$1290 ( \1667 , \1419 , \1462 );
xor \U$1291 ( \1668 , \1667 , \1588 );
and \U$1292 ( \1669 , \1666 , \1668 );
and \U$1293 ( \1670 , RIc227010_13, RIc226f98_14);
nor \U$1294 ( \1671 , RIc227010_13, RIc226f98_14);
and \U$1295 ( \1672 , RIc226f98_14, RIc226f20_15);
not \U$1296 ( \1673 , RIc226f98_14);
not \U$1297 ( \1674 , RIc226f20_15);
and \U$1298 ( \1675 , \1673 , \1674 );
nor \U$1299 ( \1676 , \1672 , \1675 );
nor \U$1300 ( \1677 , \1670 , \1671 , \1676 );
buf \U$1301 ( \1678 , \1677 );
not \U$1302 ( \1679 , \1678 );
not \U$1303 ( \1680 , \1679 );
buf \U$1304 ( \1681 , \1676 );
buf \U$1305 ( \1682 , \1681 );
or \U$1306 ( \1683 , \1680 , \1682 );
nand \U$1307 ( \1684 , \1683 , RIc227010_13);
not \U$1308 ( \1685 , RIc227100_11);
and \U$1309 ( \1686 , \1685 , \1073 );
not \U$1310 ( \1687 , \1685 );
and \U$1311 ( \1688 , \1687 , \1075 );
nor \U$1312 ( \1689 , \1686 , \1688 );
or \U$1313 ( \1690 , \1689 , \1308 );
or \U$1314 ( \1691 , \1293 , \1312 );
nand \U$1315 ( \1692 , \1690 , \1691 );
xor \U$1316 ( \1693 , \1684 , \1692 );
and \U$1317 ( \1694 , \1456 , RIc2272e0_7);
and \U$1318 ( \1695 , \1455 , \1139 );
nor \U$1319 ( \1696 , \1694 , \1695 );
or \U$1320 ( \1697 , \1696 , \1117 );
or \U$1321 ( \1698 , \1493 , \1431 );
nand \U$1322 ( \1699 , \1697 , \1698 );
and \U$1323 ( \1700 , \1693 , \1699 );
and \U$1324 ( \1701 , \1684 , \1692 );
or \U$1325 ( \1702 , \1700 , \1701 );
not \U$1326 ( \1703 , \1314 );
xor \U$1327 ( \1704 , \1702 , \1703 );
not \U$1328 ( \1705 , \1597 );
not \U$1329 ( \1706 , \840 );
and \U$1330 ( \1707 , \1706 , \1351 );
not \U$1331 ( \1708 , \1706 );
and \U$1332 ( \1709 , \1708 , RIc2271f0_9);
nor \U$1333 ( \1710 , \1707 , \1709 );
not \U$1334 ( \1711 , \1710 );
or \U$1335 ( \1712 , \1705 , \1711 );
or \U$1336 ( \1713 , \1353 , \1552 );
nand \U$1337 ( \1714 , \1712 , \1713 );
nor \U$1338 ( \1715 , \902 , \1465 );
not \U$1339 ( \1716 , \1715 );
not \U$1340 ( \1717 , \688 );
or \U$1341 ( \1718 , \1716 , \1717 );
not \U$1342 ( \1719 , \1465 );
and \U$1343 ( \1720 , \763 , \1719 );
nor \U$1344 ( \1721 , \1720 , \785 );
nand \U$1345 ( \1722 , \1718 , \1721 );
nand \U$1346 ( \1723 , \1472 , \790 );
not \U$1347 ( \1724 , \1723 );
and \U$1348 ( \1725 , \1722 , \1724 );
not \U$1349 ( \1726 , \1722 );
and \U$1350 ( \1727 , \1726 , \1723 );
nor \U$1351 ( \1728 , \1725 , \1727 );
buf \U$1352 ( \1729 , \1728 );
buf \U$1353 ( \1730 , \1729 );
and \U$1354 ( \1731 , \1730 , RIc2275b0_1);
xor \U$1355 ( \1732 , \1714 , \1731 );
not \U$1356 ( \1733 , \951 );
not \U$1357 ( \1734 , \1442 );
or \U$1358 ( \1735 , \1734 , \946 );
or \U$1359 ( \1736 , \1372 , RIc2273d0_5);
nand \U$1360 ( \1737 , \1735 , \1736 );
not \U$1361 ( \1738 , \1737 );
or \U$1362 ( \1739 , \1733 , \1738 );
or \U$1363 ( \1740 , \1407 , \955 );
nand \U$1364 ( \1741 , \1739 , \1740 );
and \U$1365 ( \1742 , \1732 , \1741 );
and \U$1366 ( \1743 , \1714 , \1731 );
or \U$1367 ( \1744 , \1742 , \1743 );
and \U$1368 ( \1745 , \1704 , \1744 );
and \U$1369 ( \1746 , \1702 , \1703 );
or \U$1370 ( \1747 , \1745 , \1746 );
xor \U$1371 ( \1748 , \1314 , \1336 );
xor \U$1372 ( \1749 , \1748 , \1416 );
xor \U$1373 ( \1750 , \1747 , \1749 );
xor \U$1374 ( \1751 , \1489 , \1499 );
xor \U$1375 ( \1752 , \1751 , \1540 );
and \U$1376 ( \1753 , \932 , RIc227010_13);
and \U$1377 ( \1754 , \931 , \1296 );
nor \U$1378 ( \1755 , \1753 , \1754 );
or \U$1379 ( \1756 , \1755 , \1679 );
not \U$1380 ( \1757 , \1682 );
not \U$1381 ( \1758 , RIc227010_13);
or \U$1382 ( \1759 , \1757 , \1758 );
nand \U$1383 ( \1760 , \1756 , \1759 );
and \U$1384 ( \1761 , \1534 , RIc2274c0_3);
and \U$1385 ( \1762 , \1533 , \1032 );
nor \U$1386 ( \1763 , \1761 , \1762 );
or \U$1387 ( \1764 , \1763 , \1041 );
or \U$1388 ( \1765 , \1398 , \1083 );
nand \U$1389 ( \1766 , \1764 , \1765 );
xor \U$1390 ( \1767 , \1760 , \1766 );
and \U$1391 ( \1768 , RIc2275b0_1, \1488 );
not \U$1392 ( \1769 , RIc2275b0_1);
not \U$1393 ( \1770 , \1488 );
and \U$1394 ( \1771 , \1769 , \1770 );
nor \U$1395 ( \1772 , \1768 , \1771 );
or \U$1396 ( \1773 , \1772 , \855 );
or \U$1397 ( \1774 , \1504 , \899 );
nand \U$1398 ( \1775 , \1773 , \1774 );
and \U$1399 ( \1776 , \1767 , \1775 );
and \U$1400 ( \1777 , \1760 , \1766 );
or \U$1401 ( \1778 , \1776 , \1777 );
xor \U$1402 ( \1779 , \1752 , \1778 );
xor \U$1403 ( \1780 , \1366 , \1400 );
xor \U$1404 ( \1781 , \1780 , \1413 );
and \U$1405 ( \1782 , \1779 , \1781 );
and \U$1406 ( \1783 , \1752 , \1778 );
or \U$1407 ( \1784 , \1782 , \1783 );
and \U$1408 ( \1785 , \1750 , \1784 );
and \U$1409 ( \1786 , \1747 , \1749 );
or \U$1410 ( \1787 , \1785 , \1786 );
xor \U$1411 ( \1788 , \1419 , \1462 );
xor \U$1412 ( \1789 , \1788 , \1588 );
and \U$1413 ( \1790 , \1787 , \1789 );
and \U$1414 ( \1791 , \1666 , \1787 );
or \U$1415 ( \1792 , \1669 , \1790 , \1791 );
nor \U$1416 ( \1793 , \1664 , \1792 );
xor \U$1417 ( \1794 , \1199 , \1224 );
xor \U$1418 ( \1795 , \1794 , \1233 );
xor \U$1419 ( \1796 , \1629 , \1631 );
and \U$1420 ( \1797 , \1796 , \1638 );
and \U$1421 ( \1798 , \1629 , \1631 );
or \U$1422 ( \1799 , \1797 , \1798 );
xor \U$1423 ( \1800 , \1795 , \1799 );
or \U$1424 ( \1801 , \1627 , \1041 );
or \U$1425 ( \1802 , \1177 , \1083 );
nand \U$1426 ( \1803 , \1801 , \1802 );
xor \U$1427 ( \1804 , \1803 , \1145 );
xor \U$1428 ( \1805 , \1650 , \1655 );
and \U$1429 ( \1806 , \1805 , \1659 );
and \U$1430 ( \1807 , \1650 , \1655 );
or \U$1431 ( \1808 , \1806 , \1807 );
xor \U$1432 ( \1809 , \1804 , \1808 );
xor \U$1433 ( \1810 , \1800 , \1809 );
xor \U$1434 ( \1811 , \1647 , \1648 );
and \U$1435 ( \1812 , \1811 , \1660 );
and \U$1436 ( \1813 , \1647 , \1648 );
or \U$1437 ( \1814 , \1812 , \1813 );
xor \U$1438 ( \1815 , \1629 , \1631 );
xor \U$1439 ( \1816 , \1815 , \1638 );
and \U$1440 ( \1817 , \1643 , \1816 );
xor \U$1441 ( \1818 , \1629 , \1631 );
xor \U$1442 ( \1819 , \1818 , \1638 );
and \U$1443 ( \1820 , \1661 , \1819 );
and \U$1444 ( \1821 , \1643 , \1661 );
or \U$1445 ( \1822 , \1817 , \1820 , \1821 );
xor \U$1446 ( \1823 , \1814 , \1822 );
xor \U$1447 ( \1824 , \1810 , \1823 );
xor \U$1448 ( \1825 , \1591 , \1622 );
and \U$1449 ( \1826 , \1825 , \1663 );
and \U$1450 ( \1827 , \1591 , \1622 );
or \U$1451 ( \1828 , \1826 , \1827 );
nor \U$1452 ( \1829 , \1824 , \1828 );
nor \U$1453 ( \1830 , \1793 , \1829 );
not \U$1454 ( \1831 , \1830 );
xor \U$1455 ( \1832 , \1236 , \1238 );
xor \U$1456 ( \1833 , \1832 , \1241 );
xor \U$1457 ( \1834 , \1803 , \1145 );
and \U$1458 ( \1835 , \1834 , \1808 );
and \U$1459 ( \1836 , \1803 , \1145 );
or \U$1460 ( \1837 , \1835 , \1836 );
xor \U$1461 ( \1838 , \1795 , \1799 );
and \U$1462 ( \1839 , \1838 , \1809 );
and \U$1463 ( \1840 , \1795 , \1799 );
or \U$1464 ( \1841 , \1839 , \1840 );
xor \U$1465 ( \1842 , \1837 , \1841 );
xor \U$1466 ( \1843 , \1833 , \1842 );
xor \U$1467 ( \1844 , \1795 , \1799 );
xor \U$1468 ( \1845 , \1844 , \1809 );
and \U$1469 ( \1846 , \1814 , \1845 );
xor \U$1470 ( \1847 , \1795 , \1799 );
xor \U$1471 ( \1848 , \1847 , \1809 );
and \U$1472 ( \1849 , \1822 , \1848 );
and \U$1473 ( \1850 , \1814 , \1822 );
or \U$1474 ( \1851 , \1846 , \1849 , \1850 );
nor \U$1475 ( \1852 , \1843 , \1851 );
nor \U$1476 ( \1853 , \1831 , \1852 );
xor \U$1477 ( \1854 , \1236 , \1238 );
xor \U$1478 ( \1855 , \1854 , \1241 );
and \U$1479 ( \1856 , \1837 , \1855 );
xor \U$1480 ( \1857 , \1236 , \1238 );
xor \U$1481 ( \1858 , \1857 , \1241 );
and \U$1482 ( \1859 , \1841 , \1858 );
and \U$1483 ( \1860 , \1837 , \1841 );
or \U$1484 ( \1861 , \1856 , \1859 , \1860 );
xor \U$1485 ( \1862 , \1135 , \1136 );
xor \U$1486 ( \1863 , \1862 , \1183 );
xor \U$1487 ( \1864 , \1190 , \1244 );
xor \U$1488 ( \1865 , \1863 , \1864 );
or \U$1489 ( \1866 , \1861 , \1865 );
nand \U$1490 ( \1867 , \1853 , \1866 );
xor \U$1491 ( \1868 , \1264 , \1266 );
xor \U$1492 ( \1869 , \1868 , \1275 );
and \U$1493 ( \1870 , \1280 , \1869 );
xor \U$1494 ( \1871 , \1264 , \1266 );
xor \U$1495 ( \1872 , \1871 , \1275 );
and \U$1496 ( \1873 , \1284 , \1872 );
and \U$1497 ( \1874 , \1280 , \1284 );
or \U$1498 ( \1875 , \1870 , \1873 , \1874 );
or \U$1499 ( \1876 , \1273 , \855 );
xor \U$1500 ( \1877 , \932 , RIc2275b0_1);
or \U$1501 ( \1878 , \1877 , \899 );
nand \U$1502 ( \1879 , \1876 , \1878 );
not \U$1503 ( \1880 , \1879 );
not \U$1504 ( \1881 , \893 );
nand \U$1505 ( \1882 , \1881 , RIc2275b0_1);
and \U$1506 ( \1883 , \1041 , \1083 );
nor \U$1507 ( \1884 , \1883 , \1027 );
nand \U$1508 ( \1885 , \1882 , \1884 );
not \U$1509 ( \1886 , \1885 );
nor \U$1510 ( \1887 , \1882 , \1884 );
nor \U$1511 ( \1888 , \1886 , \1887 );
not \U$1512 ( \1889 , \1888 );
and \U$1513 ( \1890 , \1880 , \1889 );
and \U$1514 ( \1891 , \1879 , \1888 );
nor \U$1515 ( \1892 , \1890 , \1891 );
not \U$1516 ( \1893 , \1264 );
xor \U$1517 ( \1894 , \1892 , \1893 );
xor \U$1518 ( \1895 , \1264 , \1266 );
and \U$1519 ( \1896 , \1895 , \1275 );
and \U$1520 ( \1897 , \1264 , \1266 );
or \U$1521 ( \1898 , \1896 , \1897 );
xor \U$1522 ( \1899 , \1894 , \1898 );
nor \U$1523 ( \1900 , \1875 , \1899 );
nor \U$1524 ( \1901 , \1289 , \1867 , \1900 );
not \U$1525 ( \1902 , \1901 );
and \U$1526 ( \1903 , RIc226ae8_24, RIc226a70_25);
not \U$1527 ( \1904 , RIc226ae8_24);
not \U$1528 ( \1905 , RIc226a70_25);
and \U$1529 ( \1906 , \1904 , \1905 );
nor \U$1530 ( \1907 , \1903 , \1906 );
not \U$1531 ( \1908 , \1907 );
and \U$1532 ( \1909 , RIc226ae8_24, RIc226b60_23);
not \U$1533 ( \1910 , RIc226ae8_24);
not \U$1534 ( \1911 , RIc226b60_23);
and \U$1535 ( \1912 , \1910 , \1911 );
nor \U$1536 ( \1913 , \1909 , \1912 );
and \U$1537 ( \1914 , \1908 , \1913 );
buf \U$1538 ( \1915 , \1914 );
not \U$1539 ( \1916 , \1915 );
and \U$1540 ( \1917 , \1490 , RIc226b60_23);
not \U$1541 ( \1918 , \1490 );
not \U$1542 ( \1919 , RIc226b60_23);
and \U$1543 ( \1920 , \1918 , \1919 );
or \U$1544 ( \1921 , \1917 , \1920 );
not \U$1545 ( \1922 , \1921 );
or \U$1546 ( \1923 , \1916 , \1922 );
not \U$1547 ( \1924 , RIc226b60_23);
not \U$1548 ( \1925 , \1706 );
or \U$1549 ( \1926 , \1924 , \1925 );
not \U$1550 ( \1927 , RIc226b60_23);
nand \U$1551 ( \1928 , \841 , \1927 );
nand \U$1552 ( \1929 , \1926 , \1928 );
buf \U$1553 ( \1930 , \1907 );
nand \U$1554 ( \1931 , \1929 , \1930 );
nand \U$1555 ( \1932 , \1923 , \1931 );
and \U$1556 ( \1933 , RIc226db8_18, RIc226e30_17);
not \U$1557 ( \1934 , RIc226db8_18);
not \U$1558 ( \1935 , RIc226e30_17);
and \U$1559 ( \1936 , \1934 , \1935 );
nor \U$1560 ( \1937 , \1933 , \1936 );
not \U$1561 ( \1938 , \1937 );
and \U$1562 ( \1939 , RIc226db8_18, RIc226d40_19);
not \U$1563 ( \1940 , RIc226db8_18);
not \U$1564 ( \1941 , RIc226d40_19);
and \U$1565 ( \1942 , \1940 , \1941 );
nor \U$1566 ( \1943 , \1939 , \1942 );
nor \U$1567 ( \1944 , \1938 , \1943 );
buf \U$1568 ( \1945 , \1944 );
not \U$1569 ( \1946 , \1945 );
not \U$1570 ( \1947 , RIc226e30_17);
not \U$1571 ( \1948 , \1331 );
buf \U$1572 ( \1949 , \1948 );
not \U$1573 ( \1950 , \1949 );
or \U$1574 ( \1951 , \1947 , \1950 );
not \U$1575 ( \1952 , RIc226e30_17);
nand \U$1576 ( \1953 , \1335 , \1952 );
nand \U$1577 ( \1954 , \1951 , \1953 );
not \U$1578 ( \1955 , \1954 );
or \U$1579 ( \1956 , \1946 , \1955 );
not \U$1580 ( \1957 , RIc226e30_17);
not \U$1581 ( \1958 , \1602 );
or \U$1582 ( \1959 , \1957 , \1958 );
not \U$1583 ( \1960 , RIc226e30_17);
nand \U$1584 ( \1961 , \1533 , \1960 );
nand \U$1585 ( \1962 , \1959 , \1961 );
buf \U$1586 ( \1963 , \1943 );
nand \U$1587 ( \1964 , \1962 , \1963 );
nand \U$1588 ( \1965 , \1956 , \1964 );
xor \U$1589 ( \1966 , \1932 , \1965 );
not \U$1590 ( \1967 , \1121 );
not \U$1591 ( \1968 , \381 );
nand \U$1592 ( \1969 , \395 , \1968 );
not \U$1593 ( \1970 , \414 );
nor \U$1594 ( \1971 , \1969 , \1970 );
not \U$1595 ( \1972 , \1971 );
not \U$1596 ( \1973 , \688 );
or \U$1597 ( \1974 , \1972 , \1973 );
buf \U$1598 ( \1975 , \721 );
not \U$1599 ( \1976 , \1969 );
and \U$1600 ( \1977 , \1975 , \1976 );
not \U$1601 ( \1978 , \1968 );
not \U$1602 ( \1979 , \740 );
or \U$1603 ( \1980 , \1978 , \1979 );
not \U$1604 ( \1981 , \744 );
nand \U$1605 ( \1982 , \1981 , RIc224ec8_84);
nand \U$1606 ( \1983 , \1980 , \1982 );
nor \U$1607 ( \1984 , \1977 , \1983 );
nand \U$1608 ( \1985 , \1974 , \1984 );
nand \U$1609 ( \1986 , \747 , \750 );
xnor \U$1610 ( \1987 , \1985 , \1986 );
buf \U$1611 ( \1988 , \1987 );
not \U$1612 ( \1989 , \1988 );
buf \U$1613 ( \1990 , \1989 );
not \U$1614 ( \1991 , \1990 );
and \U$1615 ( \1992 , \1991 , RIc2272e0_7);
not \U$1616 ( \1993 , \1991 );
and \U$1617 ( \1994 , \1993 , \1139 );
nor \U$1618 ( \1995 , \1992 , \1994 );
not \U$1619 ( \1996 , \1995 );
or \U$1620 ( \1997 , \1967 , \1996 );
not \U$1621 ( \1998 , RIc2272e0_7);
not \U$1622 ( \1999 , \395 );
nor \U$1623 ( \2000 , \1999 , \1970 );
not \U$1624 ( \2001 , \2000 );
not \U$1625 ( \2002 , \688 );
or \U$1626 ( \2003 , \2001 , \2002 );
and \U$1627 ( \2004 , \395 , \1975 );
nor \U$1628 ( \2005 , \2004 , \740 );
nand \U$1629 ( \2006 , \2003 , \2005 );
nand \U$1630 ( \2007 , \1968 , \1982 );
not \U$1631 ( \2008 , \2007 );
and \U$1632 ( \2009 , \2006 , \2008 );
not \U$1633 ( \2010 , \2006 );
and \U$1634 ( \2011 , \2010 , \2007 );
nor \U$1635 ( \2012 , \2009 , \2011 );
buf \U$1636 ( \2013 , \2012 );
buf \U$1637 ( \2014 , \2013 );
not \U$1638 ( \2015 , \2014 );
not \U$1639 ( \2016 , \2015 );
or \U$1640 ( \2017 , \1998 , \2016 );
not \U$1641 ( \2018 , \2015 );
nand \U$1642 ( \2019 , \2018 , \1423 );
nand \U$1643 ( \2020 , \2017 , \2019 );
nand \U$1644 ( \2021 , \2020 , \1118 );
nand \U$1645 ( \2022 , \1997 , \2021 );
xor \U$1646 ( \2023 , \1966 , \2022 );
not \U$1647 ( \2024 , \854 );
nor \U$1648 ( \2025 , \404 , \411 );
not \U$1649 ( \2026 , \2025 );
not \U$1650 ( \2027 , \688 );
or \U$1651 ( \2028 , \2026 , \2027 );
nand \U$1652 ( \2029 , \708 , \714 );
not \U$1653 ( \2030 , \2029 );
and \U$1654 ( \2031 , \2030 , \717 );
not \U$1655 ( \2032 , \691 );
nor \U$1656 ( \2033 , \2031 , \2032 );
nand \U$1657 ( \2034 , \2028 , \2033 );
not \U$1658 ( \2035 , \693 );
nor \U$1659 ( \2036 , \2035 , \410 );
and \U$1660 ( \2037 , \2034 , \2036 );
not \U$1661 ( \2038 , \2034 );
not \U$1662 ( \2039 , \2036 );
and \U$1663 ( \2040 , \2038 , \2039 );
nor \U$1664 ( \2041 , \2037 , \2040 );
buf \U$1665 ( \2042 , \2041 );
not \U$1666 ( \2043 , \2042 );
not \U$1667 ( \2044 , \2043 );
xor \U$1668 ( \2045 , RIc2275b0_1, \2044 );
not \U$1669 ( \2046 , \2045 );
or \U$1670 ( \2047 , \2024 , \2046 );
not \U$1671 ( \2048 , \404 );
buf \U$1672 ( \2049 , \412 );
and \U$1673 ( \2050 , \2048 , \2049 );
not \U$1674 ( \2051 , \2050 );
not \U$1675 ( \2052 , \688 );
or \U$1676 ( \2053 , \2051 , \2052 );
and \U$1677 ( \2054 , \2030 , \2049 );
nor \U$1678 ( \2055 , \2054 , \694 );
nand \U$1679 ( \2056 , \2053 , \2055 );
nand \U$1680 ( \2057 , \716 , \696 );
not \U$1681 ( \2058 , \2057 );
and \U$1682 ( \2059 , \2056 , \2058 );
not \U$1683 ( \2060 , \2056 );
and \U$1684 ( \2061 , \2060 , \2057 );
nor \U$1685 ( \2062 , \2059 , \2061 );
not \U$1686 ( \2063 , \2062 );
not \U$1687 ( \2064 , \2063 );
buf \U$1688 ( \2065 , \2064 );
xor \U$1689 ( \2066 , RIc2275b0_1, \2065 );
nand \U$1690 ( \2067 , \2066 , \1579 );
nand \U$1691 ( \2068 , \2047 , \2067 );
not \U$1692 ( \2069 , \2068 );
and \U$1693 ( \2070 , RIc226818_30, RIc2267a0_31);
not \U$1694 ( \2071 , RIc226818_30);
not \U$1695 ( \2072 , RIc2267a0_31);
and \U$1696 ( \2073 , \2071 , \2072 );
nor \U$1697 ( \2074 , \2070 , \2073 );
not \U$1698 ( \2075 , \2074 );
xor \U$1699 ( \2076 , RIc226890_29, RIc226818_30);
nand \U$1700 ( \2077 , \2075 , \2076 );
not \U$1701 ( \2078 , \2077 );
not \U$1702 ( \2079 , \2078 );
and \U$1703 ( \2080 , RIc226890_29, \932 );
not \U$1704 ( \2081 , RIc226890_29);
and \U$1705 ( \2082 , \2081 , \931 );
or \U$1706 ( \2083 , \2080 , \2082 );
not \U$1707 ( \2084 , \2083 );
or \U$1708 ( \2085 , \2079 , \2084 );
buf \U$1709 ( \2086 , \2074 );
nand \U$1710 ( \2087 , \2086 , RIc226890_29);
nand \U$1711 ( \2088 , \2085 , \2087 );
not \U$1712 ( \2089 , \2088 );
nand \U$1713 ( \2090 , \2069 , \2089 );
not \U$1714 ( \2091 , \2090 );
and \U$1715 ( \2092 , \403 , \711 );
not \U$1716 ( \2093 , \2092 );
not \U$1717 ( \2094 , \688 );
or \U$1718 ( \2095 , \2093 , \2094 );
nand \U$1719 ( \2096 , \707 , \703 );
and \U$1720 ( \2097 , \2096 , \711 );
not \U$1721 ( \2098 , \701 );
nor \U$1722 ( \2099 , \2097 , \2098 );
nand \U$1723 ( \2100 , \2095 , \2099 );
nand \U$1724 ( \2101 , \709 , \702 );
xnor \U$1725 ( \2102 , \2100 , \2101 );
buf \U$1726 ( \2103 , \2102 );
not \U$1727 ( \2104 , \2103 );
not \U$1728 ( \2105 , \2104 );
and \U$1729 ( \2106 , RIc2275b0_1, \2105 );
not \U$1730 ( \2107 , \1915 );
not \U$1731 ( \2108 , RIc226b60_23);
not \U$1732 ( \2109 , \1404 );
or \U$1733 ( \2110 , \2108 , \2109 );
not \U$1734 ( \2111 , RIc226b60_23);
nand \U$1735 ( \2112 , \1228 , \2111 );
nand \U$1736 ( \2113 , \2110 , \2112 );
not \U$1737 ( \2114 , \2113 );
or \U$1738 ( \2115 , \2107 , \2114 );
not \U$1739 ( \2116 , RIc226b60_23);
buf \U$1740 ( \2117 , \1019 );
not \U$1741 ( \2118 , \2117 );
not \U$1742 ( \2119 , \2118 );
not \U$1743 ( \2120 , \2119 );
not \U$1744 ( \2121 , \2120 );
or \U$1745 ( \2122 , \2116 , \2121 );
nand \U$1746 ( \2123 , \1455 , \1919 );
nand \U$1747 ( \2124 , \2122 , \2123 );
nand \U$1748 ( \2125 , \2124 , \1930 );
nand \U$1749 ( \2126 , \2115 , \2125 );
xor \U$1750 ( \2127 , \2106 , \2126 );
not \U$1751 ( \2128 , RIc226908_28);
and \U$1752 ( \2129 , RIc226890_29, \2128 );
not \U$1753 ( \2130 , RIc226890_29);
and \U$1754 ( \2131 , \2130 , RIc226908_28);
nor \U$1755 ( \2132 , \2129 , \2131 );
not \U$1756 ( \2133 , RIc226980_27);
and \U$1757 ( \2134 , \2133 , \2128 );
and \U$1758 ( \2135 , RIc226980_27, RIc226908_28);
nor \U$1759 ( \2136 , \2134 , \2135 );
and \U$1760 ( \2137 , \2132 , \2136 );
buf \U$1761 ( \2138 , \2137 );
not \U$1762 ( \2139 , \2138 );
not \U$1763 ( \2140 , RIc226980_27);
not \U$1764 ( \2141 , \890 );
or \U$1765 ( \2142 , \2140 , \2141 );
nand \U$1766 ( \2143 , \891 , \2133 );
nand \U$1767 ( \2144 , \2142 , \2143 );
not \U$1768 ( \2145 , \2144 );
or \U$1769 ( \2146 , \2139 , \2145 );
not \U$1770 ( \2147 , RIc226980_27);
not \U$1771 ( \2148 , \1074 );
or \U$1772 ( \2149 , \2147 , \2148 );
not \U$1773 ( \2150 , RIc226980_27);
nand \U$1774 ( \2151 , \1073 , \2150 );
nand \U$1775 ( \2152 , \2149 , \2151 );
not \U$1776 ( \2153 , \2132 );
buf \U$1777 ( \2154 , \2153 );
not \U$1778 ( \2155 , \2154 );
not \U$1779 ( \2156 , \2155 );
nand \U$1780 ( \2157 , \2152 , \2156 );
nand \U$1781 ( \2158 , \2146 , \2157 );
and \U$1782 ( \2159 , \2127 , \2158 );
and \U$1783 ( \2160 , \2106 , \2126 );
or \U$1784 ( \2161 , \2159 , \2160 );
not \U$1785 ( \2162 , \2161 );
or \U$1786 ( \2163 , \2091 , \2162 );
nand \U$1787 ( \2164 , \2068 , \2088 );
nand \U$1788 ( \2165 , \2163 , \2164 );
xor \U$1789 ( \2166 , \2023 , \2165 );
not \U$1790 ( \2167 , RIc2269f8_26);
and \U$1791 ( \2168 , RIc226980_27, \2167 );
not \U$1792 ( \2169 , RIc226980_27);
and \U$1793 ( \2170 , \2169 , RIc2269f8_26);
nor \U$1794 ( \2171 , \2168 , \2170 );
not \U$1795 ( \2172 , \2171 );
buf \U$1796 ( \2173 , \2172 );
not \U$1797 ( \2174 , \2173 );
not \U$1798 ( \2175 , RIc226a70_25);
not \U$1799 ( \2176 , \842 );
or \U$1800 ( \2177 , \2175 , \2176 );
not \U$1801 ( \2178 , \840 );
not \U$1802 ( \2179 , \2178 );
nand \U$1803 ( \2180 , \2179 , \1905 );
nand \U$1804 ( \2181 , \2177 , \2180 );
not \U$1805 ( \2182 , \2181 );
or \U$1806 ( \2183 , \2174 , \2182 );
not \U$1807 ( \2184 , RIc226a70_25);
not \U$1808 ( \2185 , \1490 );
or \U$1809 ( \2186 , \2184 , \2185 );
not \U$1810 ( \2187 , RIc226a70_25);
nand \U$1811 ( \2188 , \984 , \2187 );
nand \U$1812 ( \2189 , \2186 , \2188 );
not \U$1813 ( \2190 , RIc226a70_25);
and \U$1814 ( \2191 , \2190 , \2167 );
and \U$1815 ( \2192 , RIc226a70_25, RIc2269f8_26);
nor \U$1816 ( \2193 , \2191 , \2192 );
and \U$1817 ( \2194 , \2171 , \2193 );
buf \U$1818 ( \2195 , \2194 );
nand \U$1819 ( \2196 , \2189 , \2195 );
nand \U$1820 ( \2197 , \2183 , \2196 );
not \U$1821 ( \2198 , \1311 );
not \U$1822 ( \2199 , RIc227100_11);
not \U$1823 ( \2200 , \382 );
nor \U$1824 ( \2201 , \2200 , \383 );
nand \U$1825 ( \2202 , \2201 , \395 );
nor \U$1826 ( \2203 , \2202 , \1970 );
not \U$1827 ( \2204 , \2203 );
not \U$1828 ( \2205 , \688 );
or \U$1829 ( \2206 , \2204 , \2205 );
not \U$1830 ( \2207 , \2202 );
and \U$1831 ( \2208 , \1975 , \2207 );
not \U$1832 ( \2209 , \2201 );
not \U$1833 ( \2210 , \740 );
or \U$1834 ( \2211 , \2209 , \2210 );
not \U$1835 ( \2212 , \383 );
and \U$1836 ( \2213 , \751 , \2212 );
not \U$1837 ( \2214 , \754 );
nor \U$1838 ( \2215 , \2213 , \2214 );
nand \U$1839 ( \2216 , \2211 , \2215 );
nor \U$1840 ( \2217 , \2208 , \2216 );
nand \U$1841 ( \2218 , \2206 , \2217 );
nor \U$1842 ( \2219 , \758 , \384 );
and \U$1843 ( \2220 , \2218 , \2219 );
not \U$1844 ( \2221 , \2218 );
not \U$1845 ( \2222 , \2219 );
and \U$1846 ( \2223 , \2221 , \2222 );
nor \U$1847 ( \2224 , \2220 , \2223 );
buf \U$1848 ( \2225 , \2224 );
not \U$1849 ( \2226 , \2225 );
buf \U$1850 ( \2227 , \2226 );
buf \U$1851 ( \2228 , \2227 );
not \U$1852 ( \2229 , \2228 );
not \U$1853 ( \2230 , \2229 );
not \U$1854 ( \2231 , \2230 );
or \U$1855 ( \2232 , \2199 , \2231 );
not \U$1856 ( \2233 , \2225 );
buf \U$1857 ( \2234 , \2233 );
not \U$1858 ( \2235 , \2234 );
nand \U$1859 ( \2236 , \2235 , \1302 );
nand \U$1860 ( \2237 , \2232 , \2236 );
not \U$1861 ( \2238 , \2237 );
or \U$1862 ( \2239 , \2198 , \2238 );
not \U$1863 ( \2240 , RIc227100_11);
nand \U$1864 ( \2241 , \395 , \382 );
nor \U$1865 ( \2242 , \2241 , \1970 );
not \U$1866 ( \2243 , \2242 );
not \U$1867 ( \2244 , \687 );
or \U$1868 ( \2245 , \2243 , \2244 );
not \U$1869 ( \2246 , \2241 );
and \U$1870 ( \2247 , \1975 , \2246 );
not \U$1871 ( \2248 , \740 );
not \U$1872 ( \2249 , \382 );
or \U$1873 ( \2250 , \2248 , \2249 );
not \U$1874 ( \2251 , \751 );
nand \U$1875 ( \2252 , \2250 , \2251 );
nor \U$1876 ( \2253 , \2247 , \2252 );
nand \U$1877 ( \2254 , \2245 , \2253 );
nand \U$1878 ( \2255 , \2212 , \754 );
xnor \U$1879 ( \2256 , \2254 , \2255 );
not \U$1880 ( \2257 , \2256 );
buf \U$1881 ( \2258 , \2257 );
not \U$1882 ( \2259 , \2258 );
or \U$1883 ( \2260 , \2240 , \2259 );
not \U$1884 ( \2261 , \2258 );
nand \U$1885 ( \2262 , \2261 , \1685 );
nand \U$1886 ( \2263 , \2260 , \2262 );
nand \U$1887 ( \2264 , \2263 , \1307 );
nand \U$1888 ( \2265 , \2239 , \2264 );
xor \U$1889 ( \2266 , \2197 , \2265 );
not \U$1890 ( \2267 , \1363 );
and \U$1891 ( \2268 , \2015 , RIc2271f0_9);
not \U$1892 ( \2269 , \2015 );
and \U$1893 ( \2270 , \2269 , \1342 );
or \U$1894 ( \2271 , \2268 , \2270 );
not \U$1895 ( \2272 , \2271 );
or \U$1896 ( \2273 , \2267 , \2272 );
not \U$1897 ( \2274 , RIc2271f0_9);
not \U$1898 ( \2275 , \1990 );
or \U$1899 ( \2276 , \2274 , \2275 );
nand \U$1900 ( \2277 , \1991 , \1351 );
nand \U$1901 ( \2278 , \2276 , \2277 );
nand \U$1902 ( \2279 , \2278 , \1340 );
nand \U$1903 ( \2280 , \2273 , \2279 );
and \U$1904 ( \2281 , \2266 , \2280 );
and \U$1905 ( \2282 , \2197 , \2265 );
or \U$1906 ( \2283 , \2281 , \2282 );
and \U$1907 ( \2284 , \416 , \428 );
not \U$1908 ( \2285 , \2284 );
not \U$1909 ( \2286 , \688 );
or \U$1910 ( \2287 , \2285 , \2286 );
and \U$1911 ( \2288 , \763 , \428 );
nor \U$1912 ( \2289 , \2288 , \776 );
nand \U$1913 ( \2290 , \2287 , \2289 );
nand \U$1914 ( \2291 , \430 , \779 );
not \U$1915 ( \2292 , \2291 );
and \U$1916 ( \2293 , \2290 , \2292 );
not \U$1917 ( \2294 , \2290 );
and \U$1918 ( \2295 , \2294 , \2291 );
nor \U$1919 ( \2296 , \2293 , \2295 );
buf \U$1920 ( \2297 , \2296 );
not \U$1921 ( \2298 , \2297 );
not \U$1922 ( \2299 , \2298 );
not \U$1923 ( \2300 , \2299 );
not \U$1924 ( \2301 , RIc226f20_15);
not \U$1925 ( \2302 , \2301 );
and \U$1926 ( \2303 , \2300 , \2302 );
not \U$1927 ( \2304 , \2297 );
not \U$1928 ( \2305 , \2304 );
buf \U$1929 ( \2306 , \2305 );
and \U$1930 ( \2307 , \2306 , \2301 );
nor \U$1931 ( \2308 , \2303 , \2307 );
not \U$1932 ( \2309 , \2308 );
and \U$1933 ( \2310 , RIc226ea8_16, RIc226f20_15);
not \U$1934 ( \2311 , RIc226ea8_16);
and \U$1935 ( \2312 , \2311 , \2301 );
nor \U$1936 ( \2313 , \2310 , \2312 );
not \U$1937 ( \2314 , \2313 );
and \U$1938 ( \2315 , RIc226ea8_16, RIc226e30_17);
not \U$1939 ( \2316 , RIc226ea8_16);
and \U$1940 ( \2317 , \2316 , \1960 );
nor \U$1941 ( \2318 , \2315 , \2317 );
nor \U$1942 ( \2319 , \2314 , \2318 );
buf \U$1943 ( \2320 , \2319 );
not \U$1944 ( \2321 , \2320 );
not \U$1945 ( \2322 , \2321 );
and \U$1946 ( \2323 , \2309 , \2322 );
not \U$1947 ( \2324 , \2301 );
not \U$1948 ( \2325 , \428 );
nor \U$1949 ( \2326 , \2325 , \770 );
and \U$1950 ( \2327 , \416 , \2326 );
not \U$1951 ( \2328 , \2327 );
not \U$1952 ( \2329 , \688 );
or \U$1953 ( \2330 , \2328 , \2329 );
and \U$1954 ( \2331 , \763 , \2326 );
not \U$1955 ( \2332 , \430 );
not \U$1956 ( \2333 , \776 );
or \U$1957 ( \2334 , \2332 , \2333 );
nand \U$1958 ( \2335 , \2334 , \779 );
nor \U$1959 ( \2336 , \2331 , \2335 );
nand \U$1960 ( \2337 , \2330 , \2336 );
and \U$1961 ( \2338 , \429 , \782 );
and \U$1962 ( \2339 , \2337 , \2338 );
not \U$1963 ( \2340 , \2337 );
not \U$1964 ( \2341 , \2338 );
and \U$1965 ( \2342 , \2340 , \2341 );
nor \U$1966 ( \2343 , \2339 , \2342 );
buf \U$1967 ( \2344 , \2343 );
not \U$1968 ( \2345 , \2344 );
not \U$1969 ( \2346 , \2345 );
not \U$1970 ( \2347 , \2346 );
not \U$1971 ( \2348 , \2347 );
not \U$1972 ( \2349 , \2348 );
or \U$1973 ( \2350 , \2324 , \2349 );
not \U$1974 ( \2351 , RIc226f20_15);
not \U$1975 ( \2352 , \2351 );
buf \U$1976 ( \2353 , \2343 );
buf \U$1977 ( \2354 , \2353 );
not \U$1978 ( \2355 , \2354 );
nand \U$1979 ( \2356 , \2352 , \2355 );
nand \U$1980 ( \2357 , \2350 , \2356 );
buf \U$1981 ( \2358 , \2318 );
and \U$1982 ( \2359 , \2357 , \2358 );
nor \U$1983 ( \2360 , \2323 , \2359 );
not \U$1984 ( \2361 , \2360 );
not \U$1985 ( \2362 , \2361 );
and \U$1986 ( \2363 , RIc226bd8_22, RIc226b60_23);
not \U$1987 ( \2364 , RIc226bd8_22);
and \U$1988 ( \2365 , \2364 , \1927 );
nor \U$1989 ( \2366 , \2363 , \2365 );
buf \U$1990 ( \2367 , \2366 );
not \U$1991 ( \2368 , \2367 );
not \U$1992 ( \2369 , \1223 );
not \U$1993 ( \2370 , RIc226c50_21);
not \U$1994 ( \2371 , \2370 );
or \U$1995 ( \2372 , \2369 , \2371 );
not \U$1996 ( \2373 , \1440 );
not \U$1997 ( \2374 , \2373 );
nand \U$1998 ( \2375 , \2374 , RIc226c50_21);
nand \U$1999 ( \2376 , \2372 , \2375 );
not \U$2000 ( \2377 , \2376 );
or \U$2001 ( \2378 , \2368 , \2377 );
not \U$2002 ( \2379 , RIc226c50_21);
not \U$2003 ( \2380 , \1391 );
not \U$2004 ( \2381 , \2380 );
or \U$2005 ( \2382 , \2379 , \2381 );
not \U$2006 ( \2383 , RIc226c50_21);
nand \U$2007 ( \2384 , \1396 , \2383 );
nand \U$2008 ( \2385 , \2382 , \2384 );
not \U$2009 ( \2386 , \2366 );
and \U$2010 ( \2387 , RIc226bd8_22, RIc226c50_21);
not \U$2011 ( \2388 , RIc226bd8_22);
and \U$2012 ( \2389 , \2388 , \2370 );
nor \U$2013 ( \2390 , \2387 , \2389 );
and \U$2014 ( \2391 , \2386 , \2390 );
buf \U$2015 ( \2392 , \2391 );
nand \U$2016 ( \2393 , \2385 , \2392 );
nand \U$2017 ( \2394 , \2378 , \2393 );
not \U$2018 ( \2395 , \2394 );
or \U$2019 ( \2396 , \2362 , \2395 );
or \U$2020 ( \2397 , \2394 , \2361 );
not \U$2021 ( \2398 , \1682 );
not \U$2022 ( \2399 , RIc227010_13);
nor \U$2023 ( \2400 , \902 , \426 );
not \U$2024 ( \2401 , \2400 );
not \U$2025 ( \2402 , \688 );
or \U$2026 ( \2403 , \2401 , \2402 );
not \U$2027 ( \2404 , \426 );
nand \U$2028 ( \2405 , \387 , \2404 , \1975 , \395 );
not \U$2029 ( \2406 , \2404 );
not \U$2030 ( \2407 , \760 );
or \U$2031 ( \2408 , \2406 , \2407 );
nand \U$2032 ( \2409 , \2408 , \773 );
not \U$2033 ( \2410 , \2409 );
nand \U$2034 ( \2411 , \387 , \740 , \2404 );
and \U$2035 ( \2412 , \2405 , \2410 , \2411 );
nand \U$2036 ( \2413 , \2403 , \2412 );
not \U$2037 ( \2414 , \775 );
nor \U$2038 ( \2415 , \2414 , \427 );
and \U$2039 ( \2416 , \2413 , \2415 );
not \U$2040 ( \2417 , \2413 );
not \U$2041 ( \2418 , \2415 );
and \U$2042 ( \2419 , \2417 , \2418 );
nor \U$2043 ( \2420 , \2416 , \2419 );
buf \U$2044 ( \2421 , \2420 );
buf \U$2045 ( \2422 , \2421 );
buf \U$2046 ( \2423 , \2422 );
not \U$2047 ( \2424 , \2423 );
not \U$2048 ( \2425 , \2424 );
or \U$2049 ( \2426 , \2399 , \2425 );
not \U$2050 ( \2427 , RIc227010_13);
nand \U$2051 ( \2428 , \2423 , \2427 );
nand \U$2052 ( \2429 , \2426 , \2428 );
not \U$2053 ( \2430 , \2429 );
or \U$2054 ( \2431 , \2398 , \2430 );
not \U$2055 ( \2432 , \416 );
not \U$2056 ( \2433 , \688 );
or \U$2057 ( \2434 , \2432 , \2433 );
not \U$2058 ( \2435 , \763 );
nand \U$2059 ( \2436 , \2434 , \2435 );
nand \U$2060 ( \2437 , \2404 , \773 );
not \U$2061 ( \2438 , \2437 );
and \U$2062 ( \2439 , \2436 , \2438 );
not \U$2063 ( \2440 , \2436 );
and \U$2064 ( \2441 , \2440 , \2437 );
nor \U$2065 ( \2442 , \2439 , \2441 );
buf \U$2066 ( \2443 , \2442 );
not \U$2067 ( \2444 , \2443 );
buf \U$2068 ( \2445 , \2444 );
and \U$2069 ( \2446 , \2445 , RIc227010_13);
not \U$2070 ( \2447 , \2445 );
and \U$2071 ( \2448 , \2447 , \1296 );
or \U$2072 ( \2449 , \2446 , \2448 );
nand \U$2073 ( \2450 , \1680 , \2449 );
nand \U$2074 ( \2451 , \2431 , \2450 );
nand \U$2075 ( \2452 , \2397 , \2451 );
nand \U$2076 ( \2453 , \2396 , \2452 );
xor \U$2077 ( \2454 , \2283 , \2453 );
not \U$2078 ( \2455 , \954 );
not \U$2079 ( \2456 , RIc2273d0_5);
nor \U$2080 ( \2457 , \1970 , \389 );
not \U$2081 ( \2458 , \2457 );
not \U$2082 ( \2459 , \688 );
or \U$2083 ( \2460 , \2458 , \2459 );
not \U$2084 ( \2461 , \389 );
not \U$2085 ( \2462 , \2461 );
not \U$2086 ( \2463 , \1975 );
or \U$2087 ( \2464 , \2462 , \2463 );
nand \U$2088 ( \2465 , \2464 , \729 );
not \U$2089 ( \2466 , \2465 );
nand \U$2090 ( \2467 , \2460 , \2466 );
not \U$2091 ( \2468 , \731 );
nor \U$2092 ( \2469 , \2468 , \388 );
and \U$2093 ( \2470 , \2467 , \2469 );
not \U$2094 ( \2471 , \2467 );
not \U$2095 ( \2472 , \2469 );
and \U$2096 ( \2473 , \2471 , \2472 );
nor \U$2097 ( \2474 , \2470 , \2473 );
buf \U$2098 ( \2475 , \2474 );
not \U$2099 ( \2476 , \2475 );
not \U$2100 ( \2477 , \2476 );
or \U$2101 ( \2478 , \2456 , \2477 );
buf \U$2102 ( \2479 , \2475 );
buf \U$2103 ( \2480 , \2479 );
nand \U$2104 ( \2481 , \2480 , \946 );
nand \U$2105 ( \2482 , \2478 , \2481 );
not \U$2106 ( \2483 , \2482 );
or \U$2107 ( \2484 , \2455 , \2483 );
not \U$2108 ( \2485 , RIc2273d0_5);
not \U$2109 ( \2486 , \1970 );
not \U$2110 ( \2487 , \2486 );
not \U$2111 ( \2488 , \688 );
or \U$2112 ( \2489 , \2487 , \2488 );
not \U$2113 ( \2490 , \1975 );
nand \U$2114 ( \2491 , \2489 , \2490 );
nand \U$2115 ( \2492 , \2461 , \729 );
not \U$2116 ( \2493 , \2492 );
and \U$2117 ( \2494 , \2491 , \2493 );
not \U$2118 ( \2495 , \2491 );
and \U$2119 ( \2496 , \2495 , \2492 );
nor \U$2120 ( \2497 , \2494 , \2496 );
buf \U$2121 ( \2498 , \2497 );
not \U$2122 ( \2499 , \2498 );
not \U$2123 ( \2500 , \2499 );
not \U$2124 ( \2501 , \2500 );
not \U$2125 ( \2502 , \2501 );
or \U$2126 ( \2503 , \2485 , \2502 );
not \U$2127 ( \2504 , \2501 );
nand \U$2128 ( \2505 , \2504 , \946 );
nand \U$2129 ( \2506 , \2503 , \2505 );
nand \U$2130 ( \2507 , \2506 , \951 );
nand \U$2131 ( \2508 , \2484 , \2507 );
not \U$2132 ( \2509 , RIc226cc8_20);
or \U$2133 ( \2510 , \2509 , RIc226c50_21);
or \U$2134 ( \2511 , \2370 , RIc226cc8_20);
nand \U$2135 ( \2512 , \2510 , \2511 );
not \U$2136 ( \2513 , \2512 );
and \U$2137 ( \2514 , \1941 , \2509 );
and \U$2138 ( \2515 , RIc226d40_19, RIc226cc8_20);
nor \U$2139 ( \2516 , \2514 , \2515 );
and \U$2140 ( \2517 , \2513 , \2516 );
buf \U$2141 ( \2518 , \2517 );
not \U$2142 ( \2519 , \2518 );
not \U$2143 ( \2520 , RIc226d40_19);
not \U$2144 ( \2521 , \1949 );
or \U$2145 ( \2522 , \2520 , \2521 );
not \U$2146 ( \2523 , RIc226d40_19);
nand \U$2147 ( \2524 , \1335 , \2523 );
nand \U$2148 ( \2525 , \2522 , \2524 );
not \U$2149 ( \2526 , \2525 );
or \U$2150 ( \2527 , \2519 , \2526 );
not \U$2151 ( \2528 , RIc226d40_19);
not \U$2152 ( \2529 , \1602 );
or \U$2153 ( \2530 , \2528 , \2529 );
nand \U$2154 ( \2531 , \1533 , \2523 );
nand \U$2155 ( \2532 , \2530 , \2531 );
not \U$2156 ( \2533 , \2513 );
buf \U$2157 ( \2534 , \2533 );
nand \U$2158 ( \2535 , \2532 , \2534 );
nand \U$2159 ( \2536 , \2527 , \2535 );
xor \U$2160 ( \2537 , \2508 , \2536 );
not \U$2161 ( \2538 , \1118 );
not \U$2162 ( \2539 , RIc2272e0_7);
not \U$2163 ( \2540 , \390 );
nor \U$2164 ( \2541 , \2540 , \1970 );
not \U$2165 ( \2542 , \2541 );
not \U$2166 ( \2543 , \688 );
or \U$2167 ( \2544 , \2542 , \2543 );
and \U$2168 ( \2545 , \1975 , \390 );
nor \U$2169 ( \2546 , \2545 , \732 );
nand \U$2170 ( \2547 , \2544 , \2546 );
nand \U$2171 ( \2548 , \393 , \735 );
not \U$2172 ( \2549 , \2548 );
and \U$2173 ( \2550 , \2547 , \2549 );
not \U$2174 ( \2551 , \2547 );
and \U$2175 ( \2552 , \2551 , \2548 );
nor \U$2176 ( \2553 , \2550 , \2552 );
not \U$2177 ( \2554 , \2553 );
buf \U$2178 ( \2555 , \2554 );
buf \U$2179 ( \2556 , \2555 );
not \U$2180 ( \2557 , \2556 );
or \U$2181 ( \2558 , \2539 , \2557 );
not \U$2182 ( \2559 , \2556 );
nand \U$2183 ( \2560 , \2559 , \1139 );
nand \U$2184 ( \2561 , \2558 , \2560 );
not \U$2185 ( \2562 , \2561 );
or \U$2186 ( \2563 , \2538 , \2562 );
not \U$2187 ( \2564 , RIc2272e0_7);
nand \U$2188 ( \2565 , \390 , \393 );
nor \U$2189 ( \2566 , \1970 , \2565 );
not \U$2190 ( \2567 , \2566 );
not \U$2191 ( \2568 , \688 );
or \U$2192 ( \2569 , \2567 , \2568 );
not \U$2193 ( \2570 , \2565 );
not \U$2194 ( \2571 , \2570 );
not \U$2195 ( \2572 , \1975 );
or \U$2196 ( \2573 , \2571 , \2572 );
and \U$2197 ( \2574 , \732 , \393 );
nor \U$2198 ( \2575 , \2574 , \736 );
nand \U$2199 ( \2576 , \2573 , \2575 );
not \U$2200 ( \2577 , \2576 );
nand \U$2201 ( \2578 , \2569 , \2577 );
nor \U$2202 ( \2579 , \726 , \738 );
and \U$2203 ( \2580 , \2578 , \2579 );
not \U$2204 ( \2581 , \2578 );
not \U$2205 ( \2582 , \2579 );
and \U$2206 ( \2583 , \2581 , \2582 );
nor \U$2207 ( \2584 , \2580 , \2583 );
buf \U$2208 ( \2585 , \2584 );
not \U$2209 ( \2586 , \2585 );
buf \U$2210 ( \2587 , \2586 );
not \U$2211 ( \2588 , \2587 );
or \U$2212 ( \2589 , \2564 , \2588 );
buf \U$2213 ( \2590 , \2584 );
not \U$2214 ( \2591 , \2590 );
buf \U$2215 ( \2592 , \2591 );
not \U$2216 ( \2593 , \2592 );
nand \U$2217 ( \2594 , \2593 , \1139 );
nand \U$2218 ( \2595 , \2589 , \2594 );
nand \U$2219 ( \2596 , \2595 , \1121 );
nand \U$2220 ( \2597 , \2563 , \2596 );
and \U$2221 ( \2598 , \2537 , \2597 );
and \U$2222 ( \2599 , \2508 , \2536 );
or \U$2223 ( \2600 , \2598 , \2599 );
and \U$2224 ( \2601 , \2454 , \2600 );
and \U$2225 ( \2602 , \2283 , \2453 );
or \U$2226 ( \2603 , \2601 , \2602 );
xor \U$2227 ( \2604 , \2166 , \2603 );
not \U$2228 ( \2605 , \1963 );
not \U$2229 ( \2606 , RIc226e30_17);
not \U$2230 ( \2607 , \1488 );
or \U$2231 ( \2608 , \2606 , \2607 );
not \U$2232 ( \2609 , \1487 );
nand \U$2233 ( \2610 , \2609 , \1935 );
nand \U$2234 ( \2611 , \2608 , \2610 );
not \U$2235 ( \2612 , \2611 );
or \U$2236 ( \2613 , \2605 , \2612 );
not \U$2237 ( \2614 , RIc226e30_17);
not \U$2238 ( \2615 , \1730 );
buf \U$2239 ( \2616 , \2615 );
not \U$2240 ( \2617 , \2616 );
or \U$2241 ( \2618 , \2614 , \2617 );
nand \U$2242 ( \2619 , \1730 , \1935 );
nand \U$2243 ( \2620 , \2618 , \2619 );
nand \U$2244 ( \2621 , \2620 , \1945 );
nand \U$2245 ( \2622 , \2613 , \2621 );
not \U$2246 ( \2623 , \854 );
not \U$2247 ( \2624 , \2048 );
not \U$2248 ( \2625 , \688 );
or \U$2249 ( \2626 , \2624 , \2625 );
nand \U$2250 ( \2627 , \2626 , \2029 );
nand \U$2251 ( \2628 , \717 , \691 );
not \U$2252 ( \2629 , \2628 );
and \U$2253 ( \2630 , \2627 , \2629 );
not \U$2254 ( \2631 , \2627 );
and \U$2255 ( \2632 , \2631 , \2628 );
nor \U$2256 ( \2633 , \2630 , \2632 );
buf \U$2257 ( \2634 , \2633 );
not \U$2258 ( \2635 , \2634 );
not \U$2259 ( \2636 , \2635 );
xor \U$2260 ( \2637 , RIc2275b0_1, \2636 );
not \U$2261 ( \2638 , \2637 );
or \U$2262 ( \2639 , \2623 , \2638 );
nand \U$2263 ( \2640 , \2045 , \1579 );
nand \U$2264 ( \2641 , \2639 , \2640 );
xor \U$2265 ( \2642 , \2622 , \2641 );
not \U$2266 ( \2643 , \1040 );
not \U$2267 ( \2644 , RIc2274c0_3);
not \U$2268 ( \2645 , \2065 );
not \U$2269 ( \2646 , \2645 );
or \U$2270 ( \2647 , \2644 , \2646 );
nand \U$2271 ( \2648 , \2065 , \1078 );
nand \U$2272 ( \2649 , \2647 , \2648 );
not \U$2273 ( \2650 , \2649 );
or \U$2274 ( \2651 , \2643 , \2650 );
not \U$2275 ( \2652 , RIc2274c0_3);
and \U$2276 ( \2653 , \2049 , \716 );
and \U$2277 ( \2654 , \2048 , \2653 );
not \U$2278 ( \2655 , \2654 );
not \U$2279 ( \2656 , \688 );
or \U$2280 ( \2657 , \2655 , \2656 );
and \U$2281 ( \2658 , \2030 , \2653 );
nand \U$2282 ( \2659 , \694 , \716 );
nand \U$2283 ( \2660 , \2659 , \696 );
nor \U$2284 ( \2661 , \2658 , \2660 );
nand \U$2285 ( \2662 , \2657 , \2661 );
not \U$2286 ( \2663 , \698 );
nor \U$2287 ( \2664 , \2663 , \408 );
and \U$2288 ( \2665 , \2662 , \2664 );
not \U$2289 ( \2666 , \2662 );
not \U$2290 ( \2667 , \2664 );
and \U$2291 ( \2668 , \2666 , \2667 );
nor \U$2292 ( \2669 , \2665 , \2668 );
not \U$2293 ( \2670 , \2669 );
buf \U$2294 ( \2671 , \2670 );
buf \U$2295 ( \2672 , \2671 );
not \U$2296 ( \2673 , \2672 );
or \U$2297 ( \2674 , \2652 , \2673 );
not \U$2298 ( \2675 , \2672 );
nand \U$2299 ( \2676 , \2675 , \1027 );
nand \U$2300 ( \2677 , \2674 , \2676 );
nand \U$2301 ( \2678 , \2677 , \1082 );
nand \U$2302 ( \2679 , \2651 , \2678 );
xor \U$2303 ( \2680 , \2642 , \2679 );
xor \U$2304 ( \2681 , \2106 , \2126 );
xor \U$2305 ( \2682 , \2681 , \2158 );
nor \U$2306 ( \2683 , \2680 , \2682 );
xor \U$2307 ( \2684 , \2394 , \2360 );
xor \U$2308 ( \2685 , \2684 , \2451 );
or \U$2309 ( \2686 , \2683 , \2685 );
nand \U$2310 ( \2687 , \2680 , \2682 );
nand \U$2311 ( \2688 , \2686 , \2687 );
and \U$2312 ( \2689 , RIc2267a0_31, RIc226728_32);
and \U$2313 ( \2690 , RIc226728_32, RIc2266b0_33);
not \U$2314 ( \2691 , RIc226728_32);
not \U$2315 ( \2692 , RIc2266b0_33);
and \U$2316 ( \2693 , \2691 , \2692 );
nor \U$2317 ( \2694 , \2690 , \2693 );
nor \U$2318 ( \2695 , RIc2267a0_31, RIc226728_32);
nor \U$2319 ( \2696 , \2689 , \2694 , \2695 );
buf \U$2320 ( \2697 , \2696 );
not \U$2321 ( \2698 , \2697 );
not \U$2322 ( \2699 , RIc2267a0_31);
not \U$2323 ( \2700 , \930 );
buf \U$2324 ( \2701 , \2700 );
not \U$2325 ( \2702 , \2701 );
or \U$2326 ( \2703 , \2699 , \2702 );
not \U$2327 ( \2704 , \2701 );
not \U$2328 ( \2705 , RIc2267a0_31);
nand \U$2329 ( \2706 , \2704 , \2705 );
nand \U$2330 ( \2707 , \2703 , \2706 );
not \U$2331 ( \2708 , \2707 );
or \U$2332 ( \2709 , \2698 , \2708 );
buf \U$2333 ( \2710 , \2694 );
buf \U$2334 ( \2711 , \2710 );
nand \U$2335 ( \2712 , \2711 , RIc2267a0_31);
nand \U$2336 ( \2713 , \2709 , \2712 );
not \U$2337 ( \2714 , \954 );
not \U$2338 ( \2715 , \2506 );
or \U$2339 ( \2716 , \2714 , \2715 );
not \U$2340 ( \2717 , RIc2273d0_5);
not \U$2341 ( \2718 , \2672 );
or \U$2342 ( \2719 , \2717 , \2718 );
buf \U$2343 ( \2720 , \2669 );
nand \U$2344 ( \2721 , \2720 , \946 );
nand \U$2345 ( \2722 , \2719 , \2721 );
nand \U$2346 ( \2723 , \2722 , \951 );
nand \U$2347 ( \2724 , \2716 , \2723 );
xor \U$2348 ( \2725 , \2713 , \2724 );
not \U$2349 ( \2726 , \1040 );
not \U$2350 ( \2727 , RIc2274c0_3);
not \U$2351 ( \2728 , \2043 );
or \U$2352 ( \2729 , \2727 , \2728 );
buf \U$2353 ( \2730 , \2042 );
not \U$2354 ( \2731 , \2730 );
not \U$2355 ( \2732 , \2731 );
nand \U$2356 ( \2733 , \1032 , \2732 );
nand \U$2357 ( \2734 , \2729 , \2733 );
not \U$2358 ( \2735 , \2734 );
or \U$2359 ( \2736 , \2726 , \2735 );
nand \U$2360 ( \2737 , \2649 , \1082 );
nand \U$2361 ( \2738 , \2736 , \2737 );
and \U$2362 ( \2739 , \2725 , \2738 );
and \U$2363 ( \2740 , \2713 , \2724 );
or \U$2364 ( \2741 , \2739 , \2740 );
xor \U$2365 ( \2742 , \2197 , \2265 );
xor \U$2366 ( \2743 , \2742 , \2280 );
xor \U$2367 ( \2744 , \2741 , \2743 );
xor \U$2368 ( \2745 , \2508 , \2536 );
xor \U$2369 ( \2746 , \2745 , \2597 );
and \U$2370 ( \2747 , \2744 , \2746 );
and \U$2371 ( \2748 , \2741 , \2743 );
or \U$2372 ( \2749 , \2747 , \2748 );
xor \U$2373 ( \2750 , \2688 , \2749 );
xor \U$2374 ( \2751 , \2283 , \2453 );
xor \U$2375 ( \2752 , \2751 , \2600 );
and \U$2376 ( \2753 , \2750 , \2752 );
and \U$2377 ( \2754 , \2688 , \2749 );
or \U$2378 ( \2755 , \2753 , \2754 );
xor \U$2379 ( \2756 , \2604 , \2755 );
and \U$2380 ( \2757 , RIc2275b0_1, \2636 );
not \U$2381 ( \2758 , \2358 );
not \U$2382 ( \2759 , RIc226f20_15);
not \U$2383 ( \2760 , \2615 );
or \U$2384 ( \2761 , \2759 , \2760 );
not \U$2385 ( \2762 , \2616 );
nand \U$2386 ( \2763 , \2762 , \2351 );
nand \U$2387 ( \2764 , \2761 , \2763 );
not \U$2388 ( \2765 , \2764 );
or \U$2389 ( \2766 , \2758 , \2765 );
nand \U$2390 ( \2767 , \2357 , \2320 );
nand \U$2391 ( \2768 , \2766 , \2767 );
xor \U$2392 ( \2769 , \2757 , \2768 );
not \U$2393 ( \2770 , \1680 );
not \U$2394 ( \2771 , \2429 );
or \U$2395 ( \2772 , \2770 , \2771 );
not \U$2396 ( \2773 , RIc227010_13);
not \U$2397 ( \2774 , \2306 );
not \U$2398 ( \2775 , \2774 );
or \U$2399 ( \2776 , \2773 , \2775 );
nand \U$2400 ( \2777 , \2306 , \1758 );
nand \U$2401 ( \2778 , \2776 , \2777 );
nand \U$2402 ( \2779 , \2778 , \1682 );
nand \U$2403 ( \2780 , \2772 , \2779 );
and \U$2404 ( \2781 , \2769 , \2780 );
and \U$2405 ( \2782 , \2757 , \2768 );
or \U$2406 ( \2783 , \2781 , \2782 );
buf \U$2407 ( \2784 , \2078 );
or \U$2408 ( \2785 , \2784 , \2086 );
nand \U$2409 ( \2786 , \2785 , RIc226890_29);
not \U$2410 ( \2787 , \1930 );
not \U$2411 ( \2788 , \1921 );
or \U$2412 ( \2789 , \2787 , \2788 );
nand \U$2413 ( \2790 , \1915 , \2124 );
nand \U$2414 ( \2791 , \2789 , \2790 );
xor \U$2415 ( \2792 , \2786 , \2791 );
not \U$2416 ( \2793 , \2138 );
not \U$2417 ( \2794 , \2152 );
or \U$2418 ( \2795 , \2793 , \2794 );
not \U$2419 ( \2796 , RIc226980_27);
not \U$2420 ( \2797 , \932 );
or \U$2421 ( \2798 , \2796 , \2797 );
not \U$2422 ( \2799 , RIc226980_27);
nand \U$2423 ( \2800 , \931 , \2799 );
nand \U$2424 ( \2801 , \2798 , \2800 );
nand \U$2425 ( \2802 , \2801 , \2156 );
nand \U$2426 ( \2803 , \2795 , \2802 );
and \U$2427 ( \2804 , \2792 , \2803 );
and \U$2428 ( \2805 , \2786 , \2791 );
or \U$2429 ( \2806 , \2804 , \2805 );
xor \U$2430 ( \2807 , \2783 , \2806 );
not \U$2431 ( \2808 , \1340 );
and \U$2432 ( \2809 , \2258 , RIc2271f0_9);
not \U$2433 ( \2810 , \2258 );
and \U$2434 ( \2811 , \2810 , \1351 );
or \U$2435 ( \2812 , \2809 , \2811 );
not \U$2436 ( \2813 , \2812 );
or \U$2437 ( \2814 , \2808 , \2813 );
nand \U$2438 ( \2815 , \2278 , \1363 );
nand \U$2439 ( \2816 , \2814 , \2815 );
not \U$2440 ( \2817 , \2367 );
not \U$2441 ( \2818 , RIc226c50_21);
not \U$2442 ( \2819 , \1171 );
or \U$2443 ( \2820 , \2818 , \2819 );
nand \U$2444 ( \2821 , \1228 , \2370 );
nand \U$2445 ( \2822 , \2820 , \2821 );
not \U$2446 ( \2823 , \2822 );
or \U$2447 ( \2824 , \2817 , \2823 );
nand \U$2448 ( \2825 , \2376 , \2392 );
nand \U$2449 ( \2826 , \2824 , \2825 );
xor \U$2450 ( \2827 , \2816 , \2826 );
not \U$2451 ( \2828 , \1307 );
not \U$2452 ( \2829 , \2237 );
or \U$2453 ( \2830 , \2828 , \2829 );
not \U$2454 ( \2831 , RIc227100_11);
buf \U$2455 ( \2832 , \2442 );
not \U$2456 ( \2833 , \2832 );
buf \U$2457 ( \2834 , \2833 );
not \U$2458 ( \2835 , \2834 );
or \U$2459 ( \2836 , \2831 , \2835 );
not \U$2460 ( \2837 , \2834 );
nand \U$2461 ( \2838 , \2837 , \1291 );
nand \U$2462 ( \2839 , \2836 , \2838 );
nand \U$2463 ( \2840 , \2839 , \1311 );
nand \U$2464 ( \2841 , \2830 , \2840 );
and \U$2465 ( \2842 , \2827 , \2841 );
and \U$2466 ( \2843 , \2816 , \2826 );
or \U$2467 ( \2844 , \2842 , \2843 );
xor \U$2468 ( \2845 , \2807 , \2844 );
not \U$2469 ( \2846 , \2155 );
not \U$2470 ( \2847 , \2799 );
and \U$2471 ( \2848 , \2846 , \2847 );
and \U$2472 ( \2849 , \2801 , \2138 );
nor \U$2473 ( \2850 , \2848 , \2849 );
and \U$2474 ( \2851 , RIc2275b0_1, \2044 );
xor \U$2475 ( \2852 , \2850 , \2851 );
not \U$2476 ( \2853 , \1579 );
xor \U$2477 ( \2854 , RIc2275b0_1, \2675 );
not \U$2478 ( \2855 , \2854 );
or \U$2479 ( \2856 , \2853 , \2855 );
nand \U$2480 ( \2857 , \2066 , \854 );
nand \U$2481 ( \2858 , \2856 , \2857 );
xor \U$2482 ( \2859 , \2852 , \2858 );
buf \U$2483 ( \2860 , \2195 );
not \U$2484 ( \2861 , \2860 );
not \U$2485 ( \2862 , \2181 );
or \U$2486 ( \2863 , \2861 , \2862 );
not \U$2487 ( \2864 , RIc226a70_25);
not \U$2488 ( \2865 , \889 );
not \U$2489 ( \2866 , \2865 );
or \U$2490 ( \2867 , \2864 , \2866 );
nand \U$2491 ( \2868 , \891 , \1905 );
nand \U$2492 ( \2869 , \2867 , \2868 );
nand \U$2493 ( \2870 , \2869 , \2173 );
nand \U$2494 ( \2871 , \2863 , \2870 );
not \U$2495 ( \2872 , \2534 );
not \U$2496 ( \2873 , RIc226d40_19);
not \U$2497 ( \2874 , \1396 );
not \U$2498 ( \2875 , \2874 );
or \U$2499 ( \2876 , \2873 , \2875 );
nand \U$2500 ( \2877 , \1396 , \1941 );
nand \U$2501 ( \2878 , \2876 , \2877 );
not \U$2502 ( \2879 , \2878 );
or \U$2503 ( \2880 , \2872 , \2879 );
nand \U$2504 ( \2881 , \2532 , \2518 );
nand \U$2505 ( \2882 , \2880 , \2881 );
xor \U$2506 ( \2883 , \2871 , \2882 );
not \U$2507 ( \2884 , \1121 );
not \U$2508 ( \2885 , \2020 );
or \U$2509 ( \2886 , \2884 , \2885 );
nand \U$2510 ( \2887 , \2595 , \1118 );
nand \U$2511 ( \2888 , \2886 , \2887 );
and \U$2512 ( \2889 , \2883 , \2888 );
and \U$2513 ( \2890 , \2871 , \2882 );
or \U$2514 ( \2891 , \2889 , \2890 );
xor \U$2515 ( \2892 , \2859 , \2891 );
not \U$2516 ( \2893 , \1082 );
not \U$2517 ( \2894 , \2498 );
not \U$2518 ( \2895 , \2894 );
not \U$2519 ( \2896 , RIc2274c0_3);
and \U$2520 ( \2897 , \2895 , \2896 );
not \U$2521 ( \2898 , \2895 );
and \U$2522 ( \2899 , \2898 , RIc2274c0_3);
or \U$2523 ( \2900 , \2897 , \2899 );
not \U$2524 ( \2901 , \2900 );
or \U$2525 ( \2902 , \2893 , \2901 );
nand \U$2526 ( \2903 , \2677 , \1040 );
nand \U$2527 ( \2904 , \2902 , \2903 );
not \U$2528 ( \2905 , \951 );
not \U$2529 ( \2906 , \2482 );
or \U$2530 ( \2907 , \2905 , \2906 );
not \U$2531 ( \2908 , RIc2273d0_5);
not \U$2532 ( \2909 , \2556 );
or \U$2533 ( \2910 , \2908 , \2909 );
nand \U$2534 ( \2911 , \2559 , \946 );
nand \U$2535 ( \2912 , \2910 , \2911 );
nand \U$2536 ( \2913 , \2912 , \954 );
nand \U$2537 ( \2914 , \2907 , \2913 );
xor \U$2538 ( \2915 , \2904 , \2914 );
not \U$2539 ( \2916 , \1945 );
not \U$2540 ( \2917 , \2611 );
or \U$2541 ( \2918 , \2916 , \2917 );
nand \U$2542 ( \2919 , \1963 , \1954 );
nand \U$2543 ( \2920 , \2918 , \2919 );
and \U$2544 ( \2921 , \2915 , \2920 );
and \U$2545 ( \2922 , \2904 , \2914 );
or \U$2546 ( \2923 , \2921 , \2922 );
xor \U$2547 ( \2924 , \2892 , \2923 );
xor \U$2548 ( \2925 , \2845 , \2924 );
xor \U$2549 ( \2926 , \2871 , \2882 );
xor \U$2550 ( \2927 , \2926 , \2888 );
xor \U$2551 ( \2928 , \2816 , \2826 );
xor \U$2552 ( \2929 , \2928 , \2841 );
xor \U$2553 ( \2930 , \2927 , \2929 );
xor \U$2554 ( \2931 , \2904 , \2914 );
xor \U$2555 ( \2932 , \2931 , \2920 );
and \U$2556 ( \2933 , \2930 , \2932 );
and \U$2557 ( \2934 , \2927 , \2929 );
or \U$2558 ( \2935 , \2933 , \2934 );
xor \U$2559 ( \2936 , \2925 , \2935 );
xor \U$2560 ( \2937 , \2756 , \2936 );
xor \U$2561 ( \2938 , \2786 , \2791 );
xor \U$2562 ( \2939 , \2938 , \2803 );
xor \U$2563 ( \2940 , \2622 , \2641 );
and \U$2564 ( \2941 , \2940 , \2679 );
and \U$2565 ( \2942 , \2622 , \2641 );
or \U$2566 ( \2943 , \2941 , \2942 );
xor \U$2567 ( \2944 , \2939 , \2943 );
xor \U$2568 ( \2945 , \2757 , \2768 );
xor \U$2569 ( \2946 , \2945 , \2780 );
xor \U$2570 ( \2947 , \2944 , \2946 );
xor \U$2571 ( \2948 , \2927 , \2929 );
xor \U$2572 ( \2949 , \2948 , \2932 );
xor \U$2573 ( \2950 , \2947 , \2949 );
not \U$2574 ( \2951 , \2860 );
not \U$2575 ( \2952 , RIc226a70_25);
not \U$2576 ( \2953 , \1402 );
or \U$2577 ( \2954 , \2952 , \2953 );
nand \U$2578 ( \2955 , \1403 , \1905 );
nand \U$2579 ( \2956 , \2954 , \2955 );
not \U$2580 ( \2957 , \2956 );
or \U$2581 ( \2958 , \2951 , \2957 );
not \U$2582 ( \2959 , RIc226a70_25);
not \U$2583 ( \2960 , \1021 );
or \U$2584 ( \2961 , \2959 , \2960 );
not \U$2585 ( \2962 , \1021 );
nand \U$2586 ( \2963 , \2962 , \2187 );
nand \U$2587 ( \2964 , \2961 , \2963 );
nand \U$2588 ( \2965 , \2964 , \2173 );
nand \U$2589 ( \2966 , \2958 , \2965 );
not \U$2590 ( \2967 , \2966 );
not \U$2591 ( \2968 , \402 );
not \U$2592 ( \2969 , \2968 );
not \U$2593 ( \2970 , \688 );
or \U$2594 ( \2971 , \2969 , \2970 );
nand \U$2595 ( \2972 , \2971 , \706 );
not \U$2596 ( \2973 , \401 );
nand \U$2597 ( \2974 , \2973 , \703 );
not \U$2598 ( \2975 , \2974 );
and \U$2599 ( \2976 , \2972 , \2975 );
not \U$2600 ( \2977 , \2972 );
and \U$2601 ( \2978 , \2977 , \2974 );
nor \U$2602 ( \2979 , \2976 , \2978 );
buf \U$2603 ( \2980 , \2979 );
buf \U$2604 ( \2981 , \2980 );
nand \U$2605 ( \2982 , \2981 , RIc2275b0_1);
nand \U$2606 ( \2983 , \2967 , \2982 );
not \U$2607 ( \2984 , \2358 );
not \U$2608 ( \2985 , RIc226f20_15);
not \U$2609 ( \2986 , \2424 );
or \U$2610 ( \2987 , \2985 , \2986 );
nand \U$2611 ( \2988 , \2423 , \2301 );
nand \U$2612 ( \2989 , \2987 , \2988 );
not \U$2613 ( \2990 , \2989 );
or \U$2614 ( \2991 , \2984 , \2990 );
and \U$2615 ( \2992 , \2445 , RIc226f20_15);
not \U$2616 ( \2993 , \2445 );
and \U$2617 ( \2994 , \2993 , \2301 );
or \U$2618 ( \2995 , \2992 , \2994 );
nand \U$2619 ( \2996 , \2995 , \2320 );
nand \U$2620 ( \2997 , \2991 , \2996 );
and \U$2621 ( \2998 , \2983 , \2997 );
not \U$2622 ( \2999 , \2966 );
nor \U$2623 ( \3000 , \2999 , \2982 );
nor \U$2624 ( \3001 , \2998 , \3000 );
not \U$2625 ( \3002 , \3001 );
not \U$2626 ( \3003 , \3002 );
not \U$2627 ( \3004 , \951 );
not \U$2628 ( \3005 , RIc2273d0_5);
not \U$2629 ( \3006 , \2645 );
or \U$2630 ( \3007 , \3005 , \3006 );
buf \U$2631 ( \3008 , \2062 );
not \U$2632 ( \3009 , \3008 );
buf \U$2633 ( \3010 , \3009 );
buf \U$2634 ( \3011 , \3010 );
not \U$2635 ( \3012 , \3011 );
nand \U$2636 ( \3013 , \3012 , \946 );
nand \U$2637 ( \3014 , \3007 , \3013 );
not \U$2638 ( \3015 , \3014 );
or \U$2639 ( \3016 , \3004 , \3015 );
nand \U$2640 ( \3017 , \2722 , \954 );
nand \U$2641 ( \3018 , \3016 , \3017 );
not \U$2642 ( \3019 , \1118 );
not \U$2643 ( \3020 , RIc2272e0_7);
not \U$2644 ( \3021 , \2498 );
buf \U$2645 ( \3022 , \3021 );
buf \U$2646 ( \3023 , \3022 );
not \U$2647 ( \3024 , \3023 );
or \U$2648 ( \3025 , \3020 , \3024 );
not \U$2649 ( \3026 , \3023 );
not \U$2650 ( \3027 , RIc2272e0_7);
nand \U$2651 ( \3028 , \3026 , \3027 );
nand \U$2652 ( \3029 , \3025 , \3028 );
not \U$2653 ( \3030 , \3029 );
or \U$2654 ( \3031 , \3019 , \3030 );
not \U$2655 ( \3032 , RIc2272e0_7);
not \U$2656 ( \3033 , \2476 );
or \U$2657 ( \3034 , \3032 , \3033 );
not \U$2658 ( \3035 , \2475 );
not \U$2659 ( \3036 , \3035 );
nand \U$2660 ( \3037 , \3036 , \3027 );
nand \U$2661 ( \3038 , \3034 , \3037 );
nand \U$2662 ( \3039 , \3038 , \1121 );
nand \U$2663 ( \3040 , \3031 , \3039 );
or \U$2664 ( \3041 , \3018 , \3040 );
not \U$2665 ( \3042 , \2534 );
buf \U$2666 ( \3043 , \1484 );
not \U$2667 ( \3044 , \3043 );
and \U$2668 ( \3045 , \3044 , RIc226d40_19);
not \U$2669 ( \3046 , \3044 );
and \U$2670 ( \3047 , \3046 , \2523 );
or \U$2671 ( \3048 , \3045 , \3047 );
not \U$2672 ( \3049 , \3048 );
or \U$2673 ( \3050 , \3042 , \3049 );
not \U$2674 ( \3051 , RIc226d40_19);
not \U$2675 ( \3052 , \2615 );
or \U$2676 ( \3053 , \3051 , \3052 );
nand \U$2677 ( \3054 , \1730 , \2523 );
nand \U$2678 ( \3055 , \3053 , \3054 );
nand \U$2679 ( \3056 , \3055 , \2518 );
nand \U$2680 ( \3057 , \3050 , \3056 );
and \U$2681 ( \3058 , \3041 , \3057 );
and \U$2682 ( \3059 , \3040 , \3018 );
nor \U$2683 ( \3060 , \3058 , \3059 );
not \U$2684 ( \3061 , \3060 );
not \U$2685 ( \3062 , \3061 );
or \U$2686 ( \3063 , \3003 , \3062 );
not \U$2687 ( \3064 , \3060 );
not \U$2688 ( \3065 , \3001 );
or \U$2689 ( \3066 , \3064 , \3065 );
not \U$2690 ( \3067 , \2086 );
not \U$2691 ( \3068 , RIc226890_29);
not \U$2692 ( \3069 , \1074 );
or \U$2693 ( \3070 , \3068 , \3069 );
not \U$2694 ( \3071 , \1072 );
or \U$2695 ( \3072 , \3071 , RIc226890_29);
nand \U$2696 ( \3073 , \3070 , \3072 );
not \U$2697 ( \3074 , \3073 );
or \U$2698 ( \3075 , \3067 , \3074 );
not \U$2699 ( \3076 , \890 );
xor \U$2700 ( \3077 , RIc226890_29, \3076 );
nand \U$2701 ( \3078 , \3077 , \2078 );
nand \U$2702 ( \3079 , \3075 , \3078 );
not \U$2703 ( \3080 , \1963 );
not \U$2704 ( \3081 , RIc226e30_17);
not \U$2705 ( \3082 , \2355 );
or \U$2706 ( \3083 , \3081 , \3082 );
nand \U$2707 ( \3084 , \2354 , \1960 );
nand \U$2708 ( \3085 , \3083 , \3084 );
not \U$2709 ( \3086 , \3085 );
or \U$2710 ( \3087 , \3080 , \3086 );
not \U$2711 ( \3088 , RIc226e30_17);
not \U$2712 ( \3089 , \2298 );
or \U$2713 ( \3090 , \3088 , \3089 );
not \U$2714 ( \3091 , \2296 );
buf \U$2715 ( \3092 , \3091 );
buf \U$2716 ( \3093 , \3092 );
not \U$2717 ( \3094 , \3093 );
nand \U$2718 ( \3095 , \3094 , \1960 );
nand \U$2719 ( \3096 , \3090 , \3095 );
nand \U$2720 ( \3097 , \3096 , \1945 );
nand \U$2721 ( \3098 , \3087 , \3097 );
xor \U$2722 ( \3099 , \3079 , \3098 );
not \U$2723 ( \3100 , \1579 );
xor \U$2724 ( \3101 , RIc2275b0_1, \2105 );
not \U$2725 ( \3102 , \3101 );
or \U$2726 ( \3103 , \3100 , \3102 );
not \U$2727 ( \3104 , \403 );
not \U$2728 ( \3105 , \688 );
or \U$2729 ( \3106 , \3104 , \3105 );
not \U$2730 ( \3107 , \2096 );
nand \U$2731 ( \3108 , \3106 , \3107 );
nand \U$2732 ( \3109 , \711 , \701 );
not \U$2733 ( \3110 , \3109 );
and \U$2734 ( \3111 , \3108 , \3110 );
not \U$2735 ( \3112 , \3108 );
and \U$2736 ( \3113 , \3112 , \3109 );
nor \U$2737 ( \3114 , \3111 , \3113 );
buf \U$2738 ( \3115 , \3114 );
not \U$2739 ( \3116 , \3115 );
and \U$2740 ( \3117 , RIc2275b0_1, \3116 );
not \U$2741 ( \3118 , RIc2275b0_1);
not \U$2742 ( \3119 , \3115 );
not \U$2743 ( \3120 , \3119 );
not \U$2744 ( \3121 , \3120 );
not \U$2745 ( \3122 , \3121 );
and \U$2746 ( \3123 , \3118 , \3122 );
or \U$2747 ( \3124 , \3117 , \3123 );
nand \U$2748 ( \3125 , \854 , \3124 );
nand \U$2749 ( \3126 , \3103 , \3125 );
and \U$2750 ( \3127 , \3099 , \3126 );
and \U$2751 ( \3128 , \3079 , \3098 );
or \U$2752 ( \3129 , \3127 , \3128 );
nand \U$2753 ( \3130 , \3066 , \3129 );
nand \U$2754 ( \3131 , \3063 , \3130 );
or \U$2755 ( \3132 , \2697 , \2711 );
nand \U$2756 ( \3133 , \3132 , RIc2267a0_31);
not \U$2757 ( \3134 , \2078 );
not \U$2758 ( \3135 , \3073 );
or \U$2759 ( \3136 , \3134 , \3135 );
nand \U$2760 ( \3137 , \2083 , \2086 );
nand \U$2761 ( \3138 , \3136 , \3137 );
xor \U$2762 ( \3139 , \3133 , \3138 );
not \U$2763 ( \3140 , \2173 );
not \U$2764 ( \3141 , \2189 );
or \U$2765 ( \3142 , \3140 , \3141 );
nand \U$2766 ( \3143 , \2964 , \2195 );
nand \U$2767 ( \3144 , \3142 , \3143 );
and \U$2768 ( \3145 , \3139 , \3144 );
and \U$2769 ( \3146 , \3133 , \3138 );
or \U$2770 ( \3147 , \3145 , \3146 );
xor \U$2771 ( \3148 , \2088 , \3147 );
not \U$2772 ( \3149 , \3116 );
nand \U$2773 ( \3150 , \3149 , RIc2275b0_1);
not \U$2774 ( \3151 , \3150 );
not \U$2775 ( \3152 , \1579 );
not \U$2776 ( \3153 , \2637 );
or \U$2777 ( \3154 , \3152 , \3153 );
nand \U$2778 ( \3155 , \3101 , \854 );
nand \U$2779 ( \3156 , \3154 , \3155 );
not \U$2780 ( \3157 , \3156 );
not \U$2781 ( \3158 , \3157 );
or \U$2782 ( \3159 , \3151 , \3158 );
not \U$2783 ( \3160 , \1963 );
not \U$2784 ( \3161 , \2620 );
or \U$2785 ( \3162 , \3160 , \3161 );
nand \U$2786 ( \3163 , \3085 , \1945 );
nand \U$2787 ( \3164 , \3162 , \3163 );
nand \U$2788 ( \3165 , \3159 , \3164 );
not \U$2789 ( \3166 , \3150 );
nand \U$2790 ( \3167 , \3166 , \3156 );
nand \U$2791 ( \3168 , \3165 , \3167 );
xnor \U$2792 ( \3169 , \3148 , \3168 );
xor \U$2793 ( \3170 , \3131 , \3169 );
not \U$2794 ( \3171 , \1121 );
not \U$2795 ( \3172 , \2561 );
or \U$2796 ( \3173 , \3171 , \3172 );
nand \U$2797 ( \3174 , \3038 , \1118 );
nand \U$2798 ( \3175 , \3173 , \3174 );
not \U$2799 ( \3176 , \3175 );
not \U$2800 ( \3177 , \1340 );
not \U$2801 ( \3178 , \2271 );
or \U$2802 ( \3179 , \3177 , \3178 );
not \U$2803 ( \3180 , RIc2271f0_9);
not \U$2804 ( \3181 , \2592 );
or \U$2805 ( \3182 , \3180 , \3181 );
not \U$2806 ( \3183 , \2586 );
nand \U$2807 ( \3184 , \3183 , \1351 );
nand \U$2808 ( \3185 , \3182 , \3184 );
nand \U$2809 ( \3186 , \3185 , \1597 );
nand \U$2810 ( \3187 , \3179 , \3186 );
not \U$2811 ( \3188 , \3187 );
or \U$2812 ( \3189 , \3176 , \3188 );
or \U$2813 ( \3190 , \3175 , \3187 );
not \U$2814 ( \3191 , \2534 );
not \U$2815 ( \3192 , \2525 );
or \U$2816 ( \3193 , \3191 , \3192 );
nand \U$2817 ( \3194 , \3048 , \2518 );
nand \U$2818 ( \3195 , \3193 , \3194 );
nand \U$2819 ( \3196 , \3190 , \3195 );
nand \U$2820 ( \3197 , \3189 , \3196 );
not \U$2821 ( \3198 , \2367 );
not \U$2822 ( \3199 , \2385 );
or \U$2823 ( \3200 , \3198 , \3199 );
not \U$2824 ( \3201 , RIc226c50_21);
not \U$2825 ( \3202 , \1531 );
or \U$2826 ( \3203 , \3201 , \3202 );
not \U$2827 ( \3204 , RIc226c50_21);
nand \U$2828 ( \3205 , \1532 , \3204 );
nand \U$2829 ( \3206 , \3203 , \3205 );
nand \U$2830 ( \3207 , \2392 , \3206 );
nand \U$2831 ( \3208 , \3200 , \3207 );
not \U$2832 ( \3209 , \1311 );
not \U$2833 ( \3210 , \2263 );
or \U$2834 ( \3211 , \3209 , \3210 );
not \U$2835 ( \3212 , RIc227100_11);
not \U$2836 ( \3213 , \1990 );
or \U$2837 ( \3214 , \3212 , \3213 );
nand \U$2838 ( \3215 , \1991 , \1291 );
nand \U$2839 ( \3216 , \3214 , \3215 );
nand \U$2840 ( \3217 , \3216 , \1307 );
nand \U$2841 ( \3218 , \3211 , \3217 );
or \U$2842 ( \3219 , \3208 , \3218 );
not \U$2843 ( \3220 , \2156 );
not \U$2844 ( \3221 , \2144 );
or \U$2845 ( \3222 , \3220 , \3221 );
not \U$2846 ( \3223 , RIc226980_27);
not \U$2847 ( \3224 , \842 );
or \U$2848 ( \3225 , \3223 , \3224 );
nand \U$2849 ( \3226 , \2179 , \2150 );
nand \U$2850 ( \3227 , \3225 , \3226 );
nand \U$2851 ( \3228 , \3227 , \2138 );
nand \U$2852 ( \3229 , \3222 , \3228 );
nand \U$2853 ( \3230 , \3219 , \3229 );
nand \U$2854 ( \3231 , \3218 , \3208 );
nand \U$2855 ( \3232 , \3230 , \3231 );
and \U$2856 ( \3233 , \3197 , \3232 );
not \U$2857 ( \3234 , \3197 );
not \U$2858 ( \3235 , \3232 );
and \U$2859 ( \3236 , \3234 , \3235 );
nor \U$2860 ( \3237 , \3233 , \3236 );
not \U$2861 ( \3238 , \1915 );
not \U$2862 ( \3239 , RIc226b60_23);
not \U$2863 ( \3240 , \1222 );
or \U$2864 ( \3241 , \3239 , \3240 );
not \U$2865 ( \3242 , \1372 );
nand \U$2866 ( \3243 , \3242 , \1927 );
nand \U$2867 ( \3244 , \3241 , \3243 );
not \U$2868 ( \3245 , \3244 );
or \U$2869 ( \3246 , \3238 , \3245 );
nand \U$2870 ( \3247 , \2113 , \1930 );
nand \U$2871 ( \3248 , \3246 , \3247 );
not \U$2872 ( \3249 , \3248 );
not \U$2873 ( \3250 , \1679 );
not \U$2874 ( \3251 , \3250 );
not \U$2875 ( \3252 , RIc227010_13);
not \U$2876 ( \3253 , \2234 );
or \U$2877 ( \3254 , \3252 , \3253 );
nand \U$2878 ( \3255 , \2229 , \1758 );
nand \U$2879 ( \3256 , \3254 , \3255 );
not \U$2880 ( \3257 , \3256 );
or \U$2881 ( \3258 , \3251 , \3257 );
nand \U$2882 ( \3259 , \2449 , \1682 );
nand \U$2883 ( \3260 , \3258 , \3259 );
not \U$2884 ( \3261 , \3260 );
nand \U$2885 ( \3262 , \3249 , \3261 );
not \U$2886 ( \3263 , \2320 );
not \U$2887 ( \3264 , \2989 );
or \U$2888 ( \3265 , \3263 , \3264 );
not \U$2889 ( \3266 , \2308 );
nand \U$2890 ( \3267 , \3266 , \2358 );
nand \U$2891 ( \3268 , \3265 , \3267 );
and \U$2892 ( \3269 , \3262 , \3268 );
nor \U$2893 ( \3270 , \3261 , \3249 );
nor \U$2894 ( \3271 , \3269 , \3270 );
not \U$2895 ( \3272 , \3271 );
and \U$2896 ( \3273 , \3237 , \3272 );
not \U$2897 ( \3274 , \3237 );
and \U$2898 ( \3275 , \3274 , \3271 );
nor \U$2899 ( \3276 , \3273 , \3275 );
and \U$2900 ( \3277 , \3170 , \3276 );
and \U$2901 ( \3278 , \3131 , \3169 );
or \U$2902 ( \3279 , \3277 , \3278 );
and \U$2903 ( \3280 , \2950 , \3279 );
and \U$2904 ( \3281 , \2947 , \2949 );
or \U$2905 ( \3282 , \3280 , \3281 );
xor \U$2906 ( \3283 , \2939 , \2943 );
and \U$2907 ( \3284 , \3283 , \2946 );
and \U$2908 ( \3285 , \2939 , \2943 );
or \U$2909 ( \3286 , \3284 , \3285 );
not \U$2910 ( \3287 , \951 );
not \U$2911 ( \3288 , \2912 );
or \U$2912 ( \3289 , \3287 , \3288 );
not \U$2913 ( \3290 , RIc2273d0_5);
buf \U$2914 ( \3291 , \2590 );
not \U$2915 ( \3292 , \3291 );
not \U$2916 ( \3293 , \3292 );
or \U$2917 ( \3294 , \3290 , \3293 );
nand \U$2918 ( \3295 , \2593 , \946 );
nand \U$2919 ( \3296 , \3294 , \3295 );
nand \U$2920 ( \3297 , \3296 , \954 );
nand \U$2921 ( \3298 , \3289 , \3297 );
not \U$2922 ( \3299 , \3044 );
and \U$2923 ( \3300 , \2351 , \3299 );
not \U$2924 ( \3301 , \2351 );
and \U$2925 ( \3302 , \3301 , \1488 );
nor \U$2926 ( \3303 , \3300 , \3302 );
not \U$2927 ( \3304 , \3303 );
not \U$2928 ( \3305 , \2358 );
not \U$2929 ( \3306 , \3305 );
and \U$2930 ( \3307 , \3304 , \3306 );
and \U$2931 ( \3308 , \2764 , \2320 );
nor \U$2932 ( \3309 , \3307 , \3308 );
xor \U$2933 ( \3310 , \3298 , \3309 );
not \U$2934 ( \3311 , \1082 );
not \U$2935 ( \3312 , RIc2274c0_3);
not \U$2936 ( \3313 , \2480 );
not \U$2937 ( \3314 , \3313 );
or \U$2938 ( \3315 , \3312 , \3314 );
nand \U$2939 ( \3316 , \2480 , \2896 );
nand \U$2940 ( \3317 , \3315 , \3316 );
not \U$2941 ( \3318 , \3317 );
or \U$2942 ( \3319 , \3311 , \3318 );
nand \U$2943 ( \3320 , \2900 , \1040 );
nand \U$2944 ( \3321 , \3319 , \3320 );
xor \U$2945 ( \3322 , \3310 , \3321 );
not \U$2946 ( \3323 , \1597 );
not \U$2947 ( \3324 , \2812 );
or \U$2948 ( \3325 , \3323 , \3324 );
not \U$2949 ( \3326 , RIc2271f0_9);
not \U$2950 ( \3327 , \2230 );
or \U$2951 ( \3328 , \3326 , \3327 );
nand \U$2952 ( \3329 , \2235 , \1351 );
nand \U$2953 ( \3330 , \3328 , \3329 );
nand \U$2954 ( \3331 , \3330 , \1340 );
nand \U$2955 ( \3332 , \3325 , \3331 );
not \U$2956 ( \3333 , \2534 );
not \U$2957 ( \3334 , RIc226d40_19);
not \U$2958 ( \3335 , \1222 );
or \U$2959 ( \3336 , \3334 , \3335 );
not \U$2960 ( \3337 , \1441 );
not \U$2961 ( \3338 , RIc226d40_19);
nand \U$2962 ( \3339 , \3337 , \3338 );
nand \U$2963 ( \3340 , \3336 , \3339 );
not \U$2964 ( \3341 , \3340 );
or \U$2965 ( \3342 , \3333 , \3341 );
nand \U$2966 ( \3343 , \2518 , \2878 );
nand \U$2967 ( \3344 , \3342 , \3343 );
xor \U$2968 ( \3345 , \3332 , \3344 );
not \U$2969 ( \3346 , \1311 );
not \U$2970 ( \3347 , RIc227100_11);
buf \U$2971 ( \3348 , \2424 );
not \U$2972 ( \3349 , \3348 );
or \U$2973 ( \3350 , \3347 , \3349 );
not \U$2974 ( \3351 , RIc227100_11);
nand \U$2975 ( \3352 , \2423 , \3351 );
nand \U$2976 ( \3353 , \3350 , \3352 );
not \U$2977 ( \3354 , \3353 );
or \U$2978 ( \3355 , \3346 , \3354 );
nand \U$2979 ( \3356 , \2839 , \1307 );
nand \U$2980 ( \3357 , \3355 , \3356 );
xor \U$2981 ( \3358 , \3345 , \3357 );
xor \U$2982 ( \3359 , \3322 , \3358 );
not \U$2983 ( \3360 , \2173 );
and \U$2984 ( \3361 , RIc226a70_25, \1074 );
not \U$2985 ( \3362 , RIc226a70_25);
and \U$2986 ( \3363 , \3362 , \1073 );
or \U$2987 ( \3364 , \3361 , \3363 );
not \U$2988 ( \3365 , \3364 );
or \U$2989 ( \3366 , \3360 , \3365 );
nand \U$2990 ( \3367 , \2869 , \2860 );
nand \U$2991 ( \3368 , \3366 , \3367 );
not \U$2992 ( \3369 , \2392 );
not \U$2993 ( \3370 , \2822 );
or \U$2994 ( \3371 , \3369 , \3370 );
and \U$2995 ( \3372 , \3204 , \1022 );
not \U$2996 ( \3373 , \3204 );
and \U$2997 ( \3374 , \3373 , \1455 );
nor \U$2998 ( \3375 , \3372 , \3374 );
nand \U$2999 ( \3376 , \3375 , \2367 );
nand \U$3000 ( \3377 , \3371 , \3376 );
xor \U$3001 ( \3378 , \3368 , \3377 );
not \U$3002 ( \3379 , \1682 );
not \U$3003 ( \3380 , RIc227010_13);
not \U$3004 ( \3381 , \2355 );
or \U$3005 ( \3382 , \3380 , \3381 );
nand \U$3006 ( \3383 , \2348 , \1758 );
nand \U$3007 ( \3384 , \3382 , \3383 );
not \U$3008 ( \3385 , \3384 );
or \U$3009 ( \3386 , \3379 , \3385 );
nand \U$3010 ( \3387 , \1680 , \2778 );
nand \U$3011 ( \3388 , \3386 , \3387 );
xnor \U$3012 ( \3389 , \3378 , \3388 );
xor \U$3013 ( \3390 , \3359 , \3389 );
xor \U$3014 ( \3391 , \3286 , \3390 );
or \U$3015 ( \3392 , \3168 , \2089 );
nand \U$3016 ( \3393 , \3392 , \3147 );
nand \U$3017 ( \3394 , \2089 , \3168 );
and \U$3018 ( \3395 , \3393 , \3394 );
not \U$3019 ( \3396 , \3395 );
not \U$3020 ( \3397 , \3396 );
xor \U$3021 ( \3398 , \2068 , \2089 );
xor \U$3022 ( \3399 , \2161 , \3398 );
not \U$3023 ( \3400 , \3399 );
not \U$3024 ( \3401 , \3400 );
or \U$3025 ( \3402 , \3397 , \3401 );
not \U$3026 ( \3403 , \3399 );
not \U$3027 ( \3404 , \3395 );
or \U$3028 ( \3405 , \3403 , \3404 );
not \U$3029 ( \3406 , \3232 );
not \U$3030 ( \3407 , \3272 );
or \U$3031 ( \3408 , \3406 , \3407 );
not \U$3032 ( \3409 , \3235 );
not \U$3033 ( \3410 , \3271 );
or \U$3034 ( \3411 , \3409 , \3410 );
nand \U$3035 ( \3412 , \3411 , \3197 );
nand \U$3036 ( \3413 , \3408 , \3412 );
nand \U$3037 ( \3414 , \3405 , \3413 );
nand \U$3038 ( \3415 , \3402 , \3414 );
xor \U$3039 ( \3416 , \3391 , \3415 );
xor \U$3040 ( \3417 , \3282 , \3416 );
xor \U$3041 ( \3418 , \2688 , \2749 );
xor \U$3042 ( \3419 , \3418 , \2752 );
not \U$3043 ( \3420 , \3400 );
not \U$3044 ( \3421 , \3413 );
not \U$3045 ( \3422 , \3421 );
or \U$3046 ( \3423 , \3420 , \3422 );
nand \U$3047 ( \3424 , \3413 , \3399 );
nand \U$3048 ( \3425 , \3423 , \3424 );
and \U$3049 ( \3426 , \3425 , \3395 );
not \U$3050 ( \3427 , \3425 );
and \U$3051 ( \3428 , \3427 , \3396 );
nor \U$3052 ( \3429 , \3426 , \3428 );
not \U$3053 ( \3430 , \3429 );
or \U$3054 ( \3431 , \3419 , \3430 );
not \U$3055 ( \3432 , \2367 );
not \U$3056 ( \3433 , \3206 );
or \U$3057 ( \3434 , \3432 , \3433 );
not \U$3058 ( \3435 , RIc226c50_21);
not \U$3059 ( \3436 , \1333 );
or \U$3060 ( \3437 , \3435 , \3436 );
not \U$3061 ( \3438 , \1331 );
not \U$3062 ( \3439 , \3438 );
nand \U$3063 ( \3440 , \3439 , \2370 );
nand \U$3064 ( \3441 , \3437 , \3440 );
nand \U$3065 ( \3442 , \3441 , \2392 );
nand \U$3066 ( \3443 , \3434 , \3442 );
not \U$3067 ( \3444 , \1363 );
not \U$3068 ( \3445 , RIc2271f0_9);
buf \U$3069 ( \3446 , \2553 );
not \U$3070 ( \3447 , \3446 );
not \U$3071 ( \3448 , \3447 );
or \U$3072 ( \3449 , \3445 , \3448 );
not \U$3073 ( \3450 , \3447 );
nand \U$3074 ( \3451 , \3450 , \1342 );
nand \U$3075 ( \3452 , \3449 , \3451 );
not \U$3076 ( \3453 , \3452 );
or \U$3077 ( \3454 , \3444 , \3453 );
nand \U$3078 ( \3455 , \3185 , \1340 );
nand \U$3079 ( \3456 , \3454 , \3455 );
xor \U$3080 ( \3457 , \3443 , \3456 );
not \U$3081 ( \3458 , \2156 );
not \U$3082 ( \3459 , \3227 );
or \U$3083 ( \3460 , \3458 , \3459 );
not \U$3084 ( \3461 , RIc226980_27);
not \U$3085 ( \3462 , \1558 );
or \U$3086 ( \3463 , \3461 , \3462 );
not \U$3087 ( \3464 , \1557 );
nand \U$3088 ( \3465 , \3464 , \2133 );
nand \U$3089 ( \3466 , \3463 , \3465 );
nand \U$3090 ( \3467 , \3466 , \2138 );
nand \U$3091 ( \3468 , \3460 , \3467 );
and \U$3092 ( \3469 , \3457 , \3468 );
and \U$3093 ( \3470 , \3443 , \3456 );
or \U$3094 ( \3471 , \3469 , \3470 );
not \U$3095 ( \3472 , \3471 );
xor \U$3096 ( \3473 , \3150 , \3164 );
xor \U$3097 ( \3474 , \3473 , \3156 );
not \U$3098 ( \3475 , \3474 );
not \U$3099 ( \3476 , \3475 );
or \U$3100 ( \3477 , \3472 , \3476 );
not \U$3101 ( \3478 , \3471 );
not \U$3102 ( \3479 , \3478 );
not \U$3103 ( \3480 , \3474 );
or \U$3104 ( \3481 , \3479 , \3480 );
not \U$3105 ( \3482 , \1682 );
not \U$3106 ( \3483 , \3256 );
or \U$3107 ( \3484 , \3482 , \3483 );
not \U$3108 ( \3485 , RIc227010_13);
not \U$3109 ( \3486 , \2258 );
or \U$3110 ( \3487 , \3485 , \3486 );
nand \U$3111 ( \3488 , \2261 , \1296 );
nand \U$3112 ( \3489 , \3487 , \3488 );
nand \U$3113 ( \3490 , \3489 , \1680 );
nand \U$3114 ( \3491 , \3484 , \3490 );
not \U$3115 ( \3492 , \1930 );
not \U$3116 ( \3493 , \3244 );
or \U$3117 ( \3494 , \3492 , \3493 );
not \U$3118 ( \3495 , RIc226b60_23);
not \U$3119 ( \3496 , \1391 );
buf \U$3120 ( \3497 , \3496 );
not \U$3121 ( \3498 , \3497 );
or \U$3122 ( \3499 , \3495 , \3498 );
not \U$3123 ( \3500 , \3497 );
nand \U$3124 ( \3501 , \3500 , \1911 );
nand \U$3125 ( \3502 , \3499 , \3501 );
nand \U$3126 ( \3503 , \3502 , \1915 );
nand \U$3127 ( \3504 , \3494 , \3503 );
xor \U$3128 ( \3505 , \3491 , \3504 );
not \U$3129 ( \3506 , \1307 );
not \U$3130 ( \3507 , RIc227100_11);
buf \U$3131 ( \3508 , \2013 );
not \U$3132 ( \3509 , \3508 );
not \U$3133 ( \3510 , \3509 );
or \U$3134 ( \3511 , \3507 , \3510 );
nand \U$3135 ( \3512 , \3508 , \1291 );
nand \U$3136 ( \3513 , \3511 , \3512 );
not \U$3137 ( \3514 , \3513 );
or \U$3138 ( \3515 , \3506 , \3514 );
nand \U$3139 ( \3516 , \3216 , \1311 );
nand \U$3140 ( \3517 , \3515 , \3516 );
and \U$3141 ( \3518 , \3505 , \3517 );
and \U$3142 ( \3519 , \3491 , \3504 );
or \U$3143 ( \3520 , \3518 , \3519 );
nand \U$3144 ( \3521 , \3481 , \3520 );
nand \U$3145 ( \3522 , \3477 , \3521 );
xor \U$3146 ( \3523 , \2713 , \2724 );
xor \U$3147 ( \3524 , \3523 , \2738 );
not \U$3148 ( \3525 , \3524 );
xor \U$3149 ( \3526 , \3268 , \3260 );
xnor \U$3150 ( \3527 , \3526 , \3249 );
not \U$3151 ( \3528 , \3527 );
or \U$3152 ( \3529 , \3525 , \3528 );
or \U$3153 ( \3530 , \3527 , \3524 );
xor \U$3154 ( \3531 , \3133 , \3138 );
xor \U$3155 ( \3532 , \3531 , \3144 );
nand \U$3156 ( \3533 , \3530 , \3532 );
nand \U$3157 ( \3534 , \3529 , \3533 );
xor \U$3158 ( \3535 , \3522 , \3534 );
not \U$3159 ( \3536 , \2682 );
not \U$3160 ( \3537 , \2685 );
or \U$3161 ( \3538 , \3536 , \3537 );
or \U$3162 ( \3539 , \2685 , \2682 );
nand \U$3163 ( \3540 , \3538 , \3539 );
and \U$3164 ( \3541 , \3540 , \2680 );
not \U$3165 ( \3542 , \3540 );
not \U$3166 ( \3543 , \2680 );
and \U$3167 ( \3544 , \3542 , \3543 );
nor \U$3168 ( \3545 , \3541 , \3544 );
and \U$3169 ( \3546 , \3535 , \3545 );
and \U$3170 ( \3547 , \3522 , \3534 );
or \U$3171 ( \3548 , \3546 , \3547 );
nand \U$3172 ( \3549 , \3431 , \3548 );
nand \U$3173 ( \3550 , \3419 , \3430 );
nand \U$3174 ( \3551 , \3549 , \3550 );
xor \U$3175 ( \3552 , \3417 , \3551 );
xor \U$3176 ( \3553 , \2937 , \3552 );
xor \U$3177 ( \3554 , \3218 , \3229 );
xor \U$3178 ( \3555 , \3554 , \3208 );
xor \U$3179 ( \3556 , \3175 , \3187 );
xor \U$3180 ( \3557 , \3556 , \3195 );
xor \U$3181 ( \3558 , \3555 , \3557 );
not \U$3182 ( \3559 , \2713 );
not \U$3183 ( \3560 , \1082 );
not \U$3184 ( \3561 , \2734 );
or \U$3185 ( \3562 , \3560 , \3561 );
not \U$3186 ( \3563 , RIc2274c0_3);
not \U$3187 ( \3564 , \2636 );
not \U$3188 ( \3565 , \3564 );
or \U$3189 ( \3566 , \3563 , \3565 );
nand \U$3190 ( \3567 , \2636 , \1027 );
nand \U$3191 ( \3568 , \3566 , \3567 );
nand \U$3192 ( \3569 , \3568 , \1040 );
nand \U$3193 ( \3570 , \3562 , \3569 );
xor \U$3194 ( \3571 , \3559 , \3570 );
not \U$3195 ( \3572 , \1930 );
not \U$3196 ( \3573 , \3502 );
or \U$3197 ( \3574 , \3572 , \3573 );
not \U$3198 ( \3575 , RIc226b60_23);
not \U$3199 ( \3576 , \1530 );
or \U$3200 ( \3577 , \3575 , \3576 );
not \U$3201 ( \3578 , \1528 );
not \U$3202 ( \3579 , \3578 );
not \U$3203 ( \3580 , \3579 );
not \U$3204 ( \3581 , \3580 );
nand \U$3205 ( \3582 , \3581 , \2111 );
nand \U$3206 ( \3583 , \3577 , \3582 );
nand \U$3207 ( \3584 , \3583 , \1915 );
nand \U$3208 ( \3585 , \3574 , \3584 );
not \U$3209 ( \3586 , \1340 );
not \U$3210 ( \3587 , \3452 );
or \U$3211 ( \3588 , \3586 , \3587 );
not \U$3212 ( \3589 , \1351 );
not \U$3213 ( \3590 , \3036 );
or \U$3214 ( \3591 , \3589 , \3590 );
not \U$3215 ( \3592 , \2480 );
nand \U$3216 ( \3593 , \3592 , RIc2271f0_9);
nand \U$3217 ( \3594 , \3591 , \3593 );
nand \U$3218 ( \3595 , \3594 , \1597 );
nand \U$3219 ( \3596 , \3588 , \3595 );
xor \U$3220 ( \3597 , \3585 , \3596 );
not \U$3221 ( \3598 , \1311 );
not \U$3222 ( \3599 , \3513 );
or \U$3223 ( \3600 , \3598 , \3599 );
not \U$3224 ( \3601 , RIc227100_11);
not \U$3225 ( \3602 , \2587 );
or \U$3226 ( \3603 , \3601 , \3602 );
nand \U$3227 ( \3604 , \3183 , \3351 );
nand \U$3228 ( \3605 , \3603 , \3604 );
nand \U$3229 ( \3606 , \3605 , \1307 );
nand \U$3230 ( \3607 , \3600 , \3606 );
and \U$3231 ( \3608 , \3597 , \3607 );
and \U$3232 ( \3609 , \3585 , \3596 );
or \U$3233 ( \3610 , \3608 , \3609 );
and \U$3234 ( \3611 , \3571 , \3610 );
and \U$3235 ( \3612 , \3559 , \3570 );
or \U$3236 ( \3613 , \3611 , \3612 );
and \U$3237 ( \3614 , \3558 , \3613 );
and \U$3238 ( \3615 , \3555 , \3557 );
or \U$3239 ( \3616 , \3614 , \3615 );
xor \U$3240 ( \3617 , \2741 , \2743 );
xor \U$3241 ( \3618 , \3617 , \2746 );
xor \U$3242 ( \3619 , \3616 , \3618 );
not \U$3243 ( \3620 , RIc2265c0_35);
and \U$3244 ( \3621 , \3620 , RIc226638_34);
not \U$3245 ( \3622 , RIc226638_34);
and \U$3246 ( \3623 , \3622 , RIc2265c0_35);
nor \U$3247 ( \3624 , \3621 , \3623 );
and \U$3248 ( \3625 , \2692 , \3622 );
and \U$3249 ( \3626 , RIc2266b0_33, RIc226638_34);
nor \U$3250 ( \3627 , \3625 , \3626 );
and \U$3251 ( \3628 , \3624 , \3627 );
buf \U$3252 ( \3629 , \3628 );
not \U$3253 ( \3630 , \3624 );
buf \U$3254 ( \3631 , \3630 );
or \U$3255 ( \3632 , \3629 , \3631 );
nand \U$3256 ( \3633 , \3632 , RIc2266b0_33);
nand \U$3257 ( \3634 , \2968 , \706 );
not \U$3258 ( \3635 , \3634 );
not \U$3259 ( \3636 , \688 );
or \U$3260 ( \3637 , \3635 , \3636 );
or \U$3261 ( \3638 , \688 , \3634 );
nand \U$3262 ( \3639 , \3637 , \3638 );
buf \U$3263 ( \3640 , \3639 );
buf \U$3264 ( \3641 , \3640 );
and \U$3265 ( \3642 , \3641 , RIc2275b0_1);
xor \U$3266 ( \3643 , \3633 , \3642 );
not \U$3267 ( \3644 , \2697 );
not \U$3268 ( \3645 , RIc2267a0_31);
not \U$3269 ( \3646 , \3071 );
or \U$3270 ( \3647 , \3645 , \3646 );
not \U$3271 ( \3648 , RIc2267a0_31);
nand \U$3272 ( \3649 , \1072 , \3648 );
nand \U$3273 ( \3650 , \3647 , \3649 );
not \U$3274 ( \3651 , \3650 );
or \U$3275 ( \3652 , \3644 , \3651 );
buf \U$3276 ( \3653 , \2710 );
nand \U$3277 ( \3654 , \2707 , \3653 );
nand \U$3278 ( \3655 , \3652 , \3654 );
and \U$3279 ( \3656 , \3643 , \3655 );
and \U$3280 ( \3657 , \3633 , \3642 );
or \U$3281 ( \3658 , \3656 , \3657 );
not \U$3282 ( \3659 , \2154 );
not \U$3283 ( \3660 , \3466 );
or \U$3284 ( \3661 , \3659 , \3660 );
not \U$3285 ( \3662 , RIc226980_27);
not \U$3286 ( \3663 , \2120 );
or \U$3287 ( \3664 , \3662 , \3663 );
nand \U$3288 ( \3665 , \2962 , \2150 );
nand \U$3289 ( \3666 , \3664 , \3665 );
nand \U$3290 ( \3667 , \3666 , \2138 );
nand \U$3291 ( \3668 , \3661 , \3667 );
not \U$3292 ( \3669 , \2860 );
not \U$3293 ( \3670 , \1371 );
and \U$3294 ( \3671 , \3670 , RIc226a70_25);
not \U$3295 ( \3672 , \3670 );
and \U$3296 ( \3673 , \3672 , \1905 );
or \U$3297 ( \3674 , \3671 , \3673 );
not \U$3298 ( \3675 , \3674 );
or \U$3299 ( \3676 , \3669 , \3675 );
and \U$3300 ( \3677 , \1403 , \1905 );
not \U$3301 ( \3678 , \1403 );
and \U$3302 ( \3679 , \3678 , RIc226a70_25);
or \U$3303 ( \3680 , \3677 , \3679 );
nand \U$3304 ( \3681 , \3680 , \2173 );
nand \U$3305 ( \3682 , \3676 , \3681 );
xor \U$3306 ( \3683 , \3668 , \3682 );
not \U$3307 ( \3684 , \1945 );
not \U$3308 ( \3685 , RIc226e30_17);
not \U$3309 ( \3686 , \2421 );
not \U$3310 ( \3687 , \3686 );
or \U$3311 ( \3688 , \3685 , \3687 );
nand \U$3312 ( \3689 , \2423 , \1935 );
nand \U$3313 ( \3690 , \3688 , \3689 );
not \U$3314 ( \3691 , \3690 );
or \U$3315 ( \3692 , \3684 , \3691 );
nand \U$3316 ( \3693 , \3096 , \1963 );
nand \U$3317 ( \3694 , \3692 , \3693 );
and \U$3318 ( \3695 , \3683 , \3694 );
and \U$3319 ( \3696 , \3668 , \3682 );
or \U$3320 ( \3697 , \3695 , \3696 );
xor \U$3321 ( \3698 , \3658 , \3697 );
not \U$3322 ( \3699 , \2534 );
not \U$3323 ( \3700 , \3055 );
or \U$3324 ( \3701 , \3699 , \3700 );
not \U$3325 ( \3702 , RIc226d40_19);
not \U$3326 ( \3703 , \2347 );
or \U$3327 ( \3704 , \3702 , \3703 );
nand \U$3328 ( \3705 , \2348 , \2523 );
nand \U$3329 ( \3706 , \3704 , \3705 );
nand \U$3330 ( \3707 , \3706 , \2518 );
nand \U$3331 ( \3708 , \3701 , \3707 );
not \U$3332 ( \3709 , \1082 );
not \U$3333 ( \3710 , \3568 );
or \U$3334 ( \3711 , \3709 , \3710 );
not \U$3335 ( \3712 , RIc2274c0_3);
not \U$3336 ( \3713 , \2104 );
or \U$3337 ( \3714 , \3712 , \3713 );
not \U$3338 ( \3715 , \2103 );
not \U$3339 ( \3716 , \3715 );
nand \U$3340 ( \3717 , \3716 , \1027 );
nand \U$3341 ( \3718 , \3714 , \3717 );
nand \U$3342 ( \3719 , \3718 , \1040 );
nand \U$3343 ( \3720 , \3711 , \3719 );
xor \U$3344 ( \3721 , \3708 , \3720 );
not \U$3345 ( \3722 , \1579 );
not \U$3346 ( \3723 , \3124 );
or \U$3347 ( \3724 , \3722 , \3723 );
buf \U$3348 ( \3725 , \2979 );
not \U$3349 ( \3726 , \3725 );
buf \U$3350 ( \3727 , \3726 );
not \U$3351 ( \3728 , \3727 );
not \U$3352 ( \3729 , \3728 );
and \U$3353 ( \3730 , RIc2275b0_1, \3729 );
not \U$3354 ( \3731 , RIc2275b0_1);
buf \U$3355 ( \3732 , \3725 );
and \U$3356 ( \3733 , \3731 , \3732 );
or \U$3357 ( \3734 , \3730 , \3733 );
nand \U$3358 ( \3735 , \3734 , \854 );
nand \U$3359 ( \3736 , \3724 , \3735 );
and \U$3360 ( \3737 , \3721 , \3736 );
and \U$3361 ( \3738 , \3708 , \3720 );
or \U$3362 ( \3739 , \3737 , \3738 );
and \U$3363 ( \3740 , \3698 , \3739 );
and \U$3364 ( \3741 , \3658 , \3697 );
or \U$3365 ( \3742 , \3740 , \3741 );
not \U$3366 ( \3743 , \3742 );
not \U$3367 ( \3744 , \3520 );
not \U$3368 ( \3745 , \3478 );
or \U$3369 ( \3746 , \3744 , \3745 );
not \U$3370 ( \3747 , \3520 );
nand \U$3371 ( \3748 , \3747 , \3471 );
nand \U$3372 ( \3749 , \3746 , \3748 );
and \U$3373 ( \3750 , \3749 , \3475 );
not \U$3374 ( \3751 , \3749 );
and \U$3375 ( \3752 , \3751 , \3474 );
nor \U$3376 ( \3753 , \3750 , \3752 );
not \U$3377 ( \3754 , \3753 );
or \U$3378 ( \3755 , \3743 , \3754 );
or \U$3379 ( \3756 , \3753 , \3742 );
and \U$3380 ( \3757 , \3129 , \3060 );
not \U$3381 ( \3758 , \3129 );
and \U$3382 ( \3759 , \3758 , \3061 );
or \U$3383 ( \3760 , \3757 , \3759 );
and \U$3384 ( \3761 , \3760 , \3002 );
not \U$3385 ( \3762 , \3760 );
and \U$3386 ( \3763 , \3762 , \3001 );
nor \U$3387 ( \3764 , \3761 , \3763 );
nand \U$3388 ( \3765 , \3756 , \3764 );
nand \U$3389 ( \3766 , \3755 , \3765 );
and \U$3390 ( \3767 , \3619 , \3766 );
and \U$3391 ( \3768 , \3616 , \3618 );
or \U$3392 ( \3769 , \3767 , \3768 );
xor \U$3393 ( \3770 , \2947 , \2949 );
xor \U$3394 ( \3771 , \3770 , \3279 );
xor \U$3395 ( \3772 , \3769 , \3771 );
xor \U$3396 ( \3773 , \3131 , \3169 );
xor \U$3397 ( \3774 , \3773 , \3276 );
not \U$3398 ( \3775 , \3774 );
xor \U$3399 ( \3776 , \3522 , \3534 );
xor \U$3400 ( \3777 , \3776 , \3545 );
not \U$3401 ( \3778 , \3777 );
or \U$3402 ( \3779 , \3775 , \3778 );
or \U$3403 ( \3780 , \3774 , \3777 );
not \U$3404 ( \3781 , \2392 );
not \U$3405 ( \3782 , RIc226c50_21);
not \U$3406 ( \3783 , \3043 );
not \U$3407 ( \3784 , \3783 );
or \U$3408 ( \3785 , \3782 , \3784 );
nand \U$3409 ( \3786 , \3043 , \2383 );
nand \U$3410 ( \3787 , \3785 , \3786 );
not \U$3411 ( \3788 , \3787 );
or \U$3412 ( \3789 , \3781 , \3788 );
nand \U$3413 ( \3790 , \3441 , \2367 );
nand \U$3414 ( \3791 , \3789 , \3790 );
not \U$3415 ( \3792 , \954 );
not \U$3416 ( \3793 , \3014 );
or \U$3417 ( \3794 , \3792 , \3793 );
not \U$3418 ( \3795 , RIc2273d0_5);
not \U$3419 ( \3796 , \2731 );
or \U$3420 ( \3797 , \3795 , \3796 );
not \U$3421 ( \3798 , \2042 );
buf \U$3422 ( \3799 , \3798 );
not \U$3423 ( \3800 , \3799 );
nand \U$3424 ( \3801 , \3800 , \935 );
nand \U$3425 ( \3802 , \3797 , \3801 );
nand \U$3426 ( \3803 , \951 , \3802 );
nand \U$3427 ( \3804 , \3794 , \3803 );
xor \U$3428 ( \3805 , \3791 , \3804 );
not \U$3429 ( \3806 , \1121 );
not \U$3430 ( \3807 , \3029 );
or \U$3431 ( \3808 , \3806 , \3807 );
not \U$3432 ( \3809 , RIc2272e0_7);
not \U$3433 ( \3810 , \2720 );
not \U$3434 ( \3811 , \3810 );
or \U$3435 ( \3812 , \3809 , \3811 );
not \U$3436 ( \3813 , \2671 );
nand \U$3437 ( \3814 , \3813 , \1139 );
nand \U$3438 ( \3815 , \3812 , \3814 );
nand \U$3439 ( \3816 , \3815 , \1118 );
nand \U$3440 ( \3817 , \3808 , \3816 );
and \U$3441 ( \3818 , \3805 , \3817 );
and \U$3442 ( \3819 , \3791 , \3804 );
or \U$3443 ( \3820 , \3818 , \3819 );
not \U$3444 ( \3821 , \2086 );
not \U$3445 ( \3822 , \3077 );
or \U$3446 ( \3823 , \3821 , \3822 );
and \U$3447 ( \3824 , RIc226890_29, \1706 );
not \U$3448 ( \3825 , RIc226890_29);
and \U$3449 ( \3826 , \3825 , \841 );
or \U$3450 ( \3827 , \3824 , \3826 );
nand \U$3451 ( \3828 , \3827 , \2078 );
nand \U$3452 ( \3829 , \3823 , \3828 );
not \U$3453 ( \3830 , \1682 );
not \U$3454 ( \3831 , \3489 );
or \U$3455 ( \3832 , \3830 , \3831 );
not \U$3456 ( \3833 , RIc227010_13);
buf \U$3457 ( \3834 , \1988 );
not \U$3458 ( \3835 , \3834 );
not \U$3459 ( \3836 , \3835 );
or \U$3460 ( \3837 , \3833 , \3836 );
buf \U$3461 ( \3838 , \1988 );
not \U$3462 ( \3839 , \3838 );
not \U$3463 ( \3840 , \3839 );
not \U$3464 ( \3841 , RIc227010_13);
nand \U$3465 ( \3842 , \3840 , \3841 );
nand \U$3466 ( \3843 , \3837 , \3842 );
nand \U$3467 ( \3844 , \3843 , \3250 );
nand \U$3468 ( \3845 , \3832 , \3844 );
xor \U$3469 ( \3846 , \3829 , \3845 );
not \U$3470 ( \3847 , \2320 );
not \U$3471 ( \3848 , RIc226f20_15);
not \U$3472 ( \3849 , \2234 );
or \U$3473 ( \3850 , \3848 , \3849 );
not \U$3474 ( \3851 , \2234 );
nand \U$3475 ( \3852 , \3851 , \2351 );
nand \U$3476 ( \3853 , \3850 , \3852 );
not \U$3477 ( \3854 , \3853 );
or \U$3478 ( \3855 , \3847 , \3854 );
nand \U$3479 ( \3856 , \2995 , \2358 );
nand \U$3480 ( \3857 , \3855 , \3856 );
and \U$3481 ( \3858 , \3846 , \3857 );
and \U$3482 ( \3859 , \3829 , \3845 );
or \U$3483 ( \3860 , \3858 , \3859 );
xor \U$3484 ( \3861 , \3820 , \3860 );
xor \U$3485 ( \3862 , \3079 , \3098 );
xor \U$3486 ( \3863 , \3862 , \3126 );
and \U$3487 ( \3864 , \3861 , \3863 );
and \U$3488 ( \3865 , \3820 , \3860 );
or \U$3489 ( \3866 , \3864 , \3865 );
xor \U$3490 ( \3867 , \2982 , \2966 );
xnor \U$3491 ( \3868 , \3867 , \2997 );
xor \U$3492 ( \3869 , \3491 , \3504 );
xor \U$3493 ( \3870 , \3869 , \3517 );
xor \U$3494 ( \3871 , \3868 , \3870 );
xor \U$3495 ( \3872 , \3040 , \3018 );
xor \U$3496 ( \3873 , \3872 , \3057 );
and \U$3497 ( \3874 , \3871 , \3873 );
and \U$3498 ( \3875 , \3868 , \3870 );
or \U$3499 ( \3876 , \3874 , \3875 );
xor \U$3500 ( \3877 , \3866 , \3876 );
xor \U$3501 ( \3878 , \3532 , \3524 );
xor \U$3502 ( \3879 , \3878 , \3527 );
and \U$3503 ( \3880 , \3877 , \3879 );
and \U$3504 ( \3881 , \3866 , \3876 );
or \U$3505 ( \3882 , \3880 , \3881 );
nand \U$3506 ( \3883 , \3780 , \3882 );
nand \U$3507 ( \3884 , \3779 , \3883 );
and \U$3508 ( \3885 , \3772 , \3884 );
and \U$3509 ( \3886 , \3769 , \3771 );
or \U$3510 ( \3887 , \3885 , \3886 );
and \U$3511 ( \3888 , \3553 , \3887 );
not \U$3512 ( \3889 , \3553 );
not \U$3513 ( \3890 , \3887 );
and \U$3514 ( \3891 , \3889 , \3890 );
nor \U$3515 ( \3892 , \3888 , \3891 );
not \U$3516 ( \3893 , \3419 );
xor \U$3517 ( \3894 , \3548 , \3429 );
not \U$3518 ( \3895 , \3894 );
or \U$3519 ( \3896 , \3893 , \3895 );
or \U$3520 ( \3897 , \3894 , \3419 );
nand \U$3521 ( \3898 , \3896 , \3897 );
xor \U$3522 ( \3899 , \3769 , \3771 );
xor \U$3523 ( \3900 , \3899 , \3884 );
xor \U$3524 ( \3901 , \3898 , \3900 );
xor \U$3525 ( \3902 , \3616 , \3618 );
xor \U$3526 ( \3903 , \3902 , \3766 );
xor \U$3527 ( \3904 , \3555 , \3557 );
xor \U$3528 ( \3905 , \3904 , \3613 );
xor \U$3529 ( \3906 , \3443 , \3456 );
xor \U$3530 ( \3907 , \3906 , \3468 );
not \U$3531 ( \3908 , \3907 );
xor \U$3532 ( \3909 , \3559 , \3570 );
xor \U$3533 ( \3910 , \3909 , \3610 );
not \U$3534 ( \3911 , \3910 );
or \U$3535 ( \3912 , \3908 , \3911 );
or \U$3536 ( \3913 , \3910 , \3907 );
not \U$3537 ( \3914 , \1915 );
not \U$3538 ( \3915 , RIc226b60_23);
not \U$3539 ( \3916 , \1949 );
or \U$3540 ( \3917 , \3915 , \3916 );
not \U$3541 ( \3918 , \1948 );
nand \U$3542 ( \3919 , \3918 , \2111 );
nand \U$3543 ( \3920 , \3917 , \3919 );
not \U$3544 ( \3921 , \3920 );
or \U$3545 ( \3922 , \3914 , \3921 );
nand \U$3546 ( \3923 , \3583 , \1930 );
nand \U$3547 ( \3924 , \3922 , \3923 );
not \U$3548 ( \3925 , \3924 );
not \U$3549 ( \3926 , \1558 );
xor \U$3550 ( \3927 , RIc226890_29, \3926 );
not \U$3551 ( \3928 , \3927 );
not \U$3552 ( \3929 , \3928 );
not \U$3553 ( \3930 , \2784 );
not \U$3554 ( \3931 , \3930 );
and \U$3555 ( \3932 , \3929 , \3931 );
and \U$3556 ( \3933 , \3827 , \2086 );
nor \U$3557 ( \3934 , \3932 , \3933 );
not \U$3558 ( \3935 , \3934 );
not \U$3559 ( \3936 , \3935 );
or \U$3560 ( \3937 , \3925 , \3936 );
not \U$3561 ( \3938 , \3934 );
not \U$3562 ( \3939 , \3924 );
not \U$3563 ( \3940 , \3939 );
or \U$3564 ( \3941 , \3938 , \3940 );
not \U$3565 ( \3942 , \3250 );
not \U$3566 ( \3943 , RIc227010_13);
not \U$3567 ( \3944 , \2015 );
or \U$3568 ( \3945 , \3943 , \3944 );
nand \U$3569 ( \3946 , \2013 , \1296 );
nand \U$3570 ( \3947 , \3945 , \3946 );
not \U$3571 ( \3948 , \3947 );
or \U$3572 ( \3949 , \3942 , \3948 );
nand \U$3573 ( \3950 , \3843 , \1682 );
nand \U$3574 ( \3951 , \3949 , \3950 );
nand \U$3575 ( \3952 , \3941 , \3951 );
nand \U$3576 ( \3953 , \3937 , \3952 );
xor \U$3577 ( \3954 , \3633 , \3642 );
xor \U$3578 ( \3955 , \3954 , \3655 );
not \U$3579 ( \3956 , \3955 );
not \U$3580 ( \3957 , \2700 );
not \U$3581 ( \3958 , \3957 );
not \U$3582 ( \3959 , \2692 );
and \U$3583 ( \3960 , \3958 , \3959 );
and \U$3584 ( \3961 , \2704 , \2692 );
nor \U$3585 ( \3962 , \3960 , \3961 );
not \U$3586 ( \3963 , \3962 );
and \U$3587 ( \3964 , \3963 , \3629 );
not \U$3588 ( \3965 , \3631 );
nor \U$3589 ( \3966 , \3965 , \2692 );
nor \U$3590 ( \3967 , \3964 , \3966 );
nand \U$3591 ( \3968 , \3956 , \3967 );
and \U$3592 ( \3969 , \3953 , \3968 );
nor \U$3593 ( \3970 , \3956 , \3967 );
nor \U$3594 ( \3971 , \3969 , \3970 );
not \U$3595 ( \3972 , \3971 );
nand \U$3596 ( \3973 , \3913 , \3972 );
nand \U$3597 ( \3974 , \3912 , \3973 );
xor \U$3598 ( \3975 , \3905 , \3974 );
not \U$3599 ( \3976 , \2173 );
not \U$3600 ( \3977 , \3674 );
or \U$3601 ( \3978 , \3976 , \3977 );
not \U$3602 ( \3979 , RIc226a70_25);
not \U$3603 ( \3980 , \2380 );
or \U$3604 ( \3981 , \3979 , \3980 );
not \U$3605 ( \3982 , RIc226a70_25);
nand \U$3606 ( \3983 , \1396 , \3982 );
nand \U$3607 ( \3984 , \3981 , \3983 );
nand \U$3608 ( \3985 , \3984 , \2195 );
nand \U$3609 ( \3986 , \3978 , \3985 );
not \U$3610 ( \3987 , \3986 );
not \U$3611 ( \3988 , \3987 );
not \U$3612 ( \3989 , \2138 );
not \U$3613 ( \3990 , RIc226980_27);
not \U$3614 ( \3991 , \1402 );
or \U$3615 ( \3992 , \3990 , \3991 );
not \U$3616 ( \3993 , \1169 );
not \U$3617 ( \3994 , \3993 );
nand \U$3618 ( \3995 , \3994 , \2799 );
nand \U$3619 ( \3996 , \3992 , \3995 );
not \U$3620 ( \3997 , \3996 );
or \U$3621 ( \3998 , \3989 , \3997 );
nand \U$3622 ( \3999 , \3666 , \2154 );
nand \U$3623 ( \4000 , \3998 , \3999 );
not \U$3624 ( \4001 , \4000 );
not \U$3625 ( \4002 , \4001 );
or \U$3626 ( \4003 , \3988 , \4002 );
not \U$3627 ( \4004 , \2358 );
not \U$3628 ( \4005 , \3853 );
or \U$3629 ( \4006 , \4004 , \4005 );
not \U$3630 ( \4007 , RIc226f20_15);
buf \U$3631 ( \4008 , \2256 );
not \U$3632 ( \4009 , \4008 );
not \U$3633 ( \4010 , \4009 );
or \U$3634 ( \4011 , \4007 , \4010 );
nand \U$3635 ( \4012 , \4008 , \2301 );
nand \U$3636 ( \4013 , \4011 , \4012 );
nand \U$3637 ( \4014 , \4013 , \2320 );
nand \U$3638 ( \4015 , \4006 , \4014 );
nand \U$3639 ( \4016 , \4003 , \4015 );
nand \U$3640 ( \4017 , \4000 , \3986 );
nand \U$3641 ( \4018 , \4016 , \4017 );
not \U$3642 ( \4019 , \4018 );
not \U$3643 ( \4020 , \2711 );
not \U$3644 ( \4021 , \3650 );
or \U$3645 ( \4022 , \4020 , \4021 );
not \U$3646 ( \4023 , RIc2267a0_31);
not \U$3647 ( \4024 , \888 );
not \U$3648 ( \4025 , \4024 );
or \U$3649 ( \4026 , \4023 , \4025 );
nand \U$3650 ( \4027 , \889 , \2705 );
nand \U$3651 ( \4028 , \4026 , \4027 );
nand \U$3652 ( \4029 , \4028 , \2697 );
nand \U$3653 ( \4030 , \4022 , \4029 );
not \U$3654 ( \4031 , \1963 );
not \U$3655 ( \4032 , \3690 );
or \U$3656 ( \4033 , \4031 , \4032 );
not \U$3657 ( \4034 , RIc226e30_17);
not \U$3658 ( \4035 , \2834 );
or \U$3659 ( \4036 , \4034 , \4035 );
not \U$3660 ( \4037 , \2834 );
nand \U$3661 ( \4038 , \4037 , \1935 );
nand \U$3662 ( \4039 , \4036 , \4038 );
nand \U$3663 ( \4040 , \4039 , \1945 );
nand \U$3664 ( \4041 , \4033 , \4040 );
xor \U$3665 ( \4042 , \4030 , \4041 );
not \U$3666 ( \4043 , \1579 );
not \U$3667 ( \4044 , \3734 );
or \U$3668 ( \4045 , \4043 , \4044 );
not \U$3669 ( \4046 , \3641 );
and \U$3670 ( \4047 , RIc2275b0_1, \4046 );
not \U$3671 ( \4048 , RIc2275b0_1);
not \U$3672 ( \4049 , \3640 );
not \U$3673 ( \4050 , \4049 );
and \U$3674 ( \4051 , \4048 , \4050 );
or \U$3675 ( \4052 , \4047 , \4051 );
nand \U$3676 ( \4053 , \4052 , \854 );
nand \U$3677 ( \4054 , \4045 , \4053 );
and \U$3678 ( \4055 , \4042 , \4054 );
and \U$3679 ( \4056 , \4030 , \4041 );
or \U$3680 ( \4057 , \4055 , \4056 );
not \U$3681 ( \4058 , \4057 );
or \U$3682 ( \4059 , \4019 , \4058 );
or \U$3683 ( \4060 , \4018 , \4057 );
not \U$3684 ( \4061 , \555 );
nor \U$3685 ( \4062 , \4061 , \551 );
not \U$3686 ( \4063 , \4062 );
not \U$3687 ( \4064 , \648 );
not \U$3688 ( \4065 , \531 );
or \U$3689 ( \4066 , \4064 , \4065 );
not \U$3690 ( \4067 , \530 );
not \U$3691 ( \4068 , \652 );
and \U$3692 ( \4069 , \4067 , \4068 );
not \U$3693 ( \4070 , \651 );
nor \U$3694 ( \4071 , \4069 , \4070 );
nand \U$3695 ( \4072 , \4066 , \4071 );
not \U$3696 ( \4073 , \4072 );
or \U$3697 ( \4074 , \4063 , \4073 );
not \U$3698 ( \4075 , \551 );
and \U$3699 ( \4076 , \660 , \4075 );
not \U$3700 ( \4077 , \662 );
nor \U$3701 ( \4078 , \4076 , \4077 );
nand \U$3702 ( \4079 , \4074 , \4078 );
not \U$3703 ( \4080 , \4079 );
and \U$3704 ( \4081 , \594 , \596 );
and \U$3705 ( \4082 , \592 , \4081 );
nand \U$3706 ( \4083 , \521 , \477 , \4082 , \584 );
buf \U$3707 ( \4084 , \4083 );
nand \U$3708 ( \4085 , \532 , \4062 );
buf \U$3709 ( \4086 , \549 );
not \U$3710 ( \4087 , \4086 );
nor \U$3711 ( \4088 , \4085 , \4087 );
nand \U$3712 ( \4089 , \4084 , \4088 );
not \U$3713 ( \4090 , \4085 );
not \U$3714 ( \4091 , \636 );
not \U$3715 ( \4092 , \604 );
not \U$3716 ( \4093 , \595 );
not \U$3717 ( \4094 , \4093 );
and \U$3718 ( \4095 , \4092 , \4094 );
and \U$3719 ( \4096 , \607 , \595 , \608 );
not \U$3720 ( \4097 , \601 );
and \U$3721 ( \4098 , \4096 , \4097 );
nor \U$3722 ( \4099 , \4095 , \4098 );
not \U$3723 ( \4100 , \4099 );
or \U$3724 ( \4101 , \4091 , \4100 );
not \U$3725 ( \4102 , RIc224478_106);
not \U$3726 ( \4103 , RIc22a8c8_170);
and \U$3727 ( \4104 , \4102 , \4103 );
nor \U$3728 ( \4105 , \4104 , \634 );
not \U$3729 ( \4106 , \4105 );
not \U$3730 ( \4107 , \675 );
or \U$3731 ( \4108 , \4106 , \4107 );
nand \U$3732 ( \4109 , \4108 , \683 );
not \U$3733 ( \4110 , \4109 );
nand \U$3734 ( \4111 , \4101 , \4110 );
nand \U$3735 ( \4112 , \4090 , \4111 );
nand \U$3736 ( \4113 , \4080 , \4089 , \4112 );
not \U$3737 ( \4114 , \664 );
nor \U$3738 ( \4115 , \4114 , \550 );
and \U$3739 ( \4116 , \4113 , \4115 );
not \U$3740 ( \4117 , \4113 );
not \U$3741 ( \4118 , \4115 );
and \U$3742 ( \4119 , \4117 , \4118 );
nor \U$3743 ( \4120 , \4116 , \4119 );
buf \U$3744 ( \4121 , \4120 );
not \U$3745 ( \4122 , \4121 );
buf \U$3746 ( \4123 , \4122 );
not \U$3747 ( \4124 , \4123 );
and \U$3748 ( \4125 , \4124 , RIc2275b0_1);
not \U$3749 ( \4126 , \1082 );
not \U$3750 ( \4127 , \3718 );
or \U$3751 ( \4128 , \4126 , \4127 );
not \U$3752 ( \4129 , RIc2274c0_3);
not \U$3753 ( \4130 , \3116 );
or \U$3754 ( \4131 , \4129 , \4130 );
nand \U$3755 ( \4132 , \3120 , \2896 );
nand \U$3756 ( \4133 , \4131 , \4132 );
nand \U$3757 ( \4134 , \4133 , \1040 );
nand \U$3758 ( \4135 , \4128 , \4134 );
xor \U$3759 ( \4136 , \4125 , \4135 );
not \U$3760 ( \4137 , \2534 );
not \U$3761 ( \4138 , \3706 );
or \U$3762 ( \4139 , \4137 , \4138 );
not \U$3763 ( \4140 , RIc226d40_19);
not \U$3764 ( \4141 , \3093 );
or \U$3765 ( \4142 , \4140 , \4141 );
nand \U$3766 ( \4143 , \3094 , \3338 );
nand \U$3767 ( \4144 , \4142 , \4143 );
nand \U$3768 ( \4145 , \4144 , \2518 );
nand \U$3769 ( \4146 , \4139 , \4145 );
and \U$3770 ( \4147 , \4136 , \4146 );
and \U$3771 ( \4148 , \4125 , \4135 );
or \U$3772 ( \4149 , \4147 , \4148 );
nand \U$3773 ( \4150 , \4060 , \4149 );
nand \U$3774 ( \4151 , \4059 , \4150 );
xor \U$3775 ( \4152 , \3658 , \3697 );
xor \U$3776 ( \4153 , \4152 , \3739 );
xor \U$3777 ( \4154 , \4151 , \4153 );
xor \U$3778 ( \4155 , \3820 , \3860 );
xor \U$3779 ( \4156 , \4155 , \3863 );
and \U$3780 ( \4157 , \4154 , \4156 );
and \U$3781 ( \4158 , \4151 , \4153 );
or \U$3782 ( \4159 , \4157 , \4158 );
and \U$3783 ( \4160 , \3975 , \4159 );
and \U$3784 ( \4161 , \3905 , \3974 );
or \U$3785 ( \4162 , \4160 , \4161 );
xor \U$3786 ( \4163 , \3903 , \4162 );
xor \U$3787 ( \4164 , \3742 , \3753 );
buf \U$3788 ( \4165 , \3764 );
xor \U$3789 ( \4166 , \4164 , \4165 );
not \U$3790 ( \4167 , \4166 );
xor \U$3791 ( \4168 , \3866 , \3876 );
xor \U$3792 ( \4169 , \4168 , \3879 );
not \U$3793 ( \4170 , \4169 );
or \U$3794 ( \4171 , \4167 , \4170 );
or \U$3795 ( \4172 , \4169 , \4166 );
xor \U$3796 ( \4173 , \3668 , \3682 );
xor \U$3797 ( \4174 , \4173 , \3694 );
not \U$3798 ( \4175 , \2392 );
not \U$3799 ( \4176 , RIc226c50_21);
not \U$3800 ( \4177 , \1729 );
buf \U$3801 ( \4178 , \4177 );
not \U$3802 ( \4179 , \4178 );
or \U$3803 ( \4180 , \4176 , \4179 );
not \U$3804 ( \4181 , \1728 );
buf \U$3805 ( \4182 , \4181 );
not \U$3806 ( \4183 , \4182 );
nand \U$3807 ( \4184 , \4183 , \3204 );
nand \U$3808 ( \4185 , \4180 , \4184 );
not \U$3809 ( \4186 , \4185 );
or \U$3810 ( \4187 , \4175 , \4186 );
nand \U$3811 ( \4188 , \3787 , \2367 );
nand \U$3812 ( \4189 , \4187 , \4188 );
not \U$3813 ( \4190 , \4189 );
not \U$3814 ( \4191 , RIc2271f0_9);
not \U$3815 ( \4192 , \3022 );
or \U$3816 ( \4193 , \4191 , \4192 );
buf \U$3817 ( \4194 , \2497 );
not \U$3818 ( \4195 , \4194 );
not \U$3819 ( \4196 , \4195 );
nand \U$3820 ( \4197 , \4196 , \1342 );
nand \U$3821 ( \4198 , \4193 , \4197 );
and \U$3822 ( \4199 , \4198 , \1363 );
and \U$3823 ( \4200 , \3594 , \1340 );
nor \U$3824 ( \4201 , \4199 , \4200 );
nand \U$3825 ( \4202 , \4190 , \4201 );
not \U$3826 ( \4203 , \1307 );
not \U$3827 ( \4204 , RIc227100_11);
not \U$3828 ( \4205 , \3447 );
or \U$3829 ( \4206 , \4204 , \4205 );
nand \U$3830 ( \4207 , \3450 , \3351 );
nand \U$3831 ( \4208 , \4206 , \4207 );
not \U$3832 ( \4209 , \4208 );
or \U$3833 ( \4210 , \4203 , \4209 );
nand \U$3834 ( \4211 , \3605 , \1311 );
nand \U$3835 ( \4212 , \4210 , \4211 );
and \U$3836 ( \4213 , \4202 , \4212 );
nor \U$3837 ( \4214 , \4201 , \4190 );
nor \U$3838 ( \4215 , \4213 , \4214 );
not \U$3839 ( \4216 , \4215 );
or \U$3840 ( \4217 , \4174 , \4216 );
xor \U$3841 ( \4218 , \3708 , \3720 );
xor \U$3842 ( \4219 , \4218 , \3736 );
nand \U$3843 ( \4220 , \4217 , \4219 );
nand \U$3844 ( \4221 , \4174 , \4216 );
nand \U$3845 ( \4222 , \4220 , \4221 );
not \U$3846 ( \4223 , \954 );
not \U$3847 ( \4224 , \3802 );
or \U$3848 ( \4225 , \4223 , \4224 );
not \U$3849 ( \4226 , RIc2273d0_5);
not \U$3850 ( \4227 , \2634 );
buf \U$3851 ( \4228 , \4227 );
not \U$3852 ( \4229 , \4228 );
or \U$3853 ( \4230 , \4226 , \4229 );
nand \U$3854 ( \4231 , \2636 , \935 );
nand \U$3855 ( \4232 , \4230 , \4231 );
nand \U$3856 ( \4233 , \4232 , \951 );
nand \U$3857 ( \4234 , \4225 , \4233 );
xor \U$3858 ( \4235 , \3967 , \4234 );
not \U$3859 ( \4236 , \1118 );
not \U$3860 ( \4237 , RIc2272e0_7);
not \U$3861 ( \4238 , \3011 );
or \U$3862 ( \4239 , \4237 , \4238 );
buf \U$3863 ( \4240 , \3008 );
not \U$3864 ( \4241 , RIc2272e0_7);
nand \U$3865 ( \4242 , \4240 , \4241 );
nand \U$3866 ( \4243 , \4239 , \4242 );
not \U$3867 ( \4244 , \4243 );
or \U$3868 ( \4245 , \4236 , \4244 );
nand \U$3869 ( \4246 , \3815 , \1121 );
nand \U$3870 ( \4247 , \4245 , \4246 );
and \U$3871 ( \4248 , \4235 , \4247 );
and \U$3872 ( \4249 , \3967 , \4234 );
or \U$3873 ( \4250 , \4248 , \4249 );
xor \U$3874 ( \4251 , \3829 , \3845 );
xor \U$3875 ( \4252 , \4251 , \3857 );
xor \U$3876 ( \4253 , \4250 , \4252 );
xor \U$3877 ( \4254 , \3791 , \3804 );
xor \U$3878 ( \4255 , \4254 , \3817 );
and \U$3879 ( \4256 , \4253 , \4255 );
and \U$3880 ( \4257 , \4250 , \4252 );
or \U$3881 ( \4258 , \4256 , \4257 );
xor \U$3882 ( \4259 , \4222 , \4258 );
xor \U$3883 ( \4260 , \3868 , \3870 );
xor \U$3884 ( \4261 , \4260 , \3873 );
and \U$3885 ( \4262 , \4259 , \4261 );
and \U$3886 ( \4263 , \4222 , \4258 );
or \U$3887 ( \4264 , \4262 , \4263 );
nand \U$3888 ( \4265 , \4172 , \4264 );
nand \U$3889 ( \4266 , \4171 , \4265 );
and \U$3890 ( \4267 , \4163 , \4266 );
and \U$3891 ( \4268 , \3903 , \4162 );
or \U$3892 ( \4269 , \4267 , \4268 );
and \U$3893 ( \4270 , \3901 , \4269 );
and \U$3894 ( \4271 , \3898 , \3900 );
or \U$3895 ( \4272 , \4270 , \4271 );
nor \U$3896 ( \4273 , \3892 , \4272 );
not \U$3897 ( \4274 , \4273 );
xor \U$3898 ( \4275 , \3898 , \3900 );
xor \U$3899 ( \4276 , \4275 , \4269 );
xor \U$3900 ( \4277 , \3903 , \4162 );
xor \U$3901 ( \4278 , \4277 , \4266 );
xor \U$3902 ( \4279 , \3777 , \3882 );
xor \U$3903 ( \4280 , \4279 , \3774 );
or \U$3904 ( \4281 , \4278 , \4280 );
xor \U$3905 ( \4282 , \4222 , \4258 );
xor \U$3906 ( \4283 , \4282 , \4261 );
buf \U$3907 ( \4284 , \4283 );
not \U$3908 ( \4285 , \4284 );
xor \U$3909 ( \4286 , \4151 , \4153 );
xor \U$3910 ( \4287 , \4286 , \4156 );
not \U$3911 ( \4288 , \4287 );
or \U$3912 ( \4289 , \4285 , \4288 );
or \U$3913 ( \4290 , \4284 , \4287 );
xor \U$3914 ( \4291 , \4215 , \4174 );
xor \U$3915 ( \4292 , \4291 , \4219 );
xor \U$3916 ( \4293 , \4125 , \4135 );
xor \U$3917 ( \4294 , \4293 , \4146 );
xor \U$3918 ( \4295 , \3967 , \4234 );
xor \U$3919 ( \4296 , \4295 , \4247 );
xor \U$3920 ( \4297 , \4294 , \4296 );
xor \U$3921 ( \4298 , \4030 , \4041 );
xor \U$3922 ( \4299 , \4298 , \4054 );
and \U$3923 ( \4300 , \4297 , \4299 );
and \U$3924 ( \4301 , \4294 , \4296 );
or \U$3925 ( \4302 , \4300 , \4301 );
not \U$3926 ( \4303 , \4302 );
nand \U$3927 ( \4304 , \4292 , \4303 );
xor \U$3928 ( \4305 , \4250 , \4252 );
xor \U$3929 ( \4306 , \4305 , \4255 );
and \U$3930 ( \4307 , \4304 , \4306 );
nor \U$3931 ( \4308 , \4292 , \4303 );
nor \U$3932 ( \4309 , \4307 , \4308 );
not \U$3933 ( \4310 , \4309 );
nand \U$3934 ( \4311 , \4290 , \4310 );
nand \U$3935 ( \4312 , \4289 , \4311 );
not \U$3936 ( \4313 , \4312 );
xor \U$3937 ( \4314 , \3905 , \3974 );
xor \U$3938 ( \4315 , \4314 , \4159 );
not \U$3939 ( \4316 , \4315 );
or \U$3940 ( \4317 , \4313 , \4316 );
or \U$3941 ( \4318 , \4312 , \4315 );
not \U$3942 ( \4319 , \3971 );
not \U$3943 ( \4320 , \3907 );
and \U$3944 ( \4321 , \4319 , \4320 );
and \U$3945 ( \4322 , \3971 , \3907 );
nor \U$3946 ( \4323 , \4321 , \4322 );
and \U$3947 ( \4324 , \4323 , \3910 );
not \U$3948 ( \4325 , \4323 );
not \U$3949 ( \4326 , \3910 );
and \U$3950 ( \4327 , \4325 , \4326 );
nor \U$3951 ( \4328 , \4324 , \4327 );
not \U$3952 ( \4329 , \4328 );
xor \U$3953 ( \4330 , \3955 , \3967 );
xnor \U$3954 ( \4331 , \4330 , \3953 );
not \U$3955 ( \4332 , \3939 );
not \U$3956 ( \4333 , \3951 );
or \U$3957 ( \4334 , \4332 , \4333 );
or \U$3958 ( \4335 , \3951 , \3939 );
nand \U$3959 ( \4336 , \4334 , \4335 );
and \U$3960 ( \4337 , \4336 , \3934 );
not \U$3961 ( \4338 , \4336 );
and \U$3962 ( \4339 , \4338 , \3935 );
nor \U$3963 ( \4340 , \4337 , \4339 );
not \U$3964 ( \4341 , \4340 );
not \U$3965 ( \4342 , \4015 );
not \U$3966 ( \4343 , \4001 );
or \U$3967 ( \4344 , \4342 , \4343 );
or \U$3968 ( \4345 , \4015 , \4001 );
nand \U$3969 ( \4346 , \4344 , \4345 );
and \U$3970 ( \4347 , \4346 , \3987 );
not \U$3971 ( \4348 , \4346 );
and \U$3972 ( \4349 , \4348 , \3986 );
nor \U$3973 ( \4350 , \4347 , \4349 );
not \U$3974 ( \4351 , \4350 );
or \U$3975 ( \4352 , \4341 , \4351 );
xor \U$3976 ( \4353 , \4212 , \4190 );
xor \U$3977 ( \4354 , \4353 , \4201 );
nand \U$3978 ( \4355 , \4352 , \4354 );
not \U$3979 ( \4356 , \4350 );
not \U$3980 ( \4357 , \4340 );
nand \U$3981 ( \4358 , \4356 , \4357 );
nand \U$3982 ( \4359 , \4355 , \4358 );
xor \U$3983 ( \4360 , \4331 , \4359 );
xor \U$3984 ( \4361 , \4149 , \4018 );
xor \U$3985 ( \4362 , \4361 , \4057 );
and \U$3986 ( \4363 , \4360 , \4362 );
and \U$3987 ( \4364 , \4331 , \4359 );
or \U$3988 ( \4365 , \4363 , \4364 );
not \U$3989 ( \4366 , \4365 );
not \U$3990 ( \4367 , \4366 );
or \U$3991 ( \4368 , \4329 , \4367 );
xor \U$3992 ( \4369 , \3585 , \3596 );
xor \U$3993 ( \4370 , \4369 , \3607 );
not \U$3994 ( \4371 , RIc2264d0_37);
and \U$3995 ( \4372 , \4371 , RIc226548_36);
not \U$3996 ( \4373 , RIc226548_36);
and \U$3997 ( \4374 , \4373 , RIc2264d0_37);
nor \U$3998 ( \4375 , \4372 , \4374 );
not \U$3999 ( \4376 , RIc2265c0_35);
and \U$4000 ( \4377 , \4376 , \4373 );
and \U$4001 ( \4378 , RIc2265c0_35, RIc226548_36);
nor \U$4002 ( \4379 , \4377 , \4378 );
and \U$4003 ( \4380 , \4375 , \4379 );
buf \U$4004 ( \4381 , \4380 );
not \U$4005 ( \4382 , \4375 );
buf \U$4006 ( \4383 , \4382 );
or \U$4007 ( \4384 , \4381 , \4383 );
nand \U$4008 ( \4385 , \4384 , RIc2265c0_35);
not \U$4009 ( \4386 , \532 );
not \U$4010 ( \4387 , \4386 );
and \U$4011 ( \4388 , \4387 , \4086 , \555 );
nand \U$4012 ( \4389 , \4084 , \4388 );
not \U$4013 ( \4390 , \636 );
not \U$4014 ( \4391 , \4099 );
or \U$4015 ( \4392 , \4390 , \4391 );
nand \U$4016 ( \4393 , \4392 , \4110 );
not \U$4017 ( \4394 , \685 );
nor \U$4018 ( \4395 , \4394 , \4061 );
nand \U$4019 ( \4396 , \4393 , \4395 );
and \U$4020 ( \4397 , \555 , \4072 );
nor \U$4021 ( \4398 , \4397 , \660 );
nand \U$4022 ( \4399 , \4389 , \4396 , \4398 );
nand \U$4023 ( \4400 , \4075 , \662 );
not \U$4024 ( \4401 , \4400 );
and \U$4025 ( \4402 , \4399 , \4401 );
not \U$4026 ( \4403 , \4399 );
and \U$4027 ( \4404 , \4403 , \4400 );
nor \U$4028 ( \4405 , \4402 , \4404 );
buf \U$4029 ( \4406 , \4405 );
buf \U$4030 ( \4407 , \4406 );
and \U$4031 ( \4408 , RIc2275b0_1, \4407 );
xor \U$4032 ( \4409 , \4385 , \4408 );
not \U$4033 ( \4410 , \1579 );
not \U$4034 ( \4411 , \4052 );
or \U$4035 ( \4412 , \4410 , \4411 );
not \U$4036 ( \4413 , \4120 );
buf \U$4037 ( \4414 , \4413 );
and \U$4038 ( \4415 , RIc2275b0_1, \4414 );
not \U$4039 ( \4416 , RIc2275b0_1);
not \U$4040 ( \4417 , \4121 );
not \U$4041 ( \4418 , \4417 );
and \U$4042 ( \4419 , \4416 , \4418 );
or \U$4043 ( \4420 , \4415 , \4419 );
nand \U$4044 ( \4421 , \4420 , \854 );
nand \U$4045 ( \4422 , \4412 , \4421 );
and \U$4046 ( \4423 , \4409 , \4422 );
and \U$4047 ( \4424 , \4385 , \4408 );
or \U$4048 ( \4425 , \4423 , \4424 );
not \U$4049 ( \4426 , \2086 );
not \U$4050 ( \4427 , \3927 );
or \U$4051 ( \4428 , \4426 , \4427 );
not \U$4052 ( \4429 , RIc226890_29);
not \U$4053 ( \4430 , \1021 );
or \U$4054 ( \4431 , \4429 , \4430 );
not \U$4055 ( \4432 , \1020 );
or \U$4056 ( \4433 , \4432 , RIc226890_29);
nand \U$4057 ( \4434 , \4431 , \4433 );
nand \U$4058 ( \4435 , \4434 , \2078 );
nand \U$4059 ( \4436 , \4428 , \4435 );
buf \U$4060 ( \4437 , \4436 );
not \U$4061 ( \4438 , \4437 );
not \U$4062 ( \4439 , \3962 );
not \U$4063 ( \4440 , \3631 );
not \U$4064 ( \4441 , \4440 );
and \U$4065 ( \4442 , \4439 , \4441 );
and \U$4066 ( \4443 , \1072 , \2692 );
not \U$4067 ( \4444 , \1072 );
and \U$4068 ( \4445 , \4444 , RIc2266b0_33);
or \U$4069 ( \4446 , \4443 , \4445 );
and \U$4070 ( \4447 , \4446 , \3629 );
nor \U$4071 ( \4448 , \4442 , \4447 );
not \U$4072 ( \4449 , \4448 );
not \U$4073 ( \4450 , \4449 );
or \U$4074 ( \4451 , \4438 , \4450 );
or \U$4075 ( \4452 , \4437 , \4449 );
not \U$4076 ( \4453 , \2518 );
not \U$4077 ( \4454 , RIc226d40_19);
not \U$4078 ( \4455 , \3686 );
or \U$4079 ( \4456 , \4454 , \4455 );
not \U$4080 ( \4457 , \3686 );
nand \U$4081 ( \4458 , \4457 , \1941 );
nand \U$4082 ( \4459 , \4456 , \4458 );
not \U$4083 ( \4460 , \4459 );
or \U$4084 ( \4461 , \4453 , \4460 );
nand \U$4085 ( \4462 , \4144 , \2534 );
nand \U$4086 ( \4463 , \4461 , \4462 );
nand \U$4087 ( \4464 , \4452 , \4463 );
nand \U$4088 ( \4465 , \4451 , \4464 );
xor \U$4089 ( \4466 , \4425 , \4465 );
not \U$4090 ( \4467 , \2367 );
not \U$4091 ( \4468 , \4185 );
or \U$4092 ( \4469 , \4467 , \4468 );
not \U$4093 ( \4470 , RIc226c50_21);
not \U$4094 ( \4471 , \2345 );
or \U$4095 ( \4472 , \4470 , \4471 );
not \U$4096 ( \4473 , \2353 );
not \U$4097 ( \4474 , \4473 );
not \U$4098 ( \4475 , RIc226c50_21);
nand \U$4099 ( \4476 , \4474 , \4475 );
nand \U$4100 ( \4477 , \4472 , \4476 );
nand \U$4101 ( \4478 , \4477 , \2392 );
nand \U$4102 ( \4479 , \4469 , \4478 );
not \U$4103 ( \4480 , \4479 );
not \U$4104 ( \4481 , \1040 );
not \U$4105 ( \4482 , RIc2274c0_3);
not \U$4106 ( \4483 , \3727 );
or \U$4107 ( \4484 , \4482 , \4483 );
nand \U$4108 ( \4485 , \3732 , \2896 );
nand \U$4109 ( \4486 , \4484 , \4485 );
not \U$4110 ( \4487 , \4486 );
or \U$4111 ( \4488 , \4481 , \4487 );
nand \U$4112 ( \4489 , \4133 , \1082 );
nand \U$4113 ( \4490 , \4488 , \4489 );
not \U$4114 ( \4491 , \4490 );
or \U$4115 ( \4492 , \4480 , \4491 );
or \U$4116 ( \4493 , \4490 , \4479 );
not \U$4117 ( \4494 , \954 );
not \U$4118 ( \4495 , \4232 );
or \U$4119 ( \4496 , \4494 , \4495 );
not \U$4120 ( \4497 , RIc2273d0_5);
not \U$4121 ( \4498 , \2104 );
or \U$4122 ( \4499 , \4497 , \4498 );
buf \U$4123 ( \4500 , \2103 );
buf \U$4124 ( \4501 , \4500 );
nand \U$4125 ( \4502 , \4501 , \946 );
nand \U$4126 ( \4503 , \4499 , \4502 );
nand \U$4127 ( \4504 , \4503 , \951 );
nand \U$4128 ( \4505 , \4496 , \4504 );
nand \U$4129 ( \4506 , \4493 , \4505 );
nand \U$4130 ( \4507 , \4492 , \4506 );
and \U$4131 ( \4508 , \4466 , \4507 );
and \U$4132 ( \4509 , \4425 , \4465 );
or \U$4133 ( \4510 , \4508 , \4509 );
xor \U$4134 ( \4511 , \4370 , \4510 );
not \U$4135 ( \4512 , \2358 );
not \U$4136 ( \4513 , \4013 );
or \U$4137 ( \4514 , \4512 , \4513 );
not \U$4138 ( \4515 , RIc226f20_15);
not \U$4139 ( \4516 , \1989 );
or \U$4140 ( \4517 , \4515 , \4516 );
nand \U$4141 ( \4518 , \3838 , \1674 );
nand \U$4142 ( \4519 , \4517 , \4518 );
nand \U$4143 ( \4520 , \4519 , \2320 );
nand \U$4144 ( \4521 , \4514 , \4520 );
not \U$4145 ( \4522 , \2154 );
not \U$4146 ( \4523 , \3996 );
or \U$4147 ( \4524 , \4522 , \4523 );
not \U$4148 ( \4525 , RIc226980_27);
not \U$4149 ( \4526 , \1372 );
or \U$4150 ( \4527 , \4525 , \4526 );
not \U$4151 ( \4528 , RIc226980_27);
nand \U$4152 ( \4529 , \1223 , \4528 );
nand \U$4153 ( \4530 , \4527 , \4529 );
nand \U$4154 ( \4531 , \4530 , \2138 );
nand \U$4155 ( \4532 , \4524 , \4531 );
or \U$4156 ( \4533 , \4521 , \4532 );
not \U$4157 ( \4534 , \1945 );
not \U$4158 ( \4535 , RIc226e30_17);
not \U$4159 ( \4536 , \2228 );
or \U$4160 ( \4537 , \4535 , \4536 );
nand \U$4161 ( \4538 , \3851 , \1935 );
nand \U$4162 ( \4539 , \4537 , \4538 );
not \U$4163 ( \4540 , \4539 );
or \U$4164 ( \4541 , \4534 , \4540 );
nand \U$4165 ( \4542 , \4039 , \1963 );
nand \U$4166 ( \4543 , \4541 , \4542 );
nand \U$4167 ( \4544 , \4533 , \4543 );
nand \U$4168 ( \4545 , \4521 , \4532 );
nand \U$4169 ( \4546 , \4544 , \4545 );
not \U$4170 ( \4547 , \4546 );
not \U$4171 ( \4548 , \4547 );
not \U$4172 ( \4549 , \1930 );
not \U$4173 ( \4550 , \3920 );
or \U$4174 ( \4551 , \4549 , \4550 );
not \U$4175 ( \4552 , RIc226b60_23);
not \U$4176 ( \4553 , \3044 );
or \U$4177 ( \4554 , \4552 , \4553 );
nand \U$4178 ( \4555 , \1486 , \1927 );
nand \U$4179 ( \4556 , \4554 , \4555 );
nand \U$4180 ( \4557 , \4556 , \1915 );
nand \U$4181 ( \4558 , \4551 , \4557 );
not \U$4182 ( \4559 , \4558 );
not \U$4183 ( \4560 , \1363 );
not \U$4184 ( \4561 , RIc2271f0_9);
not \U$4185 ( \4562 , \3810 );
or \U$4186 ( \4563 , \4561 , \4562 );
not \U$4187 ( \4564 , \2670 );
nand \U$4188 ( \4565 , \4564 , \1351 );
nand \U$4189 ( \4566 , \4563 , \4565 );
not \U$4190 ( \4567 , \4566 );
or \U$4191 ( \4568 , \4560 , \4567 );
nand \U$4192 ( \4569 , \4198 , \1340 );
nand \U$4193 ( \4570 , \4568 , \4569 );
not \U$4194 ( \4571 , \4570 );
or \U$4195 ( \4572 , \4559 , \4571 );
or \U$4196 ( \4573 , \4570 , \4558 );
not \U$4197 ( \4574 , \1311 );
not \U$4198 ( \4575 , \4208 );
or \U$4199 ( \4576 , \4574 , \4575 );
not \U$4200 ( \4577 , \1308 );
not \U$4201 ( \4578 , RIc227100_11);
not \U$4202 ( \4579 , \3035 );
or \U$4203 ( \4580 , \4578 , \4579 );
nand \U$4204 ( \4581 , \2479 , \1302 );
nand \U$4205 ( \4582 , \4580 , \4581 );
nand \U$4206 ( \4583 , \4577 , \4582 );
nand \U$4207 ( \4584 , \4576 , \4583 );
nand \U$4208 ( \4585 , \4573 , \4584 );
nand \U$4209 ( \4586 , \4572 , \4585 );
not \U$4210 ( \4587 , \4586 );
not \U$4211 ( \4588 , \4587 );
or \U$4212 ( \4589 , \4548 , \4588 );
buf \U$4213 ( \4590 , \3578 );
not \U$4214 ( \4591 , \4590 );
not \U$4215 ( \4592 , \4591 );
not \U$4216 ( \4593 , \3982 );
and \U$4217 ( \4594 , \4592 , \4593 );
not \U$4218 ( \4595 , \1530 );
and \U$4219 ( \4596 , \4595 , \2190 );
nor \U$4220 ( \4597 , \4594 , \4596 );
not \U$4221 ( \4598 , \4597 );
not \U$4222 ( \4599 , \2860 );
not \U$4223 ( \4600 , \4599 );
and \U$4224 ( \4601 , \4598 , \4600 );
and \U$4225 ( \4602 , \3984 , \2173 );
nor \U$4226 ( \4603 , \4601 , \4602 );
not \U$4227 ( \4604 , \4603 );
not \U$4228 ( \4605 , \4604 );
not \U$4229 ( \4606 , \2697 );
not \U$4230 ( \4607 , RIc2267a0_31);
not \U$4231 ( \4608 , \840 );
not \U$4232 ( \4609 , \4608 );
or \U$4233 ( \4610 , \4607 , \4609 );
nand \U$4234 ( \4611 , \840 , \2072 );
nand \U$4235 ( \4612 , \4610 , \4611 );
not \U$4236 ( \4613 , \4612 );
or \U$4237 ( \4614 , \4606 , \4613 );
nand \U$4238 ( \4615 , \4028 , \3653 );
nand \U$4239 ( \4616 , \4614 , \4615 );
not \U$4240 ( \4617 , \4616 );
or \U$4241 ( \4618 , \4605 , \4617 );
not \U$4242 ( \4619 , \4616 );
not \U$4243 ( \4620 , \4619 );
not \U$4244 ( \4621 , \4603 );
or \U$4245 ( \4622 , \4620 , \4621 );
not \U$4246 ( \4623 , \1682 );
not \U$4247 ( \4624 , \3947 );
or \U$4248 ( \4625 , \4623 , \4624 );
not \U$4249 ( \4626 , RIc227010_13);
not \U$4250 ( \4627 , \2592 );
or \U$4251 ( \4628 , \4626 , \4627 );
nand \U$4252 ( \4629 , \3291 , \3841 );
nand \U$4253 ( \4630 , \4628 , \4629 );
nand \U$4254 ( \4631 , \4630 , \1680 );
nand \U$4255 ( \4632 , \4625 , \4631 );
nand \U$4256 ( \4633 , \4622 , \4632 );
nand \U$4257 ( \4634 , \4618 , \4633 );
nand \U$4258 ( \4635 , \4589 , \4634 );
nand \U$4259 ( \4636 , \4586 , \4546 );
nand \U$4260 ( \4637 , \4635 , \4636 );
and \U$4261 ( \4638 , \4511 , \4637 );
and \U$4262 ( \4639 , \4370 , \4510 );
or \U$4263 ( \4640 , \4638 , \4639 );
nand \U$4264 ( \4641 , \4368 , \4640 );
not \U$4265 ( \4642 , \4328 );
nand \U$4266 ( \4643 , \4365 , \4642 );
nand \U$4267 ( \4644 , \4641 , \4643 );
nand \U$4268 ( \4645 , \4318 , \4644 );
nand \U$4269 ( \4646 , \4317 , \4645 );
nand \U$4270 ( \4647 , \4281 , \4646 );
nand \U$4271 ( \4648 , \4278 , \4280 );
nand \U$4272 ( \4649 , \4647 , \4648 );
or \U$4273 ( \4650 , \4276 , \4649 );
nand \U$4274 ( \4651 , \4274 , \4650 );
or \U$4275 ( \4652 , \2165 , \2023 );
nand \U$4276 ( \4653 , \4652 , \2603 );
nand \U$4277 ( \4654 , \2165 , \2023 );
and \U$4278 ( \4655 , \4653 , \4654 );
or \U$4279 ( \4656 , \2924 , \2845 );
and \U$4280 ( \4657 , \4656 , \2935 );
and \U$4281 ( \4658 , \2845 , \2924 );
nor \U$4282 ( \4659 , \4657 , \4658 );
xor \U$4283 ( \4660 , \4655 , \4659 );
xor \U$4284 ( \4661 , \2859 , \2891 );
and \U$4285 ( \4662 , \4661 , \2923 );
and \U$4286 ( \4663 , \2859 , \2891 );
or \U$4287 ( \4664 , \4662 , \4663 );
not \U$4288 ( \4665 , \2850 );
xor \U$4289 ( \4666 , \3332 , \3344 );
and \U$4290 ( \4667 , \4666 , \3357 );
and \U$4291 ( \4668 , \3332 , \3344 );
or \U$4292 ( \4669 , \4667 , \4668 );
xor \U$4293 ( \4670 , \4665 , \4669 );
not \U$4294 ( \4671 , \3368 );
not \U$4295 ( \4672 , \3377 );
or \U$4296 ( \4673 , \4671 , \4672 );
or \U$4297 ( \4674 , \3377 , \3368 );
nand \U$4298 ( \4675 , \4674 , \3388 );
nand \U$4299 ( \4676 , \4673 , \4675 );
xor \U$4300 ( \4677 , \4670 , \4676 );
xor \U$4301 ( \4678 , \4664 , \4677 );
xor \U$4302 ( \4679 , \1932 , \1965 );
and \U$4303 ( \4680 , \4679 , \2022 );
and \U$4304 ( \4681 , \1932 , \1965 );
or \U$4305 ( \4682 , \4680 , \4681 );
not \U$4306 ( \4683 , \3298 );
not \U$4307 ( \4684 , \3321 );
or \U$4308 ( \4685 , \4683 , \4684 );
or \U$4309 ( \4686 , \3321 , \3298 );
not \U$4310 ( \4687 , \3309 );
nand \U$4311 ( \4688 , \4686 , \4687 );
nand \U$4312 ( \4689 , \4685 , \4688 );
xor \U$4313 ( \4690 , \4682 , \4689 );
not \U$4314 ( \4691 , \1682 );
not \U$4315 ( \4692 , RIc227010_13);
not \U$4316 ( \4693 , \2615 );
or \U$4317 ( \4694 , \4692 , \4693 );
nand \U$4318 ( \4695 , \1730 , \1758 );
nand \U$4319 ( \4696 , \4694 , \4695 );
not \U$4320 ( \4697 , \4696 );
or \U$4321 ( \4698 , \4691 , \4697 );
nand \U$4322 ( \4699 , \3384 , \1680 );
nand \U$4323 ( \4700 , \4698 , \4699 );
not \U$4324 ( \4701 , \1307 );
not \U$4325 ( \4702 , \3353 );
or \U$4326 ( \4703 , \4701 , \4702 );
not \U$4327 ( \4704 , RIc227100_11);
not \U$4328 ( \4705 , \2774 );
or \U$4329 ( \4706 , \4704 , \4705 );
nand \U$4330 ( \4707 , \2306 , \3351 );
nand \U$4331 ( \4708 , \4706 , \4707 );
nand \U$4332 ( \4709 , \4708 , \1311 );
nand \U$4333 ( \4710 , \4703 , \4709 );
xor \U$4334 ( \4711 , \4700 , \4710 );
not \U$4335 ( \4712 , \2534 );
not \U$4336 ( \4713 , RIc226d40_19);
not \U$4337 ( \4714 , \1404 );
or \U$4338 ( \4715 , \4713 , \4714 );
nand \U$4339 ( \4716 , \1228 , \2523 );
nand \U$4340 ( \4717 , \4715 , \4716 );
not \U$4341 ( \4718 , \4717 );
or \U$4342 ( \4719 , \4712 , \4718 );
nand \U$4343 ( \4720 , \3340 , \2518 );
nand \U$4344 ( \4721 , \4719 , \4720 );
xor \U$4345 ( \4722 , \4711 , \4721 );
xor \U$4346 ( \4723 , \4690 , \4722 );
xnor \U$4347 ( \4724 , \4678 , \4723 );
and \U$4348 ( \4725 , \4660 , \4724 );
and \U$4349 ( \4726 , \4655 , \4659 );
or \U$4350 ( \4727 , \4725 , \4726 );
xor \U$4351 ( \4728 , \3286 , \3390 );
and \U$4352 ( \4729 , \4728 , \3415 );
and \U$4353 ( \4730 , \3286 , \3390 );
or \U$4354 ( \4731 , \4729 , \4730 );
not \U$4355 ( \4732 , \4731 );
not \U$4356 ( \4733 , \3358 );
nand \U$4357 ( \4734 , \4733 , \3389 );
not \U$4358 ( \4735 , \3322 );
and \U$4359 ( \4736 , \4734 , \4735 );
nor \U$4360 ( \4737 , \4733 , \3389 );
nor \U$4361 ( \4738 , \4736 , \4737 );
not \U$4362 ( \4739 , \4738 );
not \U$4363 ( \4740 , \4739 );
or \U$4364 ( \4741 , \2138 , \2154 );
nand \U$4365 ( \4742 , \4741 , RIc226980_27);
not \U$4366 ( \4743 , \2860 );
not \U$4367 ( \4744 , \3364 );
or \U$4368 ( \4745 , \4743 , \4744 );
not \U$4369 ( \4746 , \931 );
not \U$4370 ( \4747 , \3982 );
and \U$4371 ( \4748 , \4746 , \4747 );
and \U$4372 ( \4749 , \931 , \2190 );
nor \U$4373 ( \4750 , \4748 , \4749 );
not \U$4374 ( \4751 , \4750 );
nand \U$4375 ( \4752 , \4751 , \2173 );
nand \U$4376 ( \4753 , \4745 , \4752 );
xor \U$4377 ( \4754 , \4742 , \4753 );
not \U$4378 ( \4755 , \2392 );
not \U$4379 ( \4756 , \3375 );
or \U$4380 ( \4757 , \4755 , \4756 );
not \U$4381 ( \4758 , RIc226c50_21);
not \U$4382 ( \4759 , \1490 );
or \U$4383 ( \4760 , \4758 , \4759 );
nand \U$4384 ( \4761 , \985 , \3204 );
nand \U$4385 ( \4762 , \4760 , \4761 );
nand \U$4386 ( \4763 , \4762 , \2367 );
nand \U$4387 ( \4764 , \4757 , \4763 );
xor \U$4388 ( \4765 , \4754 , \4764 );
and \U$4389 ( \4766 , RIc2275b0_1, \2065 );
not \U$4390 ( \4767 , \1579 );
xor \U$4391 ( \4768 , RIc2275b0_1, \3026 );
not \U$4392 ( \4769 , \4768 );
or \U$4393 ( \4770 , \4767 , \4769 );
nand \U$4394 ( \4771 , \2854 , \854 );
nand \U$4395 ( \4772 , \4770 , \4771 );
xor \U$4396 ( \4773 , \4766 , \4772 );
not \U$4397 ( \4774 , \2358 );
not \U$4398 ( \4775 , RIc226f20_15);
not \U$4399 ( \4776 , \1334 );
or \U$4400 ( \4777 , \4775 , \4776 );
not \U$4401 ( \4778 , \1949 );
nand \U$4402 ( \4779 , \4778 , \2301 );
nand \U$4403 ( \4780 , \4777 , \4779 );
not \U$4404 ( \4781 , \4780 );
or \U$4405 ( \4782 , \4774 , \4781 );
not \U$4406 ( \4783 , \3303 );
nand \U$4407 ( \4784 , \4783 , \2320 );
nand \U$4408 ( \4785 , \4782 , \4784 );
xor \U$4409 ( \4786 , \4773 , \4785 );
xor \U$4410 ( \4787 , \4765 , \4786 );
not \U$4411 ( \4788 , \954 );
not \U$4412 ( \4789 , RIc2273d0_5);
not \U$4413 ( \4790 , \2015 );
or \U$4414 ( \4791 , \4789 , \4790 );
nand \U$4415 ( \4792 , \3508 , \956 );
nand \U$4416 ( \4793 , \4791 , \4792 );
not \U$4417 ( \4794 , \4793 );
or \U$4418 ( \4795 , \4788 , \4794 );
nand \U$4419 ( \4796 , \3296 , \951 );
nand \U$4420 ( \4797 , \4795 , \4796 );
not \U$4421 ( \4798 , \1040 );
not \U$4422 ( \4799 , \3317 );
or \U$4423 ( \4800 , \4798 , \4799 );
not \U$4424 ( \4801 , RIc2274c0_3);
not \U$4425 ( \4802 , \3446 );
buf \U$4426 ( \4803 , \4802 );
not \U$4427 ( \4804 , \4803 );
or \U$4428 ( \4805 , \4801 , \4804 );
nand \U$4429 ( \4806 , \2559 , \2896 );
nand \U$4430 ( \4807 , \4805 , \4806 );
nand \U$4431 ( \4808 , \4807 , \1082 );
nand \U$4432 ( \4809 , \4800 , \4808 );
xor \U$4433 ( \4810 , \4797 , \4809 );
not \U$4434 ( \4811 , \1945 );
not \U$4435 ( \4812 , \1962 );
or \U$4436 ( \4813 , \4811 , \4812 );
not \U$4437 ( \4814 , RIc226e30_17);
not \U$4438 ( \4815 , \1393 );
or \U$4439 ( \4816 , \4814 , \4815 );
nand \U$4440 ( \4817 , \1396 , \1952 );
nand \U$4441 ( \4818 , \4816 , \4817 );
nand \U$4442 ( \4819 , \4818 , \1963 );
nand \U$4443 ( \4820 , \4813 , \4819 );
xor \U$4444 ( \4821 , \4810 , \4820 );
xor \U$4445 ( \4822 , \4787 , \4821 );
not \U$4446 ( \4823 , \4822 );
not \U$4447 ( \4824 , \4823 );
or \U$4448 ( \4825 , \4740 , \4824 );
nand \U$4449 ( \4826 , \4822 , \4738 );
nand \U$4450 ( \4827 , \4825 , \4826 );
xor \U$4451 ( \4828 , \2850 , \2851 );
and \U$4452 ( \4829 , \4828 , \2858 );
and \U$4453 ( \4830 , \2850 , \2851 );
or \U$4454 ( \4831 , \4829 , \4830 );
not \U$4455 ( \4832 , \1340 );
not \U$4456 ( \4833 , RIc2271f0_9);
not \U$4457 ( \4834 , \2834 );
or \U$4458 ( \4835 , \4833 , \4834 );
nand \U$4459 ( \4836 , \2837 , \1351 );
nand \U$4460 ( \4837 , \4835 , \4836 );
not \U$4461 ( \4838 , \4837 );
or \U$4462 ( \4839 , \4832 , \4838 );
nand \U$4463 ( \4840 , \3330 , \1597 );
nand \U$4464 ( \4841 , \4839 , \4840 );
not \U$4465 ( \4842 , \1930 );
not \U$4466 ( \4843 , RIc226b60_23);
not \U$4467 ( \4844 , \2865 );
or \U$4468 ( \4845 , \4843 , \4844 );
not \U$4469 ( \4846 , \890 );
nand \U$4470 ( \4847 , \4846 , \1927 );
nand \U$4471 ( \4848 , \4845 , \4847 );
not \U$4472 ( \4849 , \4848 );
or \U$4473 ( \4850 , \4842 , \4849 );
nand \U$4474 ( \4851 , \1929 , \1915 );
nand \U$4475 ( \4852 , \4850 , \4851 );
xor \U$4476 ( \4853 , \4841 , \4852 );
not \U$4477 ( \4854 , \1118 );
not \U$4478 ( \4855 , \1995 );
or \U$4479 ( \4856 , \4854 , \4855 );
and \U$4480 ( \4857 , \1139 , \2258 );
not \U$4481 ( \4858 , \1139 );
and \U$4482 ( \4859 , \4858 , \2261 );
nor \U$4483 ( \4860 , \4857 , \4859 );
nand \U$4484 ( \4861 , \4860 , \1121 );
nand \U$4485 ( \4862 , \4856 , \4861 );
xor \U$4486 ( \4863 , \4853 , \4862 );
xor \U$4487 ( \4864 , \4831 , \4863 );
xor \U$4488 ( \4865 , \2783 , \2806 );
and \U$4489 ( \4866 , \4865 , \2844 );
and \U$4490 ( \4867 , \2783 , \2806 );
or \U$4491 ( \4868 , \4866 , \4867 );
xor \U$4492 ( \4869 , \4864 , \4868 );
and \U$4493 ( \4870 , \4827 , \4869 );
not \U$4494 ( \4871 , \4827 );
not \U$4495 ( \4872 , \4869 );
and \U$4496 ( \4873 , \4871 , \4872 );
nor \U$4497 ( \4874 , \4870 , \4873 );
not \U$4498 ( \4875 , \4874 );
or \U$4499 ( \4876 , \4732 , \4875 );
xor \U$4500 ( \4877 , \2604 , \2755 );
and \U$4501 ( \4878 , \4877 , \2936 );
and \U$4502 ( \4879 , \2604 , \2755 );
or \U$4503 ( \4880 , \4878 , \4879 );
not \U$4504 ( \4881 , \4731 );
not \U$4505 ( \4882 , \4874 );
nand \U$4506 ( \4883 , \4881 , \4882 );
nand \U$4507 ( \4884 , \4880 , \4883 );
nand \U$4508 ( \4885 , \4876 , \4884 );
not \U$4509 ( \4886 , \4885 );
xor \U$4510 ( \4887 , \4727 , \4886 );
nand \U$4511 ( \4888 , \4872 , \4823 );
and \U$4512 ( \4889 , \4888 , \4739 );
nor \U$4513 ( \4890 , \4872 , \4823 );
nor \U$4514 ( \4891 , \4889 , \4890 );
xor \U$4515 ( \4892 , \4682 , \4689 );
and \U$4516 ( \4893 , \4892 , \4722 );
and \U$4517 ( \4894 , \4682 , \4689 );
or \U$4518 ( \4895 , \4893 , \4894 );
xor \U$4519 ( \4896 , \4766 , \4772 );
and \U$4520 ( \4897 , \4896 , \4785 );
and \U$4521 ( \4898 , \4766 , \4772 );
or \U$4522 ( \4899 , \4897 , \4898 );
and \U$4523 ( \4900 , RIc2275b0_1, \2675 );
not \U$4524 ( \4901 , \2367 );
not \U$4525 ( \4902 , RIc226c50_21);
not \U$4526 ( \4903 , \1706 );
or \U$4527 ( \4904 , \4902 , \4903 );
nand \U$4528 ( \4905 , \841 , \3204 );
nand \U$4529 ( \4906 , \4904 , \4905 );
not \U$4530 ( \4907 , \4906 );
or \U$4531 ( \4908 , \4901 , \4907 );
nand \U$4532 ( \4909 , \4762 , \2392 );
nand \U$4533 ( \4910 , \4908 , \4909 );
xor \U$4534 ( \4911 , \4900 , \4910 );
not \U$4535 ( \4912 , \854 );
not \U$4536 ( \4913 , \4768 );
or \U$4537 ( \4914 , \4912 , \4913 );
xor \U$4538 ( \4915 , RIc2275b0_1, \2480 );
nand \U$4539 ( \4916 , \4915 , \1579 );
nand \U$4540 ( \4917 , \4914 , \4916 );
xor \U$4541 ( \4918 , \4911 , \4917 );
xor \U$4542 ( \4919 , \4899 , \4918 );
not \U$4543 ( \4920 , \2534 );
and \U$4544 ( \4921 , \1456 , RIc226d40_19);
not \U$4545 ( \4922 , \1456 );
and \U$4546 ( \4923 , \4922 , \3338 );
or \U$4547 ( \4924 , \4921 , \4923 );
not \U$4548 ( \4925 , \4924 );
or \U$4549 ( \4926 , \4920 , \4925 );
nand \U$4550 ( \4927 , \4717 , \2518 );
nand \U$4551 ( \4928 , \4926 , \4927 );
not \U$4552 ( \4929 , \1915 );
not \U$4553 ( \4930 , \4848 );
or \U$4554 ( \4931 , \4929 , \4930 );
not \U$4555 ( \4932 , RIc226b60_23);
not \U$4556 ( \4933 , \1074 );
or \U$4557 ( \4934 , \4932 , \4933 );
nand \U$4558 ( \4935 , \1073 , \2111 );
nand \U$4559 ( \4936 , \4934 , \4935 );
nand \U$4560 ( \4937 , \4936 , \1930 );
nand \U$4561 ( \4938 , \4931 , \4937 );
xor \U$4562 ( \4939 , \4928 , \4938 );
not \U$4563 ( \4940 , \1311 );
and \U$4564 ( \4941 , \2348 , RIc227100_11);
not \U$4565 ( \4942 , \2348 );
and \U$4566 ( \4943 , \4942 , \3351 );
nor \U$4567 ( \4944 , \4941 , \4943 );
not \U$4568 ( \4945 , \4944 );
or \U$4569 ( \4946 , \4940 , \4945 );
nand \U$4570 ( \4947 , \4708 , \1307 );
nand \U$4571 ( \4948 , \4946 , \4947 );
xor \U$4572 ( \4949 , \4939 , \4948 );
xor \U$4573 ( \4950 , \4919 , \4949 );
xor \U$4574 ( \4951 , \4895 , \4950 );
not \U$4575 ( \4952 , \2320 );
not \U$4576 ( \4953 , \4780 );
or \U$4577 ( \4954 , \4952 , \4953 );
not \U$4578 ( \4955 , RIc226f20_15);
not \U$4579 ( \4956 , \1602 );
or \U$4580 ( \4957 , \4955 , \4956 );
nand \U$4581 ( \4958 , \1533 , \2351 );
nand \U$4582 ( \4959 , \4957 , \4958 );
nand \U$4583 ( \4960 , \4959 , \2358 );
nand \U$4584 ( \4961 , \4954 , \4960 );
not \U$4585 ( \4962 , \1082 );
and \U$4586 ( \4963 , \2593 , \1032 );
not \U$4587 ( \4964 , \2593 );
and \U$4588 ( \4965 , \4964 , RIc2274c0_3);
or \U$4589 ( \4966 , \4963 , \4965 );
not \U$4590 ( \4967 , \4966 );
or \U$4591 ( \4968 , \4962 , \4967 );
nand \U$4592 ( \4969 , \4807 , \1040 );
nand \U$4593 ( \4970 , \4968 , \4969 );
xor \U$4594 ( \4971 , \4961 , \4970 );
not \U$4595 ( \4972 , \951 );
not \U$4596 ( \4973 , \4793 );
or \U$4597 ( \4974 , \4972 , \4973 );
not \U$4598 ( \4975 , RIc2273d0_5);
not \U$4599 ( \4976 , \1990 );
or \U$4600 ( \4977 , \4975 , \4976 );
nand \U$4601 ( \4978 , \1991 , \946 );
nand \U$4602 ( \4979 , \4977 , \4978 );
nand \U$4603 ( \4980 , \4979 , \954 );
nand \U$4604 ( \4981 , \4974 , \4980 );
xor \U$4605 ( \4982 , \4971 , \4981 );
not \U$4606 ( \4983 , \1963 );
not \U$4607 ( \4984 , RIc226e30_17);
not \U$4608 ( \4985 , \1441 );
or \U$4609 ( \4986 , \4984 , \4985 );
nand \U$4610 ( \4987 , \3242 , \1960 );
nand \U$4611 ( \4988 , \4986 , \4987 );
not \U$4612 ( \4989 , \4988 );
or \U$4613 ( \4990 , \4983 , \4989 );
nand \U$4614 ( \4991 , \4818 , \1945 );
nand \U$4615 ( \4992 , \4990 , \4991 );
not \U$4616 ( \4993 , \1340 );
not \U$4617 ( \4994 , RIc2271f0_9);
not \U$4618 ( \4995 , \2424 );
or \U$4619 ( \4996 , \4994 , \4995 );
nand \U$4620 ( \4997 , \2423 , \1342 );
nand \U$4621 ( \4998 , \4996 , \4997 );
not \U$4622 ( \4999 , \4998 );
or \U$4623 ( \5000 , \4993 , \4999 );
nand \U$4624 ( \5001 , \4837 , \1363 );
nand \U$4625 ( \5002 , \5000 , \5001 );
xor \U$4626 ( \5003 , \4992 , \5002 );
not \U$4627 ( \5004 , \1118 );
not \U$4628 ( \5005 , \4860 );
or \U$4629 ( \5006 , \5004 , \5005 );
and \U$4630 ( \5007 , RIc2272e0_7, \2235 );
not \U$4631 ( \5008 , RIc2272e0_7);
and \U$4632 ( \5009 , \5008 , \2230 );
nor \U$4633 ( \5010 , \5007 , \5009 );
nand \U$4634 ( \5011 , \5010 , \1121 );
nand \U$4635 ( \5012 , \5006 , \5011 );
xor \U$4636 ( \5013 , \5003 , \5012 );
xor \U$4637 ( \5014 , \4982 , \5013 );
xor \U$4638 ( \5015 , \4665 , \4669 );
and \U$4639 ( \5016 , \5015 , \4676 );
and \U$4640 ( \5017 , \4665 , \4669 );
or \U$4641 ( \5018 , \5016 , \5017 );
xor \U$4642 ( \5019 , \5014 , \5018 );
xor \U$4643 ( \5020 , \4951 , \5019 );
xor \U$4644 ( \5021 , \4891 , \5020 );
xor \U$4645 ( \5022 , \4831 , \4863 );
and \U$4646 ( \5023 , \5022 , \4868 );
and \U$4647 ( \5024 , \4831 , \4863 );
or \U$4648 ( \5025 , \5023 , \5024 );
not \U$4649 ( \5026 , \4677 );
not \U$4650 ( \5027 , \4723 );
or \U$4651 ( \5028 , \5026 , \5027 );
or \U$4652 ( \5029 , \4723 , \4677 );
nand \U$4653 ( \5030 , \5029 , \4664 );
nand \U$4654 ( \5031 , \5028 , \5030 );
xor \U$4655 ( \5032 , \5025 , \5031 );
not \U$4656 ( \5033 , \2195 );
or \U$4657 ( \5034 , \4750 , \5033 );
not \U$4658 ( \5035 , \2173 );
or \U$4659 ( \5036 , \5035 , \3982 );
nand \U$4660 ( \5037 , \5034 , \5036 );
not \U$4661 ( \5038 , \5037 );
not \U$4662 ( \5039 , \4696 );
or \U$4663 ( \5040 , \5039 , \1679 );
not \U$4664 ( \5041 , RIc227010_13);
not \U$4665 ( \5042 , \3044 );
or \U$4666 ( \5043 , \5041 , \5042 );
nand \U$4667 ( \5044 , \3299 , \1296 );
nand \U$4668 ( \5045 , \5043 , \5044 );
not \U$4669 ( \5046 , \5045 );
or \U$4670 ( \5047 , \5046 , \1757 );
nand \U$4671 ( \5048 , \5040 , \5047 );
xor \U$4672 ( \5049 , \5038 , \5048 );
xor \U$4673 ( \5050 , \4797 , \4809 );
and \U$4674 ( \5051 , \5050 , \4820 );
and \U$4675 ( \5052 , \4797 , \4809 );
or \U$4676 ( \5053 , \5051 , \5052 );
xor \U$4677 ( \5054 , \5049 , \5053 );
not \U$4678 ( \5055 , \4700 );
not \U$4679 ( \5056 , \4710 );
or \U$4680 ( \5057 , \5055 , \5056 );
or \U$4681 ( \5058 , \4710 , \4700 );
nand \U$4682 ( \5059 , \5058 , \4721 );
nand \U$4683 ( \5060 , \5057 , \5059 );
xor \U$4684 ( \5061 , \4742 , \4753 );
and \U$4685 ( \5062 , \5061 , \4764 );
and \U$4686 ( \5063 , \4742 , \4753 );
or \U$4687 ( \5064 , \5062 , \5063 );
xor \U$4688 ( \5065 , \5060 , \5064 );
xor \U$4689 ( \5066 , \4841 , \4852 );
and \U$4690 ( \5067 , \5066 , \4862 );
and \U$4691 ( \5068 , \4841 , \4852 );
or \U$4692 ( \5069 , \5067 , \5068 );
xor \U$4693 ( \5070 , \5065 , \5069 );
xor \U$4694 ( \5071 , \5054 , \5070 );
xor \U$4695 ( \5072 , \4765 , \4786 );
and \U$4696 ( \5073 , \5072 , \4821 );
and \U$4697 ( \5074 , \4765 , \4786 );
or \U$4698 ( \5075 , \5073 , \5074 );
xor \U$4699 ( \5076 , \5071 , \5075 );
xor \U$4700 ( \5077 , \5032 , \5076 );
xor \U$4701 ( \5078 , \5021 , \5077 );
xor \U$4702 ( \5079 , \4887 , \5078 );
xor \U$4703 ( \5080 , \4655 , \4659 );
xor \U$4704 ( \5081 , \5080 , \4724 );
xor \U$4705 ( \5082 , \3282 , \3416 );
and \U$4706 ( \5083 , \5082 , \3551 );
and \U$4707 ( \5084 , \3282 , \3416 );
or \U$4708 ( \5085 , \5083 , \5084 );
not \U$4709 ( \5086 , \5085 );
xor \U$4710 ( \5087 , \5081 , \5086 );
not \U$4711 ( \5088 , \4880 );
and \U$4712 ( \5089 , \4731 , \4882 );
not \U$4713 ( \5090 , \4731 );
and \U$4714 ( \5091 , \5090 , \4874 );
nor \U$4715 ( \5092 , \5089 , \5091 );
not \U$4716 ( \5093 , \5092 );
and \U$4717 ( \5094 , \5088 , \5093 );
and \U$4718 ( \5095 , \4880 , \5092 );
nor \U$4719 ( \5096 , \5094 , \5095 );
and \U$4720 ( \5097 , \5087 , \5096 );
and \U$4721 ( \5098 , \5081 , \5086 );
or \U$4722 ( \5099 , \5097 , \5098 );
nand \U$4723 ( \5100 , \5079 , \5099 );
xor \U$4724 ( \5101 , \5081 , \5086 );
xor \U$4725 ( \5102 , \5101 , \5096 );
or \U$4726 ( \5103 , \3552 , \2937 );
and \U$4727 ( \5104 , \5103 , \3887 );
and \U$4728 ( \5105 , \2937 , \3552 );
nor \U$4729 ( \5106 , \5104 , \5105 );
nand \U$4730 ( \5107 , \5102 , \5106 );
nand \U$4731 ( \5108 , \5100 , \5107 );
nor \U$4732 ( \5109 , \4651 , \5108 );
not \U$4733 ( \5110 , \5109 );
xor \U$4734 ( \5111 , \4166 , \4169 );
not \U$4735 ( \5112 , \4264 );
xor \U$4736 ( \5113 , \5111 , \5112 );
xor \U$4737 ( \5114 , \4315 , \4644 );
xnor \U$4738 ( \5115 , \5114 , \4312 );
xor \U$4739 ( \5116 , \5113 , \5115 );
not \U$4740 ( \5117 , \4642 );
not \U$4741 ( \5118 , \4640 );
not \U$4742 ( \5119 , \5118 );
or \U$4743 ( \5120 , \5117 , \5119 );
nand \U$4744 ( \5121 , \4640 , \4328 );
nand \U$4745 ( \5122 , \5120 , \5121 );
and \U$4746 ( \5123 , \5122 , \4366 );
not \U$4747 ( \5124 , \5122 );
and \U$4748 ( \5125 , \5124 , \4365 );
nor \U$4749 ( \5126 , \5123 , \5125 );
not \U$4750 ( \5127 , \4381 );
not \U$4751 ( \5128 , RIc2265c0_35);
not \U$4752 ( \5129 , \932 );
or \U$4753 ( \5130 , \5128 , \5129 );
nand \U$4754 ( \5131 , \2704 , \3620 );
nand \U$4755 ( \5132 , \5130 , \5131 );
not \U$4756 ( \5133 , \5132 );
or \U$4757 ( \5134 , \5127 , \5133 );
buf \U$4758 ( \5135 , \4382 );
nand \U$4759 ( \5136 , \5135 , RIc2265c0_35);
nand \U$4760 ( \5137 , \5134 , \5136 );
xor \U$4761 ( \5138 , \4385 , \4408 );
xor \U$4762 ( \5139 , \5138 , \4422 );
xor \U$4763 ( \5140 , \5137 , \5139 );
not \U$4764 ( \5141 , \1121 );
not \U$4765 ( \5142 , \4243 );
or \U$4766 ( \5143 , \5141 , \5142 );
not \U$4767 ( \5144 , RIc2272e0_7);
not \U$4768 ( \5145 , \2043 );
or \U$4769 ( \5146 , \5144 , \5145 );
nand \U$4770 ( \5147 , \3800 , \1139 );
nand \U$4771 ( \5148 , \5146 , \5147 );
nand \U$4772 ( \5149 , \1118 , \5148 );
nand \U$4773 ( \5150 , \5143 , \5149 );
and \U$4774 ( \5151 , \5140 , \5150 );
and \U$4775 ( \5152 , \5137 , \5139 );
or \U$4776 ( \5153 , \5151 , \5152 );
not \U$4777 ( \5154 , \954 );
not \U$4778 ( \5155 , \4503 );
or \U$4779 ( \5156 , \5154 , \5155 );
not \U$4780 ( \5157 , RIc2273d0_5);
not \U$4781 ( \5158 , \3121 );
or \U$4782 ( \5159 , \5157 , \5158 );
not \U$4783 ( \5160 , \3119 );
nand \U$4784 ( \5161 , \5160 , \956 );
nand \U$4785 ( \5162 , \5159 , \5161 );
nand \U$4786 ( \5163 , \5162 , \951 );
nand \U$4787 ( \5164 , \5156 , \5163 );
not \U$4788 ( \5165 , \5164 );
not \U$4789 ( \5166 , \1082 );
not \U$4790 ( \5167 , \4486 );
or \U$4791 ( \5168 , \5166 , \5167 );
not \U$4792 ( \5169 , RIc2274c0_3);
not \U$4793 ( \5170 , \4046 );
or \U$4794 ( \5171 , \5169 , \5170 );
nand \U$4795 ( \5172 , \4050 , \1078 );
nand \U$4796 ( \5173 , \5171 , \5172 );
nand \U$4797 ( \5174 , \5173 , \1040 );
nand \U$4798 ( \5175 , \5168 , \5174 );
not \U$4799 ( \5176 , \5175 );
or \U$4800 ( \5177 , \5165 , \5176 );
or \U$4801 ( \5178 , \5175 , \5164 );
not \U$4802 ( \5179 , RIc2266b0_33);
and \U$4803 ( \5180 , \5179 , \889 );
not \U$4804 ( \5181 , \5179 );
and \U$4805 ( \5182 , \5181 , \890 );
nor \U$4806 ( \5183 , \5180 , \5182 );
not \U$4807 ( \5184 , \5183 );
not \U$4808 ( \5185 , \3629 );
not \U$4809 ( \5186 , \5185 );
and \U$4810 ( \5187 , \5184 , \5186 );
and \U$4811 ( \5188 , \4446 , \3631 );
nor \U$4812 ( \5189 , \5187 , \5188 );
not \U$4813 ( \5190 , \5189 );
nand \U$4814 ( \5191 , \5178 , \5190 );
nand \U$4815 ( \5192 , \5177 , \5191 );
not \U$4816 ( \5193 , \5192 );
nor \U$4817 ( \5194 , \4386 , \554 );
not \U$4818 ( \5195 , \5194 );
not \U$4819 ( \5196 , \4111 );
or \U$4820 ( \5197 , \5195 , \5196 );
not \U$4821 ( \5198 , \554 );
and \U$4822 ( \5199 , \4072 , \5198 );
not \U$4823 ( \5200 , \657 );
nor \U$4824 ( \5201 , \5199 , \5200 );
nand \U$4825 ( \5202 , \5197 , \5201 );
not \U$4826 ( \5203 , \5202 );
nand \U$4827 ( \5204 , \685 , \5198 );
nor \U$4828 ( \5205 , \4087 , \5204 );
nand \U$4829 ( \5206 , \4084 , \5205 );
nand \U$4830 ( \5207 , \5203 , \5206 );
not \U$4831 ( \5208 , \659 );
nor \U$4832 ( \5209 , \5208 , \553 );
and \U$4833 ( \5210 , \5207 , \5209 );
not \U$4834 ( \5211 , \5207 );
not \U$4835 ( \5212 , \5209 );
and \U$4836 ( \5213 , \5211 , \5212 );
nor \U$4837 ( \5214 , \5210 , \5213 );
buf \U$4838 ( \5215 , \5214 );
not \U$4839 ( \5216 , \5215 );
not \U$4840 ( \5217 , \5216 );
and \U$4841 ( \5218 , \5217 , RIc2275b0_1);
not \U$4842 ( \5219 , \1579 );
not \U$4843 ( \5220 , \4420 );
or \U$4844 ( \5221 , \5219 , \5220 );
xor \U$4845 ( \5222 , RIc2275b0_1, \4407 );
nand \U$4846 ( \5223 , \5222 , \854 );
nand \U$4847 ( \5224 , \5221 , \5223 );
xor \U$4848 ( \5225 , \5218 , \5224 );
not \U$4849 ( \5226 , \2367 );
not \U$4850 ( \5227 , \4477 );
or \U$4851 ( \5228 , \5226 , \5227 );
not \U$4852 ( \5229 , RIc226c50_21);
not \U$4853 ( \5230 , \3093 );
or \U$4854 ( \5231 , \5229 , \5230 );
nand \U$4855 ( \5232 , \2305 , \2383 );
nand \U$4856 ( \5233 , \5231 , \5232 );
nand \U$4857 ( \5234 , \5233 , \2392 );
nand \U$4858 ( \5235 , \5228 , \5234 );
and \U$4859 ( \5236 , \5225 , \5235 );
and \U$4860 ( \5237 , \5218 , \5224 );
or \U$4861 ( \5238 , \5236 , \5237 );
not \U$4862 ( \5239 , \5238 );
not \U$4863 ( \5240 , \2154 );
not \U$4864 ( \5241 , \4530 );
or \U$4865 ( \5242 , \5240 , \5241 );
not \U$4866 ( \5243 , RIc226980_27);
not \U$4867 ( \5244 , \3497 );
or \U$4868 ( \5245 , \5243 , \5244 );
not \U$4869 ( \5246 , \3496 );
buf \U$4870 ( \5247 , \5246 );
nand \U$4871 ( \5248 , \5247 , \2150 );
nand \U$4872 ( \5249 , \5245 , \5248 );
nand \U$4873 ( \5250 , \5249 , \2138 );
nand \U$4874 ( \5251 , \5242 , \5250 );
not \U$4875 ( \5252 , \5251 );
not \U$4876 ( \5253 , \2078 );
and \U$4877 ( \5254 , RIc226890_29, \1402 );
not \U$4878 ( \5255 , RIc226890_29);
and \U$4879 ( \5256 , \5255 , \3994 );
or \U$4880 ( \5257 , \5254 , \5256 );
not \U$4881 ( \5258 , \5257 );
or \U$4882 ( \5259 , \5253 , \5258 );
nand \U$4883 ( \5260 , \4434 , \2086 );
nand \U$4884 ( \5261 , \5259 , \5260 );
not \U$4885 ( \5262 , \5261 );
or \U$4886 ( \5263 , \5252 , \5262 );
or \U$4887 ( \5264 , \5251 , \5261 );
not \U$4888 ( \5265 , \2534 );
not \U$4889 ( \5266 , \4459 );
or \U$4890 ( \5267 , \5265 , \5266 );
not \U$4891 ( \5268 , RIc226d40_19);
buf \U$4892 ( \5269 , \2443 );
not \U$4893 ( \5270 , \5269 );
not \U$4894 ( \5271 , \5270 );
or \U$4895 ( \5272 , \5268 , \5271 );
nand \U$4896 ( \5273 , \4037 , \1941 );
nand \U$4897 ( \5274 , \5272 , \5273 );
nand \U$4898 ( \5275 , \5274 , \2518 );
nand \U$4899 ( \5276 , \5267 , \5275 );
nand \U$4900 ( \5277 , \5264 , \5276 );
nand \U$4901 ( \5278 , \5263 , \5277 );
not \U$4902 ( \5279 , \5278 );
nand \U$4903 ( \5280 , \5239 , \5279 );
not \U$4904 ( \5281 , \5280 );
or \U$4905 ( \5282 , \5193 , \5281 );
nand \U$4906 ( \5283 , \5238 , \5278 );
nand \U$4907 ( \5284 , \5282 , \5283 );
xor \U$4908 ( \5285 , \5153 , \5284 );
not \U$4909 ( \5286 , \1963 );
not \U$4910 ( \5287 , \4539 );
or \U$4911 ( \5288 , \5286 , \5287 );
and \U$4912 ( \5289 , \2258 , RIc226e30_17);
not \U$4913 ( \5290 , \2258 );
and \U$4914 ( \5291 , \5290 , \1960 );
or \U$4915 ( \5292 , \5289 , \5291 );
nand \U$4916 ( \5293 , \5292 , \1945 );
nand \U$4917 ( \5294 , \5288 , \5293 );
not \U$4918 ( \5295 , \2711 );
not \U$4919 ( \5296 , \4612 );
or \U$4920 ( \5297 , \5295 , \5296 );
not \U$4921 ( \5298 , RIc2267a0_31);
not \U$4922 ( \5299 , \1558 );
or \U$4923 ( \5300 , \5298 , \5299 );
not \U$4924 ( \5301 , \1558 );
nand \U$4925 ( \5302 , \5301 , \2705 );
nand \U$4926 ( \5303 , \5300 , \5302 );
nand \U$4927 ( \5304 , \5303 , \2697 );
nand \U$4928 ( \5305 , \5297 , \5304 );
or \U$4929 ( \5306 , \5294 , \5305 );
not \U$4930 ( \5307 , \2320 );
not \U$4931 ( \5308 , RIc226f20_15);
not \U$4932 ( \5309 , \3509 );
or \U$4933 ( \5310 , \5308 , \5309 );
nand \U$4934 ( \5311 , \3508 , \2301 );
nand \U$4935 ( \5312 , \5310 , \5311 );
not \U$4936 ( \5313 , \5312 );
or \U$4937 ( \5314 , \5307 , \5313 );
nand \U$4938 ( \5315 , \4519 , \2358 );
nand \U$4939 ( \5316 , \5314 , \5315 );
nand \U$4940 ( \5317 , \5306 , \5316 );
nand \U$4941 ( \5318 , \5294 , \5305 );
nand \U$4942 ( \5319 , \5317 , \5318 );
not \U$4943 ( \5320 , \1680 );
not \U$4944 ( \5321 , RIc227010_13);
not \U$4945 ( \5322 , \3447 );
or \U$4946 ( \5323 , \5321 , \5322 );
not \U$4947 ( \5324 , \2556 );
nand \U$4948 ( \5325 , \5324 , \1758 );
nand \U$4949 ( \5326 , \5323 , \5325 );
not \U$4950 ( \5327 , \5326 );
or \U$4951 ( \5328 , \5320 , \5327 );
nand \U$4952 ( \5329 , \4630 , \1682 );
nand \U$4953 ( \5330 , \5328 , \5329 );
not \U$4954 ( \5331 , RIc226a70_25);
not \U$4955 ( \5332 , \1333 );
or \U$4956 ( \5333 , \5331 , \5332 );
nand \U$4957 ( \5334 , \3439 , \1905 );
nand \U$4958 ( \5335 , \5333 , \5334 );
not \U$4959 ( \5336 , \5335 );
not \U$4960 ( \5337 , \2860 );
or \U$4961 ( \5338 , \5336 , \5337 );
not \U$4962 ( \5339 , \4597 );
nand \U$4963 ( \5340 , \5339 , \2173 );
nand \U$4964 ( \5341 , \5338 , \5340 );
or \U$4965 ( \5342 , \5330 , \5341 );
not \U$4966 ( \5343 , \1311 );
not \U$4967 ( \5344 , \4582 );
or \U$4968 ( \5345 , \5343 , \5344 );
not \U$4969 ( \5346 , RIc227100_11);
not \U$4970 ( \5347 , \3023 );
or \U$4971 ( \5348 , \5346 , \5347 );
nand \U$4972 ( \5349 , \2895 , \1302 );
nand \U$4973 ( \5350 , \5348 , \5349 );
nand \U$4974 ( \5351 , \5350 , \1307 );
nand \U$4975 ( \5352 , \5345 , \5351 );
nand \U$4976 ( \5353 , \5342 , \5352 );
nand \U$4977 ( \5354 , \5330 , \5341 );
nand \U$4978 ( \5355 , \5353 , \5354 );
or \U$4979 ( \5356 , \5319 , \5355 );
not \U$4980 ( \5357 , \1915 );
not \U$4981 ( \5358 , RIc226b60_23);
not \U$4982 ( \5359 , \4178 );
or \U$4983 ( \5360 , \5358 , \5359 );
nand \U$4984 ( \5361 , \1730 , \2111 );
nand \U$4985 ( \5362 , \5360 , \5361 );
not \U$4986 ( \5363 , \5362 );
or \U$4987 ( \5364 , \5357 , \5363 );
buf \U$4988 ( \5365 , \1930 );
nand \U$4989 ( \5366 , \4556 , \5365 );
nand \U$4990 ( \5367 , \5364 , \5366 );
not \U$4991 ( \5368 , \5367 );
not \U$4992 ( \5369 , \1340 );
not \U$4993 ( \5370 , \4566 );
or \U$4994 ( \5371 , \5369 , \5370 );
not \U$4995 ( \5372 , RIc2271f0_9);
not \U$4996 ( \5373 , \3010 );
or \U$4997 ( \5374 , \5372 , \5373 );
nand \U$4998 ( \5375 , \2065 , \1342 );
nand \U$4999 ( \5376 , \5374 , \5375 );
nand \U$5000 ( \5377 , \5376 , \1363 );
nand \U$5001 ( \5378 , \5371 , \5377 );
not \U$5002 ( \5379 , \5378 );
or \U$5003 ( \5380 , \5368 , \5379 );
or \U$5004 ( \5381 , \5378 , \5367 );
not \U$5005 ( \5382 , \1118 );
not \U$5006 ( \5383 , RIc2272e0_7);
not \U$5007 ( \5384 , \4228 );
or \U$5008 ( \5385 , \5383 , \5384 );
not \U$5009 ( \5386 , \4228 );
nand \U$5010 ( \5387 , \5386 , \940 );
nand \U$5011 ( \5388 , \5385 , \5387 );
not \U$5012 ( \5389 , \5388 );
or \U$5013 ( \5390 , \5382 , \5389 );
nand \U$5014 ( \5391 , \5148 , \1121 );
nand \U$5015 ( \5392 , \5390 , \5391 );
nand \U$5016 ( \5393 , \5381 , \5392 );
nand \U$5017 ( \5394 , \5380 , \5393 );
nand \U$5018 ( \5395 , \5356 , \5394 );
not \U$5019 ( \5396 , \5355 );
not \U$5020 ( \5397 , \5396 );
and \U$5021 ( \5398 , \5317 , \5318 );
not \U$5022 ( \5399 , \5398 );
nand \U$5023 ( \5400 , \5397 , \5399 );
nand \U$5024 ( \5401 , \5395 , \5400 );
and \U$5025 ( \5402 , \5285 , \5401 );
and \U$5026 ( \5403 , \5153 , \5284 );
or \U$5027 ( \5404 , \5402 , \5403 );
xor \U$5028 ( \5405 , \4370 , \4510 );
xor \U$5029 ( \5406 , \5405 , \4637 );
xor \U$5030 ( \5407 , \5404 , \5406 );
xor \U$5031 ( \5408 , \4425 , \4465 );
xor \U$5032 ( \5409 , \5408 , \4507 );
buf \U$5033 ( \5410 , \5409 );
not \U$5034 ( \5411 , \4587 );
not \U$5035 ( \5412 , \4634 );
or \U$5036 ( \5413 , \5411 , \5412 );
or \U$5037 ( \5414 , \4587 , \4634 );
nand \U$5038 ( \5415 , \5413 , \5414 );
and \U$5039 ( \5416 , \5415 , \4546 );
not \U$5040 ( \5417 , \5415 );
and \U$5041 ( \5418 , \5417 , \4547 );
nor \U$5042 ( \5419 , \5416 , \5418 );
or \U$5043 ( \5420 , \5410 , \5419 );
xor \U$5044 ( \5421 , \4490 , \4479 );
xor \U$5045 ( \5422 , \5421 , \4505 );
not \U$5046 ( \5423 , \5422 );
and \U$5047 ( \5424 , \4436 , \4449 );
not \U$5048 ( \5425 , \4436 );
and \U$5049 ( \5426 , \5425 , \4448 );
nor \U$5050 ( \5427 , \5424 , \5426 );
xor \U$5051 ( \5428 , \5427 , \4463 );
buf \U$5052 ( \5429 , \5428 );
not \U$5053 ( \5430 , \5429 );
or \U$5054 ( \5431 , \5423 , \5430 );
or \U$5055 ( \5432 , \5429 , \5422 );
xor \U$5056 ( \5433 , \4584 , \4570 );
xor \U$5057 ( \5434 , \5433 , \4558 );
nand \U$5058 ( \5435 , \5432 , \5434 );
nand \U$5059 ( \5436 , \5431 , \5435 );
nand \U$5060 ( \5437 , \5420 , \5436 );
nand \U$5061 ( \5438 , \5419 , \5410 );
nand \U$5062 ( \5439 , \5437 , \5438 );
and \U$5063 ( \5440 , \5407 , \5439 );
and \U$5064 ( \5441 , \5404 , \5406 );
or \U$5065 ( \5442 , \5440 , \5441 );
not \U$5066 ( \5443 , \5442 );
xor \U$5067 ( \5444 , \5126 , \5443 );
xor \U$5068 ( \5445 , \4309 , \4283 );
xor \U$5069 ( \5446 , \5445 , \4287 );
and \U$5070 ( \5447 , \5444 , \5446 );
and \U$5071 ( \5448 , \5126 , \5443 );
or \U$5072 ( \5449 , \5447 , \5448 );
xor \U$5073 ( \5450 , \5116 , \5449 );
xor \U$5074 ( \5451 , \4331 , \4359 );
xor \U$5075 ( \5452 , \5451 , \4362 );
not \U$5076 ( \5453 , \5452 );
not \U$5077 ( \5454 , \5453 );
xor \U$5078 ( \5455 , \4292 , \4302 );
xor \U$5079 ( \5456 , \5455 , \4306 );
not \U$5080 ( \5457 , \5456 );
or \U$5081 ( \5458 , \5454 , \5457 );
xor \U$5082 ( \5459 , \4521 , \4532 );
xor \U$5083 ( \5460 , \5459 , \4543 );
and \U$5084 ( \5461 , \4632 , \4619 );
not \U$5085 ( \5462 , \4632 );
and \U$5086 ( \5463 , \5462 , \4616 );
or \U$5087 ( \5464 , \5461 , \5463 );
not \U$5088 ( \5465 , \4604 );
and \U$5089 ( \5466 , \5464 , \5465 );
not \U$5090 ( \5467 , \5464 );
and \U$5091 ( \5468 , \5467 , \4604 );
nor \U$5092 ( \5469 , \5466 , \5468 );
not \U$5093 ( \5470 , \5469 );
or \U$5094 ( \5471 , \5460 , \5470 );
xor \U$5095 ( \5472 , \5137 , \5139 );
xor \U$5096 ( \5473 , \5472 , \5150 );
nand \U$5097 ( \5474 , \5471 , \5473 );
nand \U$5098 ( \5475 , \5470 , \5460 );
nand \U$5099 ( \5476 , \5474 , \5475 );
xor \U$5100 ( \5477 , \4294 , \4296 );
xor \U$5101 ( \5478 , \5477 , \4299 );
xor \U$5102 ( \5479 , \5476 , \5478 );
xnor \U$5103 ( \5480 , \4350 , \4354 );
and \U$5104 ( \5481 , \5480 , \4357 );
not \U$5105 ( \5482 , \5480 );
and \U$5106 ( \5483 , \5482 , \4340 );
nor \U$5107 ( \5484 , \5481 , \5483 );
and \U$5108 ( \5485 , \5479 , \5484 );
and \U$5109 ( \5486 , \5476 , \5478 );
or \U$5110 ( \5487 , \5485 , \5486 );
nand \U$5111 ( \5488 , \5458 , \5487 );
not \U$5112 ( \5489 , \5456 );
nand \U$5113 ( \5490 , \5489 , \5452 );
and \U$5114 ( \5491 , \5488 , \5490 );
xor \U$5115 ( \5492 , \5404 , \5406 );
xor \U$5116 ( \5493 , \5492 , \5439 );
not \U$5117 ( \5494 , \5493 );
not \U$5118 ( \5495 , \5494 );
and \U$5119 ( \5496 , RIc226458_38, RIc2263e0_39);
not \U$5120 ( \5497 , RIc226458_38);
not \U$5121 ( \5498 , RIc2263e0_39);
and \U$5122 ( \5499 , \5497 , \5498 );
nor \U$5123 ( \5500 , \5496 , \5499 );
not \U$5124 ( \5501 , \5500 );
and \U$5125 ( \5502 , RIc226458_38, RIc2264d0_37);
not \U$5126 ( \5503 , RIc226458_38);
not \U$5127 ( \5504 , RIc2264d0_37);
and \U$5128 ( \5505 , \5503 , \5504 );
nor \U$5129 ( \5506 , \5502 , \5505 );
nand \U$5130 ( \5507 , \5501 , \5506 );
not \U$5131 ( \5508 , \5507 );
buf \U$5132 ( \5509 , \5508 );
not \U$5133 ( \5510 , \5509 );
not \U$5134 ( \5511 , RIc2264d0_37);
not \U$5135 ( \5512 , \932 );
or \U$5136 ( \5513 , \5511 , \5512 );
not \U$5137 ( \5514 , RIc2264d0_37);
nand \U$5138 ( \5515 , \2704 , \5514 );
nand \U$5139 ( \5516 , \5513 , \5515 );
not \U$5140 ( \5517 , \5516 );
or \U$5141 ( \5518 , \5510 , \5517 );
buf \U$5142 ( \5519 , \5500 );
nand \U$5143 ( \5520 , \5519 , RIc2264d0_37);
nand \U$5144 ( \5521 , \5518 , \5520 );
not \U$5145 ( \5522 , \1597 );
not \U$5146 ( \5523 , RIc2271f0_9);
not \U$5147 ( \5524 , \2731 );
or \U$5148 ( \5525 , \5523 , \5524 );
not \U$5149 ( \5526 , \2042 );
buf \U$5150 ( \5527 , \5526 );
not \U$5151 ( \5528 , \5527 );
nand \U$5152 ( \5529 , \5528 , \1342 );
nand \U$5153 ( \5530 , \5525 , \5529 );
not \U$5154 ( \5531 , \5530 );
or \U$5155 ( \5532 , \5522 , \5531 );
nand \U$5156 ( \5533 , \1340 , \5376 );
nand \U$5157 ( \5534 , \5532 , \5533 );
xor \U$5158 ( \5535 , \5521 , \5534 );
not \U$5159 ( \5536 , \1307 );
not \U$5160 ( \5537 , RIc227100_11);
not \U$5161 ( \5538 , \2672 );
or \U$5162 ( \5539 , \5537 , \5538 );
nand \U$5163 ( \5540 , \2720 , \1291 );
nand \U$5164 ( \5541 , \5539 , \5540 );
not \U$5165 ( \5542 , \5541 );
or \U$5166 ( \5543 , \5536 , \5542 );
nand \U$5167 ( \5544 , \5350 , \1311 );
nand \U$5168 ( \5545 , \5543 , \5544 );
and \U$5169 ( \5546 , \5535 , \5545 );
and \U$5170 ( \5547 , \5521 , \5534 );
or \U$5171 ( \5548 , \5546 , \5547 );
not \U$5172 ( \5549 , \5548 );
xor \U$5173 ( \5550 , \5341 , \5352 );
xnor \U$5174 ( \5551 , \5550 , \5330 );
not \U$5175 ( \5552 , \5551 );
not \U$5176 ( \5553 , \5552 );
or \U$5177 ( \5554 , \5549 , \5553 );
not \U$5178 ( \5555 , \5137 );
not \U$5179 ( \5556 , \5519 );
not \U$5180 ( \5557 , \5556 );
not \U$5181 ( \5558 , \5509 );
not \U$5182 ( \5559 , \5558 );
or \U$5183 ( \5560 , \5557 , \5559 );
nand \U$5184 ( \5561 , \5560 , RIc2264d0_37);
not \U$5185 ( \5562 , \5561 );
not \U$5186 ( \5563 , \1082 );
not \U$5187 ( \5564 , \5173 );
or \U$5188 ( \5565 , \5563 , \5564 );
not \U$5189 ( \5566 , RIc2274c0_3);
not \U$5190 ( \5567 , \4123 );
or \U$5191 ( \5568 , \5566 , \5567 );
not \U$5192 ( \5569 , \4414 );
nand \U$5193 ( \5570 , \5569 , \1078 );
nand \U$5194 ( \5571 , \5568 , \5570 );
nand \U$5195 ( \5572 , \5571 , \1040 );
nand \U$5196 ( \5573 , \5565 , \5572 );
not \U$5197 ( \5574 , \5573 );
or \U$5198 ( \5575 , \5562 , \5574 );
or \U$5199 ( \5576 , \5573 , \5561 );
not \U$5200 ( \5577 , \1579 );
not \U$5201 ( \5578 , \5222 );
or \U$5202 ( \5579 , \5577 , \5578 );
and \U$5203 ( \5580 , RIc2275b0_1, \5216 );
not \U$5204 ( \5581 , RIc2275b0_1);
and \U$5205 ( \5582 , \5581 , \5217 );
or \U$5206 ( \5583 , \5580 , \5582 );
nand \U$5207 ( \5584 , \5583 , \854 );
nand \U$5208 ( \5585 , \5579 , \5584 );
nand \U$5209 ( \5586 , \5576 , \5585 );
nand \U$5210 ( \5587 , \5575 , \5586 );
xor \U$5211 ( \5588 , \5555 , \5587 );
xor \U$5212 ( \5589 , \5218 , \5224 );
xor \U$5213 ( \5590 , \5589 , \5235 );
xor \U$5214 ( \5591 , \5588 , \5590 );
not \U$5215 ( \5592 , \5548 );
nand \U$5216 ( \5593 , \5551 , \5592 );
nand \U$5217 ( \5594 , \5591 , \5593 );
nand \U$5218 ( \5595 , \5554 , \5594 );
not \U$5219 ( \5596 , \5595 );
xor \U$5220 ( \5597 , \5428 , \5434 );
xnor \U$5221 ( \5598 , \5597 , \5422 );
nand \U$5222 ( \5599 , \5596 , \5598 );
not \U$5223 ( \5600 , \5460 );
not \U$5224 ( \5601 , \5469 );
or \U$5225 ( \5602 , \5600 , \5601 );
or \U$5226 ( \5603 , \5460 , \5469 );
nand \U$5227 ( \5604 , \5602 , \5603 );
xor \U$5228 ( \5605 , \5604 , \5473 );
and \U$5229 ( \5606 , \5599 , \5605 );
nor \U$5230 ( \5607 , \5596 , \5598 );
nor \U$5231 ( \5608 , \5606 , \5607 );
not \U$5232 ( \5609 , \5608 );
not \U$5233 ( \5610 , \5609 );
xor \U$5234 ( \5611 , \5409 , \5436 );
xnor \U$5235 ( \5612 , \5611 , \5419 );
not \U$5236 ( \5613 , \5612 );
not \U$5237 ( \5614 , \5613 );
or \U$5238 ( \5615 , \5610 , \5614 );
not \U$5239 ( \5616 , \5612 );
not \U$5240 ( \5617 , \5608 );
or \U$5241 ( \5618 , \5616 , \5617 );
xor \U$5242 ( \5619 , \5476 , \5478 );
xor \U$5243 ( \5620 , \5619 , \5484 );
nand \U$5244 ( \5621 , \5618 , \5620 );
nand \U$5245 ( \5622 , \5615 , \5621 );
not \U$5246 ( \5623 , \5622 );
not \U$5247 ( \5624 , \5623 );
or \U$5248 ( \5625 , \5495 , \5624 );
not \U$5249 ( \5626 , \1118 );
not \U$5250 ( \5627 , \1139 );
not \U$5251 ( \5628 , \2105 );
or \U$5252 ( \5629 , \5627 , \5628 );
not \U$5253 ( \5630 , \4501 );
nand \U$5254 ( \5631 , \5630 , RIc2272e0_7);
nand \U$5255 ( \5632 , \5629 , \5631 );
not \U$5256 ( \5633 , \5632 );
or \U$5257 ( \5634 , \5626 , \5633 );
nand \U$5258 ( \5635 , \5388 , \1121 );
nand \U$5259 ( \5636 , \5634 , \5635 );
not \U$5260 ( \5637 , RIc226b60_23);
and \U$5261 ( \5638 , \5637 , \2354 );
not \U$5262 ( \5639 , \5637 );
and \U$5263 ( \5640 , \5639 , \2345 );
nor \U$5264 ( \5641 , \5638 , \5640 );
not \U$5265 ( \5642 , \5641 );
not \U$5266 ( \5643 , \1915 );
not \U$5267 ( \5644 , \5643 );
and \U$5268 ( \5645 , \5642 , \5644 );
and \U$5269 ( \5646 , \5362 , \1930 );
nor \U$5270 ( \5647 , \5645 , \5646 );
not \U$5271 ( \5648 , \4387 );
not \U$5272 ( \5649 , \4393 );
or \U$5273 ( \5650 , \5648 , \5649 );
not \U$5274 ( \5651 , \4072 );
nand \U$5275 ( \5652 , \5650 , \5651 );
not \U$5276 ( \5653 , \5652 );
nor \U$5277 ( \5654 , \4087 , \4394 );
nand \U$5278 ( \5655 , \4084 , \5654 );
nand \U$5279 ( \5656 , \5653 , \5655 );
nand \U$5280 ( \5657 , \5198 , \657 );
not \U$5281 ( \5658 , \5657 );
and \U$5282 ( \5659 , \5656 , \5658 );
not \U$5283 ( \5660 , \5656 );
and \U$5284 ( \5661 , \5660 , \5657 );
nor \U$5285 ( \5662 , \5659 , \5661 );
buf \U$5286 ( \5663 , \5662 );
not \U$5287 ( \5664 , \5663 );
buf \U$5288 ( \5665 , \5664 );
not \U$5289 ( \5666 , \5665 );
nand \U$5290 ( \5667 , \5666 , RIc2275b0_1);
nand \U$5291 ( \5668 , \5647 , \5667 );
and \U$5292 ( \5669 , \5636 , \5668 );
nor \U$5293 ( \5670 , \5647 , \5667 );
nor \U$5294 ( \5671 , \5669 , \5670 );
not \U$5295 ( \5672 , \5671 );
not \U$5296 ( \5673 , \2784 );
and \U$5297 ( \5674 , RIc226890_29, \1440 );
not \U$5298 ( \5675 , RIc226890_29);
and \U$5299 ( \5676 , \5675 , \1223 );
or \U$5300 ( \5677 , \5674 , \5676 );
not \U$5301 ( \5678 , \5677 );
or \U$5302 ( \5679 , \5673 , \5678 );
nand \U$5303 ( \5680 , \5257 , \2086 );
nand \U$5304 ( \5681 , \5679 , \5680 );
not \U$5305 ( \5682 , \5681 );
and \U$5306 ( \5683 , \5303 , \3653 );
and \U$5307 ( \5684 , \2119 , \2072 );
not \U$5308 ( \5685 , \2119 );
and \U$5309 ( \5686 , \5685 , RIc2267a0_31);
or \U$5310 ( \5687 , \5684 , \5686 );
and \U$5311 ( \5688 , \5687 , \2697 );
nor \U$5312 ( \5689 , \5683 , \5688 );
nand \U$5313 ( \5690 , \5682 , \5689 );
not \U$5314 ( \5691 , \5274 );
not \U$5315 ( \5692 , \2534 );
or \U$5316 ( \5693 , \5691 , \5692 );
not \U$5317 ( \5694 , \2229 );
not \U$5318 ( \5695 , \1941 );
and \U$5319 ( \5696 , \5694 , \5695 );
buf \U$5320 ( \5697 , \3851 );
and \U$5321 ( \5698 , \5697 , \1941 );
nor \U$5322 ( \5699 , \5696 , \5698 );
not \U$5323 ( \5700 , \2518 );
or \U$5324 ( \5701 , \5699 , \5700 );
nand \U$5325 ( \5702 , \5693 , \5701 );
and \U$5326 ( \5703 , \5690 , \5702 );
not \U$5327 ( \5704 , \5681 );
nor \U$5328 ( \5705 , \5704 , \5689 );
nor \U$5329 ( \5706 , \5703 , \5705 );
not \U$5330 ( \5707 , \5706 );
or \U$5331 ( \5708 , \5672 , \5707 );
not \U$5332 ( \5709 , \2392 );
not \U$5333 ( \5710 , RIc226c50_21);
not \U$5334 ( \5711 , \2424 );
or \U$5335 ( \5712 , \5710 , \5711 );
nand \U$5336 ( \5713 , \2423 , \2383 );
nand \U$5337 ( \5714 , \5712 , \5713 );
not \U$5338 ( \5715 , \5714 );
or \U$5339 ( \5716 , \5709 , \5715 );
nand \U$5340 ( \5717 , \5233 , \2367 );
nand \U$5341 ( \5718 , \5716 , \5717 );
not \U$5342 ( \5719 , \5718 );
and \U$5343 ( \5720 , \5162 , \954 );
not \U$5344 ( \5721 , RIc2273d0_5);
not \U$5345 ( \5722 , \3729 );
or \U$5346 ( \5723 , \5721 , \5722 );
nand \U$5347 ( \5724 , \3728 , \946 );
nand \U$5348 ( \5725 , \5723 , \5724 );
and \U$5349 ( \5726 , \5725 , \951 );
nor \U$5350 ( \5727 , \5720 , \5726 );
not \U$5351 ( \5728 , \5727 );
not \U$5352 ( \5729 , \5728 );
or \U$5353 ( \5730 , \5719 , \5729 );
not \U$5354 ( \5731 , \5727 );
not \U$5355 ( \5732 , \5718 );
not \U$5356 ( \5733 , \5732 );
or \U$5357 ( \5734 , \5731 , \5733 );
not \U$5358 ( \5735 , RIc2265c0_35);
not \U$5359 ( \5736 , \1074 );
or \U$5360 ( \5737 , \5735 , \5736 );
nand \U$5361 ( \5738 , \1073 , \4376 );
nand \U$5362 ( \5739 , \5737 , \5738 );
not \U$5363 ( \5740 , \4380 );
not \U$5364 ( \5741 , \5740 );
and \U$5365 ( \5742 , \5739 , \5741 );
and \U$5366 ( \5743 , \5132 , \5135 );
nor \U$5367 ( \5744 , \5742 , \5743 );
not \U$5368 ( \5745 , \5744 );
nand \U$5369 ( \5746 , \5734 , \5745 );
nand \U$5370 ( \5747 , \5730 , \5746 );
nand \U$5371 ( \5748 , \5708 , \5747 );
not \U$5372 ( \5749 , \5706 );
not \U$5373 ( \5750 , \5671 );
nand \U$5374 ( \5751 , \5749 , \5750 );
and \U$5375 ( \5752 , \5748 , \5751 );
not \U$5376 ( \5753 , \2138 );
not \U$5377 ( \5754 , RIc226980_27);
not \U$5378 ( \5755 , \1530 );
or \U$5379 ( \5756 , \5754 , \5755 );
nand \U$5380 ( \5757 , \3581 , \2150 );
nand \U$5381 ( \5758 , \5756 , \5757 );
not \U$5382 ( \5759 , \5758 );
or \U$5383 ( \5760 , \5753 , \5759 );
nand \U$5384 ( \5761 , \5249 , \2156 );
nand \U$5385 ( \5762 , \5760 , \5761 );
not \U$5386 ( \5763 , \5762 );
not \U$5387 ( \5764 , \5763 );
not \U$5388 ( \5765 , \1945 );
not \U$5389 ( \5766 , RIc226e30_17);
not \U$5390 ( \5767 , \3834 );
buf \U$5391 ( \5768 , \5767 );
not \U$5392 ( \5769 , \5768 );
or \U$5393 ( \5770 , \5766 , \5769 );
nand \U$5394 ( \5771 , \3840 , \1960 );
nand \U$5395 ( \5772 , \5770 , \5771 );
not \U$5396 ( \5773 , \5772 );
or \U$5397 ( \5774 , \5765 , \5773 );
nand \U$5398 ( \5775 , \5292 , \1963 );
nand \U$5399 ( \5776 , \5774 , \5775 );
not \U$5400 ( \5777 , \5776 );
not \U$5401 ( \5778 , \5777 );
or \U$5402 ( \5779 , \5764 , \5778 );
not \U$5403 ( \5780 , \2179 );
not \U$5404 ( \5781 , \2692 );
and \U$5405 ( \5782 , \5780 , \5781 );
and \U$5406 ( \5783 , \841 , \2692 );
nor \U$5407 ( \5784 , \5782 , \5783 );
or \U$5408 ( \5785 , \5784 , \5185 );
or \U$5409 ( \5786 , \5183 , \4440 );
nand \U$5410 ( \5787 , \5785 , \5786 );
nand \U$5411 ( \5788 , \5779 , \5787 );
nand \U$5412 ( \5789 , \5776 , \5762 );
nand \U$5413 ( \5790 , \5788 , \5789 );
not \U$5414 ( \5791 , \5790 );
not \U$5415 ( \5792 , \2195 );
not \U$5416 ( \5793 , RIc226a70_25);
not \U$5417 ( \5794 , \3044 );
or \U$5418 ( \5795 , \5793 , \5794 );
nand \U$5419 ( \5796 , \1486 , \2187 );
nand \U$5420 ( \5797 , \5795 , \5796 );
not \U$5421 ( \5798 , \5797 );
or \U$5422 ( \5799 , \5792 , \5798 );
nand \U$5423 ( \5800 , \5335 , \2173 );
nand \U$5424 ( \5801 , \5799 , \5800 );
not \U$5425 ( \5802 , \5801 );
not \U$5426 ( \5803 , \2358 );
not \U$5427 ( \5804 , \5312 );
or \U$5428 ( \5805 , \5803 , \5804 );
not \U$5429 ( \5806 , RIc226f20_15);
not \U$5430 ( \5807 , \2592 );
or \U$5431 ( \5808 , \5806 , \5807 );
not \U$5432 ( \5809 , \3292 );
nand \U$5433 ( \5810 , \5809 , \2351 );
nand \U$5434 ( \5811 , \5808 , \5810 );
nand \U$5435 ( \5812 , \5811 , \2320 );
nand \U$5436 ( \5813 , \5805 , \5812 );
not \U$5437 ( \5814 , \5813 );
or \U$5438 ( \5815 , \5802 , \5814 );
or \U$5439 ( \5816 , \5813 , \5801 );
not \U$5440 ( \5817 , \1680 );
not \U$5441 ( \5818 , RIc227010_13);
not \U$5442 ( \5819 , \2479 );
not \U$5443 ( \5820 , \5819 );
or \U$5444 ( \5821 , \5818 , \5820 );
nand \U$5445 ( \5822 , \2479 , \1296 );
nand \U$5446 ( \5823 , \5821 , \5822 );
not \U$5447 ( \5824 , \5823 );
or \U$5448 ( \5825 , \5817 , \5824 );
nand \U$5449 ( \5826 , \5326 , \1682 );
nand \U$5450 ( \5827 , \5825 , \5826 );
nand \U$5451 ( \5828 , \5816 , \5827 );
nand \U$5452 ( \5829 , \5815 , \5828 );
not \U$5453 ( \5830 , \5829 );
nand \U$5454 ( \5831 , \5791 , \5830 );
not \U$5455 ( \5832 , \5392 );
not \U$5456 ( \5833 , \5832 );
not \U$5457 ( \5834 , \5378 );
not \U$5458 ( \5835 , \5367 );
not \U$5459 ( \5836 , \5835 );
or \U$5460 ( \5837 , \5834 , \5836 );
or \U$5461 ( \5838 , \5835 , \5378 );
nand \U$5462 ( \5839 , \5837 , \5838 );
not \U$5463 ( \5840 , \5839 );
or \U$5464 ( \5841 , \5833 , \5840 );
or \U$5465 ( \5842 , \5839 , \5832 );
nand \U$5466 ( \5843 , \5841 , \5842 );
and \U$5467 ( \5844 , \5831 , \5843 );
and \U$5468 ( \5845 , \5790 , \5829 );
nor \U$5469 ( \5846 , \5844 , \5845 );
nand \U$5470 ( \5847 , \5752 , \5846 );
xor \U$5471 ( \5848 , \5555 , \5587 );
and \U$5472 ( \5849 , \5848 , \5590 );
and \U$5473 ( \5850 , \5555 , \5587 );
or \U$5474 ( \5851 , \5849 , \5850 );
and \U$5475 ( \5852 , \5847 , \5851 );
nor \U$5476 ( \5853 , \5752 , \5846 );
nor \U$5477 ( \5854 , \5852 , \5853 );
not \U$5478 ( \5855 , \5854 );
not \U$5479 ( \5856 , \5855 );
and \U$5480 ( \5857 , \5394 , \5355 );
not \U$5481 ( \5858 , \5394 );
and \U$5482 ( \5859 , \5858 , \5396 );
nor \U$5483 ( \5860 , \5857 , \5859 );
and \U$5484 ( \5861 , \5860 , \5398 );
not \U$5485 ( \5862 , \5860 );
and \U$5486 ( \5863 , \5862 , \5399 );
nor \U$5487 ( \5864 , \5861 , \5863 );
xor \U$5488 ( \5865 , \5238 , \5279 );
xor \U$5489 ( \5866 , \5865 , \5192 );
nand \U$5490 ( \5867 , \5864 , \5866 );
not \U$5491 ( \5868 , \5305 );
xor \U$5492 ( \5869 , \5294 , \5868 );
xor \U$5493 ( \5870 , \5869 , \5316 );
not \U$5494 ( \5871 , \5870 );
not \U$5495 ( \5872 , \5871 );
not \U$5496 ( \5873 , \5175 );
not \U$5497 ( \5874 , \5189 );
or \U$5498 ( \5875 , \5873 , \5874 );
or \U$5499 ( \5876 , \5189 , \5175 );
nand \U$5500 ( \5877 , \5875 , \5876 );
xnor \U$5501 ( \5878 , \5877 , \5164 );
not \U$5502 ( \5879 , \5878 );
not \U$5503 ( \5880 , \5879 );
or \U$5504 ( \5881 , \5872 , \5880 );
not \U$5505 ( \5882 , \5878 );
not \U$5506 ( \5883 , \5870 );
or \U$5507 ( \5884 , \5882 , \5883 );
xor \U$5508 ( \5885 , \5261 , \5251 );
xor \U$5509 ( \5886 , \5885 , \5276 );
nand \U$5510 ( \5887 , \5884 , \5886 );
nand \U$5511 ( \5888 , \5881 , \5887 );
and \U$5512 ( \5889 , \5867 , \5888 );
nor \U$5513 ( \5890 , \5864 , \5866 );
nor \U$5514 ( \5891 , \5889 , \5890 );
not \U$5515 ( \5892 , \5891 );
not \U$5516 ( \5893 , \5892 );
or \U$5517 ( \5894 , \5856 , \5893 );
not \U$5518 ( \5895 , \5891 );
not \U$5519 ( \5896 , \5854 );
or \U$5520 ( \5897 , \5895 , \5896 );
xor \U$5521 ( \5898 , \5153 , \5284 );
xor \U$5522 ( \5899 , \5898 , \5401 );
nand \U$5523 ( \5900 , \5897 , \5899 );
nand \U$5524 ( \5901 , \5894 , \5900 );
buf \U$5525 ( \5902 , \5901 );
nand \U$5526 ( \5903 , \5625 , \5902 );
not \U$5527 ( \5904 , \5494 );
nand \U$5528 ( \5905 , \5904 , \5622 );
and \U$5529 ( \5906 , \5903 , \5905 );
xor \U$5530 ( \5907 , \5491 , \5906 );
xor \U$5531 ( \5908 , \5126 , \5443 );
xor \U$5532 ( \5909 , \5908 , \5446 );
and \U$5533 ( \5910 , \5907 , \5909 );
and \U$5534 ( \5911 , \5491 , \5906 );
or \U$5535 ( \5912 , \5910 , \5911 );
nand \U$5536 ( \5913 , \5450 , \5912 );
not \U$5537 ( \5914 , \5913 );
xor \U$5538 ( \5915 , \5491 , \5906 );
xor \U$5539 ( \5916 , \5915 , \5909 );
xor \U$5540 ( \5917 , \5901 , \5493 );
xor \U$5541 ( \5918 , \5917 , \5623 );
buf \U$5542 ( \5919 , \5918 );
xor \U$5543 ( \5920 , \5487 , \5452 );
and \U$5544 ( \5921 , \5920 , \5489 );
not \U$5545 ( \5922 , \5920 );
and \U$5546 ( \5923 , \5922 , \5456 );
nor \U$5547 ( \5924 , \5921 , \5923 );
not \U$5548 ( \5925 , \5924 );
nand \U$5549 ( \5926 , \5919 , \5925 );
xor \U$5550 ( \5927 , \5609 , \5613 );
buf \U$5551 ( \5928 , \5620 );
xor \U$5552 ( \5929 , \5927 , \5928 );
not \U$5553 ( \5930 , \5929 );
xor \U$5554 ( \5931 , \5899 , \5855 );
xor \U$5555 ( \5932 , \5931 , \5892 );
not \U$5556 ( \5933 , \5932 );
not \U$5557 ( \5934 , \2697 );
not \U$5558 ( \5935 , RIc2267a0_31);
not \U$5559 ( \5936 , \1404 );
or \U$5560 ( \5937 , \5935 , \5936 );
nand \U$5561 ( \5938 , \1228 , \2705 );
nand \U$5562 ( \5939 , \5937 , \5938 );
not \U$5563 ( \5940 , \5939 );
or \U$5564 ( \5941 , \5934 , \5940 );
nand \U$5565 ( \5942 , \5687 , \3653 );
nand \U$5566 ( \5943 , \5941 , \5942 );
not \U$5567 ( \5944 , \5943 );
and \U$5568 ( \5945 , \5714 , \2367 );
not \U$5569 ( \5946 , RIc226c50_21);
not \U$5570 ( \5947 , \2834 );
or \U$5571 ( \5948 , \5946 , \5947 );
not \U$5572 ( \5949 , \2444 );
nand \U$5573 ( \5950 , \5949 , \2370 );
nand \U$5574 ( \5951 , \5948 , \5950 );
and \U$5575 ( \5952 , \5951 , \2392 );
nor \U$5576 ( \5953 , \5945 , \5952 );
not \U$5577 ( \5954 , \5953 );
not \U$5578 ( \5955 , \5954 );
or \U$5579 ( \5956 , \5944 , \5955 );
not \U$5580 ( \5957 , \5953 );
not \U$5581 ( \5958 , \5943 );
not \U$5582 ( \5959 , \5958 );
or \U$5583 ( \5960 , \5957 , \5959 );
not \U$5584 ( \5961 , \5741 );
not \U$5585 ( \5962 , RIc2265c0_35);
not \U$5586 ( \5963 , \890 );
or \U$5587 ( \5964 , \5962 , \5963 );
nand \U$5588 ( \5965 , \889 , \3620 );
nand \U$5589 ( \5966 , \5964 , \5965 );
not \U$5590 ( \5967 , \5966 );
or \U$5591 ( \5968 , \5961 , \5967 );
nand \U$5592 ( \5969 , \5739 , \5135 );
nand \U$5593 ( \5970 , \5968 , \5969 );
nand \U$5594 ( \5971 , \5960 , \5970 );
nand \U$5595 ( \5972 , \5956 , \5971 );
not \U$5596 ( \5973 , \5972 );
not \U$5597 ( \5974 , \2078 );
and \U$5598 ( \5975 , RIc226890_29, \1393 );
not \U$5599 ( \5976 , RIc226890_29);
and \U$5600 ( \5977 , \5976 , \1396 );
or \U$5601 ( \5978 , \5975 , \5977 );
not \U$5602 ( \5979 , \5978 );
or \U$5603 ( \5980 , \5974 , \5979 );
nand \U$5604 ( \5981 , \5677 , \2086 );
nand \U$5605 ( \5982 , \5980 , \5981 );
not \U$5606 ( \5983 , \5982 );
not \U$5607 ( \5984 , \1945 );
not \U$5608 ( \5985 , RIc226e30_17);
not \U$5609 ( \5986 , \2015 );
or \U$5610 ( \5987 , \5985 , \5986 );
nand \U$5611 ( \5988 , \3508 , \1935 );
nand \U$5612 ( \5989 , \5987 , \5988 );
not \U$5613 ( \5990 , \5989 );
or \U$5614 ( \5991 , \5984 , \5990 );
nand \U$5615 ( \5992 , \5772 , \1963 );
nand \U$5616 ( \5993 , \5991 , \5992 );
not \U$5617 ( \5994 , \5993 );
or \U$5618 ( \5995 , \5983 , \5994 );
or \U$5619 ( \5996 , \5982 , \5993 );
not \U$5620 ( \5997 , \2518 );
not \U$5621 ( \5998 , RIc226d40_19);
not \U$5622 ( \5999 , \2258 );
or \U$5623 ( \6000 , \5998 , \5999 );
nand \U$5624 ( \6001 , \2261 , \2523 );
nand \U$5625 ( \6002 , \6000 , \6001 );
not \U$5626 ( \6003 , \6002 );
or \U$5627 ( \6004 , \5997 , \6003 );
not \U$5628 ( \6005 , \5699 );
nand \U$5629 ( \6006 , \6005 , \2534 );
nand \U$5630 ( \6007 , \6004 , \6006 );
nand \U$5631 ( \6008 , \5996 , \6007 );
nand \U$5632 ( \6009 , \5995 , \6008 );
not \U$5633 ( \6010 , \6009 );
nand \U$5634 ( \6011 , \5973 , \6010 );
not \U$5635 ( \6012 , \5725 );
not \U$5636 ( \6013 , \954 );
or \U$5637 ( \6014 , \6012 , \6013 );
not \U$5638 ( \6015 , RIc2273d0_5);
not \U$5639 ( \6016 , \4046 );
or \U$5640 ( \6017 , \6015 , \6016 );
nand \U$5641 ( \6018 , \3641 , \935 );
nand \U$5642 ( \6019 , \6017 , \6018 );
nand \U$5643 ( \6020 , \6019 , \951 );
nand \U$5644 ( \6021 , \6014 , \6020 );
not \U$5645 ( \6022 , \1118 );
not \U$5646 ( \6023 , RIc2272e0_7);
not \U$5647 ( \6024 , \3121 );
or \U$5648 ( \6025 , \6023 , \6024 );
nand \U$5649 ( \6026 , \3122 , \1139 );
nand \U$5650 ( \6027 , \6025 , \6026 );
not \U$5651 ( \6028 , \6027 );
or \U$5652 ( \6029 , \6022 , \6028 );
nand \U$5653 ( \6030 , \5632 , \1121 );
nand \U$5654 ( \6031 , \6029 , \6030 );
xor \U$5655 ( \6032 , \6021 , \6031 );
not \U$5656 ( \6033 , \1915 );
not \U$5657 ( \6034 , RIc226b60_23);
not \U$5658 ( \6035 , \2774 );
or \U$5659 ( \6036 , \6034 , \6035 );
nand \U$5660 ( \6037 , \2306 , \2111 );
nand \U$5661 ( \6038 , \6036 , \6037 );
not \U$5662 ( \6039 , \6038 );
or \U$5663 ( \6040 , \6033 , \6039 );
not \U$5664 ( \6041 , \5641 );
nand \U$5665 ( \6042 , \6041 , \1930 );
nand \U$5666 ( \6043 , \6040 , \6042 );
and \U$5667 ( \6044 , \6032 , \6043 );
and \U$5668 ( \6045 , \6021 , \6031 );
or \U$5669 ( \6046 , \6044 , \6045 );
and \U$5670 ( \6047 , \6011 , \6046 );
nor \U$5671 ( \6048 , \5973 , \6010 );
nor \U$5672 ( \6049 , \6047 , \6048 );
not \U$5673 ( \6050 , \6049 );
not \U$5674 ( \6051 , \6050 );
xor \U$5675 ( \6052 , \5829 , \5790 );
xor \U$5676 ( \6053 , \6052 , \5843 );
not \U$5677 ( \6054 , \6053 );
or \U$5678 ( \6055 , \6051 , \6054 );
or \U$5679 ( \6056 , \6053 , \6050 );
nand \U$5680 ( \6057 , \528 , \649 );
nor \U$5681 ( \6058 , \6057 , \4087 );
nand \U$5682 ( \6059 , \4084 , \6058 );
not \U$5683 ( \6060 , \6057 );
nand \U$5684 ( \6061 , \6060 , \4393 );
and \U$5685 ( \6062 , \650 , \652 );
nand \U$5686 ( \6063 , \6059 , \6061 , \6062 );
nand \U$5687 ( \6064 , \651 , \4067 );
not \U$5688 ( \6065 , \6064 );
and \U$5689 ( \6066 , \6063 , \6065 );
not \U$5690 ( \6067 , \6063 );
and \U$5691 ( \6068 , \6067 , \6064 );
nor \U$5692 ( \6069 , \6066 , \6068 );
buf \U$5693 ( \6070 , \6069 );
buf \U$5694 ( \6071 , \6070 );
and \U$5695 ( \6072 , RIc2275b0_1, \6071 );
not \U$5696 ( \6073 , \6072 );
not \U$5697 ( \6074 , \6073 );
not \U$5698 ( \6075 , RIc2274c0_3);
not \U$5699 ( \6076 , \4406 );
not \U$5700 ( \6077 , \6076 );
or \U$5701 ( \6078 , \6075 , \6077 );
not \U$5702 ( \6079 , \6076 );
nand \U$5703 ( \6080 , \6079 , \1078 );
nand \U$5704 ( \6081 , \6078 , \6080 );
and \U$5705 ( \6082 , \6081 , \1040 );
and \U$5706 ( \6083 , \5571 , \1082 );
nor \U$5707 ( \6084 , \6082 , \6083 );
not \U$5708 ( \6085 , \6084 );
or \U$5709 ( \6086 , \6074 , \6085 );
not \U$5710 ( \6087 , \854 );
and \U$5711 ( \6088 , RIc2275b0_1, \5665 );
not \U$5712 ( \6089 , RIc2275b0_1);
and \U$5713 ( \6090 , \6089 , \5666 );
or \U$5714 ( \6091 , \6088 , \6090 );
not \U$5715 ( \6092 , \6091 );
or \U$5716 ( \6093 , \6087 , \6092 );
nand \U$5717 ( \6094 , \5583 , \1579 );
nand \U$5718 ( \6095 , \6093 , \6094 );
nand \U$5719 ( \6096 , \6086 , \6095 );
not \U$5720 ( \6097 , \6084 );
nand \U$5721 ( \6098 , \6097 , \6072 );
nand \U$5722 ( \6099 , \6096 , \6098 );
xor \U$5723 ( \6100 , \5585 , \5573 );
xor \U$5724 ( \6101 , \6100 , \5561 );
xor \U$5725 ( \6102 , \6099 , \6101 );
not \U$5726 ( \6103 , \2195 );
not \U$5727 ( \6104 , \1730 );
not \U$5728 ( \6105 , \2190 );
and \U$5729 ( \6106 , \6104 , \6105 );
not \U$5730 ( \6107 , RIc226a70_25);
and \U$5731 ( \6108 , \1730 , \6107 );
nor \U$5732 ( \6109 , \6106 , \6108 );
not \U$5733 ( \6110 , \6109 );
not \U$5734 ( \6111 , \6110 );
or \U$5735 ( \6112 , \6103 , \6111 );
nand \U$5736 ( \6113 , \5797 , \2173 );
nand \U$5737 ( \6114 , \6112 , \6113 );
not \U$5738 ( \6115 , \6114 );
not \U$5739 ( \6116 , \1307 );
not \U$5740 ( \6117 , RIc227100_11);
not \U$5741 ( \6118 , \2645 );
or \U$5742 ( \6119 , \6117 , \6118 );
not \U$5743 ( \6120 , \3011 );
nand \U$5744 ( \6121 , \6120 , \3351 );
nand \U$5745 ( \6122 , \6119 , \6121 );
not \U$5746 ( \6123 , \6122 );
or \U$5747 ( \6124 , \6116 , \6123 );
nand \U$5748 ( \6125 , \5541 , \1311 );
nand \U$5749 ( \6126 , \6124 , \6125 );
not \U$5750 ( \6127 , \6126 );
or \U$5751 ( \6128 , \6115 , \6127 );
or \U$5752 ( \6129 , \6126 , \6114 );
xnor \U$5753 ( \6130 , \1758 , \2501 );
not \U$5754 ( \6131 , \6130 );
not \U$5755 ( \6132 , \1679 );
and \U$5756 ( \6133 , \6131 , \6132 );
and \U$5757 ( \6134 , \5823 , \1682 );
nor \U$5758 ( \6135 , \6133 , \6134 );
not \U$5759 ( \6136 , \6135 );
nand \U$5760 ( \6137 , \6129 , \6136 );
nand \U$5761 ( \6138 , \6128 , \6137 );
and \U$5762 ( \6139 , \6102 , \6138 );
and \U$5763 ( \6140 , \6099 , \6101 );
or \U$5764 ( \6141 , \6139 , \6140 );
nand \U$5765 ( \6142 , \6056 , \6141 );
nand \U$5766 ( \6143 , \6055 , \6142 );
not \U$5767 ( \6144 , \6143 );
xor \U$5768 ( \6145 , \5851 , \5752 );
xnor \U$5769 ( \6146 , \6145 , \5846 );
not \U$5770 ( \6147 , \6146 );
not \U$5771 ( \6148 , \6147 );
or \U$5772 ( \6149 , \6144 , \6148 );
not \U$5773 ( \6150 , \6146 );
not \U$5774 ( \6151 , \6143 );
not \U$5775 ( \6152 , \6151 );
or \U$5776 ( \6153 , \6150 , \6152 );
xor \U$5777 ( \6154 , \5521 , \5534 );
xor \U$5778 ( \6155 , \6154 , \5545 );
not \U$5779 ( \6156 , \6155 );
and \U$5780 ( \6157 , \5777 , \5762 );
not \U$5781 ( \6158 , \5777 );
and \U$5782 ( \6159 , \6158 , \5763 );
or \U$5783 ( \6160 , \6157 , \6159 );
xor \U$5784 ( \6161 , \6160 , \5787 );
not \U$5785 ( \6162 , \6161 );
or \U$5786 ( \6163 , \6156 , \6162 );
or \U$5787 ( \6164 , \6161 , \6155 );
xor \U$5788 ( \6165 , \5667 , \5647 );
xor \U$5789 ( \6166 , \6165 , \5636 );
nand \U$5790 ( \6167 , \6164 , \6166 );
nand \U$5791 ( \6168 , \6163 , \6167 );
not \U$5792 ( \6169 , \6168 );
not \U$5793 ( \6170 , \5706 );
not \U$5794 ( \6171 , \5750 );
or \U$5795 ( \6172 , \6170 , \6171 );
nand \U$5796 ( \6173 , \5749 , \5671 );
nand \U$5797 ( \6174 , \6172 , \6173 );
xor \U$5798 ( \6175 , \6174 , \5747 );
not \U$5799 ( \6176 , \6175 );
or \U$5800 ( \6177 , \6169 , \6176 );
or \U$5801 ( \6178 , \6168 , \6175 );
xor \U$5802 ( \6179 , \5681 , \5689 );
xnor \U$5803 ( \6180 , \6179 , \5702 );
not \U$5804 ( \6181 , \6180 );
not \U$5805 ( \6182 , \2320 );
not \U$5806 ( \6183 , RIc226f20_15);
not \U$5807 ( \6184 , \4803 );
or \U$5808 ( \6185 , \6183 , \6184 );
nand \U$5809 ( \6186 , \2559 , \1674 );
nand \U$5810 ( \6187 , \6185 , \6186 );
not \U$5811 ( \6188 , \6187 );
or \U$5812 ( \6189 , \6182 , \6188 );
nand \U$5813 ( \6190 , \5811 , \2358 );
nand \U$5814 ( \6191 , \6189 , \6190 );
not \U$5815 ( \6192 , \2138 );
not \U$5816 ( \6193 , RIc226980_27);
not \U$5817 ( \6194 , \1949 );
or \U$5818 ( \6195 , \6193 , \6194 );
nand \U$5819 ( \6196 , \4778 , \2150 );
nand \U$5820 ( \6197 , \6195 , \6196 );
not \U$5821 ( \6198 , \6197 );
or \U$5822 ( \6199 , \6192 , \6198 );
nand \U$5823 ( \6200 , \5758 , \2154 );
nand \U$5824 ( \6201 , \6199 , \6200 );
or \U$5825 ( \6202 , \6191 , \6201 );
not \U$5826 ( \6203 , \3629 );
not \U$5827 ( \6204 , RIc2266b0_33);
not \U$5828 ( \6205 , \1490 );
or \U$5829 ( \6206 , \6204 , \6205 );
nand \U$5830 ( \6207 , \984 , \5179 );
nand \U$5831 ( \6208 , \6206 , \6207 );
not \U$5832 ( \6209 , \6208 );
or \U$5833 ( \6210 , \6203 , \6209 );
not \U$5834 ( \6211 , \5784 );
nand \U$5835 ( \6212 , \6211 , \3631 );
nand \U$5836 ( \6213 , \6210 , \6212 );
and \U$5837 ( \6214 , \6202 , \6213 );
and \U$5838 ( \6215 , \6191 , \6201 );
nor \U$5839 ( \6216 , \6214 , \6215 );
nand \U$5840 ( \6217 , \6181 , \6216 );
not \U$5841 ( \6218 , \6217 );
not \U$5842 ( \6219 , \5745 );
not \U$5843 ( \6220 , \5732 );
or \U$5844 ( \6221 , \6219 , \6220 );
nand \U$5845 ( \6222 , \5718 , \5744 );
nand \U$5846 ( \6223 , \6221 , \6222 );
not \U$5847 ( \6224 , \5728 );
xnor \U$5848 ( \6225 , \6223 , \6224 );
not \U$5849 ( \6226 , \6225 );
or \U$5850 ( \6227 , \6218 , \6226 );
not \U$5851 ( \6228 , \6216 );
nand \U$5852 ( \6229 , \6180 , \6228 );
nand \U$5853 ( \6230 , \6227 , \6229 );
nand \U$5854 ( \6231 , \6178 , \6230 );
nand \U$5855 ( \6232 , \6177 , \6231 );
nand \U$5856 ( \6233 , \6153 , \6232 );
nand \U$5857 ( \6234 , \6149 , \6233 );
not \U$5858 ( \6235 , \6234 );
nand \U$5859 ( \6236 , \5933 , \6235 );
not \U$5860 ( \6237 , \6236 );
or \U$5861 ( \6238 , \5930 , \6237 );
nand \U$5862 ( \6239 , \5932 , \6234 );
nand \U$5863 ( \6240 , \6238 , \6239 );
and \U$5864 ( \6241 , \5926 , \6240 );
nor \U$5865 ( \6242 , \5919 , \5925 );
nor \U$5866 ( \6243 , \6241 , \6242 );
nand \U$5867 ( \6244 , \5916 , \6243 );
buf \U$5868 ( \6245 , \6244 );
not \U$5869 ( \6246 , \6240 );
xor \U$5870 ( \6247 , \5918 , \5924 );
not \U$5871 ( \6248 , \6247 );
or \U$5872 ( \6249 , \6246 , \6248 );
or \U$5873 ( \6250 , \6247 , \6240 );
nand \U$5874 ( \6251 , \6249 , \6250 );
not \U$5875 ( \6252 , \5878 );
not \U$5876 ( \6253 , \5871 );
or \U$5877 ( \6254 , \6252 , \6253 );
nand \U$5878 ( \6255 , \5879 , \5870 );
nand \U$5879 ( \6256 , \6254 , \6255 );
and \U$5880 ( \6257 , \6256 , \5886 );
not \U$5881 ( \6258 , \6256 );
not \U$5882 ( \6259 , \5886 );
and \U$5883 ( \6260 , \6258 , \6259 );
nor \U$5884 ( \6261 , \6257 , \6260 );
not \U$5885 ( \6262 , \6261 );
not \U$5886 ( \6263 , \6262 );
xor \U$5887 ( \6264 , \5592 , \5552 );
xor \U$5888 ( \6265 , \6264 , \5591 );
not \U$5889 ( \6266 , \6265 );
or \U$5890 ( \6267 , \6263 , \6266 );
not \U$5891 ( \6268 , \5521 );
not \U$5892 ( \6269 , \1597 );
not \U$5893 ( \6270 , RIc2271f0_9);
not \U$5894 ( \6271 , \3564 );
or \U$5895 ( \6272 , \6270 , \6271 );
nand \U$5896 ( \6273 , \2636 , \1351 );
nand \U$5897 ( \6274 , \6272 , \6273 );
not \U$5898 ( \6275 , \6274 );
or \U$5899 ( \6276 , \6269 , \6275 );
nand \U$5900 ( \6277 , \5530 , \1340 );
nand \U$5901 ( \6278 , \6276 , \6277 );
xor \U$5902 ( \6279 , \6268 , \6278 );
not \U$5903 ( \6280 , \954 );
not \U$5904 ( \6281 , \6019 );
or \U$5905 ( \6282 , \6280 , \6281 );
not \U$5906 ( \6283 , RIc2273d0_5);
not \U$5907 ( \6284 , \4123 );
or \U$5908 ( \6285 , \6283 , \6284 );
nand \U$5909 ( \6286 , \4124 , \946 );
nand \U$5910 ( \6287 , \6285 , \6286 );
nand \U$5911 ( \6288 , \6287 , \951 );
nand \U$5912 ( \6289 , \6282 , \6288 );
not \U$5913 ( \6290 , \1082 );
not \U$5914 ( \6291 , \6081 );
or \U$5915 ( \6292 , \6290 , \6291 );
not \U$5916 ( \6293 , RIc2274c0_3);
not \U$5917 ( \6294 , \5216 );
or \U$5918 ( \6295 , \6293 , \6294 );
nand \U$5919 ( \6296 , \5217 , \2896 );
nand \U$5920 ( \6297 , \6295 , \6296 );
nand \U$5921 ( \6298 , \6297 , \1040 );
nand \U$5922 ( \6299 , \6292 , \6298 );
or \U$5923 ( \6300 , \6289 , \6299 );
and \U$5924 ( \6301 , RIc226368_40, RIc2262f0_41);
not \U$5925 ( \6302 , RIc226368_40);
not \U$5926 ( \6303 , RIc2262f0_41);
and \U$5927 ( \6304 , \6302 , \6303 );
nor \U$5928 ( \6305 , \6301 , \6304 );
buf \U$5929 ( \6306 , \6305 );
buf \U$5930 ( \6307 , \6306 );
not \U$5931 ( \6308 , \6307 );
not \U$5932 ( \6309 , \6308 );
and \U$5933 ( \6310 , RIc2263e0_39, RIc226368_40);
nor \U$5934 ( \6311 , RIc2263e0_39, RIc226368_40);
nor \U$5935 ( \6312 , \6310 , \6305 , \6311 );
not \U$5936 ( \6313 , \6312 );
not \U$5937 ( \6314 , \6313 );
or \U$5938 ( \6315 , \6309 , \6314 );
nand \U$5939 ( \6316 , \6315 , RIc2263e0_39);
nand \U$5940 ( \6317 , \6300 , \6316 );
nand \U$5941 ( \6318 , \6289 , \6299 );
nand \U$5942 ( \6319 , \6317 , \6318 );
and \U$5943 ( \6320 , \6279 , \6319 );
and \U$5944 ( \6321 , \6268 , \6278 );
or \U$5945 ( \6322 , \6320 , \6321 );
xor \U$5946 ( \6323 , \5813 , \5827 );
xor \U$5947 ( \6324 , \6323 , \5801 );
xor \U$5948 ( \6325 , \6322 , \6324 );
not \U$5949 ( \6326 , \1915 );
not \U$5950 ( \6327 , RIc226b60_23);
not \U$5951 ( \6328 , \2424 );
or \U$5952 ( \6329 , \6327 , \6328 );
nand \U$5953 ( \6330 , \2423 , \5637 );
nand \U$5954 ( \6331 , \6329 , \6330 );
not \U$5955 ( \6332 , \6331 );
or \U$5956 ( \6333 , \6326 , \6332 );
nand \U$5957 ( \6334 , \6038 , \1930 );
nand \U$5958 ( \6335 , \6333 , \6334 );
not \U$5959 ( \6336 , \6335 );
not \U$5960 ( \6337 , \6336 );
not \U$5961 ( \6338 , \2392 );
not \U$5962 ( \6339 , RIc226c50_21);
not \U$5963 ( \6340 , \2234 );
or \U$5964 ( \6341 , \6339 , \6340 );
nand \U$5965 ( \6342 , \2229 , \2383 );
nand \U$5966 ( \6343 , \6341 , \6342 );
not \U$5967 ( \6344 , \6343 );
or \U$5968 ( \6345 , \6338 , \6344 );
nand \U$5969 ( \6346 , \5951 , \2367 );
nand \U$5970 ( \6347 , \6345 , \6346 );
not \U$5971 ( \6348 , \6347 );
not \U$5972 ( \6349 , \6348 );
or \U$5973 ( \6350 , \6337 , \6349 );
not \U$5974 ( \6351 , \3629 );
not \U$5975 ( \6352 , RIc2266b0_33);
not \U$5976 ( \6353 , \1022 );
or \U$5977 ( \6354 , \6352 , \6353 );
not \U$5978 ( \6355 , RIc2266b0_33);
nand \U$5979 ( \6356 , \1455 , \6355 );
nand \U$5980 ( \6357 , \6354 , \6356 );
not \U$5981 ( \6358 , \6357 );
or \U$5982 ( \6359 , \6351 , \6358 );
nand \U$5983 ( \6360 , \6208 , \3631 );
nand \U$5984 ( \6361 , \6359 , \6360 );
nand \U$5985 ( \6362 , \6350 , \6361 );
nand \U$5986 ( \6363 , \6347 , \6335 );
nand \U$5987 ( \6364 , \6362 , \6363 );
not \U$5988 ( \6365 , \6364 );
not \U$5989 ( \6366 , \5135 );
not \U$5990 ( \6367 , \5966 );
or \U$5991 ( \6368 , \6366 , \6367 );
not \U$5992 ( \6369 , RIc2265c0_35);
not \U$5993 ( \6370 , \1706 );
or \U$5994 ( \6371 , \6369 , \6370 );
nand \U$5995 ( \6372 , \841 , \4376 );
nand \U$5996 ( \6373 , \6371 , \6372 );
nand \U$5997 ( \6374 , \6373 , \5741 );
nand \U$5998 ( \6375 , \6368 , \6374 );
not \U$5999 ( \6376 , \6375 );
not \U$6000 ( \6377 , \2697 );
not \U$6001 ( \6378 , RIc2267a0_31);
not \U$6002 ( \6379 , \1222 );
or \U$6003 ( \6380 , \6378 , \6379 );
nand \U$6004 ( \6381 , \3242 , \2705 );
nand \U$6005 ( \6382 , \6380 , \6381 );
not \U$6006 ( \6383 , \6382 );
or \U$6007 ( \6384 , \6377 , \6383 );
nand \U$6008 ( \6385 , \5939 , \3653 );
nand \U$6009 ( \6386 , \6384 , \6385 );
not \U$6010 ( \6387 , \6386 );
or \U$6011 ( \6388 , \6376 , \6387 );
not \U$6012 ( \6389 , \6386 );
not \U$6013 ( \6390 , \6389 );
not \U$6014 ( \6391 , \6375 );
not \U$6015 ( \6392 , \6391 );
or \U$6016 ( \6393 , \6390 , \6392 );
not \U$6017 ( \6394 , \2534 );
not \U$6018 ( \6395 , \6002 );
or \U$6019 ( \6396 , \6394 , \6395 );
not \U$6020 ( \6397 , RIc226d40_19);
not \U$6021 ( \6398 , \3835 );
or \U$6022 ( \6399 , \6397 , \6398 );
not \U$6023 ( \6400 , \5768 );
nand \U$6024 ( \6401 , \6400 , \3338 );
nand \U$6025 ( \6402 , \6399 , \6401 );
nand \U$6026 ( \6403 , \6402 , \2518 );
nand \U$6027 ( \6404 , \6396 , \6403 );
nand \U$6028 ( \6405 , \6393 , \6404 );
nand \U$6029 ( \6406 , \6388 , \6405 );
not \U$6030 ( \6407 , \6406 );
or \U$6031 ( \6408 , \6365 , \6407 );
or \U$6032 ( \6409 , \6406 , \6364 );
not \U$6033 ( \6410 , \5509 );
not \U$6034 ( \6411 , RIc2264d0_37);
not \U$6035 ( \6412 , \3071 );
or \U$6036 ( \6413 , \6411 , \6412 );
nand \U$6037 ( \6414 , \1073 , \5514 );
nand \U$6038 ( \6415 , \6413 , \6414 );
not \U$6039 ( \6416 , \6415 );
or \U$6040 ( \6417 , \6410 , \6416 );
nand \U$6041 ( \6418 , \5516 , \5519 );
nand \U$6042 ( \6419 , \6417 , \6418 );
not \U$6043 ( \6420 , \6419 );
not \U$6044 ( \6421 , \1340 );
not \U$6045 ( \6422 , \6274 );
or \U$6046 ( \6423 , \6421 , \6422 );
not \U$6047 ( \6424 , RIc2271f0_9);
not \U$6048 ( \6425 , \4501 );
not \U$6049 ( \6426 , \6425 );
or \U$6050 ( \6427 , \6424 , \6426 );
nand \U$6051 ( \6428 , \2105 , \1351 );
nand \U$6052 ( \6429 , \6427 , \6428 );
nand \U$6053 ( \6430 , \6429 , \1597 );
nand \U$6054 ( \6431 , \6423 , \6430 );
not \U$6055 ( \6432 , \6431 );
or \U$6056 ( \6433 , \6420 , \6432 );
or \U$6057 ( \6434 , \6431 , \6419 );
not \U$6058 ( \6435 , \1121 );
not \U$6059 ( \6436 , \6027 );
or \U$6060 ( \6437 , \6435 , \6436 );
not \U$6061 ( \6438 , RIc2272e0_7);
not \U$6062 ( \6439 , \3732 );
not \U$6063 ( \6440 , \6439 );
or \U$6064 ( \6441 , \6438 , \6440 );
nand \U$6065 ( \6442 , \3732 , \1139 );
nand \U$6066 ( \6443 , \6441 , \6442 );
nand \U$6067 ( \6444 , \6443 , \1118 );
nand \U$6068 ( \6445 , \6437 , \6444 );
nand \U$6069 ( \6446 , \6434 , \6445 );
nand \U$6070 ( \6447 , \6433 , \6446 );
nand \U$6071 ( \6448 , \6409 , \6447 );
nand \U$6072 ( \6449 , \6408 , \6448 );
and \U$6073 ( \6450 , \6325 , \6449 );
and \U$6074 ( \6451 , \6322 , \6324 );
or \U$6075 ( \6452 , \6450 , \6451 );
nand \U$6076 ( \6453 , \6267 , \6452 );
not \U$6077 ( \6454 , \6265 );
nand \U$6078 ( \6455 , \6454 , \6261 );
nand \U$6079 ( \6456 , \6453 , \6455 );
xor \U$6080 ( \6457 , \5866 , \5864 );
xor \U$6081 ( \6458 , \6457 , \5888 );
or \U$6082 ( \6459 , \6456 , \6458 );
xor \U$6083 ( \6460 , \5598 , \5596 );
xor \U$6084 ( \6461 , \6460 , \5605 );
nand \U$6085 ( \6462 , \6459 , \6461 );
nand \U$6086 ( \6463 , \6456 , \6458 );
nand \U$6087 ( \6464 , \6462 , \6463 );
not \U$6088 ( \6465 , \6464 );
xor \U$6089 ( \6466 , \6126 , \6135 );
xor \U$6090 ( \6467 , \6466 , \6114 );
xor \U$6091 ( \6468 , \6191 , \6201 );
xnor \U$6092 ( \6469 , \6468 , \6213 );
nand \U$6093 ( \6470 , \6467 , \6469 );
xor \U$6094 ( \6471 , \6021 , \6031 );
xor \U$6095 ( \6472 , \6471 , \6043 );
and \U$6096 ( \6473 , \6470 , \6472 );
nor \U$6097 ( \6474 , \6467 , \6469 );
nor \U$6098 ( \6475 , \6473 , \6474 );
not \U$6099 ( \6476 , \528 );
not \U$6100 ( \6477 , \4393 );
or \U$6101 ( \6478 , \6476 , \6477 );
not \U$6102 ( \6479 , \648 );
nand \U$6103 ( \6480 , \6478 , \6479 );
not \U$6104 ( \6481 , \6480 );
not \U$6105 ( \6482 , \528 );
nor \U$6106 ( \6483 , \6482 , \4087 );
nand \U$6107 ( \6484 , \4084 , \6483 );
nand \U$6108 ( \6485 , \6481 , \6484 );
nand \U$6109 ( \6486 , \649 , \652 );
not \U$6110 ( \6487 , \6486 );
and \U$6111 ( \6488 , \6485 , \6487 );
not \U$6112 ( \6489 , \6485 );
and \U$6113 ( \6490 , \6489 , \6486 );
nor \U$6114 ( \6491 , \6488 , \6490 );
buf \U$6115 ( \6492 , \6491 );
not \U$6116 ( \6493 , \6492 );
not \U$6117 ( \6494 , \6493 );
nand \U$6118 ( \6495 , \6494 , RIc2275b0_1);
xor \U$6119 ( \6496 , RIc2275b0_1, \6071 );
not \U$6120 ( \6497 , \6496 );
not \U$6121 ( \6498 , \6497 );
not \U$6122 ( \6499 , \855 );
and \U$6123 ( \6500 , \6498 , \6499 );
and \U$6124 ( \6501 , \6091 , \1579 );
nor \U$6125 ( \6502 , \6500 , \6501 );
xor \U$6126 ( \6503 , \6495 , \6502 );
not \U$6127 ( \6504 , \2354 );
not \U$6128 ( \6505 , \1905 );
and \U$6129 ( \6506 , \6504 , \6505 );
and \U$6130 ( \6507 , \2354 , \6107 );
nor \U$6131 ( \6508 , \6506 , \6507 );
not \U$6132 ( \6509 , \6508 );
not \U$6133 ( \6510 , \4599 );
and \U$6134 ( \6511 , \6509 , \6510 );
not \U$6135 ( \6512 , \2173 );
nor \U$6136 ( \6513 , \6512 , \6109 );
nor \U$6137 ( \6514 , \6511 , \6513 );
and \U$6138 ( \6515 , \6503 , \6514 );
and \U$6139 ( \6516 , \6495 , \6502 );
or \U$6140 ( \6517 , \6515 , \6516 );
not \U$6141 ( \6518 , \6517 );
not \U$6142 ( \6519 , \2086 );
not \U$6143 ( \6520 , \5978 );
or \U$6144 ( \6521 , \6519 , \6520 );
and \U$6145 ( \6522 , RIc226890_29, \1531 );
not \U$6146 ( \6523 , RIc226890_29);
and \U$6147 ( \6524 , \6523 , \1532 );
or \U$6148 ( \6525 , \6522 , \6524 );
nand \U$6149 ( \6526 , \6525 , \2078 );
nand \U$6150 ( \6527 , \6521 , \6526 );
not \U$6151 ( \6528 , \2358 );
not \U$6152 ( \6529 , \6187 );
or \U$6153 ( \6530 , \6528 , \6529 );
not \U$6154 ( \6531 , RIc226f20_15);
not \U$6155 ( \6532 , \3313 );
or \U$6156 ( \6533 , \6531 , \6532 );
not \U$6157 ( \6534 , \2476 );
nand \U$6158 ( \6535 , \6534 , \2351 );
nand \U$6159 ( \6536 , \6533 , \6535 );
nand \U$6160 ( \6537 , \6536 , \2320 );
nand \U$6161 ( \6538 , \6530 , \6537 );
or \U$6162 ( \6539 , \6527 , \6538 );
not \U$6163 ( \6540 , RIc226e30_17);
not \U$6164 ( \6541 , \2587 );
or \U$6165 ( \6542 , \6540 , \6541 );
nand \U$6166 ( \6543 , \2593 , \1952 );
nand \U$6167 ( \6544 , \6542 , \6543 );
and \U$6168 ( \6545 , \6544 , \1945 );
and \U$6169 ( \6546 , \5989 , \1963 );
nor \U$6170 ( \6547 , \6545 , \6546 );
not \U$6171 ( \6548 , \6547 );
nand \U$6172 ( \6549 , \6539 , \6548 );
nand \U$6173 ( \6550 , \6538 , \6527 );
and \U$6174 ( \6551 , \6549 , \6550 );
not \U$6175 ( \6552 , \6551 );
or \U$6176 ( \6553 , \6518 , \6552 );
xor \U$6177 ( \6554 , \6072 , \6095 );
xnor \U$6178 ( \6555 , \6554 , \6097 );
not \U$6179 ( \6556 , \6555 );
nand \U$6180 ( \6557 , \6553 , \6556 );
not \U$6181 ( \6558 , \6551 );
not \U$6182 ( \6559 , \6517 );
nand \U$6183 ( \6560 , \6558 , \6559 );
and \U$6184 ( \6561 , \6557 , \6560 );
nand \U$6185 ( \6562 , \6475 , \6561 );
not \U$6186 ( \6563 , \1311 );
not \U$6187 ( \6564 , \6122 );
or \U$6188 ( \6565 , \6563 , \6564 );
not \U$6189 ( \6566 , RIc227100_11);
not \U$6190 ( \6567 , \2043 );
or \U$6191 ( \6568 , \6566 , \6567 );
nand \U$6192 ( \6569 , \2732 , \1685 );
nand \U$6193 ( \6570 , \6568 , \6569 );
nand \U$6194 ( \6571 , \6570 , \1307 );
nand \U$6195 ( \6572 , \6565 , \6571 );
not \U$6196 ( \6573 , \2154 );
not \U$6197 ( \6574 , \6197 );
or \U$6198 ( \6575 , \6573 , \6574 );
not \U$6199 ( \6576 , RIc226980_27);
not \U$6200 ( \6577 , \1488 );
or \U$6201 ( \6578 , \6576 , \6577 );
nand \U$6202 ( \6579 , \2609 , \2133 );
nand \U$6203 ( \6580 , \6578 , \6579 );
nand \U$6204 ( \6581 , \6580 , \2138 );
nand \U$6205 ( \6582 , \6575 , \6581 );
or \U$6206 ( \6583 , \6572 , \6582 );
not \U$6207 ( \6584 , \1682 );
not \U$6208 ( \6585 , \6130 );
not \U$6209 ( \6586 , \6585 );
or \U$6210 ( \6587 , \6584 , \6586 );
and \U$6211 ( \6588 , \2672 , RIc227010_13);
not \U$6212 ( \6589 , \2672 );
and \U$6213 ( \6590 , \6589 , \2427 );
or \U$6214 ( \6591 , \6588 , \6590 );
nand \U$6215 ( \6592 , \6591 , \1680 );
nand \U$6216 ( \6593 , \6587 , \6592 );
nand \U$6217 ( \6594 , \6583 , \6593 );
nand \U$6218 ( \6595 , \6572 , \6582 );
nand \U$6219 ( \6596 , \6594 , \6595 );
not \U$6220 ( \6597 , \6596 );
xor \U$6221 ( \6598 , \5970 , \5958 );
and \U$6222 ( \6599 , \6598 , \5954 );
not \U$6223 ( \6600 , \6598 );
and \U$6224 ( \6601 , \6600 , \5953 );
nor \U$6225 ( \6602 , \6599 , \6601 );
nand \U$6226 ( \6603 , \6597 , \6602 );
not \U$6227 ( \6604 , \6603 );
xor \U$6228 ( \6605 , \6007 , \5993 );
xor \U$6229 ( \6606 , \6605 , \5982 );
not \U$6230 ( \6607 , \6606 );
or \U$6231 ( \6608 , \6604 , \6607 );
not \U$6232 ( \6609 , \6602 );
nand \U$6233 ( \6610 , \6609 , \6596 );
nand \U$6234 ( \6611 , \6608 , \6610 );
and \U$6235 ( \6612 , \6562 , \6611 );
nor \U$6236 ( \6613 , \6475 , \6561 );
nor \U$6237 ( \6614 , \6612 , \6613 );
not \U$6238 ( \6615 , \6614 );
not \U$6239 ( \6616 , \6141 );
not \U$6240 ( \6617 , \6616 );
not \U$6241 ( \6618 , \6050 );
or \U$6242 ( \6619 , \6617 , \6618 );
nand \U$6243 ( \6620 , \6049 , \6141 );
nand \U$6244 ( \6621 , \6619 , \6620 );
not \U$6245 ( \6622 , \6053 );
and \U$6246 ( \6623 , \6621 , \6622 );
not \U$6247 ( \6624 , \6621 );
and \U$6248 ( \6625 , \6624 , \6053 );
nor \U$6249 ( \6626 , \6623 , \6625 );
not \U$6250 ( \6627 , \6626 );
or \U$6251 ( \6628 , \6615 , \6627 );
xor \U$6252 ( \6629 , \5972 , \6010 );
xor \U$6253 ( \6630 , \6629 , \6046 );
not \U$6254 ( \6631 , \6630 );
not \U$6255 ( \6632 , \6225 );
not \U$6256 ( \6633 , \6216 );
and \U$6257 ( \6634 , \6632 , \6633 );
and \U$6258 ( \6635 , \6225 , \6216 );
nor \U$6259 ( \6636 , \6634 , \6635 );
not \U$6260 ( \6637 , \6636 );
not \U$6261 ( \6638 , \6180 );
and \U$6262 ( \6639 , \6637 , \6638 );
and \U$6263 ( \6640 , \6636 , \6180 );
nor \U$6264 ( \6641 , \6639 , \6640 );
not \U$6265 ( \6642 , \6641 );
or \U$6266 ( \6643 , \6631 , \6642 );
xor \U$6267 ( \6644 , \6099 , \6101 );
xor \U$6268 ( \6645 , \6644 , \6138 );
nand \U$6269 ( \6646 , \6643 , \6645 );
not \U$6270 ( \6647 , \6641 );
not \U$6271 ( \6648 , \6630 );
nand \U$6272 ( \6649 , \6647 , \6648 );
nand \U$6273 ( \6650 , \6646 , \6649 );
nand \U$6274 ( \6651 , \6628 , \6650 );
not \U$6275 ( \6652 , \6626 );
not \U$6276 ( \6653 , \6614 );
nand \U$6277 ( \6654 , \6652 , \6653 );
and \U$6278 ( \6655 , \6651 , \6654 );
and \U$6279 ( \6656 , \6232 , \6143 );
not \U$6280 ( \6657 , \6232 );
and \U$6281 ( \6658 , \6657 , \6151 );
nor \U$6282 ( \6659 , \6656 , \6658 );
not \U$6283 ( \6660 , \6659 );
not \U$6284 ( \6661 , \6147 );
not \U$6285 ( \6662 , \6661 );
and \U$6286 ( \6663 , \6660 , \6662 );
and \U$6287 ( \6664 , \6659 , \6661 );
nor \U$6288 ( \6665 , \6663 , \6664 );
nand \U$6289 ( \6666 , \6655 , \6665 );
xor \U$6290 ( \6667 , \6168 , \6175 );
xnor \U$6291 ( \6668 , \6667 , \6230 );
not \U$6292 ( \6669 , \6668 );
xor \U$6293 ( \6670 , \6261 , \6265 );
xor \U$6294 ( \6671 , \6670 , \6452 );
not \U$6295 ( \6672 , \6671 );
or \U$6296 ( \6673 , \6669 , \6672 );
xnor \U$6297 ( \6674 , \6155 , \6166 );
not \U$6298 ( \6675 , \6161 );
and \U$6299 ( \6676 , \6674 , \6675 );
not \U$6300 ( \6677 , \6674 );
and \U$6301 ( \6678 , \6677 , \6161 );
nor \U$6302 ( \6679 , \6676 , \6678 );
not \U$6303 ( \6680 , \6679 );
xor \U$6304 ( \6681 , \6322 , \6324 );
xor \U$6305 ( \6682 , \6681 , \6449 );
not \U$6306 ( \6683 , \6682 );
or \U$6307 ( \6684 , \6680 , \6683 );
or \U$6308 ( \6685 , \6682 , \6679 );
xor \U$6309 ( \6686 , \6268 , \6278 );
xor \U$6310 ( \6687 , \6686 , \6319 );
not \U$6311 ( \6688 , \6313 );
buf \U$6312 ( \6689 , \6688 );
not \U$6313 ( \6690 , \6689 );
not \U$6314 ( \6691 , RIc2263e0_39);
not \U$6315 ( \6692 , \932 );
or \U$6316 ( \6693 , \6691 , \6692 );
not \U$6317 ( \6694 , RIc2263e0_39);
nand \U$6318 ( \6695 , \931 , \6694 );
nand \U$6319 ( \6696 , \6693 , \6695 );
not \U$6320 ( \6697 , \6696 );
or \U$6321 ( \6698 , \6690 , \6697 );
nand \U$6322 ( \6699 , \6307 , RIc2263e0_39);
nand \U$6323 ( \6700 , \6698 , \6699 );
not \U$6324 ( \6701 , \6700 );
not \U$6325 ( \6702 , \527 );
not \U$6326 ( \6703 , \6702 );
not \U$6327 ( \6704 , \4111 );
or \U$6328 ( \6705 , \6703 , \6704 );
nand \U$6329 ( \6706 , RIc224568_104, RIc22a7d8_168);
nand \U$6330 ( \6707 , \6705 , \6706 );
not \U$6331 ( \6708 , \6707 );
nor \U$6332 ( \6709 , \4087 , \527 );
nand \U$6333 ( \6710 , \4084 , \6709 );
nand \U$6334 ( \6711 , \6708 , \6710 );
nand \U$6335 ( \6712 , \644 , \647 );
not \U$6336 ( \6713 , \6712 );
and \U$6337 ( \6714 , \6711 , \6713 );
not \U$6338 ( \6715 , \6711 );
and \U$6339 ( \6716 , \6715 , \6712 );
nor \U$6340 ( \6717 , \6714 , \6716 );
buf \U$6341 ( \6718 , \6717 );
not \U$6342 ( \6719 , \6718 );
not \U$6343 ( \6720 , \6719 );
and \U$6344 ( \6721 , \6720 , RIc2275b0_1);
not \U$6345 ( \6722 , \6721 );
not \U$6346 ( \6723 , \1082 );
not \U$6347 ( \6724 , \6297 );
or \U$6348 ( \6725 , \6723 , \6724 );
buf \U$6349 ( \6726 , \5663 );
and \U$6350 ( \6727 , \6726 , \1027 );
not \U$6351 ( \6728 , \6726 );
and \U$6352 ( \6729 , \6728 , RIc2274c0_3);
or \U$6353 ( \6730 , \6727 , \6729 );
nand \U$6354 ( \6731 , \6730 , \1040 );
nand \U$6355 ( \6732 , \6725 , \6731 );
not \U$6356 ( \6733 , \6732 );
or \U$6357 ( \6734 , \6722 , \6733 );
or \U$6358 ( \6735 , \6732 , \6721 );
not \U$6359 ( \6736 , \951 );
not \U$6360 ( \6737 , \946 );
not \U$6361 ( \6738 , \6079 );
or \U$6362 ( \6739 , \6737 , \6738 );
not \U$6363 ( \6740 , \4407 );
nand \U$6364 ( \6741 , \6740 , RIc2273d0_5);
nand \U$6365 ( \6742 , \6739 , \6741 );
not \U$6366 ( \6743 , \6742 );
or \U$6367 ( \6744 , \6736 , \6743 );
nand \U$6368 ( \6745 , \6287 , \954 );
nand \U$6369 ( \6746 , \6744 , \6745 );
nand \U$6370 ( \6747 , \6735 , \6746 );
nand \U$6371 ( \6748 , \6734 , \6747 );
not \U$6372 ( \6749 , \6748 );
or \U$6373 ( \6750 , \6701 , \6749 );
not \U$6374 ( \6751 , \6700 );
not \U$6375 ( \6752 , \6751 );
not \U$6376 ( \6753 , \6748 );
not \U$6377 ( \6754 , \6753 );
or \U$6378 ( \6755 , \6752 , \6754 );
not \U$6379 ( \6756 , \2086 );
not \U$6380 ( \6757 , \6525 );
or \U$6381 ( \6758 , \6756 , \6757 );
and \U$6382 ( \6759 , RIc226890_29, \3438 );
not \U$6383 ( \6760 , RIc226890_29);
and \U$6384 ( \6761 , \6760 , \1332 );
or \U$6385 ( \6762 , \6759 , \6761 );
nand \U$6386 ( \6763 , \6762 , \2078 );
nand \U$6387 ( \6764 , \6758 , \6763 );
not \U$6388 ( \6765 , \6764 );
not \U$6389 ( \6766 , \2534 );
not \U$6390 ( \6767 , \6402 );
or \U$6391 ( \6768 , \6766 , \6767 );
not \U$6392 ( \6769 , RIc226d40_19);
not \U$6393 ( \6770 , \3509 );
or \U$6394 ( \6771 , \6769 , \6770 );
nand \U$6395 ( \6772 , \3508 , \3338 );
nand \U$6396 ( \6773 , \6771 , \6772 );
nand \U$6397 ( \6774 , \6773 , \2518 );
nand \U$6398 ( \6775 , \6768 , \6774 );
not \U$6399 ( \6776 , \6775 );
or \U$6400 ( \6777 , \6765 , \6776 );
or \U$6401 ( \6778 , \6775 , \6764 );
not \U$6402 ( \6779 , \5135 );
not \U$6403 ( \6780 , \6373 );
or \U$6404 ( \6781 , \6779 , \6780 );
not \U$6405 ( \6782 , RIc2265c0_35);
not \U$6406 ( \6783 , \1559 );
or \U$6407 ( \6784 , \6782 , \6783 );
nand \U$6408 ( \6785 , \984 , \3620 );
nand \U$6409 ( \6786 , \6784 , \6785 );
nand \U$6410 ( \6787 , \6786 , \5741 );
nand \U$6411 ( \6788 , \6781 , \6787 );
nand \U$6412 ( \6789 , \6778 , \6788 );
nand \U$6413 ( \6790 , \6777 , \6789 );
nand \U$6414 ( \6791 , \6755 , \6790 );
nand \U$6415 ( \6792 , \6750 , \6791 );
or \U$6416 ( \6793 , \6687 , \6792 );
not \U$6417 ( \6794 , \5519 );
not \U$6418 ( \6795 , \6415 );
or \U$6419 ( \6796 , \6794 , \6795 );
not \U$6420 ( \6797 , RIc2264d0_37);
not \U$6421 ( \6798 , \2865 );
or \U$6422 ( \6799 , \6797 , \6798 );
nand \U$6423 ( \6800 , \889 , \4371 );
nand \U$6424 ( \6801 , \6799 , \6800 );
nand \U$6425 ( \6802 , \6801 , \5509 );
nand \U$6426 ( \6803 , \6796 , \6802 );
not \U$6427 ( \6804 , \6803 );
not \U$6428 ( \6805 , \6804 );
not \U$6429 ( \6806 , \1930 );
not \U$6430 ( \6807 , \6331 );
or \U$6431 ( \6808 , \6806 , \6807 );
not \U$6432 ( \6809 , RIc226b60_23);
not \U$6433 ( \6810 , \2834 );
or \U$6434 ( \6811 , \6809 , \6810 );
nand \U$6435 ( \6812 , \5949 , \5637 );
nand \U$6436 ( \6813 , \6811 , \6812 );
nand \U$6437 ( \6814 , \6813 , \1915 );
nand \U$6438 ( \6815 , \6808 , \6814 );
not \U$6439 ( \6816 , \6815 );
not \U$6440 ( \6817 , \6816 );
or \U$6441 ( \6818 , \6805 , \6817 );
not \U$6442 ( \6819 , \1121 );
not \U$6443 ( \6820 , \6443 );
or \U$6444 ( \6821 , \6819 , \6820 );
not \U$6445 ( \6822 , RIc2272e0_7);
not \U$6446 ( \6823 , \4046 );
or \U$6447 ( \6824 , \6822 , \6823 );
nand \U$6448 ( \6825 , \3641 , \940 );
nand \U$6449 ( \6826 , \6824 , \6825 );
nand \U$6450 ( \6827 , \6826 , \1118 );
nand \U$6451 ( \6828 , \6821 , \6827 );
nand \U$6452 ( \6829 , \6818 , \6828 );
nand \U$6453 ( \6830 , \6815 , \6803 );
nand \U$6454 ( \6831 , \6829 , \6830 );
not \U$6455 ( \6832 , \6831 );
not \U$6456 ( \6833 , \1945 );
not \U$6457 ( \6834 , RIc226e30_17);
not \U$6458 ( \6835 , \4803 );
or \U$6459 ( \6836 , \6834 , \6835 );
nand \U$6460 ( \6837 , \3450 , \1952 );
nand \U$6461 ( \6838 , \6836 , \6837 );
not \U$6462 ( \6839 , \6838 );
or \U$6463 ( \6840 , \6833 , \6839 );
nand \U$6464 ( \6841 , \6544 , \1963 );
nand \U$6465 ( \6842 , \6840 , \6841 );
not \U$6466 ( \6843 , \6842 );
not \U$6467 ( \6844 , \2156 );
not \U$6468 ( \6845 , \6580 );
or \U$6469 ( \6846 , \6844 , \6845 );
and \U$6470 ( \6847 , \2150 , \1730 );
not \U$6471 ( \6848 , \2150 );
and \U$6472 ( \6849 , \6848 , \4178 );
nor \U$6473 ( \6850 , \6847 , \6849 );
not \U$6474 ( \6851 , \6850 );
nand \U$6475 ( \6852 , \6851 , \2138 );
nand \U$6476 ( \6853 , \6846 , \6852 );
not \U$6477 ( \6854 , \6853 );
nand \U$6478 ( \6855 , \6843 , \6854 );
not \U$6479 ( \6856 , \6855 );
not \U$6480 ( \6857 , \2358 );
not \U$6481 ( \6858 , \6536 );
or \U$6482 ( \6859 , \6857 , \6858 );
not \U$6483 ( \6860 , RIc226f20_15);
not \U$6484 ( \6861 , \3023 );
or \U$6485 ( \6862 , \6860 , \6861 );
nand \U$6486 ( \6863 , \2504 , \1674 );
nand \U$6487 ( \6864 , \6862 , \6863 );
nand \U$6488 ( \6865 , \6864 , \2320 );
nand \U$6489 ( \6866 , \6859 , \6865 );
not \U$6490 ( \6867 , \6866 );
or \U$6491 ( \6868 , \6856 , \6867 );
nand \U$6492 ( \6869 , \6853 , \6842 );
nand \U$6493 ( \6870 , \6868 , \6869 );
not \U$6494 ( \6871 , \6870 );
or \U$6495 ( \6872 , \6832 , \6871 );
or \U$6496 ( \6873 , \6870 , \6831 );
not \U$6497 ( \6874 , \2367 );
not \U$6498 ( \6875 , \6343 );
or \U$6499 ( \6876 , \6874 , \6875 );
not \U$6500 ( \6877 , RIc226c50_21);
not \U$6501 ( \6878 , \2258 );
or \U$6502 ( \6879 , \6877 , \6878 );
nand \U$6503 ( \6880 , \2261 , \2383 );
nand \U$6504 ( \6881 , \6879 , \6880 );
nand \U$6505 ( \6882 , \6881 , \2392 );
nand \U$6506 ( \6883 , \6876 , \6882 );
not \U$6507 ( \6884 , \3631 );
not \U$6508 ( \6885 , \6357 );
or \U$6509 ( \6886 , \6884 , \6885 );
not \U$6510 ( \6887 , RIc2266b0_33);
not \U$6511 ( \6888 , \1171 );
or \U$6512 ( \6889 , \6887 , \6888 );
not \U$6513 ( \6890 , RIc2266b0_33);
nand \U$6514 ( \6891 , \1228 , \6890 );
nand \U$6515 ( \6892 , \6889 , \6891 );
nand \U$6516 ( \6893 , \6892 , \3629 );
nand \U$6517 ( \6894 , \6886 , \6893 );
xor \U$6518 ( \6895 , \6883 , \6894 );
not \U$6519 ( \6896 , \3653 );
not \U$6520 ( \6897 , \6382 );
or \U$6521 ( \6898 , \6896 , \6897 );
not \U$6522 ( \6899 , RIc2267a0_31);
not \U$6523 ( \6900 , \3497 );
or \U$6524 ( \6901 , \6899 , \6900 );
not \U$6525 ( \6902 , RIc2267a0_31);
nand \U$6526 ( \6903 , \3500 , \6902 );
nand \U$6527 ( \6904 , \6901 , \6903 );
nand \U$6528 ( \6905 , \6904 , \2697 );
nand \U$6529 ( \6906 , \6898 , \6905 );
and \U$6530 ( \6907 , \6895 , \6906 );
and \U$6531 ( \6908 , \6883 , \6894 );
or \U$6532 ( \6909 , \6907 , \6908 );
nand \U$6533 ( \6910 , \6873 , \6909 );
nand \U$6534 ( \6911 , \6872 , \6910 );
nand \U$6535 ( \6912 , \6793 , \6911 );
nand \U$6536 ( \6913 , \6792 , \6687 );
nand \U$6537 ( \6914 , \6912 , \6913 );
nand \U$6538 ( \6915 , \6685 , \6914 );
nand \U$6539 ( \6916 , \6684 , \6915 );
nand \U$6540 ( \6917 , \6673 , \6916 );
not \U$6541 ( \6918 , \6668 );
not \U$6542 ( \6919 , \6671 );
nand \U$6543 ( \6920 , \6918 , \6919 );
nand \U$6544 ( \6921 , \6917 , \6920 );
and \U$6545 ( \6922 , \6666 , \6921 );
nor \U$6546 ( \6923 , \6655 , \6665 );
nor \U$6547 ( \6924 , \6922 , \6923 );
not \U$6548 ( \6925 , \6924 );
not \U$6549 ( \6926 , \6925 );
or \U$6550 ( \6927 , \6465 , \6926 );
not \U$6551 ( \6928 , \6234 );
not \U$6552 ( \6929 , \5933 );
or \U$6553 ( \6930 , \6928 , \6929 );
nand \U$6554 ( \6931 , \5932 , \6235 );
nand \U$6555 ( \6932 , \6930 , \6931 );
xor \U$6556 ( \6933 , \6932 , \5929 );
not \U$6557 ( \6934 , \6464 );
nand \U$6558 ( \6935 , \6934 , \6924 );
nand \U$6559 ( \6936 , \6933 , \6935 );
nand \U$6560 ( \6937 , \6927 , \6936 );
or \U$6561 ( \6938 , \6251 , \6937 );
nand \U$6562 ( \6939 , \6245 , \6938 );
nor \U$6563 ( \6940 , \5914 , \6939 );
xor \U$6564 ( \6941 , \4280 , \4646 );
xnor \U$6565 ( \6942 , \6941 , \4278 );
xor \U$6566 ( \6943 , \5113 , \5115 );
and \U$6567 ( \6944 , \6943 , \5449 );
and \U$6568 ( \6945 , \5113 , \5115 );
or \U$6569 ( \6946 , \6944 , \6945 );
nand \U$6570 ( \6947 , \6942 , \6946 );
nand \U$6571 ( \6948 , \6940 , \6947 );
nor \U$6572 ( \6949 , \5110 , \6948 );
not \U$6573 ( \6950 , \2358 );
and \U$6574 ( \6951 , \2301 , \1022 );
not \U$6575 ( \6952 , \2301 );
and \U$6576 ( \6953 , \6952 , \1127 );
nor \U$6577 ( \6954 , \6951 , \6953 );
not \U$6578 ( \6955 , \6954 );
or \U$6579 ( \6956 , \6950 , \6955 );
and \U$6580 ( \6957 , RIc226f20_15, \1404 );
not \U$6581 ( \6958 , RIc226f20_15);
and \U$6582 ( \6959 , \6958 , \1403 );
or \U$6583 ( \6960 , \6957 , \6959 );
not \U$6584 ( \6961 , \6960 );
or \U$6585 ( \6962 , \6961 , \2321 );
nand \U$6586 ( \6963 , \6956 , \6962 );
not \U$6587 ( \6964 , \1121 );
and \U$6588 ( \6965 , \2354 , RIc2272e0_7);
not \U$6589 ( \6966 , \2354 );
and \U$6590 ( \6967 , \6966 , \1139 );
nor \U$6591 ( \6968 , \6965 , \6967 );
not \U$6592 ( \6969 , \6968 );
or \U$6593 ( \6970 , \6964 , \6969 );
and \U$6594 ( \6971 , \2774 , RIc2272e0_7);
and \U$6595 ( \6972 , \2306 , \940 );
nor \U$6596 ( \6973 , \6971 , \6972 );
or \U$6597 ( \6974 , \6973 , \1117 );
nand \U$6598 ( \6975 , \6970 , \6974 );
xor \U$6599 ( \6976 , \6963 , \6975 );
not \U$6600 ( \6977 , \2534 );
not \U$6601 ( \6978 , RIc226d40_19);
not \U$6602 ( \6979 , \1074 );
or \U$6603 ( \6980 , \6978 , \6979 );
nand \U$6604 ( \6981 , \1073 , \1941 );
nand \U$6605 ( \6982 , \6980 , \6981 );
not \U$6606 ( \6983 , \6982 );
or \U$6607 ( \6984 , \6977 , \6983 );
and \U$6608 ( \6985 , \889 , RIc226d40_19);
not \U$6609 ( \6986 , \889 );
and \U$6610 ( \6987 , \6986 , \2523 );
nor \U$6611 ( \6988 , \6985 , \6987 );
not \U$6612 ( \6989 , \6988 );
or \U$6613 ( \6990 , \6989 , \5700 );
nand \U$6614 ( \6991 , \6984 , \6990 );
xor \U$6615 ( \6992 , \6976 , \6991 );
not \U$6616 ( \6993 , \1082 );
and \U$6617 ( \6994 , \2235 , RIc2274c0_3);
not \U$6618 ( \6995 , \2235 );
and \U$6619 ( \6996 , \6995 , \1027 );
nor \U$6620 ( \6997 , \6994 , \6996 );
not \U$6621 ( \6998 , \6997 );
or \U$6622 ( \6999 , \6993 , \6998 );
not \U$6623 ( \7000 , RIc2274c0_3);
not \U$6624 ( \7001 , \2258 );
or \U$6625 ( \7002 , \7000 , \7001 );
nand \U$6626 ( \7003 , \2261 , \1078 );
nand \U$6627 ( \7004 , \7002 , \7003 );
not \U$6628 ( \7005 , \7004 );
or \U$6629 ( \7006 , \7005 , \1041 );
nand \U$6630 ( \7007 , \6999 , \7006 );
not \U$6631 ( \7008 , \954 );
not \U$6632 ( \7009 , \3348 );
and \U$6633 ( \7010 , \7009 , RIc2273d0_5);
not \U$6634 ( \7011 , \7009 );
and \U$6635 ( \7012 , \7011 , \946 );
nor \U$6636 ( \7013 , \7010 , \7012 );
not \U$6637 ( \7014 , \7013 );
or \U$6638 ( \7015 , \7008 , \7014 );
and \U$6639 ( \7016 , \2834 , RIc2273d0_5);
and \U$6640 ( \7017 , \2837 , \935 );
nor \U$6641 ( \7018 , \7016 , \7017 );
or \U$6642 ( \7019 , \7018 , \952 );
nand \U$6643 ( \7020 , \7015 , \7019 );
xor \U$6644 ( \7021 , \7007 , \7020 );
and \U$6645 ( \7022 , \1393 , RIc227010_13);
and \U$6646 ( \7023 , \1396 , \1296 );
nor \U$6647 ( \7024 , \7022 , \7023 );
or \U$6648 ( \7025 , \7024 , \1679 );
and \U$6649 ( \7026 , \1442 , RIc227010_13);
and \U$6650 ( \7027 , \1223 , \1296 );
nor \U$6651 ( \7028 , \7026 , \7027 );
or \U$6652 ( \7029 , \7028 , \1757 );
nand \U$6653 ( \7030 , \7025 , \7029 );
xor \U$6654 ( \7031 , \7021 , \7030 );
xor \U$6655 ( \7032 , \6992 , \7031 );
and \U$6656 ( \7033 , \5637 , \931 );
not \U$6657 ( \7034 , \5637 );
and \U$6658 ( \7035 , \7034 , \932 );
nor \U$6659 ( \7036 , \7033 , \7035 );
or \U$6660 ( \7037 , \7036 , \5643 );
not \U$6661 ( \7038 , \1930 );
or \U$6662 ( \7039 , \7038 , \1911 );
nand \U$6663 ( \7040 , \7037 , \7039 );
not \U$6664 ( \7041 , RIc227100_11);
not \U$6665 ( \7042 , \1488 );
or \U$6666 ( \7043 , \7041 , \7042 );
nand \U$6667 ( \7044 , \3299 , \1291 );
nand \U$6668 ( \7045 , \7043 , \7044 );
not \U$6669 ( \7046 , \7045 );
or \U$6670 ( \7047 , \7046 , \1308 );
and \U$6671 ( \7048 , \1949 , RIc227100_11);
and \U$6672 ( \7049 , \4778 , \1302 );
nor \U$6673 ( \7050 , \7048 , \7049 );
or \U$6674 ( \7051 , \7050 , \1312 );
nand \U$6675 ( \7052 , \7047 , \7051 );
xor \U$6676 ( \7053 , \7040 , \7052 );
not \U$6677 ( \7054 , \951 );
and \U$6678 ( \7055 , \2261 , RIc2273d0_5);
not \U$6679 ( \7056 , \2261 );
and \U$6680 ( \7057 , \7056 , \935 );
nor \U$6681 ( \7058 , \7055 , \7057 );
not \U$6682 ( \7059 , \7058 );
or \U$6683 ( \7060 , \7054 , \7059 );
and \U$6684 ( \7061 , \2229 , RIc2273d0_5);
not \U$6685 ( \7062 , \2229 );
and \U$6686 ( \7063 , \7062 , \946 );
nor \U$6687 ( \7064 , \7061 , \7063 );
nand \U$6688 ( \7065 , \7064 , \954 );
nand \U$6689 ( \7066 , \7060 , \7065 );
not \U$6690 ( \7067 , RIc226f20_15);
not \U$6691 ( \7068 , \2874 );
or \U$6692 ( \7069 , \7067 , \7068 );
nand \U$6693 ( \7070 , \1396 , \1674 );
nand \U$6694 ( \7071 , \7069 , \7070 );
not \U$6695 ( \7072 , \7071 );
or \U$6696 ( \7073 , \7072 , \2321 );
and \U$6697 ( \7074 , \1674 , \1442 );
not \U$6698 ( \7075 , \1674 );
and \U$6699 ( \7076 , \7075 , \1223 );
nor \U$6700 ( \7077 , \7074 , \7076 );
not \U$6701 ( \7078 , \7077 );
or \U$6702 ( \7079 , \7078 , \3305 );
nand \U$6703 ( \7080 , \7073 , \7079 );
xor \U$6704 ( \7081 , \7066 , \7080 );
and \U$6705 ( \7082 , \2837 , RIc2272e0_7);
not \U$6706 ( \7083 , \2837 );
and \U$6707 ( \7084 , \7083 , \1423 );
nor \U$6708 ( \7085 , \7082 , \7084 );
not \U$6709 ( \7086 , \7085 );
or \U$6710 ( \7087 , \7086 , \1117 );
and \U$6711 ( \7088 , \3348 , RIc2272e0_7);
and \U$6712 ( \7089 , \7009 , \1423 );
nor \U$6713 ( \7090 , \7088 , \7089 );
or \U$6714 ( \7091 , \7090 , \1431 );
nand \U$6715 ( \7092 , \7087 , \7091 );
and \U$6716 ( \7093 , \7081 , \7092 );
and \U$6717 ( \7094 , \7066 , \7080 );
or \U$6718 ( \7095 , \7093 , \7094 );
and \U$6719 ( \7096 , \7053 , \7095 );
and \U$6720 ( \7097 , \7040 , \7052 );
or \U$6721 ( \7098 , \7096 , \7097 );
xor \U$6722 ( \7099 , \7032 , \7098 );
not \U$6723 ( \7100 , \1597 );
not \U$6724 ( \7101 , RIc2271f0_9);
not \U$6725 ( \7102 , \2355 );
or \U$6726 ( \7103 , \7101 , \7102 );
nand \U$6727 ( \7104 , \2348 , \1351 );
nand \U$6728 ( \7105 , \7103 , \7104 );
not \U$6729 ( \7106 , \7105 );
or \U$6730 ( \7107 , \7100 , \7106 );
not \U$6731 ( \7108 , RIc2271f0_9);
not \U$6732 ( \7109 , \2616 );
or \U$6733 ( \7110 , \7108 , \7109 );
not \U$6734 ( \7111 , \2616 );
nand \U$6735 ( \7112 , \7111 , \1342 );
nand \U$6736 ( \7113 , \7110 , \7112 );
nand \U$6737 ( \7114 , \7113 , \1340 );
nand \U$6738 ( \7115 , \7107 , \7114 );
not \U$6739 ( \7116 , \2320 );
not \U$6740 ( \7117 , \7077 );
or \U$6741 ( \7118 , \7116 , \7117 );
nand \U$6742 ( \7119 , \6960 , \2358 );
nand \U$6743 ( \7120 , \7118 , \7119 );
xor \U$6744 ( \7121 , \7115 , \7120 );
or \U$6745 ( \7122 , \7090 , \1117 );
or \U$6746 ( \7123 , \6973 , \1431 );
nand \U$6747 ( \7124 , \7122 , \7123 );
and \U$6748 ( \7125 , \7121 , \7124 );
and \U$6749 ( \7126 , \7115 , \7120 );
or \U$6750 ( \7127 , \7125 , \7126 );
and \U$6751 ( \7128 , \2593 , RIc2275b0_1);
not \U$6752 ( \7129 , \1579 );
xor \U$6753 ( \7130 , RIc2275b0_1, \1991 );
not \U$6754 ( \7131 , \7130 );
or \U$6755 ( \7132 , \7129 , \7131 );
xor \U$6756 ( \7133 , RIc2275b0_1, \2018 );
nand \U$6757 ( \7134 , \7133 , \854 );
nand \U$6758 ( \7135 , \7132 , \7134 );
xor \U$6759 ( \7136 , \7128 , \7135 );
and \U$6760 ( \7137 , \986 , RIc226e30_17);
and \U$6761 ( \7138 , \985 , \1960 );
nor \U$6762 ( \7139 , \7137 , \7138 );
not \U$6763 ( \7140 , \1945 );
or \U$6764 ( \7141 , \7139 , \7140 );
and \U$6765 ( \7142 , \842 , RIc226e30_17);
and \U$6766 ( \7143 , \841 , \1960 );
nor \U$6767 ( \7144 , \7142 , \7143 );
not \U$6768 ( \7145 , \1963 );
or \U$6769 ( \7146 , \7144 , \7145 );
nand \U$6770 ( \7147 , \7141 , \7146 );
xor \U$6771 ( \7148 , \7136 , \7147 );
xor \U$6772 ( \7149 , \7127 , \7148 );
and \U$6773 ( \7150 , RIc226c50_21, \931 );
not \U$6774 ( \7151 , RIc226c50_21);
and \U$6775 ( \7152 , \7151 , \932 );
nor \U$6776 ( \7153 , \7150 , \7152 );
and \U$6777 ( \7154 , \7153 , \2392 );
and \U$6778 ( \7155 , \2367 , RIc226c50_21);
nor \U$6779 ( \7156 , \7154 , \7155 );
not \U$6780 ( \7157 , \1340 );
and \U$6781 ( \7158 , \1770 , RIc2271f0_9);
not \U$6782 ( \7159 , \1770 );
and \U$6783 ( \7160 , \7159 , \1342 );
nor \U$6784 ( \7161 , \7158 , \7160 );
not \U$6785 ( \7162 , \7161 );
or \U$6786 ( \7163 , \7157 , \7162 );
not \U$6787 ( \7164 , \7113 );
or \U$6788 ( \7165 , \7164 , \1364 );
nand \U$6789 ( \7166 , \7163 , \7165 );
xor \U$6790 ( \7167 , \7156 , \7166 );
or \U$6791 ( \7168 , \7050 , \1308 );
and \U$6792 ( \7169 , \1602 , RIc227100_11);
and \U$6793 ( \7170 , \1533 , \1302 );
nor \U$6794 ( \7171 , \7169 , \7170 );
or \U$6795 ( \7172 , \7171 , \1312 );
nand \U$6796 ( \7173 , \7168 , \7172 );
xor \U$6797 ( \7174 , \7167 , \7173 );
xor \U$6798 ( \7175 , \7149 , \7174 );
xor \U$6799 ( \7176 , \7099 , \7175 );
not \U$6800 ( \7177 , \4803 );
and \U$6801 ( \7178 , RIc2275b0_1, \7177 );
and \U$6802 ( \7179 , \1758 , \1533 );
not \U$6803 ( \7180 , \1758 );
and \U$6804 ( \7181 , \7180 , \1534 );
nor \U$6805 ( \7182 , \7179 , \7181 );
or \U$6806 ( \7183 , \7182 , \1679 );
or \U$6807 ( \7184 , \7024 , \1757 );
nand \U$6808 ( \7185 , \7183 , \7184 );
xor \U$6809 ( \7186 , \7178 , \7185 );
xnor \U$6810 ( \7187 , \2593 , RIc2275b0_1);
or \U$6811 ( \7188 , \7187 , \855 );
not \U$6812 ( \7189 , \7133 );
or \U$6813 ( \7190 , \7189 , \899 );
nand \U$6814 ( \7191 , \7188 , \7190 );
xor \U$6815 ( \7192 , \7186 , \7191 );
xor \U$6816 ( \7193 , \7040 , \7052 );
xor \U$6817 ( \7194 , \7193 , \7095 );
xor \U$6818 ( \7195 , \7192 , \7194 );
not \U$6819 ( \7196 , \7040 );
not \U$6820 ( \7197 , \1311 );
and \U$6821 ( \7198 , \7111 , RIc227100_11);
not \U$6822 ( \7199 , \7111 );
and \U$6823 ( \7200 , \7199 , \1685 );
nor \U$6824 ( \7201 , \7198 , \7200 );
not \U$6825 ( \7202 , \7201 );
or \U$6826 ( \7203 , \7197 , \7202 );
nand \U$6827 ( \7204 , \4944 , \1307 );
nand \U$6828 ( \7205 , \7203 , \7204 );
not \U$6829 ( \7206 , \1597 );
not \U$6830 ( \7207 , \4998 );
or \U$6831 ( \7208 , \7206 , \7207 );
and \U$6832 ( \7209 , \2774 , RIc2271f0_9);
and \U$6833 ( \7210 , \2306 , \1351 );
nor \U$6834 ( \7211 , \7209 , \7210 );
or \U$6835 ( \7212 , \7211 , \1552 );
nand \U$6836 ( \7213 , \7208 , \7212 );
xor \U$6837 ( \7214 , \7205 , \7213 );
not \U$6838 ( \7215 , \1945 );
not \U$6839 ( \7216 , \4988 );
or \U$6840 ( \7217 , \7215 , \7216 );
and \U$6841 ( \7218 , \1171 , RIc226e30_17);
and \U$6842 ( \7219 , \1403 , \1960 );
nor \U$6843 ( \7220 , \7218 , \7219 );
or \U$6844 ( \7221 , \7220 , \7145 );
nand \U$6845 ( \7222 , \7217 , \7221 );
and \U$6846 ( \7223 , \7214 , \7222 );
and \U$6847 ( \7224 , \7205 , \7213 );
or \U$6848 ( \7225 , \7223 , \7224 );
xor \U$6849 ( \7226 , \7196 , \7225 );
not \U$6850 ( \7227 , \2367 );
not \U$6851 ( \7228 , RIc226c50_21);
not \U$6852 ( \7229 , \2865 );
or \U$6853 ( \7230 , \7228 , \7229 );
nand \U$6854 ( \7231 , \891 , \3204 );
nand \U$6855 ( \7232 , \7230 , \7231 );
not \U$6856 ( \7233 , \7232 );
or \U$6857 ( \7234 , \7227 , \7233 );
nand \U$6858 ( \7235 , \4906 , \2392 );
nand \U$6859 ( \7236 , \7234 , \7235 );
not \U$6860 ( \7237 , \954 );
not \U$6861 ( \7238 , \7058 );
or \U$6862 ( \7239 , \7237 , \7238 );
nand \U$6863 ( \7240 , \4979 , \951 );
nand \U$6864 ( \7241 , \7239 , \7240 );
xor \U$6865 ( \7242 , \7236 , \7241 );
not \U$6866 ( \7243 , \1118 );
not \U$6867 ( \7244 , \5010 );
or \U$6868 ( \7245 , \7243 , \7244 );
nand \U$6869 ( \7246 , \7085 , \1121 );
nand \U$6870 ( \7247 , \7245 , \7246 );
and \U$6871 ( \7248 , \7242 , \7247 );
and \U$6872 ( \7249 , \7236 , \7241 );
or \U$6873 ( \7250 , \7248 , \7249 );
and \U$6874 ( \7251 , \7226 , \7250 );
and \U$6875 ( \7252 , \7196 , \7225 );
or \U$6876 ( \7253 , \7251 , \7252 );
and \U$6877 ( \7254 , \7195 , \7253 );
and \U$6878 ( \7255 , \7192 , \7194 );
or \U$6879 ( \7256 , \7254 , \7255 );
and \U$6880 ( \7257 , \7176 , \7256 );
and \U$6881 ( \7258 , \7099 , \7175 );
or \U$6882 ( \7259 , \7257 , \7258 );
xor \U$6883 ( \7260 , \7127 , \7148 );
and \U$6884 ( \7261 , \7260 , \7174 );
and \U$6885 ( \7262 , \7127 , \7148 );
or \U$6886 ( \7263 , \7261 , \7262 );
not \U$6887 ( \7264 , \7156 );
xor \U$6888 ( \7265 , \7128 , \7135 );
and \U$6889 ( \7266 , \7265 , \7147 );
and \U$6890 ( \7267 , \7128 , \7135 );
or \U$6891 ( \7268 , \7266 , \7267 );
xor \U$6892 ( \7269 , \7264 , \7268 );
xor \U$6893 ( \7270 , \6963 , \6975 );
and \U$6894 ( \7271 , \7270 , \6991 );
and \U$6895 ( \7272 , \6963 , \6975 );
or \U$6896 ( \7273 , \7271 , \7272 );
xor \U$6897 ( \7274 , \7269 , \7273 );
xor \U$6898 ( \7275 , \7263 , \7274 );
or \U$6899 ( \7276 , \1915 , \1930 );
nand \U$6900 ( \7277 , \7276 , RIc226b60_23);
not \U$6901 ( \7278 , \2392 );
and \U$6902 ( \7279 , \1073 , RIc226c50_21);
not \U$6903 ( \7280 , \1073 );
and \U$6904 ( \7281 , \7280 , \2370 );
nor \U$6905 ( \7282 , \7279 , \7281 );
not \U$6906 ( \7283 , \7282 );
or \U$6907 ( \7284 , \7278 , \7283 );
nand \U$6908 ( \7285 , \7153 , \2367 );
nand \U$6909 ( \7286 , \7284 , \7285 );
xor \U$6910 ( \7287 , \7277 , \7286 );
and \U$6911 ( \7288 , \1022 , RIc226e30_17);
and \U$6912 ( \7289 , \1127 , \1952 );
nor \U$6913 ( \7290 , \7288 , \7289 );
or \U$6914 ( \7291 , \7290 , \7140 );
or \U$6915 ( \7292 , \7139 , \7145 );
nand \U$6916 ( \7293 , \7291 , \7292 );
and \U$6917 ( \7294 , \7287 , \7293 );
and \U$6918 ( \7295 , \7277 , \7286 );
or \U$6919 ( \7296 , \7294 , \7295 );
xor \U$6920 ( \7297 , \7178 , \7185 );
and \U$6921 ( \7298 , \7297 , \7191 );
and \U$6922 ( \7299 , \7178 , \7185 );
or \U$6923 ( \7300 , \7298 , \7299 );
xor \U$6924 ( \7301 , \7296 , \7300 );
not \U$6925 ( \7302 , \1040 );
and \U$6926 ( \7303 , \1990 , \1078 );
not \U$6927 ( \7304 , \1990 );
and \U$6928 ( \7305 , \7304 , RIc2274c0_3);
nor \U$6929 ( \7306 , \7303 , \7305 );
not \U$6930 ( \7307 , \7306 );
or \U$6931 ( \7308 , \7302 , \7307 );
nand \U$6932 ( \7309 , \7004 , \1082 );
nand \U$6933 ( \7310 , \7308 , \7309 );
not \U$6934 ( \7311 , \2534 );
not \U$6935 ( \7312 , \6988 );
or \U$6936 ( \7313 , \7311 , \7312 );
and \U$6937 ( \7314 , \841 , RIc226d40_19);
not \U$6938 ( \7315 , \841 );
and \U$6939 ( \7316 , \7315 , \1941 );
nor \U$6940 ( \7317 , \7314 , \7316 );
nand \U$6941 ( \7318 , \2518 , \7317 );
nand \U$6942 ( \7319 , \7313 , \7318 );
xor \U$6943 ( \7320 , \7310 , \7319 );
not \U$6944 ( \7321 , \7064 );
or \U$6945 ( \7322 , \7321 , \952 );
or \U$6946 ( \7323 , \7018 , \955 );
nand \U$6947 ( \7324 , \7322 , \7323 );
and \U$6948 ( \7325 , \7320 , \7324 );
and \U$6949 ( \7326 , \7310 , \7319 );
or \U$6950 ( \7327 , \7325 , \7326 );
and \U$6951 ( \7328 , \7301 , \7327 );
and \U$6952 ( \7329 , \7296 , \7300 );
or \U$6953 ( \7330 , \7328 , \7329 );
xor \U$6954 ( \7331 , \7275 , \7330 );
and \U$6955 ( \7332 , RIc2275b0_1, \2480 );
not \U$6956 ( \7333 , \2534 );
not \U$6957 ( \7334 , \7317 );
or \U$6958 ( \7335 , \7333 , \7334 );
not \U$6959 ( \7336 , RIc226d40_19);
not \U$6960 ( \7337 , \1490 );
or \U$6961 ( \7338 , \7336 , \7337 );
not \U$6962 ( \7339 , \1559 );
nand \U$6963 ( \7340 , \7339 , \1941 );
nand \U$6964 ( \7341 , \7338 , \7340 );
nand \U$6965 ( \7342 , \7341 , \2518 );
nand \U$6966 ( \7343 , \7335 , \7342 );
xor \U$6967 ( \7344 , \7332 , \7343 );
not \U$6968 ( \7345 , \1307 );
not \U$6969 ( \7346 , \7201 );
or \U$6970 ( \7347 , \7345 , \7346 );
nand \U$6971 ( \7348 , \7045 , \1311 );
nand \U$6972 ( \7349 , \7347 , \7348 );
and \U$6973 ( \7350 , \7344 , \7349 );
and \U$6974 ( \7351 , \7332 , \7343 );
or \U$6975 ( \7352 , \7350 , \7351 );
not \U$6976 ( \7353 , RIc227010_13);
not \U$6977 ( \7354 , \1949 );
or \U$6978 ( \7355 , \7353 , \7354 );
nand \U$6979 ( \7356 , \1335 , \1758 );
nand \U$6980 ( \7357 , \7355 , \7356 );
not \U$6981 ( \7358 , \7357 );
or \U$6982 ( \7359 , \7358 , \1679 );
or \U$6983 ( \7360 , \7182 , \1757 );
nand \U$6984 ( \7361 , \7359 , \7360 );
xor \U$6985 ( \7362 , RIc2275b0_1, \7177 );
not \U$6986 ( \7363 , \7362 );
or \U$6987 ( \7364 , \7363 , \855 );
or \U$6988 ( \7365 , \7187 , \899 );
nand \U$6989 ( \7366 , \7364 , \7365 );
xor \U$6990 ( \7367 , \7361 , \7366 );
and \U$6991 ( \7368 , \2015 , RIc2274c0_3);
and \U$6992 ( \7369 , \2018 , \1078 );
nor \U$6993 ( \7370 , \7368 , \7369 );
or \U$6994 ( \7371 , \7370 , \1041 );
not \U$6995 ( \7372 , \7306 );
or \U$6996 ( \7373 , \7372 , \1083 );
nand \U$6997 ( \7374 , \7371 , \7373 );
and \U$6998 ( \7375 , \7367 , \7374 );
and \U$6999 ( \7376 , \7361 , \7366 );
or \U$7000 ( \7377 , \7375 , \7376 );
xor \U$7001 ( \7378 , \7352 , \7377 );
or \U$7002 ( \7379 , \7220 , \7140 );
or \U$7003 ( \7380 , \7290 , \7145 );
nand \U$7004 ( \7381 , \7379 , \7380 );
not \U$7005 ( \7382 , \2367 );
not \U$7006 ( \7383 , \7282 );
or \U$7007 ( \7384 , \7382 , \7383 );
nand \U$7008 ( \7385 , \7232 , \2392 );
nand \U$7009 ( \7386 , \7384 , \7385 );
xor \U$7010 ( \7387 , \7381 , \7386 );
not \U$7011 ( \7388 , \1340 );
not \U$7012 ( \7389 , \7105 );
or \U$7013 ( \7390 , \7388 , \7389 );
or \U$7014 ( \7391 , \7211 , \1364 );
nand \U$7015 ( \7392 , \7390 , \7391 );
and \U$7016 ( \7393 , \7387 , \7392 );
and \U$7017 ( \7394 , \7381 , \7386 );
or \U$7018 ( \7395 , \7393 , \7394 );
and \U$7019 ( \7396 , \7378 , \7395 );
and \U$7020 ( \7397 , \7352 , \7377 );
or \U$7021 ( \7398 , \7396 , \7397 );
not \U$7022 ( \7399 , \7398 );
xor \U$7023 ( \7400 , \7296 , \7300 );
xor \U$7024 ( \7401 , \7400 , \7327 );
not \U$7025 ( \7402 , \7401 );
or \U$7026 ( \7403 , \7399 , \7402 );
or \U$7027 ( \7404 , \7401 , \7398 );
xor \U$7028 ( \7405 , \7277 , \7286 );
xor \U$7029 ( \7406 , \7405 , \7293 );
xor \U$7030 ( \7407 , \7310 , \7319 );
xor \U$7031 ( \7408 , \7407 , \7324 );
xor \U$7032 ( \7409 , \7406 , \7408 );
xor \U$7033 ( \7410 , \7115 , \7120 );
xor \U$7034 ( \7411 , \7410 , \7124 );
and \U$7035 ( \7412 , \7409 , \7411 );
and \U$7036 ( \7413 , \7406 , \7408 );
or \U$7037 ( \7414 , \7412 , \7413 );
nand \U$7038 ( \7415 , \7404 , \7414 );
nand \U$7039 ( \7416 , \7403 , \7415 );
xor \U$7040 ( \7417 , \7331 , \7416 );
xor \U$7041 ( \7418 , \7007 , \7020 );
and \U$7042 ( \7419 , \7418 , \7030 );
and \U$7043 ( \7420 , \7007 , \7020 );
or \U$7044 ( \7421 , \7419 , \7420 );
xor \U$7045 ( \7422 , \7156 , \7166 );
and \U$7046 ( \7423 , \7422 , \7173 );
and \U$7047 ( \7424 , \7156 , \7166 );
or \U$7048 ( \7425 , \7423 , \7424 );
xor \U$7049 ( \7426 , \7421 , \7425 );
and \U$7050 ( \7427 , RIc2275b0_1, \2018 );
not \U$7051 ( \7428 , \1597 );
not \U$7052 ( \7429 , \7161 );
or \U$7053 ( \7430 , \7428 , \7429 );
and \U$7054 ( \7431 , \1342 , \1949 );
not \U$7055 ( \7432 , \1342 );
and \U$7056 ( \7433 , \7432 , \4778 );
nor \U$7057 ( \7434 , \7431 , \7433 );
nand \U$7058 ( \7435 , \7434 , \1340 );
nand \U$7059 ( \7436 , \7430 , \7435 );
xor \U$7060 ( \7437 , \7427 , \7436 );
or \U$7061 ( \7438 , \7171 , \1308 );
and \U$7062 ( \7439 , \1685 , \1393 );
not \U$7063 ( \7440 , \1685 );
and \U$7064 ( \7441 , \7440 , \1396 );
nor \U$7065 ( \7442 , \7439 , \7441 );
not \U$7066 ( \7443 , \7442 );
or \U$7067 ( \7444 , \7443 , \1312 );
nand \U$7068 ( \7445 , \7438 , \7444 );
xor \U$7069 ( \7446 , \7437 , \7445 );
xor \U$7070 ( \7447 , \7426 , \7446 );
xor \U$7071 ( \7448 , \6992 , \7031 );
and \U$7072 ( \7449 , \7448 , \7098 );
and \U$7073 ( \7450 , \6992 , \7031 );
or \U$7074 ( \7451 , \7449 , \7450 );
xor \U$7075 ( \7452 , \7447 , \7451 );
or \U$7076 ( \7453 , \2392 , \2367 );
nand \U$7077 ( \7454 , \7453 , RIc226c50_21);
not \U$7078 ( \7455 , \2518 );
not \U$7079 ( \7456 , \6982 );
or \U$7080 ( \7457 , \7455 , \7456 );
and \U$7081 ( \7458 , \932 , RIc226d40_19);
and \U$7082 ( \7459 , \931 , \2523 );
nor \U$7083 ( \7460 , \7458 , \7459 );
not \U$7084 ( \7461 , \2534 );
or \U$7085 ( \7462 , \7460 , \7461 );
nand \U$7086 ( \7463 , \7457 , \7462 );
xor \U$7087 ( \7464 , \7454 , \7463 );
not \U$7088 ( \7465 , \6954 );
or \U$7089 ( \7466 , \7465 , \2321 );
not \U$7090 ( \7467 , RIc226f20_15);
not \U$7091 ( \7468 , \1559 );
or \U$7092 ( \7469 , \7467 , \7468 );
nand \U$7093 ( \7470 , \7339 , \1674 );
nand \U$7094 ( \7471 , \7469 , \7470 );
not \U$7095 ( \7472 , \7471 );
or \U$7096 ( \7473 , \7472 , \3305 );
nand \U$7097 ( \7474 , \7466 , \7473 );
xor \U$7098 ( \7475 , \7464 , \7474 );
not \U$7099 ( \7476 , \1118 );
not \U$7100 ( \7477 , \6968 );
or \U$7101 ( \7478 , \7476 , \7477 );
and \U$7102 ( \7479 , \2616 , RIc2272e0_7);
and \U$7103 ( \7480 , \7111 , \1139 );
nor \U$7104 ( \7481 , \7479 , \7480 );
or \U$7105 ( \7482 , \7481 , \1431 );
nand \U$7106 ( \7483 , \7478 , \7482 );
not \U$7107 ( \7484 , \951 );
not \U$7108 ( \7485 , \7013 );
or \U$7109 ( \7486 , \7484 , \7485 );
and \U$7110 ( \7487 , \2774 , RIc2273d0_5);
and \U$7111 ( \7488 , \2306 , \946 );
nor \U$7112 ( \7489 , \7487 , \7488 );
or \U$7113 ( \7490 , \7489 , \955 );
nand \U$7114 ( \7491 , \7486 , \7490 );
xor \U$7115 ( \7492 , \7483 , \7491 );
or \U$7116 ( \7493 , \7028 , \1679 );
and \U$7117 ( \7494 , \1171 , RIc227010_13);
and \U$7118 ( \7495 , \1228 , \1758 );
nor \U$7119 ( \7496 , \7494 , \7495 );
or \U$7120 ( \7497 , \7496 , \1757 );
nand \U$7121 ( \7498 , \7493 , \7497 );
xor \U$7122 ( \7499 , \7492 , \7498 );
xor \U$7123 ( \7500 , \7475 , \7499 );
not \U$7124 ( \7501 , \1040 );
not \U$7125 ( \7502 , \6997 );
or \U$7126 ( \7503 , \7501 , \7502 );
and \U$7127 ( \7504 , \2837 , RIc2274c0_3);
not \U$7128 ( \7505 , \2837 );
and \U$7129 ( \7506 , \7505 , \1032 );
nor \U$7130 ( \7507 , \7504 , \7506 );
nand \U$7131 ( \7508 , \7507 , \1082 );
nand \U$7132 ( \7509 , \7503 , \7508 );
not \U$7133 ( \7510 , \854 );
not \U$7134 ( \7511 , \7130 );
or \U$7135 ( \7512 , \7510 , \7511 );
xor \U$7136 ( \7513 , RIc2275b0_1, \2261 );
nand \U$7137 ( \7514 , \7513 , \1579 );
nand \U$7138 ( \7515 , \7512 , \7514 );
xor \U$7139 ( \7516 , \7509 , \7515 );
or \U$7140 ( \7517 , \7144 , \7140 );
and \U$7141 ( \7518 , \889 , RIc226e30_17);
not \U$7142 ( \7519 , \889 );
and \U$7143 ( \7520 , \7519 , \1960 );
nor \U$7144 ( \7521 , \7518 , \7520 );
not \U$7145 ( \7522 , \7521 );
or \U$7146 ( \7523 , \7522 , \7145 );
nand \U$7147 ( \7524 , \7517 , \7523 );
xor \U$7148 ( \7525 , \7516 , \7524 );
xor \U$7149 ( \7526 , \7500 , \7525 );
xor \U$7150 ( \7527 , \7452 , \7526 );
xor \U$7151 ( \7528 , \7417 , \7527 );
xor \U$7152 ( \7529 , \7259 , \7528 );
or \U$7153 ( \7530 , \2860 , \2173 );
nand \U$7154 ( \7531 , \7530 , RIc226a70_25);
not \U$7155 ( \7532 , \1915 );
not \U$7156 ( \7533 , \4936 );
or \U$7157 ( \7534 , \7532 , \7533 );
or \U$7158 ( \7535 , \7036 , \7038 );
nand \U$7159 ( \7536 , \7534 , \7535 );
xor \U$7160 ( \7537 , \7531 , \7536 );
not \U$7161 ( \7538 , \2518 );
not \U$7162 ( \7539 , \4924 );
or \U$7163 ( \7540 , \7538 , \7539 );
not \U$7164 ( \7541 , \7341 );
or \U$7165 ( \7542 , \7541 , \7461 );
nand \U$7166 ( \7543 , \7540 , \7542 );
and \U$7167 ( \7544 , \7537 , \7543 );
and \U$7168 ( \7545 , \7531 , \7536 );
or \U$7169 ( \7546 , \7544 , \7545 );
xor \U$7170 ( \7547 , \7332 , \7343 );
xor \U$7171 ( \7548 , \7547 , \7349 );
xor \U$7172 ( \7549 , \7546 , \7548 );
not \U$7173 ( \7550 , \2358 );
not \U$7174 ( \7551 , \7071 );
or \U$7175 ( \7552 , \7550 , \7551 );
nand \U$7176 ( \7553 , \4959 , \2320 );
nand \U$7177 ( \7554 , \7552 , \7553 );
not \U$7178 ( \7555 , \854 );
not \U$7179 ( \7556 , \4915 );
or \U$7180 ( \7557 , \7555 , \7556 );
nand \U$7181 ( \7558 , \7362 , \1579 );
nand \U$7182 ( \7559 , \7557 , \7558 );
xor \U$7183 ( \7560 , \7554 , \7559 );
not \U$7184 ( \7561 , \1040 );
not \U$7185 ( \7562 , \4966 );
or \U$7186 ( \7563 , \7561 , \7562 );
or \U$7187 ( \7564 , \7370 , \1083 );
nand \U$7188 ( \7565 , \7563 , \7564 );
and \U$7189 ( \7566 , \7560 , \7565 );
and \U$7190 ( \7567 , \7554 , \7559 );
or \U$7191 ( \7568 , \7566 , \7567 );
and \U$7192 ( \7569 , \7549 , \7568 );
and \U$7193 ( \7570 , \7546 , \7548 );
or \U$7194 ( \7571 , \7569 , \7570 );
xor \U$7195 ( \7572 , \7352 , \7377 );
xor \U$7196 ( \7573 , \7572 , \7395 );
xor \U$7197 ( \7574 , \7571 , \7573 );
xor \U$7198 ( \7575 , \7381 , \7386 );
xor \U$7199 ( \7576 , \7575 , \7392 );
xor \U$7200 ( \7577 , \7361 , \7366 );
xor \U$7201 ( \7578 , \7577 , \7374 );
xor \U$7202 ( \7579 , \7576 , \7578 );
xor \U$7203 ( \7580 , \7066 , \7080 );
xor \U$7204 ( \7581 , \7580 , \7092 );
and \U$7205 ( \7582 , \7579 , \7581 );
and \U$7206 ( \7583 , \7576 , \7578 );
or \U$7207 ( \7584 , \7582 , \7583 );
and \U$7208 ( \7585 , \7574 , \7584 );
and \U$7209 ( \7586 , \7571 , \7573 );
or \U$7210 ( \7587 , \7585 , \7586 );
not \U$7211 ( \7588 , \7587 );
xor \U$7212 ( \7589 , \7398 , \7414 );
not \U$7213 ( \7590 , \7401 );
and \U$7214 ( \7591 , \7589 , \7590 );
not \U$7215 ( \7592 , \7589 );
and \U$7216 ( \7593 , \7592 , \7401 );
nor \U$7217 ( \7594 , \7591 , \7593 );
not \U$7218 ( \7595 , \7594 );
not \U$7219 ( \7596 , \7595 );
or \U$7220 ( \7597 , \7588 , \7596 );
or \U$7221 ( \7598 , \7595 , \7587 );
xor \U$7222 ( \7599 , \7406 , \7408 );
xor \U$7223 ( \7600 , \7599 , \7411 );
and \U$7224 ( \7601 , RIc2275b0_1, \3026 );
xor \U$7225 ( \7602 , \5037 , \7601 );
nand \U$7226 ( \7603 , \7357 , \1682 );
nand \U$7227 ( \7604 , \5045 , \1680 );
nand \U$7228 ( \7605 , \7603 , \7604 );
and \U$7229 ( \7606 , \7602 , \7605 );
and \U$7230 ( \7607 , \5037 , \7601 );
or \U$7231 ( \7608 , \7606 , \7607 );
not \U$7232 ( \7609 , \4938 );
not \U$7233 ( \7610 , \4928 );
or \U$7234 ( \7611 , \7609 , \7610 );
or \U$7235 ( \7612 , \4928 , \4938 );
nand \U$7236 ( \7613 , \7612 , \4948 );
nand \U$7237 ( \7614 , \7611 , \7613 );
xor \U$7238 ( \7615 , \4992 , \5002 );
and \U$7239 ( \7616 , \7615 , \5012 );
and \U$7240 ( \7617 , \4992 , \5002 );
or \U$7241 ( \7618 , \7616 , \7617 );
xor \U$7242 ( \7619 , \7614 , \7618 );
xor \U$7243 ( \7620 , \4961 , \4970 );
and \U$7244 ( \7621 , \7620 , \4981 );
and \U$7245 ( \7622 , \4961 , \4970 );
or \U$7246 ( \7623 , \7621 , \7622 );
and \U$7247 ( \7624 , \7619 , \7623 );
and \U$7248 ( \7625 , \7614 , \7618 );
or \U$7249 ( \7626 , \7624 , \7625 );
xor \U$7250 ( \7627 , \7608 , \7626 );
xor \U$7251 ( \7628 , \7196 , \7225 );
xor \U$7252 ( \7629 , \7628 , \7250 );
and \U$7253 ( \7630 , \7627 , \7629 );
and \U$7254 ( \7631 , \7608 , \7626 );
or \U$7255 ( \7632 , \7630 , \7631 );
xor \U$7256 ( \7633 , \7600 , \7632 );
xor \U$7257 ( \7634 , \7546 , \7548 );
xor \U$7258 ( \7635 , \7634 , \7568 );
xor \U$7259 ( \7636 , \7531 , \7536 );
xor \U$7260 ( \7637 , \7636 , \7543 );
xor \U$7261 ( \7638 , \7236 , \7241 );
xor \U$7262 ( \7639 , \7638 , \7247 );
xor \U$7263 ( \7640 , \7637 , \7639 );
xor \U$7264 ( \7641 , \7554 , \7559 );
xor \U$7265 ( \7642 , \7641 , \7565 );
and \U$7266 ( \7643 , \7640 , \7642 );
and \U$7267 ( \7644 , \7637 , \7639 );
or \U$7268 ( \7645 , \7643 , \7644 );
xor \U$7269 ( \7646 , \7635 , \7645 );
xor \U$7270 ( \7647 , \5037 , \7601 );
xor \U$7271 ( \7648 , \7647 , \7605 );
xor \U$7272 ( \7649 , \4900 , \4910 );
and \U$7273 ( \7650 , \7649 , \4917 );
and \U$7274 ( \7651 , \4900 , \4910 );
or \U$7275 ( \7652 , \7650 , \7651 );
xor \U$7276 ( \7653 , \7648 , \7652 );
xor \U$7277 ( \7654 , \7205 , \7213 );
xor \U$7278 ( \7655 , \7654 , \7222 );
and \U$7279 ( \7656 , \7653 , \7655 );
and \U$7280 ( \7657 , \7648 , \7652 );
or \U$7281 ( \7658 , \7656 , \7657 );
and \U$7282 ( \7659 , \7646 , \7658 );
and \U$7283 ( \7660 , \7635 , \7645 );
or \U$7284 ( \7661 , \7659 , \7660 );
and \U$7285 ( \7662 , \7633 , \7661 );
and \U$7286 ( \7663 , \7600 , \7632 );
or \U$7287 ( \7664 , \7662 , \7663 );
nand \U$7288 ( \7665 , \7598 , \7664 );
nand \U$7289 ( \7666 , \7597 , \7665 );
xor \U$7290 ( \7667 , \7529 , \7666 );
not \U$7291 ( \7668 , \7667 );
xor \U$7292 ( \7669 , \7099 , \7175 );
xor \U$7293 ( \7670 , \7669 , \7256 );
not \U$7294 ( \7671 , \7670 );
xor \U$7295 ( \7672 , \7594 , \7587 );
xor \U$7296 ( \7673 , \7672 , \7664 );
xor \U$7297 ( \7674 , \7671 , \7673 );
xor \U$7298 ( \7675 , \7192 , \7194 );
xor \U$7299 ( \7676 , \7675 , \7253 );
not \U$7300 ( \7677 , \7676 );
xor \U$7301 ( \7678 , \7571 , \7573 );
xor \U$7302 ( \7679 , \7678 , \7584 );
not \U$7303 ( \7680 , \7679 );
or \U$7304 ( \7681 , \7677 , \7680 );
or \U$7305 ( \7682 , \7679 , \7676 );
xor \U$7306 ( \7683 , \7576 , \7578 );
xor \U$7307 ( \7684 , \7683 , \7581 );
not \U$7308 ( \7685 , \7684 );
xor \U$7309 ( \7686 , \7608 , \7626 );
xor \U$7310 ( \7687 , \7686 , \7629 );
not \U$7311 ( \7688 , \7687 );
or \U$7312 ( \7689 , \7685 , \7688 );
or \U$7313 ( \7690 , \7687 , \7684 );
xor \U$7314 ( \7691 , \5038 , \5048 );
and \U$7315 ( \7692 , \7691 , \5053 );
and \U$7316 ( \7693 , \5038 , \5048 );
or \U$7317 ( \7694 , \7692 , \7693 );
xor \U$7318 ( \7695 , \5060 , \5064 );
and \U$7319 ( \7696 , \7695 , \5069 );
and \U$7320 ( \7697 , \5060 , \5064 );
or \U$7321 ( \7698 , \7696 , \7697 );
xor \U$7322 ( \7699 , \7694 , \7698 );
xor \U$7323 ( \7700 , \7614 , \7618 );
xor \U$7324 ( \7701 , \7700 , \7623 );
and \U$7325 ( \7702 , \7699 , \7701 );
and \U$7326 ( \7703 , \7694 , \7698 );
or \U$7327 ( \7704 , \7702 , \7703 );
nand \U$7328 ( \7705 , \7690 , \7704 );
nand \U$7329 ( \7706 , \7689 , \7705 );
nand \U$7330 ( \7707 , \7682 , \7706 );
nand \U$7331 ( \7708 , \7681 , \7707 );
not \U$7332 ( \7709 , \7708 );
and \U$7333 ( \7710 , \7674 , \7709 );
and \U$7334 ( \7711 , \7671 , \7673 );
or \U$7335 ( \7712 , \7710 , \7711 );
nand \U$7336 ( \7713 , \7668 , \7712 );
xor \U$7337 ( \7714 , \7447 , \7451 );
and \U$7338 ( \7715 , \7714 , \7526 );
and \U$7339 ( \7716 , \7447 , \7451 );
or \U$7340 ( \7717 , \7715 , \7716 );
xor \U$7341 ( \7718 , \7331 , \7416 );
and \U$7342 ( \7719 , \7718 , \7527 );
and \U$7343 ( \7720 , \7331 , \7416 );
or \U$7344 ( \7721 , \7719 , \7720 );
xor \U$7345 ( \7722 , \7717 , \7721 );
xor \U$7346 ( \7723 , \7263 , \7274 );
and \U$7347 ( \7724 , \7723 , \7330 );
and \U$7348 ( \7725 , \7263 , \7274 );
or \U$7349 ( \7726 , \7724 , \7725 );
or \U$7350 ( \7727 , \7460 , \5700 );
or \U$7351 ( \7728 , \7461 , \1941 );
nand \U$7352 ( \7729 , \7727 , \7728 );
not \U$7353 ( \7730 , \7729 );
or \U$7354 ( \7731 , \7481 , \1117 );
and \U$7355 ( \7732 , \1488 , RIc2272e0_7);
and \U$7356 ( \7733 , \1770 , \1423 );
nor \U$7357 ( \7734 , \7732 , \7733 );
or \U$7358 ( \7735 , \7734 , \1431 );
nand \U$7359 ( \7736 , \7731 , \7735 );
xor \U$7360 ( \7737 , \7730 , \7736 );
xor \U$7361 ( \7738 , \7509 , \7515 );
and \U$7362 ( \7739 , \7738 , \7524 );
and \U$7363 ( \7740 , \7509 , \7515 );
or \U$7364 ( \7741 , \7739 , \7740 );
xor \U$7365 ( \7742 , \7737 , \7741 );
xor \U$7366 ( \7743 , \7264 , \7268 );
and \U$7367 ( \7744 , \7743 , \7273 );
and \U$7368 ( \7745 , \7264 , \7268 );
or \U$7369 ( \7746 , \7744 , \7745 );
xor \U$7370 ( \7747 , \7742 , \7746 );
xor \U$7371 ( \7748 , \7475 , \7499 );
and \U$7372 ( \7749 , \7748 , \7525 );
and \U$7373 ( \7750 , \7475 , \7499 );
or \U$7374 ( \7751 , \7749 , \7750 );
xor \U$7375 ( \7752 , \7747 , \7751 );
xor \U$7376 ( \7753 , \7726 , \7752 );
xor \U$7377 ( \7754 , \7421 , \7425 );
and \U$7378 ( \7755 , \7754 , \7446 );
and \U$7379 ( \7756 , \7421 , \7425 );
or \U$7380 ( \7757 , \7755 , \7756 );
xor \U$7381 ( \7758 , \7454 , \7463 );
and \U$7382 ( \7759 , \7758 , \7474 );
and \U$7383 ( \7760 , \7454 , \7463 );
or \U$7384 ( \7761 , \7759 , \7760 );
xor \U$7385 ( \7762 , \7427 , \7436 );
and \U$7386 ( \7763 , \7762 , \7445 );
and \U$7387 ( \7764 , \7427 , \7436 );
or \U$7388 ( \7765 , \7763 , \7764 );
xor \U$7389 ( \7766 , \7761 , \7765 );
xor \U$7390 ( \7767 , \7483 , \7491 );
and \U$7391 ( \7768 , \7767 , \7498 );
and \U$7392 ( \7769 , \7483 , \7491 );
or \U$7393 ( \7770 , \7768 , \7769 );
xor \U$7394 ( \7771 , \7766 , \7770 );
xor \U$7395 ( \7772 , \7757 , \7771 );
and \U$7396 ( \7773 , RIc2275b0_1, \1991 );
not \U$7397 ( \7774 , \1363 );
not \U$7398 ( \7775 , \7434 );
or \U$7399 ( \7776 , \7774 , \7775 );
not \U$7400 ( \7777 , RIc2271f0_9);
not \U$7401 ( \7778 , \1602 );
or \U$7402 ( \7779 , \7777 , \7778 );
nand \U$7403 ( \7780 , \1533 , \1342 );
nand \U$7404 ( \7781 , \7779 , \7780 );
nand \U$7405 ( \7782 , \7781 , \1340 );
nand \U$7406 ( \7783 , \7776 , \7782 );
xor \U$7407 ( \7784 , \7773 , \7783 );
and \U$7408 ( \7785 , \2301 , \1706 );
not \U$7409 ( \7786 , \2301 );
and \U$7410 ( \7787 , \7786 , \841 );
nor \U$7411 ( \7788 , \7785 , \7787 );
and \U$7412 ( \7789 , \7788 , \2358 );
and \U$7413 ( \7790 , \7471 , \2320 );
nor \U$7414 ( \7791 , \7789 , \7790 );
not \U$7415 ( \7792 , \7791 );
xor \U$7416 ( \7793 , \7784 , \7792 );
not \U$7417 ( \7794 , \1311 );
and \U$7418 ( \7795 , \3337 , RIc227100_11);
not \U$7419 ( \7796 , \3337 );
and \U$7420 ( \7797 , \7796 , \1685 );
nor \U$7421 ( \7798 , \7795 , \7797 );
not \U$7422 ( \7799 , \7798 );
or \U$7423 ( \7800 , \7794 , \7799 );
nand \U$7424 ( \7801 , \7442 , \1307 );
nand \U$7425 ( \7802 , \7800 , \7801 );
not \U$7426 ( \7803 , \1040 );
not \U$7427 ( \7804 , \7507 );
or \U$7428 ( \7805 , \7803 , \7804 );
not \U$7429 ( \7806 , RIc2274c0_3);
not \U$7430 ( \7807 , \2424 );
or \U$7431 ( \7808 , \7806 , \7807 );
nand \U$7432 ( \7809 , \2423 , \1032 );
nand \U$7433 ( \7810 , \7808 , \7809 );
nand \U$7434 ( \7811 , \7810 , \1082 );
nand \U$7435 ( \7812 , \7805 , \7811 );
xor \U$7436 ( \7813 , \7802 , \7812 );
not \U$7437 ( \7814 , \1579 );
xor \U$7438 ( \7815 , RIc2275b0_1, \2235 );
not \U$7439 ( \7816 , \7815 );
or \U$7440 ( \7817 , \7814 , \7816 );
not \U$7441 ( \7818 , \7513 );
or \U$7442 ( \7819 , \7818 , \855 );
nand \U$7443 ( \7820 , \7817 , \7819 );
xor \U$7444 ( \7821 , \7813 , \7820 );
xor \U$7445 ( \7822 , \7793 , \7821 );
not \U$7446 ( \7823 , \1963 );
and \U$7447 ( \7824 , \1073 , RIc226e30_17);
not \U$7448 ( \7825 , \1073 );
and \U$7449 ( \7826 , \7825 , \1960 );
nor \U$7450 ( \7827 , \7824 , \7826 );
not \U$7451 ( \7828 , \7827 );
or \U$7452 ( \7829 , \7823 , \7828 );
nand \U$7453 ( \7830 , \7521 , \1945 );
nand \U$7454 ( \7831 , \7829 , \7830 );
or \U$7455 ( \7832 , \7496 , \1679 );
and \U$7456 ( \7833 , \1456 , RIc227010_13);
and \U$7457 ( \7834 , \1455 , \1758 );
nor \U$7458 ( \7835 , \7833 , \7834 );
or \U$7459 ( \7836 , \7835 , \1757 );
nand \U$7460 ( \7837 , \7832 , \7836 );
xor \U$7461 ( \7838 , \7831 , \7837 );
not \U$7462 ( \7839 , \954 );
and \U$7463 ( \7840 , RIc2273d0_5, \2348 );
not \U$7464 ( \7841 , RIc2273d0_5);
and \U$7465 ( \7842 , \7841 , \2355 );
nor \U$7466 ( \7843 , \7840 , \7842 );
not \U$7467 ( \7844 , \7843 );
or \U$7468 ( \7845 , \7839 , \7844 );
or \U$7469 ( \7846 , \7489 , \952 );
nand \U$7470 ( \7847 , \7845 , \7846 );
xor \U$7471 ( \7848 , \7838 , \7847 );
xor \U$7472 ( \7849 , \7822 , \7848 );
xor \U$7473 ( \7850 , \7772 , \7849 );
xor \U$7474 ( \7851 , \7753 , \7850 );
xor \U$7475 ( \7852 , \7722 , \7851 );
xor \U$7476 ( \7853 , \7259 , \7528 );
and \U$7477 ( \7854 , \7853 , \7666 );
and \U$7478 ( \7855 , \7259 , \7528 );
or \U$7479 ( \7856 , \7854 , \7855 );
or \U$7480 ( \7857 , \7852 , \7856 );
nand \U$7481 ( \7858 , \7713 , \7857 );
xor \U$7482 ( \7859 , \7757 , \7771 );
and \U$7483 ( \7860 , \7859 , \7849 );
and \U$7484 ( \7861 , \7757 , \7771 );
or \U$7485 ( \7862 , \7860 , \7861 );
not \U$7486 ( \7863 , \7781 );
or \U$7487 ( \7864 , \7863 , \1364 );
and \U$7488 ( \7865 , \1396 , RIc2271f0_9);
not \U$7489 ( \7866 , \1396 );
and \U$7490 ( \7867 , \7866 , \1342 );
nor \U$7491 ( \7868 , \7865 , \7867 );
not \U$7492 ( \7869 , \7868 );
or \U$7493 ( \7870 , \7869 , \1552 );
nand \U$7494 ( \7871 , \7864 , \7870 );
xor \U$7495 ( \7872 , \7871 , \7729 );
or \U$7496 ( \7873 , \7734 , \1117 );
and \U$7497 ( \7874 , \940 , \4778 );
not \U$7498 ( \7875 , \940 );
and \U$7499 ( \7876 , \7875 , \1334 );
nor \U$7500 ( \7877 , \7874 , \7876 );
or \U$7501 ( \7878 , \7877 , \1431 );
nand \U$7502 ( \7879 , \7873 , \7878 );
xor \U$7503 ( \7880 , \7872 , \7879 );
xor \U$7504 ( \7881 , \7730 , \7736 );
and \U$7505 ( \7882 , \7881 , \7741 );
and \U$7506 ( \7883 , \7730 , \7736 );
or \U$7507 ( \7884 , \7882 , \7883 );
xor \U$7508 ( \7885 , \7880 , \7884 );
xor \U$7509 ( \7886 , \7761 , \7765 );
and \U$7510 ( \7887 , \7886 , \7770 );
and \U$7511 ( \7888 , \7761 , \7765 );
or \U$7512 ( \7889 , \7887 , \7888 );
xor \U$7513 ( \7890 , \7885 , \7889 );
xor \U$7514 ( \7891 , \7742 , \7746 );
and \U$7515 ( \7892 , \7891 , \7751 );
and \U$7516 ( \7893 , \7742 , \7746 );
or \U$7517 ( \7894 , \7892 , \7893 );
xor \U$7518 ( \7895 , \7890 , \7894 );
xor \U$7519 ( \7896 , \7793 , \7821 );
and \U$7520 ( \7897 , \7896 , \7848 );
and \U$7521 ( \7898 , \7793 , \7821 );
or \U$7522 ( \7899 , \7897 , \7898 );
xor \U$7523 ( \7900 , \7773 , \7783 );
and \U$7524 ( \7901 , \7900 , \7792 );
and \U$7525 ( \7902 , \7773 , \7783 );
or \U$7526 ( \7903 , \7901 , \7902 );
xor \U$7527 ( \7904 , \7802 , \7812 );
and \U$7528 ( \7905 , \7904 , \7820 );
and \U$7529 ( \7906 , \7802 , \7812 );
or \U$7530 ( \7907 , \7905 , \7906 );
xor \U$7531 ( \7908 , \7903 , \7907 );
xor \U$7532 ( \7909 , \7831 , \7837 );
and \U$7533 ( \7910 , \7909 , \7847 );
and \U$7534 ( \7911 , \7831 , \7837 );
or \U$7535 ( \7912 , \7910 , \7911 );
xor \U$7536 ( \7913 , \7908 , \7912 );
xor \U$7537 ( \7914 , \7899 , \7913 );
or \U$7538 ( \7915 , \2518 , \2534 );
nand \U$7539 ( \7916 , \7915 , RIc226d40_19);
not \U$7540 ( \7917 , \1945 );
not \U$7541 ( \7918 , \7827 );
or \U$7542 ( \7919 , \7917 , \7918 );
and \U$7543 ( \7920 , \932 , RIc226e30_17);
and \U$7544 ( \7921 , \931 , \1960 );
nor \U$7545 ( \7922 , \7920 , \7921 );
or \U$7546 ( \7923 , \7922 , \7145 );
nand \U$7547 ( \7924 , \7919 , \7923 );
xor \U$7548 ( \7925 , \7916 , \7924 );
or \U$7549 ( \7926 , \7835 , \1679 );
and \U$7550 ( \7927 , \986 , RIc227010_13);
and \U$7551 ( \7928 , \985 , \1758 );
nor \U$7552 ( \7929 , \7927 , \7928 );
or \U$7553 ( \7930 , \7929 , \1757 );
nand \U$7554 ( \7931 , \7926 , \7930 );
xor \U$7555 ( \7932 , \7925 , \7931 );
and \U$7556 ( \7933 , RIc2275b0_1, \2261 );
not \U$7557 ( \7934 , \854 );
not \U$7558 ( \7935 , \7815 );
or \U$7559 ( \7936 , \7934 , \7935 );
xor \U$7560 ( \7937 , RIc2275b0_1, \2837 );
nand \U$7561 ( \7938 , \7937 , \1579 );
nand \U$7562 ( \7939 , \7936 , \7938 );
xor \U$7563 ( \7940 , \7933 , \7939 );
not \U$7564 ( \7941 , \7788 );
or \U$7565 ( \7942 , \7941 , \2321 );
and \U$7566 ( \7943 , \2865 , RIc226f20_15);
and \U$7567 ( \7944 , \889 , \2351 );
nor \U$7568 ( \7945 , \7943 , \7944 );
or \U$7569 ( \7946 , \7945 , \3305 );
nand \U$7570 ( \7947 , \7942 , \7946 );
xor \U$7571 ( \7948 , \7940 , \7947 );
not \U$7572 ( \7949 , \1082 );
and \U$7573 ( \7950 , \2306 , RIc2274c0_3);
not \U$7574 ( \7951 , \2306 );
and \U$7575 ( \7952 , \7951 , \1032 );
nor \U$7576 ( \7953 , \7950 , \7952 );
not \U$7577 ( \7954 , \7953 );
or \U$7578 ( \7955 , \7949 , \7954 );
nand \U$7579 ( \7956 , \7810 , \1040 );
nand \U$7580 ( \7957 , \7955 , \7956 );
not \U$7581 ( \7958 , \951 );
not \U$7582 ( \7959 , \7843 );
or \U$7583 ( \7960 , \7958 , \7959 );
and \U$7584 ( \7961 , \956 , \2616 );
not \U$7585 ( \7962 , \956 );
and \U$7586 ( \7963 , \7962 , \1730 );
nor \U$7587 ( \7964 , \7961 , \7963 );
nand \U$7588 ( \7965 , \7964 , \954 );
nand \U$7589 ( \7966 , \7960 , \7965 );
xor \U$7590 ( \7967 , \7957 , \7966 );
not \U$7591 ( \7968 , \7798 );
or \U$7592 ( \7969 , \7968 , \1308 );
and \U$7593 ( \7970 , \1171 , RIc227100_11);
and \U$7594 ( \7971 , \1228 , \1291 );
nor \U$7595 ( \7972 , \7970 , \7971 );
or \U$7596 ( \7973 , \7972 , \1312 );
nand \U$7597 ( \7974 , \7969 , \7973 );
xor \U$7598 ( \7975 , \7967 , \7974 );
xor \U$7599 ( \7976 , \7948 , \7975 );
xor \U$7600 ( \7977 , \7932 , \7976 );
xor \U$7601 ( \7978 , \7914 , \7977 );
xor \U$7602 ( \7979 , \7895 , \7978 );
xor \U$7603 ( \7980 , \7862 , \7979 );
xor \U$7604 ( \7981 , \7726 , \7752 );
and \U$7605 ( \7982 , \7981 , \7850 );
and \U$7606 ( \7983 , \7726 , \7752 );
or \U$7607 ( \7984 , \7982 , \7983 );
xor \U$7608 ( \7985 , \7980 , \7984 );
xor \U$7609 ( \7986 , \7717 , \7721 );
and \U$7610 ( \7987 , \7986 , \7851 );
and \U$7611 ( \7988 , \7717 , \7721 );
or \U$7612 ( \7989 , \7987 , \7988 );
nor \U$7613 ( \7990 , \7985 , \7989 );
nor \U$7614 ( \7991 , \7858 , \7990 );
xor \U$7615 ( \7992 , \7684 , \7704 );
xnor \U$7616 ( \7993 , \7992 , \7687 );
xor \U$7617 ( \7994 , \4899 , \4918 );
and \U$7618 ( \7995 , \7994 , \4949 );
and \U$7619 ( \7996 , \4899 , \4918 );
or \U$7620 ( \7997 , \7995 , \7996 );
xor \U$7621 ( \7998 , \7637 , \7639 );
xor \U$7622 ( \7999 , \7998 , \7642 );
xor \U$7623 ( \8000 , \7997 , \7999 );
xor \U$7624 ( \8001 , \7648 , \7652 );
xor \U$7625 ( \8002 , \8001 , \7655 );
and \U$7626 ( \8003 , \8000 , \8002 );
and \U$7627 ( \8004 , \7997 , \7999 );
or \U$7628 ( \8005 , \8003 , \8004 );
not \U$7629 ( \8006 , \8005 );
xor \U$7630 ( \8007 , \7635 , \7645 );
xor \U$7631 ( \8008 , \8007 , \7658 );
and \U$7632 ( \8009 , \8006 , \8008 );
not \U$7633 ( \8010 , \8006 );
not \U$7634 ( \8011 , \8008 );
and \U$7635 ( \8012 , \8010 , \8011 );
nor \U$7636 ( \8013 , \8009 , \8012 );
not \U$7637 ( \8014 , \8013 );
not \U$7638 ( \8015 , \8014 );
xor \U$7639 ( \8016 , \4982 , \5013 );
and \U$7640 ( \8017 , \8016 , \5018 );
and \U$7641 ( \8018 , \4982 , \5013 );
or \U$7642 ( \8019 , \8017 , \8018 );
not \U$7643 ( \8020 , \8019 );
not \U$7644 ( \8021 , \8020 );
xor \U$7645 ( \8022 , \7694 , \7698 );
xor \U$7646 ( \8023 , \8022 , \7701 );
not \U$7647 ( \8024 , \8023 );
not \U$7648 ( \8025 , \8024 );
or \U$7649 ( \8026 , \8021 , \8025 );
xor \U$7650 ( \8027 , \5054 , \5070 );
and \U$7651 ( \8028 , \8027 , \5075 );
and \U$7652 ( \8029 , \5054 , \5070 );
or \U$7653 ( \8030 , \8028 , \8029 );
nand \U$7654 ( \8031 , \8026 , \8030 );
not \U$7655 ( \8032 , \8024 );
nand \U$7656 ( \8033 , \8032 , \8019 );
nand \U$7657 ( \8034 , \8031 , \8033 );
not \U$7658 ( \8035 , \8034 );
not \U$7659 ( \8036 , \8035 );
or \U$7660 ( \8037 , \8015 , \8036 );
nand \U$7661 ( \8038 , \8034 , \8013 );
nand \U$7662 ( \8039 , \8037 , \8038 );
xor \U$7663 ( \8040 , \7993 , \8039 );
xor \U$7664 ( \8041 , \7997 , \7999 );
xor \U$7665 ( \8042 , \8041 , \8002 );
not \U$7666 ( \8043 , \8042 );
not \U$7667 ( \8044 , \8019 );
not \U$7668 ( \8045 , \8024 );
or \U$7669 ( \8046 , \8044 , \8045 );
nand \U$7670 ( \8047 , \8023 , \8020 );
nand \U$7671 ( \8048 , \8046 , \8047 );
not \U$7672 ( \8049 , \8030 );
and \U$7673 ( \8050 , \8048 , \8049 );
not \U$7674 ( \8051 , \8048 );
and \U$7675 ( \8052 , \8051 , \8030 );
nor \U$7676 ( \8053 , \8050 , \8052 );
not \U$7677 ( \8054 , \8053 );
not \U$7678 ( \8055 , \8054 );
or \U$7679 ( \8056 , \8043 , \8055 );
not \U$7680 ( \8057 , \8042 );
not \U$7681 ( \8058 , \8057 );
not \U$7682 ( \8059 , \8053 );
or \U$7683 ( \8060 , \8058 , \8059 );
xor \U$7684 ( \8061 , \4895 , \4950 );
and \U$7685 ( \8062 , \8061 , \5019 );
and \U$7686 ( \8063 , \4895 , \4950 );
or \U$7687 ( \8064 , \8062 , \8063 );
nand \U$7688 ( \8065 , \8060 , \8064 );
nand \U$7689 ( \8066 , \8056 , \8065 );
xor \U$7690 ( \8067 , \8040 , \8066 );
or \U$7691 ( \8068 , \5025 , \5076 );
nand \U$7692 ( \8069 , \8068 , \5031 );
nand \U$7693 ( \8070 , \5076 , \5025 );
and \U$7694 ( \8071 , \8069 , \8070 );
and \U$7695 ( \8072 , \8064 , \8057 );
not \U$7696 ( \8073 , \8064 );
and \U$7697 ( \8074 , \8073 , \8042 );
or \U$7698 ( \8075 , \8072 , \8074 );
xor \U$7699 ( \8076 , \8075 , \8053 );
xor \U$7700 ( \8077 , \8071 , \8076 );
not \U$7701 ( \8078 , \5020 );
nand \U$7702 ( \8079 , \8078 , \4891 );
not \U$7703 ( \8080 , \8079 );
not \U$7704 ( \8081 , \5077 );
or \U$7705 ( \8082 , \8080 , \8081 );
not \U$7706 ( \8083 , \4891 );
nand \U$7707 ( \8084 , \8083 , \5020 );
nand \U$7708 ( \8085 , \8082 , \8084 );
not \U$7709 ( \8086 , \8085 );
and \U$7710 ( \8087 , \8077 , \8086 );
and \U$7711 ( \8088 , \8071 , \8076 );
or \U$7712 ( \8089 , \8087 , \8088 );
nand \U$7713 ( \8090 , \8067 , \8089 );
xor \U$7714 ( \8091 , \8071 , \8076 );
xor \U$7715 ( \8092 , \8091 , \8086 );
xor \U$7716 ( \8093 , \4727 , \4886 );
and \U$7717 ( \8094 , \8093 , \5078 );
and \U$7718 ( \8095 , \4727 , \4886 );
or \U$7719 ( \8096 , \8094 , \8095 );
nand \U$7720 ( \8097 , \8092 , \8096 );
nand \U$7721 ( \8098 , \8090 , \8097 );
not \U$7722 ( \8099 , \8039 );
nand \U$7723 ( \8100 , \8099 , \7993 );
not \U$7724 ( \8101 , \8100 );
not \U$7725 ( \8102 , \8066 );
or \U$7726 ( \8103 , \8101 , \8102 );
not \U$7727 ( \8104 , \7993 );
nand \U$7728 ( \8105 , \8104 , \8039 );
nand \U$7729 ( \8106 , \8103 , \8105 );
not \U$7730 ( \8107 , \8106 );
xor \U$7731 ( \8108 , \7600 , \7632 );
xor \U$7732 ( \8109 , \8108 , \7661 );
not \U$7733 ( \8110 , \8109 );
xor \U$7734 ( \8111 , \7679 , \7676 );
xnor \U$7735 ( \8112 , \8111 , \7706 );
xor \U$7736 ( \8113 , \8110 , \8112 );
nand \U$7737 ( \8114 , \8011 , \8006 );
and \U$7738 ( \8115 , \8034 , \8114 );
and \U$7739 ( \8116 , \8008 , \8005 );
nor \U$7740 ( \8117 , \8115 , \8116 );
xor \U$7741 ( \8118 , \8113 , \8117 );
nand \U$7742 ( \8119 , \8107 , \8118 );
xor \U$7743 ( \8120 , \7671 , \7673 );
xor \U$7744 ( \8121 , \8120 , \7709 );
xor \U$7745 ( \8122 , \8110 , \8112 );
and \U$7746 ( \8123 , \8122 , \8117 );
and \U$7747 ( \8124 , \8110 , \8112 );
or \U$7748 ( \8125 , \8123 , \8124 );
nand \U$7749 ( \8126 , \8121 , \8125 );
nand \U$7750 ( \8127 , \8119 , \8126 );
nor \U$7751 ( \8128 , \8098 , \8127 );
nand \U$7752 ( \8129 , \7991 , \8128 );
xor \U$7753 ( \8130 , \7862 , \7979 );
and \U$7754 ( \8131 , \8130 , \7984 );
and \U$7755 ( \8132 , \7862 , \7979 );
or \U$7756 ( \8133 , \8131 , \8132 );
or \U$7757 ( \8134 , \7922 , \7140 );
or \U$7758 ( \8135 , \7145 , \1960 );
nand \U$7759 ( \8136 , \8134 , \8135 );
not \U$7760 ( \8137 , \8136 );
xor \U$7761 ( \8138 , \7916 , \7924 );
and \U$7762 ( \8139 , \8138 , \7931 );
and \U$7763 ( \8140 , \7916 , \7924 );
or \U$7764 ( \8141 , \8139 , \8140 );
xor \U$7765 ( \8142 , \8137 , \8141 );
xor \U$7766 ( \8143 , \7957 , \7966 );
and \U$7767 ( \8144 , \8143 , \7974 );
and \U$7768 ( \8145 , \7957 , \7966 );
or \U$7769 ( \8146 , \8144 , \8145 );
xor \U$7770 ( \8147 , \8142 , \8146 );
xor \U$7771 ( \8148 , \7916 , \7924 );
xor \U$7772 ( \8149 , \8148 , \7931 );
and \U$7773 ( \8150 , \7948 , \8149 );
xor \U$7774 ( \8151 , \7916 , \7924 );
xor \U$7775 ( \8152 , \8151 , \7931 );
and \U$7776 ( \8153 , \7975 , \8152 );
and \U$7777 ( \8154 , \7948 , \7975 );
or \U$7778 ( \8155 , \8150 , \8153 , \8154 );
xor \U$7779 ( \8156 , \8147 , \8155 );
and \U$7780 ( \8157 , RIc2275b0_1, \2235 );
not \U$7781 ( \8158 , \1340 );
and \U$7782 ( \8159 , \3242 , RIc2271f0_9);
not \U$7783 ( \8160 , \3242 );
and \U$7784 ( \8161 , \8160 , \1351 );
nor \U$7785 ( \8162 , \8159 , \8161 );
not \U$7786 ( \8163 , \8162 );
or \U$7787 ( \8164 , \8158 , \8163 );
nand \U$7788 ( \8165 , \7868 , \1597 );
nand \U$7789 ( \8166 , \8164 , \8165 );
xor \U$7790 ( \8167 , \8157 , \8166 );
not \U$7791 ( \8168 , \2358 );
and \U$7792 ( \8169 , \1073 , RIc226f20_15);
not \U$7793 ( \8170 , \1073 );
and \U$7794 ( \8171 , \8170 , \2301 );
nor \U$7795 ( \8172 , \8169 , \8171 );
not \U$7796 ( \8173 , \8172 );
or \U$7797 ( \8174 , \8168 , \8173 );
or \U$7798 ( \8175 , \7945 , \2321 );
nand \U$7799 ( \8176 , \8174 , \8175 );
xor \U$7800 ( \8177 , \8167 , \8176 );
xor \U$7801 ( \8178 , \7933 , \7939 );
and \U$7802 ( \8179 , \8178 , \7947 );
and \U$7803 ( \8180 , \7933 , \7939 );
or \U$7804 ( \8181 , \8179 , \8180 );
not \U$7805 ( \8182 , \1040 );
not \U$7806 ( \8183 , \7953 );
or \U$7807 ( \8184 , \8182 , \8183 );
and \U$7808 ( \8185 , \2355 , RIc2274c0_3);
and \U$7809 ( \8186 , \2348 , \1032 );
nor \U$7810 ( \8187 , \8185 , \8186 );
or \U$7811 ( \8188 , \8187 , \1083 );
nand \U$7812 ( \8189 , \8184 , \8188 );
or \U$7813 ( \8190 , \7972 , \1308 );
and \U$7814 ( \8191 , \1022 , RIc227100_11);
and \U$7815 ( \8192 , \1455 , \3351 );
nor \U$7816 ( \8193 , \8191 , \8192 );
or \U$7817 ( \8194 , \8193 , \1312 );
nand \U$7818 ( \8195 , \8190 , \8194 );
xor \U$7819 ( \8196 , \8189 , \8195 );
not \U$7820 ( \8197 , \7937 );
or \U$7821 ( \8198 , \8197 , \855 );
and \U$7822 ( \8199 , RIc2275b0_1, \3348 );
not \U$7823 ( \8200 , RIc2275b0_1);
and \U$7824 ( \8201 , \8200 , \7009 );
nor \U$7825 ( \8202 , \8199 , \8201 );
or \U$7826 ( \8203 , \8202 , \899 );
nand \U$7827 ( \8204 , \8198 , \8203 );
xor \U$7828 ( \8205 , \8196 , \8204 );
xor \U$7829 ( \8206 , \8181 , \8205 );
xor \U$7830 ( \8207 , \8177 , \8206 );
xor \U$7831 ( \8208 , \8156 , \8207 );
xor \U$7832 ( \8209 , \7871 , \7729 );
and \U$7833 ( \8210 , \8209 , \7879 );
and \U$7834 ( \8211 , \7871 , \7729 );
or \U$7835 ( \8212 , \8210 , \8211 );
or \U$7836 ( \8213 , \7877 , \1117 );
and \U$7837 ( \8214 , \1534 , RIc2272e0_7);
and \U$7838 ( \8215 , \1533 , \1423 );
nor \U$7839 ( \8216 , \8214 , \8215 );
or \U$7840 ( \8217 , \8216 , \1431 );
nand \U$7841 ( \8218 , \8213 , \8217 );
not \U$7842 ( \8219 , \7964 );
or \U$7843 ( \8220 , \8219 , \952 );
and \U$7844 ( \8221 , \1488 , RIc2273d0_5);
and \U$7845 ( \8222 , \1770 , \946 );
nor \U$7846 ( \8223 , \8221 , \8222 );
or \U$7847 ( \8224 , \8223 , \955 );
nand \U$7848 ( \8225 , \8220 , \8224 );
xor \U$7849 ( \8226 , \8218 , \8225 );
or \U$7850 ( \8227 , \7929 , \1679 );
and \U$7851 ( \8228 , RIc227010_13, \1706 );
not \U$7852 ( \8229 , RIc227010_13);
and \U$7853 ( \8230 , \8229 , \841 );
nor \U$7854 ( \8231 , \8228 , \8230 );
or \U$7855 ( \8232 , \8231 , \1757 );
nand \U$7856 ( \8233 , \8227 , \8232 );
xor \U$7857 ( \8234 , \8226 , \8233 );
xor \U$7858 ( \8235 , \8212 , \8234 );
xor \U$7859 ( \8236 , \7903 , \7907 );
and \U$7860 ( \8237 , \8236 , \7912 );
and \U$7861 ( \8238 , \7903 , \7907 );
or \U$7862 ( \8239 , \8237 , \8238 );
xor \U$7863 ( \8240 , \8235 , \8239 );
xor \U$7864 ( \8241 , \7880 , \7884 );
and \U$7865 ( \8242 , \8241 , \7889 );
and \U$7866 ( \8243 , \7880 , \7884 );
or \U$7867 ( \8244 , \8242 , \8243 );
xor \U$7868 ( \8245 , \8240 , \8244 );
xor \U$7869 ( \8246 , \7899 , \7913 );
and \U$7870 ( \8247 , \8246 , \7977 );
and \U$7871 ( \8248 , \7899 , \7913 );
or \U$7872 ( \8249 , \8247 , \8248 );
xor \U$7873 ( \8250 , \8245 , \8249 );
xor \U$7874 ( \8251 , \8208 , \8250 );
xor \U$7875 ( \8252 , \7890 , \7894 );
and \U$7876 ( \8253 , \8252 , \7978 );
and \U$7877 ( \8254 , \7890 , \7894 );
or \U$7878 ( \8255 , \8253 , \8254 );
xor \U$7879 ( \8256 , \8251 , \8255 );
nor \U$7880 ( \8257 , \8133 , \8256 );
nor \U$7881 ( \8258 , \8129 , \8257 );
nand \U$7882 ( \8259 , \6949 , \8258 );
xor \U$7883 ( \8260 , \8137 , \8141 );
and \U$7884 ( \8261 , \8260 , \8146 );
and \U$7885 ( \8262 , \8137 , \8141 );
or \U$7886 ( \8263 , \8261 , \8262 );
xor \U$7887 ( \8264 , \8157 , \8166 );
xor \U$7888 ( \8265 , \8264 , \8176 );
and \U$7889 ( \8266 , \8181 , \8265 );
xor \U$7890 ( \8267 , \8157 , \8166 );
xor \U$7891 ( \8268 , \8267 , \8176 );
and \U$7892 ( \8269 , \8205 , \8268 );
and \U$7893 ( \8270 , \8181 , \8205 );
or \U$7894 ( \8271 , \8266 , \8269 , \8270 );
xor \U$7895 ( \8272 , \8263 , \8271 );
xor \U$7896 ( \8273 , \8157 , \8166 );
and \U$7897 ( \8274 , \8273 , \8176 );
and \U$7898 ( \8275 , \8157 , \8166 );
or \U$7899 ( \8276 , \8274 , \8275 );
xor \U$7900 ( \8277 , \8218 , \8225 );
and \U$7901 ( \8278 , \8277 , \8233 );
and \U$7902 ( \8279 , \8218 , \8225 );
or \U$7903 ( \8280 , \8278 , \8279 );
xor \U$7904 ( \8281 , \8276 , \8280 );
and \U$7905 ( \8282 , RIc2275b0_1, \2837 );
or \U$7906 ( \8283 , \8231 , \1679 );
and \U$7907 ( \8284 , \1349 , RIc227010_13);
and \U$7908 ( \8285 , \889 , \1758 );
nor \U$7909 ( \8286 , \8284 , \8285 );
or \U$7910 ( \8287 , \8286 , \1757 );
nand \U$7911 ( \8288 , \8283 , \8287 );
xor \U$7912 ( \8289 , \8282 , \8288 );
or \U$7913 ( \8290 , \8216 , \1117 );
and \U$7914 ( \8291 , \1396 , \1139 );
not \U$7915 ( \8292 , \1396 );
and \U$7916 ( \8293 , \8292 , RIc2272e0_7);
nor \U$7917 ( \8294 , \8291 , \8293 );
or \U$7918 ( \8295 , \8294 , \1431 );
nand \U$7919 ( \8296 , \8290 , \8295 );
xor \U$7920 ( \8297 , \8289 , \8296 );
xor \U$7921 ( \8298 , \8281 , \8297 );
xor \U$7922 ( \8299 , \8272 , \8298 );
xor \U$7923 ( \8300 , \8212 , \8234 );
and \U$7924 ( \8301 , \8300 , \8239 );
and \U$7925 ( \8302 , \8212 , \8234 );
or \U$7926 ( \8303 , \8301 , \8302 );
or \U$7927 ( \8304 , \1945 , \1963 );
nand \U$7928 ( \8305 , \8304 , RIc226e30_17);
not \U$7929 ( \8306 , \2320 );
not \U$7930 ( \8307 , \8172 );
or \U$7931 ( \8308 , \8306 , \8307 );
and \U$7932 ( \8309 , RIc226f20_15, \932 );
not \U$7933 ( \8310 , RIc226f20_15);
and \U$7934 ( \8311 , \8310 , \931 );
nor \U$7935 ( \8312 , \8309 , \8311 );
or \U$7936 ( \8313 , \8312 , \3305 );
nand \U$7937 ( \8314 , \8308 , \8313 );
xor \U$7938 ( \8315 , \8305 , \8314 );
or \U$7939 ( \8316 , \8193 , \1308 );
and \U$7940 ( \8317 , \1559 , RIc227100_11);
and \U$7941 ( \8318 , \7339 , \1291 );
nor \U$7942 ( \8319 , \8317 , \8318 );
or \U$7943 ( \8320 , \8319 , \1312 );
nand \U$7944 ( \8321 , \8316 , \8320 );
xor \U$7945 ( \8322 , \8315 , \8321 );
not \U$7946 ( \8323 , \1597 );
not \U$7947 ( \8324 , \8162 );
or \U$7948 ( \8325 , \8323 , \8324 );
and \U$7949 ( \8326 , \1351 , \1404 );
not \U$7950 ( \8327 , \1351 );
and \U$7951 ( \8328 , \8327 , \1228 );
nor \U$7952 ( \8329 , \8326 , \8328 );
not \U$7953 ( \8330 , \8329 );
or \U$7954 ( \8331 , \8330 , \1552 );
nand \U$7955 ( \8332 , \8325 , \8331 );
or \U$7956 ( \8333 , \8187 , \1041 );
and \U$7957 ( \8334 , \2615 , RIc2274c0_3);
and \U$7958 ( \8335 , \7111 , \1032 );
nor \U$7959 ( \8336 , \8334 , \8335 );
or \U$7960 ( \8337 , \8336 , \1083 );
nand \U$7961 ( \8338 , \8333 , \8337 );
xor \U$7962 ( \8339 , \8332 , \8338 );
not \U$7963 ( \8340 , \1579 );
xor \U$7964 ( \8341 , RIc2275b0_1, \2306 );
not \U$7965 ( \8342 , \8341 );
or \U$7966 ( \8343 , \8340 , \8342 );
or \U$7967 ( \8344 , \8202 , \855 );
nand \U$7968 ( \8345 , \8343 , \8344 );
xor \U$7969 ( \8346 , \8339 , \8345 );
xor \U$7970 ( \8347 , \8322 , \8346 );
or \U$7971 ( \8348 , \8223 , \952 );
and \U$7972 ( \8349 , \1334 , RIc2273d0_5);
and \U$7973 ( \8350 , \1335 , \946 );
nor \U$7974 ( \8351 , \8349 , \8350 );
or \U$7975 ( \8352 , \8351 , \955 );
nand \U$7976 ( \8353 , \8348 , \8352 );
xor \U$7977 ( \8354 , \8353 , \8136 );
xor \U$7978 ( \8355 , \8189 , \8195 );
and \U$7979 ( \8356 , \8355 , \8204 );
and \U$7980 ( \8357 , \8189 , \8195 );
or \U$7981 ( \8358 , \8356 , \8357 );
xor \U$7982 ( \8359 , \8354 , \8358 );
xor \U$7983 ( \8360 , \8347 , \8359 );
xor \U$7984 ( \8361 , \8303 , \8360 );
xor \U$7985 ( \8362 , \8147 , \8155 );
and \U$7986 ( \8363 , \8362 , \8207 );
and \U$7987 ( \8364 , \8147 , \8155 );
or \U$7988 ( \8365 , \8363 , \8364 );
xor \U$7989 ( \8366 , \8361 , \8365 );
xor \U$7990 ( \8367 , \8299 , \8366 );
xor \U$7991 ( \8368 , \8240 , \8244 );
and \U$7992 ( \8369 , \8368 , \8249 );
and \U$7993 ( \8370 , \8240 , \8244 );
or \U$7994 ( \8371 , \8369 , \8370 );
xor \U$7995 ( \8372 , \8367 , \8371 );
xor \U$7996 ( \8373 , \8208 , \8250 );
and \U$7997 ( \8374 , \8373 , \8255 );
and \U$7998 ( \8375 , \8208 , \8250 );
or \U$7999 ( \8376 , \8374 , \8375 );
nor \U$8000 ( \8377 , \8372 , \8376 );
xor \U$8001 ( \8378 , \8353 , \8136 );
and \U$8002 ( \8379 , \8378 , \8358 );
and \U$8003 ( \8380 , \8353 , \8136 );
or \U$8004 ( \8381 , \8379 , \8380 );
xor \U$8005 ( \8382 , \8276 , \8280 );
and \U$8006 ( \8383 , \8382 , \8297 );
and \U$8007 ( \8384 , \8276 , \8280 );
or \U$8008 ( \8385 , \8383 , \8384 );
xor \U$8009 ( \8386 , \8381 , \8385 );
xor \U$8010 ( \8387 , \8282 , \8288 );
and \U$8011 ( \8388 , \8387 , \8296 );
and \U$8012 ( \8389 , \8282 , \8288 );
or \U$8013 ( \8390 , \8388 , \8389 );
xor \U$8014 ( \8391 , \8305 , \8314 );
and \U$8015 ( \8392 , \8391 , \8321 );
and \U$8016 ( \8393 , \8305 , \8314 );
or \U$8017 ( \8394 , \8392 , \8393 );
xor \U$8018 ( \8395 , \8390 , \8394 );
xor \U$8019 ( \8396 , \8332 , \8338 );
and \U$8020 ( \8397 , \8396 , \8345 );
and \U$8021 ( \8398 , \8332 , \8338 );
or \U$8022 ( \8399 , \8397 , \8398 );
xor \U$8023 ( \8400 , \8395 , \8399 );
xor \U$8024 ( \8401 , \8386 , \8400 );
xor \U$8025 ( \8402 , \8303 , \8360 );
and \U$8026 ( \8403 , \8402 , \8365 );
and \U$8027 ( \8404 , \8303 , \8360 );
or \U$8028 ( \8405 , \8403 , \8404 );
xor \U$8029 ( \8406 , \8401 , \8405 );
xor \U$8030 ( \8407 , \8322 , \8346 );
and \U$8031 ( \8408 , \8407 , \8359 );
and \U$8032 ( \8409 , \8322 , \8346 );
or \U$8033 ( \8410 , \8408 , \8409 );
not \U$8034 ( \8411 , RIc2275b0_1);
nor \U$8035 ( \8412 , \8411 , \3348 );
not \U$8036 ( \8413 , \1340 );
and \U$8037 ( \8414 , RIc2271f0_9, \1455 );
not \U$8038 ( \8415 , RIc2271f0_9);
and \U$8039 ( \8416 , \8415 , \1456 );
nor \U$8040 ( \8417 , \8414 , \8416 );
not \U$8041 ( \8418 , \8417 );
or \U$8042 ( \8419 , \8413 , \8418 );
nand \U$8043 ( \8420 , \8329 , \1597 );
nand \U$8044 ( \8421 , \8419 , \8420 );
xor \U$8045 ( \8422 , \8412 , \8421 );
not \U$8046 ( \8423 , \854 );
not \U$8047 ( \8424 , \8341 );
or \U$8048 ( \8425 , \8423 , \8424 );
not \U$8049 ( \8426 , \2348 );
and \U$8050 ( \8427 , RIc2275b0_1, \8426 );
not \U$8051 ( \8428 , RIc2275b0_1);
and \U$8052 ( \8429 , \8428 , \2348 );
nor \U$8053 ( \8430 , \8427 , \8429 );
or \U$8054 ( \8431 , \8430 , \899 );
nand \U$8055 ( \8432 , \8425 , \8431 );
xor \U$8056 ( \8433 , \8422 , \8432 );
not \U$8057 ( \8434 , \8312 );
and \U$8058 ( \8435 , \8434 , \2320 );
and \U$8059 ( \8436 , \2358 , RIc226f20_15);
nor \U$8060 ( \8437 , \8435 , \8436 );
or \U$8061 ( \8438 , \8351 , \952 );
and \U$8062 ( \8439 , \1534 , RIc2273d0_5);
and \U$8063 ( \8440 , \1533 , \946 );
nor \U$8064 ( \8441 , \8439 , \8440 );
or \U$8065 ( \8442 , \8441 , \955 );
nand \U$8066 ( \8443 , \8438 , \8442 );
xor \U$8067 ( \8444 , \8437 , \8443 );
or \U$8068 ( \8445 , \8336 , \1041 );
and \U$8069 ( \8446 , \1488 , RIc2274c0_3);
and \U$8070 ( \8447 , \1770 , \1032 );
nor \U$8071 ( \8448 , \8446 , \8447 );
or \U$8072 ( \8449 , \8448 , \1083 );
nand \U$8073 ( \8450 , \8445 , \8449 );
xor \U$8074 ( \8451 , \8444 , \8450 );
xor \U$8075 ( \8452 , \8433 , \8451 );
or \U$8076 ( \8453 , \8319 , \1308 );
and \U$8077 ( \8454 , \842 , RIc227100_11);
and \U$8078 ( \8455 , \841 , \1302 );
nor \U$8079 ( \8456 , \8454 , \8455 );
or \U$8080 ( \8457 , \8456 , \1312 );
nand \U$8081 ( \8458 , \8453 , \8457 );
or \U$8082 ( \8459 , \8286 , \1679 );
and \U$8083 ( \8460 , \1075 , RIc227010_13);
and \U$8084 ( \8461 , \1073 , \1758 );
nor \U$8085 ( \8462 , \8460 , \8461 );
or \U$8086 ( \8463 , \8462 , \1757 );
nand \U$8087 ( \8464 , \8459 , \8463 );
xor \U$8088 ( \8465 , \8458 , \8464 );
or \U$8089 ( \8466 , \8294 , \1117 );
and \U$8090 ( \8467 , \1222 , RIc2272e0_7);
and \U$8091 ( \8468 , \1223 , \940 );
nor \U$8092 ( \8469 , \8467 , \8468 );
or \U$8093 ( \8470 , \8469 , \1431 );
nand \U$8094 ( \8471 , \8466 , \8470 );
xor \U$8095 ( \8472 , \8465 , \8471 );
xor \U$8096 ( \8473 , \8452 , \8472 );
xor \U$8097 ( \8474 , \8410 , \8473 );
xor \U$8098 ( \8475 , \8263 , \8271 );
and \U$8099 ( \8476 , \8475 , \8298 );
and \U$8100 ( \8477 , \8263 , \8271 );
or \U$8101 ( \8478 , \8476 , \8477 );
xor \U$8102 ( \8479 , \8474 , \8478 );
xor \U$8103 ( \8480 , \8406 , \8479 );
xor \U$8104 ( \8481 , \8299 , \8366 );
and \U$8105 ( \8482 , \8481 , \8371 );
and \U$8106 ( \8483 , \8299 , \8366 );
or \U$8107 ( \8484 , \8482 , \8483 );
nor \U$8108 ( \8485 , \8480 , \8484 );
nor \U$8109 ( \8486 , \8377 , \8485 );
not \U$8110 ( \8487 , \8437 );
xor \U$8111 ( \8488 , \8412 , \8421 );
and \U$8112 ( \8489 , \8488 , \8432 );
and \U$8113 ( \8490 , \8412 , \8421 );
or \U$8114 ( \8491 , \8489 , \8490 );
xor \U$8115 ( \8492 , \8487 , \8491 );
xor \U$8116 ( \8493 , \8458 , \8464 );
and \U$8117 ( \8494 , \8493 , \8471 );
and \U$8118 ( \8495 , \8458 , \8464 );
or \U$8119 ( \8496 , \8494 , \8495 );
xor \U$8120 ( \8497 , \8492 , \8496 );
and \U$8121 ( \8498 , RIc2275b0_1, \2306 );
or \U$8122 ( \8499 , \8430 , \855 );
and \U$8123 ( \8500 , RIc2275b0_1, \2616 );
not \U$8124 ( \8501 , RIc2275b0_1);
and \U$8125 ( \8502 , \8501 , \1730 );
nor \U$8126 ( \8503 , \8500 , \8502 );
or \U$8127 ( \8504 , \8503 , \899 );
nand \U$8128 ( \8505 , \8499 , \8504 );
xor \U$8129 ( \8506 , \8498 , \8505 );
or \U$8130 ( \8507 , \8469 , \1117 );
and \U$8131 ( \8508 , \1171 , RIc2272e0_7);
and \U$8132 ( \8509 , \1228 , \1139 );
nor \U$8133 ( \8510 , \8508 , \8509 );
or \U$8134 ( \8511 , \8510 , \1431 );
nand \U$8135 ( \8512 , \8507 , \8511 );
xor \U$8136 ( \8513 , \8506 , \8512 );
xor \U$8137 ( \8514 , \8390 , \8394 );
and \U$8138 ( \8515 , \8514 , \8399 );
and \U$8139 ( \8516 , \8390 , \8394 );
or \U$8140 ( \8517 , \8515 , \8516 );
xor \U$8141 ( \8518 , \8513 , \8517 );
xor \U$8142 ( \8519 , \8497 , \8518 );
xor \U$8143 ( \8520 , \8433 , \8451 );
and \U$8144 ( \8521 , \8520 , \8472 );
and \U$8145 ( \8522 , \8433 , \8451 );
or \U$8146 ( \8523 , \8521 , \8522 );
xor \U$8147 ( \8524 , \8437 , \8443 );
and \U$8148 ( \8525 , \8524 , \8450 );
and \U$8149 ( \8526 , \8437 , \8443 );
or \U$8150 ( \8527 , \8525 , \8526 );
or \U$8151 ( \8528 , \2320 , \2358 );
nand \U$8152 ( \8529 , \8528 , RIc226f20_15);
not \U$8153 ( \8530 , \1597 );
not \U$8154 ( \8531 , \8417 );
or \U$8155 ( \8532 , \8530 , \8531 );
and \U$8156 ( \8533 , \1351 , \986 );
not \U$8157 ( \8534 , \1351 );
and \U$8158 ( \8535 , \8534 , \7339 );
nor \U$8159 ( \8536 , \8533 , \8535 );
nand \U$8160 ( \8537 , \8536 , \1340 );
nand \U$8161 ( \8538 , \8532 , \8537 );
xor \U$8162 ( \8539 , \8529 , \8538 );
or \U$8163 ( \8540 , \8462 , \1679 );
or \U$8164 ( \8541 , \1755 , \1757 );
nand \U$8165 ( \8542 , \8540 , \8541 );
xor \U$8166 ( \8543 , \8539 , \8542 );
xor \U$8167 ( \8544 , \8527 , \8543 );
or \U$8168 ( \8545 , \8441 , \952 );
and \U$8169 ( \8546 , RIc2273d0_5, \1393 );
not \U$8170 ( \8547 , RIc2273d0_5);
and \U$8171 ( \8548 , \8547 , \1396 );
nor \U$8172 ( \8549 , \8546 , \8548 );
or \U$8173 ( \8550 , \8549 , \955 );
nand \U$8174 ( \8551 , \8545 , \8550 );
or \U$8175 ( \8552 , \8448 , \1041 );
and \U$8176 ( \8553 , \1949 , RIc2274c0_3);
and \U$8177 ( \8554 , \4778 , \1027 );
nor \U$8178 ( \8555 , \8553 , \8554 );
or \U$8179 ( \8556 , \8555 , \1083 );
nand \U$8180 ( \8557 , \8552 , \8556 );
xor \U$8181 ( \8558 , \8551 , \8557 );
or \U$8182 ( \8559 , \8456 , \1308 );
and \U$8183 ( \8560 , \893 , RIc227100_11);
and \U$8184 ( \8561 , \892 , \1291 );
nor \U$8185 ( \8562 , \8560 , \8561 );
or \U$8186 ( \8563 , \8562 , \1312 );
nand \U$8187 ( \8564 , \8559 , \8563 );
xor \U$8188 ( \8565 , \8558 , \8564 );
xor \U$8189 ( \8566 , \8544 , \8565 );
xor \U$8190 ( \8567 , \8523 , \8566 );
xor \U$8191 ( \8568 , \8381 , \8385 );
and \U$8192 ( \8569 , \8568 , \8400 );
and \U$8193 ( \8570 , \8381 , \8385 );
or \U$8194 ( \8571 , \8569 , \8570 );
xor \U$8195 ( \8572 , \8567 , \8571 );
xor \U$8196 ( \8573 , \8519 , \8572 );
xor \U$8197 ( \8574 , \8410 , \8473 );
and \U$8198 ( \8575 , \8574 , \8478 );
and \U$8199 ( \8576 , \8410 , \8473 );
or \U$8200 ( \8577 , \8575 , \8576 );
xor \U$8201 ( \8578 , \8573 , \8577 );
xor \U$8202 ( \8579 , \8401 , \8405 );
and \U$8203 ( \8580 , \8579 , \8479 );
and \U$8204 ( \8581 , \8401 , \8405 );
or \U$8205 ( \8582 , \8580 , \8581 );
or \U$8206 ( \8583 , \8578 , \8582 );
xor \U$8207 ( \8584 , \8519 , \8572 );
and \U$8208 ( \8585 , \8584 , \8577 );
and \U$8209 ( \8586 , \8519 , \8572 );
or \U$8210 ( \8587 , \8585 , \8586 );
xor \U$8211 ( \8588 , \8487 , \8491 );
xor \U$8212 ( \8589 , \8588 , \8496 );
and \U$8213 ( \8590 , \8513 , \8589 );
xor \U$8214 ( \8591 , \8487 , \8491 );
xor \U$8215 ( \8592 , \8591 , \8496 );
and \U$8216 ( \8593 , \8517 , \8592 );
and \U$8217 ( \8594 , \8513 , \8517 );
or \U$8218 ( \8595 , \8590 , \8593 , \8594 );
xor \U$8219 ( \8596 , \8527 , \8543 );
and \U$8220 ( \8597 , \8596 , \8565 );
and \U$8221 ( \8598 , \8527 , \8543 );
or \U$8222 ( \8599 , \8597 , \8598 );
xor \U$8223 ( \8600 , \8498 , \8505 );
and \U$8224 ( \8601 , \8600 , \8512 );
and \U$8225 ( \8602 , \8498 , \8505 );
or \U$8226 ( \8603 , \8601 , \8602 );
xor \U$8227 ( \8604 , \8551 , \8557 );
and \U$8228 ( \8605 , \8604 , \8564 );
and \U$8229 ( \8606 , \8551 , \8557 );
or \U$8230 ( \8607 , \8605 , \8606 );
xor \U$8231 ( \8608 , \8603 , \8607 );
not \U$8232 ( \8609 , \1340 );
not \U$8233 ( \8610 , \1710 );
or \U$8234 ( \8611 , \8609 , \8610 );
not \U$8235 ( \8612 , \8536 );
or \U$8236 ( \8613 , \8612 , \1364 );
nand \U$8237 ( \8614 , \8611 , \8613 );
not \U$8238 ( \8615 , \954 );
not \U$8239 ( \8616 , \1737 );
or \U$8240 ( \8617 , \8615 , \8616 );
not \U$8241 ( \8618 , \8549 );
nand \U$8242 ( \8619 , \8618 , \951 );
nand \U$8243 ( \8620 , \8617 , \8619 );
xor \U$8244 ( \8621 , \8614 , \8620 );
or \U$8245 ( \8622 , \8555 , \1041 );
or \U$8246 ( \8623 , \1763 , \1083 );
nand \U$8247 ( \8624 , \8622 , \8623 );
xor \U$8248 ( \8625 , \8621 , \8624 );
xor \U$8249 ( \8626 , \8608 , \8625 );
xor \U$8250 ( \8627 , \8599 , \8626 );
not \U$8251 ( \8628 , RIc2275b0_1);
nor \U$8252 ( \8629 , \8628 , \8426 );
or \U$8253 ( \8630 , \8562 , \1308 );
or \U$8254 ( \8631 , \1689 , \1312 );
nand \U$8255 ( \8632 , \8630 , \8631 );
xor \U$8256 ( \8633 , \8629 , \8632 );
or \U$8257 ( \8634 , \8510 , \1117 );
or \U$8258 ( \8635 , \1696 , \1431 );
nand \U$8259 ( \8636 , \8634 , \8635 );
xor \U$8260 ( \8637 , \8633 , \8636 );
or \U$8261 ( \8638 , \8503 , \855 );
or \U$8262 ( \8639 , \1772 , \899 );
nand \U$8263 ( \8640 , \8638 , \8639 );
not \U$8264 ( \8641 , \1760 );
xor \U$8265 ( \8642 , \8640 , \8641 );
xor \U$8266 ( \8643 , \8529 , \8538 );
and \U$8267 ( \8644 , \8643 , \8542 );
and \U$8268 ( \8645 , \8529 , \8538 );
or \U$8269 ( \8646 , \8644 , \8645 );
xor \U$8270 ( \8647 , \8642 , \8646 );
xor \U$8271 ( \8648 , \8637 , \8647 );
xor \U$8272 ( \8649 , \8487 , \8491 );
and \U$8273 ( \8650 , \8649 , \8496 );
and \U$8274 ( \8651 , \8487 , \8491 );
or \U$8275 ( \8652 , \8650 , \8651 );
xor \U$8276 ( \8653 , \8648 , \8652 );
xor \U$8277 ( \8654 , \8627 , \8653 );
xor \U$8278 ( \8655 , \8595 , \8654 );
xor \U$8279 ( \8656 , \8523 , \8566 );
and \U$8280 ( \8657 , \8656 , \8571 );
and \U$8281 ( \8658 , \8523 , \8566 );
or \U$8282 ( \8659 , \8657 , \8658 );
xor \U$8283 ( \8660 , \8655 , \8659 );
or \U$8284 ( \8661 , \8587 , \8660 );
and \U$8285 ( \8662 , \8486 , \8583 , \8661 );
xor \U$8286 ( \8663 , \1714 , \1731 );
xor \U$8287 ( \8664 , \8663 , \1741 );
xor \U$8288 ( \8665 , \1760 , \1766 );
xor \U$8289 ( \8666 , \8665 , \1775 );
xor \U$8290 ( \8667 , \8640 , \8641 );
and \U$8291 ( \8668 , \8667 , \8646 );
and \U$8292 ( \8669 , \8640 , \8641 );
or \U$8293 ( \8670 , \8668 , \8669 );
xor \U$8294 ( \8671 , \8666 , \8670 );
xor \U$8295 ( \8672 , \8664 , \8671 );
xor \U$8296 ( \8673 , \8603 , \8607 );
and \U$8297 ( \8674 , \8673 , \8625 );
and \U$8298 ( \8675 , \8603 , \8607 );
or \U$8299 ( \8676 , \8674 , \8675 );
xor \U$8300 ( \8677 , \8629 , \8632 );
and \U$8301 ( \8678 , \8677 , \8636 );
and \U$8302 ( \8679 , \8629 , \8632 );
or \U$8303 ( \8680 , \8678 , \8679 );
xor \U$8304 ( \8681 , \8614 , \8620 );
and \U$8305 ( \8682 , \8681 , \8624 );
and \U$8306 ( \8683 , \8614 , \8620 );
or \U$8307 ( \8684 , \8682 , \8683 );
xor \U$8308 ( \8685 , \8680 , \8684 );
xor \U$8309 ( \8686 , \1684 , \1692 );
xor \U$8310 ( \8687 , \8686 , \1699 );
xor \U$8311 ( \8688 , \8685 , \8687 );
xor \U$8312 ( \8689 , \8676 , \8688 );
xor \U$8313 ( \8690 , \8637 , \8647 );
and \U$8314 ( \8691 , \8690 , \8652 );
and \U$8315 ( \8692 , \8637 , \8647 );
or \U$8316 ( \8693 , \8691 , \8692 );
xor \U$8317 ( \8694 , \8689 , \8693 );
xor \U$8318 ( \8695 , \8672 , \8694 );
xor \U$8319 ( \8696 , \8599 , \8626 );
and \U$8320 ( \8697 , \8696 , \8653 );
and \U$8321 ( \8698 , \8599 , \8626 );
or \U$8322 ( \8699 , \8697 , \8698 );
xor \U$8323 ( \8700 , \8695 , \8699 );
xor \U$8324 ( \8701 , \8595 , \8654 );
and \U$8325 ( \8702 , \8701 , \8659 );
and \U$8326 ( \8703 , \8595 , \8654 );
or \U$8327 ( \8704 , \8702 , \8703 );
nor \U$8328 ( \8705 , \8700 , \8704 );
xor \U$8329 ( \8706 , \1714 , \1731 );
xor \U$8330 ( \8707 , \8706 , \1741 );
and \U$8331 ( \8708 , \8666 , \8707 );
xor \U$8332 ( \8709 , \1714 , \1731 );
xor \U$8333 ( \8710 , \8709 , \1741 );
and \U$8334 ( \8711 , \8670 , \8710 );
and \U$8335 ( \8712 , \8666 , \8670 );
or \U$8336 ( \8713 , \8708 , \8711 , \8712 );
xor \U$8337 ( \8714 , \1702 , \1703 );
xor \U$8338 ( \8715 , \8714 , \1744 );
xor \U$8339 ( \8716 , \8680 , \8684 );
and \U$8340 ( \8717 , \8716 , \8687 );
and \U$8341 ( \8718 , \8680 , \8684 );
or \U$8342 ( \8719 , \8717 , \8718 );
xor \U$8343 ( \8720 , \8715 , \8719 );
xor \U$8344 ( \8721 , \1752 , \1778 );
xor \U$8345 ( \8722 , \8721 , \1781 );
xor \U$8346 ( \8723 , \8720 , \8722 );
xor \U$8347 ( \8724 , \8713 , \8723 );
xor \U$8348 ( \8725 , \8676 , \8688 );
and \U$8349 ( \8726 , \8725 , \8693 );
and \U$8350 ( \8727 , \8676 , \8688 );
or \U$8351 ( \8728 , \8726 , \8727 );
xor \U$8352 ( \8729 , \8724 , \8728 );
xor \U$8353 ( \8730 , \8672 , \8694 );
and \U$8354 ( \8731 , \8730 , \8699 );
and \U$8355 ( \8732 , \8672 , \8694 );
or \U$8356 ( \8733 , \8731 , \8732 );
nor \U$8357 ( \8734 , \8729 , \8733 );
nor \U$8358 ( \8735 , \8705 , \8734 );
xor \U$8359 ( \8736 , \1747 , \1749 );
xor \U$8360 ( \8737 , \8736 , \1784 );
xor \U$8361 ( \8738 , \1543 , \1566 );
xor \U$8362 ( \8739 , \8738 , \1585 );
xor \U$8363 ( \8740 , \8715 , \8719 );
and \U$8364 ( \8741 , \8740 , \8722 );
and \U$8365 ( \8742 , \8715 , \8719 );
or \U$8366 ( \8743 , \8741 , \8742 );
xor \U$8367 ( \8744 , \8739 , \8743 );
xor \U$8368 ( \8745 , \8737 , \8744 );
xor \U$8369 ( \8746 , \8713 , \8723 );
and \U$8370 ( \8747 , \8746 , \8728 );
and \U$8371 ( \8748 , \8713 , \8723 );
or \U$8372 ( \8749 , \8747 , \8748 );
or \U$8373 ( \8750 , \8745 , \8749 );
xor \U$8374 ( \8751 , \1747 , \1749 );
xor \U$8375 ( \8752 , \8751 , \1784 );
and \U$8376 ( \8753 , \8739 , \8752 );
xor \U$8377 ( \8754 , \1747 , \1749 );
xor \U$8378 ( \8755 , \8754 , \1784 );
and \U$8379 ( \8756 , \8743 , \8755 );
and \U$8380 ( \8757 , \8739 , \8743 );
or \U$8381 ( \8758 , \8753 , \8756 , \8757 );
xor \U$8382 ( \8759 , \1419 , \1462 );
xor \U$8383 ( \8760 , \8759 , \1588 );
xor \U$8384 ( \8761 , \1666 , \1787 );
xor \U$8385 ( \8762 , \8760 , \8761 );
or \U$8386 ( \8763 , \8758 , \8762 );
nand \U$8387 ( \8764 , \8662 , \8735 , \8750 , \8763 );
nor \U$8388 ( \8765 , \8259 , \8764 );
not \U$8389 ( \8766 , \8765 );
not \U$8390 ( \8767 , RIc225c60_55);
and \U$8391 ( \8768 , \8767 , RIc225cd8_54);
not \U$8392 ( \8769 , RIc225cd8_54);
and \U$8393 ( \8770 , \8769 , RIc225c60_55);
nor \U$8394 ( \8771 , \8768 , \8770 );
not \U$8395 ( \8772 , RIc225d50_53);
and \U$8396 ( \8773 , \8772 , \8769 );
and \U$8397 ( \8774 , RIc225d50_53, RIc225cd8_54);
nor \U$8398 ( \8775 , \8773 , \8774 );
nand \U$8399 ( \8776 , \8771 , \8775 );
not \U$8400 ( \8777 , \8776 );
not \U$8401 ( \8778 , \8777 );
not \U$8402 ( \8779 , RIc225d50_53);
not \U$8403 ( \8780 , \2700 );
or \U$8404 ( \8781 , \8779 , \8780 );
not \U$8405 ( \8782 , RIc225d50_53);
nand \U$8406 ( \8783 , \930 , \8782 );
nand \U$8407 ( \8784 , \8781 , \8783 );
not \U$8408 ( \8785 , \8784 );
or \U$8409 ( \8786 , \8778 , \8785 );
buf \U$8410 ( \8787 , \8771 );
not \U$8411 ( \8788 , \8787 );
nand \U$8412 ( \8789 , \8788 , RIc225d50_53);
nand \U$8413 ( \8790 , \8786 , \8789 );
not \U$8414 ( \8791 , \1363 );
not \U$8415 ( \8792 , RIc2271f0_9);
not \U$8416 ( \8793 , \618 );
not \U$8417 ( \8794 , \8793 );
not \U$8418 ( \8795 , \4084 );
or \U$8419 ( \8796 , \8794 , \8795 );
buf \U$8420 ( \8797 , \4099 );
not \U$8421 ( \8798 , \8797 );
nand \U$8422 ( \8799 , \8796 , \8798 );
nor \U$8423 ( \8800 , \540 , \670 );
and \U$8424 ( \8801 , \8799 , \8800 );
not \U$8425 ( \8802 , \8799 );
not \U$8426 ( \8803 , \8800 );
and \U$8427 ( \8804 , \8802 , \8803 );
nor \U$8428 ( \8805 , \8801 , \8804 );
buf \U$8429 ( \8806 , \8805 );
not \U$8430 ( \8807 , \8806 );
not \U$8431 ( \8808 , \8807 );
or \U$8432 ( \8809 , \8792 , \8808 );
not \U$8433 ( \8810 , \8806 );
not \U$8434 ( \8811 , \8810 );
nand \U$8435 ( \8812 , \8811 , \1342 );
nand \U$8436 ( \8813 , \8809 , \8812 );
not \U$8437 ( \8814 , \8813 );
or \U$8438 ( \8815 , \8791 , \8814 );
nor \U$8439 ( \8816 , \618 , \540 );
not \U$8440 ( \8817 , \8816 );
not \U$8441 ( \8818 , \4084 );
or \U$8442 ( \8819 , \8817 , \8818 );
and \U$8443 ( \8820 , \8797 , \541 );
nor \U$8444 ( \8821 , \8820 , \670 );
nand \U$8445 ( \8822 , \8819 , \8821 );
nand \U$8446 ( \8823 , \547 , \674 );
not \U$8447 ( \8824 , \8823 );
and \U$8448 ( \8825 , \8822 , \8824 );
not \U$8449 ( \8826 , \8822 );
and \U$8450 ( \8827 , \8826 , \8823 );
nor \U$8451 ( \8828 , \8825 , \8827 );
buf \U$8452 ( \8829 , \8828 );
not \U$8453 ( \8830 , \8829 );
not \U$8454 ( \8831 , \8830 );
and \U$8455 ( \8832 , \8831 , \1351 );
not \U$8456 ( \8833 , \8831 );
and \U$8457 ( \8834 , \8833 , RIc2271f0_9);
or \U$8458 ( \8835 , \8832 , \8834 );
nand \U$8459 ( \8836 , \8835 , \1340 );
nand \U$8460 ( \8837 , \8815 , \8836 );
xor \U$8461 ( \8838 , \8790 , \8837 );
not \U$8462 ( \8839 , \1307 );
not \U$8463 ( \8840 , RIc227100_11);
not \U$8464 ( \8841 , \630 );
nor \U$8465 ( \8842 , \618 , \8841 );
not \U$8466 ( \8843 , \8842 );
not \U$8467 ( \8844 , \4084 );
or \U$8468 ( \8845 , \8843 , \8844 );
not \U$8469 ( \8846 , \4099 );
nor \U$8470 ( \8847 , \8846 , \8841 );
nor \U$8471 ( \8848 , \8847 , \675 );
nand \U$8472 ( \8849 , \8845 , \8848 );
nand \U$8473 ( \8850 , \545 , \679 );
not \U$8474 ( \8851 , \8850 );
and \U$8475 ( \8852 , \8849 , \8851 );
not \U$8476 ( \8853 , \8849 );
and \U$8477 ( \8854 , \8853 , \8850 );
nor \U$8478 ( \8855 , \8852 , \8854 );
buf \U$8479 ( \8856 , \8855 );
not \U$8480 ( \8857 , \8856 );
not \U$8481 ( \8858 , \8857 );
or \U$8482 ( \8859 , \8840 , \8858 );
nand \U$8483 ( \8860 , \8856 , \3351 );
nand \U$8484 ( \8861 , \8859 , \8860 );
not \U$8485 ( \8862 , \8861 );
or \U$8486 ( \8863 , \8839 , \8862 );
not \U$8487 ( \8864 , RIc227100_11);
not \U$8488 ( \8865 , \8841 );
nand \U$8489 ( \8866 , \8865 , \545 );
nor \U$8490 ( \8867 , \8866 , \618 );
not \U$8491 ( \8868 , \8867 );
not \U$8492 ( \8869 , \4084 );
or \U$8493 ( \8870 , \8868 , \8869 );
not \U$8494 ( \8871 , \8866 );
and \U$8495 ( \8872 , \8871 , \8797 );
not \U$8496 ( \8873 , \545 );
not \U$8497 ( \8874 , \675 );
or \U$8498 ( \8875 , \8873 , \8874 );
nand \U$8499 ( \8876 , \8875 , \679 );
nor \U$8500 ( \8877 , \8872 , \8876 );
nand \U$8501 ( \8878 , \8870 , \8877 );
nor \U$8502 ( \8879 , \682 , \634 );
and \U$8503 ( \8880 , \8878 , \8879 );
not \U$8504 ( \8881 , \8878 );
not \U$8505 ( \8882 , \8879 );
and \U$8506 ( \8883 , \8881 , \8882 );
nor \U$8507 ( \8884 , \8880 , \8883 );
buf \U$8508 ( \8885 , \8884 );
buf \U$8509 ( \8886 , \8885 );
not \U$8510 ( \8887 , \8886 );
not \U$8511 ( \8888 , \8887 );
or \U$8512 ( \8889 , \8864 , \8888 );
nand \U$8513 ( \8890 , \8886 , \1302 );
nand \U$8514 ( \8891 , \8889 , \8890 );
nand \U$8515 ( \8892 , \8891 , \1311 );
nand \U$8516 ( \8893 , \8863 , \8892 );
xor \U$8517 ( \8894 , \8838 , \8893 );
not \U$8518 ( \8895 , \954 );
not \U$8519 ( \8896 , RIc2273d0_5);
not \U$8520 ( \8897 , \543 );
not \U$8521 ( \8898 , \8897 );
not \U$8522 ( \8899 , \4084 );
or \U$8523 ( \8900 , \8898 , \8899 );
nand \U$8524 ( \8901 , \8900 , \600 );
not \U$8525 ( \8902 , \599 );
nand \U$8526 ( \8903 , \8902 , \607 );
not \U$8527 ( \8904 , \8903 );
and \U$8528 ( \8905 , \8901 , \8904 );
not \U$8529 ( \8906 , \8901 );
and \U$8530 ( \8907 , \8906 , \8903 );
nor \U$8531 ( \8908 , \8905 , \8907 );
not \U$8532 ( \8909 , \8908 );
buf \U$8533 ( \8910 , \8909 );
not \U$8534 ( \8911 , \8910 );
or \U$8535 ( \8912 , \8896 , \8911 );
not \U$8536 ( \8913 , \8909 );
nand \U$8537 ( \8914 , \8913 , \935 );
nand \U$8538 ( \8915 , \8912 , \8914 );
not \U$8539 ( \8916 , \8915 );
or \U$8540 ( \8917 , \8895 , \8916 );
not \U$8541 ( \8918 , RIc2273d0_5);
not \U$8542 ( \8919 , \4084 );
and \U$8543 ( \8920 , \8897 , \600 );
or \U$8544 ( \8921 , \8919 , \8920 );
nand \U$8545 ( \8922 , \8919 , \8920 );
nand \U$8546 ( \8923 , \8921 , \8922 );
buf \U$8547 ( \8924 , \8923 );
not \U$8548 ( \8925 , \8924 );
not \U$8549 ( \8926 , \8925 );
or \U$8550 ( \8927 , \8918 , \8926 );
nand \U$8551 ( \8928 , \8924 , \946 );
nand \U$8552 ( \8929 , \8927 , \8928 );
nand \U$8553 ( \8930 , \8929 , \950 );
nand \U$8554 ( \8931 , \8917 , \8930 );
not \U$8555 ( \8932 , \1120 );
not \U$8556 ( \8933 , RIc2272e0_7);
not \U$8557 ( \8934 , \534 );
nand \U$8558 ( \8935 , \8897 , \8902 );
nor \U$8559 ( \8936 , \8934 , \8935 );
not \U$8560 ( \8937 , \8936 );
not \U$8561 ( \8938 , \4084 );
or \U$8562 ( \8939 , \8937 , \8938 );
nand \U$8563 ( \8940 , \4097 , \607 );
and \U$8564 ( \8941 , \8940 , \534 );
not \U$8565 ( \8942 , \608 );
nor \U$8566 ( \8943 , \8941 , \8942 );
nand \U$8567 ( \8944 , \8939 , \8943 );
nand \U$8568 ( \8945 , \621 , \595 );
not \U$8569 ( \8946 , \8945 );
and \U$8570 ( \8947 , \8944 , \8946 );
not \U$8571 ( \8948 , \8944 );
and \U$8572 ( \8949 , \8948 , \8945 );
nor \U$8573 ( \8950 , \8947 , \8949 );
buf \U$8574 ( \8951 , \8950 );
buf \U$8575 ( \8952 , \8951 );
not \U$8576 ( \8953 , \8952 );
not \U$8577 ( \8954 , \8953 );
or \U$8578 ( \8955 , \8933 , \8954 );
nand \U$8579 ( \8956 , \8952 , \4241 );
nand \U$8580 ( \8957 , \8955 , \8956 );
not \U$8581 ( \8958 , \8957 );
or \U$8582 ( \8959 , \8932 , \8958 );
not \U$8583 ( \8960 , RIc2272e0_7);
not \U$8584 ( \8961 , \8935 );
not \U$8585 ( \8962 , \8961 );
not \U$8586 ( \8963 , \4084 );
or \U$8587 ( \8964 , \8962 , \8963 );
not \U$8588 ( \8965 , \8940 );
nand \U$8589 ( \8966 , \8964 , \8965 );
and \U$8590 ( \8967 , \534 , \608 );
and \U$8591 ( \8968 , \8966 , \8967 );
not \U$8592 ( \8969 , \8966 );
not \U$8593 ( \8970 , \8967 );
and \U$8594 ( \8971 , \8969 , \8970 );
nor \U$8595 ( \8972 , \8968 , \8971 );
not \U$8596 ( \8973 , \8972 );
not \U$8597 ( \8974 , \8973 );
not \U$8598 ( \8975 , \8974 );
not \U$8599 ( \8976 , \8975 );
or \U$8600 ( \8977 , \8960 , \8976 );
not \U$8601 ( \8978 , \8972 );
not \U$8602 ( \8979 , \8978 );
nand \U$8603 ( \8980 , \8979 , \4241 );
nand \U$8604 ( \8981 , \8977 , \8980 );
nand \U$8605 ( \8982 , \8981 , \1118 );
nand \U$8606 ( \8983 , \8959 , \8982 );
xor \U$8607 ( \8984 , \8931 , \8983 );
not \U$8608 ( \8985 , \6689 );
not \U$8609 ( \8986 , RIc2263e0_39);
not \U$8610 ( \8987 , \3092 );
or \U$8611 ( \8988 , \8986 , \8987 );
not \U$8612 ( \8989 , \3091 );
not \U$8613 ( \8990 , RIc2263e0_39);
nand \U$8614 ( \8991 , \8989 , \8990 );
nand \U$8615 ( \8992 , \8988 , \8991 );
not \U$8616 ( \8993 , \8992 );
or \U$8617 ( \8994 , \8985 , \8993 );
not \U$8618 ( \8995 , RIc2263e0_39);
not \U$8619 ( \8996 , \4473 );
or \U$8620 ( \8997 , \8995 , \8996 );
not \U$8621 ( \8998 , RIc2263e0_39);
nand \U$8622 ( \8999 , \2344 , \8998 );
nand \U$8623 ( \9000 , \8997 , \8999 );
nand \U$8624 ( \9001 , \9000 , \6307 );
nand \U$8625 ( \9002 , \8994 , \9001 );
xor \U$8626 ( \9003 , \8984 , \9002 );
xor \U$8627 ( \9004 , \8894 , \9003 );
not \U$8628 ( \9005 , \954 );
not \U$8629 ( \9006 , RIc2273d0_5);
not \U$8630 ( \9007 , \504 );
buf \U$8631 ( \9008 , \466 );
nor \U$8632 ( \9009 , \9007 , \9008 );
not \U$8633 ( \9010 , \9009 );
buf \U$8634 ( \9011 , \562 );
nor \U$8635 ( \9012 , \9010 , \9011 );
not \U$8636 ( \9013 , \9012 );
not \U$8637 ( \9014 , \573 );
not \U$8638 ( \9015 , \518 );
nor \U$8639 ( \9016 , \9014 , \9015 );
not \U$8640 ( \9017 , \9016 );
not \U$8641 ( \9018 , \502 );
or \U$8642 ( \9019 , \9017 , \9018 );
not \U$8643 ( \9020 , \583 );
nand \U$8644 ( \9021 , \9019 , \9020 );
not \U$8645 ( \9022 , \9021 );
or \U$8646 ( \9023 , \9013 , \9022 );
not \U$8647 ( \9024 , \9009 );
not \U$8648 ( \9025 , \474 );
nand \U$8649 ( \9026 , \9025 , \457 );
not \U$8650 ( \9027 , \455 );
or \U$8651 ( \9028 , \9026 , \9027 );
not \U$8652 ( \9029 , \474 );
not \U$8653 ( \9030 , \448 );
and \U$8654 ( \9031 , \9029 , \9030 );
not \U$8655 ( \9032 , \447 );
nor \U$8656 ( \9033 , \9031 , \9032 );
nand \U$8657 ( \9034 , \9028 , \9033 );
not \U$8658 ( \9035 , \9034 );
or \U$8659 ( \9036 , \9024 , \9035 );
buf \U$8660 ( \9037 , \591 );
and \U$8661 ( \9038 , \9037 , \504 );
and \U$8662 ( \9039 , RIc2240b8_114, RIc22ac88_178);
nor \U$8663 ( \9040 , \9038 , \9039 );
nand \U$8664 ( \9041 , \9036 , \9040 );
not \U$8665 ( \9042 , \9041 );
nand \U$8666 ( \9043 , \9023 , \9042 );
nand \U$8667 ( \9044 , \510 , \596 );
xnor \U$8668 ( \9045 , \9043 , \9044 );
not \U$8669 ( \9046 , \9045 );
not \U$8670 ( \9047 , \9046 );
or \U$8671 ( \9048 , \9006 , \9047 );
not \U$8672 ( \9049 , \9045 );
not \U$8673 ( \9050 , \9049 );
buf \U$8674 ( \9051 , \9050 );
nand \U$8675 ( \9052 , \9051 , \956 );
nand \U$8676 ( \9053 , \9048 , \9052 );
not \U$8677 ( \9054 , \9053 );
or \U$8678 ( \9055 , \9005 , \9054 );
not \U$8679 ( \9056 , RIc2273d0_5);
nor \U$8680 ( \9057 , \9011 , \9008 );
not \U$8681 ( \9058 , \9057 );
not \U$8682 ( \9059 , \9021 );
or \U$8683 ( \9060 , \9058 , \9059 );
not \U$8684 ( \9061 , \9034 );
or \U$8685 ( \9062 , \9061 , \9008 );
not \U$8686 ( \9063 , \9037 );
nand \U$8687 ( \9064 , \9062 , \9063 );
not \U$8688 ( \9065 , \9064 );
nand \U$8689 ( \9066 , \9060 , \9065 );
not \U$8690 ( \9067 , \9039 );
nand \U$8691 ( \9068 , \9067 , \504 );
or \U$8692 ( \9069 , \9066 , \9068 );
nand \U$8693 ( \9070 , \9066 , \9068 );
nand \U$8694 ( \9071 , \9069 , \9070 );
buf \U$8695 ( \9072 , \9071 );
not \U$8696 ( \9073 , \9072 );
not \U$8697 ( \9074 , \9073 );
or \U$8698 ( \9075 , \9056 , \9074 );
not \U$8699 ( \9076 , \9071 );
not \U$8700 ( \9077 , \9076 );
nand \U$8701 ( \9078 , \9077 , \956 );
nand \U$8702 ( \9079 , \9075 , \9078 );
nand \U$8703 ( \9080 , \9079 , \951 );
nand \U$8704 ( \9081 , \9055 , \9080 );
not \U$8705 ( \9082 , \2138 );
not \U$8706 ( \9083 , RIc226980_27);
not \U$8707 ( \9084 , \3798 );
or \U$8708 ( \9085 , \9083 , \9084 );
nand \U$8709 ( \9086 , \2730 , \2133 );
nand \U$8710 ( \9087 , \9085 , \9086 );
not \U$8711 ( \9088 , \9087 );
or \U$8712 ( \9089 , \9082 , \9088 );
not \U$8713 ( \9090 , RIc226980_27);
not \U$8714 ( \9091 , \2063 );
or \U$8715 ( \9092 , \9090 , \9091 );
nand \U$8716 ( \9093 , \3008 , \2150 );
nand \U$8717 ( \9094 , \9092 , \9093 );
nand \U$8718 ( \9095 , \9094 , \2154 );
nand \U$8719 ( \9096 , \9089 , \9095 );
xor \U$8720 ( \9097 , \9081 , \9096 );
and \U$8721 ( \9098 , RIc226188_44, RIc226110_45);
not \U$8722 ( \9099 , RIc226188_44);
not \U$8723 ( \9100 , RIc226110_45);
and \U$8724 ( \9101 , \9099 , \9100 );
nor \U$8725 ( \9102 , \9098 , \9101 );
not \U$8726 ( \9103 , \9102 );
and \U$8727 ( \9104 , RIc226188_44, RIc226200_43);
not \U$8728 ( \9105 , RIc226188_44);
not \U$8729 ( \9106 , RIc226200_43);
and \U$8730 ( \9107 , \9105 , \9106 );
nor \U$8731 ( \9108 , \9104 , \9107 );
nand \U$8732 ( \9109 , \9103 , \9108 );
not \U$8733 ( \9110 , \9109 );
not \U$8734 ( \9111 , \9110 );
not \U$8735 ( \9112 , RIc226200_43);
not \U$8736 ( \9113 , \1487 );
or \U$8737 ( \9114 , \9112 , \9113 );
not \U$8738 ( \9115 , \1485 );
not \U$8739 ( \9116 , \9115 );
not \U$8740 ( \9117 , RIc226200_43);
nand \U$8741 ( \9118 , \9116 , \9117 );
nand \U$8742 ( \9119 , \9114 , \9118 );
not \U$8743 ( \9120 , \9119 );
or \U$8744 ( \9121 , \9111 , \9120 );
not \U$8745 ( \9122 , RIc226200_43);
not \U$8746 ( \9123 , \3438 );
or \U$8747 ( \9124 , \9122 , \9123 );
not \U$8748 ( \9125 , RIc226200_43);
nand \U$8749 ( \9126 , \1331 , \9125 );
nand \U$8750 ( \9127 , \9124 , \9126 );
buf \U$8751 ( \9128 , \9102 );
buf \U$8752 ( \9129 , \9128 );
nand \U$8753 ( \9130 , \9127 , \9129 );
nand \U$8754 ( \9131 , \9121 , \9130 );
and \U$8755 ( \9132 , \9097 , \9131 );
and \U$8756 ( \9133 , \9081 , \9096 );
or \U$8757 ( \9134 , \9132 , \9133 );
xor \U$8758 ( \9135 , \9004 , \9134 );
not \U$8759 ( \9136 , \9135 );
and \U$8760 ( \9137 , RIc226890_29, \3810 );
not \U$8761 ( \9138 , RIc226890_29);
not \U$8762 ( \9139 , \2670 );
and \U$8763 ( \9140 , \9138 , \9139 );
or \U$8764 ( \9141 , \9137 , \9140 );
buf \U$8765 ( \9142 , \2086 );
and \U$8766 ( \9143 , \9141 , \9142 );
not \U$8767 ( \9144 , RIc226890_29);
not \U$8768 ( \9145 , \9144 );
not \U$8769 ( \9146 , \2064 );
or \U$8770 ( \9147 , \9145 , \9146 );
not \U$8771 ( \9148 , \3008 );
nand \U$8772 ( \9149 , \9148 , RIc226890_29);
nand \U$8773 ( \9150 , \9147 , \9149 );
and \U$8774 ( \9151 , \9150 , \2784 );
nor \U$8775 ( \9152 , \9143 , \9151 );
not \U$8776 ( \9153 , \9152 );
not \U$8777 ( \9154 , \2697 );
not \U$8778 ( \9155 , RIc2267a0_31);
not \U$8779 ( \9156 , \2894 );
or \U$8780 ( \9157 , \9155 , \9156 );
not \U$8781 ( \9158 , \3021 );
not \U$8782 ( \9159 , RIc2267a0_31);
nand \U$8783 ( \9160 , \9158 , \9159 );
nand \U$8784 ( \9161 , \9157 , \9160 );
not \U$8785 ( \9162 , \9161 );
or \U$8786 ( \9163 , \9154 , \9162 );
not \U$8787 ( \9164 , RIc2267a0_31);
not \U$8788 ( \9165 , \5819 );
or \U$8789 ( \9166 , \9164 , \9165 );
nand \U$8790 ( \9167 , \2479 , \2705 );
nand \U$8791 ( \9168 , \9166 , \9167 );
nand \U$8792 ( \9169 , \9168 , \2711 );
nand \U$8793 ( \9170 , \9163 , \9169 );
not \U$8794 ( \9171 , \9170 );
not \U$8795 ( \9172 , \9171 );
or \U$8796 ( \9173 , \9153 , \9172 );
not \U$8797 ( \9174 , \9081 );
nand \U$8798 ( \9175 , \9173 , \9174 );
not \U$8799 ( \9176 , \9152 );
nand \U$8800 ( \9177 , \9176 , \9170 );
nand \U$8801 ( \9178 , \9175 , \9177 );
xor \U$8802 ( \9179 , \9081 , \9096 );
xor \U$8803 ( \9180 , \9179 , \9131 );
or \U$8804 ( \9181 , \9178 , \9180 );
not \U$8805 ( \9182 , \2154 );
not \U$8806 ( \9183 , \9087 );
or \U$8807 ( \9184 , \9182 , \9183 );
not \U$8808 ( \9185 , RIc226980_27);
not \U$8809 ( \9186 , \2635 );
or \U$8810 ( \9187 , \9185 , \9186 );
not \U$8811 ( \9188 , \2634 );
not \U$8812 ( \9189 , \9188 );
nand \U$8813 ( \9190 , \9189 , \2133 );
nand \U$8814 ( \9191 , \9187 , \9190 );
nand \U$8815 ( \9192 , \9191 , \2138 );
nand \U$8816 ( \9193 , \9184 , \9192 );
not \U$8817 ( \9194 , \9110 );
not \U$8818 ( \9195 , RIc226200_43);
not \U$8819 ( \9196 , \4181 );
not \U$8820 ( \9197 , \9196 );
not \U$8821 ( \9198 , \9197 );
or \U$8822 ( \9199 , \9195 , \9198 );
not \U$8823 ( \9200 , \4177 );
nand \U$8824 ( \9201 , \9200 , \9117 );
nand \U$8825 ( \9202 , \9199 , \9201 );
not \U$8826 ( \9203 , \9202 );
or \U$8827 ( \9204 , \9194 , \9203 );
buf \U$8828 ( \9205 , \9129 );
nand \U$8829 ( \9206 , \9119 , \9205 );
nand \U$8830 ( \9207 , \9204 , \9206 );
nor \U$8831 ( \9208 , \9193 , \9207 );
not \U$8832 ( \9209 , \1120 );
not \U$8833 ( \9210 , RIc2272e0_7);
buf \U$8834 ( \9211 , \8924 );
not \U$8835 ( \9212 , \9211 );
not \U$8836 ( \9213 , \9212 );
or \U$8837 ( \9214 , \9210 , \9213 );
not \U$8838 ( \9215 , \8924 );
not \U$8839 ( \9216 , \9215 );
nand \U$8840 ( \9217 , \9216 , \940 );
nand \U$8841 ( \9218 , \9214 , \9217 );
not \U$8842 ( \9219 , \9218 );
or \U$8843 ( \9220 , \9209 , \9219 );
not \U$8844 ( \9221 , RIc2272e0_7);
not \U$8845 ( \9222 , \9046 );
or \U$8846 ( \9223 , \9221 , \9222 );
not \U$8847 ( \9224 , \9045 );
not \U$8848 ( \9225 , \9224 );
nand \U$8849 ( \9226 , \9225 , \1139 );
nand \U$8850 ( \9227 , \9223 , \9226 );
nand \U$8851 ( \9228 , \9227 , \1118 );
nand \U$8852 ( \9229 , \9220 , \9228 );
not \U$8853 ( \9230 , \9229 );
not \U$8854 ( \9231 , \1082 );
not \U$8855 ( \9232 , RIc2274c0_3);
nand \U$8856 ( \9233 , RIc223fc8_116, RIc22ad78_180);
nand \U$8857 ( \9234 , \505 , \9233 );
not \U$8858 ( \9235 , \9234 );
not \U$8859 ( \9236 , \9011 );
not \U$8860 ( \9237 , \9236 );
buf \U$8861 ( \9238 , \9021 );
not \U$8862 ( \9239 , \9238 );
or \U$8863 ( \9240 , \9237 , \9239 );
nand \U$8864 ( \9241 , \9240 , \9061 );
not \U$8865 ( \9242 , \9241 );
or \U$8866 ( \9243 , \9235 , \9242 );
not \U$8867 ( \9244 , \9236 );
not \U$8868 ( \9245 , \9238 );
or \U$8869 ( \9246 , \9244 , \9245 );
nand \U$8870 ( \9247 , \9246 , \9061 );
or \U$8871 ( \9248 , \9247 , \9234 );
nand \U$8872 ( \9249 , \9243 , \9248 );
not \U$8873 ( \9250 , \9249 );
buf \U$8874 ( \9251 , \9250 );
not \U$8875 ( \9252 , \9251 );
or \U$8876 ( \9253 , \9232 , \9252 );
buf \U$8877 ( \9254 , \9249 );
not \U$8878 ( \9255 , \9254 );
not \U$8879 ( \9256 , \9255 );
nand \U$8880 ( \9257 , \9256 , \2896 );
nand \U$8881 ( \9258 , \9253 , \9257 );
not \U$8882 ( \9259 , \9258 );
or \U$8883 ( \9260 , \9231 , \9259 );
not \U$8884 ( \9261 , RIc2274c0_3);
and \U$8885 ( \9262 , \560 , \457 );
not \U$8886 ( \9263 , \9262 );
not \U$8887 ( \9264 , \9021 );
or \U$8888 ( \9265 , \9263 , \9264 );
and \U$8889 ( \9266 , \458 , \448 );
nand \U$8890 ( \9267 , \9265 , \9266 );
and \U$8891 ( \9268 , \9025 , \447 );
and \U$8892 ( \9269 , \9267 , \9268 );
not \U$8893 ( \9270 , \9267 );
not \U$8894 ( \9271 , \9268 );
and \U$8895 ( \9272 , \9270 , \9271 );
nor \U$8896 ( \9273 , \9269 , \9272 );
buf \U$8897 ( \9274 , \9273 );
buf \U$8898 ( \9275 , \9274 );
not \U$8899 ( \9276 , \9275 );
not \U$8900 ( \9277 , \9276 );
or \U$8901 ( \9278 , \9261 , \9277 );
nand \U$8902 ( \9279 , \9275 , \2896 );
nand \U$8903 ( \9280 , \9278 , \9279 );
nand \U$8904 ( \9281 , \9280 , \1040 );
nand \U$8905 ( \9282 , \9260 , \9281 );
not \U$8906 ( \9283 , \9282 );
nand \U$8907 ( \9284 , \9230 , \9283 );
not \U$8908 ( \9285 , \1579 );
nand \U$8909 ( \9286 , \457 , \448 );
not \U$8910 ( \9287 , \9286 );
not \U$8911 ( \9288 , \560 );
not \U$8912 ( \9289 , \9021 );
or \U$8913 ( \9290 , \9288 , \9289 );
buf \U$8914 ( \9291 , \9027 );
nand \U$8915 ( \9292 , \9290 , \9291 );
not \U$8916 ( \9293 , \9292 );
or \U$8917 ( \9294 , \9287 , \9293 );
or \U$8918 ( \9295 , \9292 , \9286 );
nand \U$8919 ( \9296 , \9294 , \9295 );
not \U$8920 ( \9297 , \9296 );
not \U$8921 ( \9298 , \9297 );
buf \U$8922 ( \9299 , \9298 );
not \U$8923 ( \9300 , \9299 );
and \U$8924 ( \9301 , RIc2275b0_1, \9300 );
not \U$8925 ( \9302 , RIc2275b0_1);
and \U$8926 ( \9303 , \9302 , \9299 );
or \U$8927 ( \9304 , \9301 , \9303 );
not \U$8928 ( \9305 , \9304 );
or \U$8929 ( \9306 , \9285 , \9305 );
not \U$8930 ( \9307 , \451 );
nand \U$8931 ( \9308 , \9307 , \454 );
not \U$8932 ( \9309 , \9308 );
not \U$8933 ( \9310 , \512 );
not \U$8934 ( \9311 , \9310 );
not \U$8935 ( \9312 , \9021 );
or \U$8936 ( \9313 , \9311 , \9312 );
buf \U$8937 ( \9314 , \452 );
nand \U$8938 ( \9315 , \9313 , \9314 );
not \U$8939 ( \9316 , \9315 );
or \U$8940 ( \9317 , \9309 , \9316 );
or \U$8941 ( \9318 , \9315 , \9308 );
nand \U$8942 ( \9319 , \9317 , \9318 );
buf \U$8943 ( \9320 , \9319 );
not \U$8944 ( \9321 , \9320 );
and \U$8945 ( \9322 , RIc2275b0_1, \9321 );
not \U$8946 ( \9323 , RIc2275b0_1);
buf \U$8947 ( \9324 , \9319 );
and \U$8948 ( \9325 , \9323 , \9324 );
or \U$8949 ( \9326 , \9322 , \9325 );
nand \U$8950 ( \9327 , \9326 , \854 );
nand \U$8951 ( \9328 , \9306 , \9327 );
and \U$8952 ( \9329 , \9284 , \9328 );
and \U$8953 ( \9330 , \9229 , \9282 );
nor \U$8954 ( \9331 , \9329 , \9330 );
or \U$8955 ( \9332 , \9208 , \9331 );
nand \U$8956 ( \9333 , \9193 , \9207 );
nand \U$8957 ( \9334 , \9332 , \9333 );
nand \U$8958 ( \9335 , \9181 , \9334 );
nand \U$8959 ( \9336 , \9180 , \9178 );
and \U$8960 ( \9337 , \9335 , \9336 );
not \U$8961 ( \9338 , \9337 );
not \U$8962 ( \9339 , \9338 );
or \U$8963 ( \9340 , \9136 , \9339 );
not \U$8964 ( \9341 , \9337 );
not \U$8965 ( \9342 , \9135 );
not \U$8966 ( \9343 , \9342 );
or \U$8967 ( \9344 , \9341 , \9343 );
not \U$8968 ( \9345 , \2784 );
not \U$8969 ( \9346 , \9141 );
or \U$8970 ( \9347 , \9345 , \9346 );
not \U$8971 ( \9348 , RIc226890_29);
not \U$8972 ( \9349 , \3021 );
or \U$8973 ( \9350 , \9348 , \9349 );
not \U$8974 ( \9351 , RIc226890_29);
nand \U$8975 ( \9352 , \9351 , \2498 );
nand \U$8976 ( \9353 , \9350 , \9352 );
nand \U$8977 ( \9354 , \9353 , \2086 );
nand \U$8978 ( \9355 , \9347 , \9354 );
not \U$8979 ( \9356 , \2697 );
not \U$8980 ( \9357 , \9168 );
or \U$8981 ( \9358 , \9356 , \9357 );
not \U$8982 ( \9359 , RIc2267a0_31);
not \U$8983 ( \9360 , \2554 );
not \U$8984 ( \9361 , \9360 );
not \U$8985 ( \9362 , \9361 );
or \U$8986 ( \9363 , \9359 , \9362 );
not \U$8987 ( \9364 , \4802 );
nand \U$8988 ( \9365 , \9364 , \2705 );
nand \U$8989 ( \9366 , \9363 , \9365 );
nand \U$8990 ( \9367 , \9366 , \2710 );
nand \U$8991 ( \9368 , \9358 , \9367 );
not \U$8992 ( \9369 , \9368 );
xor \U$8993 ( \9370 , \9355 , \9369 );
and \U$8994 ( \9371 , RIc226098_46, RIc226020_47);
not \U$8995 ( \9372 , RIc226098_46);
not \U$8996 ( \9373 , RIc226020_47);
and \U$8997 ( \9374 , \9372 , \9373 );
nor \U$8998 ( \9375 , \9371 , \9374 );
not \U$8999 ( \9376 , \9375 );
and \U$9000 ( \9377 , RIc226098_46, RIc226110_45);
not \U$9001 ( \9378 , RIc226098_46);
not \U$9002 ( \9379 , RIc226110_45);
and \U$9003 ( \9380 , \9378 , \9379 );
nor \U$9004 ( \9381 , \9377 , \9380 );
and \U$9005 ( \9382 , \9376 , \9381 );
not \U$9006 ( \9383 , \9382 );
not \U$9007 ( \9384 , \9383 );
not \U$9008 ( \9385 , \9384 );
not \U$9009 ( \9386 , RIc226110_45);
not \U$9010 ( \9387 , \3580 );
or \U$9011 ( \9388 , \9386 , \9387 );
nand \U$9012 ( \9389 , \4595 , \9379 );
nand \U$9013 ( \9390 , \9388 , \9389 );
not \U$9014 ( \9391 , \9390 );
or \U$9015 ( \9392 , \9385 , \9391 );
not \U$9016 ( \9393 , RIc226110_45);
not \U$9017 ( \9394 , \1392 );
or \U$9018 ( \9395 , \9393 , \9394 );
nand \U$9019 ( \9396 , \5246 , \9100 );
nand \U$9020 ( \9397 , \9395 , \9396 );
buf \U$9021 ( \9398 , \9375 );
nand \U$9022 ( \9399 , \9397 , \9398 );
nand \U$9023 ( \9400 , \9392 , \9399 );
xor \U$9024 ( \9401 , \9370 , \9400 );
not \U$9025 ( \9402 , \9401 );
not \U$9026 ( \9403 , \9402 );
not \U$9027 ( \9404 , \5741 );
not \U$9028 ( \9405 , RIc2265c0_35);
not \U$9029 ( \9406 , \1989 );
or \U$9030 ( \9407 , \9405 , \9406 );
not \U$9031 ( \9408 , \1988 );
not \U$9032 ( \9409 , \9408 );
nand \U$9033 ( \9410 , \9409 , \4376 );
nand \U$9034 ( \9411 , \9407 , \9410 );
not \U$9035 ( \9412 , \9411 );
or \U$9036 ( \9413 , \9404 , \9412 );
not \U$9037 ( \9414 , RIc2265c0_35);
not \U$9038 ( \9415 , \2257 );
or \U$9039 ( \9416 , \9414 , \9415 );
nand \U$9040 ( \9417 , \4008 , \3620 );
nand \U$9041 ( \9418 , \9416 , \9417 );
nand \U$9042 ( \9419 , \9418 , \4383 );
nand \U$9043 ( \9420 , \9413 , \9419 );
not \U$9044 ( \9421 , \3629 );
not \U$9045 ( \9422 , \2585 );
and \U$9046 ( \9423 , \9422 , RIc2266b0_33);
not \U$9047 ( \9424 , \9422 );
not \U$9048 ( \9425 , RIc2266b0_33);
and \U$9049 ( \9426 , \9424 , \9425 );
or \U$9050 ( \9427 , \9423 , \9426 );
not \U$9051 ( \9428 , \9427 );
or \U$9052 ( \9429 , \9421 , \9428 );
not \U$9053 ( \9430 , RIc2266b0_33);
not \U$9054 ( \9431 , \3509 );
or \U$9055 ( \9432 , \9430 , \9431 );
not \U$9056 ( \9433 , \2013 );
not \U$9057 ( \9434 , \9433 );
nand \U$9058 ( \9435 , \9434 , \2692 );
nand \U$9059 ( \9436 , \9432 , \9435 );
nand \U$9060 ( \9437 , \9436 , \3631 );
nand \U$9061 ( \9438 , \9429 , \9437 );
xor \U$9062 ( \9439 , \9420 , \9438 );
and \U$9063 ( \9440 , RIc225dc8_52, RIc225d50_53);
not \U$9064 ( \9441 , RIc225dc8_52);
and \U$9065 ( \9442 , \9441 , \8782 );
nor \U$9066 ( \9443 , \9440 , \9442 );
buf \U$9067 ( \9444 , \9443 );
buf \U$9068 ( \9445 , \9444 );
not \U$9069 ( \9446 , \9445 );
not \U$9070 ( \9447 , RIc225e40_51);
not \U$9071 ( \9448 , \4024 );
or \U$9072 ( \9449 , \9447 , \9448 );
not \U$9073 ( \9450 , RIc225e40_51);
nand \U$9074 ( \9451 , \889 , \9450 );
nand \U$9075 ( \9452 , \9449 , \9451 );
not \U$9076 ( \9453 , \9452 );
or \U$9077 ( \9454 , \9446 , \9453 );
and \U$9078 ( \9455 , RIc225e40_51, RIc225dc8_52);
nor \U$9079 ( \9456 , RIc225e40_51, RIc225dc8_52);
nor \U$9080 ( \9457 , \9455 , \9443 , \9456 );
buf \U$9081 ( \9458 , \9457 );
buf \U$9082 ( \9459 , \9458 );
and \U$9083 ( \9460 , RIc225e40_51, \4608 );
not \U$9084 ( \9461 , RIc225e40_51);
and \U$9085 ( \9462 , \9461 , \840 );
or \U$9086 ( \9463 , \9460 , \9462 );
nand \U$9087 ( \9464 , \9459 , \9463 );
nand \U$9088 ( \9465 , \9454 , \9464 );
and \U$9089 ( \9466 , \9439 , \9465 );
not \U$9090 ( \9467 , \9439 );
not \U$9091 ( \9468 , \9465 );
and \U$9092 ( \9469 , \9467 , \9468 );
nor \U$9093 ( \9470 , \9466 , \9469 );
not \U$9094 ( \9471 , \9470 );
or \U$9095 ( \9472 , \9403 , \9471 );
not \U$9096 ( \9473 , \9470 );
not \U$9097 ( \9474 , \9473 );
not \U$9098 ( \9475 , \9401 );
or \U$9099 ( \9476 , \9474 , \9475 );
not \U$9100 ( \9477 , \6688 );
not \U$9101 ( \9478 , RIc2263e0_39);
not \U$9102 ( \9479 , \2422 );
not \U$9103 ( \9480 , \9479 );
or \U$9104 ( \9481 , \9478 , \9480 );
nand \U$9105 ( \9482 , \4457 , \5498 );
nand \U$9106 ( \9483 , \9481 , \9482 );
not \U$9107 ( \9484 , \9483 );
or \U$9108 ( \9485 , \9477 , \9484 );
nand \U$9109 ( \9486 , \8992 , \6307 );
nand \U$9110 ( \9487 , \9485 , \9486 );
not \U$9111 ( \9488 , \8776 );
not \U$9112 ( \9489 , \9488 );
not \U$9113 ( \9490 , RIc225d50_53);
not \U$9114 ( \9491 , \1072 );
not \U$9115 ( \9492 , \9491 );
or \U$9116 ( \9493 , \9490 , \9492 );
nand \U$9117 ( \9494 , \1072 , \8782 );
nand \U$9118 ( \9495 , \9493 , \9494 );
not \U$9119 ( \9496 , \9495 );
or \U$9120 ( \9497 , \9489 , \9496 );
nand \U$9121 ( \9498 , \8784 , \8788 );
nand \U$9122 ( \9499 , \9497 , \9498 );
and \U$9123 ( \9500 , \9487 , \9499 );
not \U$9124 ( \9501 , \9487 );
not \U$9125 ( \9502 , \9499 );
and \U$9126 ( \9503 , \9501 , \9502 );
nor \U$9127 ( \9504 , \9500 , \9503 );
not \U$9128 ( \9505 , \1915 );
not \U$9129 ( \9506 , RIc226b60_23);
not \U$9130 ( \9507 , \3726 );
or \U$9131 ( \9508 , \9506 , \9507 );
nand \U$9132 ( \9509 , \2980 , \2111 );
nand \U$9133 ( \9510 , \9508 , \9509 );
not \U$9134 ( \9511 , \9510 );
or \U$9135 ( \9512 , \9505 , \9511 );
not \U$9136 ( \9513 , \3115 );
and \U$9137 ( \9514 , \5637 , \9513 );
not \U$9138 ( \9515 , \5637 );
and \U$9139 ( \9516 , \9515 , \3115 );
or \U$9140 ( \9517 , \9514 , \9516 );
not \U$9141 ( \9518 , \9517 );
nand \U$9142 ( \9519 , \9518 , \5365 );
nand \U$9143 ( \9520 , \9512 , \9519 );
xor \U$9144 ( \9521 , \9504 , \9520 );
nand \U$9145 ( \9522 , \9476 , \9521 );
nand \U$9146 ( \9523 , \9472 , \9522 );
nand \U$9147 ( \9524 , \9344 , \9523 );
nand \U$9148 ( \9525 , \9340 , \9524 );
and \U$9149 ( \9526 , RIc225f30_49, RIc225eb8_50);
and \U$9150 ( \9527 , RIc225eb8_50, RIc225e40_51);
not \U$9151 ( \9528 , RIc225eb8_50);
and \U$9152 ( \9529 , \9528 , \9450 );
nor \U$9153 ( \9530 , \9527 , \9529 );
nor \U$9154 ( \9531 , RIc225f30_49, RIc225eb8_50);
nor \U$9155 ( \9532 , \9526 , \9530 , \9531 );
not \U$9156 ( \9533 , \9532 );
not \U$9157 ( \9534 , \9533 );
not \U$9158 ( \9535 , \9534 );
not \U$9159 ( \9536 , RIc225f30_49);
not \U$9160 ( \9537 , \1402 );
or \U$9161 ( \9538 , \9536 , \9537 );
not \U$9162 ( \9539 , \1169 );
not \U$9163 ( \9540 , \9539 );
not \U$9164 ( \9541 , RIc225f30_49);
nand \U$9165 ( \9542 , \9540 , \9541 );
nand \U$9166 ( \9543 , \9538 , \9542 );
not \U$9167 ( \9544 , \9543 );
or \U$9168 ( \9545 , \9535 , \9544 );
not \U$9169 ( \9546 , RIc225f30_49);
not \U$9170 ( \9547 , \1021 );
or \U$9171 ( \9548 , \9546 , \9547 );
not \U$9172 ( \9549 , RIc225f30_49);
nand \U$9173 ( \9550 , \2119 , \9549 );
nand \U$9174 ( \9551 , \9548 , \9550 );
buf \U$9175 ( \9552 , \9530 );
nand \U$9176 ( \9553 , \9551 , \9552 );
nand \U$9177 ( \9554 , \9545 , \9553 );
buf \U$9178 ( \9555 , \8788 );
not \U$9179 ( \9556 , \9555 );
not \U$9180 ( \9557 , \9495 );
or \U$9181 ( \9558 , \9556 , \9557 );
and \U$9182 ( \9559 , RIc225d50_53, \4024 );
not \U$9183 ( \9560 , RIc225d50_53);
and \U$9184 ( \9561 , \9560 , \888 );
or \U$9185 ( \9562 , \9559 , \9561 );
nand \U$9186 ( \9563 , \9562 , \9488 );
nand \U$9187 ( \9564 , \9558 , \9563 );
or \U$9188 ( \9565 , \9554 , \9564 );
not \U$9189 ( \9566 , \6307 );
not \U$9190 ( \9567 , \9483 );
or \U$9191 ( \9568 , \9566 , \9567 );
not \U$9192 ( \9569 , RIc2263e0_39);
not \U$9193 ( \9570 , \2443 );
not \U$9194 ( \9571 , \9570 );
or \U$9195 ( \9572 , \9569 , \9571 );
not \U$9196 ( \9573 , RIc2263e0_39);
nand \U$9197 ( \9574 , \5949 , \9573 );
nand \U$9198 ( \9575 , \9572 , \9574 );
nand \U$9199 ( \9576 , \9575 , \6689 );
nand \U$9200 ( \9577 , \9568 , \9576 );
and \U$9201 ( \9578 , \9565 , \9577 );
and \U$9202 ( \9579 , \9564 , \9554 );
nor \U$9203 ( \9580 , \9578 , \9579 );
not \U$9204 ( \9581 , \9580 );
not \U$9205 ( \9582 , \5741 );
not \U$9206 ( \9583 , RIc2265c0_35);
not \U$9207 ( \9584 , \2013 );
not \U$9208 ( \9585 , \9584 );
or \U$9209 ( \9586 , \9583 , \9585 );
not \U$9210 ( \9587 , RIc2265c0_35);
nand \U$9211 ( \9588 , \3508 , \9587 );
nand \U$9212 ( \9589 , \9586 , \9588 );
not \U$9213 ( \9590 , \9589 );
or \U$9214 ( \9591 , \9582 , \9590 );
nand \U$9215 ( \9592 , \9411 , \5135 );
nand \U$9216 ( \9593 , \9591 , \9592 );
not \U$9217 ( \9594 , \9593 );
not \U$9218 ( \9595 , \5519 );
not \U$9219 ( \9596 , RIc2264d0_37);
not \U$9220 ( \9597 , \2227 );
or \U$9221 ( \9598 , \9596 , \9597 );
not \U$9222 ( \9599 , \2225 );
not \U$9223 ( \9600 , \9599 );
nand \U$9224 ( \9601 , \9600 , \5504 );
nand \U$9225 ( \9602 , \9598 , \9601 );
not \U$9226 ( \9603 , \9602 );
or \U$9227 ( \9604 , \9595 , \9603 );
not \U$9228 ( \9605 , RIc2264d0_37);
not \U$9229 ( \9606 , \2258 );
or \U$9230 ( \9607 , \9605 , \9606 );
not \U$9231 ( \9608 , \2257 );
nand \U$9232 ( \9609 , \9608 , \5514 );
nand \U$9233 ( \9610 , \9607 , \9609 );
nand \U$9234 ( \9611 , \9610 , \5509 );
nand \U$9235 ( \9612 , \9604 , \9611 );
not \U$9236 ( \9613 , \9612 );
nand \U$9237 ( \9614 , \9594 , \9613 );
and \U$9238 ( \9615 , RIc225fa8_48, RIc225f30_49);
not \U$9239 ( \9616 , RIc225fa8_48);
and \U$9240 ( \9617 , \9616 , \9549 );
nor \U$9241 ( \9618 , \9615 , \9617 );
buf \U$9242 ( \9619 , \9618 );
not \U$9243 ( \9620 , \9619 );
not \U$9244 ( \9621 , RIc226020_47);
not \U$9245 ( \9622 , \1372 );
or \U$9246 ( \9623 , \9621 , \9622 );
not \U$9247 ( \9624 , RIc226020_47);
nand \U$9248 ( \9625 , \2373 , \9624 );
nand \U$9249 ( \9626 , \9623 , \9625 );
not \U$9250 ( \9627 , \9626 );
or \U$9251 ( \9628 , \9620 , \9627 );
not \U$9252 ( \9629 , RIc226020_47);
not \U$9253 ( \9630 , \3496 );
or \U$9254 ( \9631 , \9629 , \9630 );
nand \U$9255 ( \9632 , \5246 , \9624 );
nand \U$9256 ( \9633 , \9631 , \9632 );
not \U$9257 ( \9634 , \9618 );
and \U$9258 ( \9635 , RIc225fa8_48, RIc226020_47);
not \U$9259 ( \9636 , RIc225fa8_48);
and \U$9260 ( \9637 , \9636 , \9624 );
nor \U$9261 ( \9638 , \9635 , \9637 );
and \U$9262 ( \9639 , \9634 , \9638 );
not \U$9263 ( \9640 , \9639 );
not \U$9264 ( \9641 , \9640 );
nand \U$9265 ( \9642 , \9633 , \9641 );
nand \U$9266 ( \9643 , \9628 , \9642 );
and \U$9267 ( \9644 , \9614 , \9643 );
nor \U$9268 ( \9645 , \9594 , \9613 );
nor \U$9269 ( \9646 , \9644 , \9645 );
not \U$9270 ( \9647 , \9646 );
or \U$9271 ( \9648 , \9581 , \9647 );
not \U$9272 ( \9649 , \2172 );
not \U$9273 ( \9650 , RIc226a70_25);
not \U$9274 ( \9651 , \4500 );
not \U$9275 ( \9652 , \9651 );
or \U$9276 ( \9653 , \9650 , \9652 );
buf \U$9277 ( \9654 , \2103 );
nand \U$9278 ( \9655 , \9654 , \1905 );
nand \U$9279 ( \9656 , \9653 , \9655 );
not \U$9280 ( \9657 , \9656 );
or \U$9281 ( \9658 , \9649 , \9657 );
not \U$9282 ( \9659 , RIc226a70_25);
not \U$9283 ( \9660 , \3116 );
or \U$9284 ( \9661 , \9659 , \9660 );
not \U$9285 ( \9662 , RIc226a70_25);
nand \U$9286 ( \9663 , \5160 , \9662 );
nand \U$9287 ( \9664 , \9661 , \9663 );
nand \U$9288 ( \9665 , \9664 , \2860 );
nand \U$9289 ( \9666 , \9658 , \9665 );
not \U$9290 ( \9667 , \9666 );
not \U$9291 ( \9668 , \1930 );
not \U$9292 ( \9669 , \9510 );
or \U$9293 ( \9670 , \9668 , \9669 );
not \U$9294 ( \9671 , RIc226b60_23);
not \U$9295 ( \9672 , \4049 );
or \U$9296 ( \9673 , \9671 , \9672 );
not \U$9297 ( \9674 , \3640 );
not \U$9298 ( \9675 , \9674 );
nand \U$9299 ( \9676 , \9675 , \2111 );
nand \U$9300 ( \9677 , \9673 , \9676 );
nand \U$9301 ( \9678 , \9677 , \1915 );
nand \U$9302 ( \9679 , \9670 , \9678 );
not \U$9303 ( \9680 , \9679 );
or \U$9304 ( \9681 , \9667 , \9680 );
or \U$9305 ( \9682 , \9679 , \9666 );
and \U$9306 ( \9683 , RIc2262f0_41, RIc226278_42);
and \U$9307 ( \9684 , RIc226278_42, RIc226200_43);
not \U$9308 ( \9685 , RIc226278_42);
and \U$9309 ( \9686 , \9685 , \9106 );
nor \U$9310 ( \9687 , \9684 , \9686 );
nor \U$9311 ( \9688 , RIc2262f0_41, RIc226278_42);
nor \U$9312 ( \9689 , \9683 , \9687 , \9688 );
buf \U$9313 ( \9690 , \9689 );
not \U$9314 ( \9691 , \9690 );
not \U$9315 ( \9692 , RIc2262f0_41);
not \U$9316 ( \9693 , \2298 );
or \U$9317 ( \9694 , \9692 , \9693 );
or \U$9318 ( \9695 , \3092 , RIc2262f0_41);
nand \U$9319 ( \9696 , \9694 , \9695 );
not \U$9320 ( \9697 , \9696 );
or \U$9321 ( \9698 , \9691 , \9697 );
not \U$9322 ( \9699 , RIc2262f0_41);
not \U$9323 ( \9700 , \2353 );
not \U$9324 ( \9701 , \9700 );
or \U$9325 ( \9702 , \9699 , \9701 );
nand \U$9326 ( \9703 , \2353 , \6303 );
nand \U$9327 ( \9704 , \9702 , \9703 );
buf \U$9328 ( \9705 , \9687 );
nand \U$9329 ( \9706 , \9704 , \9705 );
nand \U$9330 ( \9707 , \9698 , \9706 );
nand \U$9331 ( \9708 , \9682 , \9707 );
nand \U$9332 ( \9709 , \9681 , \9708 );
nand \U$9333 ( \9710 , \9648 , \9709 );
not \U$9334 ( \9711 , \9646 );
not \U$9335 ( \9712 , \9580 );
nand \U$9336 ( \9713 , \9711 , \9712 );
nand \U$9337 ( \9714 , \9710 , \9713 );
not \U$9338 ( \9715 , \9714 );
not \U$9339 ( \9716 , RIc227010_13);
not \U$9340 ( \9717 , \4086 );
not \U$9341 ( \9718 , \4084 );
or \U$9342 ( \9719 , \9717 , \9718 );
not \U$9343 ( \9720 , \4111 );
nand \U$9344 ( \9721 , \9719 , \9720 );
nand \U$9345 ( \9722 , \6702 , \6706 );
not \U$9346 ( \9723 , \9722 );
and \U$9347 ( \9724 , \9721 , \9723 );
not \U$9348 ( \9725 , \9721 );
and \U$9349 ( \9726 , \9725 , \9722 );
nor \U$9350 ( \9727 , \9724 , \9726 );
not \U$9351 ( \9728 , \9727 );
not \U$9352 ( \9729 , \9728 );
or \U$9353 ( \9730 , \9716 , \9729 );
buf \U$9354 ( \9731 , \9727 );
nand \U$9355 ( \9732 , \9731 , \3841 );
nand \U$9356 ( \9733 , \9730 , \9732 );
not \U$9357 ( \9734 , \9733 );
nor \U$9358 ( \9735 , \9734 , \1679 );
not \U$9359 ( \9736 , \1682 );
not \U$9360 ( \9737 , \6718 );
not \U$9361 ( \9738 , \1296 );
and \U$9362 ( \9739 , \9737 , \9738 );
buf \U$9363 ( \9740 , \6718 );
and \U$9364 ( \9741 , \9740 , \1296 );
nor \U$9365 ( \9742 , \9739 , \9741 );
nor \U$9366 ( \9743 , \9736 , \9742 );
nor \U$9367 ( \9744 , \9735 , \9743 );
not \U$9368 ( \9745 , \1945 );
not \U$9369 ( \9746 , RIc226e30_17);
not \U$9370 ( \9747 , \5664 );
or \U$9371 ( \9748 , \9746 , \9747 );
nand \U$9372 ( \9749 , \5663 , \1960 );
nand \U$9373 ( \9750 , \9748 , \9749 );
not \U$9374 ( \9751 , \9750 );
or \U$9375 ( \9752 , \9745 , \9751 );
not \U$9376 ( \9753 , RIc226e30_17);
not \U$9377 ( \9754 , \5215 );
not \U$9378 ( \9755 , \9754 );
or \U$9379 ( \9756 , \9753 , \9755 );
buf \U$9380 ( \9757 , \5215 );
nand \U$9381 ( \9758 , \9757 , \1935 );
nand \U$9382 ( \9759 , \9756 , \9758 );
nand \U$9383 ( \9760 , \9759 , \1963 );
nand \U$9384 ( \9761 , \9752 , \9760 );
not \U$9385 ( \9762 , \9761 );
xor \U$9386 ( \9763 , \9744 , \9762 );
not \U$9387 ( \9764 , RIc226f20_15);
not \U$9388 ( \9765 , \6071 );
not \U$9389 ( \9766 , \9765 );
or \U$9390 ( \9767 , \9764 , \9766 );
not \U$9391 ( \9768 , \6070 );
not \U$9392 ( \9769 , \9768 );
buf \U$9393 ( \9770 , \9769 );
nand \U$9394 ( \9771 , \9770 , \1674 );
nand \U$9395 ( \9772 , \9767 , \9771 );
and \U$9396 ( \9773 , \9772 , \2358 );
not \U$9397 ( \9774 , RIc226f20_15);
not \U$9398 ( \9775 , \6492 );
not \U$9399 ( \9776 , \9775 );
or \U$9400 ( \9777 , \9774 , \9776 );
nand \U$9401 ( \9778 , \6492 , \2301 );
nand \U$9402 ( \9779 , \9777 , \9778 );
not \U$9403 ( \9780 , \9779 );
nor \U$9404 ( \9781 , \9780 , \2321 );
nor \U$9405 ( \9782 , \9773 , \9781 );
xor \U$9406 ( \9783 , \9763 , \9782 );
not \U$9407 ( \9784 , \1118 );
not \U$9408 ( \9785 , RIc2272e0_7);
not \U$9409 ( \9786 , \8910 );
not \U$9410 ( \9787 , \9786 );
not \U$9411 ( \9788 , \9787 );
or \U$9412 ( \9789 , \9785 , \9788 );
not \U$9413 ( \9790 , \8910 );
nand \U$9414 ( \9791 , \9790 , \940 );
nand \U$9415 ( \9792 , \9789 , \9791 );
not \U$9416 ( \9793 , \9792 );
or \U$9417 ( \9794 , \9784 , \9793 );
nand \U$9418 ( \9795 , \8981 , \1120 );
nand \U$9419 ( \9796 , \9794 , \9795 );
not \U$9420 ( \9797 , \9796 );
not \U$9421 ( \9798 , \2195 );
not \U$9422 ( \9799 , \9656 );
or \U$9423 ( \9800 , \9798 , \9799 );
not \U$9424 ( \9801 , RIc226a70_25);
not \U$9425 ( \9802 , \2635 );
or \U$9426 ( \9803 , \9801 , \9802 );
not \U$9427 ( \9804 , \2634 );
not \U$9428 ( \9805 , \9804 );
nand \U$9429 ( \9806 , \9805 , \6107 );
nand \U$9430 ( \9807 , \9803 , \9806 );
nand \U$9431 ( \9808 , \9807 , \2173 );
nand \U$9432 ( \9809 , \9800 , \9808 );
not \U$9433 ( \9810 , \9809 );
or \U$9434 ( \9811 , \9797 , \9810 );
or \U$9435 ( \9812 , \9809 , \9796 );
not \U$9436 ( \9813 , \9690 );
not \U$9437 ( \9814 , \9704 );
or \U$9438 ( \9815 , \9813 , \9814 );
buf \U$9439 ( \9816 , \9705 );
not \U$9440 ( \9817 , \9816 );
not \U$9441 ( \9818 , \9817 );
not \U$9442 ( \9819 , RIc2262f0_41);
not \U$9443 ( \9820 , \4177 );
or \U$9444 ( \9821 , \9819 , \9820 );
not \U$9445 ( \9822 , RIc2262f0_41);
nand \U$9446 ( \9823 , \1729 , \9822 );
nand \U$9447 ( \9824 , \9821 , \9823 );
nand \U$9448 ( \9825 , \9818 , \9824 );
nand \U$9449 ( \9826 , \9815 , \9825 );
nand \U$9450 ( \9827 , \9812 , \9826 );
nand \U$9451 ( \9828 , \9811 , \9827 );
xor \U$9452 ( \9829 , \9783 , \9828 );
or \U$9453 ( \9830 , \9520 , \9487 );
nand \U$9454 ( \9831 , \9830 , \9499 );
nand \U$9455 ( \9832 , \9520 , \9487 );
nand \U$9456 ( \9833 , \9831 , \9832 );
not \U$9457 ( \9834 , \9833 );
xnor \U$9458 ( \9835 , \9829 , \9834 );
not \U$9459 ( \9836 , \9835 );
not \U$9460 ( \9837 , \9836 );
or \U$9461 ( \9838 , \9715 , \9837 );
or \U$9462 ( \9839 , \9836 , \9714 );
not \U$9463 ( \9840 , \2534 );
not \U$9464 ( \9841 , RIc226d40_19);
not \U$9465 ( \9842 , \4406 );
not \U$9466 ( \9843 , \9842 );
or \U$9467 ( \9844 , \9841 , \9843 );
nand \U$9468 ( \9845 , \4406 , \2523 );
nand \U$9469 ( \9846 , \9844 , \9845 );
not \U$9470 ( \9847 , \9846 );
or \U$9471 ( \9848 , \9840 , \9847 );
not \U$9472 ( \9849 , RIc226d40_19);
not \U$9473 ( \9850 , \5215 );
not \U$9474 ( \9851 , \9850 );
or \U$9475 ( \9852 , \9849 , \9851 );
nand \U$9476 ( \9853 , \5215 , \3338 );
nand \U$9477 ( \9854 , \9852 , \9853 );
nand \U$9478 ( \9855 , \9854 , \2518 );
nand \U$9479 ( \9856 , \9848 , \9855 );
not \U$9480 ( \9857 , \2320 );
not \U$9481 ( \9858 , RIc226f20_15);
not \U$9482 ( \9859 , \6718 );
not \U$9483 ( \9860 , \9859 );
or \U$9484 ( \9861 , \9858 , \9860 );
nand \U$9485 ( \9862 , \6718 , \1674 );
nand \U$9486 ( \9863 , \9861 , \9862 );
not \U$9487 ( \9864 , \9863 );
or \U$9488 ( \9865 , \9857 , \9864 );
nand \U$9489 ( \9866 , \9779 , \2358 );
nand \U$9490 ( \9867 , \9865 , \9866 );
xor \U$9491 ( \9868 , \9856 , \9867 );
not \U$9492 ( \9869 , \1963 );
not \U$9493 ( \9870 , \9750 );
or \U$9494 ( \9871 , \9869 , \9870 );
not \U$9495 ( \9872 , RIc226e30_17);
not \U$9496 ( \9873 , \9765 );
or \U$9497 ( \9874 , \9872 , \9873 );
not \U$9498 ( \9875 , \9768 );
nand \U$9499 ( \9876 , \9875 , \1935 );
nand \U$9500 ( \9877 , \9874 , \9876 );
nand \U$9501 ( \9878 , \9877 , \1945 );
nand \U$9502 ( \9879 , \9871 , \9878 );
xor \U$9503 ( \9880 , \9868 , \9879 );
not \U$9504 ( \9881 , \9880 );
not \U$9505 ( \9882 , \3250 );
not \U$9506 ( \9883 , RIc227010_13);
not \U$9507 ( \9884 , \8885 );
not \U$9508 ( \9885 , \9884 );
or \U$9509 ( \9886 , \9883 , \9885 );
nand \U$9510 ( \9887 , \8885 , \1296 );
nand \U$9511 ( \9888 , \9886 , \9887 );
not \U$9512 ( \9889 , \9888 );
or \U$9513 ( \9890 , \9882 , \9889 );
nand \U$9514 ( \9891 , \9733 , \1682 );
nand \U$9515 ( \9892 , \9890 , \9891 );
not \U$9516 ( \9893 , \1311 );
not \U$9517 ( \9894 , \8861 );
or \U$9518 ( \9895 , \9893 , \9894 );
not \U$9519 ( \9896 , RIc227100_11);
not \U$9520 ( \9897 , \8829 );
not \U$9521 ( \9898 , \9897 );
or \U$9522 ( \9899 , \9896 , \9898 );
not \U$9523 ( \9900 , \8829 );
not \U$9524 ( \9901 , \9900 );
nand \U$9525 ( \9902 , \9901 , \1685 );
nand \U$9526 ( \9903 , \9899 , \9902 );
buf \U$9527 ( \9904 , \1306 );
nand \U$9528 ( \9905 , \9903 , \9904 );
nand \U$9529 ( \9906 , \9895 , \9905 );
xor \U$9530 ( \9907 , \9892 , \9906 );
not \U$9531 ( \9908 , \1340 );
not \U$9532 ( \9909 , \8813 );
or \U$9533 ( \9910 , \9908 , \9909 );
not \U$9534 ( \9911 , RIc2271f0_9);
not \U$9535 ( \9912 , \8951 );
not \U$9536 ( \9913 , \9912 );
or \U$9537 ( \9914 , \9911 , \9913 );
not \U$9538 ( \9915 , \8951 );
not \U$9539 ( \9916 , \9915 );
nand \U$9540 ( \9917 , \9916 , \1351 );
nand \U$9541 ( \9918 , \9914 , \9917 );
nand \U$9542 ( \9919 , \9918 , \1363 );
nand \U$9543 ( \9920 , \9910 , \9919 );
xnor \U$9544 ( \9921 , \9907 , \9920 );
not \U$9545 ( \9922 , \9921 );
not \U$9546 ( \9923 , \9922 );
or \U$9547 ( \9924 , \9881 , \9923 );
or \U$9548 ( \9925 , \9922 , \9880 );
not \U$9549 ( \9926 , \9398 );
not \U$9550 ( \9927 , \9390 );
or \U$9551 ( \9928 , \9926 , \9927 );
not \U$9552 ( \9929 , RIc226110_45);
not \U$9553 ( \9930 , \3438 );
or \U$9554 ( \9931 , \9929 , \9930 );
nand \U$9555 ( \9932 , \1332 , \9379 );
nand \U$9556 ( \9933 , \9931 , \9932 );
buf \U$9557 ( \9934 , \9382 );
nand \U$9558 ( \9935 , \9933 , \9934 );
nand \U$9559 ( \9936 , \9928 , \9935 );
not \U$9560 ( \9937 , \9936 );
not \U$9561 ( \9938 , \3629 );
not \U$9562 ( \9939 , RIc2266b0_33);
not \U$9563 ( \9940 , \9361 );
or \U$9564 ( \9941 , \9939 , \9940 );
not \U$9565 ( \9942 , \2555 );
not \U$9566 ( \9943 , RIc2266b0_33);
nand \U$9567 ( \9944 , \9942 , \9943 );
nand \U$9568 ( \9945 , \9941 , \9944 );
not \U$9569 ( \9946 , \9945 );
or \U$9570 ( \9947 , \9938 , \9946 );
nand \U$9571 ( \9948 , \9427 , \3631 );
nand \U$9572 ( \9949 , \9947 , \9948 );
not \U$9573 ( \9950 , \9949 );
or \U$9574 ( \9951 , \9937 , \9950 );
or \U$9575 ( \9952 , \9949 , \9936 );
not \U$9576 ( \9953 , \9459 );
not \U$9577 ( \9954 , RIc225e40_51);
not \U$9578 ( \9955 , \1558 );
or \U$9579 ( \9956 , \9954 , \9955 );
nand \U$9580 ( \9957 , \3464 , \9450 );
nand \U$9581 ( \9958 , \9956 , \9957 );
not \U$9582 ( \9959 , \9958 );
or \U$9583 ( \9960 , \9953 , \9959 );
nand \U$9584 ( \9961 , \9463 , \9444 );
nand \U$9585 ( \9962 , \9960 , \9961 );
nand \U$9586 ( \9963 , \9952 , \9962 );
nand \U$9587 ( \9964 , \9951 , \9963 );
nand \U$9588 ( \9965 , \9925 , \9964 );
nand \U$9589 ( \9966 , \9924 , \9965 );
nand \U$9590 ( \9967 , \9839 , \9966 );
nand \U$9591 ( \9968 , \9838 , \9967 );
xor \U$9592 ( \9969 , \9525 , \9968 );
xor \U$9593 ( \9970 , \8894 , \9003 );
and \U$9594 ( \9971 , \9970 , \9134 );
and \U$9595 ( \9972 , \8894 , \9003 );
or \U$9596 ( \9973 , \9971 , \9972 );
not \U$9597 ( \9974 , \9783 );
not \U$9598 ( \9975 , \9834 );
or \U$9599 ( \9976 , \9974 , \9975 );
nand \U$9600 ( \9977 , \9976 , \9828 );
not \U$9601 ( \9978 , \9783 );
nand \U$9602 ( \9979 , \9978 , \9833 );
nand \U$9603 ( \9980 , \9977 , \9979 );
xor \U$9604 ( \9981 , \9973 , \9980 );
not \U$9605 ( \9982 , \9420 );
not \U$9606 ( \9983 , \9438 );
or \U$9607 ( \9984 , \9982 , \9983 );
or \U$9608 ( \9985 , \9438 , \9420 );
nand \U$9609 ( \9986 , \9985 , \9465 );
nand \U$9610 ( \9987 , \9984 , \9986 );
not \U$9611 ( \9988 , \9987 );
not \U$9612 ( \9989 , \9532 );
not \U$9613 ( \9990 , \9551 );
or \U$9614 ( \9991 , \9989 , \9990 );
not \U$9615 ( \9992 , RIc225f30_49);
not \U$9616 ( \9993 , \1558 );
or \U$9617 ( \9994 , \9992 , \9993 );
buf \U$9618 ( \9995 , \981 );
not \U$9619 ( \9996 , RIc225f30_49);
nand \U$9620 ( \9997 , \9995 , \9996 );
nand \U$9621 ( \9998 , \9994 , \9997 );
nand \U$9622 ( \9999 , \9998 , \9552 );
nand \U$9623 ( \10000 , \9991 , \9999 );
buf \U$9624 ( \10001 , \9639 );
not \U$9625 ( \10002 , \10001 );
not \U$9626 ( \10003 , \9626 );
or \U$9627 ( \10004 , \10002 , \10003 );
not \U$9628 ( \10005 , RIc226020_47);
not \U$9629 ( \10006 , \3993 );
or \U$9630 ( \10007 , \10005 , \10006 );
nand \U$9631 ( \10008 , \9540 , \9373 );
nand \U$9632 ( \10009 , \10007 , \10008 );
nand \U$9633 ( \10010 , \10009 , \9619 );
nand \U$9634 ( \10011 , \10004 , \10010 );
or \U$9635 ( \10012 , \10000 , \10011 );
not \U$9636 ( \10013 , \5509 );
not \U$9637 ( \10014 , \9602 );
or \U$9638 ( \10015 , \10013 , \10014 );
not \U$9639 ( \10016 , RIc2264d0_37);
not \U$9640 ( \10017 , \2833 );
or \U$9641 ( \10018 , \10016 , \10017 );
nand \U$9642 ( \10019 , \2832 , \5504 );
nand \U$9643 ( \10020 , \10018 , \10019 );
nand \U$9644 ( \10021 , \10020 , \5519 );
nand \U$9645 ( \10022 , \10015 , \10021 );
and \U$9646 ( \10023 , \10012 , \10022 );
and \U$9647 ( \10024 , \10000 , \10011 );
nor \U$9648 ( \10025 , \10023 , \10024 );
not \U$9649 ( \10026 , \10025 );
not \U$9650 ( \10027 , \10026 );
or \U$9651 ( \10028 , \9988 , \10027 );
not \U$9652 ( \10029 , \10025 );
not \U$9653 ( \10030 , \9987 );
not \U$9654 ( \10031 , \10030 );
or \U$9655 ( \10032 , \10029 , \10031 );
not \U$9656 ( \10033 , \9400 );
not \U$9657 ( \10034 , \9355 );
nand \U$9658 ( \10035 , \10034 , \9369 );
not \U$9659 ( \10036 , \10035 );
or \U$9660 ( \10037 , \10033 , \10036 );
nand \U$9661 ( \10038 , \9368 , \9355 );
nand \U$9662 ( \10039 , \10037 , \10038 );
nand \U$9663 ( \10040 , \10032 , \10039 );
nand \U$9664 ( \10041 , \10028 , \10040 );
xor \U$9665 ( \10042 , \9981 , \10041 );
xor \U$9666 ( \10043 , \9969 , \10042 );
not \U$9667 ( \10044 , \9523 );
not \U$9668 ( \10045 , \10044 );
not \U$9669 ( \10046 , \9135 );
not \U$9670 ( \10047 , \9337 );
or \U$9671 ( \10048 , \10046 , \10047 );
or \U$9672 ( \10049 , \9337 , \9135 );
nand \U$9673 ( \10050 , \10048 , \10049 );
not \U$9674 ( \10051 , \10050 );
or \U$9675 ( \10052 , \10045 , \10051 );
or \U$9676 ( \10053 , \10044 , \10050 );
nand \U$9677 ( \10054 , \10052 , \10053 );
not \U$9678 ( \10055 , \9473 );
not \U$9679 ( \10056 , \9402 );
or \U$9680 ( \10057 , \10055 , \10056 );
nand \U$9681 ( \10058 , \9470 , \9401 );
nand \U$9682 ( \10059 , \10057 , \10058 );
xnor \U$9683 ( \10060 , \10059 , \9521 );
not \U$9684 ( \10061 , \10060 );
not \U$9685 ( \10062 , \10061 );
xor \U$9686 ( \10063 , \9796 , \9826 );
xor \U$9687 ( \10064 , \10063 , \9809 );
xor \U$9688 ( \10065 , \10000 , \10011 );
xor \U$9689 ( \10066 , \10065 , \10022 );
xor \U$9690 ( \10067 , \10064 , \10066 );
not \U$9691 ( \10068 , RIc225af8_58);
and \U$9692 ( \10069 , RIc225a80_59, \10068 );
not \U$9693 ( \10070 , RIc225a80_59);
and \U$9694 ( \10071 , \10070 , RIc225af8_58);
or \U$9695 ( \10072 , \10069 , \10071 );
and \U$9696 ( \10073 , \10068 , RIc225b70_57);
not \U$9697 ( \10074 , RIc225b70_57);
and \U$9698 ( \10075 , \10074 , RIc225af8_58);
nor \U$9699 ( \10076 , \10073 , \10075 );
nor \U$9700 ( \10077 , \10076 , \10072 );
or \U$9701 ( \10078 , \10072 , \10077 );
nand \U$9702 ( \10079 , \10078 , RIc225b70_57);
nand \U$9703 ( \10080 , \9310 , \9314 );
and \U$9704 ( \10081 , \9238 , \10080 );
not \U$9705 ( \10082 , \9238 );
not \U$9706 ( \10083 , \10080 );
and \U$9707 ( \10084 , \10082 , \10083 );
or \U$9708 ( \10085 , \10081 , \10084 );
buf \U$9709 ( \10086 , \10085 );
and \U$9710 ( \10087 , \10086 , RIc2275b0_1);
xor \U$9711 ( \10088 , \10079 , \10087 );
not \U$9712 ( \10089 , \954 );
not \U$9713 ( \10090 , \9079 );
or \U$9714 ( \10091 , \10089 , \10090 );
not \U$9715 ( \10092 , RIc2273d0_5);
nand \U$9716 ( \10093 , \590 , \462 );
not \U$9717 ( \10094 , \10093 );
not \U$9718 ( \10095 , \505 );
nor \U$9719 ( \10096 , \10095 , \9011 );
not \U$9720 ( \10097 , \10096 );
not \U$9721 ( \10098 , \9021 );
or \U$9722 ( \10099 , \10097 , \10098 );
not \U$9723 ( \10100 , \505 );
not \U$9724 ( \10101 , \9034 );
or \U$9725 ( \10102 , \10100 , \10101 );
nand \U$9726 ( \10103 , \10102 , \9233 );
not \U$9727 ( \10104 , \10103 );
nand \U$9728 ( \10105 , \10099 , \10104 );
not \U$9729 ( \10106 , \10105 );
or \U$9730 ( \10107 , \10094 , \10106 );
or \U$9731 ( \10108 , \10105 , \10093 );
nand \U$9732 ( \10109 , \10107 , \10108 );
buf \U$9733 ( \10110 , \10109 );
not \U$9734 ( \10111 , \10110 );
not \U$9735 ( \10112 , \10111 );
or \U$9736 ( \10113 , \10092 , \10112 );
nand \U$9737 ( \10114 , \10110 , \946 );
nand \U$9738 ( \10115 , \10113 , \10114 );
nand \U$9739 ( \10116 , \10115 , \951 );
nand \U$9740 ( \10117 , \10091 , \10116 );
and \U$9741 ( \10118 , \10088 , \10117 );
and \U$9742 ( \10119 , \10079 , \10087 );
or \U$9743 ( \10120 , \10118 , \10119 );
not \U$9744 ( \10121 , \1963 );
not \U$9745 ( \10122 , RIc226e30_17);
not \U$9746 ( \10123 , \6493 );
or \U$9747 ( \10124 , \10122 , \10123 );
not \U$9748 ( \10125 , \6492 );
not \U$9749 ( \10126 , \10125 );
nand \U$9750 ( \10127 , \10126 , \1935 );
nand \U$9751 ( \10128 , \10124 , \10127 );
not \U$9752 ( \10129 , \10128 );
or \U$9753 ( \10130 , \10121 , \10129 );
not \U$9754 ( \10131 , RIc226e30_17);
not \U$9755 ( \10132 , \9859 );
or \U$9756 ( \10133 , \10131 , \10132 );
nand \U$9757 ( \10134 , \9740 , \1952 );
nand \U$9758 ( \10135 , \10133 , \10134 );
nand \U$9759 ( \10136 , \10135 , \1945 );
nand \U$9760 ( \10137 , \10130 , \10136 );
not \U$9761 ( \10138 , \10137 );
not \U$9762 ( \10139 , \2358 );
not \U$9763 ( \10140 , RIc226f20_15);
buf \U$9764 ( \10141 , \9727 );
not \U$9765 ( \10142 , \10141 );
not \U$9766 ( \10143 , \10142 );
or \U$9767 ( \10144 , \10140 , \10143 );
nand \U$9768 ( \10145 , \9731 , \2351 );
nand \U$9769 ( \10146 , \10144 , \10145 );
not \U$9770 ( \10147 , \10146 );
or \U$9771 ( \10148 , \10139 , \10147 );
not \U$9772 ( \10149 , RIc226f20_15);
not \U$9773 ( \10150 , \9884 );
or \U$9774 ( \10151 , \10149 , \10150 );
nand \U$9775 ( \10152 , \8885 , \1674 );
nand \U$9776 ( \10153 , \10151 , \10152 );
nand \U$9777 ( \10154 , \10153 , \2320 );
nand \U$9778 ( \10155 , \10148 , \10154 );
not \U$9779 ( \10156 , \10155 );
or \U$9780 ( \10157 , \10138 , \10156 );
or \U$9781 ( \10158 , \10155 , \10137 );
not \U$9782 ( \10159 , \2534 );
not \U$9783 ( \10160 , RIc226d40_19);
not \U$9784 ( \10161 , \5663 );
not \U$9785 ( \10162 , \10161 );
or \U$9786 ( \10163 , \10160 , \10162 );
not \U$9787 ( \10164 , \5664 );
nand \U$9788 ( \10165 , \10164 , \3338 );
nand \U$9789 ( \10166 , \10163 , \10165 );
not \U$9790 ( \10167 , \10166 );
or \U$9791 ( \10168 , \10159 , \10167 );
not \U$9792 ( \10169 , RIc226d40_19);
not \U$9793 ( \10170 , \6071 );
not \U$9794 ( \10171 , \10170 );
or \U$9795 ( \10172 , \10169 , \10171 );
nand \U$9796 ( \10173 , \9875 , \1941 );
nand \U$9797 ( \10174 , \10172 , \10173 );
nand \U$9798 ( \10175 , \10174 , \2518 );
nand \U$9799 ( \10176 , \10168 , \10175 );
nand \U$9800 ( \10177 , \10158 , \10176 );
nand \U$9801 ( \10178 , \10157 , \10177 );
xor \U$9802 ( \10179 , \10120 , \10178 );
not \U$9803 ( \10180 , \507 );
nand \U$9804 ( \10181 , \10180 , \580 );
not \U$9805 ( \10182 , \10181 );
and \U$9806 ( \10183 , \518 , \503 );
not \U$9807 ( \10184 , \10183 );
buf \U$9808 ( \10185 , \502 );
not \U$9809 ( \10186 , \10185 );
or \U$9810 ( \10187 , \10184 , \10186 );
buf \U$9811 ( \10188 , \568 );
and \U$9812 ( \10189 , \10188 , \503 );
not \U$9813 ( \10190 , \577 );
nor \U$9814 ( \10191 , \10189 , \10190 );
nand \U$9815 ( \10192 , \10187 , \10191 );
not \U$9816 ( \10193 , \10192 );
or \U$9817 ( \10194 , \10182 , \10193 );
or \U$9818 ( \10195 , \10192 , \10181 );
nand \U$9819 ( \10196 , \10194 , \10195 );
buf \U$9820 ( \10197 , \10196 );
not \U$9821 ( \10198 , \10197 );
buf \U$9822 ( \10199 , \10198 );
not \U$9823 ( \10200 , \10199 );
nand \U$9824 ( \10201 , \10200 , RIc2275b0_1);
not \U$9825 ( \10202 , \10201 );
not \U$9826 ( \10203 , \1930 );
not \U$9827 ( \10204 , \9677 );
or \U$9828 ( \10205 , \10203 , \10204 );
not \U$9829 ( \10206 , RIc226b60_23);
not \U$9830 ( \10207 , \4417 );
or \U$9831 ( \10208 , \10206 , \10207 );
not \U$9832 ( \10209 , \4414 );
not \U$9833 ( \10210 , RIc226b60_23);
nand \U$9834 ( \10211 , \10209 , \10210 );
nand \U$9835 ( \10212 , \10208 , \10211 );
not \U$9836 ( \10213 , \1914 );
not \U$9837 ( \10214 , \10213 );
nand \U$9838 ( \10215 , \10212 , \10214 );
nand \U$9839 ( \10216 , \10205 , \10215 );
xor \U$9840 ( \10217 , \10202 , \10216 );
not \U$9841 ( \10218 , \2367 );
not \U$9842 ( \10219 , RIc226c50_21);
not \U$9843 ( \10220 , \4406 );
not \U$9844 ( \10221 , \10220 );
or \U$9845 ( \10222 , \10219 , \10221 );
nand \U$9846 ( \10223 , \4406 , \2370 );
nand \U$9847 ( \10224 , \10222 , \10223 );
not \U$9848 ( \10225 , \10224 );
or \U$9849 ( \10226 , \10218 , \10225 );
not \U$9850 ( \10227 , RIc226c50_21);
not \U$9851 ( \10228 , \9850 );
or \U$9852 ( \10229 , \10227 , \10228 );
not \U$9853 ( \10230 , \5215 );
not \U$9854 ( \10231 , \10230 );
nand \U$9855 ( \10232 , \10231 , \2370 );
nand \U$9856 ( \10233 , \10229 , \10232 );
nand \U$9857 ( \10234 , \10233 , \2392 );
nand \U$9858 ( \10235 , \10226 , \10234 );
and \U$9859 ( \10236 , \10217 , \10235 );
and \U$9860 ( \10237 , \10202 , \10216 );
or \U$9861 ( \10238 , \10236 , \10237 );
and \U$9862 ( \10239 , \10179 , \10238 );
and \U$9863 ( \10240 , \10120 , \10178 );
or \U$9864 ( \10241 , \10239 , \10240 );
xor \U$9865 ( \10242 , \10067 , \10241 );
not \U$9866 ( \10243 , \10242 );
or \U$9867 ( \10244 , \10062 , \10243 );
not \U$9868 ( \10245 , \10060 );
not \U$9869 ( \10246 , \10242 );
not \U$9870 ( \10247 , \10246 );
or \U$9871 ( \10248 , \10245 , \10247 );
not \U$9872 ( \10249 , \9593 );
not \U$9873 ( \10250 , \9613 );
or \U$9874 ( \10251 , \10249 , \10250 );
or \U$9875 ( \10252 , \9613 , \9593 );
nand \U$9876 ( \10253 , \10251 , \10252 );
xor \U$9877 ( \10254 , \10253 , \9643 );
not \U$9878 ( \10255 , \10254 );
xor \U$9879 ( \10256 , \9679 , \9707 );
xnor \U$9880 ( \10257 , \10256 , \9666 );
nand \U$9881 ( \10258 , \10255 , \10257 );
not \U$9882 ( \10259 , \1082 );
not \U$9883 ( \10260 , \9280 );
or \U$9884 ( \10261 , \10259 , \10260 );
not \U$9885 ( \10262 , RIc2274c0_3);
not \U$9886 ( \10263 , \9296 );
not \U$9887 ( \10264 , \10263 );
or \U$9888 ( \10265 , \10262 , \10264 );
not \U$9889 ( \10266 , \10263 );
nand \U$9890 ( \10267 , \10266 , \1027 );
nand \U$9891 ( \10268 , \10265 , \10267 );
nand \U$9892 ( \10269 , \10268 , \1040 );
nand \U$9893 ( \10270 , \10261 , \10269 );
xor \U$9894 ( \10271 , \10201 , \10270 );
not \U$9895 ( \10272 , \1930 );
not \U$9896 ( \10273 , \10212 );
or \U$9897 ( \10274 , \10272 , \10273 );
and \U$9898 ( \10275 , RIc226b60_23, \4406 );
not \U$9899 ( \10276 , RIc226b60_23);
not \U$9900 ( \10277 , \4405 );
and \U$9901 ( \10278 , \10276 , \10277 );
nor \U$9902 ( \10279 , \10275 , \10278 );
nand \U$9903 ( \10280 , \10279 , \1915 );
nand \U$9904 ( \10281 , \10274 , \10280 );
and \U$9905 ( \10282 , \10271 , \10281 );
and \U$9906 ( \10283 , \10201 , \10270 );
or \U$9907 ( \10284 , \10282 , \10283 );
not \U$9908 ( \10285 , \1682 );
not \U$9909 ( \10286 , RIc227010_13);
not \U$9910 ( \10287 , \9900 );
or \U$9911 ( \10288 , \10286 , \10287 );
not \U$9912 ( \10289 , \9897 );
nand \U$9913 ( \10290 , \10289 , \1296 );
nand \U$9914 ( \10291 , \10288 , \10290 );
not \U$9915 ( \10292 , \10291 );
or \U$9916 ( \10293 , \10285 , \10292 );
not \U$9917 ( \10294 , RIc227010_13);
not \U$9918 ( \10295 , \8806 );
not \U$9919 ( \10296 , \10295 );
or \U$9920 ( \10297 , \10294 , \10296 );
nand \U$9921 ( \10298 , \8806 , \1758 );
nand \U$9922 ( \10299 , \10297 , \10298 );
nand \U$9923 ( \10300 , \10299 , \3250 );
nand \U$9924 ( \10301 , \10293 , \10300 );
not \U$9925 ( \10302 , \10301 );
not \U$9926 ( \10303 , \1963 );
not \U$9927 ( \10304 , \10135 );
or \U$9928 ( \10305 , \10303 , \10304 );
not \U$9929 ( \10306 , RIc226e30_17);
not \U$9930 ( \10307 , \9731 );
not \U$9931 ( \10308 , \10307 );
or \U$9932 ( \10309 , \10306 , \10308 );
buf \U$9933 ( \10310 , \9731 );
nand \U$9934 ( \10311 , \10310 , \1952 );
nand \U$9935 ( \10312 , \10309 , \10311 );
nand \U$9936 ( \10313 , \10312 , \1945 );
nand \U$9937 ( \10314 , \10305 , \10313 );
not \U$9938 ( \10315 , \10314 );
or \U$9939 ( \10316 , \10302 , \10315 );
or \U$9940 ( \10317 , \10314 , \10301 );
not \U$9941 ( \10318 , \2358 );
not \U$9942 ( \10319 , \10153 );
or \U$9943 ( \10320 , \10318 , \10319 );
not \U$9944 ( \10321 , RIc226f20_15);
not \U$9945 ( \10322 , \8856 );
not \U$9946 ( \10323 , \10322 );
or \U$9947 ( \10324 , \10321 , \10323 );
nand \U$9948 ( \10325 , \8856 , \2301 );
nand \U$9949 ( \10326 , \10324 , \10325 );
nand \U$9950 ( \10327 , \10326 , \2320 );
nand \U$9951 ( \10328 , \10320 , \10327 );
nand \U$9952 ( \10329 , \10317 , \10328 );
nand \U$9953 ( \10330 , \10316 , \10329 );
xor \U$9954 ( \10331 , \10284 , \10330 );
not \U$9955 ( \10332 , RIc225a08_60);
and \U$9956 ( \10333 , RIc225a80_59, \10332 );
not \U$9957 ( \10334 , RIc225a80_59);
and \U$9958 ( \10335 , \10334 , RIc225a08_60);
nor \U$9959 ( \10336 , \10333 , \10335 );
or \U$9960 ( \10337 , \10332 , RIc225990_61);
not \U$9961 ( \10338 , RIc225990_61);
or \U$9962 ( \10339 , \10338 , RIc225a08_60);
nand \U$9963 ( \10340 , \10337 , \10339 );
nor \U$9964 ( \10341 , \10336 , \10340 );
buf \U$9965 ( \10342 , \10340 );
or \U$9966 ( \10343 , \10341 , \10342 );
nand \U$9967 ( \10344 , \10343 , RIc225a80_59);
not \U$9968 ( \10345 , \518 );
not \U$9969 ( \10346 , \10185 );
or \U$9970 ( \10347 , \10345 , \10346 );
not \U$9971 ( \10348 , \10188 );
nand \U$9972 ( \10349 , \10347 , \10348 );
and \U$9973 ( \10350 , \503 , \577 );
and \U$9974 ( \10351 , \10349 , \10350 );
not \U$9975 ( \10352 , \10349 );
not \U$9976 ( \10353 , \10350 );
and \U$9977 ( \10354 , \10352 , \10353 );
nor \U$9978 ( \10355 , \10351 , \10354 );
buf \U$9979 ( \10356 , \10355 );
and \U$9980 ( \10357 , RIc2275b0_1, \10356 );
xor \U$9981 ( \10358 , \10344 , \10357 );
not \U$9982 ( \10359 , \1579 );
not \U$9983 ( \10360 , \10086 );
and \U$9984 ( \10361 , RIc2275b0_1, \10360 );
not \U$9985 ( \10362 , RIc2275b0_1);
and \U$9986 ( \10363 , \10362 , \10086 );
or \U$9987 ( \10364 , \10361 , \10363 );
not \U$9988 ( \10365 , \10364 );
or \U$9989 ( \10366 , \10359 , \10365 );
and \U$9990 ( \10367 , RIc2275b0_1, \10198 );
not \U$9991 ( \10368 , RIc2275b0_1);
not \U$9992 ( \10369 , \10196 );
not \U$9993 ( \10370 , \10369 );
and \U$9994 ( \10371 , \10368 , \10370 );
or \U$9995 ( \10372 , \10367 , \10371 );
nand \U$9996 ( \10373 , \10372 , \854 );
nand \U$9997 ( \10374 , \10366 , \10373 );
and \U$9998 ( \10375 , \10358 , \10374 );
and \U$9999 ( \10376 , \10344 , \10357 );
or \U$10000 ( \10377 , \10375 , \10376 );
not \U$10001 ( \10378 , \2534 );
not \U$10002 ( \10379 , \10174 );
or \U$10003 ( \10380 , \10378 , \10379 );
not \U$10004 ( \10381 , RIc226d40_19);
not \U$10005 ( \10382 , \9775 );
or \U$10006 ( \10383 , \10381 , \10382 );
nand \U$10007 ( \10384 , \6492 , \3338 );
nand \U$10008 ( \10385 , \10383 , \10384 );
nand \U$10009 ( \10386 , \10385 , \2518 );
nand \U$10010 ( \10387 , \10380 , \10386 );
xor \U$10011 ( \10388 , \10377 , \10387 );
not \U$10012 ( \10389 , \2367 );
not \U$10013 ( \10390 , \10233 );
or \U$10014 ( \10391 , \10389 , \10390 );
and \U$10015 ( \10392 , \5663 , \3204 );
not \U$10016 ( \10393 , \5663 );
and \U$10017 ( \10394 , \10393 , RIc226c50_21);
or \U$10018 ( \10395 , \10392 , \10394 );
nand \U$10019 ( \10396 , \10395 , \2392 );
nand \U$10020 ( \10397 , \10391 , \10396 );
and \U$10021 ( \10398 , \10388 , \10397 );
and \U$10022 ( \10399 , \10377 , \10387 );
or \U$10023 ( \10400 , \10398 , \10399 );
and \U$10024 ( \10401 , \10331 , \10400 );
and \U$10025 ( \10402 , \10284 , \10330 );
or \U$10026 ( \10403 , \10401 , \10402 );
and \U$10027 ( \10404 , \10258 , \10403 );
nor \U$10028 ( \10405 , \10255 , \10257 );
nor \U$10029 ( \10406 , \10404 , \10405 );
not \U$10030 ( \10407 , \10406 );
nand \U$10031 ( \10408 , \10248 , \10407 );
nand \U$10032 ( \10409 , \10244 , \10408 );
xor \U$10033 ( \10410 , \10054 , \10409 );
xor \U$10034 ( \10411 , \10064 , \10066 );
and \U$10035 ( \10412 , \10411 , \10241 );
and \U$10036 ( \10413 , \10064 , \10066 );
or \U$10037 ( \10414 , \10412 , \10413 );
not \U$10038 ( \10415 , \10039 );
not \U$10039 ( \10416 , \10030 );
or \U$10040 ( \10417 , \10415 , \10416 );
not \U$10041 ( \10418 , \10039 );
nand \U$10042 ( \10419 , \10418 , \9987 );
nand \U$10043 ( \10420 , \10417 , \10419 );
xor \U$10044 ( \10421 , \10026 , \10420 );
xor \U$10045 ( \10422 , \10414 , \10421 );
not \U$10046 ( \10423 , \9398 );
not \U$10047 ( \10424 , RIc226110_45);
not \U$10048 ( \10425 , \1222 );
or \U$10049 ( \10426 , \10424 , \10425 );
not \U$10050 ( \10427 , \1370 );
not \U$10051 ( \10428 , \10427 );
not \U$10052 ( \10429 , RIc226110_45);
nand \U$10053 ( \10430 , \10428 , \10429 );
nand \U$10054 ( \10431 , \10426 , \10430 );
not \U$10055 ( \10432 , \10431 );
or \U$10056 ( \10433 , \10423 , \10432 );
nand \U$10057 ( \10434 , \9397 , \9934 );
nand \U$10058 ( \10435 , \10433 , \10434 );
not \U$10059 ( \10436 , \3629 );
not \U$10060 ( \10437 , \9436 );
or \U$10061 ( \10438 , \10436 , \10437 );
and \U$10062 ( \10439 , \1988 , \2692 );
not \U$10063 ( \10440 , \1988 );
and \U$10064 ( \10441 , \10440 , RIc2266b0_33);
or \U$10065 ( \10442 , \10439 , \10441 );
nand \U$10066 ( \10443 , \10442 , \3631 );
nand \U$10067 ( \10444 , \10438 , \10443 );
not \U$10068 ( \10445 , \9533 );
not \U$10069 ( \10446 , \10445 );
not \U$10070 ( \10447 , \9998 );
or \U$10071 ( \10448 , \10446 , \10447 );
not \U$10072 ( \10449 , RIc225f30_49);
not \U$10073 ( \10450 , \840 );
not \U$10074 ( \10451 , \10450 );
or \U$10075 ( \10452 , \10449 , \10451 );
nand \U$10076 ( \10453 , \840 , \9549 );
nand \U$10077 ( \10454 , \10452 , \10453 );
nand \U$10078 ( \10455 , \10454 , \9552 );
nand \U$10079 ( \10456 , \10448 , \10455 );
xor \U$10080 ( \10457 , \10444 , \10456 );
xor \U$10081 ( \10458 , \10435 , \10457 );
not \U$10082 ( \10459 , \10458 );
not \U$10083 ( \10460 , \10459 );
not \U$10084 ( \10461 , \2697 );
not \U$10085 ( \10462 , \9366 );
or \U$10086 ( \10463 , \10461 , \10462 );
not \U$10087 ( \10464 , RIc2267a0_31);
not \U$10088 ( \10465 , \9422 );
or \U$10089 ( \10466 , \10464 , \10465 );
nand \U$10090 ( \10467 , \2590 , \2072 );
nand \U$10091 ( \10468 , \10466 , \10467 );
nand \U$10092 ( \10469 , \10468 , \2711 );
nand \U$10093 ( \10470 , \10463 , \10469 );
not \U$10094 ( \10471 , \2784 );
not \U$10095 ( \10472 , \9353 );
or \U$10096 ( \10473 , \10471 , \10472 );
not \U$10097 ( \10474 , RIc226890_29);
not \U$10098 ( \10475 , \3035 );
or \U$10099 ( \10476 , \10474 , \10475 );
not \U$10100 ( \10477 , RIc226890_29);
nand \U$10101 ( \10478 , \10477 , \2475 );
nand \U$10102 ( \10479 , \10476 , \10478 );
nand \U$10103 ( \10480 , \10479 , \9142 );
nand \U$10104 ( \10481 , \10473 , \10480 );
xor \U$10105 ( \10482 , \10470 , \10481 );
not \U$10106 ( \10483 , \9110 );
not \U$10107 ( \10484 , \9127 );
or \U$10108 ( \10485 , \10483 , \10484 );
not \U$10109 ( \10486 , RIc226200_43);
not \U$10110 ( \10487 , \4590 );
or \U$10111 ( \10488 , \10486 , \10487 );
nand \U$10112 ( \10489 , \3579 , \9106 );
nand \U$10113 ( \10490 , \10488 , \10489 );
nand \U$10114 ( \10491 , \10490 , \9129 );
nand \U$10115 ( \10492 , \10485 , \10491 );
xnor \U$10116 ( \10493 , \10482 , \10492 );
not \U$10117 ( \10494 , \2367 );
not \U$10118 ( \10495 , RIc226c50_21);
not \U$10119 ( \10496 , \2980 );
not \U$10120 ( \10497 , \10496 );
or \U$10121 ( \10498 , \10495 , \10497 );
nand \U$10122 ( \10499 , \2980 , \2370 );
nand \U$10123 ( \10500 , \10498 , \10499 );
not \U$10124 ( \10501 , \10500 );
or \U$10125 ( \10502 , \10494 , \10501 );
not \U$10126 ( \10503 , RIc226c50_21);
not \U$10127 ( \10504 , \4049 );
or \U$10128 ( \10505 , \10503 , \10504 );
nand \U$10129 ( \10506 , \3640 , \2383 );
nand \U$10130 ( \10507 , \10505 , \10506 );
nand \U$10131 ( \10508 , \10507 , \2392 );
nand \U$10132 ( \10509 , \10502 , \10508 );
not \U$10133 ( \10510 , \10509 );
not \U$10134 ( \10511 , \10510 );
not \U$10135 ( \10512 , \9459 );
not \U$10136 ( \10513 , \9452 );
or \U$10137 ( \10514 , \10512 , \10513 );
not \U$10138 ( \10515 , RIc225e40_51);
not \U$10139 ( \10516 , \3071 );
or \U$10140 ( \10517 , \10515 , \10516 );
nand \U$10141 ( \10518 , \1072 , \9450 );
nand \U$10142 ( \10519 , \10517 , \10518 );
nand \U$10143 ( \10520 , \10519 , \9445 );
nand \U$10144 ( \10521 , \10514 , \10520 );
not \U$10145 ( \10522 , \10521 );
or \U$10146 ( \10523 , \10511 , \10522 );
or \U$10147 ( \10524 , \10510 , \10521 );
nand \U$10148 ( \10525 , \10523 , \10524 );
not \U$10149 ( \10526 , \9517 );
not \U$10150 ( \10527 , \5643 );
and \U$10151 ( \10528 , \10526 , \10527 );
not \U$10152 ( \10529 , RIc226b60_23);
not \U$10153 ( \10530 , \9651 );
or \U$10154 ( \10531 , \10529 , \10530 );
not \U$10155 ( \10532 , \2103 );
not \U$10156 ( \10533 , \10532 );
nand \U$10157 ( \10534 , \10533 , \1911 );
nand \U$10158 ( \10535 , \10531 , \10534 );
and \U$10159 ( \10536 , \10535 , \1930 );
nor \U$10160 ( \10537 , \10528 , \10536 );
not \U$10161 ( \10538 , \10537 );
and \U$10162 ( \10539 , \10525 , \10538 );
not \U$10163 ( \10540 , \10525 );
and \U$10164 ( \10541 , \10540 , \10537 );
nor \U$10165 ( \10542 , \10539 , \10541 );
xnor \U$10166 ( \10543 , \10493 , \10542 );
not \U$10167 ( \10544 , \10543 );
or \U$10168 ( \10545 , \10460 , \10544 );
or \U$10169 ( \10546 , \10543 , \10459 );
nand \U$10170 ( \10547 , \10545 , \10546 );
xor \U$10171 ( \10548 , \10422 , \10547 );
and \U$10172 ( \10549 , \10410 , \10548 );
and \U$10173 ( \10550 , \10054 , \10409 );
or \U$10174 ( \10551 , \10549 , \10550 );
xor \U$10175 ( \10552 , \10043 , \10551 );
not \U$10176 ( \10553 , \10414 );
not \U$10177 ( \10554 , \10421 );
nand \U$10178 ( \10555 , \10553 , \10554 );
and \U$10179 ( \10556 , \10555 , \10547 );
and \U$10180 ( \10557 , \10414 , \10421 );
nor \U$10181 ( \10558 , \10556 , \10557 );
not \U$10182 ( \10559 , \10492 );
not \U$10183 ( \10560 , \10481 );
or \U$10184 ( \10561 , \10559 , \10560 );
or \U$10185 ( \10562 , \10481 , \10492 );
nand \U$10186 ( \10563 , \10562 , \10470 );
nand \U$10187 ( \10564 , \10561 , \10563 );
xor \U$10188 ( \10565 , \8931 , \8983 );
and \U$10189 ( \10566 , \10565 , \9002 );
and \U$10190 ( \10567 , \8931 , \8983 );
or \U$10191 ( \10568 , \10566 , \10567 );
xor \U$10192 ( \10569 , \10564 , \10568 );
nand \U$10193 ( \10570 , \10537 , \10510 );
and \U$10194 ( \10571 , \10570 , \10521 );
nor \U$10195 ( \10572 , \10537 , \10510 );
nor \U$10196 ( \10573 , \10571 , \10572 );
xor \U$10197 ( \10574 , \10569 , \10573 );
not \U$10198 ( \10575 , RIc2275b0_1);
nor \U$10199 ( \10576 , \10575 , \9251 );
not \U$10200 ( \10577 , \1945 );
not \U$10201 ( \10578 , \9759 );
or \U$10202 ( \10579 , \10577 , \10578 );
not \U$10203 ( \10580 , RIc226e30_17);
not \U$10204 ( \10581 , \10277 );
or \U$10205 ( \10582 , \10580 , \10581 );
nand \U$10206 ( \10583 , \4405 , \1935 );
nand \U$10207 ( \10584 , \10582 , \10583 );
nand \U$10208 ( \10585 , \10584 , \1963 );
nand \U$10209 ( \10586 , \10579 , \10585 );
xor \U$10210 ( \10587 , \10576 , \10586 );
not \U$10211 ( \10588 , \2534 );
not \U$10212 ( \10589 , RIc226d40_19);
not \U$10213 ( \10590 , \9674 );
or \U$10214 ( \10591 , \10589 , \10590 );
nand \U$10215 ( \10592 , \3640 , \2523 );
nand \U$10216 ( \10593 , \10591 , \10592 );
not \U$10217 ( \10594 , \10593 );
or \U$10218 ( \10595 , \10588 , \10594 );
not \U$10219 ( \10596 , RIc226d40_19);
not \U$10220 ( \10597 , \4122 );
or \U$10221 ( \10598 , \10596 , \10597 );
not \U$10222 ( \10599 , \4414 );
nand \U$10223 ( \10600 , \10599 , \2523 );
nand \U$10224 ( \10601 , \10598 , \10600 );
nand \U$10225 ( \10602 , \10601 , \2518 );
nand \U$10226 ( \10603 , \10595 , \10602 );
xor \U$10227 ( \10604 , \10587 , \10603 );
not \U$10228 ( \10605 , \9904 );
not \U$10229 ( \10606 , \8891 );
or \U$10230 ( \10607 , \10605 , \10606 );
not \U$10231 ( \10608 , RIc227100_11);
not \U$10232 ( \10609 , \9731 );
not \U$10233 ( \10610 , \10609 );
or \U$10234 ( \10611 , \10608 , \10610 );
not \U$10235 ( \10612 , \10307 );
nand \U$10236 ( \10613 , \10612 , \3351 );
nand \U$10237 ( \10614 , \10611 , \10613 );
nand \U$10238 ( \10615 , \10614 , \1311 );
nand \U$10239 ( \10616 , \10607 , \10615 );
not \U$10240 ( \10617 , \2320 );
not \U$10241 ( \10618 , \9772 );
or \U$10242 ( \10619 , \10617 , \10618 );
not \U$10243 ( \10620 , \5663 );
not \U$10244 ( \10621 , \2301 );
and \U$10245 ( \10622 , \10620 , \10621 );
and \U$10246 ( \10623 , \5663 , \2301 );
nor \U$10247 ( \10624 , \10622 , \10623 );
not \U$10248 ( \10625 , \10624 );
nand \U$10249 ( \10626 , \10625 , \2358 );
nand \U$10250 ( \10627 , \10619 , \10626 );
xor \U$10251 ( \10628 , \10616 , \10627 );
not \U$10252 ( \10629 , \1682 );
not \U$10253 ( \10630 , RIc227010_13);
not \U$10254 ( \10631 , \9775 );
or \U$10255 ( \10632 , \10630 , \10631 );
nand \U$10256 ( \10633 , \6492 , \1296 );
nand \U$10257 ( \10634 , \10632 , \10633 );
not \U$10258 ( \10635 , \10634 );
or \U$10259 ( \10636 , \10629 , \10635 );
not \U$10260 ( \10637 , \9742 );
nand \U$10261 ( \10638 , \10637 , \3250 );
nand \U$10262 ( \10639 , \10636 , \10638 );
xor \U$10263 ( \10640 , \10628 , \10639 );
xor \U$10264 ( \10641 , \10604 , \10640 );
not \U$10265 ( \10642 , RIc2274c0_3);
not \U$10266 ( \10643 , \9045 );
not \U$10267 ( \10644 , \10643 );
not \U$10268 ( \10645 , \10644 );
not \U$10269 ( \10646 , \10645 );
or \U$10270 ( \10647 , \10642 , \10646 );
nand \U$10271 ( \10648 , \9225 , \2896 );
nand \U$10272 ( \10649 , \10647 , \10648 );
and \U$10273 ( \10650 , \10649 , \1082 );
not \U$10274 ( \10651 , RIc2274c0_3);
not \U$10275 ( \10652 , \9071 );
not \U$10276 ( \10653 , \10652 );
not \U$10277 ( \10654 , \10653 );
not \U$10278 ( \10655 , \10654 );
or \U$10279 ( \10656 , \10651 , \10655 );
nand \U$10280 ( \10657 , \9072 , \2896 );
nand \U$10281 ( \10658 , \10656 , \10657 );
and \U$10282 ( \10659 , \10658 , \1040 );
nor \U$10283 ( \10660 , \10650 , \10659 );
not \U$10284 ( \10661 , \2138 );
not \U$10285 ( \10662 , \9094 );
or \U$10286 ( \10663 , \10661 , \10662 );
and \U$10287 ( \10664 , RIc226980_27, \2670 );
not \U$10288 ( \10665 , RIc226980_27);
and \U$10289 ( \10666 , \10665 , \2720 );
or \U$10290 ( \10667 , \10664 , \10666 );
nand \U$10291 ( \10668 , \10667 , \2154 );
nand \U$10292 ( \10669 , \10663 , \10668 );
xor \U$10293 ( \10670 , \10660 , \10669 );
not \U$10294 ( \10671 , \9690 );
not \U$10295 ( \10672 , \9824 );
or \U$10296 ( \10673 , \10671 , \10672 );
not \U$10297 ( \10674 , RIc2262f0_41);
not \U$10298 ( \10675 , \3783 );
or \U$10299 ( \10676 , \10674 , \10675 );
not \U$10300 ( \10677 , \1485 );
not \U$10301 ( \10678 , \10677 );
not \U$10302 ( \10679 , RIc2262f0_41);
nand \U$10303 ( \10680 , \10678 , \10679 );
nand \U$10304 ( \10681 , \10676 , \10680 );
nand \U$10305 ( \10682 , \10681 , \9705 );
nand \U$10306 ( \10683 , \10673 , \10682 );
and \U$10307 ( \10684 , \10670 , \10683 );
and \U$10308 ( \10685 , \10660 , \10669 );
or \U$10309 ( \10686 , \10684 , \10685 );
xor \U$10310 ( \10687 , \10641 , \10686 );
xor \U$10311 ( \10688 , \10574 , \10687 );
not \U$10312 ( \10689 , \10493 );
not \U$10313 ( \10690 , \10689 );
not \U$10314 ( \10691 , \10542 );
or \U$10315 ( \10692 , \10690 , \10691 );
not \U$10316 ( \10693 , \10542 );
nand \U$10317 ( \10694 , \10693 , \10493 );
nand \U$10318 ( \10695 , \10694 , \10458 );
nand \U$10319 ( \10696 , \10692 , \10695 );
xor \U$10320 ( \10697 , \10688 , \10696 );
and \U$10321 ( \10698 , \10558 , \10697 );
not \U$10322 ( \10699 , \10558 );
not \U$10323 ( \10700 , \10697 );
and \U$10324 ( \10701 , \10699 , \10700 );
nor \U$10325 ( \10702 , \10698 , \10701 );
not \U$10326 ( \10703 , \10435 );
not \U$10327 ( \10704 , \10456 );
or \U$10328 ( \10705 , \10703 , \10704 );
or \U$10329 ( \10706 , \10456 , \10435 );
nand \U$10330 ( \10707 , \10706 , \10444 );
nand \U$10331 ( \10708 , \10705 , \10707 );
not \U$10332 ( \10709 , \10708 );
not \U$10333 ( \10710 , \9639 );
not \U$10334 ( \10711 , \10009 );
or \U$10335 ( \10712 , \10710 , \10711 );
not \U$10336 ( \10713 , RIc226020_47);
not \U$10337 ( \10714 , \2118 );
or \U$10338 ( \10715 , \10713 , \10714 );
nand \U$10339 ( \10716 , \1020 , \9624 );
nand \U$10340 ( \10717 , \10715 , \10716 );
nand \U$10341 ( \10718 , \10717 , \9619 );
nand \U$10342 ( \10719 , \10712 , \10718 );
not \U$10343 ( \10720 , \10719 );
not \U$10344 ( \10721 , \4381 );
not \U$10345 ( \10722 , \9418 );
or \U$10346 ( \10723 , \10721 , \10722 );
and \U$10347 ( \10724 , \2225 , \4376 );
not \U$10348 ( \10725 , \2225 );
and \U$10349 ( \10726 , \10725 , RIc2265c0_35);
or \U$10350 ( \10727 , \10724 , \10726 );
nand \U$10351 ( \10728 , \10727 , \4383 );
nand \U$10352 ( \10729 , \10723 , \10728 );
not \U$10353 ( \10730 , \10729 );
or \U$10354 ( \10731 , \10720 , \10730 );
or \U$10355 ( \10732 , \10719 , \10729 );
not \U$10356 ( \10733 , \5509 );
not \U$10357 ( \10734 , \10020 );
or \U$10358 ( \10735 , \10733 , \10734 );
and \U$10359 ( \10736 , \2421 , \4371 );
not \U$10360 ( \10737 , \2421 );
and \U$10361 ( \10738 , \10737 , RIc2264d0_37);
or \U$10362 ( \10739 , \10736 , \10738 );
nand \U$10363 ( \10740 , \10739 , \5519 );
nand \U$10364 ( \10741 , \10735 , \10740 );
nand \U$10365 ( \10742 , \10732 , \10741 );
nand \U$10366 ( \10743 , \10731 , \10742 );
not \U$10367 ( \10744 , \10743 );
not \U$10368 ( \10745 , \951 );
not \U$10369 ( \10746 , \8915 );
or \U$10370 ( \10747 , \10745 , \10746 );
xor \U$10371 ( \10748 , \8966 , \8967 );
and \U$10372 ( \10749 , \10748 , \946 );
not \U$10373 ( \10750 , \10748 );
and \U$10374 ( \10751 , \10750 , RIc2273d0_5);
or \U$10375 ( \10752 , \10749 , \10751 );
nand \U$10376 ( \10753 , \10752 , \954 );
nand \U$10377 ( \10754 , \10747 , \10753 );
not \U$10378 ( \10755 , \1339 );
and \U$10379 ( \10756 , \8856 , \1351 );
not \U$10380 ( \10757 , \8856 );
and \U$10381 ( \10758 , \10757 , RIc2271f0_9);
or \U$10382 ( \10759 , \10756 , \10758 );
not \U$10383 ( \10760 , \10759 );
or \U$10384 ( \10761 , \10755 , \10760 );
nand \U$10385 ( \10762 , \8835 , \1363 );
nand \U$10386 ( \10763 , \10761 , \10762 );
xor \U$10387 ( \10764 , \10754 , \10763 );
not \U$10388 ( \10765 , \1118 );
not \U$10389 ( \10766 , \8957 );
or \U$10390 ( \10767 , \10765 , \10766 );
and \U$10391 ( \10768 , \8807 , RIc2272e0_7);
not \U$10392 ( \10769 , \8807 );
and \U$10393 ( \10770 , \10769 , \3027 );
or \U$10394 ( \10771 , \10768 , \10770 );
nand \U$10395 ( \10772 , \10771 , \1120 );
nand \U$10396 ( \10773 , \10767 , \10772 );
xor \U$10397 ( \10774 , \10764 , \10773 );
not \U$10398 ( \10775 , \10774 );
not \U$10399 ( \10776 , \10775 );
and \U$10400 ( \10777 , \10744 , \10776 );
and \U$10401 ( \10778 , \10743 , \10775 );
nor \U$10402 ( \10779 , \10777 , \10778 );
not \U$10403 ( \10780 , \10779 );
or \U$10404 ( \10781 , \10709 , \10780 );
not \U$10405 ( \10782 , \10779 );
not \U$10406 ( \10783 , \10708 );
nand \U$10407 ( \10784 , \10782 , \10783 );
nand \U$10408 ( \10785 , \10781 , \10784 );
xor \U$10409 ( \10786 , \10660 , \10669 );
xor \U$10410 ( \10787 , \10786 , \10683 );
not \U$10411 ( \10788 , \10787 );
xor \U$10412 ( \10789 , \10741 , \10729 );
xnor \U$10413 ( \10790 , \10789 , \10719 );
not \U$10414 ( \10791 , \10790 );
not \U$10415 ( \10792 , \10791 );
or \U$10416 ( \10793 , \10788 , \10792 );
not \U$10417 ( \10794 , \10787 );
not \U$10418 ( \10795 , \10794 );
not \U$10419 ( \10796 , \10790 );
or \U$10420 ( \10797 , \10795 , \10796 );
and \U$10421 ( \10798 , \9320 , RIc2275b0_1);
not \U$10422 ( \10799 , \1579 );
not \U$10423 ( \10800 , \9274 );
and \U$10424 ( \10801 , RIc2275b0_1, \10800 );
not \U$10425 ( \10802 , RIc2275b0_1);
and \U$10426 ( \10803 , \10802 , \9275 );
or \U$10427 ( \10804 , \10801 , \10803 );
not \U$10428 ( \10805 , \10804 );
or \U$10429 ( \10806 , \10799 , \10805 );
nand \U$10430 ( \10807 , \9304 , \854 );
nand \U$10431 ( \10808 , \10806 , \10807 );
xor \U$10432 ( \10809 , \10798 , \10808 );
not \U$10433 ( \10810 , \1040 );
not \U$10434 ( \10811 , \9258 );
or \U$10435 ( \10812 , \10810 , \10811 );
not \U$10436 ( \10813 , RIc2274c0_3);
not \U$10437 ( \10814 , \10110 );
not \U$10438 ( \10815 , \10814 );
or \U$10439 ( \10816 , \10813 , \10815 );
nand \U$10440 ( \10817 , \10110 , \1078 );
nand \U$10441 ( \10818 , \10816 , \10817 );
nand \U$10442 ( \10819 , \10818 , \1082 );
nand \U$10443 ( \10820 , \10812 , \10819 );
and \U$10444 ( \10821 , \10809 , \10820 );
and \U$10445 ( \10822 , \10798 , \10808 );
or \U$10446 ( \10823 , \10821 , \10822 );
not \U$10447 ( \10824 , \1963 );
not \U$10448 ( \10825 , \9877 );
or \U$10449 ( \10826 , \10824 , \10825 );
nand \U$10450 ( \10827 , \10128 , \1945 );
nand \U$10451 ( \10828 , \10826 , \10827 );
not \U$10452 ( \10829 , \10828 );
not \U$10453 ( \10830 , \2367 );
not \U$10454 ( \10831 , RIc226c50_21);
not \U$10455 ( \10832 , \4414 );
or \U$10456 ( \10833 , \10831 , \10832 );
not \U$10457 ( \10834 , RIc226c50_21);
nand \U$10458 ( \10835 , \4418 , \10834 );
nand \U$10459 ( \10836 , \10833 , \10835 );
not \U$10460 ( \10837 , \10836 );
or \U$10461 ( \10838 , \10830 , \10837 );
nand \U$10462 ( \10839 , \10224 , \2392 );
nand \U$10463 ( \10840 , \10838 , \10839 );
not \U$10464 ( \10841 , \10840 );
or \U$10465 ( \10842 , \10829 , \10841 );
or \U$10466 ( \10843 , \10840 , \10828 );
not \U$10467 ( \10844 , \2518 );
not \U$10468 ( \10845 , \10166 );
or \U$10469 ( \10846 , \10844 , \10845 );
nand \U$10470 ( \10847 , \9854 , \2534 );
nand \U$10471 ( \10848 , \10846 , \10847 );
nand \U$10472 ( \10849 , \10843 , \10848 );
nand \U$10473 ( \10850 , \10842 , \10849 );
xor \U$10474 ( \10851 , \10823 , \10850 );
not \U$10475 ( \10852 , \1311 );
not \U$10476 ( \10853 , \9903 );
or \U$10477 ( \10854 , \10852 , \10853 );
not \U$10478 ( \10855 , RIc227100_11);
not \U$10479 ( \10856 , \8807 );
or \U$10480 ( \10857 , \10855 , \10856 );
not \U$10481 ( \10858 , \8806 );
not \U$10482 ( \10859 , \10858 );
nand \U$10483 ( \10860 , \10859 , \1291 );
nand \U$10484 ( \10861 , \10857 , \10860 );
nand \U$10485 ( \10862 , \10861 , \9904 );
nand \U$10486 ( \10863 , \10854 , \10862 );
not \U$10487 ( \10864 , \10863 );
not \U$10488 ( \10865 , \2320 );
not \U$10489 ( \10866 , \10146 );
or \U$10490 ( \10867 , \10865 , \10866 );
nand \U$10491 ( \10868 , \9863 , \2358 );
nand \U$10492 ( \10869 , \10867 , \10868 );
not \U$10493 ( \10870 , \10869 );
or \U$10494 ( \10871 , \10864 , \10870 );
or \U$10495 ( \10872 , \10869 , \10863 );
not \U$10496 ( \10873 , \1682 );
not \U$10497 ( \10874 , \9888 );
or \U$10498 ( \10875 , \10873 , \10874 );
not \U$10499 ( \10876 , \1679 );
not \U$10500 ( \10877 , RIc227010_13);
not \U$10501 ( \10878 , \10322 );
or \U$10502 ( \10879 , \10877 , \10878 );
nand \U$10503 ( \10880 , \8856 , \2427 );
nand \U$10504 ( \10881 , \10879 , \10880 );
nand \U$10505 ( \10882 , \10876 , \10881 );
nand \U$10506 ( \10883 , \10875 , \10882 );
nand \U$10507 ( \10884 , \10872 , \10883 );
nand \U$10508 ( \10885 , \10871 , \10884 );
and \U$10509 ( \10886 , \10851 , \10885 );
and \U$10510 ( \10887 , \10823 , \10850 );
or \U$10511 ( \10888 , \10886 , \10887 );
nand \U$10512 ( \10889 , \10797 , \10888 );
nand \U$10513 ( \10890 , \10793 , \10889 );
xor \U$10514 ( \10891 , \10785 , \10890 );
not \U$10515 ( \10892 , \2784 );
not \U$10516 ( \10893 , \10479 );
or \U$10517 ( \10894 , \10892 , \10893 );
not \U$10518 ( \10895 , RIc226890_29);
not \U$10519 ( \10896 , \3446 );
not \U$10520 ( \10897 , \10896 );
or \U$10521 ( \10898 , \10895 , \10897 );
not \U$10522 ( \10899 , \2554 );
not \U$10523 ( \10900 , RIc226890_29);
nand \U$10524 ( \10901 , \10899 , \10900 );
nand \U$10525 ( \10902 , \10898 , \10901 );
nand \U$10526 ( \10903 , \10902 , \9142 );
nand \U$10527 ( \10904 , \10894 , \10903 );
not \U$10528 ( \10905 , \9690 );
not \U$10529 ( \10906 , \10681 );
or \U$10530 ( \10907 , \10905 , \10906 );
not \U$10531 ( \10908 , RIc2262f0_41);
not \U$10532 ( \10909 , \1331 );
not \U$10533 ( \10910 , \10909 );
or \U$10534 ( \10911 , \10908 , \10910 );
nand \U$10535 ( \10912 , \1331 , \6303 );
nand \U$10536 ( \10913 , \10911 , \10912 );
nand \U$10537 ( \10914 , \10913 , \9705 );
nand \U$10538 ( \10915 , \10907 , \10914 );
xor \U$10539 ( \10916 , \10904 , \10915 );
not \U$10540 ( \10917 , \2138 );
not \U$10541 ( \10918 , \10667 );
or \U$10542 ( \10919 , \10917 , \10918 );
and \U$10543 ( \10920 , \4194 , \2133 );
not \U$10544 ( \10921 , \4194 );
and \U$10545 ( \10922 , \10921 , RIc226980_27);
or \U$10546 ( \10923 , \10920 , \10922 );
nand \U$10547 ( \10924 , \10923 , \2154 );
nand \U$10548 ( \10925 , \10919 , \10924 );
xnor \U$10549 ( \10926 , \10916 , \10925 );
not \U$10550 ( \10927 , \10926 );
not \U$10551 ( \10928 , \5519 );
not \U$10552 ( \10929 , RIc2264d0_37);
not \U$10553 ( \10930 , \8989 );
not \U$10554 ( \10931 , \10930 );
or \U$10555 ( \10932 , \10929 , \10931 );
buf \U$10556 ( \10933 , \2296 );
not \U$10557 ( \10934 , \10933 );
not \U$10558 ( \10935 , \10934 );
not \U$10559 ( \10936 , \10935 );
not \U$10560 ( \10937 , \10936 );
nand \U$10561 ( \10938 , \10937 , \4371 );
nand \U$10562 ( \10939 , \10932 , \10938 );
not \U$10563 ( \10940 , \10939 );
or \U$10564 ( \10941 , \10928 , \10940 );
nand \U$10565 ( \10942 , \10739 , \5509 );
nand \U$10566 ( \10943 , \10941 , \10942 );
not \U$10567 ( \10944 , \9459 );
not \U$10568 ( \10945 , \10519 );
or \U$10569 ( \10946 , \10944 , \10945 );
and \U$10570 ( \10947 , \930 , \9450 );
not \U$10571 ( \10948 , \930 );
and \U$10572 ( \10949 , \10948 , RIc225e40_51);
or \U$10573 ( \10950 , \10947 , \10949 );
nand \U$10574 ( \10951 , \10950 , \9444 );
nand \U$10575 ( \10952 , \10946 , \10951 );
buf \U$10576 ( \10953 , \9619 );
not \U$10577 ( \10954 , \10953 );
not \U$10578 ( \10955 , RIc226020_47);
not \U$10579 ( \10956 , \1557 );
or \U$10580 ( \10957 , \10955 , \10956 );
nand \U$10581 ( \10958 , \981 , \9624 );
nand \U$10582 ( \10959 , \10957 , \10958 );
not \U$10583 ( \10960 , \10959 );
or \U$10584 ( \10961 , \10954 , \10960 );
nand \U$10585 ( \10962 , \10717 , \9641 );
nand \U$10586 ( \10963 , \10961 , \10962 );
xor \U$10587 ( \10964 , \10952 , \10963 );
xor \U$10588 ( \10965 , \10943 , \10964 );
not \U$10589 ( \10966 , \10965 );
or \U$10590 ( \10967 , \10927 , \10966 );
or \U$10591 ( \10968 , \10926 , \10965 );
nand \U$10592 ( \10969 , \10967 , \10968 );
not \U$10593 ( \10970 , \2518 );
not \U$10594 ( \10971 , \9846 );
or \U$10595 ( \10972 , \10970 , \10971 );
nand \U$10596 ( \10973 , \10601 , \2534 );
nand \U$10597 ( \10974 , \10972 , \10973 );
not \U$10598 ( \10975 , \9274 );
not \U$10599 ( \10976 , \10975 );
nand \U$10600 ( \10977 , \10976 , RIc2275b0_1);
not \U$10601 ( \10978 , \10977 );
not \U$10602 ( \10979 , \10978 );
not \U$10603 ( \10980 , \1579 );
xor \U$10604 ( \10981 , RIc2275b0_1, \10110 );
not \U$10605 ( \10982 , \10981 );
or \U$10606 ( \10983 , \10980 , \10982 );
and \U$10607 ( \10984 , RIc2275b0_1, \9255 );
not \U$10608 ( \10985 , RIc2275b0_1);
not \U$10609 ( \10986 , \9250 );
and \U$10610 ( \10987 , \10985 , \10986 );
or \U$10611 ( \10988 , \10984 , \10987 );
nand \U$10612 ( \10989 , \10988 , \854 );
nand \U$10613 ( \10990 , \10983 , \10989 );
not \U$10614 ( \10991 , \10990 );
not \U$10615 ( \10992 , \10991 );
or \U$10616 ( \10993 , \10979 , \10992 );
nand \U$10617 ( \10994 , \10990 , \10977 );
nand \U$10618 ( \10995 , \10993 , \10994 );
xor \U$10619 ( \10996 , \10974 , \10995 );
not \U$10620 ( \10997 , \2367 );
not \U$10621 ( \10998 , \10507 );
or \U$10622 ( \10999 , \10997 , \10998 );
nand \U$10623 ( \11000 , \10836 , \2392 );
nand \U$10624 ( \11001 , \10999 , \11000 );
nand \U$10625 ( \11002 , \10266 , RIc2275b0_1);
not \U$10626 ( \11003 , \11002 );
or \U$10627 ( \11004 , \11001 , \11003 );
not \U$10628 ( \11005 , \854 );
not \U$10629 ( \11006 , \10804 );
or \U$10630 ( \11007 , \11005 , \11006 );
nand \U$10631 ( \11008 , \10988 , \1579 );
nand \U$10632 ( \11009 , \11007 , \11008 );
nand \U$10633 ( \11010 , \11004 , \11009 );
nand \U$10634 ( \11011 , \11001 , \11003 );
nand \U$10635 ( \11012 , \11010 , \11011 );
xor \U$10636 ( \11013 , \10996 , \11012 );
or \U$10637 ( \11014 , \9920 , \9906 );
nand \U$10638 ( \11015 , \11014 , \9892 );
nand \U$10639 ( \11016 , \9920 , \9906 );
nand \U$10640 ( \11017 , \11015 , \11016 );
and \U$10641 ( \11018 , \11013 , \11017 );
and \U$10642 ( \11019 , \10996 , \11012 );
or \U$10643 ( \11020 , \11018 , \11019 );
and \U$10644 ( \11021 , \10969 , \11020 );
not \U$10645 ( \11022 , \10969 );
not \U$10646 ( \11023 , \11020 );
and \U$10647 ( \11024 , \11022 , \11023 );
nor \U$10648 ( \11025 , \11021 , \11024 );
xnor \U$10649 ( \11026 , \10891 , \11025 );
not \U$10650 ( \11027 , \11026 );
and \U$10651 ( \11028 , \10702 , \11027 );
not \U$10652 ( \11029 , \10702 );
and \U$10653 ( \11030 , \11029 , \11026 );
nor \U$10654 ( \11031 , \11028 , \11030 );
xor \U$10655 ( \11032 , \10552 , \11031 );
not \U$10656 ( \11033 , RIc225b70_57);
and \U$10657 ( \11034 , \11033 , RIc225be8_56);
not \U$10658 ( \11035 , RIc225be8_56);
and \U$10659 ( \11036 , \11035 , RIc225b70_57);
nor \U$10660 ( \11037 , \11034 , \11036 );
not \U$10661 ( \11038 , \11037 );
not \U$10662 ( \11039 , \11038 );
not \U$10663 ( \11040 , \11039 );
not \U$10664 ( \11041 , RIc225c60_55);
and \U$10665 ( \11042 , \11041 , \11035 );
and \U$10666 ( \11043 , RIc225c60_55, RIc225be8_56);
nor \U$10667 ( \11044 , \11042 , \11043 );
and \U$10668 ( \11045 , \11037 , \11044 );
not \U$10669 ( \11046 , \11045 );
not \U$10670 ( \11047 , \11046 );
or \U$10671 ( \11048 , \11040 , \11047 );
nand \U$10672 ( \11049 , \11048 , RIc225c60_55);
not \U$10673 ( \11050 , \1082 );
not \U$10674 ( \11051 , \10658 );
or \U$10675 ( \11052 , \11050 , \11051 );
nand \U$10676 ( \11053 , \10818 , \1040 );
nand \U$10677 ( \11054 , \11052 , \11053 );
xor \U$10678 ( \11055 , \11049 , \11054 );
not \U$10679 ( \11056 , \954 );
not \U$10680 ( \11057 , \8929 );
or \U$10681 ( \11058 , \11056 , \11057 );
nand \U$10682 ( \11059 , \9053 , \950 );
nand \U$10683 ( \11060 , \11058 , \11059 );
and \U$10684 ( \11061 , \11055 , \11060 );
and \U$10685 ( \11062 , \11049 , \11054 );
or \U$10686 ( \11063 , \11061 , \11062 );
not \U$10687 ( \11064 , \2860 );
not \U$10688 ( \11065 , \9807 );
or \U$10689 ( \11066 , \11064 , \11065 );
not \U$10690 ( \11067 , RIc226a70_25);
not \U$10691 ( \11068 , \2042 );
not \U$10692 ( \11069 , \11068 );
or \U$10693 ( \11070 , \11067 , \11069 );
nand \U$10694 ( \11071 , \2730 , \2187 );
nand \U$10695 ( \11072 , \11070 , \11071 );
nand \U$10696 ( \11073 , \11072 , \2173 );
nand \U$10697 ( \11074 , \11066 , \11073 );
xor \U$10698 ( \11075 , \11063 , \11074 );
xor \U$10699 ( \11076 , \9856 , \9867 );
and \U$10700 ( \11077 , \11076 , \9879 );
and \U$10701 ( \11078 , \9856 , \9867 );
or \U$10702 ( \11079 , \11077 , \11078 );
xor \U$10703 ( \11080 , \11075 , \11079 );
not \U$10704 ( \11081 , \11080 );
not \U$10705 ( \11082 , \1120 );
not \U$10706 ( \11083 , \9792 );
or \U$10707 ( \11084 , \11082 , \11083 );
nand \U$10708 ( \11085 , \9218 , \1118 );
nand \U$10709 ( \11086 , \11084 , \11085 );
not \U$10710 ( \11087 , \11086 );
not \U$10711 ( \11088 , \1340 );
not \U$10712 ( \11089 , \9918 );
or \U$10713 ( \11090 , \11088 , \11089 );
not \U$10714 ( \11091 , RIc2271f0_9);
not \U$10715 ( \11092 , \8975 );
or \U$10716 ( \11093 , \11091 , \11092 );
not \U$10717 ( \11094 , \10748 );
not \U$10718 ( \11095 , \11094 );
nand \U$10719 ( \11096 , \11095 , \1351 );
nand \U$10720 ( \11097 , \11093 , \11096 );
nand \U$10721 ( \11098 , \11097 , \1363 );
nand \U$10722 ( \11099 , \11090 , \11098 );
not \U$10723 ( \11100 , \11099 );
or \U$10724 ( \11101 , \11087 , \11100 );
not \U$10725 ( \11102 , \11099 );
not \U$10726 ( \11103 , \11102 );
not \U$10727 ( \11104 , \11086 );
not \U$10728 ( \11105 , \11104 );
or \U$10729 ( \11106 , \11103 , \11105 );
not \U$10730 ( \11107 , \11039 );
not \U$10731 ( \11108 , RIc225c60_55);
not \U$10732 ( \11109 , \11108 );
and \U$10733 ( \11110 , \11107 , \11109 );
not \U$10734 ( \11111 , RIc225c60_55);
not \U$10735 ( \11112 , \930 );
not \U$10736 ( \11113 , \11112 );
or \U$10737 ( \11114 , \11111 , \11113 );
nand \U$10738 ( \11115 , \3957 , \8767 );
nand \U$10739 ( \11116 , \11114 , \11115 );
not \U$10740 ( \11117 , \11046 );
buf \U$10741 ( \11118 , \11117 );
and \U$10742 ( \11119 , \11116 , \11118 );
nor \U$10743 ( \11120 , \11110 , \11119 );
not \U$10744 ( \11121 , \11120 );
nand \U$10745 ( \11122 , \11106 , \11121 );
nand \U$10746 ( \11123 , \11101 , \11122 );
not \U$10747 ( \11124 , \11123 );
not \U$10748 ( \11125 , \11001 );
not \U$10749 ( \11126 , \11009 );
not \U$10750 ( \11127 , \11002 );
and \U$10751 ( \11128 , \11126 , \11127 );
and \U$10752 ( \11129 , \11009 , \11002 );
nor \U$10753 ( \11130 , \11128 , \11129 );
not \U$10754 ( \11131 , \11130 );
and \U$10755 ( \11132 , \11125 , \11131 );
and \U$10756 ( \11133 , \11130 , \11001 );
nor \U$10757 ( \11134 , \11132 , \11133 );
not \U$10758 ( \11135 , \11134 );
not \U$10759 ( \11136 , \11135 );
or \U$10760 ( \11137 , \11124 , \11136 );
or \U$10761 ( \11138 , \11123 , \11135 );
xor \U$10762 ( \11139 , \11049 , \11054 );
xor \U$10763 ( \11140 , \11139 , \11060 );
nand \U$10764 ( \11141 , \11138 , \11140 );
nand \U$10765 ( \11142 , \11137 , \11141 );
not \U$10766 ( \11143 , \11142 );
not \U$10767 ( \11144 , \11143 );
or \U$10768 ( \11145 , \11081 , \11144 );
or \U$10769 ( \11146 , \11143 , \11080 );
nand \U$10770 ( \11147 , \11145 , \11146 );
xor \U$10771 ( \11148 , \10996 , \11012 );
xor \U$10772 ( \11149 , \11148 , \11017 );
not \U$10773 ( \11150 , \11149 );
and \U$10774 ( \11151 , \11147 , \11150 );
not \U$10775 ( \11152 , \11147 );
and \U$10776 ( \11153 , \11152 , \11149 );
nor \U$10777 ( \11154 , \11151 , \11153 );
xor \U$10778 ( \11155 , \10787 , \10790 );
xor \U$10779 ( \11156 , \11155 , \10888 );
nand \U$10780 ( \11157 , \11154 , \11156 );
not \U$10781 ( \11158 , \11157 );
xor \U$10782 ( \11159 , \10823 , \10850 );
xor \U$10783 ( \11160 , \11159 , \10885 );
xor \U$10784 ( \11161 , \11140 , \11134 );
xnor \U$10785 ( \11162 , \11161 , \11123 );
xor \U$10786 ( \11163 , \11160 , \11162 );
not \U$10787 ( \11164 , \9398 );
not \U$10788 ( \11165 , \9933 );
or \U$10789 ( \11166 , \11164 , \11165 );
not \U$10790 ( \11167 , RIc226110_45);
not \U$10791 ( \11168 , \3783 );
or \U$10792 ( \11169 , \11167 , \11168 );
nand \U$10793 ( \11170 , \3043 , \9100 );
nand \U$10794 ( \11171 , \11169 , \11170 );
nand \U$10795 ( \11172 , \11171 , \9384 );
nand \U$10796 ( \11173 , \11166 , \11172 );
not \U$10797 ( \11174 , \11173 );
not \U$10798 ( \11175 , RIc2267a0_31);
not \U$10799 ( \11176 , \2670 );
or \U$10800 ( \11177 , \11175 , \11176 );
nand \U$10801 ( \11178 , \9139 , \2072 );
nand \U$10802 ( \11179 , \11177 , \11178 );
not \U$10803 ( \11180 , \11179 );
not \U$10804 ( \11181 , \11180 );
not \U$10805 ( \11182 , \2697 );
not \U$10806 ( \11183 , \11182 );
and \U$10807 ( \11184 , \11181 , \11183 );
and \U$10808 ( \11185 , \9161 , \2710 );
nor \U$10809 ( \11186 , \11184 , \11185 );
not \U$10810 ( \11187 , \11186 );
not \U$10811 ( \11188 , \11187 );
or \U$10812 ( \11189 , \11174 , \11188 );
not \U$10813 ( \11190 , \11173 );
not \U$10814 ( \11191 , \11190 );
not \U$10815 ( \11192 , \11186 );
or \U$10816 ( \11193 , \11191 , \11192 );
not \U$10817 ( \11194 , \3631 );
not \U$10818 ( \11195 , \9945 );
or \U$10819 ( \11196 , \11194 , \11195 );
not \U$10820 ( \11197 , \5185 );
not \U$10821 ( \11198 , RIc2266b0_33);
not \U$10822 ( \11199 , \2476 );
or \U$10823 ( \11200 , \11198 , \11199 );
nand \U$10824 ( \11201 , \3036 , \2692 );
nand \U$10825 ( \11202 , \11200 , \11201 );
nand \U$10826 ( \11203 , \11197 , \11202 );
nand \U$10827 ( \11204 , \11196 , \11203 );
nand \U$10828 ( \11205 , \11193 , \11204 );
nand \U$10829 ( \11206 , \11189 , \11205 );
not \U$10830 ( \11207 , \11121 );
not \U$10831 ( \11208 , \11104 );
or \U$10832 ( \11209 , \11207 , \11208 );
nand \U$10833 ( \11210 , \11086 , \11120 );
nand \U$10834 ( \11211 , \11209 , \11210 );
and \U$10835 ( \11212 , \11211 , \11099 );
not \U$10836 ( \11213 , \11211 );
and \U$10837 ( \11214 , \11213 , \11102 );
nor \U$10838 ( \11215 , \11212 , \11214 );
nor \U$10839 ( \11216 , \11206 , \11215 );
xor \U$10840 ( \11217 , \10883 , \10869 );
xnor \U$10841 ( \11218 , \11217 , \10863 );
or \U$10842 ( \11219 , \11216 , \11218 );
nand \U$10843 ( \11220 , \11206 , \11215 );
nand \U$10844 ( \11221 , \11219 , \11220 );
and \U$10845 ( \11222 , \11163 , \11221 );
and \U$10846 ( \11223 , \11160 , \11162 );
or \U$10847 ( \11224 , \11222 , \11223 );
not \U$10848 ( \11225 , \11224 );
or \U$10849 ( \11226 , \11158 , \11225 );
not \U$10850 ( \11227 , \11156 );
not \U$10851 ( \11228 , \11154 );
nand \U$10852 ( \11229 , \11227 , \11228 );
nand \U$10853 ( \11230 , \11226 , \11229 );
not \U$10854 ( \11231 , \4381 );
not \U$10855 ( \11232 , \10727 );
or \U$10856 ( \11233 , \11231 , \11232 );
not \U$10857 ( \11234 , RIc2265c0_35);
not \U$10858 ( \11235 , \2833 );
or \U$10859 ( \11236 , \11234 , \11235 );
nand \U$10860 ( \11237 , \2832 , \3620 );
nand \U$10861 ( \11238 , \11236 , \11237 );
nand \U$10862 ( \11239 , \11238 , \4383 );
nand \U$10863 ( \11240 , \11233 , \11239 );
not \U$10864 ( \11241 , \11240 );
not \U$10865 ( \11242 , \2256 );
not \U$10866 ( \11243 , \2692 );
and \U$10867 ( \11244 , \11242 , \11243 );
and \U$10868 ( \11245 , \4008 , \2692 );
nor \U$10869 ( \11246 , \11244 , \11245 );
not \U$10870 ( \11247 , \11246 );
not \U$10871 ( \11248 , \4440 );
and \U$10872 ( \11249 , \11247 , \11248 );
and \U$10873 ( \11250 , \10442 , \3629 );
nor \U$10874 ( \11251 , \11249 , \11250 );
not \U$10875 ( \11252 , \11251 );
or \U$10876 ( \11253 , \11241 , \11252 );
or \U$10877 ( \11254 , \11240 , \11251 );
nand \U$10878 ( \11255 , \11253 , \11254 );
not \U$10879 ( \11256 , \9398 );
not \U$10880 ( \11257 , RIc226110_45);
not \U$10881 ( \11258 , \9539 );
or \U$10882 ( \11259 , \11257 , \11258 );
not \U$10883 ( \11260 , \1169 );
not \U$10884 ( \11261 , \11260 );
nand \U$10885 ( \11262 , \11261 , \10429 );
nand \U$10886 ( \11263 , \11259 , \11262 );
not \U$10887 ( \11264 , \11263 );
or \U$10888 ( \11265 , \11256 , \11264 );
nand \U$10889 ( \11266 , \10431 , \9934 );
nand \U$10890 ( \11267 , \11265 , \11266 );
not \U$10891 ( \11268 , \11267 );
and \U$10892 ( \11269 , \11255 , \11268 );
not \U$10893 ( \11270 , \11255 );
and \U$10894 ( \11271 , \11270 , \11267 );
nor \U$10895 ( \11272 , \11269 , \11271 );
not \U$10896 ( \11273 , \9129 );
not \U$10897 ( \11274 , RIc226200_43);
not \U$10898 ( \11275 , \1392 );
or \U$10899 ( \11276 , \11274 , \11275 );
nand \U$10900 ( \11277 , \1391 , \9125 );
nand \U$10901 ( \11278 , \11276 , \11277 );
not \U$10902 ( \11279 , \11278 );
or \U$10903 ( \11280 , \11273 , \11279 );
nand \U$10904 ( \11281 , \10490 , \9110 );
nand \U$10905 ( \11282 , \11280 , \11281 );
not \U$10906 ( \11283 , \10445 );
not \U$10907 ( \11284 , \10454 );
or \U$10908 ( \11285 , \11283 , \11284 );
not \U$10909 ( \11286 , RIc225f30_49);
not \U$10910 ( \11287 , \4024 );
or \U$10911 ( \11288 , \11286 , \11287 );
not \U$10912 ( \11289 , RIc225f30_49);
nand \U$10913 ( \11290 , \888 , \11289 );
nand \U$10914 ( \11291 , \11288 , \11290 );
nand \U$10915 ( \11292 , \11291 , \9552 );
nand \U$10916 ( \11293 , \11285 , \11292 );
xor \U$10917 ( \11294 , \11282 , \11293 );
not \U$10918 ( \11295 , \2697 );
not \U$10919 ( \11296 , \10468 );
or \U$10920 ( \11297 , \11295 , \11296 );
not \U$10921 ( \11298 , RIc2267a0_31);
not \U$10922 ( \11299 , \9584 );
or \U$10923 ( \11300 , \11298 , \11299 );
nand \U$10924 ( \11301 , \2014 , \3648 );
nand \U$10925 ( \11302 , \11300 , \11301 );
nand \U$10926 ( \11303 , \11302 , \2710 );
nand \U$10927 ( \11304 , \11297 , \11303 );
xor \U$10928 ( \11305 , \11294 , \11304 );
xor \U$10929 ( \11306 , \11272 , \11305 );
not \U$10930 ( \11307 , \6689 );
not \U$10931 ( \11308 , \9000 );
or \U$10932 ( \11309 , \11307 , \11308 );
not \U$10933 ( \11310 , RIc2263e0_39);
not \U$10934 ( \11311 , \4181 );
or \U$10935 ( \11312 , \11310 , \11311 );
nand \U$10936 ( \11313 , \1729 , \8990 );
nand \U$10937 ( \11314 , \11312 , \11313 );
nand \U$10938 ( \11315 , \11314 , \6307 );
nand \U$10939 ( \11316 , \11309 , \11315 );
not \U$10940 ( \11317 , \2367 );
not \U$10941 ( \11318 , RIc226c50_21);
not \U$10942 ( \11319 , \3114 );
not \U$10943 ( \11320 , \11319 );
not \U$10944 ( \11321 , \11320 );
not \U$10945 ( \11322 , \11321 );
or \U$10946 ( \11323 , \11318 , \11322 );
not \U$10947 ( \11324 , \11319 );
nand \U$10948 ( \11325 , \11324 , \2370 );
nand \U$10949 ( \11326 , \11323 , \11325 );
not \U$10950 ( \11327 , \11326 );
or \U$10951 ( \11328 , \11317 , \11327 );
nand \U$10952 ( \11329 , \10500 , \2392 );
nand \U$10953 ( \11330 , \11328 , \11329 );
xor \U$10954 ( \11331 , \11316 , \11330 );
not \U$10955 ( \11332 , \1915 );
not \U$10956 ( \11333 , \10535 );
or \U$10957 ( \11334 , \11332 , \11333 );
not \U$10958 ( \11335 , RIc226b60_23);
not \U$10959 ( \11336 , \9188 );
or \U$10960 ( \11337 , \11335 , \11336 );
nand \U$10961 ( \11338 , \9805 , \1927 );
nand \U$10962 ( \11339 , \11337 , \11338 );
nand \U$10963 ( \11340 , \11339 , \5365 );
nand \U$10964 ( \11341 , \11334 , \11340 );
xnor \U$10965 ( \11342 , \11331 , \11341 );
xor \U$10966 ( \11343 , \11306 , \11342 );
not \U$10967 ( \11344 , \11143 );
not \U$10968 ( \11345 , \11344 );
buf \U$10969 ( \11346 , \11080 );
not \U$10970 ( \11347 , \11346 );
or \U$10971 ( \11348 , \11345 , \11347 );
or \U$10972 ( \11349 , \11344 , \11346 );
nand \U$10973 ( \11350 , \11349 , \11149 );
nand \U$10974 ( \11351 , \11348 , \11350 );
xor \U$10975 ( \11352 , \11343 , \11351 );
not \U$10976 ( \11353 , \10660 );
not \U$10977 ( \11354 , \11353 );
not \U$10978 ( \11355 , \2195 );
not \U$10979 ( \11356 , \11072 );
or \U$10980 ( \11357 , \11355 , \11356 );
not \U$10981 ( \11358 , RIc226a70_25);
not \U$10982 ( \11359 , \3009 );
or \U$10983 ( \11360 , \11358 , \11359 );
nand \U$10984 ( \11361 , \2064 , \1905 );
nand \U$10985 ( \11362 , \11360 , \11361 );
nand \U$10986 ( \11363 , \11362 , \2173 );
nand \U$10987 ( \11364 , \11357 , \11363 );
not \U$10988 ( \11365 , \11364 );
not \U$10989 ( \11366 , \11365 );
or \U$10990 ( \11367 , \11354 , \11366 );
nand \U$10991 ( \11368 , \11364 , \10660 );
nand \U$10992 ( \11369 , \11367 , \11368 );
xor \U$10993 ( \11370 , \8790 , \8837 );
and \U$10994 ( \11371 , \11370 , \8893 );
and \U$10995 ( \11372 , \8790 , \8837 );
or \U$10996 ( \11373 , \11371 , \11372 );
not \U$10997 ( \11374 , \11373 );
and \U$10998 ( \11375 , \11369 , \11374 );
not \U$10999 ( \11376 , \11369 );
and \U$11000 ( \11377 , \11376 , \11373 );
nor \U$11001 ( \11378 , \11375 , \11377 );
not \U$11002 ( \11379 , \11378 );
not \U$11003 ( \11380 , \11379 );
xor \U$11004 ( \11381 , \11063 , \11074 );
and \U$11005 ( \11382 , \11381 , \11079 );
and \U$11006 ( \11383 , \11063 , \11074 );
or \U$11007 ( \11384 , \11382 , \11383 );
not \U$11008 ( \11385 , \11384 );
not \U$11009 ( \11386 , \11385 );
or \U$11010 ( \11387 , \11380 , \11386 );
nand \U$11011 ( \11388 , \11384 , \11378 );
nand \U$11012 ( \11389 , \11387 , \11388 );
and \U$11013 ( \11390 , \8776 , \8787 );
not \U$11014 ( \11391 , RIc225d50_53);
nor \U$11015 ( \11392 , \11390 , \11391 );
not \U$11016 ( \11393 , \1579 );
not \U$11017 ( \11394 , \9072 );
and \U$11018 ( \11395 , RIc2275b0_1, \11394 );
not \U$11019 ( \11396 , RIc2275b0_1);
and \U$11020 ( \11397 , \11396 , \9072 );
or \U$11021 ( \11398 , \11395 , \11397 );
not \U$11022 ( \11399 , \11398 );
or \U$11023 ( \11400 , \11393 , \11399 );
nand \U$11024 ( \11401 , \854 , \10981 );
nand \U$11025 ( \11402 , \11400 , \11401 );
xor \U$11026 ( \11403 , \11392 , \11402 );
not \U$11027 ( \11404 , \1082 );
not \U$11028 ( \11405 , \8924 );
not \U$11029 ( \11406 , \11405 );
and \U$11030 ( \11407 , RIc2274c0_3, \11406 );
not \U$11031 ( \11408 , RIc2274c0_3);
and \U$11032 ( \11409 , \11408 , \11405 );
nor \U$11033 ( \11410 , \11407 , \11409 );
not \U$11034 ( \11411 , \11410 );
or \U$11035 ( \11412 , \11404 , \11411 );
nand \U$11036 ( \11413 , \10649 , \1040 );
nand \U$11037 ( \11414 , \11412 , \11413 );
xor \U$11038 ( \11415 , \11403 , \11414 );
not \U$11039 ( \11416 , \11415 );
not \U$11040 ( \11417 , \11416 );
nand \U$11041 ( \11418 , \10991 , \10977 );
not \U$11042 ( \11419 , \11418 );
not \U$11043 ( \11420 , \10974 );
or \U$11044 ( \11421 , \11419 , \11420 );
nand \U$11045 ( \11422 , \10990 , \10978 );
nand \U$11046 ( \11423 , \11421 , \11422 );
not \U$11047 ( \11424 , \11423 );
not \U$11048 ( \11425 , \11424 );
or \U$11049 ( \11426 , \11417 , \11425 );
nand \U$11050 ( \11427 , \11415 , \11423 );
nand \U$11051 ( \11428 , \11426 , \11427 );
xor \U$11052 ( \11429 , \9744 , \9762 );
and \U$11053 ( \11430 , \11429 , \9782 );
and \U$11054 ( \11431 , \9744 , \9762 );
or \U$11055 ( \11432 , \11430 , \11431 );
and \U$11056 ( \11433 , \11428 , \11432 );
not \U$11057 ( \11434 , \11428 );
not \U$11058 ( \11435 , \11432 );
and \U$11059 ( \11436 , \11434 , \11435 );
nor \U$11060 ( \11437 , \11433 , \11436 );
buf \U$11061 ( \11438 , \11437 );
not \U$11062 ( \11439 , \11438 );
and \U$11063 ( \11440 , \11389 , \11439 );
not \U$11064 ( \11441 , \11389 );
and \U$11065 ( \11442 , \11441 , \11438 );
nor \U$11066 ( \11443 , \11440 , \11442 );
xor \U$11067 ( \11444 , \11352 , \11443 );
xor \U$11068 ( \11445 , \11230 , \11444 );
xor \U$11069 ( \11446 , \9966 , \9714 );
xor \U$11070 ( \11447 , \11446 , \9835 );
not \U$11071 ( \11448 , \11447 );
not \U$11072 ( \11449 , \11448 );
xor \U$11073 ( \11450 , \9880 , \9921 );
xor \U$11074 ( \11451 , \11450 , \9964 );
not \U$11075 ( \11452 , \11451 );
not \U$11076 ( \11453 , \11452 );
not \U$11077 ( \11454 , \9962 );
xor \U$11078 ( \11455 , \9949 , \11454 );
xor \U$11079 ( \11456 , \11455 , \9936 );
xor \U$11080 ( \11457 , \9564 , \9554 );
xnor \U$11081 ( \11458 , \11457 , \9577 );
nand \U$11082 ( \11459 , \11456 , \11458 );
xor \U$11083 ( \11460 , \9081 , \9170 );
xnor \U$11084 ( \11461 , \11460 , \9152 );
not \U$11085 ( \11462 , \11461 );
and \U$11086 ( \11463 , \11459 , \11462 );
nor \U$11087 ( \11464 , \11458 , \11456 );
nor \U$11088 ( \11465 , \11463 , \11464 );
not \U$11089 ( \11466 , \11465 );
not \U$11090 ( \11467 , \11466 );
or \U$11091 ( \11468 , \11453 , \11467 );
not \U$11092 ( \11469 , \11451 );
not \U$11093 ( \11470 , \11465 );
or \U$11094 ( \11471 , \11469 , \11470 );
xor \U$11095 ( \11472 , \10848 , \10840 );
xor \U$11096 ( \11473 , \11472 , \10828 );
not \U$11097 ( \11474 , \1120 );
not \U$11098 ( \11475 , \9227 );
or \U$11099 ( \11476 , \11474 , \11475 );
not \U$11100 ( \11477 , RIc2272e0_7);
buf \U$11101 ( \11478 , \9076 );
not \U$11102 ( \11479 , \11478 );
or \U$11103 ( \11480 , \11477 , \11479 );
nand \U$11104 ( \11481 , \9077 , \1139 );
nand \U$11105 ( \11482 , \11480 , \11481 );
nand \U$11106 ( \11483 , \11482 , \1118 );
nand \U$11107 ( \11484 , \11476 , \11483 );
not \U$11108 ( \11485 , \11484 );
not \U$11109 ( \11486 , \951 );
not \U$11110 ( \11487 , RIc2273d0_5);
not \U$11111 ( \11488 , \9254 );
not \U$11112 ( \11489 , \11488 );
or \U$11113 ( \11490 , \11487 , \11489 );
nand \U$11114 ( \11491 , \10986 , \946 );
nand \U$11115 ( \11492 , \11490 , \11491 );
not \U$11116 ( \11493 , \11492 );
or \U$11117 ( \11494 , \11486 , \11493 );
nand \U$11118 ( \11495 , \10115 , \954 );
nand \U$11119 ( \11496 , \11494 , \11495 );
not \U$11120 ( \11497 , \11496 );
or \U$11121 ( \11498 , \11485 , \11497 );
or \U$11122 ( \11499 , \11484 , \11496 );
not \U$11123 ( \11500 , \1579 );
not \U$11124 ( \11501 , \9326 );
or \U$11125 ( \11502 , \11500 , \11501 );
nand \U$11126 ( \11503 , \10364 , \854 );
nand \U$11127 ( \11504 , \11502 , \11503 );
nand \U$11128 ( \11505 , \11499 , \11504 );
nand \U$11129 ( \11506 , \11498 , \11505 );
xor \U$11130 ( \11507 , \10079 , \10087 );
xor \U$11131 ( \11508 , \11507 , \10117 );
xor \U$11132 ( \11509 , \11506 , \11508 );
not \U$11133 ( \11510 , \2086 );
not \U$11134 ( \11511 , \9150 );
or \U$11135 ( \11512 , \11510 , \11511 );
and \U$11136 ( \11513 , RIc226890_29, \3798 );
not \U$11137 ( \11514 , RIc226890_29);
not \U$11138 ( \11515 , \3798 );
and \U$11139 ( \11516 , \11514 , \11515 );
or \U$11140 ( \11517 , \11513 , \11516 );
nand \U$11141 ( \11518 , \11517 , \2784 );
nand \U$11142 ( \11519 , \11512 , \11518 );
and \U$11143 ( \11520 , \11509 , \11519 );
and \U$11144 ( \11521 , \11506 , \11508 );
or \U$11145 ( \11522 , \11520 , \11521 );
xor \U$11146 ( \11523 , \11473 , \11522 );
not \U$11147 ( \11524 , \9207 );
not \U$11148 ( \11525 , \9193 );
not \U$11149 ( \11526 , \11525 );
or \U$11150 ( \11527 , \11524 , \11526 );
or \U$11151 ( \11528 , \11525 , \9207 );
nand \U$11152 ( \11529 , \11527 , \11528 );
not \U$11153 ( \11530 , \11529 );
xor \U$11154 ( \11531 , \9331 , \11530 );
and \U$11155 ( \11532 , \11523 , \11531 );
and \U$11156 ( \11533 , \11473 , \11522 );
or \U$11157 ( \11534 , \11532 , \11533 );
nand \U$11158 ( \11535 , \11471 , \11534 );
nand \U$11159 ( \11536 , \11468 , \11535 );
not \U$11160 ( \11537 , \11536 );
or \U$11161 ( \11538 , \11449 , \11537 );
not \U$11162 ( \11539 , \11536 );
not \U$11163 ( \11540 , \11539 );
not \U$11164 ( \11541 , \11447 );
or \U$11165 ( \11542 , \11540 , \11541 );
xor \U$11166 ( \11543 , \10798 , \10808 );
xor \U$11167 ( \11544 , \11543 , \10820 );
not \U$11168 ( \11545 , \1682 );
not \U$11169 ( \11546 , \10881 );
or \U$11170 ( \11547 , \11545 , \11546 );
nand \U$11171 ( \11548 , \10291 , \1678 );
nand \U$11172 ( \11549 , \11547 , \11548 );
not \U$11173 ( \11550 , \1340 );
not \U$11174 ( \11551 , \11097 );
or \U$11175 ( \11552 , \11550 , \11551 );
not \U$11176 ( \11553 , RIc2271f0_9);
not \U$11177 ( \11554 , \9787 );
or \U$11178 ( \11555 , \11553 , \11554 );
nand \U$11179 ( \11556 , \9790 , \1342 );
nand \U$11180 ( \11557 , \11555 , \11556 );
nand \U$11181 ( \11558 , \11557 , \1363 );
nand \U$11182 ( \11559 , \11552 , \11558 );
xor \U$11183 ( \11560 , \11549 , \11559 );
not \U$11184 ( \11561 , \1311 );
not \U$11185 ( \11562 , \10861 );
or \U$11186 ( \11563 , \11561 , \11562 );
not \U$11187 ( \11564 , RIc227100_11);
not \U$11188 ( \11565 , \8951 );
buf \U$11189 ( \11566 , \11565 );
not \U$11190 ( \11567 , \11566 );
or \U$11191 ( \11568 , \11564 , \11567 );
nand \U$11192 ( \11569 , \8952 , \1291 );
nand \U$11193 ( \11570 , \11568 , \11569 );
nand \U$11194 ( \11571 , \11570 , \1307 );
nand \U$11195 ( \11572 , \11563 , \11571 );
and \U$11196 ( \11573 , \11560 , \11572 );
and \U$11197 ( \11574 , \11549 , \11559 );
or \U$11198 ( \11575 , \11573 , \11574 );
xor \U$11199 ( \11576 , \11544 , \11575 );
buf \U$11200 ( \11577 , \8788 );
not \U$11201 ( \11578 , \11577 );
not \U$11202 ( \11579 , \9562 );
or \U$11203 ( \11580 , \11578 , \11579 );
not \U$11204 ( \11581 , RIc225d50_53);
not \U$11205 ( \11582 , \840 );
not \U$11206 ( \11583 , \11582 );
or \U$11207 ( \11584 , \11581 , \11583 );
not \U$11208 ( \11585 , RIc225d50_53);
nand \U$11209 ( \11586 , \840 , \11585 );
nand \U$11210 ( \11587 , \11584 , \11586 );
nand \U$11211 ( \11588 , \11587 , \8777 );
nand \U$11212 ( \11589 , \11580 , \11588 );
not \U$11213 ( \11590 , \11589 );
not \U$11214 ( \11591 , \4383 );
not \U$11215 ( \11592 , \9589 );
or \U$11216 ( \11593 , \11591 , \11592 );
not \U$11217 ( \11594 , RIc2265c0_35);
not \U$11218 ( \11595 , \2586 );
or \U$11219 ( \11596 , \11594 , \11595 );
nand \U$11220 ( \11597 , \3183 , \3620 );
nand \U$11221 ( \11598 , \11596 , \11597 );
nand \U$11222 ( \11599 , \11598 , \4381 );
nand \U$11223 ( \11600 , \11593 , \11599 );
not \U$11224 ( \11601 , \9619 );
not \U$11225 ( \11602 , \9633 );
or \U$11226 ( \11603 , \11601 , \11602 );
not \U$11227 ( \11604 , RIc226020_47);
not \U$11228 ( \11605 , \1530 );
or \U$11229 ( \11606 , \11604 , \11605 );
not \U$11230 ( \11607 , RIc226020_47);
nand \U$11231 ( \11608 , \1529 , \11607 );
nand \U$11232 ( \11609 , \11606 , \11608 );
nand \U$11233 ( \11610 , \11609 , \9641 );
nand \U$11234 ( \11611 , \11603 , \11610 );
nor \U$11235 ( \11612 , \11600 , \11611 );
or \U$11236 ( \11613 , \11590 , \11612 );
nand \U$11237 ( \11614 , \11611 , \11600 );
nand \U$11238 ( \11615 , \11613 , \11614 );
and \U$11239 ( \11616 , \11576 , \11615 );
and \U$11240 ( \11617 , \11544 , \11575 );
or \U$11241 ( \11618 , \11616 , \11617 );
not \U$11242 ( \11619 , \5509 );
not \U$11243 ( \11620 , RIc2264d0_37);
not \U$11244 ( \11621 , \9408 );
or \U$11245 ( \11622 , \11620 , \11621 );
not \U$11246 ( \11623 , RIc2264d0_37);
nand \U$11247 ( \11624 , \11623 , \3838 );
nand \U$11248 ( \11625 , \11622 , \11624 );
not \U$11249 ( \11626 , \11625 );
or \U$11250 ( \11627 , \11619 , \11626 );
nand \U$11251 ( \11628 , \9610 , \5519 );
nand \U$11252 ( \11629 , \11627 , \11628 );
not \U$11253 ( \11630 , \9552 );
not \U$11254 ( \11631 , \9543 );
or \U$11255 ( \11632 , \11630 , \11631 );
not \U$11256 ( \11633 , RIc225f30_49);
not \U$11257 ( \11634 , \10427 );
or \U$11258 ( \11635 , \11633 , \11634 );
not \U$11259 ( \11636 , \1222 );
nand \U$11260 ( \11637 , \11636 , \9996 );
nand \U$11261 ( \11638 , \11635 , \11637 );
nand \U$11262 ( \11639 , \11638 , \9534 );
nand \U$11263 ( \11640 , \11632 , \11639 );
xor \U$11264 ( \11641 , \11629 , \11640 );
not \U$11265 ( \11642 , \6307 );
not \U$11266 ( \11643 , \9575 );
or \U$11267 ( \11644 , \11642 , \11643 );
not \U$11268 ( \11645 , RIc2263e0_39);
not \U$11269 ( \11646 , \2233 );
or \U$11270 ( \11647 , \11645 , \11646 );
buf \U$11271 ( \11648 , \2225 );
nand \U$11272 ( \11649 , \11648 , \8998 );
nand \U$11273 ( \11650 , \11647 , \11649 );
nand \U$11274 ( \11651 , \11650 , \6689 );
nand \U$11275 ( \11652 , \11644 , \11651 );
and \U$11276 ( \11653 , \11641 , \11652 );
and \U$11277 ( \11654 , \11629 , \11640 );
or \U$11278 ( \11655 , \11653 , \11654 );
not \U$11279 ( \11656 , \11655 );
not \U$11280 ( \11657 , \11656 );
not \U$11281 ( \11658 , \9129 );
not \U$11282 ( \11659 , \9202 );
or \U$11283 ( \11660 , \11658 , \11659 );
not \U$11284 ( \11661 , RIc226200_43);
not \U$11285 ( \11662 , \4473 );
or \U$11286 ( \11663 , \11661 , \11662 );
nand \U$11287 ( \11664 , \2353 , \9125 );
nand \U$11288 ( \11665 , \11663 , \11664 );
nand \U$11289 ( \11666 , \11665 , \9110 );
nand \U$11290 ( \11667 , \11660 , \11666 );
not \U$11291 ( \11668 , \11667 );
not \U$11292 ( \11669 , \2172 );
not \U$11293 ( \11670 , \9664 );
or \U$11294 ( \11671 , \11669 , \11670 );
not \U$11295 ( \11672 , \2980 );
and \U$11296 ( \11673 , \11672 , RIc226a70_25);
not \U$11297 ( \11674 , \11672 );
and \U$11298 ( \11675 , \11674 , \1905 );
or \U$11299 ( \11676 , \11673 , \11675 );
nand \U$11300 ( \11677 , \11676 , \2860 );
nand \U$11301 ( \11678 , \11671 , \11677 );
not \U$11302 ( \11679 , \11678 );
or \U$11303 ( \11680 , \11668 , \11679 );
or \U$11304 ( \11681 , \11667 , \11678 );
not \U$11305 ( \11682 , \2154 );
not \U$11306 ( \11683 , \9191 );
or \U$11307 ( \11684 , \11682 , \11683 );
not \U$11308 ( \11685 , RIc226980_27);
not \U$11309 ( \11686 , \3715 );
or \U$11310 ( \11687 , \11685 , \11686 );
nand \U$11311 ( \11688 , \9654 , \2150 );
nand \U$11312 ( \11689 , \11687 , \11688 );
nand \U$11313 ( \11690 , \11689 , \2138 );
nand \U$11314 ( \11691 , \11684 , \11690 );
nand \U$11315 ( \11692 , \11681 , \11691 );
nand \U$11316 ( \11693 , \11680 , \11692 );
not \U$11317 ( \11694 , \11693 );
not \U$11318 ( \11695 , \11694 );
or \U$11319 ( \11696 , \11657 , \11695 );
buf \U$11320 ( \11697 , \11045 );
not \U$11321 ( \11698 , \11697 );
not \U$11322 ( \11699 , RIc225c60_55);
not \U$11323 ( \11700 , \9491 );
or \U$11324 ( \11701 , \11699 , \11700 );
nand \U$11325 ( \11702 , \1072 , \8767 );
nand \U$11326 ( \11703 , \11701 , \11702 );
not \U$11327 ( \11704 , \11703 );
or \U$11328 ( \11705 , \11698 , \11704 );
nand \U$11329 ( \11706 , \11116 , \11038 );
nand \U$11330 ( \11707 , \11705 , \11706 );
buf \U$11331 ( \11708 , \9445 );
not \U$11332 ( \11709 , \11708 );
not \U$11333 ( \11710 , \9958 );
or \U$11334 ( \11711 , \11709 , \11710 );
and \U$11335 ( \11712 , RIc225e40_51, \2118 );
not \U$11336 ( \11713 , RIc225e40_51);
not \U$11337 ( \11714 , \2117 );
not \U$11338 ( \11715 , \11714 );
and \U$11339 ( \11716 , \11713 , \11715 );
or \U$11340 ( \11717 , \11712 , \11716 );
nand \U$11341 ( \11718 , \11717 , \9459 );
nand \U$11342 ( \11719 , \11711 , \11718 );
xor \U$11343 ( \11720 , \11707 , \11719 );
not \U$11344 ( \11721 , \9705 );
not \U$11345 ( \11722 , \9696 );
or \U$11346 ( \11723 , \11721 , \11722 );
not \U$11347 ( \11724 , RIc2262f0_41);
not \U$11348 ( \11725 , \9479 );
or \U$11349 ( \11726 , \11724 , \11725 );
nand \U$11350 ( \11727 , \2422 , \6303 );
nand \U$11351 ( \11728 , \11726 , \11727 );
nand \U$11352 ( \11729 , \11728 , \9690 );
nand \U$11353 ( \11730 , \11723 , \11729 );
and \U$11354 ( \11731 , \11720 , \11730 );
and \U$11355 ( \11732 , \11707 , \11719 );
or \U$11356 ( \11733 , \11731 , \11732 );
nand \U$11357 ( \11734 , \11696 , \11733 );
nand \U$11358 ( \11735 , \11693 , \11655 );
nand \U$11359 ( \11736 , \11734 , \11735 );
xor \U$11360 ( \11737 , \11618 , \11736 );
not \U$11361 ( \11738 , \9709 );
xor \U$11362 ( \11739 , \9646 , \11738 );
xor \U$11363 ( \11740 , \9712 , \11739 );
and \U$11364 ( \11741 , \11737 , \11740 );
and \U$11365 ( \11742 , \11618 , \11736 );
or \U$11366 ( \11743 , \11741 , \11742 );
nand \U$11367 ( \11744 , \11542 , \11743 );
nand \U$11368 ( \11745 , \11538 , \11744 );
xor \U$11369 ( \11746 , \11445 , \11745 );
xor \U$11370 ( \11747 , \11156 , \11224 );
xor \U$11371 ( \11748 , \11747 , \11228 );
not \U$11372 ( \11749 , \11748 );
not \U$11373 ( \11750 , \11749 );
xor \U$11374 ( \11751 , \10120 , \10178 );
xor \U$11375 ( \11752 , \11751 , \10238 );
xor \U$11376 ( \11753 , \11544 , \11575 );
xor \U$11377 ( \11754 , \11753 , \11615 );
xor \U$11378 ( \11755 , \11752 , \11754 );
not \U$11379 ( \11756 , \5135 );
not \U$11380 ( \11757 , \11598 );
or \U$11381 ( \11758 , \11756 , \11757 );
not \U$11382 ( \11759 , RIc2265c0_35);
not \U$11383 ( \11760 , \10896 );
or \U$11384 ( \11761 , \11759 , \11760 );
nand \U$11385 ( \11762 , \3446 , \3620 );
nand \U$11386 ( \11763 , \11761 , \11762 );
nand \U$11387 ( \11764 , \11763 , \5741 );
nand \U$11388 ( \11765 , \11758 , \11764 );
not \U$11389 ( \11766 , \9641 );
not \U$11390 ( \11767 , RIc226020_47);
not \U$11391 ( \11768 , \3438 );
or \U$11392 ( \11769 , \11767 , \11768 );
nand \U$11393 ( \11770 , \1332 , \9624 );
nand \U$11394 ( \11771 , \11769 , \11770 );
not \U$11395 ( \11772 , \11771 );
or \U$11396 ( \11773 , \11766 , \11772 );
nand \U$11397 ( \11774 , \11609 , \10953 );
nand \U$11398 ( \11775 , \11773 , \11774 );
or \U$11399 ( \11776 , \11765 , \11775 );
not \U$11400 ( \11777 , \11577 );
not \U$11401 ( \11778 , \11587 );
or \U$11402 ( \11779 , \11777 , \11778 );
and \U$11403 ( \11780 , RIc225d50_53, \1557 );
not \U$11404 ( \11781 , RIc225d50_53);
and \U$11405 ( \11782 , \11781 , \981 );
or \U$11406 ( \11783 , \11780 , \11782 );
nand \U$11407 ( \11784 , \11783 , \8777 );
nand \U$11408 ( \11785 , \11779 , \11784 );
nand \U$11409 ( \11786 , \11776 , \11785 );
nand \U$11410 ( \11787 , \11765 , \11775 );
nand \U$11411 ( \11788 , \11786 , \11787 );
not \U$11412 ( \11789 , \11717 );
not \U$11413 ( \11790 , \11708 );
or \U$11414 ( \11791 , \11789 , \11790 );
not \U$11415 ( \11792 , RIc225e40_51);
not \U$11416 ( \11793 , \9539 );
or \U$11417 ( \11794 , \11792 , \11793 );
not \U$11418 ( \11795 , RIc225e40_51);
nand \U$11419 ( \11796 , \1169 , \11795 );
nand \U$11420 ( \11797 , \11794 , \11796 );
nand \U$11421 ( \11798 , \11797 , \9458 );
nand \U$11422 ( \11799 , \11791 , \11798 );
not \U$11423 ( \11800 , \11118 );
not \U$11424 ( \11801 , RIc225c60_55);
not \U$11425 ( \11802 , \4024 );
or \U$11426 ( \11803 , \11801 , \11802 );
nand \U$11427 ( \11804 , \888 , \11041 );
nand \U$11428 ( \11805 , \11803 , \11804 );
not \U$11429 ( \11806 , \11805 );
or \U$11430 ( \11807 , \11800 , \11806 );
nand \U$11431 ( \11808 , \11703 , \11038 );
nand \U$11432 ( \11809 , \11807 , \11808 );
xor \U$11433 ( \11810 , \11799 , \11809 );
not \U$11434 ( \11811 , \9816 );
not \U$11435 ( \11812 , \11728 );
or \U$11436 ( \11813 , \11811 , \11812 );
not \U$11437 ( \11814 , RIc2262f0_41);
not \U$11438 ( \11815 , \2444 );
or \U$11439 ( \11816 , \11814 , \11815 );
nand \U$11440 ( \11817 , \2443 , \6303 );
nand \U$11441 ( \11818 , \11816 , \11817 );
nand \U$11442 ( \11819 , \11818 , \9690 );
nand \U$11443 ( \11820 , \11813 , \11819 );
and \U$11444 ( \11821 , \11810 , \11820 );
and \U$11445 ( \11822 , \11799 , \11809 );
or \U$11446 ( \11823 , \11821 , \11822 );
xor \U$11447 ( \11824 , \11788 , \11823 );
buf \U$11448 ( \11825 , \9398 );
not \U$11449 ( \11826 , \11825 );
not \U$11450 ( \11827 , \11171 );
or \U$11451 ( \11828 , \11826 , \11827 );
and \U$11452 ( \11829 , RIc226110_45, \1729 );
not \U$11453 ( \11830 , RIc226110_45);
not \U$11454 ( \11831 , \1728 );
and \U$11455 ( \11832 , \11830 , \11831 );
nor \U$11456 ( \11833 , \11829 , \11832 );
nand \U$11457 ( \11834 , \11833 , \9384 );
nand \U$11458 ( \11835 , \11828 , \11834 );
not \U$11459 ( \11836 , \11179 );
not \U$11460 ( \11837 , \2710 );
or \U$11461 ( \11838 , \11836 , \11837 );
not \U$11462 ( \11839 , \11182 );
not \U$11463 ( \11840 , RIc2267a0_31);
not \U$11464 ( \11841 , \3008 );
not \U$11465 ( \11842 , \11841 );
or \U$11466 ( \11843 , \11840 , \11842 );
not \U$11467 ( \11844 , \2063 );
nand \U$11468 ( \11845 , \11844 , \3648 );
nand \U$11469 ( \11846 , \11843 , \11845 );
nand \U$11470 ( \11847 , \11839 , \11846 );
nand \U$11471 ( \11848 , \11838 , \11847 );
xor \U$11472 ( \11849 , \11835 , \11848 );
not \U$11473 ( \11850 , \3631 );
not \U$11474 ( \11851 , \11202 );
or \U$11475 ( \11852 , \11850 , \11851 );
not \U$11476 ( \11853 , RIc2266b0_33);
not \U$11477 ( \11854 , \2498 );
not \U$11478 ( \11855 , \11854 );
or \U$11479 ( \11856 , \11853 , \11855 );
nand \U$11480 ( \11857 , \4196 , \6890 );
nand \U$11481 ( \11858 , \11856 , \11857 );
nand \U$11482 ( \11859 , \11858 , \3629 );
nand \U$11483 ( \11860 , \11852 , \11859 );
and \U$11484 ( \11861 , \11849 , \11860 );
and \U$11485 ( \11862 , \11835 , \11848 );
or \U$11486 ( \11863 , \11861 , \11862 );
and \U$11487 ( \11864 , \11824 , \11863 );
and \U$11488 ( \11865 , \11788 , \11823 );
or \U$11489 ( \11866 , \11864 , \11865 );
and \U$11490 ( \11867 , \11755 , \11866 );
and \U$11491 ( \11868 , \11752 , \11754 );
or \U$11492 ( \11869 , \11867 , \11868 );
xnor \U$11493 ( \11870 , \9180 , \9178 );
buf \U$11494 ( \11871 , \9334 );
xor \U$11495 ( \11872 , \11870 , \11871 );
not \U$11496 ( \11873 , \11872 );
or \U$11497 ( \11874 , \11869 , \11873 );
not \U$11498 ( \11875 , \6307 );
not \U$11499 ( \11876 , \11650 );
or \U$11500 ( \11877 , \11875 , \11876 );
not \U$11501 ( \11878 , RIc2263e0_39);
not \U$11502 ( \11879 , \4009 );
or \U$11503 ( \11880 , \11878 , \11879 );
nand \U$11504 ( \11881 , \9608 , \5498 );
nand \U$11505 ( \11882 , \11880 , \11881 );
nand \U$11506 ( \11883 , \11882 , \6689 );
nand \U$11507 ( \11884 , \11877 , \11883 );
not \U$11508 ( \11885 , \11884 );
not \U$11509 ( \11886 , \5519 );
not \U$11510 ( \11887 , \11625 );
or \U$11511 ( \11888 , \11886 , \11887 );
not \U$11512 ( \11889 , RIc2264d0_37);
not \U$11513 ( \11890 , \2013 );
not \U$11514 ( \11891 , \11890 );
or \U$11515 ( \11892 , \11889 , \11891 );
nand \U$11516 ( \11893 , \2013 , \4371 );
nand \U$11517 ( \11894 , \11892 , \11893 );
nand \U$11518 ( \11895 , \11894 , \5509 );
nand \U$11519 ( \11896 , \11888 , \11895 );
not \U$11520 ( \11897 , \11896 );
or \U$11521 ( \11898 , \11885 , \11897 );
not \U$11522 ( \11899 , \11896 );
not \U$11523 ( \11900 , \11899 );
not \U$11524 ( \11901 , \11884 );
not \U$11525 ( \11902 , \11901 );
or \U$11526 ( \11903 , \11900 , \11902 );
not \U$11527 ( \11904 , \9552 );
not \U$11528 ( \11905 , \11638 );
or \U$11529 ( \11906 , \11904 , \11905 );
xor \U$11530 ( \11907 , RIc225f30_49, \1391 );
nand \U$11531 ( \11908 , \11907 , \9534 );
nand \U$11532 ( \11909 , \11906 , \11908 );
nand \U$11533 ( \11910 , \11903 , \11909 );
nand \U$11534 ( \11911 , \11898 , \11910 );
not \U$11535 ( \11912 , \11911 );
not \U$11536 ( \11913 , \11190 );
not \U$11537 ( \11914 , \11204 );
or \U$11538 ( \11915 , \11913 , \11914 );
or \U$11539 ( \11916 , \11190 , \11204 );
nand \U$11540 ( \11917 , \11915 , \11916 );
and \U$11541 ( \11918 , \11917 , \11186 );
not \U$11542 ( \11919 , \11917 );
and \U$11543 ( \11920 , \11919 , \11187 );
nor \U$11544 ( \11921 , \11918 , \11920 );
nand \U$11545 ( \11922 , \11912 , \11921 );
xor \U$11546 ( \11923 , \11611 , \11590 );
xnor \U$11547 ( \11924 , \11923 , \11600 );
and \U$11548 ( \11925 , \11922 , \11924 );
not \U$11549 ( \11926 , \11911 );
nor \U$11550 ( \11927 , \11921 , \11926 );
nor \U$11551 ( \11928 , \11925 , \11927 );
not \U$11552 ( \11929 , \11928 );
not \U$11553 ( \11930 , \11929 );
xor \U$11554 ( \11931 , \11629 , \11640 );
xor \U$11555 ( \11932 , \11931 , \11652 );
xor \U$11556 ( \11933 , \11707 , \11719 );
xor \U$11557 ( \11934 , \11933 , \11730 );
or \U$11558 ( \11935 , \11932 , \11934 );
xor \U$11559 ( \11936 , \11667 , \11678 );
and \U$11560 ( \11937 , \11936 , \11691 );
not \U$11561 ( \11938 , \11936 );
not \U$11562 ( \11939 , \11691 );
and \U$11563 ( \11940 , \11938 , \11939 );
nor \U$11564 ( \11941 , \11937 , \11940 );
and \U$11565 ( \11942 , \11935 , \11941 );
and \U$11566 ( \11943 , \11934 , \11932 );
nor \U$11567 ( \11944 , \11942 , \11943 );
not \U$11568 ( \11945 , \11944 );
not \U$11569 ( \11946 , \11945 );
or \U$11570 ( \11947 , \11930 , \11946 );
not \U$11571 ( \11948 , \11944 );
not \U$11572 ( \11949 , \11928 );
or \U$11573 ( \11950 , \11948 , \11949 );
xor \U$11574 ( \11951 , \11218 , \11215 );
xor \U$11575 ( \11952 , \11951 , \11206 );
not \U$11576 ( \11953 , \11952 );
nand \U$11577 ( \11954 , \11950 , \11953 );
nand \U$11578 ( \11955 , \11947 , \11954 );
nand \U$11579 ( \11956 , \11874 , \11955 );
not \U$11580 ( \11957 , \11872 );
nand \U$11581 ( \11958 , \11957 , \11869 );
and \U$11582 ( \11959 , \11956 , \11958 );
not \U$11583 ( \11960 , \11959 );
not \U$11584 ( \11961 , \11960 );
or \U$11585 ( \11962 , \11750 , \11961 );
xor \U$11586 ( \11963 , \11160 , \11162 );
xor \U$11587 ( \11964 , \11963 , \11221 );
buf \U$11588 ( \11965 , \10077 );
not \U$11589 ( \11966 , \11965 );
not \U$11590 ( \11967 , \11033 );
not \U$11591 ( \11968 , \930 );
or \U$11592 ( \11969 , \11967 , \11968 );
nand \U$11593 ( \11970 , \11112 , RIc225b70_57);
nand \U$11594 ( \11971 , \11969 , \11970 );
not \U$11595 ( \11972 , \11971 );
or \U$11596 ( \11973 , \11966 , \11972 );
buf \U$11597 ( \11974 , \10072 );
nand \U$11598 ( \11975 , \11974 , RIc225b70_57);
nand \U$11599 ( \11976 , \11973 , \11975 );
not \U$11600 ( \11977 , \1339 );
not \U$11601 ( \11978 , \11557 );
or \U$11602 ( \11979 , \11977 , \11978 );
not \U$11603 ( \11980 , RIc2271f0_9);
not \U$11604 ( \11981 , \9215 );
or \U$11605 ( \11982 , \11980 , \11981 );
nand \U$11606 ( \11983 , \8924 , \1351 );
nand \U$11607 ( \11984 , \11982 , \11983 );
nand \U$11608 ( \11985 , \11984 , \1363 );
nand \U$11609 ( \11986 , \11979 , \11985 );
xor \U$11610 ( \11987 , \11976 , \11986 );
not \U$11611 ( \11988 , \1311 );
not \U$11612 ( \11989 , \11570 );
or \U$11613 ( \11990 , \11988 , \11989 );
not \U$11614 ( \11991 , RIc227100_11);
not \U$11615 ( \11992 , \11094 );
or \U$11616 ( \11993 , \11991 , \11992 );
not \U$11617 ( \11994 , \8973 );
nand \U$11618 ( \11995 , \11994 , \3351 );
nand \U$11619 ( \11996 , \11993 , \11995 );
nand \U$11620 ( \11997 , \11996 , \9904 );
nand \U$11621 ( \11998 , \11990 , \11997 );
and \U$11622 ( \11999 , \11987 , \11998 );
and \U$11623 ( \12000 , \11976 , \11986 );
or \U$11624 ( \12001 , \11999 , \12000 );
not \U$11625 ( \12002 , \12001 );
xor \U$11626 ( \12003 , \9328 , \9283 );
xnor \U$11627 ( \12004 , \12003 , \9229 );
not \U$11628 ( \12005 , \12004 );
nand \U$11629 ( \12006 , \12002 , \12005 );
not \U$11630 ( \12007 , \12006 );
not \U$11631 ( \12008 , \9205 );
not \U$11632 ( \12009 , \11665 );
or \U$11633 ( \12010 , \12008 , \12009 );
and \U$11634 ( \12011 , \2297 , \9117 );
not \U$11635 ( \12012 , \2297 );
and \U$11636 ( \12013 , \12012 , RIc226200_43);
or \U$11637 ( \12014 , \12011 , \12013 );
nand \U$11638 ( \12015 , \12014 , \9110 );
nand \U$11639 ( \12016 , \12010 , \12015 );
not \U$11640 ( \12017 , \2172 );
not \U$11641 ( \12018 , \11676 );
or \U$11642 ( \12019 , \12017 , \12018 );
not \U$11643 ( \12020 , RIc226a70_25);
not \U$11644 ( \12021 , \9674 );
or \U$11645 ( \12022 , \12020 , \12021 );
nand \U$11646 ( \12023 , \3640 , \1905 );
nand \U$11647 ( \12024 , \12022 , \12023 );
nand \U$11648 ( \12025 , \12024 , \2195 );
nand \U$11649 ( \12026 , \12019 , \12025 );
xor \U$11650 ( \12027 , \12016 , \12026 );
not \U$11651 ( \12028 , \2154 );
not \U$11652 ( \12029 , \11689 );
or \U$11653 ( \12030 , \12028 , \12029 );
not \U$11654 ( \12031 , RIc226980_27);
not \U$11655 ( \12032 , \11321 );
or \U$11656 ( \12033 , \12031 , \12032 );
nand \U$11657 ( \12034 , \3120 , \2799 );
nand \U$11658 ( \12035 , \12033 , \12034 );
nand \U$11659 ( \12036 , \12035 , \2138 );
nand \U$11660 ( \12037 , \12030 , \12036 );
and \U$11661 ( \12038 , \12027 , \12037 );
and \U$11662 ( \12039 , \12016 , \12026 );
or \U$11663 ( \12040 , \12038 , \12039 );
not \U$11664 ( \12041 , \12040 );
or \U$11665 ( \12042 , \12007 , \12041 );
nand \U$11666 ( \12043 , \12001 , \12004 );
nand \U$11667 ( \12044 , \12042 , \12043 );
not \U$11668 ( \12045 , \12044 );
not \U$11669 ( \12046 , \12045 );
not \U$11670 ( \12047 , \11733 );
not \U$11671 ( \12048 , \11694 );
or \U$11672 ( \12049 , \12047 , \12048 );
not \U$11673 ( \12050 , \11733 );
nand \U$11674 ( \12051 , \12050 , \11693 );
nand \U$11675 ( \12052 , \12049 , \12051 );
xor \U$11676 ( \12053 , \12052 , \11656 );
not \U$11677 ( \12054 , \12053 );
or \U$11678 ( \12055 , \12046 , \12054 );
xor \U$11679 ( \12056 , \10202 , \10216 );
xor \U$11680 ( \12057 , \12056 , \10235 );
xor \U$11681 ( \12058 , \11549 , \11559 );
xor \U$11682 ( \12059 , \12058 , \11572 );
xor \U$11683 ( \12060 , \12057 , \12059 );
xor \U$11684 ( \12061 , \10137 , \10176 );
xor \U$11685 ( \12062 , \12061 , \10155 );
and \U$11686 ( \12063 , \12060 , \12062 );
and \U$11687 ( \12064 , \12057 , \12059 );
or \U$11688 ( \12065 , \12063 , \12064 );
nand \U$11689 ( \12066 , \12055 , \12065 );
not \U$11690 ( \12067 , \12053 );
nand \U$11691 ( \12068 , \12067 , \12044 );
nand \U$11692 ( \12069 , \12066 , \12068 );
xor \U$11693 ( \12070 , \11964 , \12069 );
xor \U$11694 ( \12071 , \11618 , \11736 );
xor \U$11695 ( \12072 , \12071 , \11740 );
and \U$11696 ( \12073 , \12070 , \12072 );
and \U$11697 ( \12074 , \11964 , \12069 );
or \U$11698 ( \12075 , \12073 , \12074 );
nand \U$11699 ( \12076 , \11959 , \11748 );
nand \U$11700 ( \12077 , \12075 , \12076 );
nand \U$11701 ( \12078 , \11962 , \12077 );
xor \U$11702 ( \12079 , \11746 , \12078 );
xor \U$11703 ( \12080 , \11473 , \11522 );
xor \U$11704 ( \12081 , \12080 , \11531 );
not \U$11705 ( \12082 , \12081 );
xor \U$11706 ( \12083 , \10254 , \10257 );
xnor \U$11707 ( \12084 , \12083 , \10403 );
not \U$11708 ( \12085 , \12084 );
or \U$11709 ( \12086 , \12082 , \12085 );
or \U$11710 ( \12087 , \12084 , \12081 );
xor \U$11711 ( \12088 , \11506 , \11508 );
xor \U$11712 ( \12089 , \12088 , \11519 );
not \U$11713 ( \12090 , \854 );
xor \U$11714 ( \12091 , RIc2275b0_1, \10356 );
not \U$11715 ( \12092 , \12091 );
or \U$11716 ( \12093 , \12090 , \12092 );
nand \U$11717 ( \12094 , \10372 , \1579 );
nand \U$11718 ( \12095 , \12093 , \12094 );
not \U$11719 ( \12096 , \1082 );
not \U$11720 ( \12097 , \10268 );
or \U$11721 ( \12098 , \12096 , \12097 );
not \U$11722 ( \12099 , RIc2274c0_3);
not \U$11723 ( \12100 , \9320 );
not \U$11724 ( \12101 , \12100 );
or \U$11725 ( \12102 , \12099 , \12101 );
nand \U$11726 ( \12103 , \9324 , \1032 );
nand \U$11727 ( \12104 , \12102 , \12103 );
nand \U$11728 ( \12105 , \12104 , \1040 );
nand \U$11729 ( \12106 , \12098 , \12105 );
xor \U$11730 ( \12107 , \12095 , \12106 );
not \U$11731 ( \12108 , \1118 );
not \U$11732 ( \12109 , RIc2272e0_7);
not \U$11733 ( \12110 , \10814 );
or \U$11734 ( \12111 , \12109 , \12110 );
nand \U$11735 ( \12112 , \10110 , \1139 );
nand \U$11736 ( \12113 , \12111 , \12112 );
not \U$11737 ( \12114 , \12113 );
or \U$11738 ( \12115 , \12108 , \12114 );
nand \U$11739 ( \12116 , \11482 , \1121 );
nand \U$11740 ( \12117 , \12115 , \12116 );
and \U$11741 ( \12118 , \12107 , \12117 );
and \U$11742 ( \12119 , \12095 , \12106 );
or \U$11743 ( \12120 , \12118 , \12119 );
not \U$11744 ( \12121 , \9142 );
not \U$11745 ( \12122 , \11517 );
or \U$11746 ( \12123 , \12121 , \12122 );
and \U$11747 ( \12124 , RIc226890_29, \2635 );
not \U$11748 ( \12125 , RIc226890_29);
and \U$11749 ( \12126 , \12125 , \2634 );
or \U$11750 ( \12127 , \12124 , \12126 );
nand \U$11751 ( \12128 , \12127 , \2784 );
nand \U$11752 ( \12129 , \12123 , \12128 );
xor \U$11753 ( \12130 , \12120 , \12129 );
not \U$11754 ( \12131 , \950 );
not \U$11755 ( \12132 , RIc2273d0_5);
not \U$11756 ( \12133 , \10800 );
or \U$11757 ( \12134 , \12132 , \12133 );
nand \U$11758 ( \12135 , \9274 , \946 );
nand \U$11759 ( \12136 , \12134 , \12135 );
not \U$11760 ( \12137 , \12136 );
or \U$11761 ( \12138 , \12131 , \12137 );
nand \U$11762 ( \12139 , \11492 , \954 );
nand \U$11763 ( \12140 , \12138 , \12139 );
not \U$11764 ( \12141 , \1339 );
not \U$11765 ( \12142 , \11984 );
or \U$11766 ( \12143 , \12141 , \12142 );
not \U$11767 ( \12144 , RIc2271f0_9);
not \U$11768 ( \12145 , \10645 );
or \U$11769 ( \12146 , \12144 , \12145 );
nand \U$11770 ( \12147 , \9225 , \1351 );
nand \U$11771 ( \12148 , \12146 , \12147 );
nand \U$11772 ( \12149 , \12148 , \1363 );
nand \U$11773 ( \12150 , \12143 , \12149 );
xor \U$11774 ( \12151 , \12140 , \12150 );
not \U$11775 ( \12152 , \2172 );
not \U$11776 ( \12153 , \12024 );
or \U$11777 ( \12154 , \12152 , \12153 );
and \U$11778 ( \12155 , RIc226a70_25, \4121 );
not \U$11779 ( \12156 , RIc226a70_25);
and \U$11780 ( \12157 , \12156 , \4414 );
nor \U$11781 ( \12158 , \12155 , \12157 );
nand \U$11782 ( \12159 , \12158 , \2860 );
nand \U$11783 ( \12160 , \12154 , \12159 );
and \U$11784 ( \12161 , \12151 , \12160 );
and \U$11785 ( \12162 , \12140 , \12150 );
or \U$11786 ( \12163 , \12161 , \12162 );
and \U$11787 ( \12164 , \12130 , \12163 );
and \U$11788 ( \12165 , \12120 , \12129 );
or \U$11789 ( \12166 , \12164 , \12165 );
xor \U$11790 ( \12167 , \12089 , \12166 );
xor \U$11791 ( \12168 , \10201 , \10270 );
xor \U$11792 ( \12169 , \12168 , \10281 );
not \U$11793 ( \12170 , \12169 );
not \U$11794 ( \12171 , \1930 );
not \U$11795 ( \12172 , \10279 );
or \U$11796 ( \12173 , \12171 , \12172 );
and \U$11797 ( \12174 , RIc226b60_23, \5215 );
not \U$11798 ( \12175 , RIc226b60_23);
and \U$11799 ( \12176 , \12175 , \9850 );
nor \U$11800 ( \12177 , \12174 , \12176 );
nand \U$11801 ( \12178 , \12177 , \10214 );
nand \U$11802 ( \12179 , \12173 , \12178 );
not \U$11803 ( \12180 , \12179 );
and \U$11804 ( \12181 , \10395 , \2367 );
not \U$11805 ( \12182 , \2391 );
xor \U$11806 ( \12183 , \2370 , \6070 );
nor \U$11807 ( \12184 , \12182 , \12183 );
nor \U$11808 ( \12185 , \12181 , \12184 );
not \U$11809 ( \12186 , \12185 );
not \U$11810 ( \12187 , \12186 );
or \U$11811 ( \12188 , \12180 , \12187 );
not \U$11812 ( \12189 , \12185 );
not \U$11813 ( \12190 , \12179 );
not \U$11814 ( \12191 , \12190 );
or \U$11815 ( \12192 , \12189 , \12191 );
not \U$11816 ( \12193 , \2518 );
and \U$11817 ( \12194 , \6718 , \1941 );
not \U$11818 ( \12195 , \6718 );
and \U$11819 ( \12196 , \12195 , RIc226d40_19);
or \U$11820 ( \12197 , \12194 , \12196 );
not \U$11821 ( \12198 , \12197 );
or \U$11822 ( \12199 , \12193 , \12198 );
nand \U$11823 ( \12200 , \10385 , \2534 );
nand \U$11824 ( \12201 , \12199 , \12200 );
nand \U$11825 ( \12202 , \12192 , \12201 );
nand \U$11826 ( \12203 , \12188 , \12202 );
not \U$11827 ( \12204 , \12203 );
nand \U$11828 ( \12205 , \12170 , \12204 );
not \U$11829 ( \12206 , \12205 );
not \U$11830 ( \12207 , \2358 );
not \U$11831 ( \12208 , \10326 );
or \U$11832 ( \12209 , \12207 , \12208 );
not \U$11833 ( \12210 , RIc226f20_15);
not \U$11834 ( \12211 , \9900 );
or \U$11835 ( \12212 , \12210 , \12211 );
nand \U$11836 ( \12213 , \8829 , \1674 );
nand \U$11837 ( \12214 , \12212 , \12213 );
nand \U$11838 ( \12215 , \12214 , \2320 );
nand \U$11839 ( \12216 , \12209 , \12215 );
not \U$11840 ( \12217 , \1682 );
not \U$11841 ( \12218 , \10299 );
or \U$11842 ( \12219 , \12217 , \12218 );
xor \U$11843 ( \12220 , RIc227010_13, \8951 );
nand \U$11844 ( \12221 , \12220 , \3250 );
nand \U$11845 ( \12222 , \12219 , \12221 );
or \U$11846 ( \12223 , \12216 , \12222 );
not \U$11847 ( \12224 , \1963 );
not \U$11848 ( \12225 , \10312 );
or \U$11849 ( \12226 , \12224 , \12225 );
not \U$11850 ( \12227 , RIc226e30_17);
not \U$11851 ( \12228 , \8885 );
not \U$11852 ( \12229 , \12228 );
or \U$11853 ( \12230 , \12227 , \12229 );
nand \U$11854 ( \12231 , \8885 , \1952 );
nand \U$11855 ( \12232 , \12230 , \12231 );
nand \U$11856 ( \12233 , \12232 , \1945 );
nand \U$11857 ( \12234 , \12226 , \12233 );
nand \U$11858 ( \12235 , \12223 , \12234 );
nand \U$11859 ( \12236 , \12216 , \12222 );
nand \U$11860 ( \12237 , \12235 , \12236 );
not \U$11861 ( \12238 , \12237 );
or \U$11862 ( \12239 , \12206 , \12238 );
not \U$11863 ( \12240 , \12204 );
nand \U$11864 ( \12241 , \12240 , \12169 );
nand \U$11865 ( \12242 , \12239 , \12241 );
and \U$11866 ( \12243 , \12167 , \12242 );
and \U$11867 ( \12244 , \12089 , \12166 );
or \U$11868 ( \12245 , \12243 , \12244 );
nand \U$11869 ( \12246 , \12087 , \12245 );
nand \U$11870 ( \12247 , \12086 , \12246 );
not \U$11871 ( \12248 , \12247 );
and \U$11872 ( \12249 , \11465 , \11451 );
not \U$11873 ( \12250 , \11465 );
and \U$11874 ( \12251 , \12250 , \11452 );
nor \U$11875 ( \12252 , \12249 , \12251 );
xor \U$11876 ( \12253 , \12252 , \11534 );
not \U$11877 ( \12254 , \12253 );
or \U$11878 ( \12255 , \12248 , \12254 );
or \U$11879 ( \12256 , \12247 , \12253 );
xor \U$11880 ( \12257 , \10406 , \10242 );
xnor \U$11881 ( \12258 , \12257 , \10061 );
nand \U$11882 ( \12259 , \12256 , \12258 );
nand \U$11883 ( \12260 , \12255 , \12259 );
not \U$11884 ( \12261 , \12260 );
and \U$11885 ( \12262 , \11536 , \11447 );
not \U$11886 ( \12263 , \11536 );
and \U$11887 ( \12264 , \12263 , \11448 );
or \U$11888 ( \12265 , \12262 , \12264 );
buf \U$11889 ( \12266 , \11743 );
and \U$11890 ( \12267 , \12265 , \12266 );
not \U$11891 ( \12268 , \12265 );
not \U$11892 ( \12269 , \12266 );
and \U$11893 ( \12270 , \12268 , \12269 );
nor \U$11894 ( \12271 , \12267 , \12270 );
not \U$11895 ( \12272 , \12271 );
or \U$11896 ( \12273 , \12261 , \12272 );
or \U$11897 ( \12274 , \12271 , \12260 );
xor \U$11898 ( \12275 , \10054 , \10409 );
xor \U$11899 ( \12276 , \12275 , \10548 );
nand \U$11900 ( \12277 , \12274 , \12276 );
nand \U$11901 ( \12278 , \12273 , \12277 );
xnor \U$11902 ( \12279 , \12079 , \12278 );
xor \U$11903 ( \12280 , \11032 , \12279 );
and \U$11904 ( \12281 , \11458 , \11462 );
not \U$11905 ( \12282 , \11458 );
and \U$11906 ( \12283 , \12282 , \11461 );
or \U$11907 ( \12284 , \12281 , \12283 );
buf \U$11908 ( \12285 , \11456 );
not \U$11909 ( \12286 , \12285 );
and \U$11910 ( \12287 , \12284 , \12286 );
not \U$11911 ( \12288 , \12284 );
and \U$11912 ( \12289 , \12288 , \12285 );
nor \U$11913 ( \12290 , \12287 , \12289 );
xor \U$11914 ( \12291 , \10284 , \10330 );
xor \U$11915 ( \12292 , \12291 , \10400 );
xor \U$11916 ( \12293 , \10344 , \10357 );
xor \U$11917 ( \12294 , \12293 , \10374 );
not \U$11918 ( \12295 , \9641 );
not \U$11919 ( \12296 , RIc226020_47);
not \U$11920 ( \12297 , \3783 );
or \U$11921 ( \12298 , \12296 , \12297 );
not \U$11922 ( \12299 , \10677 );
nand \U$11923 ( \12300 , \12299 , \11607 );
nand \U$11924 ( \12301 , \12298 , \12300 );
not \U$11925 ( \12302 , \12301 );
or \U$11926 ( \12303 , \12295 , \12302 );
buf \U$11927 ( \12304 , \9619 );
nand \U$11928 ( \12305 , \11771 , \12304 );
nand \U$11929 ( \12306 , \12303 , \12305 );
xor \U$11930 ( \12307 , \12294 , \12306 );
not \U$11931 ( \12308 , \2697 );
not \U$11932 ( \12309 , RIc2267a0_31);
not \U$11933 ( \12310 , \11515 );
not \U$11934 ( \12311 , \12310 );
or \U$11935 ( \12312 , \12309 , \12311 );
nand \U$11936 ( \12313 , \11515 , \9159 );
nand \U$11937 ( \12314 , \12312 , \12313 );
not \U$11938 ( \12315 , \12314 );
or \U$11939 ( \12316 , \12308 , \12315 );
nand \U$11940 ( \12317 , \11846 , \3653 );
nand \U$11941 ( \12318 , \12316 , \12317 );
and \U$11942 ( \12319 , \12307 , \12318 );
and \U$11943 ( \12320 , \12294 , \12306 );
or \U$11944 ( \12321 , \12319 , \12320 );
not \U$11945 ( \12322 , \12321 );
xor \U$11946 ( \12323 , \11976 , \11986 );
xor \U$11947 ( \12324 , \12323 , \11998 );
not \U$11948 ( \12325 , \12324 );
xor \U$11949 ( \12326 , \10301 , \10328 );
not \U$11950 ( \12327 , \10314 );
and \U$11951 ( \12328 , \12326 , \12327 );
not \U$11952 ( \12329 , \12326 );
and \U$11953 ( \12330 , \12329 , \10314 );
nor \U$11954 ( \12331 , \12328 , \12330 );
nand \U$11955 ( \12332 , \12325 , \12331 );
not \U$11956 ( \12333 , \12332 );
or \U$11957 ( \12334 , \12322 , \12333 );
not \U$11958 ( \12335 , \12331 );
nand \U$11959 ( \12336 , \12335 , \12324 );
nand \U$11960 ( \12337 , \12334 , \12336 );
xor \U$11961 ( \12338 , \12292 , \12337 );
and \U$11962 ( \12339 , \12001 , \12004 );
not \U$11963 ( \12340 , \12001 );
and \U$11964 ( \12341 , \12340 , \12005 );
nor \U$11965 ( \12342 , \12339 , \12341 );
xor \U$11966 ( \12343 , \12040 , \12342 );
and \U$11967 ( \12344 , \12338 , \12343 );
and \U$11968 ( \12345 , \12292 , \12337 );
or \U$11969 ( \12346 , \12344 , \12345 );
xor \U$11970 ( \12347 , \12290 , \12346 );
xor \U$11971 ( \12348 , \12057 , \12059 );
xor \U$11972 ( \12349 , \12348 , \12062 );
xor \U$11973 ( \12350 , \10377 , \10387 );
xor \U$11974 ( \12351 , \12350 , \10397 );
xor \U$11975 ( \12352 , \11835 , \11848 );
xor \U$11976 ( \12353 , \12352 , \11860 );
xor \U$11977 ( \12354 , \12351 , \12353 );
xor \U$11978 ( \12355 , \11799 , \11809 );
xor \U$11979 ( \12356 , \12355 , \11820 );
and \U$11980 ( \12357 , \12354 , \12356 );
and \U$11981 ( \12358 , \12351 , \12353 );
or \U$11982 ( \12359 , \12357 , \12358 );
xor \U$11983 ( \12360 , \12349 , \12359 );
xor \U$11984 ( \12361 , \11788 , \11823 );
xor \U$11985 ( \12362 , \12361 , \11863 );
and \U$11986 ( \12363 , \12360 , \12362 );
and \U$11987 ( \12364 , \12349 , \12359 );
or \U$11988 ( \12365 , \12363 , \12364 );
and \U$11989 ( \12366 , \12347 , \12365 );
and \U$11990 ( \12367 , \12290 , \12346 );
or \U$11991 ( \12368 , \12366 , \12367 );
not \U$11992 ( \12369 , \12065 );
not \U$11993 ( \12370 , \12045 );
or \U$11994 ( \12371 , \12369 , \12370 );
not \U$11995 ( \12372 , \12065 );
nand \U$11996 ( \12373 , \12372 , \12044 );
nand \U$11997 ( \12374 , \12371 , \12373 );
xor \U$11998 ( \12375 , \12374 , \12053 );
not \U$11999 ( \12376 , \12375 );
not \U$12000 ( \12377 , \12376 );
xor \U$12001 ( \12378 , \11496 , \11504 );
xor \U$12002 ( \12379 , \12378 , \11484 );
not \U$12003 ( \12380 , \9934 );
not \U$12004 ( \12381 , RIc226110_45);
not \U$12005 ( \12382 , \2353 );
not \U$12006 ( \12383 , \12382 );
or \U$12007 ( \12384 , \12381 , \12383 );
nand \U$12008 ( \12385 , \2353 , \10429 );
nand \U$12009 ( \12386 , \12384 , \12385 );
not \U$12010 ( \12387 , \12386 );
or \U$12011 ( \12388 , \12380 , \12387 );
nand \U$12012 ( \12389 , \11833 , \9398 );
nand \U$12013 ( \12390 , \12388 , \12389 );
not \U$12014 ( \12391 , \2784 );
and \U$12015 ( \12392 , RIc226890_29, \3715 );
not \U$12016 ( \12393 , RIc226890_29);
and \U$12017 ( \12394 , \12393 , \3716 );
or \U$12018 ( \12395 , \12392 , \12394 );
not \U$12019 ( \12396 , \12395 );
or \U$12020 ( \12397 , \12391 , \12396 );
nand \U$12021 ( \12398 , \12127 , \2086 );
nand \U$12022 ( \12399 , \12397 , \12398 );
or \U$12023 ( \12400 , \12390 , \12399 );
not \U$12024 ( \12401 , \9904 );
not \U$12025 ( \12402 , RIc227100_11);
not \U$12026 ( \12403 , \8913 );
not \U$12027 ( \12404 , \12403 );
or \U$12028 ( \12405 , \12402 , \12404 );
buf \U$12029 ( \12406 , \8913 );
nand \U$12030 ( \12407 , \12406 , \1685 );
nand \U$12031 ( \12408 , \12405 , \12407 );
not \U$12032 ( \12409 , \12408 );
or \U$12033 ( \12410 , \12401 , \12409 );
nand \U$12034 ( \12411 , \11996 , \1311 );
nand \U$12035 ( \12412 , \12410 , \12411 );
nand \U$12036 ( \12413 , \12400 , \12412 );
nand \U$12037 ( \12414 , \12399 , \12390 );
nand \U$12038 ( \12415 , \12413 , \12414 );
xor \U$12039 ( \12416 , \12379 , \12415 );
not \U$12040 ( \12417 , \9444 );
not \U$12041 ( \12418 , \11797 );
or \U$12042 ( \12419 , \12417 , \12418 );
not \U$12043 ( \12420 , RIc225e40_51);
not \U$12044 ( \12421 , \1438 );
or \U$12045 ( \12422 , \12420 , \12421 );
not \U$12046 ( \12423 , RIc225e40_51);
nand \U$12047 ( \12424 , \1370 , \12423 );
nand \U$12048 ( \12425 , \12422 , \12424 );
nand \U$12049 ( \12426 , \12425 , \9459 );
nand \U$12050 ( \12427 , \12419 , \12426 );
not \U$12051 ( \12428 , \9488 );
not \U$12052 ( \12429 , RIc225d50_53);
not \U$12053 ( \12430 , \2118 );
or \U$12054 ( \12431 , \12429 , \12430 );
nand \U$12055 ( \12432 , \1020 , \11585 );
nand \U$12056 ( \12433 , \12431 , \12432 );
not \U$12057 ( \12434 , \12433 );
or \U$12058 ( \12435 , \12428 , \12434 );
nand \U$12059 ( \12436 , \11783 , \11577 );
nand \U$12060 ( \12437 , \12435 , \12436 );
xor \U$12061 ( \12438 , \12427 , \12437 );
not \U$12062 ( \12439 , \9816 );
not \U$12063 ( \12440 , \11818 );
or \U$12064 ( \12441 , \12439 , \12440 );
not \U$12065 ( \12442 , RIc2262f0_41);
not \U$12066 ( \12443 , \2226 );
or \U$12067 ( \12444 , \12442 , \12443 );
nand \U$12068 ( \12445 , \2225 , \6303 );
nand \U$12069 ( \12446 , \12444 , \12445 );
nand \U$12070 ( \12447 , \12446 , \9690 );
nand \U$12071 ( \12448 , \12441 , \12447 );
and \U$12072 ( \12449 , \12438 , \12448 );
and \U$12073 ( \12450 , \12427 , \12437 );
or \U$12074 ( \12451 , \12449 , \12450 );
and \U$12075 ( \12452 , \12416 , \12451 );
and \U$12076 ( \12453 , \12379 , \12415 );
or \U$12077 ( \12454 , \12452 , \12453 );
not \U$12078 ( \12455 , \9110 );
not \U$12079 ( \12456 , RIc226200_43);
and \U$12080 ( \12457 , \2421 , \12456 );
not \U$12081 ( \12458 , \2421 );
and \U$12082 ( \12459 , \12458 , RIc226200_43);
or \U$12083 ( \12460 , \12457 , \12459 );
not \U$12084 ( \12461 , \12460 );
or \U$12085 ( \12462 , \12455 , \12461 );
nand \U$12086 ( \12463 , \12014 , \9129 );
nand \U$12087 ( \12464 , \12462 , \12463 );
not \U$12088 ( \12465 , \12464 );
not \U$12089 ( \12466 , \11971 );
not \U$12090 ( \12467 , \12466 );
not \U$12091 ( \12468 , \11974 );
not \U$12092 ( \12469 , \12468 );
and \U$12093 ( \12470 , \12467 , \12469 );
not \U$12094 ( \12471 , RIc225b70_57);
not \U$12095 ( \12472 , \1072 );
not \U$12096 ( \12473 , \12472 );
or \U$12097 ( \12474 , \12471 , \12473 );
not \U$12098 ( \12475 , RIc225b70_57);
nand \U$12099 ( \12476 , \1072 , \12475 );
nand \U$12100 ( \12477 , \12474 , \12476 );
and \U$12101 ( \12478 , \12477 , \11965 );
nor \U$12102 ( \12479 , \12470 , \12478 );
not \U$12103 ( \12480 , \12479 );
not \U$12104 ( \12481 , \12480 );
or \U$12105 ( \12482 , \12465 , \12481 );
not \U$12106 ( \12483 , \9110 );
not \U$12107 ( \12484 , \12460 );
or \U$12108 ( \12485 , \12483 , \12484 );
nand \U$12109 ( \12486 , \12485 , \12463 );
not \U$12110 ( \12487 , \12486 );
not \U$12111 ( \12488 , \12487 );
not \U$12112 ( \12489 , \12479 );
or \U$12113 ( \12490 , \12488 , \12489 );
not \U$12114 ( \12491 , \2138 );
not \U$12115 ( \12492 , RIc226980_27);
not \U$12116 ( \12493 , \2980 );
not \U$12117 ( \12494 , \12493 );
or \U$12118 ( \12495 , \12492 , \12494 );
nand \U$12119 ( \12496 , \3725 , \4528 );
nand \U$12120 ( \12497 , \12495 , \12496 );
not \U$12121 ( \12498 , \12497 );
or \U$12122 ( \12499 , \12491 , \12498 );
nand \U$12123 ( \12500 , \12035 , \2154 );
nand \U$12124 ( \12501 , \12499 , \12500 );
nand \U$12125 ( \12502 , \12490 , \12501 );
nand \U$12126 ( \12503 , \12482 , \12502 );
not \U$12127 ( \12504 , \6688 );
not \U$12128 ( \12505 , RIc2263e0_39);
not \U$12129 ( \12506 , \1989 );
or \U$12130 ( \12507 , \12505 , \12506 );
not \U$12131 ( \12508 , \1988 );
not \U$12132 ( \12509 , \12508 );
nand \U$12133 ( \12510 , \12509 , \6694 );
nand \U$12134 ( \12511 , \12507 , \12510 );
not \U$12135 ( \12512 , \12511 );
or \U$12136 ( \12513 , \12504 , \12512 );
nand \U$12137 ( \12514 , \11882 , \6307 );
nand \U$12138 ( \12515 , \12513 , \12514 );
not \U$12139 ( \12516 , \12515 );
not \U$12140 ( \12517 , \5509 );
not \U$12141 ( \12518 , RIc2264d0_37);
not \U$12142 ( \12519 , \2590 );
not \U$12143 ( \12520 , \12519 );
or \U$12144 ( \12521 , \12518 , \12520 );
not \U$12145 ( \12522 , RIc2264d0_37);
nand \U$12146 ( \12523 , \2590 , \12522 );
nand \U$12147 ( \12524 , \12521 , \12523 );
not \U$12148 ( \12525 , \12524 );
or \U$12149 ( \12526 , \12517 , \12525 );
nand \U$12150 ( \12527 , \11894 , \5519 );
nand \U$12151 ( \12528 , \12526 , \12527 );
not \U$12152 ( \12529 , \12528 );
or \U$12153 ( \12530 , \12516 , \12529 );
or \U$12154 ( \12531 , \12528 , \12515 );
buf \U$12155 ( \12532 , \11038 );
not \U$12156 ( \12533 , \12532 );
not \U$12157 ( \12534 , \11805 );
or \U$12158 ( \12535 , \12533 , \12534 );
not \U$12159 ( \12536 , RIc225c60_55);
not \U$12160 ( \12537 , \839 );
not \U$12161 ( \12538 , \12537 );
or \U$12162 ( \12539 , \12536 , \12538 );
nand \U$12163 ( \12540 , \840 , \11041 );
nand \U$12164 ( \12541 , \12539 , \12540 );
nand \U$12165 ( \12542 , \12541 , \11118 );
nand \U$12166 ( \12543 , \12535 , \12542 );
nand \U$12167 ( \12544 , \12531 , \12543 );
nand \U$12168 ( \12545 , \12530 , \12544 );
xor \U$12169 ( \12546 , \12503 , \12545 );
not \U$12170 ( \12547 , RIc2266b0_33);
not \U$12171 ( \12548 , \2720 );
not \U$12172 ( \12549 , \12548 );
or \U$12173 ( \12550 , \12547 , \12549 );
not \U$12174 ( \12551 , RIc2266b0_33);
nand \U$12175 ( \12552 , \2720 , \12551 );
nand \U$12176 ( \12553 , \12550 , \12552 );
not \U$12177 ( \12554 , \12553 );
not \U$12178 ( \12555 , \12554 );
not \U$12179 ( \12556 , \5185 );
and \U$12180 ( \12557 , \12555 , \12556 );
and \U$12181 ( \12558 , \11858 , \3631 );
nor \U$12182 ( \12559 , \12557 , \12558 );
not \U$12183 ( \12560 , \12559 );
not \U$12184 ( \12561 , \4383 );
not \U$12185 ( \12562 , \11763 );
or \U$12186 ( \12563 , \12561 , \12562 );
and \U$12187 ( \12564 , \2475 , \3620 );
not \U$12188 ( \12565 , \2475 );
and \U$12189 ( \12566 , \12565 , RIc2265c0_35);
or \U$12190 ( \12567 , \12564 , \12566 );
nand \U$12191 ( \12568 , \12567 , \4381 );
nand \U$12192 ( \12569 , \12563 , \12568 );
or \U$12193 ( \12570 , \12560 , \12569 );
not \U$12194 ( \12571 , \9552 );
not \U$12195 ( \12572 , \11907 );
or \U$12196 ( \12573 , \12571 , \12572 );
not \U$12197 ( \12574 , RIc225f30_49);
not \U$12198 ( \12575 , \3578 );
or \U$12199 ( \12576 , \12574 , \12575 );
not \U$12200 ( \12577 , RIc225f30_49);
nand \U$12201 ( \12578 , \12577 , \1529 );
nand \U$12202 ( \12579 , \12576 , \12578 );
nand \U$12203 ( \12580 , \12579 , \9532 );
nand \U$12204 ( \12581 , \12573 , \12580 );
nand \U$12205 ( \12582 , \12570 , \12581 );
nand \U$12206 ( \12583 , \12569 , \12560 );
nand \U$12207 ( \12584 , \12582 , \12583 );
and \U$12208 ( \12585 , \12546 , \12584 );
and \U$12209 ( \12586 , \12503 , \12545 );
or \U$12210 ( \12587 , \12585 , \12586 );
xor \U$12211 ( \12588 , \12454 , \12587 );
xor \U$12212 ( \12589 , \11785 , \11775 );
not \U$12213 ( \12590 , \11765 );
xor \U$12214 ( \12591 , \12589 , \12590 );
not \U$12215 ( \12592 , \12591 );
not \U$12216 ( \12593 , \11909 );
not \U$12217 ( \12594 , \11901 );
or \U$12218 ( \12595 , \12593 , \12594 );
not \U$12219 ( \12596 , \11909 );
nand \U$12220 ( \12597 , \12596 , \11884 );
nand \U$12221 ( \12598 , \12595 , \12597 );
and \U$12222 ( \12599 , \12598 , \11899 );
not \U$12223 ( \12600 , \12598 );
and \U$12224 ( \12601 , \12600 , \11896 );
nor \U$12225 ( \12602 , \12599 , \12601 );
not \U$12226 ( \12603 , \12602 );
or \U$12227 ( \12604 , \12592 , \12603 );
xor \U$12228 ( \12605 , \12016 , \12026 );
xor \U$12229 ( \12606 , \12605 , \12037 );
nand \U$12230 ( \12607 , \12604 , \12606 );
not \U$12231 ( \12608 , \12602 );
not \U$12232 ( \12609 , \12591 );
nand \U$12233 ( \12610 , \12608 , \12609 );
nand \U$12234 ( \12611 , \12607 , \12610 );
and \U$12235 ( \12612 , \12588 , \12611 );
and \U$12236 ( \12613 , \12454 , \12587 );
or \U$12237 ( \12614 , \12612 , \12613 );
not \U$12238 ( \12615 , \12614 );
or \U$12239 ( \12616 , \12377 , \12615 );
not \U$12240 ( \12617 , \12614 );
not \U$12241 ( \12618 , \12617 );
not \U$12242 ( \12619 , \12375 );
or \U$12243 ( \12620 , \12618 , \12619 );
xor \U$12244 ( \12621 , \11752 , \11754 );
xor \U$12245 ( \12622 , \12621 , \11866 );
nand \U$12246 ( \12623 , \12620 , \12622 );
nand \U$12247 ( \12624 , \12616 , \12623 );
xor \U$12248 ( \12625 , \12368 , \12624 );
xor \U$12249 ( \12626 , \11872 , \11869 );
xnor \U$12250 ( \12627 , \12626 , \11955 );
and \U$12251 ( \12628 , \12625 , \12627 );
and \U$12252 ( \12629 , \12368 , \12624 );
or \U$12253 ( \12630 , \12628 , \12629 );
xor \U$12254 ( \12631 , \11749 , \11960 );
xor \U$12255 ( \12632 , \12631 , \12075 );
xor \U$12256 ( \12633 , \12630 , \12632 );
xor \U$12257 ( \12634 , \11964 , \12069 );
xor \U$12258 ( \12635 , \12634 , \12072 );
and \U$12259 ( \12636 , \11928 , \11952 );
not \U$12260 ( \12637 , \11928 );
and \U$12261 ( \12638 , \12637 , \11953 );
nor \U$12262 ( \12639 , \12636 , \12638 );
and \U$12263 ( \12640 , \12639 , \11945 );
not \U$12264 ( \12641 , \12639 );
and \U$12265 ( \12642 , \12641 , \11944 );
nor \U$12266 ( \12643 , \12640 , \12642 );
not \U$12267 ( \12644 , \12643 );
xor \U$12268 ( \12645 , \12245 , \12081 );
xnor \U$12269 ( \12646 , \12645 , \12084 );
not \U$12270 ( \12647 , \12646 );
not \U$12271 ( \12648 , \12647 );
or \U$12272 ( \12649 , \12644 , \12648 );
not \U$12273 ( \12650 , \12643 );
not \U$12274 ( \12651 , \12650 );
not \U$12275 ( \12652 , \12646 );
or \U$12276 ( \12653 , \12651 , \12652 );
xor \U$12277 ( \12654 , \11911 , \11924 );
xnor \U$12278 ( \12655 , \12654 , \11921 );
xor \U$12279 ( \12656 , \11934 , \11932 );
xor \U$12280 ( \12657 , \12656 , \11941 );
or \U$12281 ( \12658 , \12655 , \12657 );
xor \U$12282 ( \12659 , \12120 , \12129 );
xor \U$12283 ( \12660 , \12659 , \12163 );
xor \U$12284 ( \12661 , \12140 , \12150 );
xor \U$12285 ( \12662 , \12661 , \12160 );
not \U$12286 ( \12663 , \12662 );
not \U$12287 ( \12664 , \12663 );
buf \U$12288 ( \12665 , \10341 );
not \U$12289 ( \12666 , \12665 );
xor \U$12290 ( \12667 , RIc225a80_59, \930 );
not \U$12291 ( \12668 , \12667 );
or \U$12292 ( \12669 , \12666 , \12668 );
buf \U$12293 ( \12670 , \10342 );
nand \U$12294 ( \12671 , \12670 , RIc225a80_59);
nand \U$12295 ( \12672 , \12669 , \12671 );
not \U$12296 ( \12673 , \12672 );
and \U$12297 ( \12674 , \12214 , \2358 );
not \U$12298 ( \12675 , RIc226f20_15);
not \U$12299 ( \12676 , \8807 );
or \U$12300 ( \12677 , \12675 , \12676 );
nand \U$12301 ( \12678 , \8806 , \2301 );
nand \U$12302 ( \12679 , \12677 , \12678 );
and \U$12303 ( \12680 , \12679 , \2320 );
nor \U$12304 ( \12681 , \12674 , \12680 );
nand \U$12305 ( \12682 , \12673 , \12681 );
not \U$12306 ( \12683 , \3250 );
and \U$12307 ( \12684 , RIc227010_13, \11094 );
not \U$12308 ( \12685 , RIc227010_13);
and \U$12309 ( \12686 , \12685 , \8979 );
or \U$12310 ( \12687 , \12684 , \12686 );
not \U$12311 ( \12688 , \12687 );
or \U$12312 ( \12689 , \12683 , \12688 );
nand \U$12313 ( \12690 , \12220 , \1682 );
nand \U$12314 ( \12691 , \12689 , \12690 );
and \U$12315 ( \12692 , \12682 , \12691 );
nor \U$12316 ( \12693 , \12673 , \12681 );
nor \U$12317 ( \12694 , \12692 , \12693 );
not \U$12318 ( \12695 , \12694 );
or \U$12319 ( \12696 , \12664 , \12695 );
not \U$12320 ( \12697 , RIc226c50_21);
not \U$12321 ( \12698 , \6492 );
not \U$12322 ( \12699 , \12698 );
or \U$12323 ( \12700 , \12697 , \12699 );
nand \U$12324 ( \12701 , \6492 , \4475 );
nand \U$12325 ( \12702 , \12700 , \12701 );
and \U$12326 ( \12703 , \12702 , \2392 );
not \U$12327 ( \12704 , \12183 );
and \U$12328 ( \12705 , \12704 , \2367 );
nor \U$12329 ( \12706 , \12703 , \12705 );
not \U$12330 ( \12707 , \12706 );
not \U$12331 ( \12708 , \2518 );
not \U$12332 ( \12709 , RIc226d40_19);
not \U$12333 ( \12710 , \10142 );
or \U$12334 ( \12711 , \12709 , \12710 );
not \U$12335 ( \12712 , \9728 );
nand \U$12336 ( \12713 , \12712 , \2523 );
nand \U$12337 ( \12714 , \12711 , \12713 );
not \U$12338 ( \12715 , \12714 );
or \U$12339 ( \12716 , \12708 , \12715 );
nand \U$12340 ( \12717 , \12197 , \2534 );
nand \U$12341 ( \12718 , \12716 , \12717 );
not \U$12342 ( \12719 , \12718 );
not \U$12343 ( \12720 , \12719 );
or \U$12344 ( \12721 , \12707 , \12720 );
not \U$12345 ( \12722 , \1945 );
not \U$12346 ( \12723 , RIc226e30_17);
not \U$12347 ( \12724 , \8856 );
not \U$12348 ( \12725 , \12724 );
or \U$12349 ( \12726 , \12723 , \12725 );
buf \U$12350 ( \12727 , \8856 );
nand \U$12351 ( \12728 , \12727 , \1935 );
nand \U$12352 ( \12729 , \12726 , \12728 );
not \U$12353 ( \12730 , \12729 );
or \U$12354 ( \12731 , \12722 , \12730 );
nand \U$12355 ( \12732 , \12232 , \1963 );
nand \U$12356 ( \12733 , \12731 , \12732 );
nand \U$12357 ( \12734 , \12721 , \12733 );
or \U$12358 ( \12735 , \12706 , \12719 );
nand \U$12359 ( \12736 , \12734 , \12735 );
nand \U$12360 ( \12737 , \12696 , \12736 );
not \U$12361 ( \12738 , \12663 );
not \U$12362 ( \12739 , \12694 );
nand \U$12363 ( \12740 , \12738 , \12739 );
nand \U$12364 ( \12741 , \12737 , \12740 );
xor \U$12365 ( \12742 , \12660 , \12741 );
not \U$12366 ( \12743 , \517 );
not \U$12367 ( \12744 , \12743 );
not \U$12368 ( \12745 , \10185 );
or \U$12369 ( \12746 , \12744 , \12745 );
nand \U$12370 ( \12747 , \12746 , \565 );
not \U$12371 ( \12748 , \567 );
nor \U$12372 ( \12749 , \12748 , \564 );
and \U$12373 ( \12750 , \12747 , \12749 );
not \U$12374 ( \12751 , \12747 );
not \U$12375 ( \12752 , \12749 );
and \U$12376 ( \12753 , \12751 , \12752 );
nor \U$12377 ( \12754 , \12750 , \12753 );
buf \U$12378 ( \12755 , \12754 );
buf \U$12379 ( \12756 , \12755 );
and \U$12380 ( \12757 , \12756 , RIc2275b0_1);
not \U$12381 ( \12758 , \12095 );
xor \U$12382 ( \12759 , \12757 , \12758 );
not \U$12383 ( \12760 , \1339 );
not \U$12384 ( \12761 , \12148 );
or \U$12385 ( \12762 , \12760 , \12761 );
not \U$12386 ( \12763 , RIc2271f0_9);
not \U$12387 ( \12764 , \9076 );
or \U$12388 ( \12765 , \12763 , \12764 );
nand \U$12389 ( \12766 , \10653 , \1351 );
nand \U$12390 ( \12767 , \12765 , \12766 );
nand \U$12391 ( \12768 , \12767 , \1363 );
nand \U$12392 ( \12769 , \12762 , \12768 );
and \U$12393 ( \12770 , \12759 , \12769 );
and \U$12394 ( \12771 , \12757 , \12758 );
or \U$12395 ( \12772 , \12770 , \12771 );
not \U$12396 ( \12773 , \12772 );
not \U$12397 ( \12774 , \12773 );
not \U$12398 ( \12775 , \12158 );
not \U$12399 ( \12776 , \12775 );
not \U$12400 ( \12777 , \2171 );
and \U$12401 ( \12778 , \12776 , \12777 );
not \U$12402 ( \12779 , RIc226a70_25);
not \U$12403 ( \12780 , \6076 );
or \U$12404 ( \12781 , \12779 , \12780 );
nand \U$12405 ( \12782 , \4406 , \1905 );
nand \U$12406 ( \12783 , \12781 , \12782 );
and \U$12407 ( \12784 , \12783 , \2195 );
nor \U$12408 ( \12785 , \12778 , \12784 );
not \U$12409 ( \12786 , \12785 );
not \U$12410 ( \12787 , \12786 );
not \U$12411 ( \12788 , RIc226b60_23);
not \U$12412 ( \12789 , \10161 );
or \U$12413 ( \12790 , \12788 , \12789 );
not \U$12414 ( \12791 , \10161 );
nand \U$12415 ( \12792 , \12791 , \5637 );
nand \U$12416 ( \12793 , \12790 , \12792 );
and \U$12417 ( \12794 , \12793 , \10214 );
and \U$12418 ( \12795 , \12177 , \1930 );
nor \U$12419 ( \12796 , \12794 , \12795 );
not \U$12420 ( \12797 , \12796 );
not \U$12421 ( \12798 , \12797 );
or \U$12422 ( \12799 , \12787 , \12798 );
not \U$12423 ( \12800 , \12796 );
not \U$12424 ( \12801 , \12785 );
or \U$12425 ( \12802 , \12800 , \12801 );
xor \U$12426 ( \12803 , RIc225918_62, RIc2258a0_63);
not \U$12427 ( \12804 , \12803 );
not \U$12428 ( \12805 , \12804 );
not \U$12429 ( \12806 , RIc225990_61);
and \U$12430 ( \12807 , RIc225918_62, \12806 );
not \U$12431 ( \12808 , RIc225918_62);
and \U$12432 ( \12809 , \12808 , RIc225990_61);
nor \U$12433 ( \12810 , \12807 , \12809 );
nor \U$12434 ( \12811 , \12810 , \12803 );
not \U$12435 ( \12812 , \12811 );
not \U$12436 ( \12813 , \12812 );
or \U$12437 ( \12814 , \12805 , \12813 );
nand \U$12438 ( \12815 , \12814 , RIc225990_61);
not \U$12439 ( \12816 , \565 );
nor \U$12440 ( \12817 , \12816 , \517 );
not \U$12441 ( \12818 , \12817 );
not \U$12442 ( \12819 , \10185 );
not \U$12443 ( \12820 , \12819 );
or \U$12444 ( \12821 , \12818 , \12820 );
not \U$12445 ( \12822 , \12817 );
nand \U$12446 ( \12823 , \12822 , \10185 );
nand \U$12447 ( \12824 , \12821 , \12823 );
buf \U$12448 ( \12825 , \12824 );
and \U$12449 ( \12826 , \12825 , RIc2275b0_1);
xor \U$12450 ( \12827 , \12815 , \12826 );
not \U$12451 ( \12828 , \491 );
not \U$12452 ( \12829 , \482 );
not \U$12453 ( \12830 , \487 );
and \U$12454 ( \12831 , \12829 , \12830 );
and \U$12455 ( \12832 , RIc2294a0_127, RIc22b2a0_191);
nor \U$12456 ( \12833 , \12831 , \12832 );
not \U$12457 ( \12834 , \12833 );
not \U$12458 ( \12835 , \12834 );
or \U$12459 ( \12836 , \12828 , \12835 );
nand \U$12460 ( \12837 , \12836 , \493 );
nand \U$12461 ( \12838 , \497 , \499 );
not \U$12462 ( \12839 , \12838 );
and \U$12463 ( \12840 , \12837 , \12839 );
not \U$12464 ( \12841 , \12837 );
and \U$12465 ( \12842 , \12841 , \12838 );
nor \U$12466 ( \12843 , \12840 , \12842 );
buf \U$12467 ( \12844 , \12843 );
buf \U$12468 ( \12845 , \12844 );
not \U$12469 ( \12846 , \12845 );
not \U$12470 ( \12847 , \12846 );
nand \U$12471 ( \12848 , \12847 , RIc2275b0_1);
not \U$12472 ( \12849 , \12848 );
and \U$12473 ( \12850 , \12827 , \12849 );
and \U$12474 ( \12851 , \12815 , \12826 );
or \U$12475 ( \12852 , \12850 , \12851 );
nand \U$12476 ( \12853 , \12802 , \12852 );
nand \U$12477 ( \12854 , \12799 , \12853 );
not \U$12478 ( \12855 , \12854 );
not \U$12479 ( \12856 , \12855 );
or \U$12480 ( \12857 , \12774 , \12856 );
not \U$12481 ( \12858 , \1082 );
not \U$12482 ( \12859 , \12104 );
or \U$12483 ( \12860 , \12858 , \12859 );
not \U$12484 ( \12861 , RIc2274c0_3);
not \U$12485 ( \12862 , \10086 );
not \U$12486 ( \12863 , \12862 );
or \U$12487 ( \12864 , \12861 , \12863 );
nand \U$12488 ( \12865 , \10086 , \1032 );
nand \U$12489 ( \12866 , \12864 , \12865 );
nand \U$12490 ( \12867 , \12866 , \1040 );
nand \U$12491 ( \12868 , \12860 , \12867 );
not \U$12492 ( \12869 , \950 );
not \U$12493 ( \12870 , RIc2273d0_5);
not \U$12494 ( \12871 , \9297 );
or \U$12495 ( \12872 , \12870 , \12871 );
nand \U$12496 ( \12873 , \9299 , \946 );
nand \U$12497 ( \12874 , \12872 , \12873 );
not \U$12498 ( \12875 , \12874 );
or \U$12499 ( \12876 , \12869 , \12875 );
nand \U$12500 ( \12877 , \12136 , \954 );
nand \U$12501 ( \12878 , \12876 , \12877 );
or \U$12502 ( \12879 , \12868 , \12878 );
not \U$12503 ( \12880 , \1120 );
not \U$12504 ( \12881 , \12113 );
or \U$12505 ( \12882 , \12880 , \12881 );
not \U$12506 ( \12883 , RIc2272e0_7);
not \U$12507 ( \12884 , \9255 );
or \U$12508 ( \12885 , \12883 , \12884 );
nand \U$12509 ( \12886 , \10986 , \3027 );
nand \U$12510 ( \12887 , \12885 , \12886 );
nand \U$12511 ( \12888 , \1118 , \12887 );
nand \U$12512 ( \12889 , \12882 , \12888 );
nand \U$12513 ( \12890 , \12879 , \12889 );
nand \U$12514 ( \12891 , \12868 , \12878 );
nand \U$12515 ( \12892 , \12890 , \12891 );
nand \U$12516 ( \12893 , \12857 , \12892 );
nand \U$12517 ( \12894 , \12854 , \12772 );
nand \U$12518 ( \12895 , \12893 , \12894 );
and \U$12519 ( \12896 , \12742 , \12895 );
and \U$12520 ( \12897 , \12660 , \12741 );
or \U$12521 ( \12898 , \12896 , \12897 );
nand \U$12522 ( \12899 , \12658 , \12898 );
nand \U$12523 ( \12900 , \12657 , \12655 );
nand \U$12524 ( \12901 , \12899 , \12900 );
nand \U$12525 ( \12902 , \12653 , \12901 );
nand \U$12526 ( \12903 , \12649 , \12902 );
xor \U$12527 ( \12904 , \12635 , \12903 );
and \U$12528 ( \12905 , \12253 , \12247 );
not \U$12529 ( \12906 , \12253 );
not \U$12530 ( \12907 , \12247 );
and \U$12531 ( \12908 , \12906 , \12907 );
nor \U$12532 ( \12909 , \12905 , \12908 );
and \U$12533 ( \12910 , \12909 , \12258 );
not \U$12534 ( \12911 , \12909 );
not \U$12535 ( \12912 , \12258 );
and \U$12536 ( \12913 , \12911 , \12912 );
nor \U$12537 ( \12914 , \12910 , \12913 );
and \U$12538 ( \12915 , \12904 , \12914 );
and \U$12539 ( \12916 , \12635 , \12903 );
or \U$12540 ( \12917 , \12915 , \12916 );
and \U$12541 ( \12918 , \12633 , \12917 );
and \U$12542 ( \12919 , \12630 , \12632 );
or \U$12543 ( \12920 , \12918 , \12919 );
xnor \U$12544 ( \12921 , \12280 , \12920 );
not \U$12545 ( \12922 , \12921 );
xor \U$12546 ( \12923 , \12630 , \12632 );
xor \U$12547 ( \12924 , \12923 , \12917 );
not \U$12548 ( \12925 , \12924 );
xor \U$12549 ( \12926 , \12089 , \12166 );
xor \U$12550 ( \12927 , \12926 , \12242 );
not \U$12551 ( \12928 , \12927 );
xor \U$12552 ( \12929 , \12203 , \12237 );
xnor \U$12553 ( \12930 , \12929 , \12169 );
not \U$12554 ( \12931 , \12930 );
not \U$12555 ( \12932 , \12931 );
not \U$12556 ( \12933 , \9690 );
not \U$12557 ( \12934 , RIc2262f0_41);
not \U$12558 ( \12935 , \2257 );
or \U$12559 ( \12936 , \12934 , \12935 );
not \U$12560 ( \12937 , RIc2262f0_41);
nand \U$12561 ( \12938 , \4008 , \12937 );
nand \U$12562 ( \12939 , \12936 , \12938 );
not \U$12563 ( \12940 , \12939 );
or \U$12564 ( \12941 , \12933 , \12940 );
nand \U$12565 ( \12942 , \12446 , \9816 );
nand \U$12566 ( \12943 , \12941 , \12942 );
not \U$12567 ( \12944 , \12943 );
buf \U$12568 ( \12945 , \8788 );
not \U$12569 ( \12946 , \12945 );
not \U$12570 ( \12947 , \12433 );
or \U$12571 ( \12948 , \12946 , \12947 );
not \U$12572 ( \12949 , RIc225d50_53);
not \U$12573 ( \12950 , \9539 );
or \U$12574 ( \12951 , \12949 , \12950 );
nand \U$12575 ( \12952 , \1169 , \11585 );
nand \U$12576 ( \12953 , \12951 , \12952 );
nand \U$12577 ( \12954 , \12953 , \8777 );
nand \U$12578 ( \12955 , \12948 , \12954 );
not \U$12579 ( \12956 , \12955 );
or \U$12580 ( \12957 , \12944 , \12956 );
or \U$12581 ( \12958 , \12943 , \12955 );
not \U$12582 ( \12959 , \9459 );
not \U$12583 ( \12960 , RIc225e40_51);
not \U$12584 ( \12961 , \1391 );
not \U$12585 ( \12962 , \12961 );
or \U$12586 ( \12963 , \12960 , \12962 );
nand \U$12587 ( \12964 , \1391 , \9450 );
nand \U$12588 ( \12965 , \12963 , \12964 );
not \U$12589 ( \12966 , \12965 );
or \U$12590 ( \12967 , \12959 , \12966 );
nand \U$12591 ( \12968 , \12425 , \9445 );
nand \U$12592 ( \12969 , \12967 , \12968 );
nand \U$12593 ( \12970 , \12958 , \12969 );
nand \U$12594 ( \12971 , \12957 , \12970 );
not \U$12595 ( \12972 , \12971 );
not \U$12596 ( \12973 , \3631 );
not \U$12597 ( \12974 , \12553 );
or \U$12598 ( \12975 , \12973 , \12974 );
not \U$12599 ( \12976 , RIc2266b0_33);
not \U$12600 ( \12977 , \3008 );
not \U$12601 ( \12978 , \12977 );
or \U$12602 ( \12979 , \12976 , \12978 );
nand \U$12603 ( \12980 , \3008 , \5179 );
nand \U$12604 ( \12981 , \12979 , \12980 );
nand \U$12605 ( \12982 , \12981 , \3629 );
nand \U$12606 ( \12983 , \12975 , \12982 );
not \U$12607 ( \12984 , \12983 );
not \U$12608 ( \12985 , \4381 );
not \U$12609 ( \12986 , RIc2265c0_35);
not \U$12610 ( \12987 , \2499 );
or \U$12611 ( \12988 , \12986 , \12987 );
not \U$12612 ( \12989 , \4194 );
not \U$12613 ( \12990 , \12989 );
nand \U$12614 ( \12991 , \12990 , \3620 );
nand \U$12615 ( \12992 , \12988 , \12991 );
not \U$12616 ( \12993 , \12992 );
or \U$12617 ( \12994 , \12985 , \12993 );
nand \U$12618 ( \12995 , \12567 , \4383 );
nand \U$12619 ( \12996 , \12994 , \12995 );
not \U$12620 ( \12997 , \12996 );
nand \U$12621 ( \12998 , \12984 , \12997 );
not \U$12622 ( \12999 , \10445 );
not \U$12623 ( \13000 , RIc225f30_49);
not \U$12624 ( \13001 , \10909 );
or \U$12625 ( \13002 , \13000 , \13001 );
nand \U$12626 ( \13003 , \1331 , \9549 );
nand \U$12627 ( \13004 , \13002 , \13003 );
not \U$12628 ( \13005 , \13004 );
or \U$12629 ( \13006 , \12999 , \13005 );
nand \U$12630 ( \13007 , \12579 , \9552 );
nand \U$12631 ( \13008 , \13006 , \13007 );
and \U$12632 ( \13009 , \12998 , \13008 );
nand \U$12633 ( \13010 , \12983 , \12996 );
not \U$12634 ( \13011 , \13010 );
nor \U$12635 ( \13012 , \13009 , \13011 );
not \U$12636 ( \13013 , \13012 );
not \U$12637 ( \13014 , \13013 );
or \U$12638 ( \13015 , \12972 , \13014 );
not \U$12639 ( \13016 , \11117 );
not \U$12640 ( \13017 , RIc225c60_55);
not \U$12641 ( \13018 , \982 );
or \U$12642 ( \13019 , \13017 , \13018 );
nand \U$12643 ( \13020 , \981 , \11041 );
nand \U$12644 ( \13021 , \13019 , \13020 );
not \U$12645 ( \13022 , \13021 );
or \U$12646 ( \13023 , \13016 , \13022 );
not \U$12647 ( \13024 , \11039 );
buf \U$12648 ( \13025 , \13024 );
nand \U$12649 ( \13026 , \12541 , \13025 );
nand \U$12650 ( \13027 , \13023 , \13026 );
not \U$12651 ( \13028 , \13027 );
not \U$12652 ( \13029 , \13028 );
not \U$12653 ( \13030 , \6307 );
not \U$12654 ( \13031 , \12511 );
or \U$12655 ( \13032 , \13030 , \13031 );
not \U$12656 ( \13033 , RIc2263e0_39);
not \U$12657 ( \13034 , \9584 );
or \U$12658 ( \13035 , \13033 , \13034 );
nand \U$12659 ( \13036 , \2014 , \5498 );
nand \U$12660 ( \13037 , \13035 , \13036 );
nand \U$12661 ( \13038 , \13037 , \6689 );
nand \U$12662 ( \13039 , \13032 , \13038 );
not \U$12663 ( \13040 , \13039 );
not \U$12664 ( \13041 , \13040 );
or \U$12665 ( \13042 , \13029 , \13041 );
not \U$12666 ( \13043 , \5509 );
not \U$12667 ( \13044 , RIc2264d0_37);
not \U$12668 ( \13045 , \2555 );
or \U$12669 ( \13046 , \13044 , \13045 );
nand \U$12670 ( \13047 , \10899 , \5504 );
nand \U$12671 ( \13048 , \13046 , \13047 );
not \U$12672 ( \13049 , \13048 );
or \U$12673 ( \13050 , \13043 , \13049 );
nand \U$12674 ( \13051 , \12524 , \5519 );
nand \U$12675 ( \13052 , \13050 , \13051 );
nand \U$12676 ( \13053 , \13042 , \13052 );
nand \U$12677 ( \13054 , \13039 , \13027 );
nand \U$12678 ( \13055 , \13053 , \13054 );
not \U$12679 ( \13056 , \12971 );
nand \U$12680 ( \13057 , \13056 , \13012 );
nand \U$12681 ( \13058 , \13055 , \13057 );
nand \U$12682 ( \13059 , \13015 , \13058 );
not \U$12683 ( \13060 , \13059 );
or \U$12684 ( \13061 , \12932 , \13060 );
or \U$12685 ( \13062 , \12931 , \13059 );
xor \U$12686 ( \13063 , \12095 , \12106 );
xor \U$12687 ( \13064 , \13063 , \12117 );
not \U$12688 ( \13065 , \9110 );
and \U$12689 ( \13066 , \2443 , \9117 );
not \U$12690 ( \13067 , \2443 );
and \U$12691 ( \13068 , \13067 , RIc226200_43);
or \U$12692 ( \13069 , \13066 , \13068 );
not \U$12693 ( \13070 , \13069 );
or \U$12694 ( \13071 , \13065 , \13070 );
nand \U$12695 ( \13072 , \12460 , \9129 );
nand \U$12696 ( \13073 , \13071 , \13072 );
not \U$12697 ( \13074 , \13073 );
not \U$12698 ( \13075 , \11965 );
not \U$12699 ( \13076 , RIc225b70_57);
not \U$12700 ( \13077 , \888 );
not \U$12701 ( \13078 , \13077 );
or \U$12702 ( \13079 , \13076 , \13078 );
nand \U$12703 ( \13080 , \888 , \10074 );
nand \U$12704 ( \13081 , \13079 , \13080 );
not \U$12705 ( \13082 , \13081 );
or \U$12706 ( \13083 , \13075 , \13082 );
nand \U$12707 ( \13084 , \12477 , \11974 );
nand \U$12708 ( \13085 , \13083 , \13084 );
not \U$12709 ( \13086 , \13085 );
or \U$12710 ( \13087 , \13074 , \13086 );
or \U$12711 ( \13088 , \13085 , \13073 );
and \U$12712 ( \13089 , \12497 , \2154 );
not \U$12713 ( \13090 , RIc226980_27);
not \U$12714 ( \13091 , \4049 );
or \U$12715 ( \13092 , \13090 , \13091 );
nand \U$12716 ( \13093 , \3640 , \2133 );
nand \U$12717 ( \13094 , \13092 , \13093 );
and \U$12718 ( \13095 , \13094 , \2138 );
nor \U$12719 ( \13096 , \13089 , \13095 );
not \U$12720 ( \13097 , \13096 );
nand \U$12721 ( \13098 , \13088 , \13097 );
nand \U$12722 ( \13099 , \13087 , \13098 );
xor \U$12723 ( \13100 , \13064 , \13099 );
not \U$12724 ( \13101 , \2784 );
not \U$12725 ( \13102 , \3115 );
and \U$12726 ( \13103 , RIc226890_29, \13102 );
not \U$12727 ( \13104 , RIc226890_29);
and \U$12728 ( \13105 , \13104 , \11320 );
or \U$12729 ( \13106 , \13103 , \13105 );
not \U$12730 ( \13107 , \13106 );
or \U$12731 ( \13108 , \13101 , \13107 );
nand \U$12732 ( \13109 , \12395 , \9142 );
nand \U$12733 ( \13110 , \13108 , \13109 );
not \U$12734 ( \13111 , \9934 );
not \U$12735 ( \13112 , RIc226110_45);
not \U$12736 ( \13113 , \2298 );
or \U$12737 ( \13114 , \13112 , \13113 );
not \U$12738 ( \13115 , RIc226110_45);
nand \U$12739 ( \13116 , \13115 , \10935 );
nand \U$12740 ( \13117 , \13114 , \13116 );
not \U$12741 ( \13118 , \13117 );
or \U$12742 ( \13119 , \13111 , \13118 );
nand \U$12743 ( \13120 , \12386 , \9398 );
nand \U$12744 ( \13121 , \13119 , \13120 );
or \U$12745 ( \13122 , \13110 , \13121 );
not \U$12746 ( \13123 , \1311 );
not \U$12747 ( \13124 , \12408 );
or \U$12748 ( \13125 , \13123 , \13124 );
not \U$12749 ( \13126 , RIc227100_11);
not \U$12750 ( \13127 , \9215 );
or \U$12751 ( \13128 , \13126 , \13127 );
not \U$12752 ( \13129 , \8924 );
not \U$12753 ( \13130 , \13129 );
nand \U$12754 ( \13131 , \13130 , \1291 );
nand \U$12755 ( \13132 , \13128 , \13131 );
nand \U$12756 ( \13133 , \13132 , \9904 );
nand \U$12757 ( \13134 , \13125 , \13133 );
nand \U$12758 ( \13135 , \13122 , \13134 );
nand \U$12759 ( \13136 , \13110 , \13121 );
nand \U$12760 ( \13137 , \13135 , \13136 );
and \U$12761 ( \13138 , \13100 , \13137 );
and \U$12762 ( \13139 , \13064 , \13099 );
or \U$12763 ( \13140 , \13138 , \13139 );
nand \U$12764 ( \13141 , \13062 , \13140 );
nand \U$12765 ( \13142 , \13061 , \13141 );
not \U$12766 ( \13143 , \13142 );
or \U$12767 ( \13144 , \12928 , \13143 );
or \U$12768 ( \13145 , \12927 , \13142 );
xor \U$12769 ( \13146 , \12379 , \12415 );
xor \U$12770 ( \13147 , \13146 , \12451 );
not \U$12771 ( \13148 , \13147 );
not \U$12772 ( \13149 , \12331 );
not \U$12773 ( \13150 , \12324 );
or \U$12774 ( \13151 , \13149 , \13150 );
or \U$12775 ( \13152 , \12324 , \12331 );
nand \U$12776 ( \13153 , \13151 , \13152 );
xnor \U$12777 ( \13154 , \13153 , \12321 );
not \U$12778 ( \13155 , \13154 );
not \U$12779 ( \13156 , \13155 );
or \U$12780 ( \13157 , \13148 , \13156 );
not \U$12781 ( \13158 , \13154 );
not \U$12782 ( \13159 , \13147 );
not \U$12783 ( \13160 , \13159 );
or \U$12784 ( \13161 , \13158 , \13160 );
xor \U$12785 ( \13162 , \12222 , \12216 );
xnor \U$12786 ( \13163 , \13162 , \12234 );
xor \U$12787 ( \13164 , \12179 , \12186 );
xor \U$12788 ( \13165 , \13164 , \12201 );
not \U$12789 ( \13166 , \13165 );
nand \U$12790 ( \13167 , \13163 , \13166 );
not \U$12791 ( \13168 , \13167 );
xor \U$12792 ( \13169 , \12294 , \12306 );
xor \U$12793 ( \13170 , \13169 , \12318 );
not \U$12794 ( \13171 , \13170 );
or \U$12795 ( \13172 , \13168 , \13171 );
not \U$12796 ( \13173 , \13166 );
xor \U$12797 ( \13174 , \12222 , \12216 );
xor \U$12798 ( \13175 , \13174 , \12234 );
nand \U$12799 ( \13176 , \13173 , \13175 );
nand \U$12800 ( \13177 , \13172 , \13176 );
nand \U$12801 ( \13178 , \13161 , \13177 );
nand \U$12802 ( \13179 , \13157 , \13178 );
nand \U$12803 ( \13180 , \13145 , \13179 );
nand \U$12804 ( \13181 , \13144 , \13180 );
xor \U$12805 ( \13182 , \12290 , \12346 );
xor \U$12806 ( \13183 , \13182 , \12365 );
xor \U$12807 ( \13184 , \13181 , \13183 );
xor \U$12808 ( \13185 , \12454 , \12587 );
xor \U$12809 ( \13186 , \13185 , \12611 );
xor \U$12810 ( \13187 , \12292 , \12337 );
xor \U$12811 ( \13188 , \13187 , \12343 );
xor \U$12812 ( \13189 , \13186 , \13188 );
xor \U$12813 ( \13190 , \12412 , \12390 );
xnor \U$12814 ( \13191 , \13190 , \12399 );
not \U$12815 ( \13192 , \13191 );
xor \U$12816 ( \13193 , \12581 , \12569 );
xor \U$12817 ( \13194 , \13193 , \12559 );
not \U$12818 ( \13195 , \13194 );
or \U$12819 ( \13196 , \13192 , \13195 );
not \U$12820 ( \13197 , \854 );
not \U$12821 ( \13198 , \12755 );
and \U$12822 ( \13199 , RIc2275b0_1, \13198 );
not \U$12823 ( \13200 , RIc2275b0_1);
and \U$12824 ( \13201 , \13200 , \12755 );
or \U$12825 ( \13202 , \13199 , \13201 );
not \U$12826 ( \13203 , \13202 );
or \U$12827 ( \13204 , \13197 , \13203 );
nand \U$12828 ( \13205 , \12091 , \1579 );
nand \U$12829 ( \13206 , \13204 , \13205 );
not \U$12830 ( \13207 , \1081 );
not \U$12831 ( \13208 , \12866 );
or \U$12832 ( \13209 , \13207 , \13208 );
not \U$12833 ( \13210 , RIc2274c0_3);
buf \U$12834 ( \13211 , \10369 );
not \U$12835 ( \13212 , \13211 );
or \U$12836 ( \13213 , \13210 , \13212 );
nand \U$12837 ( \13214 , \10197 , \1032 );
nand \U$12838 ( \13215 , \13213 , \13214 );
nand \U$12839 ( \13216 , \1040 , \13215 );
nand \U$12840 ( \13217 , \13209 , \13216 );
xor \U$12841 ( \13218 , \13206 , \13217 );
not \U$12842 ( \13219 , \1339 );
not \U$12843 ( \13220 , \12767 );
or \U$12844 ( \13221 , \13219 , \13220 );
not \U$12845 ( \13222 , RIc2271f0_9);
not \U$12846 ( \13223 , \10110 );
not \U$12847 ( \13224 , \13223 );
or \U$12848 ( \13225 , \13222 , \13224 );
nand \U$12849 ( \13226 , \10110 , \1342 );
nand \U$12850 ( \13227 , \13225 , \13226 );
nand \U$12851 ( \13228 , \13227 , \1363 );
nand \U$12852 ( \13229 , \13221 , \13228 );
and \U$12853 ( \13230 , \13218 , \13229 );
and \U$12854 ( \13231 , \13206 , \13217 );
or \U$12855 ( \13232 , \13230 , \13231 );
not \U$12856 ( \13233 , \9641 );
not \U$12857 ( \13234 , RIc226020_47);
not \U$12858 ( \13235 , \1729 );
not \U$12859 ( \13236 , \13235 );
or \U$12860 ( \13237 , \13234 , \13236 );
nand \U$12861 ( \13238 , \9196 , \9373 );
nand \U$12862 ( \13239 , \13237 , \13238 );
not \U$12863 ( \13240 , \13239 );
or \U$12864 ( \13241 , \13233 , \13240 );
nand \U$12865 ( \13242 , \12301 , \9619 );
nand \U$12866 ( \13243 , \13241 , \13242 );
xor \U$12867 ( \13244 , \13232 , \13243 );
not \U$12868 ( \13245 , \3653 );
not \U$12869 ( \13246 , \12314 );
or \U$12870 ( \13247 , \13245 , \13246 );
not \U$12871 ( \13248 , RIc2267a0_31);
not \U$12872 ( \13249 , \4227 );
or \U$12873 ( \13250 , \13248 , \13249 );
not \U$12874 ( \13251 , \4227 );
nand \U$12875 ( \13252 , \13251 , \3648 );
nand \U$12876 ( \13253 , \13250 , \13252 );
nand \U$12877 ( \13254 , \13253 , \2697 );
nand \U$12878 ( \13255 , \13247 , \13254 );
and \U$12879 ( \13256 , \13244 , \13255 );
and \U$12880 ( \13257 , \13232 , \13243 );
or \U$12881 ( \13258 , \13256 , \13257 );
nand \U$12882 ( \13259 , \13196 , \13258 );
not \U$12883 ( \13260 , \13194 );
not \U$12884 ( \13261 , \13191 );
nand \U$12885 ( \13262 , \13260 , \13261 );
nand \U$12886 ( \13263 , \13259 , \13262 );
xor \U$12887 ( \13264 , \12503 , \12545 );
xor \U$12888 ( \13265 , \13264 , \12584 );
xor \U$12889 ( \13266 , \13263 , \13265 );
and \U$12890 ( \13267 , \12543 , \12528 );
not \U$12891 ( \13268 , \12543 );
not \U$12892 ( \13269 , \12528 );
and \U$12893 ( \13270 , \13268 , \13269 );
nor \U$12894 ( \13271 , \13267 , \13270 );
not \U$12895 ( \13272 , \12515 );
and \U$12896 ( \13273 , \13271 , \13272 );
not \U$12897 ( \13274 , \13271 );
and \U$12898 ( \13275 , \13274 , \12515 );
nor \U$12899 ( \13276 , \13273 , \13275 );
not \U$12900 ( \13277 , \13276 );
buf \U$12901 ( \13278 , \12486 );
xor \U$12902 ( \13279 , \12480 , \13278 );
xnor \U$12903 ( \13280 , \13279 , \12501 );
not \U$12904 ( \13281 , \13280 );
or \U$12905 ( \13282 , \13277 , \13281 );
xor \U$12906 ( \13283 , \12427 , \12437 );
xor \U$12907 ( \13284 , \13283 , \12448 );
nand \U$12908 ( \13285 , \13282 , \13284 );
not \U$12909 ( \13286 , \13276 );
not \U$12910 ( \13287 , \13280 );
nand \U$12911 ( \13288 , \13286 , \13287 );
nand \U$12912 ( \13289 , \13285 , \13288 );
and \U$12913 ( \13290 , \13266 , \13289 );
and \U$12914 ( \13291 , \13263 , \13265 );
or \U$12915 ( \13292 , \13290 , \13291 );
and \U$12916 ( \13293 , \13189 , \13292 );
and \U$12917 ( \13294 , \13186 , \13188 );
or \U$12918 ( \13295 , \13293 , \13294 );
and \U$12919 ( \13296 , \13184 , \13295 );
and \U$12920 ( \13297 , \13181 , \13183 );
or \U$12921 ( \13298 , \13296 , \13297 );
xor \U$12922 ( \13299 , \12368 , \12624 );
xor \U$12923 ( \13300 , \13299 , \12627 );
xor \U$12924 ( \13301 , \13298 , \13300 );
xor \U$12925 ( \13302 , \12614 , \12622 );
xor \U$12926 ( \13303 , \13302 , \12375 );
not \U$12927 ( \13304 , \13303 );
not \U$12928 ( \13305 , \13304 );
not \U$12929 ( \13306 , \12901 );
not \U$12930 ( \13307 , \12643 );
not \U$12931 ( \13308 , \13307 );
or \U$12932 ( \13309 , \13306 , \13308 );
not \U$12933 ( \13310 , \12901 );
nand \U$12934 ( \13311 , \13310 , \12643 );
nand \U$12935 ( \13312 , \13309 , \13311 );
and \U$12936 ( \13313 , \13312 , \12646 );
not \U$12937 ( \13314 , \13312 );
and \U$12938 ( \13315 , \13314 , \12647 );
nor \U$12939 ( \13316 , \13313 , \13315 );
not \U$12940 ( \13317 , \13316 );
not \U$12941 ( \13318 , \13317 );
or \U$12942 ( \13319 , \13305 , \13318 );
not \U$12943 ( \13320 , \13316 );
not \U$12944 ( \13321 , \13303 );
or \U$12945 ( \13322 , \13320 , \13321 );
xor \U$12946 ( \13323 , \12349 , \12359 );
xor \U$12947 ( \13324 , \13323 , \12362 );
not \U$12948 ( \13325 , \13324 );
xor \U$12949 ( \13326 , \12898 , \12657 );
xnor \U$12950 ( \13327 , \13326 , \12655 );
not \U$12951 ( \13328 , \13327 );
not \U$12952 ( \13329 , \13328 );
or \U$12953 ( \13330 , \13325 , \13329 );
not \U$12954 ( \13331 , \13324 );
not \U$12955 ( \13332 , \13331 );
not \U$12956 ( \13333 , \13327 );
or \U$12957 ( \13334 , \13332 , \13333 );
xor \U$12958 ( \13335 , \12351 , \12353 );
xor \U$12959 ( \13336 , \13335 , \12356 );
not \U$12960 ( \13337 , \13336 );
not \U$12961 ( \13338 , \12602 );
not \U$12962 ( \13339 , \12606 );
or \U$12963 ( \13340 , \13338 , \13339 );
or \U$12964 ( \13341 , \12602 , \12606 );
nand \U$12965 ( \13342 , \13340 , \13341 );
and \U$12966 ( \13343 , \13342 , \12591 );
not \U$12967 ( \13344 , \13342 );
and \U$12968 ( \13345 , \13344 , \12609 );
nor \U$12969 ( \13346 , \13343 , \13345 );
nand \U$12970 ( \13347 , \13337 , \13346 );
xor \U$12971 ( \13348 , \12757 , \12758 );
xor \U$12972 ( \13349 , \13348 , \12769 );
not \U$12973 ( \13350 , \13349 );
xor \U$12974 ( \13351 , \12868 , \12878 );
xnor \U$12975 ( \13352 , \13351 , \12889 );
nand \U$12976 ( \13353 , \13350 , \13352 );
not \U$12977 ( \13354 , \13353 );
xor \U$12978 ( \13355 , \12815 , \12826 );
xor \U$12979 ( \13356 , \13355 , \12849 );
not \U$12980 ( \13357 , \1963 );
not \U$12981 ( \13358 , \12729 );
or \U$12982 ( \13359 , \13357 , \13358 );
not \U$12983 ( \13360 , RIc226e30_17);
not \U$12984 ( \13361 , \8830 );
or \U$12985 ( \13362 , \13360 , \13361 );
nand \U$12986 ( \13363 , \10289 , \1952 );
nand \U$12987 ( \13364 , \13362 , \13363 );
nand \U$12988 ( \13365 , \1945 , \13364 );
nand \U$12989 ( \13366 , \13359 , \13365 );
xor \U$12990 ( \13367 , \13356 , \13366 );
not \U$12991 ( \13368 , \2320 );
not \U$12992 ( \13369 , RIc226f20_15);
not \U$12993 ( \13370 , \8952 );
not \U$12994 ( \13371 , \13370 );
or \U$12995 ( \13372 , \13369 , \13371 );
nand \U$12996 ( \13373 , \8951 , \1674 );
nand \U$12997 ( \13374 , \13372 , \13373 );
not \U$12998 ( \13375 , \13374 );
or \U$12999 ( \13376 , \13368 , \13375 );
nand \U$13000 ( \13377 , \12679 , \2358 );
nand \U$13001 ( \13378 , \13376 , \13377 );
and \U$13002 ( \13379 , \13367 , \13378 );
and \U$13003 ( \13380 , \13356 , \13366 );
or \U$13004 ( \13381 , \13379 , \13380 );
not \U$13005 ( \13382 , \13381 );
or \U$13006 ( \13383 , \13354 , \13382 );
not \U$13007 ( \13384 , \13352 );
nand \U$13008 ( \13385 , \13384 , \13349 );
nand \U$13009 ( \13386 , \13383 , \13385 );
not \U$13010 ( \13387 , \13386 );
and \U$13011 ( \13388 , \12892 , \12773 );
not \U$13012 ( \13389 , \12892 );
and \U$13013 ( \13390 , \13389 , \12772 );
or \U$13014 ( \13391 , \13388 , \13390 );
xor \U$13015 ( \13392 , \13391 , \12855 );
not \U$13016 ( \13393 , \13392 );
not \U$13017 ( \13394 , \13393 );
or \U$13018 ( \13395 , \13387 , \13394 );
not \U$13019 ( \13396 , \13386 );
not \U$13020 ( \13397 , \13396 );
not \U$13021 ( \13398 , \13392 );
or \U$13022 ( \13399 , \13397 , \13398 );
not \U$13023 ( \13400 , \2367 );
not \U$13024 ( \13401 , \12702 );
or \U$13025 ( \13402 , \13400 , \13401 );
not \U$13026 ( \13403 , RIc226c50_21);
not \U$13027 ( \13404 , \6719 );
or \U$13028 ( \13405 , \13403 , \13404 );
nand \U$13029 ( \13406 , \9740 , \4475 );
nand \U$13030 ( \13407 , \13405 , \13406 );
nand \U$13031 ( \13408 , \13407 , \2392 );
nand \U$13032 ( \13409 , \13402 , \13408 );
not \U$13033 ( \13410 , \13409 );
not \U$13034 ( \13411 , \1930 );
not \U$13035 ( \13412 , \12793 );
or \U$13036 ( \13413 , \13411 , \13412 );
not \U$13037 ( \13414 , RIc226b60_23);
not \U$13038 ( \13415 , \9765 );
or \U$13039 ( \13416 , \13414 , \13415 );
nand \U$13040 ( \13417 , \6071 , \1927 );
nand \U$13041 ( \13418 , \13416 , \13417 );
nand \U$13042 ( \13419 , \13418 , \1915 );
nand \U$13043 ( \13420 , \13413 , \13419 );
not \U$13044 ( \13421 , \13420 );
nand \U$13045 ( \13422 , \13410 , \13421 );
not \U$13046 ( \13423 , \2534 );
not \U$13047 ( \13424 , \12714 );
or \U$13048 ( \13425 , \13423 , \13424 );
not \U$13049 ( \13426 , RIc226d40_19);
not \U$13050 ( \13427 , \12228 );
or \U$13051 ( \13428 , \13426 , \13427 );
nand \U$13052 ( \13429 , \8885 , \2523 );
nand \U$13053 ( \13430 , \13428 , \13429 );
nand \U$13054 ( \13431 , \13430 , \2518 );
nand \U$13055 ( \13432 , \13425 , \13431 );
and \U$13056 ( \13433 , \13422 , \13432 );
nor \U$13057 ( \13434 , \13421 , \13410 );
nor \U$13058 ( \13435 , \13433 , \13434 );
not \U$13059 ( \13436 , \13435 );
not \U$13060 ( \13437 , \13436 );
not \U$13061 ( \13438 , \954 );
not \U$13062 ( \13439 , \12874 );
or \U$13063 ( \13440 , \13438 , \13439 );
not \U$13064 ( \13441 , RIc2273d0_5);
not \U$13065 ( \13442 , \9324 );
not \U$13066 ( \13443 , \13442 );
or \U$13067 ( \13444 , \13441 , \13443 );
nand \U$13068 ( \13445 , \9320 , \946 );
nand \U$13069 ( \13446 , \13444 , \13445 );
nand \U$13070 ( \13447 , \13446 , \950 );
nand \U$13071 ( \13448 , \13440 , \13447 );
not \U$13072 ( \13449 , \1121 );
not \U$13073 ( \13450 , \12887 );
or \U$13074 ( \13451 , \13449 , \13450 );
not \U$13075 ( \13452 , RIc2272e0_7);
not \U$13076 ( \13453 , \9275 );
not \U$13077 ( \13454 , \13453 );
or \U$13078 ( \13455 , \13452 , \13454 );
nand \U$13079 ( \13456 , \9275 , \1139 );
nand \U$13080 ( \13457 , \13455 , \13456 );
nand \U$13081 ( \13458 , \13457 , \1118 );
nand \U$13082 ( \13459 , \13451 , \13458 );
xor \U$13083 ( \13460 , \13448 , \13459 );
not \U$13084 ( \13461 , \1311 );
not \U$13085 ( \13462 , \13132 );
or \U$13086 ( \13463 , \13461 , \13462 );
not \U$13087 ( \13464 , RIc227100_11);
buf \U$13088 ( \13465 , \9224 );
not \U$13089 ( \13466 , \13465 );
or \U$13090 ( \13467 , \13464 , \13466 );
nand \U$13091 ( \13468 , \9051 , \1685 );
nand \U$13092 ( \13469 , \13467 , \13468 );
nand \U$13093 ( \13470 , \13469 , \1307 );
nand \U$13094 ( \13471 , \13463 , \13470 );
and \U$13095 ( \13472 , \13460 , \13471 );
and \U$13096 ( \13473 , \13448 , \13459 );
or \U$13097 ( \13474 , \13472 , \13473 );
not \U$13098 ( \13475 , \13474 );
or \U$13099 ( \13476 , \13437 , \13475 );
not \U$13100 ( \13477 , \13474 );
not \U$13101 ( \13478 , \13477 );
not \U$13102 ( \13479 , \13435 );
or \U$13103 ( \13480 , \13478 , \13479 );
not \U$13104 ( \13481 , RIc2275b0_1);
and \U$13105 ( \13482 , \493 , \491 );
nor \U$13106 ( \13483 , \12833 , \13482 );
not \U$13107 ( \13484 , \13483 );
nand \U$13108 ( \13485 , \12833 , \13482 );
nand \U$13109 ( \13486 , \13484 , \13485 );
buf \U$13110 ( \13487 , \13486 );
buf \U$13111 ( \13488 , \13487 );
not \U$13112 ( \13489 , \13488 );
or \U$13113 ( \13490 , \13481 , \13489 );
nand \U$13114 ( \13491 , \13490 , RIc2258a0_63);
xor \U$13115 ( \13492 , \13491 , \12848 );
not \U$13116 ( \13493 , \1081 );
not \U$13117 ( \13494 , \13215 );
or \U$13118 ( \13495 , \13493 , \13494 );
not \U$13119 ( \13496 , RIc2274c0_3);
buf \U$13120 ( \13497 , \10355 );
not \U$13121 ( \13498 , \13497 );
not \U$13122 ( \13499 , \13498 );
or \U$13123 ( \13500 , \13496 , \13499 );
nand \U$13124 ( \13501 , \13497 , \2896 );
nand \U$13125 ( \13502 , \13500 , \13501 );
nand \U$13126 ( \13503 , \13502 , \1040 );
nand \U$13127 ( \13504 , \13495 , \13503 );
and \U$13128 ( \13505 , \13492 , \13504 );
and \U$13129 ( \13506 , \13491 , \12848 );
or \U$13130 ( \13507 , \13505 , \13506 );
not \U$13131 ( \13508 , \2173 );
not \U$13132 ( \13509 , \12783 );
or \U$13133 ( \13510 , \13508 , \13509 );
not \U$13134 ( \13511 , RIc226a70_25);
not \U$13135 ( \13512 , \5215 );
not \U$13136 ( \13513 , \13512 );
or \U$13137 ( \13514 , \13511 , \13513 );
not \U$13138 ( \13515 , \9850 );
nand \U$13139 ( \13516 , \13515 , \9662 );
nand \U$13140 ( \13517 , \13514 , \13516 );
nand \U$13141 ( \13518 , \13517 , \2195 );
nand \U$13142 ( \13519 , \13510 , \13518 );
xor \U$13143 ( \13520 , \13507 , \13519 );
not \U$13144 ( \13521 , \2154 );
not \U$13145 ( \13522 , \13094 );
or \U$13146 ( \13523 , \13521 , \13522 );
not \U$13147 ( \13524 , RIc226980_27);
not \U$13148 ( \13525 , \4121 );
not \U$13149 ( \13526 , \13525 );
or \U$13150 ( \13527 , \13524 , \13526 );
not \U$13151 ( \13528 , \4122 );
nand \U$13152 ( \13529 , \13528 , \2150 );
nand \U$13153 ( \13530 , \13527 , \13529 );
nand \U$13154 ( \13531 , \13530 , \2138 );
nand \U$13155 ( \13532 , \13523 , \13531 );
and \U$13156 ( \13533 , \13520 , \13532 );
and \U$13157 ( \13534 , \13507 , \13519 );
or \U$13158 ( \13535 , \13533 , \13534 );
nand \U$13159 ( \13536 , \13480 , \13535 );
nand \U$13160 ( \13537 , \13476 , \13536 );
nand \U$13161 ( \13538 , \13399 , \13537 );
nand \U$13162 ( \13539 , \13395 , \13538 );
and \U$13163 ( \13540 , \13347 , \13539 );
nor \U$13164 ( \13541 , \13346 , \13337 );
nor \U$13165 ( \13542 , \13540 , \13541 );
not \U$13166 ( \13543 , \13542 );
nand \U$13167 ( \13544 , \13334 , \13543 );
nand \U$13168 ( \13545 , \13330 , \13544 );
nand \U$13169 ( \13546 , \13322 , \13545 );
nand \U$13170 ( \13547 , \13319 , \13546 );
and \U$13171 ( \13548 , \13301 , \13547 );
and \U$13172 ( \13549 , \13298 , \13300 );
or \U$13173 ( \13550 , \13548 , \13549 );
not \U$13174 ( \13551 , \13550 );
xor \U$13175 ( \13552 , \12271 , \12260 );
xor \U$13176 ( \13553 , \13552 , \12276 );
not \U$13177 ( \13554 , \13553 );
nand \U$13178 ( \13555 , \13551 , \13554 );
not \U$13179 ( \13556 , \13555 );
or \U$13180 ( \13557 , \12925 , \13556 );
nand \U$13181 ( \13558 , \13550 , \13553 );
nand \U$13182 ( \13559 , \13557 , \13558 );
not \U$13183 ( \13560 , \13559 );
nand \U$13184 ( \13561 , \12922 , \13560 );
not \U$13185 ( \13562 , \9973 );
not \U$13186 ( \13563 , \10041 );
or \U$13187 ( \13564 , \13562 , \13563 );
or \U$13188 ( \13565 , \10041 , \9973 );
nand \U$13189 ( \13566 , \13565 , \9980 );
nand \U$13190 ( \13567 , \13564 , \13566 );
not \U$13191 ( \13568 , \13567 );
not \U$13192 ( \13569 , \13568 );
not \U$13193 ( \13570 , \10574 );
not \U$13194 ( \13571 , \13570 );
not \U$13195 ( \13572 , \10696 );
or \U$13196 ( \13573 , \13571 , \13572 );
or \U$13197 ( \13574 , \10696 , \13570 );
nand \U$13198 ( \13575 , \13574 , \10687 );
nand \U$13199 ( \13576 , \13573 , \13575 );
not \U$13200 ( \13577 , \13576 );
or \U$13201 ( \13578 , \13569 , \13577 );
or \U$13202 ( \13579 , \13576 , \13568 );
nand \U$13203 ( \13580 , \13578 , \13579 );
nor \U$13204 ( \13581 , \10564 , \10568 );
or \U$13205 ( \13582 , \13581 , \10573 );
nand \U$13206 ( \13583 , \10564 , \10568 );
nand \U$13207 ( \13584 , \13582 , \13583 );
nor \U$13208 ( \13585 , \10743 , \10708 );
or \U$13209 ( \13586 , \13585 , \10775 );
nand \U$13210 ( \13587 , \10743 , \10708 );
nand \U$13211 ( \13588 , \13586 , \13587 );
buf \U$13212 ( \13589 , \13588 );
xor \U$13213 ( \13590 , \13584 , \13589 );
xor \U$13214 ( \13591 , \10604 , \10640 );
and \U$13215 ( \13592 , \13591 , \10686 );
and \U$13216 ( \13593 , \10604 , \10640 );
or \U$13217 ( \13594 , \13592 , \13593 );
xnor \U$13218 ( \13595 , \13590 , \13594 );
and \U$13219 ( \13596 , \13580 , \13595 );
not \U$13220 ( \13597 , \13580 );
not \U$13221 ( \13598 , \13595 );
and \U$13222 ( \13599 , \13597 , \13598 );
nor \U$13223 ( \13600 , \13596 , \13599 );
not \U$13224 ( \13601 , \11027 );
not \U$13225 ( \13602 , \10558 );
not \U$13226 ( \13603 , \13602 );
or \U$13227 ( \13604 , \13601 , \13603 );
not \U$13228 ( \13605 , \11026 );
not \U$13229 ( \13606 , \10558 );
or \U$13230 ( \13607 , \13605 , \13606 );
nand \U$13231 ( \13608 , \13607 , \10700 );
nand \U$13232 ( \13609 , \13604 , \13608 );
xor \U$13233 ( \13610 , \13600 , \13609 );
or \U$13234 ( \13611 , \10890 , \10785 );
and \U$13235 ( \13612 , \13611 , \11025 );
and \U$13236 ( \13613 , \10890 , \10785 );
nor \U$13237 ( \13614 , \13612 , \13613 );
and \U$13238 ( \13615 , RIc2275b0_1, \10110 );
not \U$13239 ( \13616 , \1963 );
and \U$13240 ( \13617 , \4413 , RIc226e30_17);
not \U$13241 ( \13618 , \4413 );
and \U$13242 ( \13619 , \13618 , \1960 );
or \U$13243 ( \13620 , \13617 , \13619 );
not \U$13244 ( \13621 , \13620 );
or \U$13245 ( \13622 , \13616 , \13621 );
nand \U$13246 ( \13623 , \10584 , \1945 );
nand \U$13247 ( \13624 , \13622 , \13623 );
xor \U$13248 ( \13625 , \13615 , \13624 );
not \U$13249 ( \13626 , \2358 );
and \U$13250 ( \13627 , \5215 , \2351 );
not \U$13251 ( \13628 , \5215 );
and \U$13252 ( \13629 , \13628 , RIc226f20_15);
or \U$13253 ( \13630 , \13627 , \13629 );
not \U$13254 ( \13631 , \13630 );
or \U$13255 ( \13632 , \13626 , \13631 );
or \U$13256 ( \13633 , \10624 , \2321 );
nand \U$13257 ( \13634 , \13632 , \13633 );
xor \U$13258 ( \13635 , \13625 , \13634 );
not \U$13259 ( \13636 , \9458 );
not \U$13260 ( \13637 , \10950 );
or \U$13261 ( \13638 , \13636 , \13637 );
nand \U$13262 ( \13639 , \9444 , RIc225e40_51);
nand \U$13263 ( \13640 , \13638 , \13639 );
not \U$13264 ( \13641 , \1118 );
not \U$13265 ( \13642 , \10771 );
or \U$13266 ( \13643 , \13641 , \13642 );
and \U$13267 ( \13644 , \8829 , \1139 );
not \U$13268 ( \13645 , \8829 );
and \U$13269 ( \13646 , \13645 , RIc2272e0_7);
or \U$13270 ( \13647 , \13644 , \13646 );
nand \U$13271 ( \13648 , \13647 , \1120 );
nand \U$13272 ( \13649 , \13643 , \13648 );
xor \U$13273 ( \13650 , \13640 , \13649 );
not \U$13274 ( \13651 , \954 );
not \U$13275 ( \13652 , RIc2273d0_5);
not \U$13276 ( \13653 , \9915 );
or \U$13277 ( \13654 , \13652 , \13653 );
nand \U$13278 ( \13655 , \8951 , \935 );
nand \U$13279 ( \13656 , \13654 , \13655 );
not \U$13280 ( \13657 , \13656 );
or \U$13281 ( \13658 , \13651 , \13657 );
nand \U$13282 ( \13659 , \10752 , \950 );
nand \U$13283 ( \13660 , \13658 , \13659 );
xnor \U$13284 ( \13661 , \13650 , \13660 );
xor \U$13285 ( \13662 , \13635 , \13661 );
not \U$13286 ( \13663 , RIc2271f0_9);
not \U$13287 ( \13664 , \12228 );
or \U$13288 ( \13665 , \13663 , \13664 );
nand \U$13289 ( \13666 , \8885 , \1342 );
nand \U$13290 ( \13667 , \13665 , \13666 );
and \U$13291 ( \13668 , \13667 , \1339 );
and \U$13292 ( \13669 , \10759 , \1363 );
nor \U$13293 ( \13670 , \13668 , \13669 );
not \U$13294 ( \13671 , \1311 );
not \U$13295 ( \13672 , RIc227100_11);
not \U$13296 ( \13673 , \6719 );
or \U$13297 ( \13674 , \13672 , \13673 );
nand \U$13298 ( \13675 , \9740 , \1685 );
nand \U$13299 ( \13676 , \13674 , \13675 );
not \U$13300 ( \13677 , \13676 );
or \U$13301 ( \13678 , \13671 , \13677 );
nand \U$13302 ( \13679 , \10614 , \9904 );
nand \U$13303 ( \13680 , \13678 , \13679 );
xor \U$13304 ( \13681 , \13670 , \13680 );
not \U$13305 ( \13682 , \1678 );
not \U$13306 ( \13683 , \10634 );
or \U$13307 ( \13684 , \13682 , \13683 );
and \U$13308 ( \13685 , RIc227010_13, \6070 );
not \U$13309 ( \13686 , RIc227010_13);
not \U$13310 ( \13687 , \6070 );
and \U$13311 ( \13688 , \13686 , \13687 );
or \U$13312 ( \13689 , \13685 , \13688 );
not \U$13313 ( \13690 , \13689 );
nand \U$13314 ( \13691 , \13690 , \1682 );
nand \U$13315 ( \13692 , \13684 , \13691 );
not \U$13316 ( \13693 , \13692 );
xor \U$13317 ( \13694 , \13681 , \13693 );
xnor \U$13318 ( \13695 , \13662 , \13694 );
nand \U$13319 ( \13696 , \11272 , \11342 );
and \U$13320 ( \13697 , \13696 , \11305 );
nor \U$13321 ( \13698 , \11272 , \11342 );
nor \U$13322 ( \13699 , \13697 , \13698 );
xor \U$13323 ( \13700 , \13695 , \13699 );
xor \U$13324 ( \13701 , \10616 , \10627 );
and \U$13325 ( \13702 , \13701 , \10639 );
and \U$13326 ( \13703 , \10616 , \10627 );
or \U$13327 ( \13704 , \13702 , \13703 );
not \U$13328 ( \13705 , \11341 );
not \U$13329 ( \13706 , \11330 );
or \U$13330 ( \13707 , \13705 , \13706 );
or \U$13331 ( \13708 , \11341 , \11330 );
nand \U$13332 ( \13709 , \13708 , \11316 );
nand \U$13333 ( \13710 , \13707 , \13709 );
xor \U$13334 ( \13711 , \13704 , \13710 );
or \U$13335 ( \13712 , \10963 , \10952 );
and \U$13336 ( \13713 , \10943 , \13712 );
and \U$13337 ( \13714 , \10952 , \10963 );
nor \U$13338 ( \13715 , \13713 , \13714 );
not \U$13339 ( \13716 , \13715 );
xnor \U$13340 ( \13717 , \13711 , \13716 );
not \U$13341 ( \13718 , \13717 );
xor \U$13342 ( \13719 , \13700 , \13718 );
xor \U$13343 ( \13720 , \13614 , \13719 );
xor \U$13344 ( \13721 , \11343 , \11351 );
and \U$13345 ( \13722 , \13721 , \11443 );
and \U$13346 ( \13723 , \11343 , \11351 );
or \U$13347 ( \13724 , \13722 , \13723 );
buf \U$13348 ( \13725 , \13724 );
and \U$13349 ( \13726 , \13720 , \13725 );
not \U$13350 ( \13727 , \13720 );
not \U$13351 ( \13728 , \13725 );
and \U$13352 ( \13729 , \13727 , \13728 );
nor \U$13353 ( \13730 , \13726 , \13729 );
xnor \U$13354 ( \13731 , \13610 , \13730 );
not \U$13355 ( \13732 , \12078 );
not \U$13356 ( \13733 , \11746 );
nand \U$13357 ( \13734 , \13732 , \13733 );
not \U$13358 ( \13735 , \13734 );
not \U$13359 ( \13736 , \12278 );
or \U$13360 ( \13737 , \13735 , \13736 );
not \U$13361 ( \13738 , \13733 );
nand \U$13362 ( \13739 , \13738 , \12078 );
nand \U$13363 ( \13740 , \13737 , \13739 );
xor \U$13364 ( \13741 , \13731 , \13740 );
not \U$13365 ( \13742 , \11267 );
not \U$13366 ( \13743 , \11251 );
not \U$13367 ( \13744 , \13743 );
or \U$13368 ( \13745 , \13742 , \13744 );
or \U$13369 ( \13746 , \13743 , \11267 );
nand \U$13370 ( \13747 , \13746 , \11240 );
nand \U$13371 ( \13748 , \13745 , \13747 );
not \U$13372 ( \13749 , \10925 );
not \U$13373 ( \13750 , \10904 );
or \U$13374 ( \13751 , \13749 , \13750 );
or \U$13375 ( \13752 , \10925 , \10904 );
nand \U$13376 ( \13753 , \13752 , \10915 );
nand \U$13377 ( \13754 , \13751 , \13753 );
and \U$13378 ( \13755 , \13748 , \13754 );
not \U$13379 ( \13756 , \13748 );
not \U$13380 ( \13757 , \13754 );
and \U$13381 ( \13758 , \13756 , \13757 );
nor \U$13382 ( \13759 , \13755 , \13758 );
xor \U$13383 ( \13760 , \11282 , \11293 );
and \U$13384 ( \13761 , \13760 , \11304 );
and \U$13385 ( \13762 , \11282 , \11293 );
or \U$13386 ( \13763 , \13761 , \13762 );
and \U$13387 ( \13764 , \13759 , \13763 );
not \U$13388 ( \13765 , \13759 );
not \U$13389 ( \13766 , \13763 );
and \U$13390 ( \13767 , \13765 , \13766 );
nor \U$13391 ( \13768 , \13764 , \13767 );
not \U$13392 ( \13769 , \13768 );
not \U$13393 ( \13770 , \13769 );
not \U$13394 ( \13771 , \854 );
not \U$13395 ( \13772 , \11398 );
or \U$13396 ( \13773 , \13771 , \13772 );
and \U$13397 ( \13774 , RIc2275b0_1, \9224 );
not \U$13398 ( \13775 , RIc2275b0_1);
and \U$13399 ( \13776 , \13775 , \10644 );
or \U$13400 ( \13777 , \13774 , \13776 );
nand \U$13401 ( \13778 , \13777 , \1579 );
nand \U$13402 ( \13779 , \13773 , \13778 );
not \U$13403 ( \13780 , \2475 );
and \U$13404 ( \13781 , RIc226980_27, \13780 );
not \U$13405 ( \13782 , RIc226980_27);
and \U$13406 ( \13783 , \13782 , \2475 );
nor \U$13407 ( \13784 , \13781 , \13783 );
not \U$13408 ( \13785 , \13784 );
not \U$13409 ( \13786 , \2155 );
and \U$13410 ( \13787 , \13785 , \13786 );
and \U$13411 ( \13788 , \10923 , \2138 );
nor \U$13412 ( \13789 , \13787 , \13788 );
xor \U$13413 ( \13790 , \13779 , \13789 );
and \U$13414 ( \13791 , \10913 , \9690 );
and \U$13415 ( \13792 , \3579 , \12937 );
not \U$13416 ( \13793 , \3579 );
and \U$13417 ( \13794 , \13793 , RIc2262f0_41);
or \U$13418 ( \13795 , \13792 , \13794 );
and \U$13419 ( \13796 , \13795 , \9705 );
nor \U$13420 ( \13797 , \13791 , \13796 );
xor \U$13421 ( \13798 , \13790 , \13797 );
not \U$13422 ( \13799 , \9110 );
not \U$13423 ( \13800 , \11278 );
or \U$13424 ( \13801 , \13799 , \13800 );
not \U$13425 ( \13802 , RIc226200_43);
not \U$13426 ( \13803 , \1221 );
or \U$13427 ( \13804 , \13802 , \13803 );
not \U$13428 ( \13805 , RIc226200_43);
nand \U$13429 ( \13806 , \13805 , \1220 );
nand \U$13430 ( \13807 , \13804 , \13806 );
nand \U$13431 ( \13808 , \13807 , \9205 );
nand \U$13432 ( \13809 , \13801 , \13808 );
not \U$13433 ( \13810 , \9384 );
not \U$13434 ( \13811 , \11263 );
or \U$13435 ( \13812 , \13810 , \13811 );
not \U$13436 ( \13813 , RIc226110_45);
not \U$13437 ( \13814 , \11714 );
or \U$13438 ( \13815 , \13813 , \13814 );
nand \U$13439 ( \13816 , \2117 , \9100 );
nand \U$13440 ( \13817 , \13815 , \13816 );
nand \U$13441 ( \13818 , \13817 , \9398 );
nand \U$13442 ( \13819 , \13812 , \13818 );
xor \U$13443 ( \13820 , \13809 , \13819 );
not \U$13444 ( \13821 , \3631 );
not \U$13445 ( \13822 , RIc2266b0_33);
not \U$13446 ( \13823 , \2233 );
or \U$13447 ( \13824 , \13822 , \13823 );
nand \U$13448 ( \13825 , \2225 , \2692 );
nand \U$13449 ( \13826 , \13824 , \13825 );
not \U$13450 ( \13827 , \13826 );
or \U$13451 ( \13828 , \13821 , \13827 );
not \U$13452 ( \13829 , \11246 );
nand \U$13453 ( \13830 , \13829 , \3629 );
nand \U$13454 ( \13831 , \13828 , \13830 );
xor \U$13455 ( \13832 , \13820 , \13831 );
xor \U$13456 ( \13833 , \13798 , \13832 );
not \U$13457 ( \13834 , \2173 );
not \U$13458 ( \13835 , RIc226a70_25);
not \U$13459 ( \13836 , \2670 );
or \U$13460 ( \13837 , \13835 , \13836 );
not \U$13461 ( \13838 , RIc226a70_25);
nand \U$13462 ( \13839 , \9139 , \13838 );
nand \U$13463 ( \13840 , \13837 , \13839 );
not \U$13464 ( \13841 , \13840 );
or \U$13465 ( \13842 , \13834 , \13841 );
nand \U$13466 ( \13843 , \11362 , \2195 );
nand \U$13467 ( \13844 , \13842 , \13843 );
not \U$13468 ( \13845 , \6307 );
not \U$13469 ( \13846 , RIc2263e0_39);
not \U$13470 ( \13847 , \3044 );
or \U$13471 ( \13848 , \13846 , \13847 );
nand \U$13472 ( \13849 , \3043 , \5498 );
nand \U$13473 ( \13850 , \13848 , \13849 );
not \U$13474 ( \13851 , \13850 );
or \U$13475 ( \13852 , \13845 , \13851 );
nand \U$13476 ( \13853 , \11314 , \6688 );
nand \U$13477 ( \13854 , \13852 , \13853 );
not \U$13478 ( \13855 , \13854 );
and \U$13479 ( \13856 , \13844 , \13855 );
not \U$13480 ( \13857 , \13844 );
and \U$13481 ( \13858 , \13857 , \13854 );
or \U$13482 ( \13859 , \13856 , \13858 );
not \U$13483 ( \13860 , \1930 );
not \U$13484 ( \13861 , RIc226b60_23);
not \U$13485 ( \13862 , \5526 );
or \U$13486 ( \13863 , \13861 , \13862 );
nand \U$13487 ( \13864 , \2042 , \2111 );
nand \U$13488 ( \13865 , \13863 , \13864 );
not \U$13489 ( \13866 , \13865 );
or \U$13490 ( \13867 , \13860 , \13866 );
nand \U$13491 ( \13868 , \11339 , \1915 );
nand \U$13492 ( \13869 , \13867 , \13868 );
buf \U$13493 ( \13870 , \13869 );
and \U$13494 ( \13871 , \13859 , \13870 );
not \U$13495 ( \13872 , \13859 );
not \U$13496 ( \13873 , \13870 );
and \U$13497 ( \13874 , \13872 , \13873 );
nor \U$13498 ( \13875 , \13871 , \13874 );
xor \U$13499 ( \13876 , \13833 , \13875 );
not \U$13500 ( \13877 , \13876 );
not \U$13501 ( \13878 , \13877 );
or \U$13502 ( \13879 , \13770 , \13878 );
nand \U$13503 ( \13880 , \13876 , \13768 );
nand \U$13504 ( \13881 , \13879 , \13880 );
not \U$13505 ( \13882 , \2534 );
and \U$13506 ( \13883 , \3725 , \1941 );
not \U$13507 ( \13884 , \3725 );
and \U$13508 ( \13885 , \13884 , RIc226d40_19);
or \U$13509 ( \13886 , \13883 , \13885 );
not \U$13510 ( \13887 , \13886 );
or \U$13511 ( \13888 , \13882 , \13887 );
nand \U$13512 ( \13889 , \10593 , \2518 );
nand \U$13513 ( \13890 , \13888 , \13889 );
not \U$13514 ( \13891 , \13890 );
not \U$13515 ( \13892 , \10445 );
not \U$13516 ( \13893 , \11291 );
or \U$13517 ( \13894 , \13892 , \13893 );
not \U$13518 ( \13895 , RIc225f30_49);
not \U$13519 ( \13896 , \12472 );
or \U$13520 ( \13897 , \13895 , \13896 );
nand \U$13521 ( \13898 , \1072 , \9549 );
nand \U$13522 ( \13899 , \13897 , \13898 );
nand \U$13523 ( \13900 , \13899 , \9552 );
nand \U$13524 ( \13901 , \13894 , \13900 );
not \U$13525 ( \13902 , \13901 );
not \U$13526 ( \13903 , \13902 );
or \U$13527 ( \13904 , \13891 , \13903 );
not \U$13528 ( \13905 , \13890 );
nand \U$13529 ( \13906 , \13905 , \13901 );
nand \U$13530 ( \13907 , \13904 , \13906 );
not \U$13531 ( \13908 , \11238 );
not \U$13532 ( \13909 , \13908 );
not \U$13533 ( \13910 , \4381 );
not \U$13534 ( \13911 , \13910 );
and \U$13535 ( \13912 , \13909 , \13911 );
not \U$13536 ( \13913 , RIc2265c0_35);
not \U$13537 ( \13914 , \2421 );
not \U$13538 ( \13915 , \13914 );
or \U$13539 ( \13916 , \13913 , \13915 );
nand \U$13540 ( \13917 , \2421 , \3620 );
nand \U$13541 ( \13918 , \13916 , \13917 );
and \U$13542 ( \13919 , \13918 , \4383 );
nor \U$13543 ( \13920 , \13912 , \13919 );
not \U$13544 ( \13921 , \13920 );
not \U$13545 ( \13922 , \13921 );
and \U$13546 ( \13923 , \13907 , \13922 );
not \U$13547 ( \13924 , \13907 );
and \U$13548 ( \13925 , \13924 , \13921 );
nor \U$13549 ( \13926 , \13923 , \13925 );
not \U$13550 ( \13927 , \10001 );
not \U$13551 ( \13928 , \10959 );
or \U$13552 ( \13929 , \13927 , \13928 );
not \U$13553 ( \13930 , RIc226020_47);
not \U$13554 ( \13931 , \12537 );
or \U$13555 ( \13932 , \13930 , \13931 );
nand \U$13556 ( \13933 , \840 , \9373 );
nand \U$13557 ( \13934 , \13932 , \13933 );
nand \U$13558 ( \13935 , \13934 , \12304 );
nand \U$13559 ( \13936 , \13929 , \13935 );
not \U$13560 ( \13937 , \2078 );
not \U$13561 ( \13938 , \10902 );
or \U$13562 ( \13939 , \13937 , \13938 );
and \U$13563 ( \13940 , RIc226890_29, \12519 );
not \U$13564 ( \13941 , RIc226890_29);
and \U$13565 ( \13942 , \13941 , \2590 );
or \U$13566 ( \13943 , \13940 , \13942 );
nand \U$13567 ( \13944 , \13943 , \9142 );
nand \U$13568 ( \13945 , \13939 , \13944 );
and \U$13569 ( \13946 , \13936 , \13945 );
not \U$13570 ( \13947 , \13936 );
not \U$13571 ( \13948 , \13945 );
and \U$13572 ( \13949 , \13947 , \13948 );
nor \U$13573 ( \13950 , \13946 , \13949 );
not \U$13574 ( \13951 , RIc2267a0_31);
not \U$13575 ( \13952 , \1988 );
not \U$13576 ( \13953 , \13952 );
or \U$13577 ( \13954 , \13951 , \13953 );
not \U$13578 ( \13955 , RIc2267a0_31);
nand \U$13579 ( \13956 , \13955 , \1988 );
nand \U$13580 ( \13957 , \13954 , \13956 );
and \U$13581 ( \13958 , \13957 , \2710 );
and \U$13582 ( \13959 , \11302 , \2697 );
nor \U$13583 ( \13960 , \13958 , \13959 );
and \U$13584 ( \13961 , \13950 , \13960 );
not \U$13585 ( \13962 , \13950 );
not \U$13586 ( \13963 , \13960 );
and \U$13587 ( \13964 , \13962 , \13963 );
nor \U$13588 ( \13965 , \13961 , \13964 );
xnor \U$13589 ( \13966 , \13926 , \13965 );
not \U$13590 ( \13967 , \1082 );
not \U$13591 ( \13968 , RIc2274c0_3);
not \U$13592 ( \13969 , \8910 );
or \U$13593 ( \13970 , \13968 , \13969 );
nand \U$13594 ( \13971 , \9790 , \1032 );
nand \U$13595 ( \13972 , \13970 , \13971 );
not \U$13596 ( \13973 , \13972 );
or \U$13597 ( \13974 , \13967 , \13973 );
nand \U$13598 ( \13975 , \11410 , \1040 );
nand \U$13599 ( \13976 , \13974 , \13975 );
not \U$13600 ( \13977 , \2367 );
not \U$13601 ( \13978 , RIc226c50_21);
not \U$13602 ( \13979 , \9651 );
or \U$13603 ( \13980 , \13978 , \13979 );
nand \U$13604 ( \13981 , \4500 , \2370 );
nand \U$13605 ( \13982 , \13980 , \13981 );
not \U$13606 ( \13983 , \13982 );
or \U$13607 ( \13984 , \13977 , \13983 );
nand \U$13608 ( \13985 , \11326 , \2392 );
nand \U$13609 ( \13986 , \13984 , \13985 );
xor \U$13610 ( \13987 , \13976 , \13986 );
not \U$13611 ( \13988 , \5509 );
not \U$13612 ( \13989 , \10939 );
or \U$13613 ( \13990 , \13988 , \13989 );
and \U$13614 ( \13991 , \2353 , \5504 );
not \U$13615 ( \13992 , \2353 );
and \U$13616 ( \13993 , \13992 , RIc2264d0_37);
or \U$13617 ( \13994 , \13991 , \13993 );
nand \U$13618 ( \13995 , \13994 , \5519 );
nand \U$13619 ( \13996 , \13990 , \13995 );
xor \U$13620 ( \13997 , \13987 , \13996 );
xor \U$13621 ( \13998 , \13966 , \13997 );
and \U$13622 ( \13999 , \13881 , \13998 );
not \U$13623 ( \14000 , \13881 );
not \U$13624 ( \14001 , \13998 );
and \U$13625 ( \14002 , \14000 , \14001 );
nor \U$13626 ( \14003 , \13999 , \14002 );
not \U$13627 ( \14004 , \14003 );
not \U$13628 ( \14005 , \14004 );
not \U$13629 ( \14006 , \11020 );
not \U$13630 ( \14007 , \10965 );
nand \U$13631 ( \14008 , \14007 , \10926 );
not \U$13632 ( \14009 , \14008 );
or \U$13633 ( \14010 , \14006 , \14009 );
not \U$13634 ( \14011 , \10926 );
nand \U$13635 ( \14012 , \14011 , \10965 );
nand \U$13636 ( \14013 , \14010 , \14012 );
not \U$13637 ( \14014 , \11379 );
not \U$13638 ( \14015 , \11437 );
not \U$13639 ( \14016 , \14015 );
or \U$13640 ( \14017 , \14014 , \14016 );
not \U$13641 ( \14018 , \11437 );
not \U$13642 ( \14019 , \11378 );
or \U$13643 ( \14020 , \14018 , \14019 );
nand \U$13644 ( \14021 , \14020 , \11384 );
nand \U$13645 ( \14022 , \14017 , \14021 );
xor \U$13646 ( \14023 , \14013 , \14022 );
not \U$13647 ( \14024 , \10660 );
not \U$13648 ( \14025 , \11365 );
or \U$13649 ( \14026 , \14024 , \14025 );
nand \U$13650 ( \14027 , \14026 , \11373 );
nand \U$13651 ( \14028 , \11364 , \11353 );
nand \U$13652 ( \14029 , \14027 , \14028 );
not \U$13653 ( \14030 , \11423 );
not \U$13654 ( \14031 , \11435 );
or \U$13655 ( \14032 , \14030 , \14031 );
or \U$13656 ( \14033 , \11435 , \11423 );
nand \U$13657 ( \14034 , \14033 , \11416 );
nand \U$13658 ( \14035 , \14032 , \14034 );
xor \U$13659 ( \14036 , \14029 , \14035 );
not \U$13660 ( \14037 , \11392 );
not \U$13661 ( \14038 , \11414 );
not \U$13662 ( \14039 , \14038 );
or \U$13663 ( \14040 , \14037 , \14039 );
nand \U$13664 ( \14041 , \14040 , \11402 );
not \U$13665 ( \14042 , \11392 );
nand \U$13666 ( \14043 , \14042 , \11414 );
nand \U$13667 ( \14044 , \14041 , \14043 );
xor \U$13668 ( \14045 , \10754 , \10763 );
and \U$13669 ( \14046 , \14045 , \10773 );
and \U$13670 ( \14047 , \10754 , \10763 );
or \U$13671 ( \14048 , \14046 , \14047 );
xor \U$13672 ( \14049 , \14044 , \14048 );
xor \U$13673 ( \14050 , \10576 , \10586 );
and \U$13674 ( \14051 , \14050 , \10603 );
and \U$13675 ( \14052 , \10576 , \10586 );
or \U$13676 ( \14053 , \14051 , \14052 );
xor \U$13677 ( \14054 , \14049 , \14053 );
xor \U$13678 ( \14055 , \14036 , \14054 );
xor \U$13679 ( \14056 , \14023 , \14055 );
not \U$13680 ( \14057 , \14056 );
not \U$13681 ( \14058 , \14057 );
or \U$13682 ( \14059 , \14005 , \14058 );
nand \U$13683 ( \14060 , \14056 , \14003 );
nand \U$13684 ( \14061 , \14059 , \14060 );
not \U$13685 ( \14062 , \10042 );
not \U$13686 ( \14063 , \9525 );
or \U$13687 ( \14064 , \14062 , \14063 );
or \U$13688 ( \14065 , \9525 , \10042 );
nand \U$13689 ( \14066 , \14065 , \9968 );
nand \U$13690 ( \14067 , \14064 , \14066 );
not \U$13691 ( \14068 , \14067 );
and \U$13692 ( \14069 , \14061 , \14068 );
not \U$13693 ( \14070 , \14061 );
and \U$13694 ( \14071 , \14070 , \14067 );
nor \U$13695 ( \14072 , \14069 , \14071 );
xor \U$13696 ( \14073 , \11230 , \11444 );
and \U$13697 ( \14074 , \14073 , \11745 );
and \U$13698 ( \14075 , \11230 , \11444 );
or \U$13699 ( \14076 , \14074 , \14075 );
xor \U$13700 ( \14077 , \14072 , \14076 );
not \U$13701 ( \14078 , \10043 );
not \U$13702 ( \14079 , \10551 );
or \U$13703 ( \14080 , \14078 , \14079 );
or \U$13704 ( \14081 , \10043 , \10551 );
nand \U$13705 ( \14082 , \14081 , \11031 );
nand \U$13706 ( \14083 , \14080 , \14082 );
xnor \U$13707 ( \14084 , \14077 , \14083 );
xor \U$13708 ( \14085 , \13741 , \14084 );
not \U$13709 ( \14086 , \14085 );
not \U$13710 ( \14087 , \11032 );
nand \U$13711 ( \14088 , \14087 , \12279 );
and \U$13712 ( \14089 , \14088 , \12920 );
nor \U$13713 ( \14090 , \12279 , \14087 );
nor \U$13714 ( \14091 , \14089 , \14090 );
nand \U$13715 ( \14092 , \14086 , \14091 );
nand \U$13716 ( \14093 , \13561 , \14092 );
nand \U$13717 ( \14094 , \13719 , \13614 );
and \U$13718 ( \14095 , \13724 , \14094 );
nor \U$13719 ( \14096 , \13719 , \13614 );
nor \U$13720 ( \14097 , \14095 , \14096 );
not \U$13721 ( \14098 , \14097 );
xor \U$13722 ( \14099 , \14029 , \14035 );
and \U$13723 ( \14100 , \14099 , \14054 );
and \U$13724 ( \14101 , \14029 , \14035 );
or \U$13725 ( \14102 , \14100 , \14101 );
not \U$13726 ( \14103 , \1915 );
not \U$13727 ( \14104 , \13865 );
or \U$13728 ( \14105 , \14103 , \14104 );
not \U$13729 ( \14106 , RIc226b60_23);
not \U$13730 ( \14107 , \2063 );
or \U$13731 ( \14108 , \14106 , \14107 );
nand \U$13732 ( \14109 , \3008 , \5637 );
nand \U$13733 ( \14110 , \14108 , \14109 );
nand \U$13734 ( \14111 , \14110 , \5365 );
nand \U$13735 ( \14112 , \14105 , \14111 );
or \U$13736 ( \14113 , \9457 , \9444 );
nand \U$13737 ( \14114 , \14113 , RIc225e40_51);
and \U$13738 ( \14115 , \10653 , RIc2275b0_1);
xor \U$13739 ( \14116 , \14114 , \14115 );
not \U$13740 ( \14117 , \1579 );
xor \U$13741 ( \14118 , RIc2275b0_1, \8924 );
not \U$13742 ( \14119 , \14118 );
or \U$13743 ( \14120 , \14117 , \14119 );
nand \U$13744 ( \14121 , \13777 , \854 );
nand \U$13745 ( \14122 , \14120 , \14121 );
xor \U$13746 ( \14123 , \14116 , \14122 );
not \U$13747 ( \14124 , \14123 );
xor \U$13748 ( \14125 , \14112 , \14124 );
xor \U$13749 ( \14126 , \13615 , \13624 );
and \U$13750 ( \14127 , \14126 , \13634 );
and \U$13751 ( \14128 , \13615 , \13624 );
or \U$13752 ( \14129 , \14127 , \14128 );
xnor \U$13753 ( \14130 , \14125 , \14129 );
not \U$13754 ( \14131 , \13635 );
nand \U$13755 ( \14132 , \13661 , \14131 );
and \U$13756 ( \14133 , \14132 , \13694 );
nor \U$13757 ( \14134 , \13661 , \14131 );
nor \U$13758 ( \14135 , \14133 , \14134 );
not \U$13759 ( \14136 , \14135 );
xor \U$13760 ( \14137 , \14130 , \14136 );
or \U$13761 ( \14138 , \13748 , \13754 );
nand \U$13762 ( \14139 , \14138 , \13763 );
nand \U$13763 ( \14140 , \13748 , \13754 );
nand \U$13764 ( \14141 , \14139 , \14140 );
xnor \U$13765 ( \14142 , \14137 , \14141 );
xor \U$13766 ( \14143 , \14102 , \14142 );
not \U$13767 ( \14144 , \13699 );
not \U$13768 ( \14145 , \14144 );
not \U$13769 ( \14146 , \13718 );
or \U$13770 ( \14147 , \14145 , \14146 );
not \U$13771 ( \14148 , \13699 );
not \U$13772 ( \14149 , \13717 );
or \U$13773 ( \14150 , \14148 , \14149 );
nand \U$13774 ( \14151 , \14150 , \13695 );
nand \U$13775 ( \14152 , \14147 , \14151 );
xor \U$13776 ( \14153 , \14143 , \14152 );
not \U$13777 ( \14154 , \14153 );
and \U$13778 ( \14155 , \14098 , \14154 );
not \U$13779 ( \14156 , \14098 );
and \U$13780 ( \14157 , \14156 , \14153 );
nor \U$13781 ( \14158 , \14155 , \14157 );
not \U$13782 ( \14159 , \13704 );
nand \U$13783 ( \14160 , \14159 , \13715 );
not \U$13784 ( \14161 , \14160 );
not \U$13785 ( \14162 , \13710 );
or \U$13786 ( \14163 , \14161 , \14162 );
nand \U$13787 ( \14164 , \13716 , \13704 );
nand \U$13788 ( \14165 , \14163 , \14164 );
nand \U$13789 ( \14166 , \13965 , \13926 );
and \U$13790 ( \14167 , \14166 , \13997 );
nor \U$13791 ( \14168 , \13965 , \13926 );
nor \U$13792 ( \14169 , \14167 , \14168 );
not \U$13793 ( \14170 , \14169 );
xor \U$13794 ( \14171 , \14165 , \14170 );
not \U$13795 ( \14172 , \13798 );
or \U$13796 ( \14173 , \14172 , \13832 );
nand \U$13797 ( \14174 , \14173 , \13875 );
nand \U$13798 ( \14175 , \13832 , \14172 );
nand \U$13799 ( \14176 , \14174 , \14175 );
xor \U$13800 ( \14177 , \14171 , \14176 );
not \U$13801 ( \14178 , \14001 );
not \U$13802 ( \14179 , \13768 );
or \U$13803 ( \14180 , \14178 , \14179 );
not \U$13804 ( \14181 , \13769 );
not \U$13805 ( \14182 , \13998 );
or \U$13806 ( \14183 , \14181 , \14182 );
not \U$13807 ( \14184 , \13876 );
nand \U$13808 ( \14185 , \14183 , \14184 );
nand \U$13809 ( \14186 , \14180 , \14185 );
xor \U$13810 ( \14187 , \14177 , \14186 );
not \U$13811 ( \14188 , \1307 );
not \U$13812 ( \14189 , \13676 );
or \U$13813 ( \14190 , \14188 , \14189 );
not \U$13814 ( \14191 , RIc227100_11);
not \U$13815 ( \14192 , \6492 );
not \U$13816 ( \14193 , \14192 );
or \U$13817 ( \14194 , \14191 , \14193 );
nand \U$13818 ( \14195 , \6492 , \3351 );
nand \U$13819 ( \14196 , \14194 , \14195 );
nand \U$13820 ( \14197 , \14196 , \1311 );
nand \U$13821 ( \14198 , \14190 , \14197 );
not \U$13822 ( \14199 , \1120 );
and \U$13823 ( \14200 , \8856 , \1139 );
not \U$13824 ( \14201 , \8856 );
and \U$13825 ( \14202 , \14201 , RIc2272e0_7);
or \U$13826 ( \14203 , \14200 , \14202 );
not \U$13827 ( \14204 , \14203 );
or \U$13828 ( \14205 , \14199 , \14204 );
nand \U$13829 ( \14206 , \13647 , \1118 );
nand \U$13830 ( \14207 , \14205 , \14206 );
not \U$13831 ( \14208 , \14207 );
and \U$13832 ( \14209 , \14198 , \14208 );
not \U$13833 ( \14210 , \14198 );
and \U$13834 ( \14211 , \14210 , \14207 );
or \U$13835 ( \14212 , \14209 , \14211 );
not \U$13836 ( \14213 , \1363 );
not \U$13837 ( \14214 , \13667 );
or \U$13838 ( \14215 , \14213 , \14214 );
not \U$13839 ( \14216 , RIc2271f0_9);
not \U$13840 ( \14217 , \9728 );
or \U$13841 ( \14218 , \14216 , \14217 );
nand \U$13842 ( \14219 , \9731 , \1342 );
nand \U$13843 ( \14220 , \14218 , \14219 );
nand \U$13844 ( \14221 , \14220 , \1340 );
nand \U$13845 ( \14222 , \14215 , \14221 );
not \U$13846 ( \14223 , \14222 );
and \U$13847 ( \14224 , \14212 , \14223 );
not \U$13848 ( \14225 , \14212 );
and \U$13849 ( \14226 , \14225 , \14222 );
nor \U$13850 ( \14227 , \14224 , \14226 );
not \U$13851 ( \14228 , \14227 );
not \U$13852 ( \14229 , \1040 );
not \U$13853 ( \14230 , \13972 );
or \U$13854 ( \14231 , \14229 , \14230 );
not \U$13855 ( \14232 , RIc2274c0_3);
not \U$13856 ( \14233 , \11094 );
or \U$13857 ( \14234 , \14232 , \14233 );
nand \U$13858 ( \14235 , \8979 , \1032 );
nand \U$13859 ( \14236 , \14234 , \14235 );
nand \U$13860 ( \14237 , \14236 , \1082 );
nand \U$13861 ( \14238 , \14231 , \14237 );
not \U$13862 ( \14239 , \950 );
not \U$13863 ( \14240 , \13656 );
or \U$13864 ( \14241 , \14239 , \14240 );
and \U$13865 ( \14242 , \8806 , \946 );
not \U$13866 ( \14243 , \8806 );
and \U$13867 ( \14244 , \14243 , RIc2273d0_5);
or \U$13868 ( \14245 , \14242 , \14244 );
nand \U$13869 ( \14246 , \14245 , \954 );
nand \U$13870 ( \14247 , \14241 , \14246 );
not \U$13871 ( \14248 , \14247 );
xor \U$13872 ( \14249 , \14238 , \14248 );
not \U$13873 ( \14250 , \5509 );
not \U$13874 ( \14251 , \13994 );
or \U$13875 ( \14252 , \14250 , \14251 );
not \U$13876 ( \14253 , RIc2264d0_37);
not \U$13877 ( \14254 , \4177 );
or \U$13878 ( \14255 , \14253 , \14254 );
nand \U$13879 ( \14256 , \1729 , \5504 );
nand \U$13880 ( \14257 , \14255 , \14256 );
nand \U$13881 ( \14258 , \14257 , \5519 );
nand \U$13882 ( \14259 , \14252 , \14258 );
xor \U$13883 ( \14260 , \14249 , \14259 );
not \U$13884 ( \14261 , \14260 );
not \U$13885 ( \14262 , \14261 );
or \U$13886 ( \14263 , \14228 , \14262 );
not \U$13887 ( \14264 , \14227 );
nand \U$13888 ( \14265 , \14264 , \14260 );
nand \U$13889 ( \14266 , \14263 , \14265 );
not \U$13890 ( \14267 , \2078 );
not \U$13891 ( \14268 , \13943 );
or \U$13892 ( \14269 , \14267 , \14268 );
xor \U$13893 ( \14270 , RIc226890_29, \2013 );
nand \U$13894 ( \14271 , \14270 , \9142 );
nand \U$13895 ( \14272 , \14269 , \14271 );
not \U$13896 ( \14273 , RIc226980_27);
not \U$13897 ( \14274 , \4802 );
or \U$13898 ( \14275 , \14273 , \14274 );
not \U$13899 ( \14276 , RIc226980_27);
nand \U$13900 ( \14277 , \14276 , \3446 );
nand \U$13901 ( \14278 , \14275 , \14277 );
not \U$13902 ( \14279 , \14278 );
not \U$13903 ( \14280 , \2154 );
or \U$13904 ( \14281 , \14279 , \14280 );
not \U$13905 ( \14282 , \13784 );
nand \U$13906 ( \14283 , \14282 , \2138 );
nand \U$13907 ( \14284 , \14281 , \14283 );
xor \U$13908 ( \14285 , \14272 , \14284 );
not \U$13909 ( \14286 , \9816 );
and \U$13910 ( \14287 , \1392 , RIc2262f0_41);
not \U$13911 ( \14288 , \1392 );
and \U$13912 ( \14289 , \14288 , \6303 );
or \U$13913 ( \14290 , \14287 , \14289 );
not \U$13914 ( \14291 , \14290 );
or \U$13915 ( \14292 , \14286 , \14291 );
nand \U$13916 ( \14293 , \13795 , \9690 );
nand \U$13917 ( \14294 , \14292 , \14293 );
xor \U$13918 ( \14295 , \14285 , \14294 );
xor \U$13919 ( \14296 , \14266 , \14295 );
not \U$13920 ( \14297 , \1963 );
not \U$13921 ( \14298 , RIc226e30_17);
not \U$13922 ( \14299 , \3640 );
not \U$13923 ( \14300 , \14299 );
or \U$13924 ( \14301 , \14298 , \14300 );
nand \U$13925 ( \14302 , \3640 , \1960 );
nand \U$13926 ( \14303 , \14301 , \14302 );
not \U$13927 ( \14304 , \14303 );
or \U$13928 ( \14305 , \14297 , \14304 );
nand \U$13929 ( \14306 , \13620 , \1945 );
nand \U$13930 ( \14307 , \14305 , \14306 );
not \U$13931 ( \14308 , \14307 );
not \U$13932 ( \14309 , \2358 );
and \U$13933 ( \14310 , RIc226f20_15, \10277 );
not \U$13934 ( \14311 , RIc226f20_15);
and \U$13935 ( \14312 , \14311 , \4406 );
or \U$13936 ( \14313 , \14310 , \14312 );
not \U$13937 ( \14314 , \14313 );
or \U$13938 ( \14315 , \14309 , \14314 );
nand \U$13939 ( \14316 , \13630 , \2320 );
nand \U$13940 ( \14317 , \14315 , \14316 );
not \U$13941 ( \14318 , \14317 );
not \U$13942 ( \14319 , \14318 );
or \U$13943 ( \14320 , \14308 , \14319 );
or \U$13944 ( \14321 , \14307 , \14318 );
nand \U$13945 ( \14322 , \14320 , \14321 );
not \U$13946 ( \14323 , \13689 );
not \U$13947 ( \14324 , \1679 );
and \U$13948 ( \14325 , \14323 , \14324 );
and \U$13949 ( \14326 , \5663 , \1296 );
not \U$13950 ( \14327 , \5663 );
and \U$13951 ( \14328 , \14327 , RIc227010_13);
or \U$13952 ( \14329 , \14326 , \14328 );
and \U$13953 ( \14330 , \14329 , \1682 );
nor \U$13954 ( \14331 , \14325 , \14330 );
not \U$13955 ( \14332 , \14331 );
and \U$13956 ( \14333 , \14322 , \14332 );
not \U$13957 ( \14334 , \14322 );
not \U$13958 ( \14335 , \14332 );
and \U$13959 ( \14336 , \14334 , \14335 );
nor \U$13960 ( \14337 , \14333 , \14336 );
xor \U$13961 ( \14338 , \13779 , \13789 );
and \U$13962 ( \14339 , \14338 , \13797 );
and \U$13963 ( \14340 , \13779 , \13789 );
or \U$13964 ( \14341 , \14339 , \14340 );
not \U$13965 ( \14342 , \14341 );
xor \U$13966 ( \14343 , \14337 , \14342 );
nor \U$13967 ( \14344 , \13844 , \13869 );
or \U$13968 ( \14345 , \14344 , \13855 );
nand \U$13969 ( \14346 , \13844 , \13869 );
nand \U$13970 ( \14347 , \14345 , \14346 );
xor \U$13971 ( \14348 , \14343 , \14347 );
xor \U$13972 ( \14349 , \14296 , \14348 );
not \U$13973 ( \14350 , \13901 );
not \U$13974 ( \14351 , \13921 );
or \U$13975 ( \14352 , \14350 , \14351 );
not \U$13976 ( \14353 , \13902 );
not \U$13977 ( \14354 , \13920 );
or \U$13978 ( \14355 , \14353 , \14354 );
nand \U$13979 ( \14356 , \14355 , \13890 );
nand \U$13980 ( \14357 , \14352 , \14356 );
not \U$13981 ( \14358 , \13945 );
not \U$13982 ( \14359 , \13963 );
or \U$13983 ( \14360 , \14358 , \14359 );
not \U$13984 ( \14361 , \13960 );
not \U$13985 ( \14362 , \13948 );
or \U$13986 ( \14363 , \14361 , \14362 );
nand \U$13987 ( \14364 , \14363 , \13936 );
nand \U$13988 ( \14365 , \14360 , \14364 );
xor \U$13989 ( \14366 , \14357 , \14365 );
xor \U$13990 ( \14367 , \13809 , \13819 );
and \U$13991 ( \14368 , \14367 , \13831 );
and \U$13992 ( \14369 , \13809 , \13819 );
or \U$13993 ( \14370 , \14368 , \14369 );
xor \U$13994 ( \14371 , \14366 , \14370 );
xor \U$13995 ( \14372 , \14349 , \14371 );
xor \U$13996 ( \14373 , \14187 , \14372 );
xnor \U$13997 ( \14374 , \14158 , \14373 );
buf \U$13998 ( \14375 , \14004 );
or \U$13999 ( \14376 , \14375 , \14067 );
nand \U$14000 ( \14377 , \14376 , \14056 );
nand \U$14001 ( \14378 , \14067 , \14375 );
nand \U$14002 ( \14379 , \14377 , \14378 );
not \U$14003 ( \14380 , \14379 );
not \U$14004 ( \14381 , \14380 );
xor \U$14005 ( \14382 , \14013 , \14022 );
and \U$14006 ( \14383 , \14382 , \14055 );
and \U$14007 ( \14384 , \14013 , \14022 );
or \U$14008 ( \14385 , \14383 , \14384 );
not \U$14009 ( \14386 , \9398 );
not \U$14010 ( \14387 , RIc226110_45);
not \U$14011 ( \14388 , \1557 );
or \U$14012 ( \14389 , \14387 , \14388 );
not \U$14013 ( \14390 , RIc226110_45);
nand \U$14014 ( \14391 , \980 , \14390 );
nand \U$14015 ( \14392 , \14389 , \14391 );
not \U$14016 ( \14393 , \14392 );
or \U$14017 ( \14394 , \14386 , \14393 );
nand \U$14018 ( \14395 , \13817 , \9934 );
nand \U$14019 ( \14396 , \14394 , \14395 );
not \U$14020 ( \14397 , \4381 );
not \U$14021 ( \14398 , \13918 );
or \U$14022 ( \14399 , \14397 , \14398 );
not \U$14023 ( \14400 , RIc2265c0_35);
not \U$14024 ( \14401 , \3092 );
or \U$14025 ( \14402 , \14400 , \14401 );
nand \U$14026 ( \14403 , \8989 , \4376 );
nand \U$14027 ( \14404 , \14402 , \14403 );
nand \U$14028 ( \14405 , \14404 , \4383 );
nand \U$14029 ( \14406 , \14399 , \14405 );
xor \U$14030 ( \14407 , \14396 , \14406 );
not \U$14031 ( \14408 , \3629 );
not \U$14032 ( \14409 , \13826 );
or \U$14033 ( \14410 , \14408 , \14409 );
not \U$14034 ( \14411 , RIc2266b0_33);
not \U$14035 ( \14412 , \9570 );
or \U$14036 ( \14413 , \14411 , \14412 );
nand \U$14037 ( \14414 , \2443 , \5179 );
nand \U$14038 ( \14415 , \14413 , \14414 );
nand \U$14039 ( \14416 , \14415 , \3631 );
nand \U$14040 ( \14417 , \14410 , \14416 );
xor \U$14041 ( \14418 , \14407 , \14417 );
not \U$14042 ( \14419 , \9205 );
not \U$14043 ( \14420 , RIc226200_43);
not \U$14044 ( \14421 , \1169 );
not \U$14045 ( \14422 , \14421 );
or \U$14046 ( \14423 , \14420 , \14422 );
nand \U$14047 ( \14424 , \1169 , \9117 );
nand \U$14048 ( \14425 , \14423 , \14424 );
not \U$14049 ( \14426 , \14425 );
or \U$14050 ( \14427 , \14419 , \14426 );
nand \U$14051 ( \14428 , \13807 , \9110 );
nand \U$14052 ( \14429 , \14427 , \14428 );
not \U$14053 ( \14430 , \9619 );
not \U$14054 ( \14431 , RIc226020_47);
not \U$14055 ( \14432 , \13077 );
or \U$14056 ( \14433 , \14431 , \14432 );
nand \U$14057 ( \14434 , \888 , \9624 );
nand \U$14058 ( \14435 , \14433 , \14434 );
not \U$14059 ( \14436 , \14435 );
or \U$14060 ( \14437 , \14430 , \14436 );
nand \U$14061 ( \14438 , \13934 , \9639 );
nand \U$14062 ( \14439 , \14437 , \14438 );
xor \U$14063 ( \14440 , \14429 , \14439 );
not \U$14064 ( \14441 , \2710 );
not \U$14065 ( \14442 , RIc2267a0_31);
not \U$14066 ( \14443 , \2257 );
or \U$14067 ( \14444 , \14442 , \14443 );
nand \U$14068 ( \14445 , \4008 , \3648 );
nand \U$14069 ( \14446 , \14444 , \14445 );
not \U$14070 ( \14447 , \14446 );
or \U$14071 ( \14448 , \14441 , \14447 );
nand \U$14072 ( \14449 , \13957 , \2697 );
nand \U$14073 ( \14450 , \14448 , \14449 );
xor \U$14074 ( \14451 , \14440 , \14450 );
xor \U$14075 ( \14452 , \14418 , \14451 );
not \U$14076 ( \14453 , \10445 );
not \U$14077 ( \14454 , \13899 );
or \U$14078 ( \14455 , \14453 , \14454 );
not \U$14079 ( \14456 , \9541 );
not \U$14080 ( \14457 , \930 );
or \U$14081 ( \14458 , \14456 , \14457 );
nand \U$14082 ( \14459 , \11112 , RIc225f30_49);
nand \U$14083 ( \14460 , \14458 , \14459 );
nand \U$14084 ( \14461 , \9552 , \14460 );
nand \U$14085 ( \14462 , \14455 , \14461 );
not \U$14086 ( \14463 , \2518 );
not \U$14087 ( \14464 , \13886 );
or \U$14088 ( \14465 , \14463 , \14464 );
not \U$14089 ( \14466 , RIc226d40_19);
not \U$14090 ( \14467 , \13102 );
or \U$14091 ( \14468 , \14466 , \14467 );
nand \U$14092 ( \14469 , \3115 , \3338 );
nand \U$14093 ( \14470 , \14468 , \14469 );
nand \U$14094 ( \14471 , \14470 , \2534 );
nand \U$14095 ( \14472 , \14465 , \14471 );
xor \U$14096 ( \14473 , \14462 , \14472 );
not \U$14097 ( \14474 , \2367 );
not \U$14098 ( \14475 , RIc226c50_21);
not \U$14099 ( \14476 , \2634 );
not \U$14100 ( \14477 , \14476 );
or \U$14101 ( \14478 , \14475 , \14477 );
nand \U$14102 ( \14479 , \2634 , \2383 );
nand \U$14103 ( \14480 , \14478 , \14479 );
not \U$14104 ( \14481 , \14480 );
or \U$14105 ( \14482 , \14474 , \14481 );
nand \U$14106 ( \14483 , \13982 , \2392 );
nand \U$14107 ( \14484 , \14482 , \14483 );
xor \U$14108 ( \14485 , \14473 , \14484 );
xor \U$14109 ( \14486 , \14452 , \14485 );
not \U$14110 ( \14487 , \13588 );
not \U$14111 ( \14488 , \13584 );
or \U$14112 ( \14489 , \14487 , \14488 );
or \U$14113 ( \14490 , \13584 , \13588 );
nand \U$14114 ( \14491 , \14490 , \13594 );
nand \U$14115 ( \14492 , \14489 , \14491 );
xor \U$14116 ( \14493 , \14486 , \14492 );
not \U$14117 ( \14494 , \6689 );
not \U$14118 ( \14495 , \13850 );
or \U$14119 ( \14496 , \14494 , \14495 );
not \U$14120 ( \14497 , RIc2263e0_39);
not \U$14121 ( \14498 , \1948 );
or \U$14122 ( \14499 , \14497 , \14498 );
not \U$14123 ( \14500 , RIc2263e0_39);
nand \U$14124 ( \14501 , \14500 , \1331 );
nand \U$14125 ( \14502 , \14499 , \14501 );
nand \U$14126 ( \14503 , \14502 , \6307 );
nand \U$14127 ( \14504 , \14496 , \14503 );
xor \U$14128 ( \14505 , \13779 , \14504 );
not \U$14129 ( \14506 , RIc226a70_25);
not \U$14130 ( \14507 , \4195 );
or \U$14131 ( \14508 , \14506 , \14507 );
nand \U$14132 ( \14509 , \2498 , \1905 );
nand \U$14133 ( \14510 , \14508 , \14509 );
not \U$14134 ( \14511 , \14510 );
not \U$14135 ( \14512 , \14511 );
not \U$14136 ( \14513 , \2171 );
and \U$14137 ( \14514 , \14512 , \14513 );
and \U$14138 ( \14515 , \13840 , \2195 );
nor \U$14139 ( \14516 , \14514 , \14515 );
not \U$14140 ( \14517 , \14516 );
xnor \U$14141 ( \14518 , \14505 , \14517 );
xor \U$14142 ( \14519 , \14044 , \14048 );
and \U$14143 ( \14520 , \14519 , \14053 );
and \U$14144 ( \14521 , \14044 , \14048 );
or \U$14145 ( \14522 , \14520 , \14521 );
xor \U$14146 ( \14523 , \14518 , \14522 );
or \U$14147 ( \14524 , \13640 , \13660 );
nand \U$14148 ( \14525 , \14524 , \13649 );
nand \U$14149 ( \14526 , \13660 , \13640 );
nand \U$14150 ( \14527 , \14525 , \14526 );
not \U$14151 ( \14528 , \13670 );
not \U$14152 ( \14529 , \13693 );
or \U$14153 ( \14530 , \14528 , \14529 );
nand \U$14154 ( \14531 , \14530 , \13680 );
not \U$14155 ( \14532 , \13670 );
nand \U$14156 ( \14533 , \14532 , \13692 );
nand \U$14157 ( \14534 , \14531 , \14533 );
xor \U$14158 ( \14535 , \14527 , \14534 );
not \U$14159 ( \14536 , \13976 );
not \U$14160 ( \14537 , \13986 );
or \U$14161 ( \14538 , \14536 , \14537 );
or \U$14162 ( \14539 , \13986 , \13976 );
nand \U$14163 ( \14540 , \14539 , \13996 );
nand \U$14164 ( \14541 , \14538 , \14540 );
xor \U$14165 ( \14542 , \14535 , \14541 );
xnor \U$14166 ( \14543 , \14523 , \14542 );
xnor \U$14167 ( \14544 , \14493 , \14543 );
not \U$14168 ( \14545 , \14544 );
xor \U$14169 ( \14546 , \14385 , \14545 );
not \U$14170 ( \14547 , \13567 );
not \U$14171 ( \14548 , \13598 );
or \U$14172 ( \14549 , \14547 , \14548 );
not \U$14173 ( \14550 , \13595 );
not \U$14174 ( \14551 , \13568 );
or \U$14175 ( \14552 , \14550 , \14551 );
nand \U$14176 ( \14553 , \14552 , \13576 );
nand \U$14177 ( \14554 , \14549 , \14553 );
not \U$14178 ( \14555 , \14554 );
xnor \U$14179 ( \14556 , \14546 , \14555 );
not \U$14180 ( \14557 , \14556 );
or \U$14181 ( \14558 , \14381 , \14557 );
or \U$14182 ( \14559 , \14380 , \14556 );
nand \U$14183 ( \14560 , \14558 , \14559 );
not \U$14184 ( \14561 , \13609 );
not \U$14185 ( \14562 , \13600 );
not \U$14186 ( \14563 , \14562 );
or \U$14187 ( \14564 , \14561 , \14563 );
or \U$14188 ( \14565 , \13609 , \14562 );
nand \U$14189 ( \14566 , \14565 , \13730 );
nand \U$14190 ( \14567 , \14564 , \14566 );
not \U$14191 ( \14568 , \14567 );
and \U$14192 ( \14569 , \14560 , \14568 );
not \U$14193 ( \14570 , \14560 );
and \U$14194 ( \14571 , \14570 , \14567 );
nor \U$14195 ( \14572 , \14569 , \14571 );
xor \U$14196 ( \14573 , \14374 , \14572 );
not \U$14197 ( \14574 , \14076 );
buf \U$14198 ( \14575 , \14072 );
nand \U$14199 ( \14576 , \14574 , \14575 );
buf \U$14200 ( \14577 , \14083 );
and \U$14201 ( \14578 , \14576 , \14577 );
nor \U$14202 ( \14579 , \14574 , \14575 );
nor \U$14203 ( \14580 , \14578 , \14579 );
and \U$14204 ( \14581 , \14573 , \14580 );
and \U$14205 ( \14582 , \14374 , \14572 );
or \U$14206 ( \14583 , \14581 , \14582 );
nand \U$14207 ( \14584 , \14097 , \14153 );
not \U$14208 ( \14585 , \14584 );
not \U$14209 ( \14586 , \14373 );
or \U$14210 ( \14587 , \14585 , \14586 );
nand \U$14211 ( \14588 , \14098 , \14154 );
nand \U$14212 ( \14589 , \14587 , \14588 );
not \U$14213 ( \14590 , \14589 );
not \U$14214 ( \14591 , \14590 );
not \U$14215 ( \14592 , \14385 );
nand \U$14216 ( \14593 , \14592 , \14544 );
not \U$14217 ( \14594 , \14593 );
not \U$14218 ( \14595 , \14554 );
or \U$14219 ( \14596 , \14594 , \14595 );
not \U$14220 ( \14597 , \14544 );
nand \U$14221 ( \14598 , \14597 , \14385 );
nand \U$14222 ( \14599 , \14596 , \14598 );
not \U$14223 ( \14600 , \14599 );
not \U$14224 ( \14601 , \14543 );
buf \U$14225 ( \14602 , \14486 );
not \U$14226 ( \14603 , \14602 );
or \U$14227 ( \14604 , \14601 , \14603 );
or \U$14228 ( \14605 , \14602 , \14543 );
nand \U$14229 ( \14606 , \14605 , \14492 );
nand \U$14230 ( \14607 , \14604 , \14606 );
not \U$14231 ( \14608 , \9046 );
nand \U$14232 ( \14609 , \14608 , RIc2275b0_1);
not \U$14233 ( \14610 , \2697 );
not \U$14234 ( \14611 , \14446 );
or \U$14235 ( \14612 , \14610 , \14611 );
and \U$14236 ( \14613 , RIc2267a0_31, \2226 );
not \U$14237 ( \14614 , RIc2267a0_31);
and \U$14238 ( \14615 , \14614 , \2225 );
or \U$14239 ( \14616 , \14613 , \14615 );
nand \U$14240 ( \14617 , \14616 , \2710 );
nand \U$14241 ( \14618 , \14612 , \14617 );
xor \U$14242 ( \14619 , \14609 , \14618 );
not \U$14243 ( \14620 , \9690 );
not \U$14244 ( \14621 , \14290 );
or \U$14245 ( \14622 , \14620 , \14621 );
not \U$14246 ( \14623 , RIc2262f0_41);
not \U$14247 ( \14624 , \1222 );
or \U$14248 ( \14625 , \14623 , \14624 );
nand \U$14249 ( \14626 , \1370 , \6303 );
nand \U$14250 ( \14627 , \14625 , \14626 );
nand \U$14251 ( \14628 , \14627 , \9705 );
nand \U$14252 ( \14629 , \14622 , \14628 );
xor \U$14253 ( \14630 , \14619 , \14629 );
not \U$14254 ( \14631 , \2784 );
not \U$14255 ( \14632 , \14270 );
or \U$14256 ( \14633 , \14631 , \14632 );
not \U$14257 ( \14634 , RIc226890_29);
not \U$14258 ( \14635 , \1988 );
not \U$14259 ( \14636 , \14635 );
or \U$14260 ( \14637 , \14634 , \14636 );
not \U$14261 ( \14638 , RIc226890_29);
nand \U$14262 ( \14639 , \14638 , \1988 );
nand \U$14263 ( \14640 , \14637 , \14639 );
nand \U$14264 ( \14641 , \14640 , \9142 );
nand \U$14265 ( \14642 , \14633 , \14641 );
not \U$14266 ( \14643 , \2138 );
not \U$14267 ( \14644 , \14278 );
or \U$14268 ( \14645 , \14643 , \14644 );
and \U$14269 ( \14646 , RIc226980_27, \2591 );
not \U$14270 ( \14647 , RIc226980_27);
and \U$14271 ( \14648 , \14647 , \2590 );
or \U$14272 ( \14649 , \14646 , \14648 );
nand \U$14273 ( \14650 , \14649 , \2154 );
nand \U$14274 ( \14651 , \14645 , \14650 );
xor \U$14275 ( \14652 , \14642 , \14651 );
not \U$14276 ( \14653 , \9384 );
not \U$14277 ( \14654 , \14392 );
or \U$14278 ( \14655 , \14653 , \14654 );
not \U$14279 ( \14656 , RIc226110_45);
not \U$14280 ( \14657 , \10450 );
or \U$14281 ( \14658 , \14656 , \14657 );
not \U$14282 ( \14659 , \12537 );
not \U$14283 ( \14660 , RIc226110_45);
nand \U$14284 ( \14661 , \14659 , \14660 );
nand \U$14285 ( \14662 , \14658 , \14661 );
nand \U$14286 ( \14663 , \14662 , \9398 );
nand \U$14287 ( \14664 , \14655 , \14663 );
xor \U$14288 ( \14665 , \14652 , \14664 );
xor \U$14289 ( \14666 , \14630 , \14665 );
not \U$14290 ( \14667 , \9619 );
not \U$14291 ( \14668 , RIc226020_47);
not \U$14292 ( \14669 , \12472 );
or \U$14293 ( \14670 , \14668 , \14669 );
nand \U$14294 ( \14671 , \1072 , \9373 );
nand \U$14295 ( \14672 , \14670 , \14671 );
not \U$14296 ( \14673 , \14672 );
or \U$14297 ( \14674 , \14667 , \14673 );
nand \U$14298 ( \14675 , \14435 , \10001 );
nand \U$14299 ( \14676 , \14674 , \14675 );
not \U$14300 ( \14677 , \9110 );
not \U$14301 ( \14678 , \14425 );
or \U$14302 ( \14679 , \14677 , \14678 );
not \U$14303 ( \14680 , RIc226200_43);
not \U$14304 ( \14681 , \4432 );
or \U$14305 ( \14682 , \14680 , \14681 );
nand \U$14306 ( \14683 , \1020 , \9106 );
nand \U$14307 ( \14684 , \14682 , \14683 );
nand \U$14308 ( \14685 , \14684 , \9129 );
nand \U$14309 ( \14686 , \14679 , \14685 );
xor \U$14310 ( \14687 , \14676 , \14686 );
not \U$14311 ( \14688 , \3631 );
not \U$14312 ( \14689 , RIc2266b0_33);
not \U$14313 ( \14690 , \3686 );
or \U$14314 ( \14691 , \14689 , \14690 );
nand \U$14315 ( \14692 , \2422 , \9943 );
nand \U$14316 ( \14693 , \14691 , \14692 );
not \U$14317 ( \14694 , \14693 );
or \U$14318 ( \14695 , \14688 , \14694 );
nand \U$14319 ( \14696 , \14415 , \3629 );
nand \U$14320 ( \14697 , \14695 , \14696 );
xor \U$14321 ( \14698 , \14687 , \14697 );
xor \U$14322 ( \14699 , \14666 , \14698 );
not \U$14323 ( \14700 , \14699 );
not \U$14324 ( \14701 , \14700 );
not \U$14325 ( \14702 , \14129 );
not \U$14326 ( \14703 , \14112 );
or \U$14327 ( \14704 , \14702 , \14703 );
or \U$14328 ( \14705 , \14129 , \14112 );
nand \U$14329 ( \14706 , \14705 , \14123 );
nand \U$14330 ( \14707 , \14704 , \14706 );
xor \U$14331 ( \14708 , \14114 , \14115 );
and \U$14332 ( \14709 , \14708 , \14122 );
and \U$14333 ( \14710 , \14114 , \14115 );
or \U$14334 ( \14711 , \14709 , \14710 );
not \U$14335 ( \14712 , \1915 );
not \U$14336 ( \14713 , \14110 );
or \U$14337 ( \14714 , \14712 , \14713 );
not \U$14338 ( \14715 , RIc226b60_23);
not \U$14339 ( \14716 , \12548 );
or \U$14340 ( \14717 , \14715 , \14716 );
nand \U$14341 ( \14718 , \2720 , \10210 );
nand \U$14342 ( \14719 , \14717 , \14718 );
nand \U$14343 ( \14720 , \14719 , \5365 );
nand \U$14344 ( \14721 , \14714 , \14720 );
xor \U$14345 ( \14722 , \14711 , \14721 );
not \U$14346 ( \14723 , \2392 );
not \U$14347 ( \14724 , \14480 );
or \U$14348 ( \14725 , \14723 , \14724 );
not \U$14349 ( \14726 , RIc226c50_21);
not \U$14350 ( \14727 , \3798 );
or \U$14351 ( \14728 , \14726 , \14727 );
nand \U$14352 ( \14729 , \2042 , \2383 );
nand \U$14353 ( \14730 , \14728 , \14729 );
nand \U$14354 ( \14731 , \14730 , \2367 );
nand \U$14355 ( \14732 , \14725 , \14731 );
xor \U$14356 ( \14733 , \14722 , \14732 );
xor \U$14357 ( \14734 , \14707 , \14733 );
not \U$14358 ( \14735 , \4381 );
not \U$14359 ( \14736 , \14404 );
or \U$14360 ( \14737 , \14735 , \14736 );
not \U$14361 ( \14738 , RIc2265c0_35);
not \U$14362 ( \14739 , \9700 );
or \U$14363 ( \14740 , \14738 , \14739 );
nand \U$14364 ( \14741 , \2353 , \4376 );
nand \U$14365 ( \14742 , \14740 , \14741 );
nand \U$14366 ( \14743 , \14742 , \5135 );
nand \U$14367 ( \14744 , \14737 , \14743 );
not \U$14368 ( \14745 , \1963 );
not \U$14369 ( \14746 , RIc226e30_17);
not \U$14370 ( \14747 , \11672 );
or \U$14371 ( \14748 , \14746 , \14747 );
nand \U$14372 ( \14749 , \2981 , \1935 );
nand \U$14373 ( \14750 , \14748 , \14749 );
not \U$14374 ( \14751 , \14750 );
or \U$14375 ( \14752 , \14745 , \14751 );
nand \U$14376 ( \14753 , \14303 , \1945 );
nand \U$14377 ( \14754 , \14752 , \14753 );
xor \U$14378 ( \14755 , \14744 , \14754 );
not \U$14379 ( \14756 , \2534 );
not \U$14380 ( \14757 , RIc226d40_19);
not \U$14381 ( \14758 , \2104 );
or \U$14382 ( \14759 , \14757 , \14758 );
nand \U$14383 ( \14760 , \9654 , \1941 );
nand \U$14384 ( \14761 , \14759 , \14760 );
not \U$14385 ( \14762 , \14761 );
or \U$14386 ( \14763 , \14756 , \14762 );
nand \U$14387 ( \14764 , \14470 , \2518 );
nand \U$14388 ( \14765 , \14763 , \14764 );
xor \U$14389 ( \14766 , \14755 , \14765 );
xnor \U$14390 ( \14767 , \14734 , \14766 );
not \U$14391 ( \14768 , \14767 );
not \U$14392 ( \14769 , \14768 );
or \U$14393 ( \14770 , \14701 , \14769 );
nand \U$14394 ( \14771 , \14767 , \14699 );
nand \U$14395 ( \14772 , \14770 , \14771 );
not \U$14396 ( \14773 , \14136 );
not \U$14397 ( \14774 , \14141 );
or \U$14398 ( \14775 , \14773 , \14774 );
or \U$14399 ( \14776 , \14141 , \14136 );
nand \U$14400 ( \14777 , \14776 , \14130 );
nand \U$14401 ( \14778 , \14775 , \14777 );
xnor \U$14402 ( \14779 , \14772 , \14778 );
and \U$14403 ( \14780 , \14607 , \14779 );
not \U$14404 ( \14781 , \14607 );
xor \U$14405 ( \14782 , \14772 , \14778 );
and \U$14406 ( \14783 , \14781 , \14782 );
nor \U$14407 ( \14784 , \14780 , \14783 );
not \U$14408 ( \14785 , \14102 );
not \U$14409 ( \14786 , \14152 );
or \U$14410 ( \14787 , \14785 , \14786 );
or \U$14411 ( \14788 , \14152 , \14102 );
not \U$14412 ( \14789 , \14142 );
nand \U$14413 ( \14790 , \14788 , \14789 );
nand \U$14414 ( \14791 , \14787 , \14790 );
xor \U$14415 ( \14792 , \14784 , \14791 );
not \U$14416 ( \14793 , \14792 );
or \U$14417 ( \14794 , \14600 , \14793 );
buf \U$14418 ( \14795 , \14599 );
or \U$14419 ( \14796 , \14795 , \14792 );
nand \U$14420 ( \14797 , \14794 , \14796 );
not \U$14421 ( \14798 , \14797 );
or \U$14422 ( \14799 , \14591 , \14798 );
or \U$14423 ( \14800 , \14590 , \14797 );
nand \U$14424 ( \14801 , \14799 , \14800 );
not \U$14425 ( \14802 , \14165 );
not \U$14426 ( \14803 , \14170 );
or \U$14427 ( \14804 , \14802 , \14803 );
not \U$14428 ( \14805 , \14169 );
not \U$14429 ( \14806 , \14165 );
not \U$14430 ( \14807 , \14806 );
or \U$14431 ( \14808 , \14805 , \14807 );
nand \U$14432 ( \14809 , \14808 , \14176 );
nand \U$14433 ( \14810 , \14804 , \14809 );
not \U$14434 ( \14811 , \14542 );
buf \U$14435 ( \14812 , \14518 );
nand \U$14436 ( \14813 , \14811 , \14812 );
and \U$14437 ( \14814 , \14813 , \14522 );
nor \U$14438 ( \14815 , \14811 , \14812 );
nor \U$14439 ( \14816 , \14814 , \14815 );
not \U$14440 ( \14817 , \14816 );
and \U$14441 ( \14818 , \14810 , \14817 );
not \U$14442 ( \14819 , \14810 );
and \U$14443 ( \14820 , \14819 , \14816 );
nor \U$14444 ( \14821 , \14818 , \14820 );
not \U$14445 ( \14822 , \14371 );
not \U$14446 ( \14823 , \14348 );
or \U$14447 ( \14824 , \14822 , \14823 );
or \U$14448 ( \14825 , \14348 , \14371 );
nand \U$14449 ( \14826 , \14825 , \14296 );
nand \U$14450 ( \14827 , \14824 , \14826 );
xor \U$14451 ( \14828 , \14821 , \14827 );
xor \U$14452 ( \14829 , \14462 , \14472 );
and \U$14453 ( \14830 , \14829 , \14484 );
and \U$14454 ( \14831 , \14462 , \14472 );
or \U$14455 ( \14832 , \14830 , \14831 );
not \U$14456 ( \14833 , \14832 );
not \U$14457 ( \14834 , \14223 );
not \U$14458 ( \14835 , \14208 );
or \U$14459 ( \14836 , \14834 , \14835 );
nand \U$14460 ( \14837 , \14836 , \14198 );
nand \U$14461 ( \14838 , \14207 , \14222 );
nand \U$14462 ( \14839 , \14837 , \14838 );
not \U$14463 ( \14840 , \14839 );
not \U$14464 ( \14841 , \14840 );
not \U$14465 ( \14842 , \14317 );
not \U$14466 ( \14843 , \14332 );
or \U$14467 ( \14844 , \14842 , \14843 );
not \U$14468 ( \14845 , \14331 );
not \U$14469 ( \14846 , \14318 );
or \U$14470 ( \14847 , \14845 , \14846 );
nand \U$14471 ( \14848 , \14847 , \14307 );
nand \U$14472 ( \14849 , \14844 , \14848 );
not \U$14473 ( \14850 , \14849 );
or \U$14474 ( \14851 , \14841 , \14850 );
or \U$14475 ( \14852 , \14840 , \14849 );
nand \U$14476 ( \14853 , \14851 , \14852 );
not \U$14477 ( \14854 , \14853 );
not \U$14478 ( \14855 , \14854 );
or \U$14479 ( \14856 , \14833 , \14855 );
not \U$14480 ( \14857 , \14832 );
nand \U$14481 ( \14858 , \14857 , \14853 );
nand \U$14482 ( \14859 , \14856 , \14858 );
not \U$14483 ( \14860 , \14337 );
not \U$14484 ( \14861 , \14342 );
or \U$14485 ( \14862 , \14860 , \14861 );
not \U$14486 ( \14863 , \14337 );
not \U$14487 ( \14864 , \14863 );
not \U$14488 ( \14865 , \14341 );
or \U$14489 ( \14866 , \14864 , \14865 );
nand \U$14490 ( \14867 , \14866 , \14347 );
nand \U$14491 ( \14868 , \14862 , \14867 );
xor \U$14492 ( \14869 , \14859 , \14868 );
or \U$14493 ( \14870 , \14370 , \14365 );
nand \U$14494 ( \14871 , \14870 , \14357 );
nand \U$14495 ( \14872 , \14365 , \14370 );
nand \U$14496 ( \14873 , \14871 , \14872 );
not \U$14497 ( \14874 , \14873 );
and \U$14498 ( \14875 , \14869 , \14874 );
not \U$14499 ( \14876 , \14869 );
and \U$14500 ( \14877 , \14876 , \14873 );
nor \U$14501 ( \14878 , \14875 , \14877 );
or \U$14502 ( \14879 , \14534 , \14527 );
and \U$14503 ( \14880 , \14879 , \14541 );
and \U$14504 ( \14881 , \14527 , \14534 );
nor \U$14505 ( \14882 , \14880 , \14881 );
not \U$14506 ( \14883 , \14261 );
not \U$14507 ( \14884 , \14264 );
or \U$14508 ( \14885 , \14883 , \14884 );
not \U$14509 ( \14886 , \14227 );
not \U$14510 ( \14887 , \14260 );
or \U$14511 ( \14888 , \14886 , \14887 );
nand \U$14512 ( \14889 , \14888 , \14295 );
nand \U$14513 ( \14890 , \14885 , \14889 );
not \U$14514 ( \14891 , \14890 );
xor \U$14515 ( \14892 , \14882 , \14891 );
not \U$14516 ( \14893 , \14247 );
not \U$14517 ( \14894 , \14238 );
or \U$14518 ( \14895 , \14893 , \14894 );
not \U$14519 ( \14896 , \14238 );
nand \U$14520 ( \14897 , \14896 , \14248 );
nand \U$14521 ( \14898 , \14897 , \14259 );
nand \U$14522 ( \14899 , \14895 , \14898 );
not \U$14523 ( \14900 , \1118 );
not \U$14524 ( \14901 , \14203 );
or \U$14525 ( \14902 , \14900 , \14901 );
not \U$14526 ( \14903 , RIc2272e0_7);
not \U$14527 ( \14904 , \9884 );
or \U$14528 ( \14905 , \14903 , \14904 );
nand \U$14529 ( \14906 , \8885 , \1139 );
nand \U$14530 ( \14907 , \14905 , \14906 );
nand \U$14531 ( \14908 , \14907 , \1121 );
nand \U$14532 ( \14909 , \14902 , \14908 );
not \U$14533 ( \14910 , \8830 );
xor \U$14534 ( \14911 , \956 , \14910 );
not \U$14535 ( \14912 , \14911 );
not \U$14536 ( \14913 , \955 );
and \U$14537 ( \14914 , \14912 , \14913 );
and \U$14538 ( \14915 , \14245 , \951 );
nor \U$14539 ( \14916 , \14914 , \14915 );
xor \U$14540 ( \14917 , \14909 , \14916 );
not \U$14541 ( \14918 , \1340 );
not \U$14542 ( \14919 , RIc2271f0_9);
not \U$14543 ( \14920 , \9859 );
or \U$14544 ( \14921 , \14919 , \14920 );
nand \U$14545 ( \14922 , \9740 , \1351 );
nand \U$14546 ( \14923 , \14921 , \14922 );
not \U$14547 ( \14924 , \14923 );
or \U$14548 ( \14925 , \14918 , \14924 );
nand \U$14549 ( \14926 , \14220 , \1363 );
nand \U$14550 ( \14927 , \14925 , \14926 );
xor \U$14551 ( \14928 , \14917 , \14927 );
xor \U$14552 ( \14929 , \14899 , \14928 );
not \U$14553 ( \14930 , \2172 );
not \U$14554 ( \14931 , RIc226a70_25);
not \U$14555 ( \14932 , \13780 );
or \U$14556 ( \14933 , \14931 , \14932 );
nand \U$14557 ( \14934 , \2475 , \9662 );
nand \U$14558 ( \14935 , \14933 , \14934 );
not \U$14559 ( \14936 , \14935 );
or \U$14560 ( \14937 , \14930 , \14936 );
nand \U$14561 ( \14938 , \14510 , \2195 );
nand \U$14562 ( \14939 , \14937 , \14938 );
not \U$14563 ( \14940 , \6307 );
not \U$14564 ( \14941 , RIc2263e0_39);
not \U$14565 ( \14942 , \1530 );
or \U$14566 ( \14943 , \14941 , \14942 );
nand \U$14567 ( \14944 , \1529 , \9573 );
nand \U$14568 ( \14945 , \14943 , \14944 );
not \U$14569 ( \14946 , \14945 );
or \U$14570 ( \14947 , \14940 , \14946 );
nand \U$14571 ( \14948 , \14502 , \6688 );
nand \U$14572 ( \14949 , \14947 , \14948 );
xor \U$14573 ( \14950 , \14939 , \14949 );
not \U$14574 ( \14951 , \5509 );
not \U$14575 ( \14952 , \14257 );
or \U$14576 ( \14953 , \14951 , \14952 );
not \U$14577 ( \14954 , RIc2264d0_37);
not \U$14578 ( \14955 , \3783 );
or \U$14579 ( \14956 , \14954 , \14955 );
nand \U$14580 ( \14957 , \3043 , \5504 );
nand \U$14581 ( \14958 , \14956 , \14957 );
nand \U$14582 ( \14959 , \14958 , \5519 );
nand \U$14583 ( \14960 , \14953 , \14959 );
xor \U$14584 ( \14961 , \14950 , \14960 );
xor \U$14585 ( \14962 , \14929 , \14961 );
xor \U$14586 ( \14963 , \14892 , \14962 );
xor \U$14587 ( \14964 , \14878 , \14963 );
not \U$14588 ( \14965 , \1579 );
and \U$14589 ( \14966 , RIc2275b0_1, \8910 );
not \U$14590 ( \14967 , RIc2275b0_1);
not \U$14591 ( \14968 , \8910 );
and \U$14592 ( \14969 , \14967 , \14968 );
or \U$14593 ( \14970 , \14966 , \14969 );
not \U$14594 ( \14971 , \14970 );
or \U$14595 ( \14972 , \14965 , \14971 );
nand \U$14596 ( \14973 , \14118 , \854 );
nand \U$14597 ( \14974 , \14972 , \14973 );
not \U$14598 ( \14975 , \9534 );
not \U$14599 ( \14976 , \14460 );
or \U$14600 ( \14977 , \14975 , \14976 );
nand \U$14601 ( \14978 , \9552 , RIc225f30_49);
nand \U$14602 ( \14979 , \14977 , \14978 );
xor \U$14603 ( \14980 , \14974 , \14979 );
not \U$14604 ( \14981 , \1082 );
not \U$14605 ( \14982 , RIc2274c0_3);
not \U$14606 ( \14983 , \11566 );
or \U$14607 ( \14984 , \14982 , \14983 );
nand \U$14608 ( \14985 , \9916 , \1032 );
nand \U$14609 ( \14986 , \14984 , \14985 );
not \U$14610 ( \14987 , \14986 );
or \U$14611 ( \14988 , \14981 , \14987 );
nand \U$14612 ( \14989 , \14236 , \1040 );
nand \U$14613 ( \14990 , \14988 , \14989 );
xor \U$14614 ( \14991 , \14980 , \14990 );
not \U$14615 ( \14992 , \1307 );
not \U$14616 ( \14993 , \14196 );
or \U$14617 ( \14994 , \14992 , \14993 );
not \U$14618 ( \14995 , RIc227100_11);
not \U$14619 ( \14996 , \13687 );
or \U$14620 ( \14997 , \14995 , \14996 );
not \U$14621 ( \14998 , \9768 );
nand \U$14622 ( \14999 , \14998 , \1291 );
nand \U$14623 ( \15000 , \14997 , \14999 );
nand \U$14624 ( \15001 , \15000 , \1311 );
nand \U$14625 ( \15002 , \14994 , \15001 );
not \U$14626 ( \15003 , \1682 );
not \U$14627 ( \15004 , RIc227010_13);
not \U$14628 ( \15005 , \13512 );
or \U$14629 ( \15006 , \15004 , \15005 );
not \U$14630 ( \15007 , \13512 );
nand \U$14631 ( \15008 , \15007 , \3841 );
nand \U$14632 ( \15009 , \15006 , \15008 );
not \U$14633 ( \15010 , \15009 );
or \U$14634 ( \15011 , \15003 , \15010 );
nand \U$14635 ( \15012 , \14329 , \1678 );
nand \U$14636 ( \15013 , \15011 , \15012 );
xor \U$14637 ( \15014 , \15002 , \15013 );
not \U$14638 ( \15015 , \2358 );
not \U$14639 ( \15016 , RIc226f20_15);
not \U$14640 ( \15017 , \4122 );
or \U$14641 ( \15018 , \15016 , \15017 );
nand \U$14642 ( \15019 , \10209 , \2301 );
nand \U$14643 ( \15020 , \15018 , \15019 );
not \U$14644 ( \15021 , \15020 );
or \U$14645 ( \15022 , \15015 , \15021 );
nand \U$14646 ( \15023 , \14313 , \2320 );
nand \U$14647 ( \15024 , \15022 , \15023 );
xor \U$14648 ( \15025 , \15014 , \15024 );
xor \U$14649 ( \15026 , \14991 , \15025 );
not \U$14650 ( \15027 , \14517 );
not \U$14651 ( \15028 , \13779 );
or \U$14652 ( \15029 , \15027 , \15028 );
not \U$14653 ( \15030 , \13779 );
not \U$14654 ( \15031 , \15030 );
not \U$14655 ( \15032 , \14516 );
or \U$14656 ( \15033 , \15031 , \15032 );
nand \U$14657 ( \15034 , \15033 , \14504 );
nand \U$14658 ( \15035 , \15029 , \15034 );
xor \U$14659 ( \15036 , \15026 , \15035 );
not \U$14660 ( \15037 , \14485 );
not \U$14661 ( \15038 , \14451 );
or \U$14662 ( \15039 , \15037 , \15038 );
or \U$14663 ( \15040 , \14485 , \14451 );
buf \U$14664 ( \15041 , \14418 );
nand \U$14665 ( \15042 , \15040 , \15041 );
nand \U$14666 ( \15043 , \15039 , \15042 );
xor \U$14667 ( \15044 , \15036 , \15043 );
xor \U$14668 ( \15045 , \14429 , \14439 );
and \U$14669 ( \15046 , \15045 , \14450 );
and \U$14670 ( \15047 , \14429 , \14439 );
or \U$14671 ( \15048 , \15046 , \15047 );
xor \U$14672 ( \15049 , \14396 , \14406 );
and \U$14673 ( \15050 , \15049 , \14417 );
and \U$14674 ( \15051 , \14396 , \14406 );
or \U$14675 ( \15052 , \15050 , \15051 );
xor \U$14676 ( \15053 , \15048 , \15052 );
buf \U$14677 ( \15054 , \14284 );
not \U$14678 ( \15055 , \15054 );
not \U$14679 ( \15056 , \14272 );
or \U$14680 ( \15057 , \15055 , \15056 );
or \U$14681 ( \15058 , \15054 , \14272 );
nand \U$14682 ( \15059 , \15058 , \14294 );
nand \U$14683 ( \15060 , \15057 , \15059 );
xor \U$14684 ( \15061 , \15053 , \15060 );
not \U$14685 ( \15062 , \15061 );
xnor \U$14686 ( \15063 , \15044 , \15062 );
not \U$14687 ( \15064 , \15063 );
and \U$14688 ( \15065 , \14964 , \15064 );
not \U$14689 ( \15066 , \14964 );
and \U$14690 ( \15067 , \15066 , \15063 );
nor \U$14691 ( \15068 , \15065 , \15067 );
not \U$14692 ( \15069 , \15068 );
xor \U$14693 ( \15070 , \14828 , \15069 );
xor \U$14694 ( \15071 , \14177 , \14186 );
and \U$14695 ( \15072 , \15071 , \14372 );
and \U$14696 ( \15073 , \14177 , \14186 );
or \U$14697 ( \15074 , \15072 , \15073 );
xor \U$14698 ( \15075 , \15070 , \15074 );
and \U$14699 ( \15076 , \14801 , \15075 );
not \U$14700 ( \15077 , \14801 );
not \U$14701 ( \15078 , \15075 );
and \U$14702 ( \15079 , \15077 , \15078 );
nor \U$14703 ( \15080 , \15076 , \15079 );
not \U$14704 ( \15081 , \14556 );
nand \U$14705 ( \15082 , \15081 , \14380 );
not \U$14706 ( \15083 , \15082 );
not \U$14707 ( \15084 , \14567 );
or \U$14708 ( \15085 , \15083 , \15084 );
nand \U$14709 ( \15086 , \14379 , \14556 );
nand \U$14710 ( \15087 , \15085 , \15086 );
buf \U$14711 ( \15088 , \15087 );
xnor \U$14712 ( \15089 , \15080 , \15088 );
nand \U$14713 ( \15090 , \14583 , \15089 );
xor \U$14714 ( \15091 , \13731 , \13740 );
and \U$14715 ( \15092 , \15091 , \14084 );
and \U$14716 ( \15093 , \13731 , \13740 );
or \U$14717 ( \15094 , \15092 , \15093 );
not \U$14718 ( \15095 , \15094 );
xor \U$14719 ( \15096 , \14374 , \14572 );
xor \U$14720 ( \15097 , \15096 , \14580 );
nand \U$14721 ( \15098 , \15095 , \15097 );
nand \U$14722 ( \15099 , \15090 , \15098 );
nor \U$14723 ( \15100 , \14093 , \15099 );
not \U$14724 ( \15101 , \15100 );
xor \U$14725 ( \15102 , \12635 , \12903 );
xor \U$14726 ( \15103 , \15102 , \12914 );
xor \U$14727 ( \15104 , \12660 , \12741 );
xor \U$14728 ( \15105 , \15104 , \12895 );
not \U$14729 ( \15106 , \15105 );
not \U$14730 ( \15107 , \12931 );
not \U$14731 ( \15108 , \13059 );
not \U$14732 ( \15109 , \15108 );
or \U$14733 ( \15110 , \15107 , \15109 );
nand \U$14734 ( \15111 , \12930 , \13059 );
nand \U$14735 ( \15112 , \15110 , \15111 );
and \U$14736 ( \15113 , \15112 , \13140 );
not \U$14737 ( \15114 , \15112 );
not \U$14738 ( \15115 , \13140 );
and \U$14739 ( \15116 , \15114 , \15115 );
nor \U$14740 ( \15117 , \15113 , \15116 );
not \U$14741 ( \15118 , \15117 );
or \U$14742 ( \15119 , \15106 , \15118 );
or \U$14743 ( \15120 , \15105 , \15117 );
not \U$14744 ( \15121 , \9488 );
not \U$14745 ( \15122 , RIc225d50_53);
not \U$14746 ( \15123 , \10427 );
or \U$14747 ( \15124 , \15122 , \15123 );
nand \U$14748 ( \15125 , \1439 , \11585 );
nand \U$14749 ( \15126 , \15124 , \15125 );
not \U$14750 ( \15127 , \15126 );
or \U$14751 ( \15128 , \15121 , \15127 );
nand \U$14752 ( \15129 , \12953 , \8788 );
nand \U$14753 ( \15130 , \15128 , \15129 );
not \U$14754 ( \15131 , \15130 );
not \U$14755 ( \15132 , RIc226200_43);
not \U$14756 ( \15133 , \2226 );
or \U$14757 ( \15134 , \15132 , \15133 );
nand \U$14758 ( \15135 , \2225 , \9117 );
nand \U$14759 ( \15136 , \15134 , \15135 );
buf \U$14760 ( \15137 , \15136 );
and \U$14761 ( \15138 , \15137 , \9110 );
and \U$14762 ( \15139 , \13069 , \9205 );
nor \U$14763 ( \15140 , \15138 , \15139 );
nand \U$14764 ( \15141 , \15131 , \15140 );
not \U$14765 ( \15142 , \11697 );
not \U$14766 ( \15143 , RIc225c60_55);
not \U$14767 ( \15144 , \2118 );
or \U$14768 ( \15145 , \15143 , \15144 );
nand \U$14769 ( \15146 , \1020 , \11108 );
nand \U$14770 ( \15147 , \15145 , \15146 );
not \U$14771 ( \15148 , \15147 );
or \U$14772 ( \15149 , \15142 , \15148 );
nand \U$14773 ( \15150 , \13021 , \11038 );
nand \U$14774 ( \15151 , \15149 , \15150 );
and \U$14775 ( \15152 , \15141 , \15151 );
not \U$14776 ( \15153 , \15130 );
nor \U$14777 ( \15154 , \15153 , \15140 );
nor \U$14778 ( \15155 , \15152 , \15154 );
not \U$14779 ( \15156 , \15155 );
not \U$14780 ( \15157 , \15156 );
not \U$14781 ( \15158 , \9142 );
not \U$14782 ( \15159 , \13106 );
or \U$14783 ( \15160 , \15158 , \15159 );
xor \U$14784 ( \15161 , RIc226890_29, \2980 );
nand \U$14785 ( \15162 , \15161 , \2784 );
nand \U$14786 ( \15163 , \15160 , \15162 );
buf \U$14787 ( \15164 , \12665 );
not \U$14788 ( \15165 , \15164 );
and \U$14789 ( \15166 , RIc225a80_59, \9491 );
not \U$14790 ( \15167 , RIc225a80_59);
and \U$14791 ( \15168 , \15167 , \1072 );
or \U$14792 ( \15169 , \15166 , \15168 );
not \U$14793 ( \15170 , \15169 );
or \U$14794 ( \15171 , \15165 , \15170 );
nand \U$14795 ( \15172 , \12667 , \12670 );
nand \U$14796 ( \15173 , \15171 , \15172 );
or \U$14797 ( \15174 , \15163 , \15173 );
not \U$14798 ( \15175 , \9934 );
not \U$14799 ( \15176 , RIc226110_45);
not \U$14800 ( \15177 , \3686 );
or \U$14801 ( \15178 , \15176 , \15177 );
nand \U$14802 ( \15179 , \2422 , \14390 );
nand \U$14803 ( \15180 , \15178 , \15179 );
not \U$14804 ( \15181 , \15180 );
or \U$14805 ( \15182 , \15175 , \15181 );
buf \U$14806 ( \15183 , \9398 );
nand \U$14807 ( \15184 , \13117 , \15183 );
nand \U$14808 ( \15185 , \15182 , \15184 );
nand \U$14809 ( \15186 , \15174 , \15185 );
nand \U$14810 ( \15187 , \15173 , \15163 );
nand \U$14811 ( \15188 , \15186 , \15187 );
not \U$14812 ( \15189 , \15188 );
or \U$14813 ( \15190 , \15157 , \15189 );
not \U$14814 ( \15191 , \15188 );
nand \U$14815 ( \15192 , \15191 , \15155 );
not \U$14816 ( \15193 , \1682 );
not \U$14817 ( \15194 , \12687 );
or \U$14818 ( \15195 , \15193 , \15194 );
and \U$14819 ( \15196 , RIc227010_13, \12403 );
not \U$14820 ( \15197 , RIc227010_13);
and \U$14821 ( \15198 , \15197 , \9786 );
or \U$14822 ( \15199 , \15196 , \15198 );
nand \U$14823 ( \15200 , \15199 , \3250 );
nand \U$14824 ( \15201 , \15195 , \15200 );
not \U$14825 ( \15202 , \9619 );
not \U$14826 ( \15203 , \13239 );
or \U$14827 ( \15204 , \15202 , \15203 );
and \U$14828 ( \15205 , \2345 , RIc226020_47);
not \U$14829 ( \15206 , \2345 );
and \U$14830 ( \15207 , \15206 , \11607 );
or \U$14831 ( \15208 , \15205 , \15207 );
nand \U$14832 ( \15209 , \15208 , \10001 );
nand \U$14833 ( \15210 , \15204 , \15209 );
xor \U$14834 ( \15211 , \15201 , \15210 );
not \U$14835 ( \15212 , \2697 );
not \U$14836 ( \15213 , RIc2267a0_31);
not \U$14837 ( \15214 , \9651 );
or \U$14838 ( \15215 , \15213 , \15214 );
not \U$14839 ( \15216 , \2103 );
not \U$14840 ( \15217 , \15216 );
nand \U$14841 ( \15218 , \15217 , \3648 );
nand \U$14842 ( \15219 , \15215 , \15218 );
not \U$14843 ( \15220 , \15219 );
or \U$14844 ( \15221 , \15212 , \15220 );
nand \U$14845 ( \15222 , \13253 , \2711 );
nand \U$14846 ( \15223 , \15221 , \15222 );
and \U$14847 ( \15224 , \15211 , \15223 );
and \U$14848 ( \15225 , \15201 , \15210 );
or \U$14849 ( \15226 , \15224 , \15225 );
nand \U$14850 ( \15227 , \15192 , \15226 );
nand \U$14851 ( \15228 , \15190 , \15227 );
and \U$14852 ( \15229 , \12702 , \2392 );
and \U$14853 ( \15230 , \12704 , \2367 );
nor \U$14854 ( \15231 , \15229 , \15230 );
not \U$14855 ( \15232 , \15231 );
not \U$14856 ( \15233 , \12718 );
or \U$14857 ( \15234 , \15232 , \15233 );
or \U$14858 ( \15235 , \12706 , \12718 );
nand \U$14859 ( \15236 , \15234 , \15235 );
not \U$14860 ( \15237 , \15236 );
not \U$14861 ( \15238 , \12733 );
not \U$14862 ( \15239 , \15238 );
and \U$14863 ( \15240 , \15237 , \15239 );
and \U$14864 ( \15241 , \15236 , \15238 );
nor \U$14865 ( \15242 , \15240 , \15241 );
not \U$14866 ( \15243 , \15242 );
not \U$14867 ( \15244 , \15243 );
not \U$14868 ( \15245 , \12672 );
not \U$14869 ( \15246 , \12691 );
not \U$14870 ( \15247 , \15246 );
or \U$14871 ( \15248 , \15245 , \15247 );
nand \U$14872 ( \15249 , \12673 , \12691 );
nand \U$14873 ( \15250 , \15248 , \15249 );
not \U$14874 ( \15251 , \12681 );
and \U$14875 ( \15252 , \15250 , \15251 );
not \U$14876 ( \15253 , \15250 );
and \U$14877 ( \15254 , \15253 , \12681 );
nor \U$14878 ( \15255 , \15252 , \15254 );
not \U$14879 ( \15256 , \15255 );
or \U$14880 ( \15257 , \15244 , \15256 );
not \U$14881 ( \15258 , \11965 );
not \U$14882 ( \15259 , RIc225b70_57);
not \U$14883 ( \15260 , \1706 );
or \U$14884 ( \15261 , \15259 , \15260 );
not \U$14885 ( \15262 , RIc225b70_57);
nand \U$14886 ( \15263 , \840 , \15262 );
nand \U$14887 ( \15264 , \15261 , \15263 );
not \U$14888 ( \15265 , \15264 );
or \U$14889 ( \15266 , \15258 , \15265 );
buf \U$14890 ( \15267 , \11974 );
nand \U$14891 ( \15268 , \15267 , \13081 );
nand \U$14892 ( \15269 , \15266 , \15268 );
not \U$14893 ( \15270 , \15269 );
not \U$14894 ( \15271 , \6688 );
and \U$14895 ( \15272 , \9422 , RIc2263e0_39);
not \U$14896 ( \15273 , \9422 );
and \U$14897 ( \15274 , \15273 , \8998 );
or \U$14898 ( \15275 , \15272 , \15274 );
not \U$14899 ( \15276 , \15275 );
or \U$14900 ( \15277 , \15271 , \15276 );
nand \U$14901 ( \15278 , \13037 , \6307 );
nand \U$14902 ( \15279 , \15277 , \15278 );
not \U$14903 ( \15280 , \15279 );
or \U$14904 ( \15281 , \15270 , \15280 );
or \U$14905 ( \15282 , \15269 , \15279 );
not \U$14906 ( \15283 , \9690 );
not \U$14907 ( \15284 , RIc2262f0_41);
not \U$14908 ( \15285 , \5767 );
or \U$14909 ( \15286 , \15284 , \15285 );
not \U$14910 ( \15287 , \9408 );
nand \U$14911 ( \15288 , \15287 , \9822 );
nand \U$14912 ( \15289 , \15286 , \15288 );
not \U$14913 ( \15290 , \15289 );
or \U$14914 ( \15291 , \15283 , \15290 );
nand \U$14915 ( \15292 , \12939 , \9705 );
nand \U$14916 ( \15293 , \15291 , \15292 );
nand \U$14917 ( \15294 , \15282 , \15293 );
nand \U$14918 ( \15295 , \15281 , \15294 );
not \U$14919 ( \15296 , \15255 );
nand \U$14920 ( \15297 , \15296 , \15242 );
nand \U$14921 ( \15298 , \15295 , \15297 );
nand \U$14922 ( \15299 , \15257 , \15298 );
or \U$14923 ( \15300 , \15228 , \15299 );
xor \U$14924 ( \15301 , \12662 , \12739 );
xnor \U$14925 ( \15302 , \15301 , \12736 );
not \U$14926 ( \15303 , \15302 );
nand \U$14927 ( \15304 , \15300 , \15303 );
nand \U$14928 ( \15305 , \15299 , \15228 );
nand \U$14929 ( \15306 , \15304 , \15305 );
nand \U$14930 ( \15307 , \15120 , \15306 );
nand \U$14931 ( \15308 , \15119 , \15307 );
not \U$14932 ( \15309 , \15308 );
xor \U$14933 ( \15310 , \12927 , \13142 );
xnor \U$14934 ( \15311 , \15310 , \13179 );
nand \U$14935 ( \15312 , \15309 , \15311 );
not \U$14936 ( \15313 , \15312 );
xor \U$14937 ( \15314 , \13186 , \13188 );
xor \U$14938 ( \15315 , \15314 , \13292 );
not \U$14939 ( \15316 , \15315 );
or \U$14940 ( \15317 , \15313 , \15316 );
not \U$14941 ( \15318 , \15311 );
nand \U$14942 ( \15319 , \15318 , \15308 );
nand \U$14943 ( \15320 , \15317 , \15319 );
xor \U$14944 ( \15321 , \13181 , \13183 );
xor \U$14945 ( \15322 , \15321 , \13295 );
xor \U$14946 ( \15323 , \15320 , \15322 );
not \U$14947 ( \15324 , \13166 );
not \U$14948 ( \15325 , \13175 );
or \U$14949 ( \15326 , \15324 , \15325 );
nand \U$14950 ( \15327 , \13163 , \13165 );
nand \U$14951 ( \15328 , \15326 , \15327 );
not \U$14952 ( \15329 , \13170 );
and \U$14953 ( \15330 , \15328 , \15329 );
not \U$14954 ( \15331 , \15328 );
and \U$14955 ( \15332 , \15331 , \13170 );
nor \U$14956 ( \15333 , \15330 , \15332 );
not \U$14957 ( \15334 , \15333 );
not \U$14958 ( \15335 , \15334 );
not \U$14959 ( \15336 , \13008 );
not \U$14960 ( \15337 , \12997 );
or \U$14961 ( \15338 , \15336 , \15337 );
or \U$14962 ( \15339 , \13008 , \12997 );
nand \U$14963 ( \15340 , \15338 , \15339 );
and \U$14964 ( \15341 , \15340 , \12984 );
not \U$14965 ( \15342 , \15340 );
and \U$14966 ( \15343 , \15342 , \12983 );
nor \U$14967 ( \15344 , \15341 , \15343 );
xor \U$14968 ( \15345 , \13134 , \13121 );
xnor \U$14969 ( \15346 , \15345 , \13110 );
nand \U$14970 ( \15347 , \15344 , \15346 );
not \U$14971 ( \15348 , \13096 );
not \U$14972 ( \15349 , \13085 );
and \U$14973 ( \15350 , \15348 , \15349 );
and \U$14974 ( \15351 , \13096 , \13085 );
nor \U$14975 ( \15352 , \15350 , \15351 );
not \U$14976 ( \15353 , \13073 );
and \U$14977 ( \15354 , \15352 , \15353 );
not \U$14978 ( \15355 , \15352 );
and \U$14979 ( \15356 , \15355 , \13073 );
nor \U$14980 ( \15357 , \15354 , \15356 );
and \U$14981 ( \15358 , \15347 , \15357 );
nor \U$14982 ( \15359 , \15346 , \15344 );
nor \U$14983 ( \15360 , \15358 , \15359 );
not \U$14984 ( \15361 , \15360 );
not \U$14985 ( \15362 , \15361 );
or \U$14986 ( \15363 , \15335 , \15362 );
not \U$14987 ( \15364 , \15360 );
not \U$14988 ( \15365 , \15333 );
or \U$14989 ( \15366 , \15364 , \15365 );
not \U$14990 ( \15367 , \12992 );
not \U$14991 ( \15368 , \15367 );
not \U$14992 ( \15369 , \4383 );
not \U$14993 ( \15370 , \15369 );
and \U$14994 ( \15371 , \15368 , \15370 );
not \U$14995 ( \15372 , RIc2265c0_35);
not \U$14996 ( \15373 , \2670 );
or \U$14997 ( \15374 , \15372 , \15373 );
nand \U$14998 ( \15375 , \9139 , \4376 );
nand \U$14999 ( \15376 , \15374 , \15375 );
and \U$15000 ( \15377 , \15376 , \5741 );
nor \U$15001 ( \15378 , \15371 , \15377 );
not \U$15002 ( \15379 , \15378 );
not \U$15003 ( \15380 , \5509 );
not \U$15004 ( \15381 , RIc2264d0_37);
not \U$15005 ( \15382 , \2475 );
not \U$15006 ( \15383 , \15382 );
or \U$15007 ( \15384 , \15381 , \15383 );
nand \U$15008 ( \15385 , \3036 , \4371 );
nand \U$15009 ( \15386 , \15384 , \15385 );
not \U$15010 ( \15387 , \15386 );
or \U$15011 ( \15388 , \15380 , \15387 );
nand \U$15012 ( \15389 , \13048 , \5519 );
nand \U$15013 ( \15390 , \15388 , \15389 );
not \U$15014 ( \15391 , \15390 );
not \U$15015 ( \15392 , \15391 );
or \U$15016 ( \15393 , \15379 , \15392 );
not \U$15017 ( \15394 , \9459 );
not \U$15018 ( \15395 , RIc225e40_51);
not \U$15019 ( \15396 , \1530 );
or \U$15020 ( \15397 , \15395 , \15396 );
nand \U$15021 ( \15398 , \3579 , \12423 );
nand \U$15022 ( \15399 , \15397 , \15398 );
not \U$15023 ( \15400 , \15399 );
or \U$15024 ( \15401 , \15394 , \15400 );
nand \U$15025 ( \15402 , \9445 , \12965 );
nand \U$15026 ( \15403 , \15401 , \15402 );
nand \U$15027 ( \15404 , \15393 , \15403 );
not \U$15028 ( \15405 , \15378 );
nand \U$15029 ( \15406 , \15405 , \15390 );
nand \U$15030 ( \15407 , \15404 , \15406 );
not \U$15031 ( \15408 , \15407 );
xor \U$15032 ( \15409 , \12852 , \12786 );
xnor \U$15033 ( \15410 , \15409 , \12797 );
nand \U$15034 ( \15411 , \15408 , \15410 );
xor \U$15035 ( \15412 , \13232 , \13243 );
xor \U$15036 ( \15413 , \15412 , \13255 );
and \U$15037 ( \15414 , \15411 , \15413 );
not \U$15038 ( \15415 , \15407 );
nor \U$15039 ( \15416 , \15415 , \15410 );
nor \U$15040 ( \15417 , \15414 , \15416 );
not \U$15041 ( \15418 , \15417 );
nand \U$15042 ( \15419 , \15366 , \15418 );
nand \U$15043 ( \15420 , \15363 , \15419 );
xor \U$15044 ( \15421 , \13064 , \13099 );
xor \U$15045 ( \15422 , \15421 , \13137 );
xor \U$15046 ( \15423 , \12971 , \13013 );
xor \U$15047 ( \15424 , \15423 , \13055 );
xor \U$15048 ( \15425 , \15422 , \15424 );
xor \U$15049 ( \15426 , \12969 , \12943 );
xnor \U$15050 ( \15427 , \15426 , \12955 );
not \U$15051 ( \15428 , \15427 );
not \U$15052 ( \15429 , \13052 );
not \U$15053 ( \15430 , \13040 );
or \U$15054 ( \15431 , \15429 , \15430 );
or \U$15055 ( \15432 , \13052 , \13040 );
nand \U$15056 ( \15433 , \15431 , \15432 );
and \U$15057 ( \15434 , \15433 , \13028 );
not \U$15058 ( \15435 , \15433 );
and \U$15059 ( \15436 , \15435 , \13027 );
nor \U$15060 ( \15437 , \15434 , \15436 );
not \U$15061 ( \15438 , \15437 );
or \U$15062 ( \15439 , \15428 , \15438 );
not \U$15063 ( \15440 , \1579 );
not \U$15064 ( \15441 , \13202 );
or \U$15065 ( \15442 , \15440 , \15441 );
buf \U$15066 ( \15443 , \12824 );
not \U$15067 ( \15444 , \15443 );
and \U$15068 ( \15445 , RIc2275b0_1, \15444 );
not \U$15069 ( \15446 , RIc2275b0_1);
and \U$15070 ( \15447 , \15446 , \15443 );
or \U$15071 ( \15448 , \15445 , \15447 );
nand \U$15072 ( \15449 , \15448 , \854 );
nand \U$15073 ( \15450 , \15442 , \15449 );
not \U$15074 ( \15451 , \954 );
not \U$15075 ( \15452 , \13446 );
or \U$15076 ( \15453 , \15451 , \15452 );
not \U$15077 ( \15454 , RIc2273d0_5);
not \U$15078 ( \15455 , \10360 );
or \U$15079 ( \15456 , \15454 , \15455 );
nand \U$15080 ( \15457 , \10086 , \956 );
nand \U$15081 ( \15458 , \15456 , \15457 );
nand \U$15082 ( \15459 , \15458 , \950 );
nand \U$15083 ( \15460 , \15453 , \15459 );
xor \U$15084 ( \15461 , \15450 , \15460 );
not \U$15085 ( \15462 , \1307 );
not \U$15086 ( \15463 , RIc227100_11);
not \U$15087 ( \15464 , \9076 );
or \U$15088 ( \15465 , \15463 , \15464 );
nand \U$15089 ( \15466 , \10653 , \1302 );
nand \U$15090 ( \15467 , \15465 , \15466 );
not \U$15091 ( \15468 , \15467 );
or \U$15092 ( \15469 , \15462 , \15468 );
nand \U$15093 ( \15470 , \13469 , \1311 );
nand \U$15094 ( \15471 , \15469 , \15470 );
and \U$15095 ( \15472 , \15461 , \15471 );
and \U$15096 ( \15473 , \15450 , \15460 );
or \U$15097 ( \15474 , \15472 , \15473 );
not \U$15098 ( \15475 , \9534 );
not \U$15099 ( \15476 , RIc225f30_49);
not \U$15100 ( \15477 , \3044 );
or \U$15101 ( \15478 , \15476 , \15477 );
nand \U$15102 ( \15479 , \3043 , \9541 );
nand \U$15103 ( \15480 , \15478 , \15479 );
not \U$15104 ( \15481 , \15480 );
or \U$15105 ( \15482 , \15475 , \15481 );
nand \U$15106 ( \15483 , \13004 , \9552 );
nand \U$15107 ( \15484 , \15482 , \15483 );
xor \U$15108 ( \15485 , \15474 , \15484 );
not \U$15109 ( \15486 , \3629 );
not \U$15110 ( \15487 , RIc2266b0_33);
not \U$15111 ( \15488 , \11068 );
or \U$15112 ( \15489 , \15487 , \15488 );
not \U$15113 ( \15490 , \5526 );
nand \U$15114 ( \15491 , \15490 , \5179 );
nand \U$15115 ( \15492 , \15489 , \15491 );
not \U$15116 ( \15493 , \15492 );
or \U$15117 ( \15494 , \15486 , \15493 );
nand \U$15118 ( \15495 , \12981 , \3631 );
nand \U$15119 ( \15496 , \15494 , \15495 );
and \U$15120 ( \15497 , \15485 , \15496 );
and \U$15121 ( \15498 , \15474 , \15484 );
or \U$15122 ( \15499 , \15497 , \15498 );
nand \U$15123 ( \15500 , \15439 , \15499 );
not \U$15124 ( \15501 , \15427 );
not \U$15125 ( \15502 , \15437 );
nand \U$15126 ( \15503 , \15501 , \15502 );
nand \U$15127 ( \15504 , \15500 , \15503 );
and \U$15128 ( \15505 , \15425 , \15504 );
and \U$15129 ( \15506 , \15422 , \15424 );
or \U$15130 ( \15507 , \15505 , \15506 );
xor \U$15131 ( \15508 , \15420 , \15507 );
and \U$15132 ( \15509 , \13177 , \13159 );
not \U$15133 ( \15510 , \13177 );
and \U$15134 ( \15511 , \15510 , \13147 );
or \U$15135 ( \15512 , \15509 , \15511 );
and \U$15136 ( \15513 , \15512 , \13155 );
not \U$15137 ( \15514 , \15512 );
and \U$15138 ( \15515 , \15514 , \13154 );
nor \U$15139 ( \15516 , \15513 , \15515 );
and \U$15140 ( \15517 , \15508 , \15516 );
and \U$15141 ( \15518 , \15420 , \15507 );
or \U$15142 ( \15519 , \15517 , \15518 );
xnor \U$15143 ( \15520 , \13284 , \13276 );
and \U$15144 ( \15521 , \15520 , \13280 );
not \U$15145 ( \15522 , \15520 );
and \U$15146 ( \15523 , \15522 , \13287 );
nor \U$15147 ( \15524 , \15521 , \15523 );
not \U$15148 ( \15525 , \15524 );
not \U$15149 ( \15526 , \13258 );
not \U$15150 ( \15527 , \13194 );
or \U$15151 ( \15528 , \15526 , \15527 );
or \U$15152 ( \15529 , \13194 , \13258 );
nand \U$15153 ( \15530 , \15528 , \15529 );
xnor \U$15154 ( \15531 , \15530 , \13261 );
not \U$15155 ( \15532 , \15531 );
or \U$15156 ( \15533 , \15525 , \15532 );
not \U$15157 ( \15534 , \13396 );
xor \U$15158 ( \15535 , \13393 , \13537 );
not \U$15159 ( \15536 , \15535 );
or \U$15160 ( \15537 , \15534 , \15536 );
or \U$15161 ( \15538 , \15535 , \13396 );
nand \U$15162 ( \15539 , \15537 , \15538 );
nand \U$15163 ( \15540 , \15533 , \15539 );
not \U$15164 ( \15541 , \15524 );
not \U$15165 ( \15542 , \15531 );
nand \U$15166 ( \15543 , \15541 , \15542 );
nand \U$15167 ( \15544 , \15540 , \15543 );
xor \U$15168 ( \15545 , \13263 , \13265 );
xor \U$15169 ( \15546 , \15545 , \13289 );
xor \U$15170 ( \15547 , \15544 , \15546 );
xor \U$15171 ( \15548 , \13539 , \13336 );
xnor \U$15172 ( \15549 , \15548 , \13346 );
and \U$15173 ( \15550 , \15547 , \15549 );
and \U$15174 ( \15551 , \15544 , \15546 );
or \U$15175 ( \15552 , \15550 , \15551 );
xor \U$15176 ( \15553 , \15519 , \15552 );
not \U$15177 ( \15554 , \13324 );
not \U$15178 ( \15555 , \13542 );
or \U$15179 ( \15556 , \15554 , \15555 );
or \U$15180 ( \15557 , \13324 , \13542 );
nand \U$15181 ( \15558 , \15556 , \15557 );
and \U$15182 ( \15559 , \15558 , \13327 );
not \U$15183 ( \15560 , \15558 );
and \U$15184 ( \15561 , \15560 , \13328 );
or \U$15185 ( \15562 , \15559 , \15561 );
and \U$15186 ( \15563 , \15553 , \15562 );
and \U$15187 ( \15564 , \15519 , \15552 );
or \U$15188 ( \15565 , \15563 , \15564 );
and \U$15189 ( \15566 , \15323 , \15565 );
and \U$15190 ( \15567 , \15320 , \15322 );
or \U$15191 ( \15568 , \15566 , \15567 );
xor \U$15192 ( \15569 , \15103 , \15568 );
xor \U$15193 ( \15570 , \13298 , \13300 );
xor \U$15194 ( \15571 , \15570 , \13547 );
xor \U$15195 ( \15572 , \15569 , \15571 );
xor \U$15196 ( \15573 , \13303 , \13545 );
xnor \U$15197 ( \15574 , \15573 , \13317 );
xor \U$15198 ( \15575 , \13206 , \13217 );
xor \U$15199 ( \15576 , \15575 , \13229 );
not \U$15200 ( \15577 , \15576 );
not \U$15201 ( \15578 , \1363 );
not \U$15202 ( \15579 , RIc2271f0_9);
not \U$15203 ( \15580 , \9255 );
or \U$15204 ( \15581 , \15579 , \15580 );
nand \U$15205 ( \15582 , \10986 , \1342 );
nand \U$15206 ( \15583 , \15581 , \15582 );
not \U$15207 ( \15584 , \15583 );
or \U$15208 ( \15585 , \15578 , \15584 );
nand \U$15209 ( \15586 , \13227 , \1339 );
nand \U$15210 ( \15587 , \15585 , \15586 );
not \U$15211 ( \15588 , \1118 );
not \U$15212 ( \15589 , RIc2272e0_7);
not \U$15213 ( \15590 , \9297 );
or \U$15214 ( \15591 , \15589 , \15590 );
nand \U$15215 ( \15592 , \9298 , \1423 );
nand \U$15216 ( \15593 , \15591 , \15592 );
not \U$15217 ( \15594 , \15593 );
or \U$15218 ( \15595 , \15588 , \15594 );
nand \U$15219 ( \15596 , \13457 , \1120 );
nand \U$15220 ( \15597 , \15595 , \15596 );
xor \U$15221 ( \15598 , \15587 , \15597 );
not \U$15222 ( \15599 , \2173 );
not \U$15223 ( \15600 , \13517 );
or \U$15224 ( \15601 , \15599 , \15600 );
not \U$15225 ( \15602 , RIc226a70_25);
not \U$15226 ( \15603 , \5663 );
not \U$15227 ( \15604 , \15603 );
or \U$15228 ( \15605 , \15602 , \15604 );
nand \U$15229 ( \15606 , \5663 , \6107 );
nand \U$15230 ( \15607 , \15605 , \15606 );
nand \U$15231 ( \15608 , \15607 , \2195 );
nand \U$15232 ( \15609 , \15601 , \15608 );
and \U$15233 ( \15610 , \15598 , \15609 );
and \U$15234 ( \15611 , \15587 , \15597 );
or \U$15235 ( \15612 , \15610 , \15611 );
not \U$15236 ( \15613 , \15612 );
or \U$15237 ( \15614 , \15577 , \15613 );
not \U$15238 ( \15615 , \15576 );
not \U$15239 ( \15616 , \15615 );
not \U$15240 ( \15617 , \15612 );
not \U$15241 ( \15618 , \15617 );
or \U$15242 ( \15619 , \15616 , \15618 );
not \U$15243 ( \15620 , RIc2258a0_63);
not \U$15244 ( \15621 , \15620 );
not \U$15245 ( \15622 , RIc2275b0_1);
not \U$15246 ( \15623 , \13488 );
nor \U$15247 ( \15624 , \15622 , \15623 );
not \U$15248 ( \15625 , \15624 );
or \U$15249 ( \15626 , \15621 , \15625 );
nand \U$15250 ( \15627 , \15626 , \13491 );
not \U$15251 ( \15628 , \854 );
not \U$15252 ( \15629 , \12843 );
buf \U$15253 ( \15630 , \15629 );
and \U$15254 ( \15631 , RIc2275b0_1, \15630 );
not \U$15255 ( \15632 , RIc2275b0_1);
not \U$15256 ( \15633 , \15630 );
and \U$15257 ( \15634 , \15632 , \15633 );
or \U$15258 ( \15635 , \15631 , \15634 );
not \U$15259 ( \15636 , \15635 );
or \U$15260 ( \15637 , \15628 , \15636 );
nand \U$15261 ( \15638 , \15448 , \1579 );
nand \U$15262 ( \15639 , \15637 , \15638 );
and \U$15263 ( \15640 , \15627 , \15639 );
not \U$15264 ( \15641 , \10214 );
not \U$15265 ( \15642 , RIc226b60_23);
not \U$15266 ( \15643 , \14192 );
or \U$15267 ( \15644 , \15642 , \15643 );
not \U$15268 ( \15645 , \14192 );
nand \U$15269 ( \15646 , \15645 , \1927 );
nand \U$15270 ( \15647 , \15644 , \15646 );
not \U$15271 ( \15648 , \15647 );
or \U$15272 ( \15649 , \15641 , \15648 );
nand \U$15273 ( \15650 , \13418 , \1930 );
nand \U$15274 ( \15651 , \15649 , \15650 );
xor \U$15275 ( \15652 , \15640 , \15651 );
not \U$15276 ( \15653 , \2138 );
not \U$15277 ( \15654 , RIc226980_27);
not \U$15278 ( \15655 , \9842 );
or \U$15279 ( \15656 , \15654 , \15655 );
nand \U$15280 ( \15657 , \4406 , \2150 );
nand \U$15281 ( \15658 , \15656 , \15657 );
not \U$15282 ( \15659 , \15658 );
or \U$15283 ( \15660 , \15653 , \15659 );
nand \U$15284 ( \15661 , \13530 , \2154 );
nand \U$15285 ( \15662 , \15660 , \15661 );
and \U$15286 ( \15663 , \15652 , \15662 );
and \U$15287 ( \15664 , \15640 , \15651 );
or \U$15288 ( \15665 , \15663 , \15664 );
nand \U$15289 ( \15666 , \15619 , \15665 );
nand \U$15290 ( \15667 , \15614 , \15666 );
xor \U$15291 ( \15668 , \13448 , \13459 );
xor \U$15292 ( \15669 , \15668 , \13471 );
not \U$15293 ( \15670 , \2518 );
not \U$15294 ( \15671 , RIc226d40_19);
not \U$15295 ( \15672 , \10322 );
or \U$15296 ( \15673 , \15671 , \15672 );
nand \U$15297 ( \15674 , \8856 , \1941 );
nand \U$15298 ( \15675 , \15673 , \15674 );
not \U$15299 ( \15676 , \15675 );
or \U$15300 ( \15677 , \15670 , \15676 );
nand \U$15301 ( \15678 , \13430 , \2534 );
nand \U$15302 ( \15679 , \15677 , \15678 );
not \U$15303 ( \15680 , \1945 );
not \U$15304 ( \15681 , RIc226e30_17);
not \U$15305 ( \15682 , \8807 );
or \U$15306 ( \15683 , \15681 , \15682 );
not \U$15307 ( \15684 , \8806 );
not \U$15308 ( \15685 , \15684 );
nand \U$15309 ( \15686 , \15685 , \1935 );
nand \U$15310 ( \15687 , \15683 , \15686 );
not \U$15311 ( \15688 , \15687 );
or \U$15312 ( \15689 , \15680 , \15688 );
nand \U$15313 ( \15690 , \1963 , \13364 );
nand \U$15314 ( \15691 , \15689 , \15690 );
xor \U$15315 ( \15692 , \15679 , \15691 );
not \U$15316 ( \15693 , \2367 );
not \U$15317 ( \15694 , \13407 );
or \U$15318 ( \15695 , \15693 , \15694 );
not \U$15319 ( \15696 , RIc226c50_21);
not \U$15320 ( \15697 , \10142 );
or \U$15321 ( \15698 , \15696 , \15697 );
buf \U$15322 ( \15699 , \9728 );
not \U$15323 ( \15700 , \15699 );
nand \U$15324 ( \15701 , \15700 , \2383 );
nand \U$15325 ( \15702 , \15698 , \15701 );
nand \U$15326 ( \15703 , \15702 , \2392 );
nand \U$15327 ( \15704 , \15695 , \15703 );
and \U$15328 ( \15705 , \15692 , \15704 );
and \U$15329 ( \15706 , \15679 , \15691 );
or \U$15330 ( \15707 , \15705 , \15706 );
xor \U$15331 ( \15708 , \15669 , \15707 );
not \U$15332 ( \15709 , \2358 );
not \U$15333 ( \15710 , \13374 );
or \U$15334 ( \15711 , \15709 , \15710 );
not \U$15335 ( \15712 , RIc226f20_15);
not \U$15336 ( \15713 , \8975 );
or \U$15337 ( \15714 , \15712 , \15713 );
nand \U$15338 ( \15715 , \11994 , \2351 );
nand \U$15339 ( \15716 , \15714 , \15715 );
nand \U$15340 ( \15717 , \15716 , \2320 );
nand \U$15341 ( \15718 , \15711 , \15717 );
buf \U$15342 ( \15719 , \12811 );
not \U$15343 ( \15720 , \15719 );
not \U$15344 ( \15721 , \12806 );
not \U$15345 ( \15722 , \931 );
or \U$15346 ( \15723 , \15721 , \15722 );
not \U$15347 ( \15724 , \930 );
nand \U$15348 ( \15725 , \15724 , RIc225990_61);
nand \U$15349 ( \15726 , \15723 , \15725 );
not \U$15350 ( \15727 , \15726 );
or \U$15351 ( \15728 , \15720 , \15727 );
buf \U$15352 ( \15729 , \12803 );
nand \U$15353 ( \15730 , \15729 , RIc225990_61);
nand \U$15354 ( \15731 , \15728 , \15730 );
nor \U$15355 ( \15732 , \15718 , \15731 );
not \U$15356 ( \15733 , \1682 );
not \U$15357 ( \15734 , \15199 );
or \U$15358 ( \15735 , \15733 , \15734 );
not \U$15359 ( \15736 , RIc227010_13);
not \U$15360 ( \15737 , \13129 );
or \U$15361 ( \15738 , \15736 , \15737 );
nand \U$15362 ( \15739 , \9211 , \1758 );
nand \U$15363 ( \15740 , \15738 , \15739 );
nand \U$15364 ( \15741 , \15740 , \3250 );
nand \U$15365 ( \15742 , \15735 , \15741 );
not \U$15366 ( \15743 , \15742 );
or \U$15367 ( \15744 , \15732 , \15743 );
nand \U$15368 ( \15745 , \15718 , \15731 );
nand \U$15369 ( \15746 , \15744 , \15745 );
and \U$15370 ( \15747 , \15708 , \15746 );
and \U$15371 ( \15748 , \15669 , \15707 );
or \U$15372 ( \15749 , \15747 , \15748 );
xor \U$15373 ( \15750 , \15667 , \15749 );
not \U$15374 ( \15751 , \2710 );
not \U$15375 ( \15752 , \15219 );
or \U$15376 ( \15753 , \15751 , \15752 );
not \U$15377 ( \15754 , RIc2267a0_31);
not \U$15378 ( \15755 , \11324 );
not \U$15379 ( \15756 , \15755 );
or \U$15380 ( \15757 , \15754 , \15756 );
nand \U$15381 ( \15758 , \3115 , \9159 );
nand \U$15382 ( \15759 , \15757 , \15758 );
nand \U$15383 ( \15760 , \15759 , \2697 );
nand \U$15384 ( \15761 , \15753 , \15760 );
not \U$15385 ( \15762 , \15761 );
not \U$15386 ( \15763 , \2086 );
not \U$15387 ( \15764 , \15161 );
or \U$15388 ( \15765 , \15763 , \15764 );
and \U$15389 ( \15766 , RIc226890_29, \14299 );
not \U$15390 ( \15767 , RIc226890_29);
not \U$15391 ( \15768 , \14299 );
and \U$15392 ( \15769 , \15767 , \15768 );
or \U$15393 ( \15770 , \15766 , \15769 );
nand \U$15394 ( \15771 , \15770 , \2784 );
nand \U$15395 ( \15772 , \15765 , \15771 );
not \U$15396 ( \15773 , \15772 );
nand \U$15397 ( \15774 , \15762 , \15773 );
not \U$15398 ( \15775 , \10001 );
not \U$15399 ( \15776 , RIc226020_47);
not \U$15400 ( \15777 , \2304 );
or \U$15401 ( \15778 , \15776 , \15777 );
nand \U$15402 ( \15779 , \10935 , \9624 );
nand \U$15403 ( \15780 , \15778 , \15779 );
not \U$15404 ( \15781 , \15780 );
or \U$15405 ( \15782 , \15775 , \15781 );
nand \U$15406 ( \15783 , \15208 , \12304 );
nand \U$15407 ( \15784 , \15782 , \15783 );
buf \U$15408 ( \15785 , \15784 );
and \U$15409 ( \15786 , \15774 , \15785 );
and \U$15410 ( \15787 , \15761 , \15772 );
nor \U$15411 ( \15788 , \15786 , \15787 );
not \U$15412 ( \15789 , \15788 );
not \U$15413 ( \15790 , \15789 );
not \U$15414 ( \15791 , \9705 );
not \U$15415 ( \15792 , \15289 );
or \U$15416 ( \15793 , \15791 , \15792 );
not \U$15417 ( \15794 , RIc2262f0_41);
not \U$15418 ( \15795 , \9433 );
or \U$15419 ( \15796 , \15794 , \15795 );
nand \U$15420 ( \15797 , \2014 , \12937 );
nand \U$15421 ( \15798 , \15796 , \15797 );
nand \U$15422 ( \15799 , \15798 , \9690 );
nand \U$15423 ( \15800 , \15793 , \15799 );
not \U$15424 ( \15801 , \15800 );
not \U$15425 ( \15802 , \9129 );
not \U$15426 ( \15803 , \15136 );
or \U$15427 ( \15804 , \15802 , \15803 );
not \U$15428 ( \15805 , RIc226200_43);
not \U$15429 ( \15806 , \2257 );
or \U$15430 ( \15807 , \15805 , \15806 );
nand \U$15431 ( \15808 , \4008 , \9125 );
nand \U$15432 ( \15809 , \15807 , \15808 );
nand \U$15433 ( \15810 , \15809 , \9110 );
nand \U$15434 ( \15811 , \15804 , \15810 );
not \U$15435 ( \15812 , \15811 );
nand \U$15436 ( \15813 , \15801 , \15812 );
not \U$15437 ( \15814 , \9555 );
not \U$15438 ( \15815 , \15126 );
or \U$15439 ( \15816 , \15814 , \15815 );
not \U$15440 ( \15817 , RIc225d50_53);
not \U$15441 ( \15818 , \12961 );
or \U$15442 ( \15819 , \15817 , \15818 );
nand \U$15443 ( \15820 , \1391 , \11585 );
nand \U$15444 ( \15821 , \15819 , \15820 );
nand \U$15445 ( \15822 , \15821 , \8777 );
nand \U$15446 ( \15823 , \15816 , \15822 );
and \U$15447 ( \15824 , \15813 , \15823 );
nor \U$15448 ( \15825 , \15801 , \15812 );
nor \U$15449 ( \15826 , \15824 , \15825 );
not \U$15450 ( \15827 , \15826 );
not \U$15451 ( \15828 , \15827 );
or \U$15452 ( \15829 , \15790 , \15828 );
not \U$15453 ( \15830 , \15826 );
not \U$15454 ( \15831 , \15788 );
or \U$15455 ( \15832 , \15830 , \15831 );
not \U$15456 ( \15833 , \12670 );
not \U$15457 ( \15834 , \15169 );
or \U$15458 ( \15835 , \15833 , \15834 );
and \U$15459 ( \15836 , RIc225a80_59, \4024 );
not \U$15460 ( \15837 , RIc225a80_59);
and \U$15461 ( \15838 , \15837 , \888 );
nor \U$15462 ( \15839 , \15836 , \15838 );
not \U$15463 ( \15840 , \15839 );
nand \U$15464 ( \15841 , \15840 , \15164 );
nand \U$15465 ( \15842 , \15835 , \15841 );
not \U$15466 ( \15843 , \9398 );
not \U$15467 ( \15844 , \15180 );
or \U$15468 ( \15845 , \15843 , \15844 );
not \U$15469 ( \15846 , RIc226110_45);
not \U$15470 ( \15847 , \9570 );
or \U$15471 ( \15848 , \15846 , \15847 );
nand \U$15472 ( \15849 , \5949 , \14660 );
nand \U$15473 ( \15850 , \15848 , \15849 );
nand \U$15474 ( \15851 , \15850 , \9934 );
nand \U$15475 ( \15852 , \15845 , \15851 );
xor \U$15476 ( \15853 , \15842 , \15852 );
not \U$15477 ( \15854 , \11118 );
not \U$15478 ( \15855 , RIc225c60_55);
not \U$15479 ( \15856 , \1170 );
or \U$15480 ( \15857 , \15855 , \15856 );
nand \U$15481 ( \15858 , \11261 , \11041 );
nand \U$15482 ( \15859 , \15857 , \15858 );
not \U$15483 ( \15860 , \15859 );
or \U$15484 ( \15861 , \15854 , \15860 );
nand \U$15485 ( \15862 , \15147 , \13025 );
nand \U$15486 ( \15863 , \15861 , \15862 );
and \U$15487 ( \15864 , \15853 , \15863 );
and \U$15488 ( \15865 , \15842 , \15852 );
or \U$15489 ( \15866 , \15864 , \15865 );
nand \U$15490 ( \15867 , \15832 , \15866 );
nand \U$15491 ( \15868 , \15829 , \15867 );
and \U$15492 ( \15869 , \15750 , \15868 );
and \U$15493 ( \15870 , \15667 , \15749 );
or \U$15494 ( \15871 , \15869 , \15870 );
not \U$15495 ( \15872 , \15871 );
not \U$15496 ( \15873 , \15872 );
xor \U$15497 ( \15874 , \15188 , \15156 );
xnor \U$15498 ( \15875 , \15874 , \15226 );
xor \U$15499 ( \15876 , \15255 , \15243 );
xnor \U$15500 ( \15877 , \15876 , \15295 );
nand \U$15501 ( \15878 , \15875 , \15877 );
xor \U$15502 ( \15879 , \13507 , \13519 );
xor \U$15503 ( \15880 , \15879 , \13532 );
not \U$15504 ( \15881 , \9459 );
not \U$15505 ( \15882 , RIc225e40_51);
not \U$15506 ( \15883 , \1948 );
or \U$15507 ( \15884 , \15882 , \15883 );
nand \U$15508 ( \15885 , \1331 , \9450 );
nand \U$15509 ( \15886 , \15884 , \15885 );
not \U$15510 ( \15887 , \15886 );
or \U$15511 ( \15888 , \15881 , \15887 );
nand \U$15512 ( \15889 , \15399 , \9445 );
nand \U$15513 ( \15890 , \15888 , \15889 );
not \U$15514 ( \15891 , \11965 );
not \U$15515 ( \15892 , RIc225b70_57);
not \U$15516 ( \15893 , \1558 );
or \U$15517 ( \15894 , \15892 , \15893 );
nand \U$15518 ( \15895 , \9995 , \15262 );
nand \U$15519 ( \15896 , \15894 , \15895 );
not \U$15520 ( \15897 , \15896 );
or \U$15521 ( \15898 , \15891 , \15897 );
nand \U$15522 ( \15899 , \15264 , \11974 );
nand \U$15523 ( \15900 , \15898 , \15899 );
xor \U$15524 ( \15901 , \15890 , \15900 );
not \U$15525 ( \15902 , \6307 );
not \U$15526 ( \15903 , \15275 );
or \U$15527 ( \15904 , \15902 , \15903 );
not \U$15528 ( \15905 , RIc2263e0_39);
not \U$15529 ( \15906 , \2556 );
or \U$15530 ( \15907 , \15905 , \15906 );
not \U$15531 ( \15908 , \10899 );
not \U$15532 ( \15909 , \15908 );
nand \U$15533 ( \15910 , \15909 , \8998 );
nand \U$15534 ( \15911 , \15907 , \15910 );
nand \U$15535 ( \15912 , \15911 , \6689 );
nand \U$15536 ( \15913 , \15904 , \15912 );
and \U$15537 ( \15914 , \15901 , \15913 );
and \U$15538 ( \15915 , \15890 , \15900 );
or \U$15539 ( \15916 , \15914 , \15915 );
xor \U$15540 ( \15917 , \15880 , \15916 );
xor \U$15541 ( \15918 , \15474 , \15484 );
xor \U$15542 ( \15919 , \15918 , \15496 );
and \U$15543 ( \15920 , \15917 , \15919 );
and \U$15544 ( \15921 , \15880 , \15916 );
or \U$15545 ( \15922 , \15920 , \15921 );
and \U$15546 ( \15923 , \15878 , \15922 );
nor \U$15547 ( \15924 , \15875 , \15877 );
nor \U$15548 ( \15925 , \15923 , \15924 );
not \U$15549 ( \15926 , \15925 );
or \U$15550 ( \15927 , \15873 , \15926 );
xor \U$15551 ( \15928 , \13356 , \13366 );
xor \U$15552 ( \15929 , \15928 , \13378 );
and \U$15553 ( \15930 , \13432 , \13410 );
not \U$15554 ( \15931 , \13432 );
and \U$15555 ( \15932 , \15931 , \13409 );
or \U$15556 ( \15933 , \15930 , \15932 );
and \U$15557 ( \15934 , \15933 , \13420 );
not \U$15558 ( \15935 , \15933 );
and \U$15559 ( \15936 , \15935 , \13421 );
nor \U$15560 ( \15937 , \15934 , \15936 );
xor \U$15561 ( \15938 , \15929 , \15937 );
not \U$15562 ( \15939 , \5519 );
not \U$15563 ( \15940 , \15386 );
or \U$15564 ( \15941 , \15939 , \15940 );
not \U$15565 ( \15942 , RIc2264d0_37);
not \U$15566 ( \15943 , \12989 );
or \U$15567 ( \15944 , \15942 , \15943 );
nand \U$15568 ( \15945 , \12990 , \4371 );
nand \U$15569 ( \15946 , \15944 , \15945 );
nand \U$15570 ( \15947 , \15946 , \5509 );
nand \U$15571 ( \15948 , \15941 , \15947 );
buf \U$15572 ( \15949 , \15948 );
not \U$15573 ( \15950 , \9552 );
not \U$15574 ( \15951 , \15480 );
or \U$15575 ( \15952 , \15950 , \15951 );
not \U$15576 ( \15953 , RIc225f30_49);
not \U$15577 ( \15954 , \4181 );
or \U$15578 ( \15955 , \15953 , \15954 );
nand \U$15579 ( \15956 , \1729 , \9549 );
nand \U$15580 ( \15957 , \15955 , \15956 );
nand \U$15581 ( \15958 , \15957 , \9534 );
nand \U$15582 ( \15959 , \15952 , \15958 );
or \U$15583 ( \15960 , \15949 , \15959 );
not \U$15584 ( \15961 , \4383 );
not \U$15585 ( \15962 , \15376 );
or \U$15586 ( \15963 , \15961 , \15962 );
and \U$15587 ( \15964 , RIc2265c0_35, \12977 );
not \U$15588 ( \15965 , RIc2265c0_35);
and \U$15589 ( \15966 , \15965 , \11844 );
or \U$15590 ( \15967 , \15964 , \15966 );
nand \U$15591 ( \15968 , \15967 , \4381 );
nand \U$15592 ( \15969 , \15963 , \15968 );
nand \U$15593 ( \15970 , \15960 , \15969 );
nand \U$15594 ( \15971 , \15949 , \15959 );
nand \U$15595 ( \15972 , \15970 , \15971 );
and \U$15596 ( \15973 , \15938 , \15972 );
and \U$15597 ( \15974 , \15929 , \15937 );
or \U$15598 ( \15975 , \15973 , \15974 );
not \U$15599 ( \15976 , \15975 );
xor \U$15600 ( \15977 , \13477 , \13535 );
xnor \U$15601 ( \15978 , \15977 , \13435 );
xor \U$15602 ( \15979 , \13349 , \13384 );
xnor \U$15603 ( \15980 , \15979 , \13381 );
nand \U$15604 ( \15981 , \15978 , \15980 );
not \U$15605 ( \15982 , \15981 );
or \U$15606 ( \15983 , \15976 , \15982 );
not \U$15607 ( \15984 , \15978 );
not \U$15608 ( \15985 , \15980 );
nand \U$15609 ( \15986 , \15984 , \15985 );
nand \U$15610 ( \15987 , \15983 , \15986 );
nand \U$15611 ( \15988 , \15927 , \15987 );
not \U$15612 ( \15989 , \15872 );
not \U$15613 ( \15990 , \15925 );
nand \U$15614 ( \15991 , \15989 , \15990 );
nand \U$15615 ( \15992 , \15988 , \15991 );
not \U$15616 ( \15993 , \15992 );
not \U$15617 ( \15994 , \15993 );
not \U$15618 ( \15995 , \15105 );
not \U$15619 ( \15996 , \15306 );
not \U$15620 ( \15997 , \15996 );
or \U$15621 ( \15998 , \15995 , \15997 );
not \U$15622 ( \15999 , \15305 );
not \U$15623 ( \16000 , \15304 );
or \U$15624 ( \16001 , \15999 , \16000 );
not \U$15625 ( \16002 , \15105 );
nand \U$15626 ( \16003 , \16001 , \16002 );
nand \U$15627 ( \16004 , \15998 , \16003 );
not \U$15628 ( \16005 , \15117 );
and \U$15629 ( \16006 , \16004 , \16005 );
not \U$15630 ( \16007 , \16004 );
and \U$15631 ( \16008 , \16007 , \15117 );
nor \U$15632 ( \16009 , \16006 , \16008 );
not \U$15633 ( \16010 , \16009 );
or \U$15634 ( \16011 , \15994 , \16010 );
not \U$15635 ( \16012 , \15303 );
not \U$15636 ( \16013 , \15299 );
not \U$15637 ( \16014 , \16013 );
or \U$15638 ( \16015 , \16012 , \16014 );
nand \U$15639 ( \16016 , \15299 , \15302 );
nand \U$15640 ( \16017 , \16015 , \16016 );
buf \U$15641 ( \16018 , \15228 );
xor \U$15642 ( \16019 , \16017 , \16018 );
not \U$15643 ( \16020 , \16019 );
and \U$15644 ( \16021 , \15417 , \15334 );
not \U$15645 ( \16022 , \15417 );
and \U$15646 ( \16023 , \16022 , \15333 );
nor \U$15647 ( \16024 , \16021 , \16023 );
xor \U$15648 ( \16025 , \16024 , \15361 );
not \U$15649 ( \16026 , \16025 );
not \U$15650 ( \16027 , \16026 );
or \U$15651 ( \16028 , \16020 , \16027 );
not \U$15652 ( \16029 , \16019 );
not \U$15653 ( \16030 , \16029 );
not \U$15654 ( \16031 , \16025 );
or \U$15655 ( \16032 , \16030 , \16031 );
xor \U$15656 ( \16033 , \15151 , \15131 );
xnor \U$15657 ( \16034 , \16033 , \15140 );
xor \U$15658 ( \16035 , \15173 , \15163 );
xnor \U$15659 ( \16036 , \16035 , \15185 );
nand \U$15660 ( \16037 , \16034 , \16036 );
xor \U$15661 ( \16038 , \13491 , \12848 );
xor \U$15662 ( \16039 , \16038 , \13504 );
not \U$15663 ( \16040 , \1040 );
not \U$15664 ( \16041 , RIc2274c0_3);
not \U$15665 ( \16042 , \12755 );
not \U$15666 ( \16043 , \16042 );
or \U$15667 ( \16044 , \16041 , \16043 );
nand \U$15668 ( \16045 , \12755 , \1032 );
nand \U$15669 ( \16046 , \16044 , \16045 );
not \U$15670 ( \16047 , \16046 );
or \U$15671 ( \16048 , \16040 , \16047 );
nand \U$15672 ( \16049 , \13502 , \1081 );
nand \U$15673 ( \16050 , \16048 , \16049 );
not \U$15674 ( \16051 , \954 );
not \U$15675 ( \16052 , \15458 );
or \U$15676 ( \16053 , \16051 , \16052 );
not \U$15677 ( \16054 , RIc2273d0_5);
not \U$15678 ( \16055 , \10198 );
or \U$15679 ( \16056 , \16054 , \16055 );
nand \U$15680 ( \16057 , \10197 , \935 );
nand \U$15681 ( \16058 , \16056 , \16057 );
nand \U$15682 ( \16059 , \16058 , \950 );
nand \U$15683 ( \16060 , \16053 , \16059 );
xor \U$15684 ( \16061 , \16050 , \16060 );
not \U$15685 ( \16062 , \9904 );
not \U$15686 ( \16063 , RIc227100_11);
not \U$15687 ( \16064 , \10814 );
or \U$15688 ( \16065 , \16063 , \16064 );
nand \U$15689 ( \16066 , \10110 , \1302 );
nand \U$15690 ( \16067 , \16065 , \16066 );
not \U$15691 ( \16068 , \16067 );
or \U$15692 ( \16069 , \16062 , \16068 );
nand \U$15693 ( \16070 , \15467 , \1310 );
nand \U$15694 ( \16071 , \16069 , \16070 );
and \U$15695 ( \16072 , \16061 , \16071 );
and \U$15696 ( \16073 , \16050 , \16060 );
or \U$15697 ( \16074 , \16072 , \16073 );
xor \U$15698 ( \16075 , \16039 , \16074 );
not \U$15699 ( \16076 , \3631 );
not \U$15700 ( \16077 , \15492 );
or \U$15701 ( \16078 , \16076 , \16077 );
and \U$15702 ( \16079 , \2634 , \5179 );
not \U$15703 ( \16080 , \2634 );
and \U$15704 ( \16081 , \16080 , RIc2266b0_33);
or \U$15705 ( \16082 , \16079 , \16081 );
nand \U$15706 ( \16083 , \16082 , \3629 );
nand \U$15707 ( \16084 , \16078 , \16083 );
and \U$15708 ( \16085 , \16075 , \16084 );
and \U$15709 ( \16086 , \16039 , \16074 );
or \U$15710 ( \16087 , \16085 , \16086 );
and \U$15711 ( \16088 , \16037 , \16087 );
nor \U$15712 ( \16089 , \16034 , \16036 );
nor \U$15713 ( \16090 , \16088 , \16089 );
not \U$15714 ( \16091 , \16090 );
xor \U$15715 ( \16092 , \15293 , \15279 );
not \U$15716 ( \16093 , \15269 );
and \U$15717 ( \16094 , \16092 , \16093 );
not \U$15718 ( \16095 , \16092 );
and \U$15719 ( \16096 , \16095 , \15269 );
nor \U$15720 ( \16097 , \16094 , \16096 );
xor \U$15721 ( \16098 , \15403 , \15391 );
xnor \U$15722 ( \16099 , \16098 , \15378 );
nand \U$15723 ( \16100 , \16097 , \16099 );
xor \U$15724 ( \16101 , \15201 , \15210 );
xor \U$15725 ( \16102 , \16101 , \15223 );
and \U$15726 ( \16103 , \16100 , \16102 );
nor \U$15727 ( \16104 , \16099 , \16097 );
nor \U$15728 ( \16105 , \16103 , \16104 );
not \U$15729 ( \16106 , \16105 );
or \U$15730 ( \16107 , \16091 , \16106 );
xor \U$15731 ( \16108 , \15410 , \15407 );
xnor \U$15732 ( \16109 , \16108 , \15413 );
nand \U$15733 ( \16110 , \16107 , \16109 );
not \U$15734 ( \16111 , \16090 );
not \U$15735 ( \16112 , \16105 );
nand \U$15736 ( \16113 , \16111 , \16112 );
nand \U$15737 ( \16114 , \16110 , \16113 );
not \U$15738 ( \16115 , \16114 );
not \U$15739 ( \16116 , \16115 );
nand \U$15740 ( \16117 , \16032 , \16116 );
nand \U$15741 ( \16118 , \16028 , \16117 );
nand \U$15742 ( \16119 , \16011 , \16118 );
not \U$15743 ( \16120 , \16009 );
nand \U$15744 ( \16121 , \16120 , \15992 );
nand \U$15745 ( \16122 , \16119 , \16121 );
not \U$15746 ( \16123 , \15308 );
not \U$15747 ( \16124 , \15311 );
or \U$15748 ( \16125 , \16123 , \16124 );
or \U$15749 ( \16126 , \15308 , \15311 );
nand \U$15750 ( \16127 , \16125 , \16126 );
and \U$15751 ( \16128 , \16127 , \15315 );
not \U$15752 ( \16129 , \16127 );
not \U$15753 ( \16130 , \15315 );
and \U$15754 ( \16131 , \16129 , \16130 );
nor \U$15755 ( \16132 , \16128 , \16131 );
xor \U$15756 ( \16133 , \16122 , \16132 );
xor \U$15757 ( \16134 , \15544 , \15546 );
xor \U$15758 ( \16135 , \16134 , \15549 );
xor \U$15759 ( \16136 , \15420 , \15507 );
xor \U$15760 ( \16137 , \16136 , \15516 );
or \U$15761 ( \16138 , \16135 , \16137 );
xor \U$15762 ( \16139 , \15422 , \15424 );
xor \U$15763 ( \16140 , \16139 , \15504 );
xor \U$15764 ( \16141 , \15667 , \15749 );
xor \U$15765 ( \16142 , \16141 , \15868 );
not \U$15766 ( \16143 , \16142 );
not \U$15767 ( \16144 , \15499 );
not \U$15768 ( \16145 , \16144 );
not \U$15769 ( \16146 , \15502 );
or \U$15770 ( \16147 , \16145 , \16146 );
nand \U$15771 ( \16148 , \15437 , \15499 );
nand \U$15772 ( \16149 , \16147 , \16148 );
and \U$15773 ( \16150 , \16149 , \15427 );
not \U$15774 ( \16151 , \16149 );
and \U$15775 ( \16152 , \16151 , \15501 );
nor \U$15776 ( \16153 , \16150 , \16152 );
not \U$15777 ( \16154 , \15344 );
not \U$15778 ( \16155 , \15357 );
or \U$15779 ( \16156 , \16154 , \16155 );
or \U$15780 ( \16157 , \15357 , \15344 );
nand \U$15781 ( \16158 , \16156 , \16157 );
buf \U$15782 ( \16159 , \15346 );
and \U$15783 ( \16160 , \16158 , \16159 );
not \U$15784 ( \16161 , \16158 );
not \U$15785 ( \16162 , \16159 );
and \U$15786 ( \16163 , \16161 , \16162 );
nor \U$15787 ( \16164 , \16160 , \16163 );
nand \U$15788 ( \16165 , \16153 , \16164 );
not \U$15789 ( \16166 , \16165 );
or \U$15790 ( \16167 , \16143 , \16166 );
not \U$15791 ( \16168 , \16153 );
not \U$15792 ( \16169 , \16164 );
nand \U$15793 ( \16170 , \16168 , \16169 );
nand \U$15794 ( \16171 , \16167 , \16170 );
xor \U$15795 ( \16172 , \16140 , \16171 );
not \U$15796 ( \16173 , \15524 );
not \U$15797 ( \16174 , \15542 );
or \U$15798 ( \16175 , \16173 , \16174 );
or \U$15799 ( \16176 , \15542 , \15524 );
nand \U$15800 ( \16177 , \16175 , \16176 );
xor \U$15801 ( \16178 , \15539 , \16177 );
and \U$15802 ( \16179 , \16172 , \16178 );
and \U$15803 ( \16180 , \16140 , \16171 );
or \U$15804 ( \16181 , \16179 , \16180 );
nand \U$15805 ( \16182 , \16138 , \16181 );
nand \U$15806 ( \16183 , \16135 , \16137 );
nand \U$15807 ( \16184 , \16182 , \16183 );
and \U$15808 ( \16185 , \16133 , \16184 );
and \U$15809 ( \16186 , \16122 , \16132 );
or \U$15810 ( \16187 , \16185 , \16186 );
xor \U$15811 ( \16188 , \15574 , \16187 );
xor \U$15812 ( \16189 , \15320 , \15322 );
xor \U$15813 ( \16190 , \16189 , \15565 );
and \U$15814 ( \16191 , \16188 , \16190 );
and \U$15815 ( \16192 , \15574 , \16187 );
or \U$15816 ( \16193 , \16191 , \16192 );
nor \U$15817 ( \16194 , \15572 , \16193 );
not \U$15818 ( \16195 , \16194 );
xor \U$15819 ( \16196 , \15574 , \16187 );
xor \U$15820 ( \16197 , \16196 , \16190 );
not \U$15821 ( \16198 , \16197 );
xor \U$15822 ( \16199 , \15519 , \15552 );
xor \U$15823 ( \16200 , \16199 , \15562 );
xor \U$15824 ( \16201 , \16122 , \16132 );
xor \U$15825 ( \16202 , \16201 , \16184 );
xor \U$15826 ( \16203 , \16200 , \16202 );
not \U$15827 ( \16204 , \15871 );
not \U$15828 ( \16205 , \15987 );
not \U$15829 ( \16206 , \16205 );
or \U$15830 ( \16207 , \16204 , \16206 );
nand \U$15831 ( \16208 , \15872 , \15987 );
nand \U$15832 ( \16209 , \16207 , \16208 );
not \U$15833 ( \16210 , \15990 );
and \U$15834 ( \16211 , \16209 , \16210 );
not \U$15835 ( \16212 , \16209 );
and \U$15836 ( \16213 , \16212 , \15990 );
nor \U$15837 ( \16214 , \16211 , \16213 );
not \U$15838 ( \16215 , \16214 );
not \U$15839 ( \16216 , \16215 );
and \U$15840 ( \16217 , \16019 , \16114 );
not \U$15841 ( \16218 , \16019 );
and \U$15842 ( \16219 , \16218 , \16115 );
nor \U$15843 ( \16220 , \16217 , \16219 );
and \U$15844 ( \16221 , \16220 , \16026 );
not \U$15845 ( \16222 , \16220 );
and \U$15846 ( \16223 , \16222 , \16025 );
nor \U$15847 ( \16224 , \16221 , \16223 );
not \U$15848 ( \16225 , \16224 );
or \U$15849 ( \16226 , \16216 , \16225 );
or \U$15850 ( \16227 , \16224 , \16215 );
xor \U$15851 ( \16228 , \15842 , \15852 );
xor \U$15852 ( \16229 , \16228 , \15863 );
not \U$15853 ( \16230 , \16229 );
xor \U$15854 ( \16231 , \15784 , \15772 );
and \U$15855 ( \16232 , \16231 , \15761 );
not \U$15856 ( \16233 , \16231 );
and \U$15857 ( \16234 , \16233 , \15762 );
nor \U$15858 ( \16235 , \16232 , \16234 );
not \U$15859 ( \16236 , \16235 );
nand \U$15860 ( \16237 , \16230 , \16236 );
not \U$15861 ( \16238 , \1081 );
not \U$15862 ( \16239 , \16046 );
or \U$15863 ( \16240 , \16238 , \16239 );
and \U$15864 ( \16241 , RIc2274c0_3, \15443 );
not \U$15865 ( \16242 , RIc2274c0_3);
and \U$15866 ( \16243 , \16242 , \15444 );
nor \U$15867 ( \16244 , \16241 , \16243 );
nand \U$15868 ( \16245 , \16244 , \1040 );
nand \U$15869 ( \16246 , \16240 , \16245 );
xor \U$15870 ( \16247 , RIc229518_128, RIc22b318_192);
buf \U$15871 ( \16248 , \16247 );
and \U$15872 ( \16249 , RIc2275b0_1, \16248 );
not \U$15873 ( \16250 , \898 );
xor \U$15874 ( \16251 , \13487 , RIc2275b0_1);
not \U$15875 ( \16252 , \16251 );
or \U$15876 ( \16253 , \16250 , \16252 );
xor \U$15877 ( \16254 , RIc2294a0_127, RIc22b2a0_191);
xnor \U$15878 ( \16255 , \16254 , \487 );
buf \U$15879 ( \16256 , \16255 );
and \U$15880 ( \16257 , RIc2275b0_1, \16256 );
not \U$15881 ( \16258 , RIc2275b0_1);
not \U$15882 ( \16259 , \16256 );
and \U$15883 ( \16260 , \16258 , \16259 );
nor \U$15884 ( \16261 , \16257 , \16260 );
nand \U$15885 ( \16262 , \16261 , \853 );
nand \U$15886 ( \16263 , \16253 , \16262 );
xor \U$15887 ( \16264 , \16249 , \16263 );
not \U$15888 ( \16265 , \1040 );
not \U$15889 ( \16266 , RIc2274c0_3);
not \U$15890 ( \16267 , \15630 );
or \U$15891 ( \16268 , \16266 , \16267 );
nand \U$15892 ( \16269 , \12845 , \2896 );
nand \U$15893 ( \16270 , \16268 , \16269 );
not \U$15894 ( \16271 , \16270 );
or \U$15895 ( \16272 , \16265 , \16271 );
nand \U$15896 ( \16273 , \16244 , \1081 );
nand \U$15897 ( \16274 , \16272 , \16273 );
and \U$15898 ( \16275 , \16264 , \16274 );
and \U$15899 ( \16276 , \16249 , \16263 );
or \U$15900 ( \16277 , \16275 , \16276 );
xor \U$15901 ( \16278 , \16246 , \16277 );
not \U$15902 ( \16279 , \1682 );
not \U$15903 ( \16280 , RIc227010_13);
not \U$15904 ( \16281 , \10643 );
or \U$15905 ( \16282 , \16280 , \16281 );
nand \U$15906 ( \16283 , \9050 , \1758 );
nand \U$15907 ( \16284 , \16282 , \16283 );
not \U$15908 ( \16285 , \16284 );
or \U$15909 ( \16286 , \16279 , \16285 );
not \U$15910 ( \16287 , RIc227010_13);
not \U$15911 ( \16288 , \9076 );
or \U$15912 ( \16289 , \16287 , \16288 );
nand \U$15913 ( \16290 , \9072 , \1296 );
nand \U$15914 ( \16291 , \16289 , \16290 );
nand \U$15915 ( \16292 , \16291 , \1678 );
nand \U$15916 ( \16293 , \16286 , \16292 );
and \U$15917 ( \16294 , \16278 , \16293 );
and \U$15918 ( \16295 , \16246 , \16277 );
or \U$15919 ( \16296 , \16294 , \16295 );
not \U$15920 ( \16297 , \9444 );
not \U$15921 ( \16298 , \15886 );
or \U$15922 ( \16299 , \16297 , \16298 );
not \U$15923 ( \16300 , RIc225e40_51);
not \U$15924 ( \16301 , \3783 );
or \U$15925 ( \16302 , \16300 , \16301 );
nand \U$15926 ( \16303 , \10678 , \9450 );
nand \U$15927 ( \16304 , \16302 , \16303 );
nand \U$15928 ( \16305 , \16304 , \9458 );
nand \U$15929 ( \16306 , \16299 , \16305 );
xor \U$15930 ( \16307 , \16296 , \16306 );
not \U$15931 ( \16308 , \5135 );
not \U$15932 ( \16309 , \15967 );
or \U$15933 ( \16310 , \16308 , \16309 );
not \U$15934 ( \16311 , RIc2265c0_35);
not \U$15935 ( \16312 , \2731 );
or \U$15936 ( \16313 , \16311 , \16312 );
not \U$15937 ( \16314 , RIc2265c0_35);
nand \U$15938 ( \16315 , \15490 , \16314 );
nand \U$15939 ( \16316 , \16313 , \16315 );
nand \U$15940 ( \16317 , \16316 , \5741 );
nand \U$15941 ( \16318 , \16310 , \16317 );
and \U$15942 ( \16319 , \16307 , \16318 );
and \U$15943 ( \16320 , \16296 , \16306 );
or \U$15944 ( \16321 , \16319 , \16320 );
and \U$15945 ( \16322 , \16237 , \16321 );
and \U$15946 ( \16323 , \16229 , \16235 );
nor \U$15947 ( \16324 , \16322 , \16323 );
not \U$15948 ( \16325 , \16324 );
xor \U$15949 ( \16326 , \15948 , \15969 );
xnor \U$15950 ( \16327 , \16326 , \15959 );
not \U$15951 ( \16328 , \15823 );
not \U$15952 ( \16329 , \15812 );
or \U$15953 ( \16330 , \16328 , \16329 );
not \U$15954 ( \16331 , \15823 );
nand \U$15955 ( \16332 , \16331 , \15811 );
nand \U$15956 ( \16333 , \16330 , \16332 );
and \U$15957 ( \16334 , \16333 , \15801 );
not \U$15958 ( \16335 , \16333 );
and \U$15959 ( \16336 , \16335 , \15800 );
nor \U$15960 ( \16337 , \16334 , \16336 );
nand \U$15961 ( \16338 , \16327 , \16337 );
xor \U$15962 ( \16339 , \15890 , \15900 );
xor \U$15963 ( \16340 , \16339 , \15913 );
and \U$15964 ( \16341 , \16338 , \16340 );
nor \U$15965 ( \16342 , \16327 , \16337 );
nor \U$15966 ( \16343 , \16341 , \16342 );
not \U$15967 ( \16344 , \16343 );
or \U$15968 ( \16345 , \16325 , \16344 );
xor \U$15969 ( \16346 , \15929 , \15937 );
xor \U$15970 ( \16347 , \16346 , \15972 );
nand \U$15971 ( \16348 , \16345 , \16347 );
not \U$15972 ( \16349 , \16343 );
not \U$15973 ( \16350 , \16324 );
nand \U$15974 ( \16351 , \16349 , \16350 );
nand \U$15975 ( \16352 , \16348 , \16351 );
not \U$15976 ( \16353 , \16352 );
xor \U$15977 ( \16354 , \15576 , \15617 );
xor \U$15978 ( \16355 , \16354 , \15665 );
not \U$15979 ( \16356 , \16355 );
not \U$15980 ( \16357 , \3631 );
not \U$15981 ( \16358 , \16082 );
or \U$15982 ( \16359 , \16357 , \16358 );
not \U$15983 ( \16360 , RIc2266b0_33);
and \U$15984 ( \16361 , \2103 , \16360 );
not \U$15985 ( \16362 , \2103 );
and \U$15986 ( \16363 , \16362 , RIc2266b0_33);
or \U$15987 ( \16364 , \16361 , \16363 );
nand \U$15988 ( \16365 , \16364 , \3629 );
nand \U$15989 ( \16366 , \16359 , \16365 );
not \U$15990 ( \16367 , \16366 );
not \U$15991 ( \16368 , \2320 );
not \U$15992 ( \16369 , RIc226f20_15);
not \U$15993 ( \16370 , \12403 );
or \U$15994 ( \16371 , \16369 , \16370 );
nand \U$15995 ( \16372 , \12406 , \1674 );
nand \U$15996 ( \16373 , \16371 , \16372 );
not \U$15997 ( \16374 , \16373 );
or \U$15998 ( \16375 , \16368 , \16374 );
nand \U$15999 ( \16376 , \15716 , \2358 );
nand \U$16000 ( \16377 , \16375 , \16376 );
not \U$16001 ( \16378 , \16377 );
nand \U$16002 ( \16379 , \16367 , \16378 );
not \U$16003 ( \16380 , \9534 );
and \U$16004 ( \16381 , \9700 , RIc225f30_49);
not \U$16005 ( \16382 , \9700 );
and \U$16006 ( \16383 , \16382 , \11289 );
or \U$16007 ( \16384 , \16381 , \16383 );
not \U$16008 ( \16385 , \16384 );
or \U$16009 ( \16386 , \16380 , \16385 );
nand \U$16010 ( \16387 , \15957 , \9552 );
nand \U$16011 ( \16388 , \16386 , \16387 );
and \U$16012 ( \16389 , \16379 , \16388 );
and \U$16013 ( \16390 , \16366 , \16377 );
nor \U$16014 ( \16391 , \16389 , \16390 );
not \U$16015 ( \16392 , \15719 );
not \U$16016 ( \16393 , RIc225990_61);
not \U$16017 ( \16394 , \9491 );
or \U$16018 ( \16395 , \16393 , \16394 );
nand \U$16019 ( \16396 , \1072 , \12806 );
nand \U$16020 ( \16397 , \16395 , \16396 );
not \U$16021 ( \16398 , \16397 );
or \U$16022 ( \16399 , \16392 , \16398 );
nand \U$16023 ( \16400 , \15726 , \15729 );
nand \U$16024 ( \16401 , \16399 , \16400 );
not \U$16025 ( \16402 , \16401 );
not \U$16026 ( \16403 , \2711 );
not \U$16027 ( \16404 , \15759 );
or \U$16028 ( \16405 , \16403 , \16404 );
not \U$16029 ( \16406 , RIc2267a0_31);
not \U$16030 ( \16407 , \3726 );
or \U$16031 ( \16408 , \16406 , \16407 );
nand \U$16032 ( \16409 , \2980 , \3648 );
nand \U$16033 ( \16410 , \16408 , \16409 );
nand \U$16034 ( \16411 , \16410 , \2697 );
nand \U$16035 ( \16412 , \16405 , \16411 );
not \U$16036 ( \16413 , \16412 );
or \U$16037 ( \16414 , \16402 , \16413 );
or \U$16038 ( \16415 , \16412 , \16401 );
not \U$16039 ( \16416 , \9641 );
not \U$16040 ( \16417 , RIc226020_47);
not \U$16041 ( \16418 , \3686 );
or \U$16042 ( \16419 , \16417 , \16418 );
not \U$16043 ( \16420 , \13914 );
nand \U$16044 ( \16421 , \16420 , \9373 );
nand \U$16045 ( \16422 , \16419 , \16421 );
not \U$16046 ( \16423 , \16422 );
or \U$16047 ( \16424 , \16416 , \16423 );
nand \U$16048 ( \16425 , \15780 , \9619 );
nand \U$16049 ( \16426 , \16424 , \16425 );
nand \U$16050 ( \16427 , \16415 , \16426 );
nand \U$16051 ( \16428 , \16414 , \16427 );
not \U$16052 ( \16429 , \16428 );
xor \U$16053 ( \16430 , \16391 , \16429 );
not \U$16054 ( \16431 , \15839 );
not \U$16055 ( \16432 , \12670 );
not \U$16056 ( \16433 , \16432 );
and \U$16057 ( \16434 , \16431 , \16433 );
and \U$16058 ( \16435 , RIc225a80_59, \4608 );
not \U$16059 ( \16436 , RIc225a80_59);
and \U$16060 ( \16437 , \16436 , \840 );
nor \U$16061 ( \16438 , \16435 , \16437 );
not \U$16062 ( \16439 , \15164 );
nor \U$16063 ( \16440 , \16438 , \16439 );
nor \U$16064 ( \16441 , \16434 , \16440 );
not \U$16065 ( \16442 , \1988 );
not \U$16066 ( \16443 , \9125 );
and \U$16067 ( \16444 , \16442 , \16443 );
and \U$16068 ( \16445 , \12509 , \12456 );
nor \U$16069 ( \16446 , \16444 , \16445 );
not \U$16070 ( \16447 , \16446 );
not \U$16071 ( \16448 , \9109 );
and \U$16072 ( \16449 , \16447 , \16448 );
and \U$16073 ( \16450 , \15809 , \9129 );
nor \U$16074 ( \16451 , \16449 , \16450 );
xor \U$16075 ( \16452 , \16441 , \16451 );
and \U$16076 ( \16453 , RIc2262f0_41, \9422 );
not \U$16077 ( \16454 , RIc2262f0_41);
not \U$16078 ( \16455 , \2591 );
and \U$16079 ( \16456 , \16454 , \16455 );
nor \U$16080 ( \16457 , \16453 , \16456 );
not \U$16081 ( \16458 , \16457 );
not \U$16082 ( \16459 , \9690 );
not \U$16083 ( \16460 , \16459 );
and \U$16084 ( \16461 , \16458 , \16460 );
and \U$16085 ( \16462 , \15798 , \9816 );
nor \U$16086 ( \16463 , \16461 , \16462 );
and \U$16087 ( \16464 , \16452 , \16463 );
and \U$16088 ( \16465 , \16441 , \16451 );
or \U$16089 ( \16466 , \16464 , \16465 );
and \U$16090 ( \16467 , \16430 , \16466 );
and \U$16091 ( \16468 , \16391 , \16429 );
or \U$16092 ( \16469 , \16467 , \16468 );
not \U$16093 ( \16470 , \16469 );
or \U$16094 ( \16471 , \16356 , \16470 );
xor \U$16095 ( \16472 , \15669 , \15707 );
xor \U$16096 ( \16473 , \16472 , \15746 );
buf \U$16097 ( \16474 , \16473 );
nand \U$16098 ( \16475 , \16471 , \16474 );
not \U$16099 ( \16476 , \16469 );
not \U$16100 ( \16477 , \16355 );
nand \U$16101 ( \16478 , \16476 , \16477 );
nand \U$16102 ( \16479 , \16475 , \16478 );
buf \U$16103 ( \16480 , \16479 );
not \U$16104 ( \16481 , \16480 );
buf \U$16105 ( \16482 , \16256 );
and \U$16106 ( \16483 , \16482 , RIc2275b0_1);
not \U$16107 ( \16484 , \898 );
not \U$16108 ( \16485 , \15635 );
or \U$16109 ( \16486 , \16484 , \16485 );
nand \U$16110 ( \16487 , \16251 , \853 );
nand \U$16111 ( \16488 , \16486 , \16487 );
xor \U$16112 ( \16489 , \16483 , \16488 );
not \U$16113 ( \16490 , \950 );
not \U$16114 ( \16491 , RIc2273d0_5);
not \U$16115 ( \16492 , \10355 );
not \U$16116 ( \16493 , \16492 );
or \U$16117 ( \16494 , \16491 , \16493 );
nand \U$16118 ( \16495 , \13497 , \946 );
nand \U$16119 ( \16496 , \16494 , \16495 );
not \U$16120 ( \16497 , \16496 );
or \U$16121 ( \16498 , \16490 , \16497 );
nand \U$16122 ( \16499 , \16058 , \954 );
nand \U$16123 ( \16500 , \16498 , \16499 );
and \U$16124 ( \16501 , \16489 , \16500 );
and \U$16125 ( \16502 , \16483 , \16488 );
or \U$16126 ( \16503 , \16501 , \16502 );
not \U$16127 ( \16504 , \2154 );
not \U$16128 ( \16505 , \15658 );
or \U$16129 ( \16506 , \16504 , \16505 );
not \U$16130 ( \16507 , RIc226980_27);
not \U$16131 ( \16508 , \10230 );
or \U$16132 ( \16509 , \16507 , \16508 );
not \U$16133 ( \16510 , RIc226980_27);
nand \U$16134 ( \16511 , \9757 , \16510 );
nand \U$16135 ( \16512 , \16509 , \16511 );
nand \U$16136 ( \16513 , \16512 , \2138 );
nand \U$16137 ( \16514 , \16506 , \16513 );
xor \U$16138 ( \16515 , \16503 , \16514 );
not \U$16139 ( \16516 , \9142 );
not \U$16140 ( \16517 , \15770 );
or \U$16141 ( \16518 , \16516 , \16517 );
not \U$16142 ( \16519 , \4413 );
xor \U$16143 ( \16520 , RIc226890_29, \16519 );
nand \U$16144 ( \16521 , \16520 , \2784 );
nand \U$16145 ( \16522 , \16518 , \16521 );
and \U$16146 ( \16523 , \16515 , \16522 );
and \U$16147 ( \16524 , \16503 , \16514 );
or \U$16148 ( \16525 , \16523 , \16524 );
not \U$16149 ( \16526 , \2367 );
not \U$16150 ( \16527 , \15702 );
or \U$16151 ( \16528 , \16526 , \16527 );
and \U$16152 ( \16529 , \3204 , \9884 );
not \U$16153 ( \16530 , \3204 );
not \U$16154 ( \16531 , \8885 );
not \U$16155 ( \16532 , \16531 );
and \U$16156 ( \16533 , \16530 , \16532 );
or \U$16157 ( \16534 , \16529 , \16533 );
not \U$16158 ( \16535 , \16534 );
nand \U$16159 ( \16536 , \16535 , \2392 );
nand \U$16160 ( \16537 , \16528 , \16536 );
not \U$16161 ( \16538 , \16537 );
not \U$16162 ( \16539 , \10214 );
not \U$16163 ( \16540 , RIc226b60_23);
not \U$16164 ( \16541 , \6719 );
or \U$16165 ( \16542 , \16540 , \16541 );
not \U$16166 ( \16543 , \9859 );
nand \U$16167 ( \16544 , \16543 , \1919 );
nand \U$16168 ( \16545 , \16542 , \16544 );
not \U$16169 ( \16546 , \16545 );
or \U$16170 ( \16547 , \16539 , \16546 );
nand \U$16171 ( \16548 , \15647 , \5365 );
nand \U$16172 ( \16549 , \16547 , \16548 );
not \U$16173 ( \16550 , \16549 );
or \U$16174 ( \16551 , \16538 , \16550 );
or \U$16175 ( \16552 , \16537 , \16549 );
not \U$16176 ( \16553 , \2195 );
not \U$16177 ( \16554 , RIc226a70_25);
not \U$16178 ( \16555 , \6070 );
not \U$16179 ( \16556 , \16555 );
or \U$16180 ( \16557 , \16554 , \16556 );
nand \U$16181 ( \16558 , \9769 , \2187 );
nand \U$16182 ( \16559 , \16557 , \16558 );
not \U$16183 ( \16560 , \16559 );
or \U$16184 ( \16561 , \16553 , \16560 );
nand \U$16185 ( \16562 , \15607 , \2172 );
nand \U$16186 ( \16563 , \16561 , \16562 );
nand \U$16187 ( \16564 , \16552 , \16563 );
nand \U$16188 ( \16565 , \16551 , \16564 );
not \U$16189 ( \16566 , \16565 );
and \U$16190 ( \16567 , \15740 , \1682 );
not \U$16191 ( \16568 , \16284 );
nor \U$16192 ( \16569 , \16568 , \1679 );
nor \U$16193 ( \16570 , \16567 , \16569 );
not \U$16194 ( \16571 , \16570 );
not \U$16195 ( \16572 , \16571 );
not \U$16196 ( \16573 , \1118 );
and \U$16197 ( \16574 , \9324 , \940 );
not \U$16198 ( \16575 , \9324 );
and \U$16199 ( \16576 , \16575 , RIc2272e0_7);
or \U$16200 ( \16577 , \16574 , \16576 );
not \U$16201 ( \16578 , \16577 );
or \U$16202 ( \16579 , \16573 , \16578 );
nand \U$16203 ( \16580 , \15593 , \1121 );
nand \U$16204 ( \16581 , \16579 , \16580 );
not \U$16205 ( \16582 , \16581 );
not \U$16206 ( \16583 , \1363 );
not \U$16207 ( \16584 , RIc2271f0_9);
not \U$16208 ( \16585 , \10800 );
or \U$16209 ( \16586 , \16584 , \16585 );
nand \U$16210 ( \16587 , \9274 , \1351 );
nand \U$16211 ( \16588 , \16586 , \16587 );
not \U$16212 ( \16589 , \16588 );
or \U$16213 ( \16590 , \16583 , \16589 );
nand \U$16214 ( \16591 , \15583 , \1339 );
nand \U$16215 ( \16592 , \16590 , \16591 );
not \U$16216 ( \16593 , \16592 );
nand \U$16217 ( \16594 , \16582 , \16593 );
not \U$16218 ( \16595 , \16594 );
or \U$16219 ( \16596 , \16572 , \16595 );
nand \U$16220 ( \16597 , \16592 , \16581 );
nand \U$16221 ( \16598 , \16596 , \16597 );
not \U$16222 ( \16599 , \16598 );
nand \U$16223 ( \16600 , \16566 , \16599 );
and \U$16224 ( \16601 , \16525 , \16600 );
nor \U$16225 ( \16602 , \16566 , \16599 );
nor \U$16226 ( \16603 , \16601 , \16602 );
xor \U$16227 ( \16604 , \15627 , \15639 );
not \U$16228 ( \16605 , \2518 );
not \U$16229 ( \16606 , RIc226d40_19);
not \U$16230 ( \16607 , \9900 );
or \U$16231 ( \16608 , \16606 , \16607 );
nand \U$16232 ( \16609 , \9901 , \3338 );
nand \U$16233 ( \16610 , \16608 , \16609 );
not \U$16234 ( \16611 , \16610 );
or \U$16235 ( \16612 , \16605 , \16611 );
nand \U$16236 ( \16613 , \2534 , \15675 );
nand \U$16237 ( \16614 , \16612 , \16613 );
xor \U$16238 ( \16615 , \16604 , \16614 );
not \U$16239 ( \16616 , \1945 );
and \U$16240 ( \16617 , RIc226e30_17, \11566 );
not \U$16241 ( \16618 , RIc226e30_17);
and \U$16242 ( \16619 , \16618 , \8952 );
or \U$16243 ( \16620 , \16617 , \16619 );
not \U$16244 ( \16621 , \16620 );
or \U$16245 ( \16622 , \16616 , \16621 );
nand \U$16246 ( \16623 , \15687 , \1963 );
nand \U$16247 ( \16624 , \16622 , \16623 );
and \U$16248 ( \16625 , \16615 , \16624 );
and \U$16249 ( \16626 , \16604 , \16614 );
or \U$16250 ( \16627 , \16625 , \16626 );
xor \U$16251 ( \16628 , \15450 , \15460 );
xor \U$16252 ( \16629 , \16628 , \15471 );
xor \U$16253 ( \16630 , \15587 , \15597 );
xor \U$16254 ( \16631 , \16630 , \15609 );
or \U$16255 ( \16632 , \16629 , \16631 );
and \U$16256 ( \16633 , \16627 , \16632 );
and \U$16257 ( \16634 , \16631 , \16629 );
nor \U$16258 ( \16635 , \16633 , \16634 );
nand \U$16259 ( \16636 , \16603 , \16635 );
not \U$16260 ( \16637 , \16636 );
not \U$16261 ( \16638 , \5509 );
not \U$16262 ( \16639 , RIc2264d0_37);
not \U$16263 ( \16640 , \3810 );
or \U$16264 ( \16641 , \16639 , \16640 );
not \U$16265 ( \16642 , \2670 );
nand \U$16266 ( \16643 , \16642 , \5504 );
nand \U$16267 ( \16644 , \16641 , \16643 );
not \U$16268 ( \16645 , \16644 );
or \U$16269 ( \16646 , \16638 , \16645 );
nand \U$16270 ( \16647 , \15946 , \5519 );
nand \U$16271 ( \16648 , \16646 , \16647 );
not \U$16272 ( \16649 , \16648 );
not \U$16273 ( \16650 , \15911 );
not \U$16274 ( \16651 , \6307 );
or \U$16275 ( \16652 , \16650 , \16651 );
not \U$16276 ( \16653 , \13780 );
not \U$16277 ( \16654 , \16653 );
not \U$16278 ( \16655 , \9573 );
and \U$16279 ( \16656 , \16654 , \16655 );
and \U$16280 ( \16657 , \2479 , \8998 );
nor \U$16281 ( \16658 , \16656 , \16657 );
not \U$16282 ( \16659 , \16658 );
nand \U$16283 ( \16660 , \16659 , \6689 );
nand \U$16284 ( \16661 , \16652 , \16660 );
not \U$16285 ( \16662 , \16661 );
or \U$16286 ( \16663 , \16649 , \16662 );
or \U$16287 ( \16664 , \16661 , \16648 );
not \U$16288 ( \16665 , \9488 );
not \U$16289 ( \16666 , RIc225d50_53);
not \U$16290 ( \16667 , \1530 );
or \U$16291 ( \16668 , \16666 , \16667 );
nand \U$16292 ( \16669 , \3579 , \8772 );
nand \U$16293 ( \16670 , \16668 , \16669 );
not \U$16294 ( \16671 , \16670 );
or \U$16295 ( \16672 , \16665 , \16671 );
nand \U$16296 ( \16673 , \12945 , \15821 );
nand \U$16297 ( \16674 , \16672 , \16673 );
nand \U$16298 ( \16675 , \16664 , \16674 );
nand \U$16299 ( \16676 , \16663 , \16675 );
not \U$16300 ( \16677 , \16676 );
xor \U$16301 ( \16678 , \15679 , \15691 );
xor \U$16302 ( \16679 , \16678 , \15704 );
not \U$16303 ( \16680 , \16679 );
nand \U$16304 ( \16681 , \16677 , \16680 );
not \U$16305 ( \16682 , \16681 );
and \U$16306 ( \16683 , \15731 , \15742 );
not \U$16307 ( \16684 , \15731 );
and \U$16308 ( \16685 , \16684 , \15743 );
nor \U$16309 ( \16686 , \16683 , \16685 );
not \U$16310 ( \16687 , \15718 );
and \U$16311 ( \16688 , \16686 , \16687 );
not \U$16312 ( \16689 , \16686 );
and \U$16313 ( \16690 , \16689 , \15718 );
nor \U$16314 ( \16691 , \16688 , \16690 );
not \U$16315 ( \16692 , \16691 );
not \U$16316 ( \16693 , \16692 );
or \U$16317 ( \16694 , \16682 , \16693 );
nand \U$16318 ( \16695 , \16676 , \16679 );
nand \U$16319 ( \16696 , \16694 , \16695 );
not \U$16320 ( \16697 , \16696 );
or \U$16321 ( \16698 , \16637 , \16697 );
not \U$16322 ( \16699 , \16603 );
not \U$16323 ( \16700 , \16635 );
nand \U$16324 ( \16701 , \16699 , \16700 );
nand \U$16325 ( \16702 , \16698 , \16701 );
buf \U$16326 ( \16703 , \16702 );
not \U$16327 ( \16704 , \16703 );
nand \U$16328 ( \16705 , \16481 , \16704 );
not \U$16329 ( \16706 , \16705 );
or \U$16330 ( \16707 , \16353 , \16706 );
nand \U$16331 ( \16708 , \16480 , \16703 );
nand \U$16332 ( \16709 , \16707 , \16708 );
nand \U$16333 ( \16710 , \16227 , \16709 );
nand \U$16334 ( \16711 , \16226 , \16710 );
not \U$16335 ( \16712 , \16711 );
not \U$16336 ( \16713 , \16009 );
not \U$16337 ( \16714 , \16713 );
not \U$16338 ( \16715 , \15993 );
or \U$16339 ( \16716 , \16714 , \16715 );
nand \U$16340 ( \16717 , \16009 , \15992 );
nand \U$16341 ( \16718 , \16716 , \16717 );
and \U$16342 ( \16719 , \16718 , \16118 );
not \U$16343 ( \16720 , \16718 );
not \U$16344 ( \16721 , \16118 );
and \U$16345 ( \16722 , \16720 , \16721 );
nor \U$16346 ( \16723 , \16719 , \16722 );
not \U$16347 ( \16724 , \16723 );
nand \U$16348 ( \16725 , \16712 , \16724 );
not \U$16349 ( \16726 , \16725 );
xor \U$16350 ( \16727 , \16137 , \16181 );
xor \U$16351 ( \16728 , \16727 , \16135 );
not \U$16352 ( \16729 , \16728 );
or \U$16353 ( \16730 , \16726 , \16729 );
not \U$16354 ( \16731 , \16712 );
not \U$16355 ( \16732 , \16724 );
nand \U$16356 ( \16733 , \16731 , \16732 );
nand \U$16357 ( \16734 , \16730 , \16733 );
and \U$16358 ( \16735 , \16203 , \16734 );
and \U$16359 ( \16736 , \16200 , \16202 );
or \U$16360 ( \16737 , \16735 , \16736 );
not \U$16361 ( \16738 , \16737 );
nand \U$16362 ( \16739 , \16198 , \16738 );
buf \U$16363 ( \16740 , \16739 );
xor \U$16364 ( \16741 , \16200 , \16202 );
xor \U$16365 ( \16742 , \16741 , \16734 );
not \U$16366 ( \16743 , \16728 );
and \U$16367 ( \16744 , \16711 , \16723 );
not \U$16368 ( \16745 , \16711 );
and \U$16369 ( \16746 , \16745 , \16724 );
nor \U$16370 ( \16747 , \16744 , \16746 );
not \U$16371 ( \16748 , \16747 );
not \U$16372 ( \16749 , \16748 );
or \U$16373 ( \16750 , \16743 , \16749 );
not \U$16374 ( \16751 , \16728 );
nand \U$16375 ( \16752 , \16751 , \16747 );
nand \U$16376 ( \16753 , \16750 , \16752 );
xor \U$16377 ( \16754 , \15640 , \15651 );
xor \U$16378 ( \16755 , \16754 , \15662 );
not \U$16379 ( \16756 , \9398 );
not \U$16380 ( \16757 , \15850 );
or \U$16381 ( \16758 , \16756 , \16757 );
not \U$16382 ( \16759 , RIc226110_45);
not \U$16383 ( \16760 , \2234 );
or \U$16384 ( \16761 , \16759 , \16760 );
not \U$16385 ( \16762 , \11648 );
not \U$16386 ( \16763 , \16762 );
nand \U$16387 ( \16764 , \16763 , \10429 );
nand \U$16388 ( \16765 , \16761 , \16764 );
nand \U$16389 ( \16766 , \16765 , \9384 );
nand \U$16390 ( \16767 , \16758 , \16766 );
not \U$16391 ( \16768 , \16767 );
not \U$16392 ( \16769 , \11974 );
not \U$16393 ( \16770 , \15896 );
or \U$16394 ( \16771 , \16769 , \16770 );
not \U$16395 ( \16772 , RIc225b70_57);
not \U$16396 ( \16773 , \2118 );
or \U$16397 ( \16774 , \16772 , \16773 );
nand \U$16398 ( \16775 , \1020 , \15262 );
nand \U$16399 ( \16776 , \16774 , \16775 );
nand \U$16400 ( \16777 , \16776 , \11965 );
nand \U$16401 ( \16778 , \16771 , \16777 );
not \U$16402 ( \16779 , \16778 );
or \U$16403 ( \16780 , \16768 , \16779 );
or \U$16404 ( \16781 , \16767 , \16778 );
not \U$16405 ( \16782 , \11038 );
not \U$16406 ( \16783 , \15859 );
or \U$16407 ( \16784 , \16782 , \16783 );
not \U$16408 ( \16785 , RIc225c60_55);
not \U$16409 ( \16786 , \1440 );
or \U$16410 ( \16787 , \16785 , \16786 );
not \U$16411 ( \16788 , RIc225c60_55);
nand \U$16412 ( \16789 , \1371 , \16788 );
nand \U$16413 ( \16790 , \16787 , \16789 );
nand \U$16414 ( \16791 , \16790 , \11118 );
nand \U$16415 ( \16792 , \16784 , \16791 );
nand \U$16416 ( \16793 , \16781 , \16792 );
nand \U$16417 ( \16794 , \16780 , \16793 );
xor \U$16418 ( \16795 , \16755 , \16794 );
xor \U$16419 ( \16796 , \16039 , \16074 );
xor \U$16420 ( \16797 , \16796 , \16084 );
and \U$16421 ( \16798 , \16795 , \16797 );
and \U$16422 ( \16799 , \16755 , \16794 );
or \U$16423 ( \16800 , \16798 , \16799 );
xor \U$16424 ( \16801 , \15880 , \15916 );
xor \U$16425 ( \16802 , \16801 , \15919 );
xor \U$16426 ( \16803 , \16800 , \16802 );
and \U$16427 ( \16804 , \15789 , \15826 );
not \U$16428 ( \16805 , \15789 );
and \U$16429 ( \16806 , \16805 , \15827 );
or \U$16430 ( \16807 , \16804 , \16806 );
xor \U$16431 ( \16808 , \16807 , \15866 );
and \U$16432 ( \16809 , \16803 , \16808 );
and \U$16433 ( \16810 , \16800 , \16802 );
or \U$16434 ( \16811 , \16809 , \16810 );
not \U$16435 ( \16812 , \15985 );
not \U$16436 ( \16813 , \15978 );
or \U$16437 ( \16814 , \16812 , \16813 );
nand \U$16438 ( \16815 , \15984 , \15980 );
nand \U$16439 ( \16816 , \16814 , \16815 );
xor \U$16440 ( \16817 , \16816 , \15975 );
xor \U$16441 ( \16818 , \16811 , \16817 );
buf \U$16442 ( \16819 , \15875 );
xor \U$16443 ( \16820 , \15877 , \15922 );
xor \U$16444 ( \16821 , \16819 , \16820 );
and \U$16445 ( \16822 , \16818 , \16821 );
and \U$16446 ( \16823 , \16811 , \16817 );
or \U$16447 ( \16824 , \16822 , \16823 );
xor \U$16448 ( \16825 , \16109 , \16090 );
xnor \U$16449 ( \16826 , \16825 , \16112 );
not \U$16450 ( \16827 , \16826 );
not \U$16451 ( \16828 , \16169 );
not \U$16452 ( \16829 , \16153 );
or \U$16453 ( \16830 , \16828 , \16829 );
nand \U$16454 ( \16831 , \16168 , \16164 );
nand \U$16455 ( \16832 , \16830 , \16831 );
and \U$16456 ( \16833 , \16832 , \16142 );
not \U$16457 ( \16834 , \16832 );
not \U$16458 ( \16835 , \16142 );
and \U$16459 ( \16836 , \16834 , \16835 );
nor \U$16460 ( \16837 , \16833 , \16836 );
not \U$16461 ( \16838 , \16837 );
or \U$16462 ( \16839 , \16827 , \16838 );
or \U$16463 ( \16840 , \16837 , \16826 );
xor \U$16464 ( \16841 , \16087 , \16036 );
xor \U$16465 ( \16842 , \16841 , \16034 );
not \U$16466 ( \16843 , \16842 );
xor \U$16467 ( \16844 , \16102 , \16097 );
xnor \U$16468 ( \16845 , \16844 , \16099 );
not \U$16469 ( \16846 , \16845 );
not \U$16470 ( \16847 , \16846 );
or \U$16471 ( \16848 , \16843 , \16847 );
or \U$16472 ( \16849 , \16846 , \16842 );
and \U$16473 ( \16850 , \16699 , \16700 );
not \U$16474 ( \16851 , \16699 );
and \U$16475 ( \16852 , \16851 , \16635 );
nor \U$16476 ( \16853 , \16850 , \16852 );
xor \U$16477 ( \16854 , \16696 , \16853 );
nand \U$16478 ( \16855 , \16849 , \16854 );
nand \U$16479 ( \16856 , \16848 , \16855 );
nand \U$16480 ( \16857 , \16840 , \16856 );
nand \U$16481 ( \16858 , \16839 , \16857 );
xor \U$16482 ( \16859 , \16824 , \16858 );
xor \U$16483 ( \16860 , \16140 , \16171 );
xor \U$16484 ( \16861 , \16860 , \16178 );
and \U$16485 ( \16862 , \16859 , \16861 );
and \U$16486 ( \16863 , \16824 , \16858 );
or \U$16487 ( \16864 , \16862 , \16863 );
or \U$16488 ( \16865 , \16753 , \16864 );
xor \U$16489 ( \16866 , \16824 , \16858 );
xor \U$16490 ( \16867 , \16866 , \16861 );
not \U$16491 ( \16868 , \16867 );
xor \U$16492 ( \16869 , \16702 , \16479 );
not \U$16493 ( \16870 , \16352 );
and \U$16494 ( \16871 , \16869 , \16870 );
not \U$16495 ( \16872 , \16869 );
and \U$16496 ( \16873 , \16872 , \16352 );
nor \U$16497 ( \16874 , \16871 , \16873 );
not \U$16498 ( \16875 , \16874 );
not \U$16499 ( \16876 , \16875 );
xor \U$16500 ( \16877 , \16581 , \16593 );
xnor \U$16501 ( \16878 , \16877 , \16570 );
not \U$16502 ( \16879 , \16878 );
not \U$16503 ( \16880 , RIc2258a0_63);
not \U$16504 ( \16881 , \16880 );
not \U$16505 ( \16882 , RIc225828_64);
not \U$16506 ( \16883 , \16882 );
and \U$16507 ( \16884 , \16881 , \16883 );
and \U$16508 ( \16885 , \930 , \15620 );
not \U$16509 ( \16886 , \930 );
and \U$16510 ( \16887 , \16886 , RIc2258a0_63);
or \U$16511 ( \16888 , \16885 , \16887 );
nand \U$16512 ( \16889 , \16882 , RIc2258a0_63);
not \U$16513 ( \16890 , \16889 );
buf \U$16514 ( \16891 , \16890 );
and \U$16515 ( \16892 , \16888 , \16891 );
nor \U$16516 ( \16893 , \16884 , \16892 );
not \U$16517 ( \16894 , \2534 );
not \U$16518 ( \16895 , \16610 );
or \U$16519 ( \16896 , \16894 , \16895 );
not \U$16520 ( \16897 , RIc226d40_19);
not \U$16521 ( \16898 , \15684 );
or \U$16522 ( \16899 , \16897 , \16898 );
nand \U$16523 ( \16900 , \8806 , \3338 );
nand \U$16524 ( \16901 , \16899 , \16900 );
nand \U$16525 ( \16902 , \16901 , \2518 );
nand \U$16526 ( \16903 , \16896 , \16902 );
not \U$16527 ( \16904 , \16903 );
xor \U$16528 ( \16905 , \16893 , \16904 );
not \U$16529 ( \16906 , \2367 );
nor \U$16530 ( \16907 , \16906 , \16534 );
and \U$16531 ( \16908 , \8856 , \2370 );
not \U$16532 ( \16909 , \8856 );
and \U$16533 ( \16910 , \16909 , RIc226c50_21);
or \U$16534 ( \16911 , \16908 , \16910 );
and \U$16535 ( \16912 , \16911 , \2392 );
nor \U$16536 ( \16913 , \16907 , \16912 );
and \U$16537 ( \16914 , \16905 , \16913 );
and \U$16538 ( \16915 , \16893 , \16904 );
or \U$16539 ( \16916 , \16914 , \16915 );
not \U$16540 ( \16917 , \16916 );
or \U$16541 ( \16918 , \16879 , \16917 );
not \U$16542 ( \16919 , \898 );
not \U$16543 ( \16920 , \16261 );
or \U$16544 ( \16921 , \16919 , \16920 );
xor \U$16545 ( \16922 , RIc2275b0_1, \16248 );
nand \U$16546 ( \16923 , \16922 , \853 );
nand \U$16547 ( \16924 , \16921 , \16923 );
not \U$16548 ( \16925 , \16924 );
or \U$16549 ( \16926 , RIc227538_2, RIc2274c0_3);
nand \U$16550 ( \16927 , \16926 , \16248 );
and \U$16551 ( \16928 , RIc227538_2, RIc2274c0_3);
not \U$16552 ( \16929 , RIc2275b0_1);
nor \U$16553 ( \16930 , \16928 , \16929 );
nand \U$16554 ( \16931 , \16927 , \16930 );
nor \U$16555 ( \16932 , \16925 , \16931 );
not \U$16556 ( \16933 , \954 );
not \U$16557 ( \16934 , \16496 );
or \U$16558 ( \16935 , \16933 , \16934 );
and \U$16559 ( \16936 , \12755 , \946 );
not \U$16560 ( \16937 , \12755 );
and \U$16561 ( \16938 , \16937 , RIc2273d0_5);
or \U$16562 ( \16939 , \16936 , \16938 );
nand \U$16563 ( \16940 , \16939 , \950 );
nand \U$16564 ( \16941 , \16935 , \16940 );
xor \U$16565 ( \16942 , \16932 , \16941 );
not \U$16566 ( \16943 , \1120 );
not \U$16567 ( \16944 , RIc2272e0_7);
not \U$16568 ( \16945 , \10085 );
not \U$16569 ( \16946 , \16945 );
or \U$16570 ( \16947 , \16944 , \16946 );
nand \U$16571 ( \16948 , \10086 , \940 );
nand \U$16572 ( \16949 , \16947 , \16948 );
not \U$16573 ( \16950 , \16949 );
or \U$16574 ( \16951 , \16943 , \16950 );
not \U$16575 ( \16952 , RIc2272e0_7);
not \U$16576 ( \16953 , \10198 );
or \U$16577 ( \16954 , \16952 , \16953 );
nand \U$16578 ( \16955 , \10370 , \1139 );
nand \U$16579 ( \16956 , \16954 , \16955 );
nand \U$16580 ( \16957 , \16956 , \1118 );
nand \U$16581 ( \16958 , \16951 , \16957 );
and \U$16582 ( \16959 , \16942 , \16958 );
and \U$16583 ( \16960 , \16932 , \16941 );
or \U$16584 ( \16961 , \16959 , \16960 );
not \U$16585 ( \16962 , \2172 );
not \U$16586 ( \16963 , \16559 );
or \U$16587 ( \16964 , \16962 , \16963 );
not \U$16588 ( \16965 , RIc226a70_25);
not \U$16589 ( \16966 , \9775 );
or \U$16590 ( \16967 , \16965 , \16966 );
nand \U$16591 ( \16968 , \6492 , \3982 );
nand \U$16592 ( \16969 , \16967 , \16968 );
nand \U$16593 ( \16970 , \16969 , \2860 );
nand \U$16594 ( \16971 , \16964 , \16970 );
xor \U$16595 ( \16972 , \16961 , \16971 );
not \U$16596 ( \16973 , \1915 );
not \U$16597 ( \16974 , RIc226b60_23);
not \U$16598 ( \16975 , \10609 );
or \U$16599 ( \16976 , \16974 , \16975 );
nand \U$16600 ( \16977 , \10612 , \2111 );
nand \U$16601 ( \16978 , \16976 , \16977 );
not \U$16602 ( \16979 , \16978 );
or \U$16603 ( \16980 , \16973 , \16979 );
nand \U$16604 ( \16981 , \16545 , \1930 );
nand \U$16605 ( \16982 , \16980 , \16981 );
and \U$16606 ( \16983 , \16972 , \16982 );
and \U$16607 ( \16984 , \16961 , \16971 );
or \U$16608 ( \16985 , \16983 , \16984 );
nand \U$16609 ( \16986 , \16918 , \16985 );
not \U$16610 ( \16987 , \16878 );
not \U$16611 ( \16988 , \16916 );
nand \U$16612 ( \16989 , \16987 , \16988 );
nand \U$16613 ( \16990 , \16986 , \16989 );
xor \U$16614 ( \16991 , \16050 , \16060 );
xor \U$16615 ( \16992 , \16991 , \16071 );
not \U$16616 ( \16993 , \16992 );
and \U$16617 ( \16994 , \16588 , \1340 );
not \U$16618 ( \16995 , RIc2271f0_9);
not \U$16619 ( \16996 , \9297 );
or \U$16620 ( \16997 , \16995 , \16996 );
not \U$16621 ( \16998 , \10263 );
nand \U$16622 ( \16999 , \16998 , \1342 );
nand \U$16623 ( \17000 , \16997 , \16999 );
not \U$16624 ( \17001 , \17000 );
nor \U$16625 ( \17002 , \17001 , \1364 );
nor \U$16626 ( \17003 , \16994 , \17002 );
not \U$16627 ( \17004 , \17003 );
and \U$16628 ( \17005 , \16577 , \1120 );
and \U$16629 ( \17006 , \16949 , \1118 );
nor \U$16630 ( \17007 , \17005 , \17006 );
not \U$16631 ( \17008 , \17007 );
or \U$16632 ( \17009 , \17004 , \17008 );
not \U$16633 ( \17010 , \1310 );
not \U$16634 ( \17011 , \16067 );
or \U$16635 ( \17012 , \17010 , \17011 );
not \U$16636 ( \17013 , RIc227100_11);
not \U$16637 ( \17014 , \9250 );
not \U$16638 ( \17015 , \17014 );
not \U$16639 ( \17016 , \17015 );
or \U$16640 ( \17017 , \17013 , \17016 );
not \U$16641 ( \17018 , \11488 );
nand \U$16642 ( \17019 , \17018 , \1685 );
nand \U$16643 ( \17020 , \17017 , \17019 );
nand \U$16644 ( \17021 , \17020 , \9904 );
nand \U$16645 ( \17022 , \17012 , \17021 );
nand \U$16646 ( \17023 , \17009 , \17022 );
or \U$16647 ( \17024 , \17007 , \17003 );
nand \U$16648 ( \17025 , \17023 , \17024 );
not \U$16649 ( \17026 , \17025 );
nand \U$16650 ( \17027 , \16993 , \17026 );
not \U$16651 ( \17028 , \17027 );
not \U$16652 ( \17029 , \2154 );
not \U$16653 ( \17030 , \16512 );
or \U$16654 ( \17031 , \17029 , \17030 );
not \U$16655 ( \17032 , RIc226980_27);
not \U$16656 ( \17033 , \15603 );
or \U$16657 ( \17034 , \17032 , \17033 );
nand \U$16658 ( \17035 , \12791 , \2150 );
nand \U$16659 ( \17036 , \17034 , \17035 );
nand \U$16660 ( \17037 , \17036 , \2138 );
nand \U$16661 ( \17038 , \17031 , \17037 );
not \U$16662 ( \17039 , \17038 );
not \U$16663 ( \17040 , \9142 );
not \U$16664 ( \17041 , \16520 );
or \U$16665 ( \17042 , \17040 , \17041 );
and \U$16666 ( \17043 , RIc226890_29, \10220 );
not \U$16667 ( \17044 , RIc226890_29);
and \U$16668 ( \17045 , \17044 , \4407 );
or \U$16669 ( \17046 , \17043 , \17045 );
nand \U$16670 ( \17047 , \17046 , \2784 );
nand \U$16671 ( \17048 , \17042 , \17047 );
not \U$16672 ( \17049 , \17048 );
or \U$16673 ( \17050 , \17039 , \17049 );
or \U$16674 ( \17051 , \17048 , \17038 );
xor \U$16675 ( \17052 , \16483 , \16488 );
xor \U$16676 ( \17053 , \17052 , \16500 );
nand \U$16677 ( \17054 , \17051 , \17053 );
nand \U$16678 ( \17055 , \17050 , \17054 );
not \U$16679 ( \17056 , \17055 );
or \U$16680 ( \17057 , \17028 , \17056 );
nand \U$16681 ( \17058 , \17025 , \16992 );
nand \U$16682 ( \17059 , \17057 , \17058 );
xor \U$16683 ( \17060 , \16990 , \17059 );
not \U$16684 ( \17061 , \16438 );
not \U$16685 ( \17062 , \16432 );
and \U$16686 ( \17063 , \17061 , \17062 );
not \U$16687 ( \17064 , RIc225a80_59);
not \U$16688 ( \17065 , \17064 );
not \U$16689 ( \17066 , \3464 );
or \U$16690 ( \17067 , \17065 , \17066 );
not \U$16691 ( \17068 , \981 );
nand \U$16692 ( \17069 , \17068 , RIc225a80_59);
nand \U$16693 ( \17070 , \17067 , \17069 );
and \U$16694 ( \17071 , \17070 , \15164 );
nor \U$16695 ( \17072 , \17063 , \17071 );
not \U$16696 ( \17073 , \17072 );
not \U$16697 ( \17074 , \16446 );
not \U$16698 ( \17075 , \9129 );
not \U$16699 ( \17076 , \17075 );
and \U$16700 ( \17077 , \17074 , \17076 );
not \U$16701 ( \17078 , RIc226200_43);
not \U$16702 ( \17079 , \9584 );
or \U$16703 ( \17080 , \17078 , \17079 );
not \U$16704 ( \17081 , \2013 );
not \U$16705 ( \17082 , \17081 );
nand \U$16706 ( \17083 , \17082 , \9106 );
nand \U$16707 ( \17084 , \17080 , \17083 );
and \U$16708 ( \17085 , \17084 , \9110 );
nor \U$16709 ( \17086 , \17077 , \17085 );
not \U$16710 ( \17087 , \17086 );
or \U$16711 ( \17088 , \17073 , \17087 );
not \U$16712 ( \17089 , \11118 );
not \U$16713 ( \17090 , RIc225c60_55);
not \U$16714 ( \17091 , \3496 );
or \U$16715 ( \17092 , \17090 , \17091 );
nand \U$16716 ( \17093 , \5246 , \8767 );
nand \U$16717 ( \17094 , \17092 , \17093 );
not \U$16718 ( \17095 , \17094 );
or \U$16719 ( \17096 , \17089 , \17095 );
nand \U$16720 ( \17097 , \16790 , \11038 );
nand \U$16721 ( \17098 , \17096 , \17097 );
nand \U$16722 ( \17099 , \17088 , \17098 );
not \U$16723 ( \17100 , \17086 );
not \U$16724 ( \17101 , \17072 );
nand \U$16725 ( \17102 , \17100 , \17101 );
nand \U$16726 ( \17103 , \17099 , \17102 );
not \U$16727 ( \17104 , \17103 );
not \U$16728 ( \17105 , \16457 );
not \U$16729 ( \17106 , \9817 );
and \U$16730 ( \17107 , \17105 , \17106 );
not \U$16731 ( \17108 , RIc2262f0_41);
not \U$16732 ( \17109 , \15908 );
or \U$16733 ( \17110 , \17108 , \17109 );
nand \U$16734 ( \17111 , \9942 , \9822 );
nand \U$16735 ( \17112 , \17110 , \17111 );
and \U$16736 ( \17113 , \17112 , \9690 );
nor \U$16737 ( \17114 , \17107 , \17113 );
not \U$16738 ( \17115 , \17114 );
not \U$16739 ( \17116 , \16658 );
not \U$16740 ( \17117 , \6308 );
and \U$16741 ( \17118 , \17116 , \17117 );
not \U$16742 ( \17119 , \12990 );
not \U$16743 ( \17120 , \8998 );
and \U$16744 ( \17121 , \17119 , \17120 );
not \U$16745 ( \17122 , \11854 );
and \U$16746 ( \17123 , \17122 , \9573 );
nor \U$16747 ( \17124 , \17121 , \17123 );
not \U$16748 ( \17125 , \6689 );
nor \U$16749 ( \17126 , \17124 , \17125 );
nor \U$16750 ( \17127 , \17118 , \17126 );
not \U$16751 ( \17128 , \17127 );
or \U$16752 ( \17129 , \17115 , \17128 );
not \U$16753 ( \17130 , \9488 );
not \U$16754 ( \17131 , RIc225d50_53);
not \U$16755 ( \17132 , \1948 );
or \U$16756 ( \17133 , \17131 , \17132 );
nand \U$16757 ( \17134 , \3439 , \8782 );
nand \U$16758 ( \17135 , \17133 , \17134 );
not \U$16759 ( \17136 , \17135 );
or \U$16760 ( \17137 , \17130 , \17136 );
nand \U$16761 ( \17138 , \16670 , \11577 );
nand \U$16762 ( \17139 , \17137 , \17138 );
nand \U$16763 ( \17140 , \17129 , \17139 );
not \U$16764 ( \17141 , \17127 );
not \U$16765 ( \17142 , \17114 );
nand \U$16766 ( \17143 , \17141 , \17142 );
nand \U$16767 ( \17144 , \17140 , \17143 );
not \U$16768 ( \17145 , \17144 );
or \U$16769 ( \17146 , \17104 , \17145 );
or \U$16770 ( \17147 , \17144 , \17103 );
xor \U$16771 ( \17148 , \16604 , \16614 );
xor \U$16772 ( \17149 , \17148 , \16624 );
nand \U$16773 ( \17150 , \17147 , \17149 );
nand \U$16774 ( \17151 , \17146 , \17150 );
and \U$16775 ( \17152 , \17060 , \17151 );
and \U$16776 ( \17153 , \16990 , \17059 );
or \U$16777 ( \17154 , \17152 , \17153 );
not \U$16778 ( \17155 , \15267 );
not \U$16779 ( \17156 , \16776 );
or \U$16780 ( \17157 , \17155 , \17156 );
not \U$16781 ( \17158 , \14421 );
not \U$16782 ( \17159 , RIc225b70_57);
and \U$16783 ( \17160 , \17158 , \17159 );
not \U$16784 ( \17161 , \1169 );
and \U$16785 ( \17162 , \17161 , RIc225b70_57);
nor \U$16786 ( \17163 , \17160 , \17162 );
not \U$16787 ( \17164 , \17163 );
nand \U$16788 ( \17165 , \17164 , \11965 );
nand \U$16789 ( \17166 , \17157 , \17165 );
not \U$16790 ( \17167 , \10001 );
not \U$16791 ( \17168 , RIc226020_47);
not \U$16792 ( \17169 , \2833 );
or \U$16793 ( \17170 , \17168 , \17169 );
nand \U$16794 ( \17171 , \2443 , \9624 );
nand \U$16795 ( \17172 , \17170 , \17171 );
not \U$16796 ( \17173 , \17172 );
or \U$16797 ( \17174 , \17167 , \17173 );
nand \U$16798 ( \17175 , \16422 , \10953 );
nand \U$16799 ( \17176 , \17174 , \17175 );
xor \U$16800 ( \17177 , \17166 , \17176 );
not \U$16801 ( \17178 , \9934 );
not \U$16802 ( \17179 , RIc226110_45);
not \U$16803 ( \17180 , \4009 );
or \U$16804 ( \17181 , \17179 , \17180 );
not \U$16805 ( \17182 , \2258 );
nand \U$16806 ( \17183 , \17182 , \9100 );
nand \U$16807 ( \17184 , \17181 , \17183 );
not \U$16808 ( \17185 , \17184 );
or \U$16809 ( \17186 , \17178 , \17185 );
nand \U$16810 ( \17187 , \16765 , \15183 );
nand \U$16811 ( \17188 , \17186 , \17187 );
and \U$16812 ( \17189 , \17177 , \17188 );
and \U$16813 ( \17190 , \17166 , \17176 );
or \U$16814 ( \17191 , \17189 , \17190 );
not \U$16815 ( \17192 , \17191 );
not \U$16816 ( \17193 , \2358 );
not \U$16817 ( \17194 , \16373 );
or \U$16818 ( \17195 , \17193 , \17194 );
not \U$16819 ( \17196 , RIc226f20_15);
not \U$16820 ( \17197 , \9215 );
or \U$16821 ( \17198 , \17196 , \17197 );
nand \U$16822 ( \17199 , \8924 , \2301 );
nand \U$16823 ( \17200 , \17198 , \17199 );
nand \U$16824 ( \17201 , \17200 , \2320 );
nand \U$16825 ( \17202 , \17195 , \17201 );
not \U$16826 ( \17203 , \1963 );
not \U$16827 ( \17204 , \16620 );
or \U$16828 ( \17205 , \17203 , \17204 );
not \U$16829 ( \17206 , RIc226e30_17);
not \U$16830 ( \17207 , \8978 );
or \U$16831 ( \17208 , \17206 , \17207 );
nand \U$16832 ( \17209 , \8974 , \1960 );
nand \U$16833 ( \17210 , \17208 , \17209 );
nand \U$16834 ( \17211 , \17210 , \1945 );
nand \U$16835 ( \17212 , \17205 , \17211 );
xor \U$16836 ( \17213 , \17202 , \17212 );
not \U$16837 ( \17214 , \3629 );
not \U$16838 ( \17215 , RIc2266b0_33);
not \U$16839 ( \17216 , \15755 );
or \U$16840 ( \17217 , \17215 , \17216 );
nand \U$16841 ( \17218 , \3115 , \6355 );
nand \U$16842 ( \17219 , \17217 , \17218 );
not \U$16843 ( \17220 , \17219 );
or \U$16844 ( \17221 , \17214 , \17220 );
nand \U$16845 ( \17222 , \16364 , \3631 );
nand \U$16846 ( \17223 , \17221 , \17222 );
and \U$16847 ( \17224 , \17213 , \17223 );
and \U$16848 ( \17225 , \17202 , \17212 );
or \U$16849 ( \17226 , \17224 , \17225 );
not \U$16850 ( \17227 , \17226 );
nand \U$16851 ( \17228 , \17192 , \17227 );
not \U$16852 ( \17229 , \9459 );
not \U$16853 ( \17230 , RIc225e40_51);
not \U$16854 ( \17231 , \13235 );
or \U$16855 ( \17232 , \17230 , \17231 );
nand \U$16856 ( \17233 , \1729 , \12423 );
nand \U$16857 ( \17234 , \17232 , \17233 );
not \U$16858 ( \17235 , \17234 );
or \U$16859 ( \17236 , \17229 , \17235 );
nand \U$16860 ( \17237 , \16304 , \9445 );
nand \U$16861 ( \17238 , \17236 , \17237 );
not \U$16862 ( \17239 , \17238 );
not \U$16863 ( \17240 , \5519 );
not \U$16864 ( \17241 , \16644 );
or \U$16865 ( \17242 , \17240 , \17241 );
not \U$16866 ( \17243 , RIc2264d0_37);
not \U$16867 ( \17244 , \11841 );
or \U$16868 ( \17245 , \17243 , \17244 );
nand \U$16869 ( \17246 , \2064 , \5504 );
nand \U$16870 ( \17247 , \17245 , \17246 );
nand \U$16871 ( \17248 , \17247 , \5509 );
nand \U$16872 ( \17249 , \17242 , \17248 );
not \U$16873 ( \17250 , \17249 );
or \U$16874 ( \17251 , \17239 , \17250 );
or \U$16875 ( \17252 , \17249 , \17238 );
not \U$16876 ( \17253 , \4381 );
not \U$16877 ( \17254 , RIc2265c0_35);
not \U$16878 ( \17255 , \9804 );
or \U$16879 ( \17256 , \17254 , \17255 );
nand \U$16880 ( \17257 , \13251 , \3620 );
nand \U$16881 ( \17258 , \17256 , \17257 );
not \U$16882 ( \17259 , \17258 );
or \U$16883 ( \17260 , \17253 , \17259 );
nand \U$16884 ( \17261 , \16316 , \5135 );
nand \U$16885 ( \17262 , \17260 , \17261 );
nand \U$16886 ( \17263 , \17252 , \17262 );
nand \U$16887 ( \17264 , \17251 , \17263 );
and \U$16888 ( \17265 , \17228 , \17264 );
and \U$16889 ( \17266 , \17191 , \17226 );
nor \U$16890 ( \17267 , \17265 , \17266 );
not \U$16891 ( \17268 , \17267 );
not \U$16892 ( \17269 , \17268 );
xor \U$16893 ( \17270 , \16631 , \16629 );
and \U$16894 ( \17271 , \17270 , \16627 );
not \U$16895 ( \17272 , \17270 );
not \U$16896 ( \17273 , \16627 );
and \U$16897 ( \17274 , \17272 , \17273 );
nor \U$16898 ( \17275 , \17271 , \17274 );
not \U$16899 ( \17276 , \17275 );
or \U$16900 ( \17277 , \17269 , \17276 );
not \U$16901 ( \17278 , \17275 );
not \U$16902 ( \17279 , \17278 );
not \U$16903 ( \17280 , \17267 );
or \U$16904 ( \17281 , \17279 , \17280 );
not \U$16905 ( \17282 , \3653 );
not \U$16906 ( \17283 , \16410 );
or \U$16907 ( \17284 , \17282 , \17283 );
and \U$16908 ( \17285 , \9674 , RIc2267a0_31);
not \U$16909 ( \17286 , \9674 );
and \U$16910 ( \17287 , \17286 , \2072 );
or \U$16911 ( \17288 , \17285 , \17287 );
nand \U$16912 ( \17289 , \17288 , \2697 );
nand \U$16913 ( \17290 , \17284 , \17289 );
not \U$16914 ( \17291 , \17290 );
not \U$16915 ( \17292 , \15719 );
not \U$16916 ( \17293 , RIc225990_61);
not \U$16917 ( \17294 , \888 );
not \U$16918 ( \17295 , \17294 );
or \U$16919 ( \17296 , \17293 , \17295 );
nand \U$16920 ( \17297 , \888 , \12806 );
nand \U$16921 ( \17298 , \17296 , \17297 );
not \U$16922 ( \17299 , \17298 );
or \U$16923 ( \17300 , \17292 , \17299 );
nand \U$16924 ( \17301 , \16397 , \15729 );
nand \U$16925 ( \17302 , \17300 , \17301 );
not \U$16926 ( \17303 , \17302 );
or \U$16927 ( \17304 , \17291 , \17303 );
or \U$16928 ( \17305 , \17302 , \17290 );
not \U$16929 ( \17306 , \9534 );
and \U$16930 ( \17307 , RIc225f30_49, \3092 );
not \U$16931 ( \17308 , RIc225f30_49);
and \U$16932 ( \17309 , \17308 , \2305 );
or \U$16933 ( \17310 , \17307 , \17309 );
not \U$16934 ( \17311 , \17310 );
or \U$16935 ( \17312 , \17306 , \17311 );
nand \U$16936 ( \17313 , \16384 , \9552 );
nand \U$16937 ( \17314 , \17312 , \17313 );
nand \U$16938 ( \17315 , \17305 , \17314 );
nand \U$16939 ( \17316 , \17304 , \17315 );
not \U$16940 ( \17317 , \17316 );
xor \U$16941 ( \17318 , \16563 , \16549 );
xor \U$16942 ( \17319 , \17318 , \16537 );
not \U$16943 ( \17320 , \17319 );
or \U$16944 ( \17321 , \17317 , \17320 );
or \U$16945 ( \17322 , \17316 , \17319 );
xor \U$16946 ( \17323 , \16503 , \16514 );
xor \U$16947 ( \17324 , \17323 , \16522 );
nand \U$16948 ( \17325 , \17322 , \17324 );
nand \U$16949 ( \17326 , \17321 , \17325 );
nand \U$16950 ( \17327 , \17281 , \17326 );
nand \U$16951 ( \17328 , \17277 , \17327 );
xor \U$16952 ( \17329 , \17154 , \17328 );
xor \U$16953 ( \17330 , \16391 , \16429 );
xor \U$16954 ( \17331 , \17330 , \16466 );
not \U$16955 ( \17332 , \17331 );
not \U$16956 ( \17333 , \17332 );
not \U$16957 ( \17334 , \16680 );
not \U$16958 ( \17335 , \16692 );
or \U$16959 ( \17336 , \17334 , \17335 );
nand \U$16960 ( \17337 , \16691 , \16679 );
nand \U$16961 ( \17338 , \17336 , \17337 );
not \U$16962 ( \17339 , \16676 );
and \U$16963 ( \17340 , \17338 , \17339 );
not \U$16964 ( \17341 , \17338 );
and \U$16965 ( \17342 , \17341 , \16676 );
nor \U$16966 ( \17343 , \17340 , \17342 );
not \U$16967 ( \17344 , \17343 );
not \U$16968 ( \17345 , \17344 );
or \U$16969 ( \17346 , \17333 , \17345 );
not \U$16970 ( \17347 , \17331 );
not \U$16971 ( \17348 , \17343 );
or \U$16972 ( \17349 , \17347 , \17348 );
xor \U$16973 ( \17350 , \16598 , \16565 );
xor \U$16974 ( \17351 , \17350 , \16525 );
nand \U$16975 ( \17352 , \17349 , \17351 );
nand \U$16976 ( \17353 , \17346 , \17352 );
and \U$16977 ( \17354 , \17329 , \17353 );
and \U$16978 ( \17355 , \17154 , \17328 );
or \U$16979 ( \17356 , \17354 , \17355 );
not \U$16980 ( \17357 , \17356 );
not \U$16981 ( \17358 , \17357 );
not \U$16982 ( \17359 , \17358 );
or \U$16983 ( \17360 , \16876 , \17359 );
not \U$16984 ( \17361 , \17357 );
not \U$16985 ( \17362 , \16874 );
or \U$16986 ( \17363 , \17361 , \17362 );
and \U$16987 ( \17364 , \16473 , \16355 );
not \U$16988 ( \17365 , \16473 );
and \U$16989 ( \17366 , \17365 , \16477 );
nor \U$16990 ( \17367 , \17364 , \17366 );
buf \U$16991 ( \17368 , \16469 );
xor \U$16992 ( \17369 , \17367 , \17368 );
xor \U$16993 ( \17370 , \16755 , \16794 );
xor \U$16994 ( \17371 , \17370 , \16797 );
buf \U$16995 ( \17372 , \16366 );
xor \U$16996 ( \17373 , \16378 , \17372 );
xor \U$16997 ( \17374 , \17373 , \16388 );
not \U$16998 ( \17375 , \17374 );
not \U$16999 ( \17376 , \17375 );
xor \U$17000 ( \17377 , \16674 , \16661 );
xnor \U$17001 ( \17378 , \17377 , \16648 );
not \U$17002 ( \17379 , \17378 );
not \U$17003 ( \17380 , \17379 );
or \U$17004 ( \17381 , \17376 , \17380 );
not \U$17005 ( \17382 , \17378 );
not \U$17006 ( \17383 , \17374 );
or \U$17007 ( \17384 , \17382 , \17383 );
xor \U$17008 ( \17385 , \16296 , \16306 );
xor \U$17009 ( \17386 , \17385 , \16318 );
nand \U$17010 ( \17387 , \17384 , \17386 );
nand \U$17011 ( \17388 , \17381 , \17387 );
xor \U$17012 ( \17389 , \17371 , \17388 );
xor \U$17013 ( \17390 , \16441 , \16451 );
xor \U$17014 ( \17391 , \17390 , \16463 );
not \U$17015 ( \17392 , \17391 );
buf \U$17016 ( \17393 , \16767 );
xor \U$17017 ( \17394 , \16778 , \16792 );
xor \U$17018 ( \17395 , \17393 , \17394 );
buf \U$17019 ( \17396 , \17395 );
or \U$17020 ( \17397 , \17392 , \17396 );
xor \U$17021 ( \17398 , \16426 , \16401 );
xor \U$17022 ( \17399 , \17398 , \16412 );
buf \U$17023 ( \17400 , \17399 );
nand \U$17024 ( \17401 , \17397 , \17400 );
nand \U$17025 ( \17402 , \17396 , \17392 );
nand \U$17026 ( \17403 , \17401 , \17402 );
and \U$17027 ( \17404 , \17389 , \17403 );
and \U$17028 ( \17405 , \17371 , \17388 );
or \U$17029 ( \17406 , \17404 , \17405 );
xor \U$17030 ( \17407 , \17369 , \17406 );
not \U$17031 ( \17408 , \16347 );
not \U$17032 ( \17409 , \17408 );
not \U$17033 ( \17410 , \16349 );
or \U$17034 ( \17411 , \17409 , \17410 );
nand \U$17035 ( \17412 , \16343 , \16347 );
nand \U$17036 ( \17413 , \17411 , \17412 );
and \U$17037 ( \17414 , \17413 , \16350 );
not \U$17038 ( \17415 , \17413 );
not \U$17039 ( \17416 , \16350 );
and \U$17040 ( \17417 , \17415 , \17416 );
nor \U$17041 ( \17418 , \17414 , \17417 );
and \U$17042 ( \17419 , \17407 , \17418 );
and \U$17043 ( \17420 , \17369 , \17406 );
or \U$17044 ( \17421 , \17419 , \17420 );
nand \U$17045 ( \17422 , \17363 , \17421 );
nand \U$17046 ( \17423 , \17360 , \17422 );
not \U$17047 ( \17424 , \17423 );
not \U$17048 ( \17425 , \16215 );
not \U$17049 ( \17426 , \16709 );
not \U$17050 ( \17427 , \17426 );
or \U$17051 ( \17428 , \17425 , \17427 );
nand \U$17052 ( \17429 , \16214 , \16709 );
nand \U$17053 ( \17430 , \17428 , \17429 );
not \U$17054 ( \17431 , \16224 );
and \U$17055 ( \17432 , \17430 , \17431 );
not \U$17056 ( \17433 , \17430 );
and \U$17057 ( \17434 , \17433 , \16224 );
nor \U$17058 ( \17435 , \17432 , \17434 );
nand \U$17059 ( \17436 , \17424 , \17435 );
not \U$17060 ( \17437 , \17436 );
or \U$17061 ( \17438 , \16868 , \17437 );
not \U$17062 ( \17439 , \17435 );
nand \U$17063 ( \17440 , \17439 , \17423 );
nand \U$17064 ( \17441 , \17438 , \17440 );
nand \U$17065 ( \17442 , \16865 , \17441 );
nand \U$17066 ( \17443 , \16753 , \16864 );
nand \U$17067 ( \17444 , \17442 , \17443 );
or \U$17068 ( \17445 , \16742 , \17444 );
not \U$17069 ( \17446 , \15103 );
not \U$17070 ( \17447 , \15571 );
nand \U$17071 ( \17448 , \17446 , \17447 );
buf \U$17072 ( \17449 , \15568 );
and \U$17073 ( \17450 , \17448 , \17449 );
not \U$17074 ( \17451 , \15103 );
nor \U$17075 ( \17452 , \17451 , \17447 );
nor \U$17076 ( \17453 , \17450 , \17452 );
xor \U$17077 ( \17454 , \13553 , \13550 );
xnor \U$17078 ( \17455 , \17454 , \12924 );
nand \U$17079 ( \17456 , \17453 , \17455 );
nand \U$17080 ( \17457 , \16195 , \16740 , \17445 , \17456 );
nor \U$17081 ( \17458 , \15101 , \17457 );
not \U$17082 ( \17459 , \17458 );
xor \U$17083 ( \17460 , \16811 , \16817 );
xor \U$17084 ( \17461 , \17460 , \16821 );
xor \U$17085 ( \17462 , \16800 , \16802 );
xor \U$17086 ( \17463 , \17462 , \16808 );
buf \U$17087 ( \17464 , \17463 );
not \U$17088 ( \17465 , \17464 );
not \U$17089 ( \17466 , \16842 );
not \U$17090 ( \17467 , \17466 );
not \U$17091 ( \17468 , \16846 );
or \U$17092 ( \17469 , \17467 , \17468 );
nand \U$17093 ( \17470 , \16845 , \16842 );
nand \U$17094 ( \17471 , \17469 , \17470 );
and \U$17095 ( \17472 , \17471 , \16854 );
not \U$17096 ( \17473 , \17471 );
not \U$17097 ( \17474 , \16854 );
and \U$17098 ( \17475 , \17473 , \17474 );
nor \U$17099 ( \17476 , \17472 , \17475 );
not \U$17100 ( \17477 , \17476 );
or \U$17101 ( \17478 , \17465 , \17477 );
or \U$17102 ( \17479 , \17464 , \17476 );
not \U$17103 ( \17480 , \16337 );
not \U$17104 ( \17481 , \16340 );
or \U$17105 ( \17482 , \17480 , \17481 );
or \U$17106 ( \17483 , \16340 , \16337 );
nand \U$17107 ( \17484 , \17482 , \17483 );
not \U$17108 ( \17485 , \16327 );
and \U$17109 ( \17486 , \17484 , \17485 );
not \U$17110 ( \17487 , \17484 );
and \U$17111 ( \17488 , \17487 , \16327 );
nor \U$17112 ( \17489 , \17486 , \17488 );
not \U$17113 ( \17490 , \17489 );
xor \U$17114 ( \17491 , \16321 , \16229 );
xnor \U$17115 ( \17492 , \17491 , \16235 );
nand \U$17116 ( \17493 , \17490 , \17492 );
xor \U$17117 ( \17494 , \16246 , \16277 );
xor \U$17118 ( \17495 , \17494 , \16293 );
xor \U$17119 ( \17496 , \16249 , \16263 );
xor \U$17120 ( \17497 , \17496 , \16274 );
not \U$17121 ( \17498 , \1340 );
not \U$17122 ( \17499 , \17000 );
or \U$17123 ( \17500 , \17498 , \17499 );
and \U$17124 ( \17501 , RIc2271f0_9, \9324 );
not \U$17125 ( \17502 , RIc2271f0_9);
and \U$17126 ( \17503 , \17502 , \12100 );
nor \U$17127 ( \17504 , \17501 , \17503 );
nand \U$17128 ( \17505 , \17504 , \1363 );
nand \U$17129 ( \17506 , \17500 , \17505 );
xor \U$17130 ( \17507 , \17497 , \17506 );
not \U$17131 ( \17508 , \1311 );
not \U$17132 ( \17509 , \17020 );
or \U$17133 ( \17510 , \17508 , \17509 );
and \U$17134 ( \17511 , RIc227100_11, \10976 );
not \U$17135 ( \17512 , RIc227100_11);
and \U$17136 ( \17513 , \17512 , \13453 );
nor \U$17137 ( \17514 , \17511 , \17513 );
nand \U$17138 ( \17515 , \17514 , \1306 );
nand \U$17139 ( \17516 , \17510 , \17515 );
and \U$17140 ( \17517 , \17507 , \17516 );
and \U$17141 ( \17518 , \17497 , \17506 );
or \U$17142 ( \17519 , \17517 , \17518 );
xor \U$17143 ( \17520 , \17495 , \17519 );
not \U$17144 ( \17521 , \1682 );
not \U$17145 ( \17522 , \16291 );
or \U$17146 ( \17523 , \17521 , \17522 );
not \U$17147 ( \17524 , RIc227010_13);
not \U$17148 ( \17525 , \13223 );
or \U$17149 ( \17526 , \17524 , \17525 );
nand \U$17150 ( \17527 , \10110 , \1758 );
nand \U$17151 ( \17528 , \17526 , \17527 );
nand \U$17152 ( \17529 , \17528 , \1678 );
nand \U$17153 ( \17530 , \17523 , \17529 );
not \U$17154 ( \17531 , \17530 );
not \U$17155 ( \17532 , \2358 );
not \U$17156 ( \17533 , \17200 );
or \U$17157 ( \17534 , \17532 , \17533 );
not \U$17158 ( \17535 , RIc226f20_15);
not \U$17159 ( \17536 , \9046 );
or \U$17160 ( \17537 , \17535 , \17536 );
nand \U$17161 ( \17538 , \10644 , \1674 );
nand \U$17162 ( \17539 , \17537 , \17538 );
nand \U$17163 ( \17540 , \17539 , \2320 );
nand \U$17164 ( \17541 , \17534 , \17540 );
not \U$17165 ( \17542 , \17541 );
or \U$17166 ( \17543 , \17531 , \17542 );
or \U$17167 ( \17544 , \17541 , \17530 );
not \U$17168 ( \17545 , \2154 );
not \U$17169 ( \17546 , \17036 );
or \U$17170 ( \17547 , \17545 , \17546 );
not \U$17171 ( \17548 , RIc226980_27);
buf \U$17172 ( \17549 , \13687 );
not \U$17173 ( \17550 , \17549 );
or \U$17174 ( \17551 , \17548 , \17550 );
nand \U$17175 ( \17552 , \9875 , \2799 );
nand \U$17176 ( \17553 , \17551 , \17552 );
nand \U$17177 ( \17554 , \17553 , \2138 );
nand \U$17178 ( \17555 , \17547 , \17554 );
nand \U$17179 ( \17556 , \17544 , \17555 );
nand \U$17180 ( \17557 , \17543 , \17556 );
and \U$17181 ( \17558 , \17520 , \17557 );
and \U$17182 ( \17559 , \17495 , \17519 );
or \U$17183 ( \17560 , \17558 , \17559 );
xor \U$17184 ( \17561 , \17026 , \16992 );
xnor \U$17185 ( \17562 , \17561 , \17055 );
xor \U$17186 ( \17563 , \17560 , \17562 );
xor \U$17187 ( \17564 , \17003 , \17007 );
xor \U$17188 ( \17565 , \17564 , \17022 );
not \U$17189 ( \17566 , \2367 );
not \U$17190 ( \17567 , \16911 );
or \U$17191 ( \17568 , \17566 , \17567 );
not \U$17192 ( \17569 , RIc226c50_21);
not \U$17193 ( \17570 , \8830 );
or \U$17194 ( \17571 , \17569 , \17570 );
nand \U$17195 ( \17572 , \10289 , \2370 );
nand \U$17196 ( \17573 , \17571 , \17572 );
nand \U$17197 ( \17574 , \17573 , \2392 );
nand \U$17198 ( \17575 , \17568 , \17574 );
not \U$17199 ( \17576 , \17575 );
not \U$17200 ( \17577 , \1915 );
not \U$17201 ( \17578 , RIc226b60_23);
not \U$17202 ( \17579 , \8885 );
not \U$17203 ( \17580 , \17579 );
or \U$17204 ( \17581 , \17578 , \17580 );
not \U$17205 ( \17582 , \17579 );
nand \U$17206 ( \17583 , \17582 , \10210 );
nand \U$17207 ( \17584 , \17581 , \17583 );
not \U$17208 ( \17585 , \17584 );
or \U$17209 ( \17586 , \17577 , \17585 );
nand \U$17210 ( \17587 , \16978 , \1930 );
nand \U$17211 ( \17588 , \17586 , \17587 );
not \U$17212 ( \17589 , \17588 );
or \U$17213 ( \17590 , \17576 , \17589 );
or \U$17214 ( \17591 , \17588 , \17575 );
not \U$17215 ( \17592 , \2534 );
not \U$17216 ( \17593 , \16901 );
or \U$17217 ( \17594 , \17592 , \17593 );
and \U$17218 ( \17595 , RIc226d40_19, \9915 );
not \U$17219 ( \17596 , RIc226d40_19);
and \U$17220 ( \17597 , \17596 , \8951 );
or \U$17221 ( \17598 , \17595 , \17597 );
nand \U$17222 ( \17599 , \17598 , \2518 );
nand \U$17223 ( \17600 , \17594 , \17599 );
nand \U$17224 ( \17601 , \17591 , \17600 );
nand \U$17225 ( \17602 , \17590 , \17601 );
xor \U$17226 ( \17603 , \17565 , \17602 );
not \U$17227 ( \17604 , \16931 );
not \U$17228 ( \17605 , \16924 );
or \U$17229 ( \17606 , \17604 , \17605 );
or \U$17230 ( \17607 , \16924 , \16931 );
nand \U$17231 ( \17608 , \17606 , \17607 );
not \U$17232 ( \17609 , \1081 );
not \U$17233 ( \17610 , \16270 );
or \U$17234 ( \17611 , \17609 , \17610 );
not \U$17235 ( \17612 , RIc2274c0_3);
not \U$17236 ( \17613 , \13487 );
not \U$17237 ( \17614 , \17613 );
or \U$17238 ( \17615 , \17612 , \17614 );
nand \U$17239 ( \17616 , \13487 , \1032 );
nand \U$17240 ( \17617 , \17615 , \17616 );
nand \U$17241 ( \17618 , \17617 , \1040 );
nand \U$17242 ( \17619 , \17611 , \17618 );
xor \U$17243 ( \17620 , \17608 , \17619 );
not \U$17244 ( \17621 , \1120 );
not \U$17245 ( \17622 , \16956 );
or \U$17246 ( \17623 , \17621 , \17622 );
not \U$17247 ( \17624 , RIc2272e0_7);
not \U$17248 ( \17625 , \13497 );
not \U$17249 ( \17626 , \17625 );
or \U$17250 ( \17627 , \17624 , \17626 );
nand \U$17251 ( \17628 , \10356 , \1139 );
nand \U$17252 ( \17629 , \17627 , \17628 );
nand \U$17253 ( \17630 , \17629 , \1118 );
nand \U$17254 ( \17631 , \17623 , \17630 );
and \U$17255 ( \17632 , \17620 , \17631 );
and \U$17256 ( \17633 , \17608 , \17619 );
or \U$17257 ( \17634 , \17632 , \17633 );
not \U$17258 ( \17635 , \2086 );
not \U$17259 ( \17636 , \17046 );
or \U$17260 ( \17637 , \17635 , \17636 );
and \U$17261 ( \17638 , RIc226890_29, \5216 );
not \U$17262 ( \17639 , RIc226890_29);
and \U$17263 ( \17640 , \17639 , \13515 );
or \U$17264 ( \17641 , \17638 , \17640 );
nand \U$17265 ( \17642 , \17641 , \2784 );
nand \U$17266 ( \17643 , \17637 , \17642 );
xor \U$17267 ( \17644 , \17634 , \17643 );
not \U$17268 ( \17645 , \2860 );
not \U$17269 ( \17646 , RIc226a70_25);
not \U$17270 ( \17647 , \6719 );
or \U$17271 ( \17648 , \17646 , \17647 );
nand \U$17272 ( \17649 , \16543 , \1905 );
nand \U$17273 ( \17650 , \17648 , \17649 );
not \U$17274 ( \17651 , \17650 );
or \U$17275 ( \17652 , \17645 , \17651 );
nand \U$17276 ( \17653 , \16969 , \2173 );
nand \U$17277 ( \17654 , \17652 , \17653 );
and \U$17278 ( \17655 , \17644 , \17654 );
and \U$17279 ( \17656 , \17634 , \17643 );
or \U$17280 ( \17657 , \17655 , \17656 );
and \U$17281 ( \17658 , \17603 , \17657 );
and \U$17282 ( \17659 , \17565 , \17602 );
or \U$17283 ( \17660 , \17658 , \17659 );
and \U$17284 ( \17661 , \17563 , \17660 );
and \U$17285 ( \17662 , \17560 , \17562 );
or \U$17286 ( \17663 , \17661 , \17662 );
and \U$17287 ( \17664 , \17493 , \17663 );
nor \U$17288 ( \17665 , \17490 , \17492 );
nor \U$17289 ( \17666 , \17664 , \17665 );
not \U$17290 ( \17667 , \17666 );
nand \U$17291 ( \17668 , \17479 , \17667 );
nand \U$17292 ( \17669 , \17478 , \17668 );
xor \U$17293 ( \17670 , \17461 , \17669 );
xor \U$17294 ( \17671 , \16856 , \16826 );
and \U$17295 ( \17672 , \17671 , \16837 );
not \U$17296 ( \17673 , \17671 );
not \U$17297 ( \17674 , \16837 );
and \U$17298 ( \17675 , \17673 , \17674 );
nor \U$17299 ( \17676 , \17672 , \17675 );
xnor \U$17300 ( \17677 , \17670 , \17676 );
xor \U$17301 ( \17678 , \17560 , \17562 );
xor \U$17302 ( \17679 , \17678 , \17660 );
xor \U$17303 ( \17680 , \17497 , \17506 );
xor \U$17304 ( \17681 , \17680 , \17516 );
not \U$17305 ( \17682 , \17681 );
xor \U$17306 ( \17683 , \17530 , \17541 );
xnor \U$17307 ( \17684 , \17683 , \17555 );
nand \U$17308 ( \17685 , \17682 , \17684 );
not \U$17309 ( \17686 , \17685 );
not \U$17310 ( \17687 , \15267 );
not \U$17311 ( \17688 , RIc225b70_57);
not \U$17312 ( \17689 , \1222 );
or \U$17313 ( \17690 , \17688 , \17689 );
nand \U$17314 ( \17691 , \1439 , \11033 );
nand \U$17315 ( \17692 , \17690 , \17691 );
not \U$17316 ( \17693 , \17692 );
or \U$17317 ( \17694 , \17687 , \17693 );
and \U$17318 ( \17695 , RIc225b70_57, \5246 );
not \U$17319 ( \17696 , RIc225b70_57);
and \U$17320 ( \17697 , \17696 , \2380 );
nor \U$17321 ( \17698 , \17695 , \17697 );
nand \U$17322 ( \17699 , \17698 , \11965 );
nand \U$17323 ( \17700 , \17694 , \17699 );
not \U$17324 ( \17701 , \17700 );
not \U$17325 ( \17702 , RIc2266b0_33);
not \U$17326 ( \17703 , \3725 );
not \U$17327 ( \17704 , \17703 );
or \U$17328 ( \17705 , \17702 , \17704 );
nand \U$17329 ( \17706 , \2980 , \16360 );
nand \U$17330 ( \17707 , \17705 , \17706 );
and \U$17331 ( \17708 , \17707 , \3631 );
and \U$17332 ( \17709 , \3640 , \12551 );
not \U$17333 ( \17710 , \3640 );
and \U$17334 ( \17711 , \17710 , RIc2266b0_33);
or \U$17335 ( \17712 , \17709 , \17711 );
and \U$17336 ( \17713 , \17712 , \3629 );
nor \U$17337 ( \17714 , \17708 , \17713 );
or \U$17338 ( \17715 , \17701 , \17714 );
not \U$17339 ( \17716 , \17714 );
not \U$17340 ( \17717 , \17701 );
or \U$17341 ( \17718 , \17716 , \17717 );
xor \U$17342 ( \17719 , \17608 , \17619 );
xor \U$17343 ( \17720 , \17719 , \17631 );
nand \U$17344 ( \17721 , \17718 , \17720 );
nand \U$17345 ( \17722 , \17715 , \17721 );
not \U$17346 ( \17723 , \17722 );
or \U$17347 ( \17724 , \17686 , \17723 );
not \U$17348 ( \17725 , \17684 );
nand \U$17349 ( \17726 , \17725 , \17681 );
nand \U$17350 ( \17727 , \17724 , \17726 );
not \U$17351 ( \17728 , \17727 );
xor \U$17352 ( \17729 , \17565 , \17602 );
xor \U$17353 ( \17730 , \17729 , \17657 );
not \U$17354 ( \17731 , \17730 );
or \U$17355 ( \17732 , \17728 , \17731 );
not \U$17356 ( \17733 , \17727 );
not \U$17357 ( \17734 , \17733 );
not \U$17358 ( \17735 , \17730 );
not \U$17359 ( \17736 , \17735 );
or \U$17360 ( \17737 , \17734 , \17736 );
not \U$17361 ( \17738 , \1963 );
not \U$17362 ( \17739 , \17210 );
or \U$17363 ( \17740 , \17738 , \17739 );
not \U$17364 ( \17741 , \1952 );
not \U$17365 ( \17742 , \14968 );
or \U$17366 ( \17743 , \17741 , \17742 );
not \U$17367 ( \17744 , \8910 );
or \U$17368 ( \17745 , \17744 , \1952 );
nand \U$17369 ( \17746 , \17743 , \17745 );
nand \U$17370 ( \17747 , \17746 , \1945 );
nand \U$17371 ( \17748 , \17740 , \17747 );
and \U$17372 ( \17749 , \2072 , \5569 );
not \U$17373 ( \17750 , \2072 );
and \U$17374 ( \17751 , \17750 , \13525 );
nor \U$17375 ( \17752 , \17749 , \17751 );
not \U$17376 ( \17753 , \17752 );
not \U$17377 ( \17754 , \11182 );
and \U$17378 ( \17755 , \17753 , \17754 );
and \U$17379 ( \17756 , \17288 , \2710 );
nor \U$17380 ( \17757 , \17755 , \17756 );
not \U$17381 ( \17758 , \17757 );
xor \U$17382 ( \17759 , \17748 , \17758 );
not \U$17383 ( \17760 , \3629 );
not \U$17384 ( \17761 , \17707 );
or \U$17385 ( \17762 , \17760 , \17761 );
nand \U$17386 ( \17763 , \17219 , \3631 );
nand \U$17387 ( \17764 , \17762 , \17763 );
xnor \U$17388 ( \17765 , \17759 , \17764 );
xor \U$17389 ( \17766 , \17600 , \17575 );
xnor \U$17390 ( \17767 , \17766 , \17588 );
nand \U$17391 ( \17768 , \17765 , \17767 );
xor \U$17392 ( \17769 , \17634 , \17643 );
xor \U$17393 ( \17770 , \17769 , \17654 );
and \U$17394 ( \17771 , \17768 , \17770 );
nor \U$17395 ( \17772 , \17765 , \17767 );
nor \U$17396 ( \17773 , \17771 , \17772 );
not \U$17397 ( \17774 , \17773 );
nand \U$17398 ( \17775 , \17737 , \17774 );
nand \U$17399 ( \17776 , \17732 , \17775 );
xor \U$17400 ( \17777 , \17679 , \17776 );
xor \U$17401 ( \17778 , \17202 , \17212 );
xor \U$17402 ( \17779 , \17778 , \17223 );
not \U$17403 ( \17780 , \5519 );
not \U$17404 ( \17781 , \17247 );
or \U$17405 ( \17782 , \17780 , \17781 );
not \U$17406 ( \17783 , RIc2264d0_37);
not \U$17407 ( \17784 , \11068 );
or \U$17408 ( \17785 , \17783 , \17784 );
nand \U$17409 ( \17786 , \2730 , \5504 );
nand \U$17410 ( \17787 , \17785 , \17786 );
nand \U$17411 ( \17788 , \17787 , \5509 );
nand \U$17412 ( \17789 , \17782 , \17788 );
not \U$17413 ( \17790 , \9459 );
not \U$17414 ( \17791 , RIc225e40_51);
not \U$17415 ( \17792 , \2345 );
or \U$17416 ( \17793 , \17791 , \17792 );
nand \U$17417 ( \17794 , \2353 , \11795 );
nand \U$17418 ( \17795 , \17793 , \17794 );
not \U$17419 ( \17796 , \17795 );
or \U$17420 ( \17797 , \17790 , \17796 );
nand \U$17421 ( \17798 , \17234 , \11708 );
nand \U$17422 ( \17799 , \17797 , \17798 );
or \U$17423 ( \17800 , \17789 , \17799 );
not \U$17424 ( \17801 , \4381 );
not \U$17425 ( \17802 , RIc2265c0_35);
not \U$17426 ( \17803 , \10532 );
or \U$17427 ( \17804 , \17802 , \17803 );
nand \U$17428 ( \17805 , \4500 , \9587 );
nand \U$17429 ( \17806 , \17804 , \17805 );
not \U$17430 ( \17807 , \17806 );
or \U$17431 ( \17808 , \17801 , \17807 );
nand \U$17432 ( \17809 , \17258 , \4383 );
nand \U$17433 ( \17810 , \17808 , \17809 );
nand \U$17434 ( \17811 , \17800 , \17810 );
nand \U$17435 ( \17812 , \17789 , \17799 );
nand \U$17436 ( \17813 , \17811 , \17812 );
xor \U$17437 ( \17814 , \17779 , \17813 );
not \U$17438 ( \17815 , \9690 );
not \U$17439 ( \17816 , RIc2262f0_41);
not \U$17440 ( \17817 , \5819 );
or \U$17441 ( \17818 , \17816 , \17817 );
not \U$17442 ( \17819 , \15382 );
not \U$17443 ( \17820 , RIc2262f0_41);
nand \U$17444 ( \17821 , \17819 , \17820 );
nand \U$17445 ( \17822 , \17818 , \17821 );
not \U$17446 ( \17823 , \17822 );
or \U$17447 ( \17824 , \17815 , \17823 );
nand \U$17448 ( \17825 , \17112 , \9816 );
nand \U$17449 ( \17826 , \17824 , \17825 );
not \U$17450 ( \17827 , \6689 );
not \U$17451 ( \17828 , RIc2263e0_39);
not \U$17452 ( \17829 , \2670 );
or \U$17453 ( \17830 , \17828 , \17829 );
buf \U$17454 ( \17831 , \2720 );
nand \U$17455 ( \17832 , \17831 , \5498 );
nand \U$17456 ( \17833 , \17830 , \17832 );
not \U$17457 ( \17834 , \17833 );
or \U$17458 ( \17835 , \17827 , \17834 );
not \U$17459 ( \17836 , \17124 );
nand \U$17460 ( \17837 , \17836 , \6307 );
nand \U$17461 ( \17838 , \17835 , \17837 );
nor \U$17462 ( \17839 , \17826 , \17838 );
not \U$17463 ( \17840 , \9488 );
not \U$17464 ( \17841 , RIc225d50_53);
not \U$17465 ( \17842 , \3783 );
or \U$17466 ( \17843 , \17841 , \17842 );
nand \U$17467 ( \17844 , \1486 , \8782 );
nand \U$17468 ( \17845 , \17843 , \17844 );
not \U$17469 ( \17846 , \17845 );
or \U$17470 ( \17847 , \17840 , \17846 );
nand \U$17471 ( \17848 , \17135 , \12945 );
nand \U$17472 ( \17849 , \17847 , \17848 );
not \U$17473 ( \17850 , \17849 );
or \U$17474 ( \17851 , \17839 , \17850 );
nand \U$17475 ( \17852 , \17826 , \17838 );
nand \U$17476 ( \17853 , \17851 , \17852 );
xor \U$17477 ( \17854 , \17814 , \17853 );
not \U$17478 ( \17855 , \17854 );
not \U$17479 ( \17856 , \11324 );
not \U$17480 ( \17857 , \3620 );
and \U$17481 ( \17858 , \17856 , \17857 );
and \U$17482 ( \17859 , \11320 , \3620 );
nor \U$17483 ( \17860 , \17858 , \17859 );
not \U$17484 ( \17861 , \17860 );
not \U$17485 ( \17862 , \13910 );
and \U$17486 ( \17863 , \17861 , \17862 );
and \U$17487 ( \17864 , \17806 , \4383 );
nor \U$17488 ( \17865 , \17863 , \17864 );
not \U$17489 ( \17866 , \888 );
xor \U$17490 ( \17867 , RIc2258a0_63, \17866 );
not \U$17491 ( \17868 , \17867 );
not \U$17492 ( \17869 , \16891 );
not \U$17493 ( \17870 , \17869 );
and \U$17494 ( \17871 , \17868 , \17870 );
not \U$17495 ( \17872 , RIc2258a0_63);
not \U$17496 ( \17873 , \12472 );
or \U$17497 ( \17874 , \17872 , \17873 );
nand \U$17498 ( \17875 , \1072 , \16880 );
nand \U$17499 ( \17876 , \17874 , \17875 );
and \U$17500 ( \17877 , \17876 , RIc225828_64);
nor \U$17501 ( \17878 , \17871 , \17877 );
nand \U$17502 ( \17879 , \17865 , \17878 );
not \U$17503 ( \17880 , \9552 );
not \U$17504 ( \17881 , RIc225f30_49);
not \U$17505 ( \17882 , \13914 );
or \U$17506 ( \17883 , \17881 , \17882 );
nand \U$17507 ( \17884 , \2421 , \9541 );
nand \U$17508 ( \17885 , \17883 , \17884 );
not \U$17509 ( \17886 , \17885 );
or \U$17510 ( \17887 , \17880 , \17886 );
not \U$17511 ( \17888 , RIc225f30_49);
not \U$17512 ( \17889 , \9570 );
or \U$17513 ( \17890 , \17888 , \17889 );
nand \U$17514 ( \17891 , \2443 , \9541 );
nand \U$17515 ( \17892 , \17890 , \17891 );
nand \U$17516 ( \17893 , \17892 , \10445 );
nand \U$17517 ( \17894 , \17887 , \17893 );
and \U$17518 ( \17895 , \17879 , \17894 );
nor \U$17519 ( \17896 , \17865 , \17878 );
nor \U$17520 ( \17897 , \17895 , \17896 );
not \U$17521 ( \17898 , \17897 );
not \U$17522 ( \17899 , \9129 );
and \U$17523 ( \17900 , \2591 , RIc226200_43);
not \U$17524 ( \17901 , \2591 );
and \U$17525 ( \17902 , \17901 , \9125 );
or \U$17526 ( \17903 , \17900 , \17902 );
not \U$17527 ( \17904 , \17903 );
or \U$17528 ( \17905 , \17899 , \17904 );
not \U$17529 ( \17906 , RIc226200_43);
not \U$17530 ( \17907 , \2554 );
or \U$17531 ( \17908 , \17906 , \17907 );
nand \U$17532 ( \17909 , \3446 , \9106 );
nand \U$17533 ( \17910 , \17908 , \17909 );
nand \U$17534 ( \17911 , \17910 , \9110 );
nand \U$17535 ( \17912 , \17905 , \17911 );
not \U$17536 ( \17913 , \12670 );
and \U$17537 ( \17914 , RIc225a80_59, \1021 );
not \U$17538 ( \17915 , RIc225a80_59);
and \U$17539 ( \17916 , \17915 , \2119 );
or \U$17540 ( \17917 , \17914 , \17916 );
not \U$17541 ( \17918 , \17917 );
or \U$17542 ( \17919 , \17913 , \17918 );
and \U$17543 ( \17920 , RIc225a80_59, \1170 );
not \U$17544 ( \17921 , RIc225a80_59);
and \U$17545 ( \17922 , \17921 , \1169 );
or \U$17546 ( \17923 , \17920 , \17922 );
nand \U$17547 ( \17924 , \17923 , \15164 );
nand \U$17548 ( \17925 , \17919 , \17924 );
or \U$17549 ( \17926 , \17912 , \17925 );
not \U$17550 ( \17927 , \12532 );
not \U$17551 ( \17928 , RIc225c60_55);
not \U$17552 ( \17929 , \1529 );
not \U$17553 ( \17930 , \17929 );
or \U$17554 ( \17931 , \17928 , \17930 );
nand \U$17555 ( \17932 , \3579 , \8767 );
nand \U$17556 ( \17933 , \17931 , \17932 );
not \U$17557 ( \17934 , \17933 );
or \U$17558 ( \17935 , \17927 , \17934 );
not \U$17559 ( \17936 , RIc225c60_55);
not \U$17560 ( \17937 , \10909 );
or \U$17561 ( \17938 , \17936 , \17937 );
not \U$17562 ( \17939 , RIc225c60_55);
nand \U$17563 ( \17940 , \17939 , \1330 );
nand \U$17564 ( \17941 , \17938 , \17940 );
nand \U$17565 ( \17942 , \17941 , \11118 );
nand \U$17566 ( \17943 , \17935 , \17942 );
and \U$17567 ( \17944 , \17926 , \17943 );
and \U$17568 ( \17945 , \17912 , \17925 );
nor \U$17569 ( \17946 , \17944 , \17945 );
not \U$17570 ( \17947 , \17946 );
or \U$17571 ( \17948 , \17898 , \17947 );
not \U$17572 ( \17949 , \9705 );
not \U$17573 ( \17950 , \17822 );
or \U$17574 ( \17951 , \17949 , \17950 );
not \U$17575 ( \17952 , RIc2262f0_41);
not \U$17576 ( \17953 , \2894 );
or \U$17577 ( \17954 , \17952 , \17953 );
nand \U$17578 ( \17955 , \2498 , \12937 );
nand \U$17579 ( \17956 , \17954 , \17955 );
nand \U$17580 ( \17957 , \17956 , \9690 );
nand \U$17581 ( \17958 , \17951 , \17957 );
not \U$17582 ( \17959 , \17958 );
not \U$17583 ( \17960 , \6307 );
not \U$17584 ( \17961 , \17833 );
or \U$17585 ( \17962 , \17960 , \17961 );
not \U$17586 ( \17963 , RIc2263e0_39);
not \U$17587 ( \17964 , \11841 );
or \U$17588 ( \17965 , \17963 , \17964 );
not \U$17589 ( \17966 , \11841 );
nand \U$17590 ( \17967 , \17966 , \8990 );
nand \U$17591 ( \17968 , \17965 , \17967 );
nand \U$17592 ( \17969 , \17968 , \6689 );
nand \U$17593 ( \17970 , \17962 , \17969 );
not \U$17594 ( \17971 , \17970 );
or \U$17595 ( \17972 , \17959 , \17971 );
or \U$17596 ( \17973 , \17970 , \17958 );
not \U$17597 ( \17974 , \12945 );
not \U$17598 ( \17975 , \17845 );
or \U$17599 ( \17976 , \17974 , \17975 );
not \U$17600 ( \17977 , \11831 );
and \U$17601 ( \17978 , RIc225d50_53, \17977 );
not \U$17602 ( \17979 , RIc225d50_53);
and \U$17603 ( \17980 , \17979 , \4177 );
nor \U$17604 ( \17981 , \17978 , \17980 );
nand \U$17605 ( \17982 , \17981 , \8777 );
nand \U$17606 ( \17983 , \17976 , \17982 );
nand \U$17607 ( \17984 , \17973 , \17983 );
nand \U$17608 ( \17985 , \17972 , \17984 );
nand \U$17609 ( \17986 , \17948 , \17985 );
not \U$17610 ( \17987 , \17946 );
not \U$17611 ( \17988 , \17897 );
nand \U$17612 ( \17989 , \17987 , \17988 );
nand \U$17613 ( \17990 , \17986 , \17989 );
not \U$17614 ( \17991 , \17990 );
not \U$17615 ( \17992 , \17748 );
not \U$17616 ( \17993 , \17992 );
not \U$17617 ( \17994 , \17993 );
not \U$17618 ( \17995 , \17758 );
or \U$17619 ( \17996 , \17994 , \17995 );
not \U$17620 ( \17997 , \17992 );
not \U$17621 ( \17998 , \17757 );
or \U$17622 ( \17999 , \17997 , \17998 );
nand \U$17623 ( \18000 , \17999 , \17764 );
nand \U$17624 ( \18001 , \17996 , \18000 );
not \U$17625 ( \18002 , \16888 );
not \U$17626 ( \18003 , \18002 );
not \U$17627 ( \18004 , \16882 );
and \U$17628 ( \18005 , \18003 , \18004 );
and \U$17629 ( \18006 , \17876 , \16891 );
nor \U$17630 ( \18007 , \18005 , \18006 );
not \U$17631 ( \18008 , \18007 );
not \U$17632 ( \18009 , \18008 );
not \U$17633 ( \18010 , \17163 );
not \U$17634 ( \18011 , \12468 );
and \U$17635 ( \18012 , \18010 , \18011 );
and \U$17636 ( \18013 , \17692 , \11965 );
nor \U$17637 ( \18014 , \18012 , \18013 );
not \U$17638 ( \18015 , \18014 );
not \U$17639 ( \18016 , \18015 );
or \U$17640 ( \18017 , \18009 , \18016 );
not \U$17641 ( \18018 , \18007 );
not \U$17642 ( \18019 , \18014 );
or \U$17643 ( \18020 , \18018 , \18019 );
not \U$17644 ( \18021 , \9552 );
not \U$17645 ( \18022 , \17310 );
or \U$17646 ( \18023 , \18021 , \18022 );
nand \U$17647 ( \18024 , \17885 , \10445 );
nand \U$17648 ( \18025 , \18023 , \18024 );
nand \U$17649 ( \18026 , \18020 , \18025 );
nand \U$17650 ( \18027 , \18017 , \18026 );
xor \U$17651 ( \18028 , \18001 , \18027 );
not \U$17652 ( \18029 , \9110 );
not \U$17653 ( \18030 , \17903 );
or \U$17654 ( \18031 , \18029 , \18030 );
nand \U$17655 ( \18032 , \17084 , \9129 );
nand \U$17656 ( \18033 , \18031 , \18032 );
not \U$17657 ( \18034 , \15164 );
not \U$17658 ( \18035 , \17917 );
or \U$17659 ( \18036 , \18034 , \18035 );
buf \U$17660 ( \18037 , \12670 );
nand \U$17661 ( \18038 , \17070 , \18037 );
nand \U$17662 ( \18039 , \18036 , \18038 );
or \U$17663 ( \18040 , \18033 , \18039 );
not \U$17664 ( \18041 , \13025 );
not \U$17665 ( \18042 , \17094 );
or \U$17666 ( \18043 , \18041 , \18042 );
nand \U$17667 ( \18044 , \17933 , \11118 );
nand \U$17668 ( \18045 , \18043 , \18044 );
nand \U$17669 ( \18046 , \18040 , \18045 );
nand \U$17670 ( \18047 , \18033 , \18039 );
nand \U$17671 ( \18048 , \18046 , \18047 );
xnor \U$17672 ( \18049 , \18028 , \18048 );
nand \U$17673 ( \18050 , \17991 , \18049 );
not \U$17674 ( \18051 , \18050 );
or \U$17675 ( \18052 , \17855 , \18051 );
not \U$17676 ( \18053 , \18049 );
nand \U$17677 ( \18054 , \18053 , \17990 );
nand \U$17678 ( \18055 , \18052 , \18054 );
and \U$17679 ( \18056 , \17777 , \18055 );
and \U$17680 ( \18057 , \17679 , \17776 );
or \U$17681 ( \18058 , \18056 , \18057 );
not \U$17682 ( \18059 , \18058 );
not \U$17683 ( \18060 , \15729 );
not \U$17684 ( \18061 , \17298 );
or \U$17685 ( \18062 , \18060 , \18061 );
and \U$17686 ( \18063 , \11582 , RIc225990_61);
not \U$17687 ( \18064 , \11582 );
and \U$17688 ( \18065 , \18064 , \10338 );
or \U$17689 ( \18066 , \18063 , \18065 );
nand \U$17690 ( \18067 , \18066 , \15719 );
nand \U$17691 ( \18068 , \18062 , \18067 );
not \U$17692 ( \18069 , \9934 );
not \U$17693 ( \18070 , RIc226110_45);
not \U$17694 ( \18071 , \5767 );
or \U$17695 ( \18072 , \18070 , \18071 );
nand \U$17696 ( \18073 , \3838 , \9379 );
nand \U$17697 ( \18074 , \18072 , \18073 );
not \U$17698 ( \18075 , \18074 );
or \U$17699 ( \18076 , \18069 , \18075 );
nand \U$17700 ( \18077 , \17184 , \9398 );
nand \U$17701 ( \18078 , \18076 , \18077 );
xor \U$17702 ( \18079 , \18068 , \18078 );
not \U$17703 ( \18080 , \9619 );
not \U$17704 ( \18081 , \17172 );
or \U$17705 ( \18082 , \18080 , \18081 );
not \U$17706 ( \18083 , RIc226020_47);
not \U$17707 ( \18084 , \2234 );
or \U$17708 ( \18085 , \18083 , \18084 );
not \U$17709 ( \18086 , \2225 );
not \U$17710 ( \18087 , \18086 );
nand \U$17711 ( \18088 , \18087 , \11607 );
nand \U$17712 ( \18089 , \18085 , \18088 );
nand \U$17713 ( \18090 , \18089 , \9641 );
nand \U$17714 ( \18091 , \18082 , \18090 );
xor \U$17715 ( \18092 , \18079 , \18091 );
not \U$17716 ( \18093 , \18092 );
and \U$17717 ( \18094 , \18074 , \15183 );
and \U$17718 ( \18095 , RIc226110_45, \17081 );
not \U$17719 ( \18096 , RIc226110_45);
and \U$17720 ( \18097 , \18096 , \2013 );
or \U$17721 ( \18098 , \18095 , \18097 );
and \U$17722 ( \18099 , \18098 , \9934 );
nor \U$17723 ( \18100 , \18094 , \18099 );
not \U$17724 ( \18101 , \18100 );
not \U$17725 ( \18102 , \15729 );
not \U$17726 ( \18103 , \18066 );
or \U$17727 ( \18104 , \18102 , \18103 );
and \U$17728 ( \18105 , RIc225990_61, \982 );
not \U$17729 ( \18106 , RIc225990_61);
and \U$17730 ( \18107 , \18106 , \981 );
or \U$17731 ( \18108 , \18105 , \18107 );
nand \U$17732 ( \18109 , \18108 , \15719 );
nand \U$17733 ( \18110 , \18104 , \18109 );
not \U$17734 ( \18111 , \18110 );
not \U$17735 ( \18112 , \18111 );
or \U$17736 ( \18113 , \18101 , \18112 );
not \U$17737 ( \18114 , \10001 );
not \U$17738 ( \18115 , RIc226020_47);
not \U$17739 ( \18116 , \4009 );
or \U$17740 ( \18117 , \18115 , \18116 );
nand \U$17741 ( \18118 , \4008 , \9373 );
nand \U$17742 ( \18119 , \18117 , \18118 );
not \U$17743 ( \18120 , \18119 );
or \U$17744 ( \18121 , \18114 , \18120 );
nand \U$17745 ( \18122 , \18089 , \9619 );
nand \U$17746 ( \18123 , \18121 , \18122 );
nand \U$17747 ( \18124 , \18113 , \18123 );
not \U$17748 ( \18125 , \18100 );
nand \U$17749 ( \18126 , \18125 , \18110 );
nand \U$17750 ( \18127 , \18124 , \18126 );
not \U$17751 ( \18128 , \18127 );
or \U$17752 ( \18129 , \18093 , \18128 );
or \U$17753 ( \18130 , \18092 , \18127 );
xor \U$17754 ( \18131 , \17799 , \17810 );
xor \U$17755 ( \18132 , \18131 , \17789 );
nand \U$17756 ( \18133 , \18130 , \18132 );
nand \U$17757 ( \18134 , \18129 , \18133 );
not \U$17758 ( \18135 , \18134 );
xor \U$17759 ( \18136 , \16893 , \16904 );
xor \U$17760 ( \18137 , \18136 , \16913 );
xor \U$17761 ( \18138 , \17053 , \17038 );
xnor \U$17762 ( \18139 , \18138 , \17048 );
and \U$17763 ( \18140 , \18137 , \18139 );
not \U$17764 ( \18141 , \18137 );
not \U$17765 ( \18142 , \18139 );
and \U$17766 ( \18143 , \18141 , \18142 );
nor \U$17767 ( \18144 , \18140 , \18143 );
xor \U$17768 ( \18145 , \16961 , \16971 );
xor \U$17769 ( \18146 , \18145 , \16982 );
buf \U$17770 ( \18147 , \18146 );
and \U$17771 ( \18148 , \18144 , \18147 );
not \U$17772 ( \18149 , \18144 );
not \U$17773 ( \18150 , \18147 );
and \U$17774 ( \18151 , \18149 , \18150 );
nor \U$17775 ( \18152 , \18148 , \18151 );
not \U$17776 ( \18153 , \18152 );
or \U$17777 ( \18154 , \18135 , \18153 );
or \U$17778 ( \18155 , \18134 , \18152 );
not \U$17779 ( \18156 , \950 );
not \U$17780 ( \18157 , RIc2273d0_5);
not \U$17781 ( \18158 , \12844 );
not \U$17782 ( \18159 , \18158 );
or \U$17783 ( \18160 , \18157 , \18159 );
not \U$17784 ( \18161 , \15629 );
nand \U$17785 ( \18162 , \18161 , \935 );
nand \U$17786 ( \18163 , \18160 , \18162 );
not \U$17787 ( \18164 , \18163 );
or \U$17788 ( \18165 , \18156 , \18164 );
not \U$17789 ( \18166 , RIc2273d0_5);
not \U$17790 ( \18167 , \12825 );
not \U$17791 ( \18168 , \18167 );
or \U$17792 ( \18169 , \18166 , \18168 );
nand \U$17793 ( \18170 , \12825 , \946 );
nand \U$17794 ( \18171 , \18169 , \18170 );
nand \U$17795 ( \18172 , \18171 , \954 );
nand \U$17796 ( \18173 , \18165 , \18172 );
not \U$17797 ( \18174 , \18173 );
and \U$17798 ( \18175 , \17617 , \1081 );
not \U$17799 ( \18176 , \1039 );
xor \U$17800 ( \18177 , \2896 , \16256 );
nor \U$17801 ( \18178 , \18176 , \18177 );
nor \U$17802 ( \18179 , \18175 , \18178 );
not \U$17803 ( \18180 , \18179 );
not \U$17804 ( \18181 , \16248 );
not \U$17805 ( \18182 , \18181 );
and \U$17806 ( \18183 , \18182 , \898 );
not \U$17807 ( \18184 , \18183 );
and \U$17808 ( \18185 , \18180 , \18184 );
and \U$17809 ( \18186 , \18179 , \18183 );
nor \U$17810 ( \18187 , \18185 , \18186 );
not \U$17811 ( \18188 , \18187 );
or \U$17812 ( \18189 , \18174 , \18188 );
or \U$17813 ( \18190 , \18173 , \18187 );
nand \U$17814 ( \18191 , \18189 , \18190 );
not \U$17815 ( \18192 , \1678 );
not \U$17816 ( \18193 , RIc227010_13);
not \U$17817 ( \18194 , \10800 );
or \U$17818 ( \18195 , \18193 , \18194 );
nand \U$17819 ( \18196 , \9275 , \3841 );
nand \U$17820 ( \18197 , \18195 , \18196 );
not \U$17821 ( \18198 , \18197 );
or \U$17822 ( \18199 , \18192 , \18198 );
not \U$17823 ( \18200 , RIc227010_13);
not \U$17824 ( \18201 , \9255 );
or \U$17825 ( \18202 , \18200 , \18201 );
nand \U$17826 ( \18203 , \10986 , \1296 );
nand \U$17827 ( \18204 , \18202 , \18203 );
nand \U$17828 ( \18205 , \18204 , \1682 );
nand \U$17829 ( \18206 , \18199 , \18205 );
xor \U$17830 ( \18207 , \18191 , \18206 );
not \U$17831 ( \18208 , \1306 );
not \U$17832 ( \18209 , RIc227100_11);
not \U$17833 ( \18210 , \9321 );
or \U$17834 ( \18211 , \18209 , \18210 );
nand \U$17835 ( \18212 , \9324 , \1302 );
nand \U$17836 ( \18213 , \18211 , \18212 );
not \U$17837 ( \18214 , \18213 );
or \U$17838 ( \18215 , \18208 , \18214 );
and \U$17839 ( \18216 , RIc227100_11, \10266 );
not \U$17840 ( \18217 , RIc227100_11);
and \U$17841 ( \18218 , \18217 , \10263 );
nor \U$17842 ( \18219 , \18216 , \18218 );
nand \U$17843 ( \18220 , \18219 , \1311 );
nand \U$17844 ( \18221 , \18215 , \18220 );
and \U$17845 ( \18222 , \18207 , \18221 );
and \U$17846 ( \18223 , \18191 , \18206 );
or \U$17847 ( \18224 , \18222 , \18223 );
not \U$17848 ( \18225 , \9445 );
not \U$17849 ( \18226 , \17795 );
or \U$17850 ( \18227 , \18225 , \18226 );
not \U$17851 ( \18228 , RIc225e40_51);
not \U$17852 ( \18229 , \2304 );
or \U$17853 ( \18230 , \18228 , \18229 );
nand \U$17854 ( \18231 , \8989 , \11795 );
nand \U$17855 ( \18232 , \18230 , \18231 );
nand \U$17856 ( \18233 , \18232 , \9459 );
nand \U$17857 ( \18234 , \18227 , \18233 );
xor \U$17858 ( \18235 , \18224 , \18234 );
not \U$17859 ( \18236 , \5509 );
not \U$17860 ( \18237 , RIc2264d0_37);
not \U$17861 ( \18238 , \9188 );
or \U$17862 ( \18239 , \18237 , \18238 );
not \U$17863 ( \18240 , \14476 );
nand \U$17864 ( \18241 , \18240 , \4371 );
nand \U$17865 ( \18242 , \18239 , \18241 );
not \U$17866 ( \18243 , \18242 );
or \U$17867 ( \18244 , \18236 , \18243 );
nand \U$17868 ( \18245 , \17787 , \5519 );
nand \U$17869 ( \18246 , \18244 , \18245 );
and \U$17870 ( \18247 , \18235 , \18246 );
and \U$17871 ( \18248 , \18224 , \18234 );
or \U$17872 ( \18249 , \18247 , \18248 );
xor \U$17873 ( \18250 , \18008 , \18015 );
xor \U$17874 ( \18251 , \18250 , \18025 );
xor \U$17875 ( \18252 , \18249 , \18251 );
xor \U$17876 ( \18253 , \18045 , \18033 );
xor \U$17877 ( \18254 , \18253 , \18039 );
and \U$17878 ( \18255 , \18252 , \18254 );
and \U$17879 ( \18256 , \18249 , \18251 );
or \U$17880 ( \18257 , \18255 , \18256 );
nand \U$17881 ( \18258 , \18155 , \18257 );
nand \U$17882 ( \18259 , \18154 , \18258 );
not \U$17883 ( \18260 , \18259 );
not \U$17884 ( \18261 , \18146 );
nand \U$17885 ( \18262 , \18261 , \18137 );
and \U$17886 ( \18263 , \18262 , \18142 );
not \U$17887 ( \18264 , \18146 );
nor \U$17888 ( \18265 , \18264 , \18137 );
nor \U$17889 ( \18266 , \18263 , \18265 );
not \U$17890 ( \18267 , \18001 );
not \U$17891 ( \18268 , \18027 );
or \U$17892 ( \18269 , \18267 , \18268 );
or \U$17893 ( \18270 , \18027 , \18001 );
nand \U$17894 ( \18271 , \18270 , \18048 );
nand \U$17895 ( \18272 , \18269 , \18271 );
xor \U$17896 ( \18273 , \18266 , \18272 );
not \U$17897 ( \18274 , \17813 );
not \U$17898 ( \18275 , \17853 );
or \U$17899 ( \18276 , \18274 , \18275 );
or \U$17900 ( \18277 , \17813 , \17853 );
nand \U$17901 ( \18278 , \18277 , \17779 );
nand \U$17902 ( \18279 , \18276 , \18278 );
xor \U$17903 ( \18280 , \18273 , \18279 );
buf \U$17904 ( \18281 , \18280 );
nand \U$17905 ( \18282 , \18260 , \18281 );
xor \U$17906 ( \18283 , \17166 , \17176 );
xor \U$17907 ( \18284 , \18283 , \17188 );
xor \U$17908 ( \18285 , \18068 , \18078 );
and \U$17909 ( \18286 , \18285 , \18091 );
and \U$17910 ( \18287 , \18068 , \18078 );
or \U$17911 ( \18288 , \18286 , \18287 );
not \U$17912 ( \18289 , \18288 );
and \U$17913 ( \18290 , \18284 , \18289 );
not \U$17914 ( \18291 , \18284 );
and \U$17915 ( \18292 , \18291 , \18288 );
nor \U$17916 ( \18293 , \18290 , \18292 );
xor \U$17917 ( \18294 , \17238 , \17249 );
xnor \U$17918 ( \18295 , \18294 , \17262 );
xor \U$17919 ( \18296 , \18293 , \18295 );
not \U$17920 ( \18297 , \18296 );
xor \U$17921 ( \18298 , \16932 , \16941 );
xor \U$17922 ( \18299 , \18298 , \16958 );
not \U$17923 ( \18300 , \954 );
not \U$17924 ( \18301 , \16939 );
or \U$17925 ( \18302 , \18300 , \18301 );
nand \U$17926 ( \18303 , \18171 , \950 );
nand \U$17927 ( \18304 , \18302 , \18303 );
not \U$17928 ( \18305 , \18304 );
not \U$17929 ( \18306 , \1310 );
not \U$17930 ( \18307 , \17514 );
or \U$17931 ( \18308 , \18306 , \18307 );
nand \U$17932 ( \18309 , \18219 , \9904 );
nand \U$17933 ( \18310 , \18308 , \18309 );
not \U$17934 ( \18311 , \18310 );
or \U$17935 ( \18312 , \18305 , \18311 );
or \U$17936 ( \18313 , \18310 , \18304 );
not \U$17937 ( \18314 , \18183 );
not \U$17938 ( \18315 , \18179 );
not \U$17939 ( \18316 , \18315 );
or \U$17940 ( \18317 , \18314 , \18316 );
not \U$17941 ( \18318 , \18183 );
nand \U$17942 ( \18319 , \18318 , \18179 );
nand \U$17943 ( \18320 , \18173 , \18319 );
nand \U$17944 ( \18321 , \18317 , \18320 );
nand \U$17945 ( \18322 , \18313 , \18321 );
nand \U$17946 ( \18323 , \18312 , \18322 );
xor \U$17947 ( \18324 , \18299 , \18323 );
not \U$17948 ( \18325 , \1339 );
not \U$17949 ( \18326 , \17504 );
or \U$17950 ( \18327 , \18325 , \18326 );
not \U$17951 ( \18328 , RIc2271f0_9);
not \U$17952 ( \18329 , \16945 );
or \U$17953 ( \18330 , \18328 , \18329 );
nand \U$17954 ( \18331 , \10086 , \1342 );
nand \U$17955 ( \18332 , \18330 , \18331 );
nand \U$17956 ( \18333 , \1363 , \18332 );
nand \U$17957 ( \18334 , \18327 , \18333 );
not \U$17958 ( \18335 , \1682 );
not \U$17959 ( \18336 , \17528 );
or \U$17960 ( \18337 , \18335 , \18336 );
nand \U$17961 ( \18338 , \18204 , \1678 );
nand \U$17962 ( \18339 , \18337 , \18338 );
xor \U$17963 ( \18340 , \18334 , \18339 );
not \U$17964 ( \18341 , \2320 );
not \U$17965 ( \18342 , RIc226f20_15);
not \U$17966 ( \18343 , \9073 );
or \U$17967 ( \18344 , \18342 , \18343 );
nand \U$17968 ( \18345 , \9072 , \2351 );
nand \U$17969 ( \18346 , \18344 , \18345 );
not \U$17970 ( \18347 , \18346 );
or \U$17971 ( \18348 , \18341 , \18347 );
nand \U$17972 ( \18349 , \17539 , \2358 );
nand \U$17973 ( \18350 , \18348 , \18349 );
and \U$17974 ( \18351 , \18340 , \18350 );
and \U$17975 ( \18352 , \18334 , \18339 );
or \U$17976 ( \18353 , \18351 , \18352 );
xor \U$17977 ( \18354 , \18324 , \18353 );
or \U$17978 ( \18355 , RIc227448_4, RIc2273d0_5);
not \U$17979 ( \18356 , \16248 );
not \U$17980 ( \18357 , \18356 );
nand \U$17981 ( \18358 , \18355 , \18357 );
and \U$17982 ( \18359 , RIc227448_4, RIc2273d0_5);
nor \U$17983 ( \18360 , \18359 , \1032 );
and \U$17984 ( \18361 , \18358 , \18360 );
not \U$17985 ( \18362 , \1081 );
not \U$17986 ( \18363 , \18177 );
not \U$17987 ( \18364 , \18363 );
or \U$17988 ( \18365 , \18362 , \18364 );
not \U$17989 ( \18366 , \16248 );
not \U$17990 ( \18367 , \18366 );
or \U$17991 ( \18368 , \18367 , \1032 );
or \U$17992 ( \18369 , \18366 , RIc2274c0_3);
nand \U$17993 ( \18370 , \18368 , \18369 );
nand \U$17994 ( \18371 , \18370 , \1039 );
nand \U$17995 ( \18372 , \18365 , \18371 );
xor \U$17996 ( \18373 , \18361 , \18372 );
not \U$17997 ( \18374 , \954 );
not \U$17998 ( \18375 , \18163 );
or \U$17999 ( \18376 , \18374 , \18375 );
xor \U$18000 ( \18377 , \946 , \13487 );
not \U$18001 ( \18378 , \18377 );
nand \U$18002 ( \18379 , \18378 , \950 );
nand \U$18003 ( \18380 , \18376 , \18379 );
xor \U$18004 ( \18381 , \18373 , \18380 );
not \U$18005 ( \18382 , \1339 );
not \U$18006 ( \18383 , RIc2271f0_9);
not \U$18007 ( \18384 , \10369 );
or \U$18008 ( \18385 , \18383 , \18384 );
nand \U$18009 ( \18386 , \10197 , \1351 );
nand \U$18010 ( \18387 , \18385 , \18386 );
not \U$18011 ( \18388 , \18387 );
or \U$18012 ( \18389 , \18382 , \18388 );
not \U$18013 ( \18390 , RIc2271f0_9);
not \U$18014 ( \18391 , \17625 );
or \U$18015 ( \18392 , \18390 , \18391 );
nand \U$18016 ( \18393 , \13497 , \1351 );
nand \U$18017 ( \18394 , \18392 , \18393 );
nand \U$18018 ( \18395 , \18394 , \1363 );
nand \U$18019 ( \18396 , \18389 , \18395 );
and \U$18020 ( \18397 , \18381 , \18396 );
and \U$18021 ( \18398 , \18373 , \18380 );
or \U$18022 ( \18399 , \18397 , \18398 );
not \U$18023 ( \18400 , \2154 );
not \U$18024 ( \18401 , RIc226980_27);
not \U$18025 ( \18402 , \14192 );
or \U$18026 ( \18403 , \18401 , \18402 );
not \U$18027 ( \18404 , RIc226980_27);
nand \U$18028 ( \18405 , \18404 , \10126 );
nand \U$18029 ( \18406 , \18403 , \18405 );
not \U$18030 ( \18407 , \18406 );
or \U$18031 ( \18408 , \18400 , \18407 );
not \U$18032 ( \18409 , RIc226980_27);
not \U$18033 ( \18410 , \6718 );
not \U$18034 ( \18411 , \18410 );
or \U$18035 ( \18412 , \18409 , \18411 );
nand \U$18036 ( \18413 , \6718 , \2133 );
nand \U$18037 ( \18414 , \18412 , \18413 );
nand \U$18038 ( \18415 , \18414 , \2138 );
nand \U$18039 ( \18416 , \18408 , \18415 );
xor \U$18040 ( \18417 , \18399 , \18416 );
not \U$18041 ( \18418 , \9142 );
xnor \U$18042 ( \18419 , RIc226890_29, \15603 );
not \U$18043 ( \18420 , \18419 );
or \U$18044 ( \18421 , \18418 , \18420 );
and \U$18045 ( \18422 , RIc226890_29, \9765 );
not \U$18046 ( \18423 , RIc226890_29);
and \U$18047 ( \18424 , \18423 , \9875 );
or \U$18048 ( \18425 , \18422 , \18424 );
nand \U$18049 ( \18426 , \18425 , \2784 );
nand \U$18050 ( \18427 , \18421 , \18426 );
and \U$18051 ( \18428 , \18417 , \18427 );
and \U$18052 ( \18429 , \18399 , \18416 );
or \U$18053 ( \18430 , \18428 , \18429 );
not \U$18054 ( \18431 , \18430 );
not \U$18055 ( \18432 , \1963 );
not \U$18056 ( \18433 , RIc226e30_17);
not \U$18057 ( \18434 , \11405 );
or \U$18058 ( \18435 , \18433 , \18434 );
not \U$18059 ( \18436 , RIc226e30_17);
nand \U$18060 ( \18437 , \18436 , \8924 );
nand \U$18061 ( \18438 , \18435 , \18437 );
not \U$18062 ( \18439 , \18438 );
or \U$18063 ( \18440 , \18432 , \18439 );
not \U$18064 ( \18441 , RIc226e30_17);
not \U$18065 ( \18442 , \10643 );
or \U$18066 ( \18443 , \18441 , \18442 );
nand \U$18067 ( \18444 , \9050 , \1960 );
nand \U$18068 ( \18445 , \18443 , \18444 );
nand \U$18069 ( \18446 , \18445 , \1945 );
nand \U$18070 ( \18447 , \18440 , \18446 );
not \U$18071 ( \18448 , \18447 );
not \U$18072 ( \18449 , \2710 );
not \U$18073 ( \18450 , \4406 );
and \U$18074 ( \18451 , RIc2267a0_31, \18450 );
not \U$18075 ( \18452 , RIc2267a0_31);
and \U$18076 ( \18453 , \18452 , \4406 );
or \U$18077 ( \18454 , \18451 , \18453 );
not \U$18078 ( \18455 , \18454 );
or \U$18079 ( \18456 , \18449 , \18455 );
and \U$18080 ( \18457 , \2072 , \13512 );
not \U$18081 ( \18458 , \2072 );
not \U$18082 ( \18459 , \9754 );
and \U$18083 ( \18460 , \18458 , \18459 );
nor \U$18084 ( \18461 , \18457 , \18460 );
nand \U$18085 ( \18462 , \18461 , \2697 );
nand \U$18086 ( \18463 , \18456 , \18462 );
not \U$18087 ( \18464 , \18463 );
or \U$18088 ( \18465 , \18448 , \18464 );
or \U$18089 ( \18466 , \18463 , \18447 );
not \U$18090 ( \18467 , \2358 );
not \U$18091 ( \18468 , \18346 );
or \U$18092 ( \18469 , \18467 , \18468 );
not \U$18093 ( \18470 , RIc226f20_15);
not \U$18094 ( \18471 , \10111 );
or \U$18095 ( \18472 , \18470 , \18471 );
nand \U$18096 ( \18473 , \10110 , \1674 );
nand \U$18097 ( \18474 , \18472 , \18473 );
nand \U$18098 ( \18475 , \18474 , \2320 );
nand \U$18099 ( \18476 , \18469 , \18475 );
nand \U$18100 ( \18477 , \18466 , \18476 );
nand \U$18101 ( \18478 , \18465 , \18477 );
not \U$18102 ( \18479 , \18478 );
xor \U$18103 ( \18480 , \18304 , \18321 );
xnor \U$18104 ( \18481 , \18480 , \18310 );
nand \U$18105 ( \18482 , \18479 , \18481 );
not \U$18106 ( \18483 , \18482 );
or \U$18107 ( \18484 , \18431 , \18483 );
not \U$18108 ( \18485 , \18481 );
nand \U$18109 ( \18486 , \18485 , \18478 );
nand \U$18110 ( \18487 , \18484 , \18486 );
xor \U$18111 ( \18488 , \18354 , \18487 );
not \U$18112 ( \18489 , \17838 );
not \U$18113 ( \18490 , \18489 );
not \U$18114 ( \18491 , \17826 );
not \U$18115 ( \18492 , \17850 );
or \U$18116 ( \18493 , \18491 , \18492 );
or \U$18117 ( \18494 , \17826 , \17850 );
nand \U$18118 ( \18495 , \18493 , \18494 );
not \U$18119 ( \18496 , \18495 );
or \U$18120 ( \18497 , \18490 , \18496 );
or \U$18121 ( \18498 , \18489 , \18495 );
nand \U$18122 ( \18499 , \18497 , \18498 );
and \U$18123 ( \18500 , \18488 , \18499 );
and \U$18124 ( \18501 , \18354 , \18487 );
or \U$18125 ( \18502 , \18500 , \18501 );
not \U$18126 ( \18503 , \18502 );
nand \U$18127 ( \18504 , \18297 , \18503 );
not \U$18128 ( \18505 , \18504 );
xor \U$18129 ( \18506 , \18299 , \18323 );
and \U$18130 ( \18507 , \18506 , \18353 );
and \U$18131 ( \18508 , \18299 , \18323 );
or \U$18132 ( \18509 , \18507 , \18508 );
and \U$18133 ( \18510 , \17314 , \17302 );
not \U$18134 ( \18511 , \17314 );
not \U$18135 ( \18512 , \17302 );
and \U$18136 ( \18513 , \18511 , \18512 );
nor \U$18137 ( \18514 , \18510 , \18513 );
and \U$18138 ( \18515 , \18514 , \17290 );
not \U$18139 ( \18516 , \18514 );
not \U$18140 ( \18517 , \17290 );
and \U$18141 ( \18518 , \18516 , \18517 );
nor \U$18142 ( \18519 , \18515 , \18518 );
xor \U$18143 ( \18520 , \18509 , \18519 );
not \U$18144 ( \18521 , \17098 );
buf \U$18145 ( \18522 , \17086 );
not \U$18146 ( \18523 , \18522 );
or \U$18147 ( \18524 , \18521 , \18523 );
or \U$18148 ( \18525 , \18522 , \17098 );
nand \U$18149 ( \18526 , \18524 , \18525 );
and \U$18150 ( \18527 , \18526 , \17101 );
not \U$18151 ( \18528 , \18526 );
and \U$18152 ( \18529 , \18528 , \17072 );
nor \U$18153 ( \18530 , \18527 , \18529 );
xor \U$18154 ( \18531 , \18520 , \18530 );
not \U$18155 ( \18532 , \18531 );
or \U$18156 ( \18533 , \18505 , \18532 );
not \U$18157 ( \18534 , \18503 );
nand \U$18158 ( \18535 , \18534 , \18296 );
nand \U$18159 ( \18536 , \18533 , \18535 );
and \U$18160 ( \18537 , \18282 , \18536 );
nor \U$18161 ( \18538 , \18281 , \18260 );
nor \U$18162 ( \18539 , \18537 , \18538 );
not \U$18163 ( \18540 , \18539 );
not \U$18164 ( \18541 , \18540 );
or \U$18165 ( \18542 , \18059 , \18541 );
not \U$18166 ( \18543 , \18539 );
not \U$18167 ( \18544 , \18058 );
not \U$18168 ( \18545 , \18544 );
or \U$18169 ( \18546 , \18543 , \18545 );
xor \U$18170 ( \18547 , \16990 , \17059 );
xor \U$18171 ( \18548 , \18547 , \17151 );
not \U$18172 ( \18549 , \18279 );
not \U$18173 ( \18550 , \18272 );
or \U$18174 ( \18551 , \18549 , \18550 );
or \U$18175 ( \18552 , \18272 , \18279 );
not \U$18176 ( \18553 , \18266 );
nand \U$18177 ( \18554 , \18552 , \18553 );
nand \U$18178 ( \18555 , \18551 , \18554 );
xor \U$18179 ( \18556 , \18548 , \18555 );
xor \U$18180 ( \18557 , \17275 , \17326 );
xnor \U$18181 ( \18558 , \18557 , \17268 );
xor \U$18182 ( \18559 , \18556 , \18558 );
not \U$18183 ( \18560 , \18559 );
buf \U$18184 ( \18561 , \18560 );
nand \U$18185 ( \18562 , \18546 , \18561 );
nand \U$18186 ( \18563 , \18542 , \18562 );
not \U$18187 ( \18564 , \18563 );
not \U$18188 ( \18565 , \18564 );
not \U$18189 ( \18566 , \18555 );
not \U$18190 ( \18567 , \18548 );
nand \U$18191 ( \18568 , \18566 , \18567 );
not \U$18192 ( \18569 , \18558 );
and \U$18193 ( \18570 , \18568 , \18569 );
nor \U$18194 ( \18571 , \18566 , \18567 );
nor \U$18195 ( \18572 , \18570 , \18571 );
not \U$18196 ( \18573 , \18572 );
xor \U$18197 ( \18574 , \17154 , \17328 );
xor \U$18198 ( \18575 , \18574 , \17353 );
not \U$18199 ( \18576 , \18575 );
or \U$18200 ( \18577 , \18573 , \18576 );
buf \U$18201 ( \18578 , \18572 );
or \U$18202 ( \18579 , \18578 , \18575 );
nand \U$18203 ( \18580 , \18577 , \18579 );
xor \U$18204 ( \18581 , \17324 , \17316 );
xor \U$18205 ( \18582 , \18581 , \17319 );
not \U$18206 ( \18583 , \18582 );
not \U$18207 ( \18584 , \18288 );
nand \U$18208 ( \18585 , \18584 , \18295 );
and \U$18209 ( \18586 , \18585 , \18284 );
nor \U$18210 ( \18587 , \18295 , \18289 );
nor \U$18211 ( \18588 , \18586 , \18587 );
not \U$18212 ( \18589 , \18588 );
not \U$18213 ( \18590 , \18589 );
or \U$18214 ( \18591 , \18583 , \18590 );
not \U$18215 ( \18592 , \18582 );
not \U$18216 ( \18593 , \18592 );
not \U$18217 ( \18594 , \18588 );
or \U$18218 ( \18595 , \18593 , \18594 );
xor \U$18219 ( \18596 , \18509 , \18519 );
and \U$18220 ( \18597 , \18596 , \18530 );
and \U$18221 ( \18598 , \18509 , \18519 );
or \U$18222 ( \18599 , \18597 , \18598 );
nand \U$18223 ( \18600 , \18595 , \18599 );
nand \U$18224 ( \18601 , \18591 , \18600 );
not \U$18225 ( \18602 , \18601 );
xor \U$18226 ( \18603 , \17371 , \17388 );
xor \U$18227 ( \18604 , \18603 , \17403 );
not \U$18228 ( \18605 , \18604 );
or \U$18229 ( \18606 , \18602 , \18605 );
or \U$18230 ( \18607 , \18604 , \18601 );
not \U$18231 ( \18608 , \17264 );
not \U$18232 ( \18609 , \17227 );
and \U$18233 ( \18610 , \18608 , \18609 );
and \U$18234 ( \18611 , \17264 , \17227 );
nor \U$18235 ( \18612 , \18610 , \18611 );
not \U$18236 ( \18613 , \17191 );
xor \U$18237 ( \18614 , \18612 , \18613 );
not \U$18238 ( \18615 , \18614 );
not \U$18239 ( \18616 , \16878 );
and \U$18240 ( \18617 , \16988 , \18616 );
not \U$18241 ( \18618 , \16988 );
and \U$18242 ( \18619 , \18618 , \16878 );
nor \U$18243 ( \18620 , \18617 , \18619 );
xor \U$18244 ( \18621 , \18620 , \16985 );
not \U$18245 ( \18622 , \18621 );
nand \U$18246 ( \18623 , \18615 , \18622 );
xor \U$18247 ( \18624 , \17149 , \17103 );
not \U$18248 ( \18625 , \17144 );
xnor \U$18249 ( \18626 , \18624 , \18625 );
and \U$18250 ( \18627 , \18623 , \18626 );
and \U$18251 ( \18628 , \18614 , \18621 );
nor \U$18252 ( \18629 , \18627 , \18628 );
not \U$18253 ( \18630 , \18629 );
nand \U$18254 ( \18631 , \18607 , \18630 );
nand \U$18255 ( \18632 , \18606 , \18631 );
not \U$18256 ( \18633 , \18632 );
and \U$18257 ( \18634 , \18580 , \18633 );
not \U$18258 ( \18635 , \18580 );
and \U$18259 ( \18636 , \18635 , \18632 );
nor \U$18260 ( \18637 , \18634 , \18636 );
not \U$18261 ( \18638 , \18637 );
or \U$18262 ( \18639 , \18565 , \18638 );
xor \U$18263 ( \18640 , \17351 , \17332 );
xor \U$18264 ( \18641 , \18640 , \17344 );
xor \U$18265 ( \18642 , \17391 , \17395 );
xor \U$18266 ( \18643 , \18642 , \17399 );
not \U$18267 ( \18644 , \18643 );
not \U$18268 ( \18645 , \18644 );
xor \U$18269 ( \18646 , \17374 , \17386 );
xor \U$18270 ( \18647 , \18646 , \17379 );
not \U$18271 ( \18648 , \18647 );
not \U$18272 ( \18649 , \18648 );
or \U$18273 ( \18650 , \18645 , \18649 );
not \U$18274 ( \18651 , \18647 );
not \U$18275 ( \18652 , \18643 );
or \U$18276 ( \18653 , \18651 , \18652 );
xor \U$18277 ( \18654 , \17495 , \17519 );
xor \U$18278 ( \18655 , \18654 , \17557 );
and \U$18279 ( \18656 , \17139 , \17114 );
not \U$18280 ( \18657 , \17139 );
and \U$18281 ( \18658 , \18657 , \17142 );
or \U$18282 ( \18659 , \18656 , \18658 );
buf \U$18283 ( \18660 , \17127 );
xnor \U$18284 ( \18661 , \18659 , \18660 );
xor \U$18285 ( \18662 , \18655 , \18661 );
not \U$18286 ( \18663 , \2173 );
not \U$18287 ( \18664 , \17650 );
or \U$18288 ( \18665 , \18663 , \18664 );
not \U$18289 ( \18666 , RIc226a70_25);
not \U$18290 ( \18667 , \10307 );
or \U$18291 ( \18668 , \18666 , \18667 );
nand \U$18292 ( \18669 , \10141 , \1905 );
nand \U$18293 ( \18670 , \18668 , \18669 );
nand \U$18294 ( \18671 , \18670 , \2860 );
nand \U$18295 ( \18672 , \18665 , \18671 );
not \U$18296 ( \18673 , \2367 );
not \U$18297 ( \18674 , \17573 );
or \U$18298 ( \18675 , \18673 , \18674 );
not \U$18299 ( \18676 , RIc226c50_21);
not \U$18300 ( \18677 , \15684 );
or \U$18301 ( \18678 , \18676 , \18677 );
nand \U$18302 ( \18679 , \8806 , \3204 );
nand \U$18303 ( \18680 , \18678 , \18679 );
nand \U$18304 ( \18681 , \18680 , \2392 );
nand \U$18305 ( \18682 , \18675 , \18681 );
xor \U$18306 ( \18683 , \18672 , \18682 );
not \U$18307 ( \18684 , \1930 );
not \U$18308 ( \18685 , \17584 );
or \U$18309 ( \18686 , \18684 , \18685 );
not \U$18310 ( \18687 , RIc226b60_23);
not \U$18311 ( \18688 , \8857 );
or \U$18312 ( \18689 , \18687 , \18688 );
nand \U$18313 ( \18690 , \8856 , \1927 );
nand \U$18314 ( \18691 , \18689 , \18690 );
nand \U$18315 ( \18692 , \18691 , \1915 );
nand \U$18316 ( \18693 , \18686 , \18692 );
and \U$18317 ( \18694 , \18683 , \18693 );
and \U$18318 ( \18695 , \18672 , \18682 );
or \U$18319 ( \18696 , \18694 , \18695 );
and \U$18320 ( \18697 , \18361 , \18372 );
not \U$18321 ( \18698 , \1118 );
not \U$18322 ( \18699 , RIc2272e0_7);
not \U$18323 ( \18700 , \13198 );
or \U$18324 ( \18701 , \18699 , \18700 );
nand \U$18325 ( \18702 , \12755 , \1139 );
nand \U$18326 ( \18703 , \18701 , \18702 );
not \U$18327 ( \18704 , \18703 );
or \U$18328 ( \18705 , \18698 , \18704 );
nand \U$18329 ( \18706 , \17629 , \1120 );
nand \U$18330 ( \18707 , \18705 , \18706 );
xor \U$18331 ( \18708 , \18697 , \18707 );
not \U$18332 ( \18709 , \1339 );
not \U$18333 ( \18710 , \18332 );
or \U$18334 ( \18711 , \18709 , \18710 );
nand \U$18335 ( \18712 , \18387 , \1363 );
nand \U$18336 ( \18713 , \18711 , \18712 );
and \U$18337 ( \18714 , \18708 , \18713 );
and \U$18338 ( \18715 , \18697 , \18707 );
or \U$18339 ( \18716 , \18714 , \18715 );
not \U$18340 ( \18717 , \2138 );
not \U$18341 ( \18718 , \18406 );
or \U$18342 ( \18719 , \18717 , \18718 );
nand \U$18343 ( \18720 , \17553 , \2154 );
nand \U$18344 ( \18721 , \18719 , \18720 );
xor \U$18345 ( \18722 , \18716 , \18721 );
not \U$18346 ( \18723 , \2784 );
not \U$18347 ( \18724 , \18419 );
or \U$18348 ( \18725 , \18723 , \18724 );
nand \U$18349 ( \18726 , \17641 , \9142 );
nand \U$18350 ( \18727 , \18725 , \18726 );
and \U$18351 ( \18728 , \18722 , \18727 );
and \U$18352 ( \18729 , \18716 , \18721 );
or \U$18353 ( \18730 , \18728 , \18729 );
xor \U$18354 ( \18731 , \18696 , \18730 );
not \U$18355 ( \18732 , \18438 );
not \U$18356 ( \18733 , \18732 );
not \U$18357 ( \18734 , \7140 );
and \U$18358 ( \18735 , \18733 , \18734 );
and \U$18359 ( \18736 , \17746 , \1963 );
nor \U$18360 ( \18737 , \18735 , \18736 );
not \U$18361 ( \18738 , \18737 );
not \U$18362 ( \18739 , \17752 );
not \U$18363 ( \18740 , \2710 );
not \U$18364 ( \18741 , \18740 );
and \U$18365 ( \18742 , \18739 , \18741 );
and \U$18366 ( \18743 , \18454 , \2697 );
nor \U$18367 ( \18744 , \18742 , \18743 );
not \U$18368 ( \18745 , \18744 );
or \U$18369 ( \18746 , \18738 , \18745 );
not \U$18370 ( \18747 , \2534 );
not \U$18371 ( \18748 , \17598 );
or \U$18372 ( \18749 , \18747 , \18748 );
and \U$18373 ( \18750 , RIc226d40_19, \8979 );
not \U$18374 ( \18751 , RIc226d40_19);
and \U$18375 ( \18752 , \18751 , \8973 );
nor \U$18376 ( \18753 , \18750 , \18752 );
nand \U$18377 ( \18754 , \18753 , \2518 );
nand \U$18378 ( \18755 , \18749 , \18754 );
nand \U$18379 ( \18756 , \18746 , \18755 );
not \U$18380 ( \18757 , \18737 );
not \U$18381 ( \18758 , \18744 );
nand \U$18382 ( \18759 , \18757 , \18758 );
nand \U$18383 ( \18760 , \18756 , \18759 );
and \U$18384 ( \18761 , \18731 , \18760 );
and \U$18385 ( \18762 , \18696 , \18730 );
or \U$18386 ( \18763 , \18761 , \18762 );
and \U$18387 ( \18764 , \18662 , \18763 );
and \U$18388 ( \18765 , \18655 , \18661 );
or \U$18389 ( \18766 , \18764 , \18765 );
nand \U$18390 ( \18767 , \18653 , \18766 );
nand \U$18391 ( \18768 , \18650 , \18767 );
xor \U$18392 ( \18769 , \18641 , \18768 );
xor \U$18393 ( \18770 , \17663 , \17489 );
xor \U$18394 ( \18771 , \16321 , \16229 );
not \U$18395 ( \18772 , \16236 );
xor \U$18396 ( \18773 , \18771 , \18772 );
xor \U$18397 ( \18774 , \18770 , \18773 );
xnor \U$18398 ( \18775 , \18769 , \18774 );
not \U$18399 ( \18776 , \18775 );
not \U$18400 ( \18777 , \18776 );
xor \U$18401 ( \18778 , \18629 , \18601 );
xor \U$18402 ( \18779 , \18778 , \18604 );
not \U$18403 ( \18780 , \18779 );
not \U$18404 ( \18781 , \18780 );
or \U$18405 ( \18782 , \18777 , \18781 );
not \U$18406 ( \18783 , \18779 );
not \U$18407 ( \18784 , \18775 );
or \U$18408 ( \18785 , \18783 , \18784 );
and \U$18409 ( \18786 , \18626 , \18622 );
not \U$18410 ( \18787 , \18626 );
and \U$18411 ( \18788 , \18787 , \18621 );
nor \U$18412 ( \18789 , \18786 , \18788 );
and \U$18413 ( \18790 , \18789 , \18614 );
not \U$18414 ( \18791 , \18789 );
and \U$18415 ( \18792 , \18791 , \18615 );
or \U$18416 ( \18793 , \18790 , \18792 );
xor \U$18417 ( \18794 , \18582 , \18589 );
xor \U$18418 ( \18795 , \18794 , \18599 );
xor \U$18419 ( \18796 , \18793 , \18795 );
not \U$18420 ( \18797 , \18644 );
not \U$18421 ( \18798 , \18766 );
not \U$18422 ( \18799 , \18798 );
or \U$18423 ( \18800 , \18797 , \18799 );
nand \U$18424 ( \18801 , \18643 , \18766 );
nand \U$18425 ( \18802 , \18800 , \18801 );
and \U$18426 ( \18803 , \18802 , \18648 );
not \U$18427 ( \18804 , \18802 );
and \U$18428 ( \18805 , \18804 , \18647 );
nor \U$18429 ( \18806 , \18803 , \18805 );
and \U$18430 ( \18807 , \18796 , \18806 );
and \U$18431 ( \18808 , \18793 , \18795 );
or \U$18432 ( \18809 , \18807 , \18808 );
nand \U$18433 ( \18810 , \18785 , \18809 );
nand \U$18434 ( \18811 , \18782 , \18810 );
nand \U$18435 ( \18812 , \18639 , \18811 );
not \U$18436 ( \18813 , \18637 );
nand \U$18437 ( \18814 , \18813 , \18563 );
and \U$18438 ( \18815 , \18812 , \18814 );
xor \U$18439 ( \18816 , \17677 , \18815 );
not \U$18440 ( \18817 , \18578 );
not \U$18441 ( \18818 , \18817 );
not \U$18442 ( \18819 , \18575 );
not \U$18443 ( \18820 , \18819 );
not \U$18444 ( \18821 , \18820 );
or \U$18445 ( \18822 , \18818 , \18821 );
nand \U$18446 ( \18823 , \18819 , \18578 );
nand \U$18447 ( \18824 , \18823 , \18632 );
nand \U$18448 ( \18825 , \18822 , \18824 );
xor \U$18449 ( \18826 , \17356 , \16874 );
xor \U$18450 ( \18827 , \18826 , \17421 );
xor \U$18451 ( \18828 , \18825 , \18827 );
not \U$18452 ( \18829 , \18774 );
not \U$18453 ( \18830 , \18641 );
or \U$18454 ( \18831 , \18829 , \18830 );
or \U$18455 ( \18832 , \18774 , \18641 );
nand \U$18456 ( \18833 , \18832 , \18768 );
nand \U$18457 ( \18834 , \18831 , \18833 );
not \U$18458 ( \18835 , \18834 );
xor \U$18459 ( \18836 , \17369 , \17406 );
xor \U$18460 ( \18837 , \18836 , \17418 );
not \U$18461 ( \18838 , \18837 );
or \U$18462 ( \18839 , \18835 , \18838 );
or \U$18463 ( \18840 , \18834 , \18837 );
not \U$18464 ( \18841 , \17463 );
not \U$18465 ( \18842 , \18841 );
not \U$18466 ( \18843 , \17667 );
or \U$18467 ( \18844 , \18842 , \18843 );
nand \U$18468 ( \18845 , \17666 , \17463 );
nand \U$18469 ( \18846 , \18844 , \18845 );
and \U$18470 ( \18847 , \18846 , \17476 );
not \U$18471 ( \18848 , \18846 );
not \U$18472 ( \18849 , \17476 );
and \U$18473 ( \18850 , \18848 , \18849 );
nor \U$18474 ( \18851 , \18847 , \18850 );
nand \U$18475 ( \18852 , \18840 , \18851 );
nand \U$18476 ( \18853 , \18839 , \18852 );
xor \U$18477 ( \18854 , \18828 , \18853 );
and \U$18478 ( \18855 , \18816 , \18854 );
and \U$18479 ( \18856 , \17677 , \18815 );
or \U$18480 ( \18857 , \18855 , \18856 );
buf \U$18481 ( \18858 , \17461 );
not \U$18482 ( \18859 , \18858 );
not \U$18483 ( \18860 , \17676 );
or \U$18484 ( \18861 , \18859 , \18860 );
or \U$18485 ( \18862 , \18858 , \17676 );
nand \U$18486 ( \18863 , \18862 , \17669 );
nand \U$18487 ( \18864 , \18861 , \18863 );
not \U$18488 ( \18865 , \18827 );
not \U$18489 ( \18866 , \18865 );
not \U$18490 ( \18867 , \18825 );
or \U$18491 ( \18868 , \18866 , \18867 );
not \U$18492 ( \18869 , \18825 );
not \U$18493 ( \18870 , \18869 );
not \U$18494 ( \18871 , \18827 );
or \U$18495 ( \18872 , \18870 , \18871 );
nand \U$18496 ( \18873 , \18872 , \18853 );
nand \U$18497 ( \18874 , \18868 , \18873 );
xor \U$18498 ( \18875 , \18864 , \18874 );
not \U$18499 ( \18876 , \16867 );
not \U$18500 ( \18877 , \17423 );
not \U$18501 ( \18878 , \17435 );
or \U$18502 ( \18879 , \18877 , \18878 );
or \U$18503 ( \18880 , \17435 , \17423 );
nand \U$18504 ( \18881 , \18879 , \18880 );
not \U$18505 ( \18882 , \18881 );
not \U$18506 ( \18883 , \18882 );
or \U$18507 ( \18884 , \18876 , \18883 );
not \U$18508 ( \18885 , \16867 );
nand \U$18509 ( \18886 , \18881 , \18885 );
nand \U$18510 ( \18887 , \18884 , \18886 );
xnor \U$18511 ( \18888 , \18875 , \18887 );
nand \U$18512 ( \18889 , \18857 , \18888 );
not \U$18513 ( \18890 , \18889 );
xor \U$18514 ( \18891 , \18837 , \18834 );
xnor \U$18515 ( \18892 , \18891 , \18851 );
xor \U$18516 ( \18893 , \17679 , \17776 );
xor \U$18517 ( \18894 , \18893 , \18055 );
not \U$18518 ( \18895 , \18894 );
not \U$18519 ( \18896 , \18895 );
not \U$18520 ( \18897 , \18737 );
not \U$18521 ( \18898 , \18755 );
or \U$18522 ( \18899 , \18897 , \18898 );
or \U$18523 ( \18900 , \18755 , \18737 );
nand \U$18524 ( \18901 , \18899 , \18900 );
and \U$18525 ( \18902 , \18901 , \18744 );
not \U$18526 ( \18903 , \18901 );
and \U$18527 ( \18904 , \18903 , \18758 );
nor \U$18528 ( \18905 , \18902 , \18904 );
not \U$18529 ( \18906 , \18905 );
not \U$18530 ( \18907 , \18906 );
not \U$18531 ( \18908 , \12670 );
not \U$18532 ( \18909 , \17923 );
or \U$18533 ( \18910 , \18908 , \18909 );
and \U$18534 ( \18911 , RIc225a80_59, \1222 );
not \U$18535 ( \18912 , RIc225a80_59);
and \U$18536 ( \18913 , \18912 , \1439 );
or \U$18537 ( \18914 , \18911 , \18913 );
nand \U$18538 ( \18915 , \18914 , \15164 );
nand \U$18539 ( \18916 , \18910 , \18915 );
not \U$18540 ( \18917 , \18916 );
not \U$18541 ( \18918 , \9110 );
and \U$18542 ( \18919 , RIc226200_43, \15382 );
not \U$18543 ( \18920 , RIc226200_43);
and \U$18544 ( \18921 , \18920 , \2475 );
or \U$18545 ( \18922 , \18919 , \18921 );
not \U$18546 ( \18923 , \18922 );
or \U$18547 ( \18924 , \18918 , \18923 );
nand \U$18548 ( \18925 , \17910 , \9129 );
nand \U$18549 ( \18926 , \18924 , \18925 );
not \U$18550 ( \18927 , \18926 );
nand \U$18551 ( \18928 , \18917 , \18927 );
not \U$18552 ( \18929 , \9690 );
not \U$18553 ( \18930 , RIc2262f0_41);
not \U$18554 ( \18931 , \12548 );
or \U$18555 ( \18932 , \18930 , \18931 );
nand \U$18556 ( \18933 , \2720 , \10679 );
nand \U$18557 ( \18934 , \18932 , \18933 );
not \U$18558 ( \18935 , \18934 );
or \U$18559 ( \18936 , \18929 , \18935 );
nand \U$18560 ( \18937 , \17956 , \9705 );
nand \U$18561 ( \18938 , \18936 , \18937 );
and \U$18562 ( \18939 , \18928 , \18938 );
and \U$18563 ( \18940 , \18916 , \18926 );
nor \U$18564 ( \18941 , \18939 , \18940 );
not \U$18565 ( \18942 , \18941 );
not \U$18566 ( \18943 , \18942 );
or \U$18567 ( \18944 , \18907 , \18943 );
not \U$18568 ( \18945 , \18905 );
not \U$18569 ( \18946 , \18941 );
or \U$18570 ( \18947 , \18945 , \18946 );
not \U$18571 ( \18948 , \6307 );
not \U$18572 ( \18949 , \17968 );
or \U$18573 ( \18950 , \18948 , \18949 );
and \U$18574 ( \18951 , RIc2263e0_39, \5526 );
not \U$18575 ( \18952 , RIc2263e0_39);
and \U$18576 ( \18953 , \18952 , \2042 );
or \U$18577 ( \18954 , \18951 , \18953 );
nand \U$18578 ( \18955 , \18954 , \6688 );
nand \U$18579 ( \18956 , \18950 , \18955 );
not \U$18580 ( \18957 , \18956 );
not \U$18581 ( \18958 , \9555 );
not \U$18582 ( \18959 , \17981 );
or \U$18583 ( \18960 , \18958 , \18959 );
not \U$18584 ( \18961 , \2344 );
and \U$18585 ( \18962 , RIc225d50_53, \18961 );
not \U$18586 ( \18963 , RIc225d50_53);
and \U$18587 ( \18964 , \18963 , \2344 );
or \U$18588 ( \18965 , \18962 , \18964 );
nand \U$18589 ( \18966 , \18965 , \9488 );
nand \U$18590 ( \18967 , \18960 , \18966 );
not \U$18591 ( \18968 , \18967 );
nand \U$18592 ( \18969 , \18957 , \18968 );
not \U$18593 ( \18970 , \18969 );
xor \U$18594 ( \18971 , \18697 , \18707 );
xor \U$18595 ( \18972 , \18971 , \18713 );
not \U$18596 ( \18973 , \18972 );
or \U$18597 ( \18974 , \18970 , \18973 );
not \U$18598 ( \18975 , \18968 );
nand \U$18599 ( \18976 , \18975 , \18956 );
nand \U$18600 ( \18977 , \18974 , \18976 );
nand \U$18601 ( \18978 , \18947 , \18977 );
nand \U$18602 ( \18979 , \18944 , \18978 );
not \U$18603 ( \18980 , \18979 );
not \U$18604 ( \18981 , \11965 );
not \U$18605 ( \18982 , RIc225b70_57);
not \U$18606 ( \18983 , \17929 );
or \U$18607 ( \18984 , \18982 , \18983 );
nand \U$18608 ( \18985 , \3579 , \15262 );
nand \U$18609 ( \18986 , \18984 , \18985 );
not \U$18610 ( \18987 , \18986 );
or \U$18611 ( \18988 , \18981 , \18987 );
nand \U$18612 ( \18989 , \17698 , \11974 );
nand \U$18613 ( \18990 , \18988 , \18989 );
not \U$18614 ( \18991 , \15719 );
not \U$18615 ( \18992 , RIc225990_61);
not \U$18616 ( \18993 , \1020 );
not \U$18617 ( \18994 , \18993 );
or \U$18618 ( \18995 , \18992 , \18994 );
nand \U$18619 ( \18996 , \11715 , \12806 );
nand \U$18620 ( \18997 , \18995 , \18996 );
not \U$18621 ( \18998 , \18997 );
or \U$18622 ( \18999 , \18991 , \18998 );
nand \U$18623 ( \19000 , \18108 , \15729 );
nand \U$18624 ( \19001 , \18999 , \19000 );
or \U$18625 ( \19002 , \18990 , \19001 );
not \U$18626 ( \19003 , \9619 );
not \U$18627 ( \19004 , \18119 );
or \U$18628 ( \19005 , \19003 , \19004 );
and \U$18629 ( \19006 , RIc226020_47, \9408 );
not \U$18630 ( \19007 , RIc226020_47);
and \U$18631 ( \19008 , \19007 , \3834 );
or \U$18632 ( \19009 , \19006 , \19008 );
nand \U$18633 ( \19010 , \19009 , \9641 );
nand \U$18634 ( \19011 , \19005 , \19010 );
nand \U$18635 ( \19012 , \19002 , \19011 );
nand \U$18636 ( \19013 , \19001 , \18990 );
nand \U$18637 ( \19014 , \19012 , \19013 );
not \U$18638 ( \19015 , \16891 );
not \U$18639 ( \19016 , RIc2258a0_63);
not \U$18640 ( \19017 , \11582 );
or \U$18641 ( \19018 , \19016 , \19017 );
nand \U$18642 ( \19019 , \14659 , \15620 );
nand \U$18643 ( \19020 , \19018 , \19019 );
not \U$18644 ( \19021 , \19020 );
or \U$18645 ( \19022 , \19015 , \19021 );
not \U$18646 ( \19023 , \17867 );
nand \U$18647 ( \19024 , \19023 , RIc225828_64);
nand \U$18648 ( \19025 , \19022 , \19024 );
not \U$18649 ( \19026 , \19025 );
not \U$18650 ( \19027 , \9398 );
not \U$18651 ( \19028 , \18098 );
or \U$18652 ( \19029 , \19027 , \19028 );
and \U$18653 ( \19030 , \2585 , \14660 );
not \U$18654 ( \19031 , \2585 );
and \U$18655 ( \19032 , \19031 , RIc226110_45);
or \U$18656 ( \19033 , \19030 , \19032 );
nand \U$18657 ( \19034 , \19033 , \9934 );
nand \U$18658 ( \19035 , \19029 , \19034 );
not \U$18659 ( \19036 , \19035 );
or \U$18660 ( \19037 , \19026 , \19036 );
or \U$18661 ( \19038 , \19025 , \19035 );
not \U$18662 ( \19039 , \11117 );
not \U$18663 ( \19040 , RIc225c60_55);
not \U$18664 ( \19041 , \9115 );
or \U$18665 ( \19042 , \19040 , \19041 );
not \U$18666 ( \19043 , RIc225c60_55);
nand \U$18667 ( \19044 , \19043 , \3043 );
nand \U$18668 ( \19045 , \19042 , \19044 );
not \U$18669 ( \19046 , \19045 );
or \U$18670 ( \19047 , \19039 , \19046 );
nand \U$18671 ( \19048 , \17941 , \12532 );
nand \U$18672 ( \19049 , \19047 , \19048 );
nand \U$18673 ( \19050 , \19038 , \19049 );
nand \U$18674 ( \19051 , \19037 , \19050 );
or \U$18675 ( \19052 , \19014 , \19051 );
not \U$18676 ( \19053 , RIc2265c0_35);
not \U$18677 ( \19054 , \10496 );
or \U$18678 ( \19055 , \19053 , \19054 );
nand \U$18679 ( \19056 , \3725 , \3620 );
nand \U$18680 ( \19057 , \19055 , \19056 );
not \U$18681 ( \19058 , \19057 );
not \U$18682 ( \19059 , \4381 );
or \U$18683 ( \19060 , \19058 , \19059 );
not \U$18684 ( \19061 , \17860 );
nand \U$18685 ( \19062 , \19061 , \5135 );
nand \U$18686 ( \19063 , \19060 , \19062 );
not \U$18687 ( \19064 , \19063 );
not \U$18688 ( \19065 , \9444 );
not \U$18689 ( \19066 , \18232 );
or \U$18690 ( \19067 , \19065 , \19066 );
not \U$18691 ( \19068 , RIc225e40_51);
not \U$18692 ( \19069 , \13914 );
or \U$18693 ( \19070 , \19068 , \19069 );
nand \U$18694 ( \19071 , \2421 , \12423 );
nand \U$18695 ( \19072 , \19070 , \19071 );
nand \U$18696 ( \19073 , \19072 , \9459 );
nand \U$18697 ( \19074 , \19067 , \19073 );
not \U$18698 ( \19075 , \19074 );
or \U$18699 ( \19076 , \19064 , \19075 );
or \U$18700 ( \19077 , \19074 , \19063 );
not \U$18701 ( \19078 , \5519 );
not \U$18702 ( \19079 , \18242 );
or \U$18703 ( \19080 , \19078 , \19079 );
and \U$18704 ( \19081 , RIc2264d0_37, \3715 );
not \U$18705 ( \19082 , RIc2264d0_37);
and \U$18706 ( \19083 , \19082 , \3716 );
or \U$18707 ( \19084 , \19081 , \19083 );
nand \U$18708 ( \19085 , \19084 , \5509 );
nand \U$18709 ( \19086 , \19080 , \19085 );
nand \U$18710 ( \19087 , \19077 , \19086 );
nand \U$18711 ( \19088 , \19076 , \19087 );
nand \U$18712 ( \19089 , \19052 , \19088 );
nand \U$18713 ( \19090 , \19014 , \19051 );
nand \U$18714 ( \19091 , \19089 , \19090 );
not \U$18715 ( \19092 , \19091 );
or \U$18716 ( \19093 , \18980 , \19092 );
or \U$18717 ( \19094 , \19091 , \18979 );
not \U$18718 ( \19095 , \17681 );
not \U$18719 ( \19096 , \17684 );
or \U$18720 ( \19097 , \19095 , \19096 );
or \U$18721 ( \19098 , \17684 , \17681 );
nand \U$18722 ( \19099 , \19097 , \19098 );
not \U$18723 ( \19100 , \19099 );
not \U$18724 ( \19101 , \17722 );
not \U$18725 ( \19102 , \19101 );
or \U$18726 ( \19103 , \19100 , \19102 );
not \U$18727 ( \19104 , \17721 );
not \U$18728 ( \19105 , \17715 );
or \U$18729 ( \19106 , \19104 , \19105 );
not \U$18730 ( \19107 , \19099 );
nand \U$18731 ( \19108 , \19106 , \19107 );
nand \U$18732 ( \19109 , \19103 , \19108 );
nand \U$18733 ( \19110 , \19094 , \19109 );
nand \U$18734 ( \19111 , \19093 , \19110 );
xor \U$18735 ( \19112 , \18655 , \18661 );
xor \U$18736 ( \19113 , \19112 , \18763 );
xor \U$18737 ( \19114 , \19111 , \19113 );
xor \U$18738 ( \19115 , \18716 , \18721 );
xor \U$18739 ( \19116 , \19115 , \18727 );
xor \U$18740 ( \19117 , \18672 , \18682 );
xor \U$18741 ( \19118 , \19117 , \18693 );
xor \U$18742 ( \19119 , \19116 , \19118 );
xor \U$18743 ( \19120 , \18224 , \18234 );
xor \U$18744 ( \19121 , \19120 , \18246 );
and \U$18745 ( \19122 , \19119 , \19121 );
and \U$18746 ( \19123 , \19116 , \19118 );
or \U$18747 ( \19124 , \19122 , \19123 );
xnor \U$18748 ( \19125 , \17770 , \17767 );
not \U$18749 ( \19126 , \17765 );
and \U$18750 ( \19127 , \19125 , \19126 );
not \U$18751 ( \19128 , \19125 );
and \U$18752 ( \19129 , \19128 , \17765 );
nor \U$18753 ( \19130 , \19127 , \19129 );
xor \U$18754 ( \19131 , \19124 , \19130 );
xnor \U$18755 ( \19132 , \17894 , \17878 );
not \U$18756 ( \19133 , \17865 );
and \U$18757 ( \19134 , \19132 , \19133 );
not \U$18758 ( \19135 , \19132 );
and \U$18759 ( \19136 , \19135 , \17865 );
nor \U$18760 ( \19137 , \19134 , \19136 );
xor \U$18761 ( \19138 , \18110 , \18123 );
xor \U$18762 ( \19139 , \19138 , \18125 );
xor \U$18763 ( \19140 , \19137 , \19139 );
xor \U$18764 ( \19141 , \17983 , \17958 );
xor \U$18765 ( \19142 , \19141 , \17970 );
and \U$18766 ( \19143 , \19140 , \19142 );
and \U$18767 ( \19144 , \19137 , \19139 );
or \U$18768 ( \19145 , \19143 , \19144 );
and \U$18769 ( \19146 , \19131 , \19145 );
and \U$18770 ( \19147 , \19124 , \19130 );
or \U$18771 ( \19148 , \19146 , \19147 );
and \U$18772 ( \19149 , \19114 , \19148 );
and \U$18773 ( \19150 , \19111 , \19113 );
or \U$18774 ( \19151 , \19149 , \19150 );
not \U$18775 ( \19152 , \19151 );
not \U$18776 ( \19153 , \19152 );
or \U$18777 ( \19154 , \18896 , \19153 );
not \U$18778 ( \19155 , \17735 );
not \U$18779 ( \19156 , \17774 );
or \U$18780 ( \19157 , \19155 , \19156 );
nand \U$18781 ( \19158 , \17773 , \17730 );
nand \U$18782 ( \19159 , \19157 , \19158 );
and \U$18783 ( \19160 , \19159 , \17727 );
not \U$18784 ( \19161 , \19159 );
and \U$18785 ( \19162 , \19161 , \17733 );
nor \U$18786 ( \19163 , \19160 , \19162 );
xor \U$18787 ( \19164 , \18334 , \18339 );
xor \U$18788 ( \19165 , \19164 , \18350 );
not \U$18789 ( \19166 , \2195 );
not \U$18790 ( \19167 , RIc226a70_25);
not \U$18791 ( \19168 , \9884 );
or \U$18792 ( \19169 , \19167 , \19168 );
nand \U$18793 ( \19170 , \8885 , \1905 );
nand \U$18794 ( \19171 , \19169 , \19170 );
not \U$18795 ( \19172 , \19171 );
or \U$18796 ( \19173 , \19166 , \19172 );
nand \U$18797 ( \19174 , \18670 , \2172 );
nand \U$18798 ( \19175 , \19173 , \19174 );
not \U$18799 ( \19176 , \19175 );
not \U$18800 ( \19177 , \2392 );
not \U$18801 ( \19178 , RIc226c50_21);
not \U$18802 ( \19179 , \11565 );
or \U$18803 ( \19180 , \19178 , \19179 );
nand \U$18804 ( \19181 , \8951 , \2370 );
nand \U$18805 ( \19182 , \19180 , \19181 );
not \U$18806 ( \19183 , \19182 );
or \U$18807 ( \19184 , \19177 , \19183 );
nand \U$18808 ( \19185 , \18680 , \2367 );
nand \U$18809 ( \19186 , \19184 , \19185 );
not \U$18810 ( \19187 , \19186 );
or \U$18811 ( \19188 , \19176 , \19187 );
or \U$18812 ( \19189 , \19186 , \19175 );
not \U$18813 ( \19190 , \1930 );
not \U$18814 ( \19191 , \18691 );
or \U$18815 ( \19192 , \19190 , \19191 );
and \U$18816 ( \19193 , \8829 , \1927 );
not \U$18817 ( \19194 , \8829 );
and \U$18818 ( \19195 , \19194 , RIc226b60_23);
or \U$18819 ( \19196 , \19193 , \19195 );
nand \U$18820 ( \19197 , \19196 , \1915 );
nand \U$18821 ( \19198 , \19192 , \19197 );
nand \U$18822 ( \19199 , \19189 , \19198 );
nand \U$18823 ( \19200 , \19188 , \19199 );
xor \U$18824 ( \19201 , \19165 , \19200 );
not \U$18825 ( \19202 , \4121 );
not \U$18826 ( \19203 , \9943 );
and \U$18827 ( \19204 , \19202 , \19203 );
and \U$18828 ( \19205 , \4121 , \5179 );
nor \U$18829 ( \19206 , \19204 , \19205 );
not \U$18830 ( \19207 , \19206 );
not \U$18831 ( \19208 , \5185 );
and \U$18832 ( \19209 , \19207 , \19208 );
and \U$18833 ( \19210 , \17712 , \3631 );
nor \U$18834 ( \19211 , \19209 , \19210 );
not \U$18835 ( \19212 , \2518 );
and \U$18836 ( \19213 , RIc226d40_19, \8913 );
not \U$18837 ( \19214 , RIc226d40_19);
and \U$18838 ( \19215 , \19214 , \8910 );
nor \U$18839 ( \19216 , \19213 , \19215 );
not \U$18840 ( \19217 , \19216 );
or \U$18841 ( \19218 , \19212 , \19217 );
nand \U$18842 ( \19219 , \18753 , \2534 );
nand \U$18843 ( \19220 , \19218 , \19219 );
not \U$18844 ( \19221 , \19220 );
nand \U$18845 ( \19222 , \19211 , \19221 );
not \U$18846 ( \19223 , \19222 );
not \U$18847 ( \19224 , \10445 );
not \U$18848 ( \19225 , RIc225f30_49);
not \U$18849 ( \19226 , \2225 );
not \U$18850 ( \19227 , \19226 );
or \U$18851 ( \19228 , \19225 , \19227 );
nand \U$18852 ( \19229 , \11648 , \11289 );
nand \U$18853 ( \19230 , \19228 , \19229 );
not \U$18854 ( \19231 , \19230 );
or \U$18855 ( \19232 , \19224 , \19231 );
nand \U$18856 ( \19233 , \17892 , \9552 );
nand \U$18857 ( \19234 , \19232 , \19233 );
not \U$18858 ( \19235 , \19234 );
or \U$18859 ( \19236 , \19223 , \19235 );
or \U$18860 ( \19237 , \19211 , \19221 );
nand \U$18861 ( \19238 , \19236 , \19237 );
and \U$18862 ( \19239 , \19201 , \19238 );
and \U$18863 ( \19240 , \19165 , \19200 );
or \U$18864 ( \19241 , \19239 , \19240 );
xor \U$18865 ( \19242 , \18696 , \18730 );
xor \U$18866 ( \19243 , \19242 , \18760 );
xor \U$18867 ( \19244 , \19241 , \19243 );
and \U$18868 ( \19245 , \17985 , \17946 );
not \U$18869 ( \19246 , \17985 );
and \U$18870 ( \19247 , \19246 , \17987 );
or \U$18871 ( \19248 , \19245 , \19247 );
and \U$18872 ( \19249 , \19248 , \17988 );
not \U$18873 ( \19250 , \19248 );
and \U$18874 ( \19251 , \19250 , \17897 );
nor \U$18875 ( \19252 , \19249 , \19251 );
and \U$18876 ( \19253 , \19244 , \19252 );
and \U$18877 ( \19254 , \19241 , \19243 );
or \U$18878 ( \19255 , \19253 , \19254 );
xor \U$18879 ( \19256 , \19163 , \19255 );
and \U$18880 ( \19257 , \18134 , \18152 );
not \U$18881 ( \19258 , \18134 );
not \U$18882 ( \19259 , \18152 );
and \U$18883 ( \19260 , \19258 , \19259 );
nor \U$18884 ( \19261 , \19257 , \19260 );
and \U$18885 ( \19262 , \19261 , \18257 );
not \U$18886 ( \19263 , \19261 );
not \U$18887 ( \19264 , \18257 );
and \U$18888 ( \19265 , \19263 , \19264 );
nor \U$18889 ( \19266 , \19262 , \19265 );
and \U$18890 ( \19267 , \19256 , \19266 );
and \U$18891 ( \19268 , \19163 , \19255 );
or \U$18892 ( \19269 , \19267 , \19268 );
nand \U$18893 ( \19270 , \19154 , \19269 );
nand \U$18894 ( \19271 , \18894 , \19151 );
nand \U$18895 ( \19272 , \19270 , \19271 );
not \U$18896 ( \19273 , \19272 );
not \U$18897 ( \19274 , \19273 );
not \U$18898 ( \19275 , \18544 );
not \U$18899 ( \19276 , \18560 );
or \U$18900 ( \19277 , \19275 , \19276 );
nand \U$18901 ( \19278 , \18559 , \18058 );
nand \U$18902 ( \19279 , \19277 , \19278 );
buf \U$18903 ( \19280 , \18539 );
and \U$18904 ( \19281 , \19279 , \19280 );
not \U$18905 ( \19282 , \19279 );
and \U$18906 ( \19283 , \19282 , \18540 );
nor \U$18907 ( \19284 , \19281 , \19283 );
not \U$18908 ( \19285 , \19284 );
or \U$18909 ( \19286 , \19274 , \19285 );
not \U$18910 ( \19287 , \18536 );
xor \U$18911 ( \19288 , \18280 , \18259 );
not \U$18912 ( \19289 , \19288 );
or \U$18913 ( \19290 , \19287 , \19289 );
or \U$18914 ( \19291 , \19288 , \18536 );
nand \U$18915 ( \19292 , \19290 , \19291 );
xor \U$18916 ( \19293 , \17990 , \18053 );
xor \U$18917 ( \19294 , \19293 , \17854 );
not \U$18918 ( \19295 , \19294 );
not \U$18919 ( \19296 , \19295 );
xor \U$18920 ( \19297 , \18502 , \18531 );
xnor \U$18921 ( \19298 , \19297 , \18296 );
not \U$18922 ( \19299 , \19298 );
or \U$18923 ( \19300 , \19296 , \19299 );
xor \U$18924 ( \19301 , \17720 , \17700 );
xnor \U$18925 ( \19302 , \19301 , \17714 );
buf \U$18926 ( \19303 , \19302 );
xor \U$18927 ( \19304 , \17943 , \17912 );
xor \U$18928 ( \19305 , \19304 , \17925 );
or \U$18929 ( \19306 , \19303 , \19305 );
xor \U$18930 ( \19307 , \18476 , \18447 );
xnor \U$18931 ( \19308 , \19307 , \18463 );
not \U$18932 ( \19309 , \19308 );
not \U$18933 ( \19310 , \2518 );
not \U$18934 ( \19311 , RIc226d40_19);
not \U$18935 ( \19312 , \9215 );
or \U$18936 ( \19313 , \19311 , \19312 );
nand \U$18937 ( \19314 , \8924 , \1941 );
nand \U$18938 ( \19315 , \19313 , \19314 );
not \U$18939 ( \19316 , \19315 );
or \U$18940 ( \19317 , \19310 , \19316 );
nand \U$18941 ( \19318 , \19216 , \2534 );
nand \U$18942 ( \19319 , \19317 , \19318 );
not \U$18943 ( \19320 , \19319 );
and \U$18944 ( \19321 , \19182 , \2367 );
not \U$18945 ( \19322 , RIc226c50_21);
not \U$18946 ( \19323 , \8975 );
or \U$18947 ( \19324 , \19322 , \19323 );
nand \U$18948 ( \19325 , \8979 , \3204 );
nand \U$18949 ( \19326 , \19324 , \19325 );
and \U$18950 ( \19327 , \19326 , \2392 );
nor \U$18951 ( \19328 , \19321 , \19327 );
not \U$18952 ( \19329 , \19328 );
not \U$18953 ( \19330 , \19329 );
or \U$18954 ( \19331 , \19320 , \19330 );
not \U$18955 ( \19332 , \19319 );
not \U$18956 ( \19333 , \19332 );
not \U$18957 ( \19334 , \19328 );
or \U$18958 ( \19335 , \19333 , \19334 );
not \U$18959 ( \19336 , \3629 );
not \U$18960 ( \19337 , RIc2266b0_33);
not \U$18961 ( \19338 , \18450 );
or \U$18962 ( \19339 , \19337 , \19338 );
nand \U$18963 ( \19340 , \4406 , \2692 );
nand \U$18964 ( \19341 , \19339 , \19340 );
not \U$18965 ( \19342 , \19341 );
or \U$18966 ( \19343 , \19336 , \19342 );
not \U$18967 ( \19344 , \19206 );
nand \U$18968 ( \19345 , \19344 , \3631 );
nand \U$18969 ( \19346 , \19343 , \19345 );
nand \U$18970 ( \19347 , \19335 , \19346 );
nand \U$18971 ( \19348 , \19331 , \19347 );
not \U$18972 ( \19349 , \19348 );
not \U$18973 ( \19350 , \19349 );
or \U$18974 ( \19351 , \19309 , \19350 );
not \U$18975 ( \19352 , RIc226a70_25);
not \U$18976 ( \19353 , \10322 );
or \U$18977 ( \19354 , \19352 , \19353 );
nand \U$18978 ( \19355 , \8856 , \2187 );
nand \U$18979 ( \19356 , \19354 , \19355 );
and \U$18980 ( \19357 , \19356 , \2195 );
and \U$18981 ( \19358 , \19171 , \2173 );
nor \U$18982 ( \19359 , \19357 , \19358 );
not \U$18983 ( \19360 , \19359 );
not \U$18984 ( \19361 , \19360 );
and \U$18985 ( \19362 , \8806 , \10210 );
not \U$18986 ( \19363 , \8806 );
and \U$18987 ( \19364 , \19363 , RIc226b60_23);
or \U$18988 ( \19365 , \19362 , \19364 );
not \U$18989 ( \19366 , \19365 );
not \U$18990 ( \19367 , \10214 );
or \U$18991 ( \19368 , \19366 , \19367 );
nand \U$18992 ( \19369 , \19196 , \1930 );
nand \U$18993 ( \19370 , \19368 , \19369 );
not \U$18994 ( \19371 , \19370 );
or \U$18995 ( \19372 , \19361 , \19371 );
not \U$18996 ( \19373 , \19370 );
not \U$18997 ( \19374 , \19373 );
not \U$18998 ( \19375 , \19359 );
or \U$18999 ( \19376 , \19374 , \19375 );
not \U$19000 ( \19377 , \2154 );
not \U$19001 ( \19378 , \18414 );
or \U$19002 ( \19379 , \19377 , \19378 );
not \U$19003 ( \19380 , RIc226980_27);
not \U$19004 ( \19381 , \10307 );
or \U$19005 ( \19382 , \19380 , \19381 );
nand \U$19006 ( \19383 , \9731 , \2799 );
nand \U$19007 ( \19384 , \19382 , \19383 );
nand \U$19008 ( \19385 , \19384 , \2138 );
nand \U$19009 ( \19386 , \19379 , \19385 );
nand \U$19010 ( \19387 , \19376 , \19386 );
nand \U$19011 ( \19388 , \19372 , \19387 );
nand \U$19012 ( \19389 , \19351 , \19388 );
not \U$19013 ( \19390 , \19308 );
nand \U$19014 ( \19391 , \19348 , \19390 );
nand \U$19015 ( \19392 , \19389 , \19391 );
nand \U$19016 ( \19393 , \19306 , \19392 );
nand \U$19017 ( \19394 , \19305 , \19303 );
nand \U$19018 ( \19395 , \19393 , \19394 );
not \U$19019 ( \19396 , \19395 );
not \U$19020 ( \19397 , \19396 );
xor \U$19021 ( \19398 , \18127 , \18132 );
xnor \U$19022 ( \19399 , \19398 , \18092 );
not \U$19023 ( \19400 , \19399 );
or \U$19024 ( \19401 , \19397 , \19400 );
xor \U$19025 ( \19402 , \18249 , \18251 );
xor \U$19026 ( \19403 , \19402 , \18254 );
nand \U$19027 ( \19404 , \19401 , \19403 );
not \U$19028 ( \19405 , \19396 );
not \U$19029 ( \19406 , \19399 );
nand \U$19030 ( \19407 , \19405 , \19406 );
nand \U$19031 ( \19408 , \19404 , \19407 );
nand \U$19032 ( \19409 , \19300 , \19408 );
not \U$19033 ( \19410 , \19295 );
not \U$19034 ( \19411 , \19298 );
nand \U$19035 ( \19412 , \19410 , \19411 );
nand \U$19036 ( \19413 , \19409 , \19412 );
xor \U$19037 ( \19414 , \19292 , \19413 );
xor \U$19038 ( \19415 , \18793 , \18795 );
xor \U$19039 ( \19416 , \19415 , \18806 );
and \U$19040 ( \19417 , \19414 , \19416 );
and \U$19041 ( \19418 , \19292 , \19413 );
or \U$19042 ( \19419 , \19417 , \19418 );
nand \U$19043 ( \19420 , \19286 , \19419 );
not \U$19044 ( \19421 , \19284 );
nand \U$19045 ( \19422 , \19421 , \19272 );
and \U$19046 ( \19423 , \19420 , \19422 );
xor \U$19047 ( \19424 , \18892 , \19423 );
not \U$19048 ( \19425 , \18563 );
not \U$19049 ( \19426 , \18637 );
or \U$19050 ( \19427 , \19425 , \19426 );
or \U$19051 ( \19428 , \18563 , \18637 );
nand \U$19052 ( \19429 , \19427 , \19428 );
not \U$19053 ( \19430 , \18811 );
and \U$19054 ( \19431 , \19429 , \19430 );
not \U$19055 ( \19432 , \19429 );
and \U$19056 ( \19433 , \19432 , \18811 );
nor \U$19057 ( \19434 , \19431 , \19433 );
xor \U$19058 ( \19435 , \19424 , \19434 );
xor \U$19059 ( \19436 , \18779 , \18809 );
buf \U$19060 ( \19437 , \18775 );
xnor \U$19061 ( \19438 , \19436 , \19437 );
xor \U$19062 ( \19439 , \19163 , \19255 );
xor \U$19063 ( \19440 , \19439 , \19266 );
not \U$19064 ( \19441 , \19440 );
not \U$19065 ( \19442 , \19441 );
not \U$19066 ( \19443 , \19294 );
not \U$19067 ( \19444 , \19408 );
not \U$19068 ( \19445 , \19444 );
or \U$19069 ( \19446 , \19443 , \19445 );
nand \U$19070 ( \19447 , \19295 , \19408 );
nand \U$19071 ( \19448 , \19446 , \19447 );
and \U$19072 ( \19449 , \19448 , \19298 );
not \U$19073 ( \19450 , \19448 );
and \U$19074 ( \19451 , \19450 , \19411 );
nor \U$19075 ( \19452 , \19449 , \19451 );
not \U$19076 ( \19453 , \19452 );
or \U$19077 ( \19454 , \19442 , \19453 );
xor \U$19078 ( \19455 , \19124 , \19130 );
xor \U$19079 ( \19456 , \19455 , \19145 );
and \U$19080 ( \19457 , \18942 , \18906 );
not \U$19081 ( \19458 , \18942 );
and \U$19082 ( \19459 , \19458 , \18905 );
nor \U$19083 ( \19460 , \19457 , \19459 );
and \U$19084 ( \19461 , \19460 , \18977 );
not \U$19085 ( \19462 , \19460 );
not \U$19086 ( \19463 , \18977 );
and \U$19087 ( \19464 , \19462 , \19463 );
nor \U$19088 ( \19465 , \19461 , \19464 );
xor \U$19089 ( \19466 , \19116 , \19118 );
xor \U$19090 ( \19467 , \19466 , \19121 );
xor \U$19091 ( \19468 , \19465 , \19467 );
xor \U$19092 ( \19469 , \19137 , \19139 );
xor \U$19093 ( \19470 , \19469 , \19142 );
and \U$19094 ( \19471 , \19468 , \19470 );
and \U$19095 ( \19472 , \19465 , \19467 );
or \U$19096 ( \19473 , \19471 , \19472 );
xor \U$19097 ( \19474 , \19456 , \19473 );
xor \U$19098 ( \19475 , \19395 , \19403 );
xor \U$19099 ( \19476 , \19475 , \19406 );
and \U$19100 ( \19477 , \19474 , \19476 );
and \U$19101 ( \19478 , \19456 , \19473 );
or \U$19102 ( \19479 , \19477 , \19478 );
nand \U$19103 ( \19480 , \19454 , \19479 );
not \U$19104 ( \19481 , \19441 );
not \U$19105 ( \19482 , \19452 );
nand \U$19106 ( \19483 , \19481 , \19482 );
nand \U$19107 ( \19484 , \19480 , \19483 );
not \U$19108 ( \19485 , \19484 );
not \U$19109 ( \19486 , \19151 );
not \U$19110 ( \19487 , \18895 );
or \U$19111 ( \19488 , \19486 , \19487 );
nand \U$19112 ( \19489 , \19152 , \18894 );
nand \U$19113 ( \19490 , \19488 , \19489 );
not \U$19114 ( \19491 , \19269 );
and \U$19115 ( \19492 , \19490 , \19491 );
not \U$19116 ( \19493 , \19490 );
and \U$19117 ( \19494 , \19493 , \19269 );
nor \U$19118 ( \19495 , \19492 , \19494 );
not \U$19119 ( \19496 , \19495 );
not \U$19120 ( \19497 , \19496 );
nand \U$19121 ( \19498 , \19485 , \19497 );
xor \U$19122 ( \19499 , \18354 , \18487 );
xor \U$19123 ( \19500 , \19499 , \18499 );
not \U$19124 ( \19501 , \19500 );
not \U$19125 ( \19502 , \18430 );
xor \U$19126 ( \19503 , \18478 , \18481 );
not \U$19127 ( \19504 , \19503 );
or \U$19128 ( \19505 , \19502 , \19504 );
or \U$19129 ( \19506 , \18430 , \19503 );
nand \U$19130 ( \19507 , \19505 , \19506 );
xor \U$19131 ( \19508 , \19165 , \19200 );
xor \U$19132 ( \19509 , \19508 , \19238 );
or \U$19133 ( \19510 , \19507 , \19509 );
xor \U$19134 ( \19511 , \18191 , \18206 );
xor \U$19135 ( \19512 , \19511 , \18221 );
not \U$19136 ( \19513 , \19512 );
not \U$19137 ( \19514 , \11974 );
not \U$19138 ( \19515 , \18986 );
or \U$19139 ( \19516 , \19514 , \19515 );
not \U$19140 ( \19517 , RIc225b70_57);
not \U$19141 ( \19518 , \10909 );
or \U$19142 ( \19519 , \19517 , \19518 );
nand \U$19143 ( \19520 , \1331 , \11033 );
nand \U$19144 ( \19521 , \19519 , \19520 );
nand \U$19145 ( \19522 , \19521 , \11965 );
nand \U$19146 ( \19523 , \19516 , \19522 );
not \U$19147 ( \19524 , \10953 );
not \U$19148 ( \19525 , \19009 );
or \U$19149 ( \19526 , \19524 , \19525 );
not \U$19150 ( \19527 , \11607 );
not \U$19151 ( \19528 , \3508 );
or \U$19152 ( \19529 , \19527 , \19528 );
not \U$19153 ( \19530 , \9434 );
nand \U$19154 ( \19531 , \19530 , RIc226020_47);
nand \U$19155 ( \19532 , \19529 , \19531 );
nand \U$19156 ( \19533 , \19532 , \9641 );
nand \U$19157 ( \19534 , \19526 , \19533 );
xor \U$19158 ( \19535 , \19523 , \19534 );
not \U$19159 ( \19536 , \9458 );
not \U$19160 ( \19537 , RIc225e40_51);
not \U$19161 ( \19538 , \2444 );
or \U$19162 ( \19539 , \19537 , \19538 );
nand \U$19163 ( \19540 , \5269 , \11795 );
nand \U$19164 ( \19541 , \19539 , \19540 );
not \U$19165 ( \19542 , \19541 );
or \U$19166 ( \19543 , \19536 , \19542 );
nand \U$19167 ( \19544 , \19072 , \9444 );
nand \U$19168 ( \19545 , \19543 , \19544 );
and \U$19169 ( \19546 , \19535 , \19545 );
and \U$19170 ( \19547 , \19523 , \19534 );
or \U$19171 ( \19548 , \19546 , \19547 );
not \U$19172 ( \19549 , \19548 );
or \U$19173 ( \19550 , \19513 , \19549 );
or \U$19174 ( \19551 , \19548 , \19512 );
xor \U$19175 ( \19552 , \18373 , \18380 );
xor \U$19176 ( \19553 , \19552 , \18396 );
not \U$19177 ( \19554 , \15719 );
and \U$19178 ( \19555 , \17161 , RIc225990_61);
not \U$19179 ( \19556 , \17161 );
and \U$19180 ( \19557 , \19556 , \12806 );
or \U$19181 ( \19558 , \19555 , \19557 );
not \U$19182 ( \19559 , \19558 );
or \U$19183 ( \19560 , \19554 , \19559 );
nand \U$19184 ( \19561 , \18997 , \15729 );
nand \U$19185 ( \19562 , \19560 , \19561 );
xor \U$19186 ( \19563 , \19553 , \19562 );
not \U$19187 ( \19564 , \9534 );
not \U$19188 ( \19565 , RIc225f30_49);
not \U$19189 ( \19566 , \4009 );
or \U$19190 ( \19567 , \19565 , \19566 );
nand \U$19191 ( \19568 , \4008 , \11289 );
nand \U$19192 ( \19569 , \19567 , \19568 );
not \U$19193 ( \19570 , \19569 );
or \U$19194 ( \19571 , \19564 , \19570 );
nand \U$19195 ( \19572 , \19230 , \9552 );
nand \U$19196 ( \19573 , \19571 , \19572 );
and \U$19197 ( \19574 , \19563 , \19573 );
and \U$19198 ( \19575 , \19553 , \19562 );
or \U$19199 ( \19576 , \19574 , \19575 );
nand \U$19200 ( \19577 , \19551 , \19576 );
nand \U$19201 ( \19578 , \19550 , \19577 );
nand \U$19202 ( \19579 , \19510 , \19578 );
nand \U$19203 ( \19580 , \19509 , \19507 );
nand \U$19204 ( \19581 , \19579 , \19580 );
not \U$19205 ( \19582 , \19581 );
or \U$19206 ( \19583 , \19501 , \19582 );
not \U$19207 ( \19584 , \19500 );
not \U$19208 ( \19585 , \19584 );
not \U$19209 ( \19586 , \19581 );
not \U$19210 ( \19587 , \19586 );
or \U$19211 ( \19588 , \19585 , \19587 );
not \U$19212 ( \19589 , \9555 );
not \U$19213 ( \19590 , \18965 );
or \U$19214 ( \19591 , \19589 , \19590 );
and \U$19215 ( \19592 , RIc225d50_53, \2297 );
not \U$19216 ( \19593 , RIc225d50_53);
and \U$19217 ( \19594 , \19593 , \10934 );
nor \U$19218 ( \19595 , \19592 , \19594 );
nand \U$19219 ( \19596 , \19595 , \8777 );
nand \U$19220 ( \19597 , \19591 , \19596 );
not \U$19221 ( \19598 , \19597 );
not \U$19222 ( \19599 , \5519 );
not \U$19223 ( \19600 , \19084 );
or \U$19224 ( \19601 , \19599 , \19600 );
not \U$19225 ( \19602 , RIc2264d0_37);
not \U$19226 ( \19603 , \13102 );
or \U$19227 ( \19604 , \19602 , \19603 );
nand \U$19228 ( \19605 , \3115 , \5504 );
nand \U$19229 ( \19606 , \19604 , \19605 );
nand \U$19230 ( \19607 , \19606 , \5509 );
nand \U$19231 ( \19608 , \19601 , \19607 );
not \U$19232 ( \19609 , \19608 );
or \U$19233 ( \19610 , \19598 , \19609 );
or \U$19234 ( \19611 , \19597 , \19608 );
not \U$19235 ( \19612 , \6689 );
xor \U$19236 ( \19613 , RIc2263e0_39, \2634 );
not \U$19237 ( \19614 , \19613 );
or \U$19238 ( \19615 , \19612 , \19614 );
nand \U$19239 ( \19616 , \18954 , \6307 );
nand \U$19240 ( \19617 , \19615 , \19616 );
nand \U$19241 ( \19618 , \19611 , \19617 );
nand \U$19242 ( \19619 , \19610 , \19618 );
not \U$19243 ( \19620 , \16891 );
not \U$19244 ( \19621 , RIc2258a0_63);
not \U$19245 ( \19622 , \1557 );
or \U$19246 ( \19623 , \19621 , \19622 );
nand \U$19247 ( \19624 , \3464 , \15620 );
nand \U$19248 ( \19625 , \19623 , \19624 );
not \U$19249 ( \19626 , \19625 );
or \U$19250 ( \19627 , \19620 , \19626 );
nand \U$19251 ( \19628 , \19020 , RIc225828_64);
nand \U$19252 ( \19629 , \19627 , \19628 );
not \U$19253 ( \19630 , \19629 );
not \U$19254 ( \19631 , \9934 );
not \U$19255 ( \19632 , RIc226110_45);
not \U$19256 ( \19633 , \10896 );
or \U$19257 ( \19634 , \19632 , \19633 );
not \U$19258 ( \19635 , RIc226110_45);
nand \U$19259 ( \19636 , \19635 , \10899 );
nand \U$19260 ( \19637 , \19634 , \19636 );
not \U$19261 ( \19638 , \19637 );
or \U$19262 ( \19639 , \19631 , \19638 );
nand \U$19263 ( \19640 , \19033 , \9398 );
nand \U$19264 ( \19641 , \19639 , \19640 );
not \U$19265 ( \19642 , \19641 );
or \U$19266 ( \19643 , \19630 , \19642 );
or \U$19267 ( \19644 , \19629 , \19641 );
not \U$19268 ( \19645 , \11118 );
and \U$19269 ( \19646 , RIc225c60_55, \11831 );
not \U$19270 ( \19647 , RIc225c60_55);
and \U$19271 ( \19648 , \19647 , \1729 );
or \U$19272 ( \19649 , \19646 , \19648 );
not \U$19273 ( \19650 , \19649 );
or \U$19274 ( \19651 , \19645 , \19650 );
nand \U$19275 ( \19652 , \19045 , \12532 );
nand \U$19276 ( \19653 , \19651 , \19652 );
nand \U$19277 ( \19654 , \19644 , \19653 );
nand \U$19278 ( \19655 , \19643 , \19654 );
nor \U$19279 ( \19656 , \19619 , \19655 );
xor \U$19280 ( \19657 , \18399 , \18416 );
xor \U$19281 ( \19658 , \19657 , \18427 );
not \U$19282 ( \19659 , \19658 );
or \U$19283 ( \19660 , \19656 , \19659 );
nand \U$19284 ( \19661 , \19619 , \19655 );
nand \U$19285 ( \19662 , \19660 , \19661 );
not \U$19286 ( \19663 , \19662 );
not \U$19287 ( \19664 , \19663 );
and \U$19288 ( \19665 , \19211 , \19221 );
not \U$19289 ( \19666 , \19211 );
and \U$19290 ( \19667 , \19666 , \19220 );
nor \U$19291 ( \19668 , \19665 , \19667 );
xnor \U$19292 ( \19669 , \19234 , \19668 );
xor \U$19293 ( \19670 , \19186 , \19198 );
xnor \U$19294 ( \19671 , \19670 , \19175 );
nand \U$19295 ( \19672 , \19669 , \19671 );
not \U$19296 ( \19673 , \12670 );
not \U$19297 ( \19674 , \18914 );
or \U$19298 ( \19675 , \19673 , \19674 );
and \U$19299 ( \19676 , RIc225a80_59, \1391 );
not \U$19300 ( \19677 , RIc225a80_59);
not \U$19301 ( \19678 , \1391 );
and \U$19302 ( \19679 , \19677 , \19678 );
nor \U$19303 ( \19680 , \19676 , \19679 );
nand \U$19304 ( \19681 , \19680 , \15164 );
nand \U$19305 ( \19682 , \19675 , \19681 );
not \U$19306 ( \19683 , \19682 );
not \U$19307 ( \19684 , \9110 );
not \U$19308 ( \19685 , RIc226200_43);
not \U$19309 ( \19686 , \2894 );
or \U$19310 ( \19687 , \19685 , \19686 );
not \U$19311 ( \19688 , \12989 );
nand \U$19312 ( \19689 , \19688 , \9117 );
nand \U$19313 ( \19690 , \19687 , \19689 );
not \U$19314 ( \19691 , \19690 );
or \U$19315 ( \19692 , \19684 , \19691 );
nand \U$19316 ( \19693 , \18922 , \9129 );
nand \U$19317 ( \19694 , \19692 , \19693 );
not \U$19318 ( \19695 , \19694 );
or \U$19319 ( \19696 , \19683 , \19695 );
or \U$19320 ( \19697 , \19694 , \19682 );
not \U$19321 ( \19698 , \9690 );
not \U$19322 ( \19699 , RIc2262f0_41);
not \U$19323 ( \19700 , \12977 );
or \U$19324 ( \19701 , \19699 , \19700 );
nand \U$19325 ( \19702 , \11844 , \9822 );
nand \U$19326 ( \19703 , \19701 , \19702 );
not \U$19327 ( \19704 , \19703 );
or \U$19328 ( \19705 , \19698 , \19704 );
nand \U$19329 ( \19706 , \18934 , \9816 );
nand \U$19330 ( \19707 , \19705 , \19706 );
nand \U$19331 ( \19708 , \19697 , \19707 );
nand \U$19332 ( \19709 , \19696 , \19708 );
and \U$19333 ( \19710 , \19672 , \19709 );
nor \U$19334 ( \19711 , \19669 , \19671 );
nor \U$19335 ( \19712 , \19710 , \19711 );
not \U$19336 ( \19713 , \19712 );
or \U$19337 ( \19714 , \19664 , \19713 );
not \U$19338 ( \19715 , \1120 );
not \U$19339 ( \19716 , \18703 );
or \U$19340 ( \19717 , \19715 , \19716 );
not \U$19341 ( \19718 , \15443 );
not \U$19342 ( \19719 , \1139 );
and \U$19343 ( \19720 , \19718 , \19719 );
buf \U$19344 ( \19721 , \15443 );
and \U$19345 ( \19722 , \19721 , \1139 );
nor \U$19346 ( \19723 , \19720 , \19722 );
not \U$19347 ( \19724 , \19723 );
nand \U$19348 ( \19725 , \19724 , \1118 );
nand \U$19349 ( \19726 , \19717 , \19725 );
and \U$19350 ( \19727 , \18367 , \1081 );
or \U$19351 ( \19728 , \18377 , \955 );
not \U$19352 ( \19729 , \16256 );
not \U$19353 ( \19730 , \946 );
and \U$19354 ( \19731 , \19729 , \19730 );
and \U$19355 ( \19732 , \16482 , \946 );
nor \U$19356 ( \19733 , \19731 , \19732 );
not \U$19357 ( \19734 , \19733 );
nand \U$19358 ( \19735 , \19734 , \950 );
nand \U$19359 ( \19736 , \19728 , \19735 );
xor \U$19360 ( \19737 , \19727 , \19736 );
not \U$19361 ( \19738 , \12845 );
not \U$19362 ( \19739 , \1139 );
and \U$19363 ( \19740 , \19738 , \19739 );
and \U$19364 ( \19741 , \12844 , \940 );
nor \U$19365 ( \19742 , \19740 , \19741 );
or \U$19366 ( \19743 , \19742 , \1117 );
or \U$19367 ( \19744 , \19723 , \1119 );
nand \U$19368 ( \19745 , \19743 , \19744 );
and \U$19369 ( \19746 , \19737 , \19745 );
and \U$19370 ( \19747 , \19727 , \19736 );
or \U$19371 ( \19748 , \19746 , \19747 );
xor \U$19372 ( \19749 , \19726 , \19748 );
not \U$19373 ( \19750 , \1682 );
not \U$19374 ( \19751 , \18197 );
or \U$19375 ( \19752 , \19750 , \19751 );
not \U$19376 ( \19753 , RIc227010_13);
not \U$19377 ( \19754 , \10263 );
or \U$19378 ( \19755 , \19753 , \19754 );
nand \U$19379 ( \19756 , \16998 , \3841 );
nand \U$19380 ( \19757 , \19755 , \19756 );
nand \U$19381 ( \19758 , \19757 , \1678 );
nand \U$19382 ( \19759 , \19752 , \19758 );
and \U$19383 ( \19760 , \19749 , \19759 );
and \U$19384 ( \19761 , \19726 , \19748 );
or \U$19385 ( \19762 , \19760 , \19761 );
not \U$19386 ( \19763 , \19762 );
not \U$19387 ( \19764 , \1311 );
not \U$19388 ( \19765 , \18213 );
or \U$19389 ( \19766 , \19764 , \19765 );
not \U$19390 ( \19767 , RIc227100_11);
not \U$19391 ( \19768 , \10360 );
or \U$19392 ( \19769 , \19767 , \19768 );
nand \U$19393 ( \19770 , \10086 , \1685 );
nand \U$19394 ( \19771 , \19769 , \19770 );
nand \U$19395 ( \19772 , \19771 , \1306 );
nand \U$19396 ( \19773 , \19766 , \19772 );
not \U$19397 ( \19774 , \2320 );
not \U$19398 ( \19775 , RIc226f20_15);
not \U$19399 ( \19776 , \11488 );
or \U$19400 ( \19777 , \19775 , \19776 );
nand \U$19401 ( \19778 , \17014 , \2351 );
nand \U$19402 ( \19779 , \19777 , \19778 );
not \U$19403 ( \19780 , \19779 );
or \U$19404 ( \19781 , \19774 , \19780 );
nand \U$19405 ( \19782 , \18474 , \2358 );
nand \U$19406 ( \19783 , \19781 , \19782 );
or \U$19407 ( \19784 , \19773 , \19783 );
not \U$19408 ( \19785 , \1945 );
not \U$19409 ( \19786 , RIc226e30_17);
not \U$19410 ( \19787 , \9073 );
or \U$19411 ( \19788 , \19786 , \19787 );
buf \U$19412 ( \19789 , \10652 );
not \U$19413 ( \19790 , \19789 );
nand \U$19414 ( \19791 , \19790 , \1935 );
nand \U$19415 ( \19792 , \19788 , \19791 );
not \U$19416 ( \19793 , \19792 );
or \U$19417 ( \19794 , \19785 , \19793 );
nand \U$19418 ( \19795 , \18445 , \1963 );
nand \U$19419 ( \19796 , \19794 , \19795 );
and \U$19420 ( \19797 , \19784 , \19796 );
and \U$19421 ( \19798 , \19783 , \19773 );
nor \U$19422 ( \19799 , \19797 , \19798 );
nand \U$19423 ( \19800 , \19763 , \19799 );
not \U$19424 ( \19801 , \19800 );
or \U$19425 ( \19802 , RIc227358_6, RIc2272e0_7);
nand \U$19426 ( \19803 , \19802 , \18367 );
and \U$19427 ( \19804 , RIc227358_6, RIc2272e0_7);
nor \U$19428 ( \19805 , \19804 , \956 );
and \U$19429 ( \19806 , \19803 , \19805 );
or \U$19430 ( \19807 , \16248 , \946 );
or \U$19431 ( \19808 , \18366 , RIc2273d0_5);
nand \U$19432 ( \19809 , \19807 , \19808 );
not \U$19433 ( \19810 , \19809 );
not \U$19434 ( \19811 , \950 );
or \U$19435 ( \19812 , \19810 , \19811 );
or \U$19436 ( \19813 , \19733 , \955 );
nand \U$19437 ( \19814 , \19812 , \19813 );
and \U$19438 ( \19815 , \19806 , \19814 );
not \U$19439 ( \19816 , \1363 );
not \U$19440 ( \19817 , \1342 );
not \U$19441 ( \19818 , \12755 );
or \U$19442 ( \19819 , \19817 , \19818 );
nand \U$19443 ( \19820 , \13198 , RIc2271f0_9);
nand \U$19444 ( \19821 , \19819 , \19820 );
not \U$19445 ( \19822 , \19821 );
or \U$19446 ( \19823 , \19816 , \19822 );
nand \U$19447 ( \19824 , \18394 , \1339 );
nand \U$19448 ( \19825 , \19823 , \19824 );
xor \U$19449 ( \19826 , \19815 , \19825 );
not \U$19450 ( \19827 , \19771 );
not \U$19451 ( \19828 , \1310 );
or \U$19452 ( \19829 , \19827 , \19828 );
not \U$19453 ( \19830 , RIc227100_11);
not \U$19454 ( \19831 , \10369 );
or \U$19455 ( \19832 , \19830 , \19831 );
nand \U$19456 ( \19833 , \10197 , \1685 );
nand \U$19457 ( \19834 , \19832 , \19833 );
nand \U$19458 ( \19835 , \19834 , \1306 );
nand \U$19459 ( \19836 , \19829 , \19835 );
and \U$19460 ( \19837 , \19826 , \19836 );
and \U$19461 ( \19838 , \19815 , \19825 );
or \U$19462 ( \19839 , \19837 , \19838 );
not \U$19463 ( \19840 , \2086 );
not \U$19464 ( \19841 , \18425 );
or \U$19465 ( \19842 , \19840 , \19841 );
not \U$19466 ( \19843 , \15645 );
not \U$19467 ( \19844 , \10900 );
and \U$19468 ( \19845 , \19843 , \19844 );
not \U$19469 ( \19846 , RIc226890_29);
and \U$19470 ( \19847 , \10126 , \19846 );
nor \U$19471 ( \19848 , \19845 , \19847 );
or \U$19472 ( \19849 , \19848 , \3930 );
nand \U$19473 ( \19850 , \19842 , \19849 );
xor \U$19474 ( \19851 , \19839 , \19850 );
not \U$19475 ( \19852 , \2710 );
not \U$19476 ( \19853 , \18461 );
or \U$19477 ( \19854 , \19852 , \19853 );
not \U$19478 ( \19855 , \11182 );
not \U$19479 ( \19856 , RIc2267a0_31);
not \U$19480 ( \19857 , \5664 );
or \U$19481 ( \19858 , \19856 , \19857 );
not \U$19482 ( \19859 , \10161 );
nand \U$19483 ( \19860 , \19859 , \2072 );
nand \U$19484 ( \19861 , \19858 , \19860 );
nand \U$19485 ( \19862 , \19855 , \19861 );
nand \U$19486 ( \19863 , \19854 , \19862 );
and \U$19487 ( \19864 , \19851 , \19863 );
and \U$19488 ( \19865 , \19839 , \19850 );
or \U$19489 ( \19866 , \19864 , \19865 );
not \U$19490 ( \19867 , \19866 );
or \U$19491 ( \19868 , \19801 , \19867 );
not \U$19492 ( \19869 , \19799 );
nand \U$19493 ( \19870 , \19869 , \19762 );
nand \U$19494 ( \19871 , \19868 , \19870 );
nand \U$19495 ( \19872 , \19714 , \19871 );
not \U$19496 ( \19873 , \19663 );
not \U$19497 ( \19874 , \19712 );
nand \U$19498 ( \19875 , \19873 , \19874 );
nand \U$19499 ( \19876 , \19872 , \19875 );
nand \U$19500 ( \19877 , \19588 , \19876 );
nand \U$19501 ( \19878 , \19583 , \19877 );
xor \U$19502 ( \19879 , \19111 , \19113 );
xor \U$19503 ( \19880 , \19879 , \19148 );
xor \U$19504 ( \19881 , \19878 , \19880 );
not \U$19505 ( \19882 , \18979 );
and \U$19506 ( \19883 , \19109 , \19882 );
not \U$19507 ( \19884 , \19109 );
and \U$19508 ( \19885 , \19884 , \18979 );
nor \U$19509 ( \19886 , \19883 , \19885 );
not \U$19510 ( \19887 , \19091 );
and \U$19511 ( \19888 , \19886 , \19887 );
not \U$19512 ( \19889 , \19886 );
and \U$19513 ( \19890 , \19889 , \19091 );
nor \U$19514 ( \19891 , \19888 , \19890 );
not \U$19515 ( \19892 , \19891 );
not \U$19516 ( \19893 , \19892 );
not \U$19517 ( \19894 , \19049 );
and \U$19518 ( \19895 , \19035 , \19894 );
not \U$19519 ( \19896 , \19035 );
and \U$19520 ( \19897 , \19896 , \19049 );
nor \U$19521 ( \19898 , \19895 , \19897 );
and \U$19522 ( \19899 , \19898 , \19025 );
not \U$19523 ( \19900 , \19898 );
not \U$19524 ( \19901 , \19025 );
and \U$19525 ( \19902 , \19900 , \19901 );
nor \U$19526 ( \19903 , \19899 , \19902 );
not \U$19527 ( \19904 , \19903 );
xor \U$19528 ( \19905 , \18938 , \18927 );
xor \U$19529 ( \19906 , \19905 , \18916 );
not \U$19530 ( \19907 , \19906 );
or \U$19531 ( \19908 , \19904 , \19907 );
xor \U$19532 ( \19909 , \18972 , \18967 );
xnor \U$19533 ( \19910 , \19909 , \18956 );
not \U$19534 ( \19911 , \19910 );
nand \U$19535 ( \19912 , \19908 , \19911 );
not \U$19536 ( \19913 , \19906 );
not \U$19537 ( \19914 , \19903 );
nand \U$19538 ( \19915 , \19913 , \19914 );
nand \U$19539 ( \19916 , \19912 , \19915 );
xor \U$19540 ( \19917 , \19088 , \19051 );
xor \U$19541 ( \19918 , \19917 , \19014 );
xor \U$19542 ( \19919 , \19916 , \19918 );
xor \U$19543 ( \19920 , \19726 , \19748 );
xor \U$19544 ( \19921 , \19920 , \19759 );
not \U$19545 ( \19922 , \4383 );
not \U$19546 ( \19923 , \19057 );
or \U$19547 ( \19924 , \19922 , \19923 );
not \U$19548 ( \19925 , RIc2265c0_35);
not \U$19549 ( \19926 , \3641 );
not \U$19550 ( \19927 , \19926 );
or \U$19551 ( \19928 , \19925 , \19927 );
not \U$19552 ( \19929 , \4049 );
nand \U$19553 ( \19930 , \19929 , \3620 );
nand \U$19554 ( \19931 , \19928 , \19930 );
nand \U$19555 ( \19932 , \19931 , \5741 );
nand \U$19556 ( \19933 , \19924 , \19932 );
xor \U$19557 ( \19934 , \19921 , \19933 );
xor \U$19558 ( \19935 , \19727 , \19736 );
xor \U$19559 ( \19936 , \19935 , \19745 );
not \U$19560 ( \19937 , \2320 );
not \U$19561 ( \19938 , RIc226f20_15);
not \U$19562 ( \19939 , \9276 );
or \U$19563 ( \19940 , \19938 , \19939 );
nand \U$19564 ( \19941 , \9275 , \2301 );
nand \U$19565 ( \19942 , \19940 , \19941 );
not \U$19566 ( \19943 , \19942 );
or \U$19567 ( \19944 , \19937 , \19943 );
nand \U$19568 ( \19945 , \19779 , \2358 );
nand \U$19569 ( \19946 , \19944 , \19945 );
xor \U$19570 ( \19947 , \19936 , \19946 );
not \U$19571 ( \19948 , \1963 );
not \U$19572 ( \19949 , \19792 );
or \U$19573 ( \19950 , \19948 , \19949 );
not \U$19574 ( \19951 , RIc226e30_17);
not \U$19575 ( \19952 , \10111 );
or \U$19576 ( \19953 , \19951 , \19952 );
nand \U$19577 ( \19954 , \10110 , \1952 );
nand \U$19578 ( \19955 , \19953 , \19954 );
nand \U$19579 ( \19956 , \19955 , \1945 );
nand \U$19580 ( \19957 , \19950 , \19956 );
and \U$19581 ( \19958 , \19947 , \19957 );
and \U$19582 ( \19959 , \19936 , \19946 );
or \U$19583 ( \19960 , \19958 , \19959 );
and \U$19584 ( \19961 , \19934 , \19960 );
and \U$19585 ( \19962 , \19921 , \19933 );
or \U$19586 ( \19963 , \19961 , \19962 );
xor \U$19587 ( \19964 , \18990 , \19001 );
xor \U$19588 ( \19965 , \19964 , \19011 );
xor \U$19589 ( \19966 , \19963 , \19965 );
xor \U$19590 ( \19967 , \19086 , \19074 );
xor \U$19591 ( \19968 , \19967 , \19063 );
and \U$19592 ( \19969 , \19966 , \19968 );
and \U$19593 ( \19970 , \19963 , \19965 );
or \U$19594 ( \19971 , \19969 , \19970 );
and \U$19595 ( \19972 , \19919 , \19971 );
and \U$19596 ( \19973 , \19916 , \19918 );
or \U$19597 ( \19974 , \19972 , \19973 );
not \U$19598 ( \19975 , \19974 );
not \U$19599 ( \19976 , \19975 );
or \U$19600 ( \19977 , \19893 , \19976 );
xor \U$19601 ( \19978 , \19241 , \19243 );
xor \U$19602 ( \19979 , \19978 , \19252 );
nand \U$19603 ( \19980 , \19977 , \19979 );
not \U$19604 ( \19981 , \19892 );
nand \U$19605 ( \19982 , \19981 , \19974 );
nand \U$19606 ( \19983 , \19980 , \19982 );
and \U$19607 ( \19984 , \19881 , \19983 );
and \U$19608 ( \19985 , \19878 , \19880 );
or \U$19609 ( \19986 , \19984 , \19985 );
and \U$19610 ( \19987 , \19498 , \19986 );
and \U$19611 ( \19988 , \19484 , \19496 );
nor \U$19612 ( \19989 , \19987 , \19988 );
nand \U$19613 ( \19990 , \19438 , \19989 );
xor \U$19614 ( \19991 , \19272 , \19284 );
xnor \U$19615 ( \19992 , \19991 , \19419 );
and \U$19616 ( \19993 , \19990 , \19992 );
nor \U$19617 ( \19994 , \19989 , \19438 );
nor \U$19618 ( \19995 , \19993 , \19994 );
nor \U$19619 ( \19996 , \19435 , \19995 );
not \U$19620 ( \19997 , \19996 );
xor \U$19621 ( \19998 , \17677 , \18815 );
xor \U$19622 ( \19999 , \19998 , \18854 );
xor \U$19623 ( \20000 , \18892 , \19423 );
and \U$19624 ( \20001 , \20000 , \19434 );
and \U$19625 ( \20002 , \18892 , \19423 );
or \U$19626 ( \20003 , \20001 , \20002 );
nand \U$19627 ( \20004 , \19999 , \20003 );
not \U$19628 ( \20005 , \20004 );
or \U$19629 ( \20006 , \19997 , \20005 );
not \U$19630 ( \20007 , \19999 );
not \U$19631 ( \20008 , \20003 );
nand \U$19632 ( \20009 , \20007 , \20008 );
nand \U$19633 ( \20010 , \20006 , \20009 );
not \U$19634 ( \20011 , \20010 );
or \U$19635 ( \20012 , \18890 , \20011 );
or \U$19636 ( \20013 , \18888 , \18857 );
nand \U$19637 ( \20014 , \20012 , \20013 );
xor \U$19638 ( \20015 , \16864 , \17441 );
xnor \U$19639 ( \20016 , \20015 , \16753 );
not \U$19640 ( \20017 , \18887 );
not \U$19641 ( \20018 , \18864 );
nand \U$19642 ( \20019 , \20017 , \20018 );
and \U$19643 ( \20020 , \20019 , \18874 );
nor \U$19644 ( \20021 , \20017 , \20018 );
nor \U$19645 ( \20022 , \20020 , \20021 );
nand \U$19646 ( \20023 , \20016 , \20022 );
buf \U$19647 ( \20024 , \20023 );
and \U$19648 ( \20025 , \20014 , \20024 );
nor \U$19649 ( \20026 , \20016 , \20022 );
nor \U$19650 ( \20027 , \20025 , \20026 );
and \U$19651 ( \20028 , \19992 , \19438 );
not \U$19652 ( \20029 , \19992 );
not \U$19653 ( \20030 , \19438 );
and \U$19654 ( \20031 , \20029 , \20030 );
nor \U$19655 ( \20032 , \20028 , \20031 );
buf \U$19656 ( \20033 , \19989 );
not \U$19657 ( \20034 , \20033 );
and \U$19658 ( \20035 , \20032 , \20034 );
not \U$19659 ( \20036 , \20032 );
and \U$19660 ( \20037 , \20036 , \20033 );
nor \U$19661 ( \20038 , \20035 , \20037 );
xor \U$19662 ( \20039 , \19292 , \19413 );
xor \U$19663 ( \20040 , \20039 , \19416 );
not \U$19664 ( \20041 , \20040 );
buf \U$19665 ( \20042 , \19484 );
not \U$19666 ( \20043 , \20042 );
not \U$19667 ( \20044 , \19495 );
not \U$19668 ( \20045 , \19986 );
and \U$19669 ( \20046 , \20044 , \20045 );
and \U$19670 ( \20047 , \19495 , \19986 );
nor \U$19671 ( \20048 , \20046 , \20047 );
not \U$19672 ( \20049 , \20048 );
or \U$19673 ( \20050 , \20043 , \20049 );
or \U$19674 ( \20051 , \20048 , \20042 );
nand \U$19675 ( \20052 , \20050 , \20051 );
not \U$19676 ( \20053 , \20052 );
nand \U$19677 ( \20054 , \20041 , \20053 );
not \U$19678 ( \20055 , \19876 );
not \U$19679 ( \20056 , \19586 );
or \U$19680 ( \20057 , \20055 , \20056 );
nand \U$19681 ( \20058 , \19872 , \19875 , \19581 );
nand \U$19682 ( \20059 , \20057 , \20058 );
and \U$19683 ( \20060 , \20059 , \19584 );
not \U$19684 ( \20061 , \20059 );
and \U$19685 ( \20062 , \20061 , \19500 );
nor \U$19686 ( \20063 , \20060 , \20062 );
not \U$19687 ( \20064 , \19390 );
not \U$19688 ( \20065 , \19388 );
not \U$19689 ( \20066 , \20065 );
or \U$19690 ( \20067 , \20064 , \20066 );
nand \U$19691 ( \20068 , \19308 , \19388 );
nand \U$19692 ( \20069 , \20067 , \20068 );
and \U$19693 ( \20070 , \20069 , \19349 );
not \U$19694 ( \20071 , \20069 );
and \U$19695 ( \20072 , \20071 , \19348 );
nor \U$19696 ( \20073 , \20070 , \20072 );
not \U$19697 ( \20074 , \20073 );
not \U$19698 ( \20075 , \20074 );
not \U$19699 ( \20076 , \11965 );
and \U$19700 ( \20077 , RIc225b70_57, \9115 );
not \U$19701 ( \20078 , RIc225b70_57);
and \U$19702 ( \20079 , \20078 , \3043 );
or \U$19703 ( \20080 , \20077 , \20079 );
not \U$19704 ( \20081 , \20080 );
or \U$19705 ( \20082 , \20076 , \20081 );
nand \U$19706 ( \20083 , \19521 , \11974 );
nand \U$19707 ( \20084 , \20082 , \20083 );
not \U$19708 ( \20085 , \15729 );
not \U$19709 ( \20086 , \19558 );
or \U$19710 ( \20087 , \20085 , \20086 );
not \U$19711 ( \20088 , RIc225990_61);
not \U$19712 ( \20089 , \1222 );
or \U$19713 ( \20090 , \20088 , \20089 );
nand \U$19714 ( \20091 , \10428 , \12806 );
nand \U$19715 ( \20092 , \20090 , \20091 );
nand \U$19716 ( \20093 , \20092 , \15719 );
nand \U$19717 ( \20094 , \20087 , \20093 );
xor \U$19718 ( \20095 , \20084 , \20094 );
not \U$19719 ( \20096 , \10001 );
not \U$19720 ( \20097 , RIc226020_47);
not \U$19721 ( \20098 , \2586 );
or \U$19722 ( \20099 , \20097 , \20098 );
or \U$19723 ( \20100 , RIc226020_47, \2592 );
nand \U$19724 ( \20101 , \20099 , \20100 );
not \U$19725 ( \20102 , \20101 );
or \U$19726 ( \20103 , \20096 , \20102 );
nand \U$19727 ( \20104 , \19532 , \9619 );
nand \U$19728 ( \20105 , \20103 , \20104 );
and \U$19729 ( \20106 , \20095 , \20105 );
and \U$19730 ( \20107 , \20084 , \20094 );
or \U$19731 ( \20108 , \20106 , \20107 );
not \U$19732 ( \20109 , \20108 );
not \U$19733 ( \20110 , \9934 );
not \U$19734 ( \20111 , RIc226110_45);
not \U$19735 ( \20112 , \2476 );
or \U$19736 ( \20113 , \20111 , \20112 );
not \U$19737 ( \20114 , \2476 );
nand \U$19738 ( \20115 , \20114 , \10429 );
nand \U$19739 ( \20116 , \20113 , \20115 );
not \U$19740 ( \20117 , \20116 );
or \U$19741 ( \20118 , \20110 , \20117 );
nand \U$19742 ( \20119 , \19637 , \9398 );
nand \U$19743 ( \20120 , \20118 , \20119 );
not \U$19744 ( \20121 , \20120 );
not \U$19745 ( \20122 , \9129 );
not \U$19746 ( \20123 , \19690 );
or \U$19747 ( \20124 , \20122 , \20123 );
not \U$19748 ( \20125 , RIc226200_43);
not \U$19749 ( \20126 , \2670 );
or \U$19750 ( \20127 , \20125 , \20126 );
nand \U$19751 ( \20128 , \2720 , \9117 );
nand \U$19752 ( \20129 , \20127 , \20128 );
nand \U$19753 ( \20130 , \20129 , \9110 );
nand \U$19754 ( \20131 , \20124 , \20130 );
not \U$19755 ( \20132 , \20131 );
or \U$19756 ( \20133 , \20121 , \20132 );
or \U$19757 ( \20134 , \20131 , \20120 );
not \U$19758 ( \20135 , \11118 );
not \U$19759 ( \20136 , RIc225c60_55);
not \U$19760 ( \20137 , \9700 );
or \U$19761 ( \20138 , \20136 , \20137 );
nand \U$19762 ( \20139 , \2353 , \11108 );
nand \U$19763 ( \20140 , \20138 , \20139 );
not \U$19764 ( \20141 , \20140 );
or \U$19765 ( \20142 , \20135 , \20141 );
nand \U$19766 ( \20143 , \19649 , \13025 );
nand \U$19767 ( \20144 , \20142 , \20143 );
nand \U$19768 ( \20145 , \20134 , \20144 );
nand \U$19769 ( \20146 , \20133 , \20145 );
not \U$19770 ( \20147 , \20146 );
nand \U$19771 ( \20148 , \20109 , \20147 );
not \U$19772 ( \20149 , \19625 );
not \U$19773 ( \20150 , \20149 );
not \U$19774 ( \20151 , \16882 );
and \U$19775 ( \20152 , \20150 , \20151 );
not \U$19776 ( \20153 , \16880 );
not \U$19777 ( \20154 , \2119 );
or \U$19778 ( \20155 , \20153 , \20154 );
not \U$19779 ( \20156 , \1020 );
nand \U$19780 ( \20157 , \20156 , RIc2258a0_63);
nand \U$19781 ( \20158 , \20155 , \20157 );
buf \U$19782 ( \20159 , \16891 );
and \U$19783 ( \20160 , \20158 , \20159 );
nor \U$19784 ( \20161 , \20152 , \20160 );
not \U$19785 ( \20162 , \20161 );
not \U$19786 ( \20163 , \20162 );
and \U$19787 ( \20164 , \19595 , \11577 );
not \U$19788 ( \20165 , RIc225d50_53);
not \U$19789 ( \20166 , \13914 );
or \U$19790 ( \20167 , \20165 , \20166 );
nand \U$19791 ( \20168 , \4457 , \11391 );
nand \U$19792 ( \20169 , \20167 , \20168 );
and \U$19793 ( \20170 , \20169 , \8777 );
nor \U$19794 ( \20171 , \20164 , \20170 );
not \U$19795 ( \20172 , \20171 );
not \U$19796 ( \20173 , \20172 );
or \U$19797 ( \20174 , \20163 , \20173 );
not \U$19798 ( \20175 , \20161 );
not \U$19799 ( \20176 , \20171 );
or \U$19800 ( \20177 , \20175 , \20176 );
not \U$19801 ( \20178 , \9705 );
not \U$19802 ( \20179 , \19703 );
or \U$19803 ( \20180 , \20178 , \20179 );
and \U$19804 ( \20181 , RIc2262f0_41, \11068 );
not \U$19805 ( \20182 , RIc2262f0_41);
not \U$19806 ( \20183 , \11068 );
and \U$19807 ( \20184 , \20182 , \20183 );
or \U$19808 ( \20185 , \20181 , \20184 );
nand \U$19809 ( \20186 , \20185 , \9690 );
nand \U$19810 ( \20187 , \20180 , \20186 );
nand \U$19811 ( \20188 , \20177 , \20187 );
nand \U$19812 ( \20189 , \20174 , \20188 );
and \U$19813 ( \20190 , \20148 , \20189 );
not \U$19814 ( \20191 , \20108 );
nor \U$19815 ( \20192 , \20191 , \20147 );
nor \U$19816 ( \20193 , \20190 , \20192 );
not \U$19817 ( \20194 , \20193 );
not \U$19818 ( \20195 , \20194 );
or \U$19819 ( \20196 , \20075 , \20195 );
not \U$19820 ( \20197 , \20193 );
not \U$19821 ( \20198 , \20073 );
or \U$19822 ( \20199 , \20197 , \20198 );
xor \U$19823 ( \20200 , \19319 , \19346 );
xnor \U$19824 ( \20201 , \20200 , \19329 );
not \U$19825 ( \20202 , \20201 );
not \U$19826 ( \20203 , \9552 );
not \U$19827 ( \20204 , \19569 );
or \U$19828 ( \20205 , \20203 , \20204 );
not \U$19829 ( \20206 , RIc225f30_49);
not \U$19830 ( \20207 , \3839 );
or \U$19831 ( \20208 , \20206 , \20207 );
nand \U$19832 ( \20209 , \15287 , \11289 );
nand \U$19833 ( \20210 , \20208 , \20209 );
nand \U$19834 ( \20211 , \20210 , \9534 );
nand \U$19835 ( \20212 , \20205 , \20211 );
not \U$19836 ( \20213 , \20212 );
not \U$19837 ( \20214 , \2195 );
not \U$19838 ( \20215 , RIc226a70_25);
buf \U$19839 ( \20216 , \8829 );
not \U$19840 ( \20217 , \20216 );
not \U$19841 ( \20218 , \20217 );
or \U$19842 ( \20219 , \20215 , \20218 );
nand \U$19843 ( \20220 , \20216 , \1905 );
nand \U$19844 ( \20221 , \20219 , \20220 );
not \U$19845 ( \20222 , \20221 );
or \U$19846 ( \20223 , \20214 , \20222 );
nand \U$19847 ( \20224 , \19356 , \2173 );
nand \U$19848 ( \20225 , \20223 , \20224 );
not \U$19849 ( \20226 , \20225 );
not \U$19850 ( \20227 , \2392 );
not \U$19851 ( \20228 , RIc226c50_21);
not \U$19852 ( \20229 , \8910 );
or \U$19853 ( \20230 , \20228 , \20229 );
nand \U$19854 ( \20231 , \9790 , \3204 );
nand \U$19855 ( \20232 , \20230 , \20231 );
not \U$19856 ( \20233 , \20232 );
or \U$19857 ( \20234 , \20227 , \20233 );
nand \U$19858 ( \20235 , \19326 , \2367 );
nand \U$19859 ( \20236 , \20234 , \20235 );
not \U$19860 ( \20237 , \20236 );
nand \U$19861 ( \20238 , \20226 , \20237 );
not \U$19862 ( \20239 , \20238 );
or \U$19863 ( \20240 , \20213 , \20239 );
nand \U$19864 ( \20241 , \20236 , \20225 );
nand \U$19865 ( \20242 , \20240 , \20241 );
not \U$19866 ( \20243 , \20242 );
not \U$19867 ( \20244 , \20243 );
or \U$19868 ( \20245 , \20202 , \20244 );
xor \U$19869 ( \20246 , \19839 , \19850 );
xor \U$19870 ( \20247 , \20246 , \19863 );
nand \U$19871 ( \20248 , \20245 , \20247 );
not \U$19872 ( \20249 , \20201 );
nand \U$19873 ( \20250 , \20249 , \20242 );
nand \U$19874 ( \20251 , \20248 , \20250 );
nand \U$19875 ( \20252 , \20199 , \20251 );
nand \U$19876 ( \20253 , \20196 , \20252 );
not \U$19877 ( \20254 , \20253 );
not \U$19878 ( \20255 , \19866 );
not \U$19879 ( \20256 , \19799 );
not \U$19880 ( \20257 , \19762 );
and \U$19881 ( \20258 , \20256 , \20257 );
and \U$19882 ( \20259 , \19799 , \19762 );
nor \U$19883 ( \20260 , \20258 , \20259 );
not \U$19884 ( \20261 , \20260 );
and \U$19885 ( \20262 , \20255 , \20261 );
and \U$19886 ( \20263 , \19866 , \20260 );
nor \U$19887 ( \20264 , \20262 , \20263 );
not \U$19888 ( \20265 , \20264 );
not \U$19889 ( \20266 , \19613 );
not \U$19890 ( \20267 , \20266 );
not \U$19891 ( \20268 , \6308 );
and \U$19892 ( \20269 , \20267 , \20268 );
not \U$19893 ( \20270 , RIc2263e0_39);
not \U$19894 ( \20271 , \10532 );
or \U$19895 ( \20272 , \20270 , \20271 );
nand \U$19896 ( \20273 , \4500 , \5498 );
nand \U$19897 ( \20274 , \20272 , \20273 );
and \U$19898 ( \20275 , \20274 , \6689 );
nor \U$19899 ( \20276 , \20269 , \20275 );
not \U$19900 ( \20277 , \20276 );
not \U$19901 ( \20278 , \20277 );
not \U$19902 ( \20279 , RIc2264d0_37);
not \U$19903 ( \20280 , \12493 );
or \U$19904 ( \20281 , \20279 , \20280 );
nand \U$19905 ( \20282 , \2980 , \4371 );
nand \U$19906 ( \20283 , \20281 , \20282 );
and \U$19907 ( \20284 , \20283 , \5509 );
and \U$19908 ( \20285 , \19606 , \5519 );
nor \U$19909 ( \20286 , \20284 , \20285 );
not \U$19910 ( \20287 , \20286 );
not \U$19911 ( \20288 , \20287 );
or \U$19912 ( \20289 , \20278 , \20288 );
not \U$19913 ( \20290 , \20276 );
not \U$19914 ( \20291 , \20286 );
or \U$19915 ( \20292 , \20290 , \20291 );
xor \U$19916 ( \20293 , \19815 , \19825 );
xor \U$19917 ( \20294 , \20293 , \19836 );
nand \U$19918 ( \20295 , \20292 , \20294 );
nand \U$19919 ( \20296 , \20289 , \20295 );
xor \U$19920 ( \20297 , \19773 , \19783 );
xor \U$19921 ( \20298 , \20297 , \19796 );
not \U$19922 ( \20299 , \20298 );
not \U$19923 ( \20300 , \19386 );
not \U$19924 ( \20301 , \19373 );
or \U$19925 ( \20302 , \20300 , \20301 );
or \U$19926 ( \20303 , \19373 , \19386 );
nand \U$19927 ( \20304 , \20302 , \20303 );
and \U$19928 ( \20305 , \20304 , \19359 );
not \U$19929 ( \20306 , \20304 );
and \U$19930 ( \20307 , \20306 , \19360 );
nor \U$19931 ( \20308 , \20305 , \20307 );
nand \U$19932 ( \20309 , \20299 , \20308 );
and \U$19933 ( \20310 , \20296 , \20309 );
not \U$19934 ( \20311 , \20298 );
nor \U$19935 ( \20312 , \20311 , \20308 );
nor \U$19936 ( \20313 , \20310 , \20312 );
not \U$19937 ( \20314 , \20313 );
or \U$19938 ( \20315 , \20265 , \20314 );
not \U$19939 ( \20316 , \1682 );
not \U$19940 ( \20317 , \19757 );
or \U$19941 ( \20318 , \20316 , \20317 );
not \U$19942 ( \20319 , RIc227010_13);
not \U$19943 ( \20320 , \13442 );
or \U$19944 ( \20321 , \20319 , \20320 );
nand \U$19945 ( \20322 , \9320 , \3841 );
nand \U$19946 ( \20323 , \20321 , \20322 );
nand \U$19947 ( \20324 , \20323 , \1678 );
nand \U$19948 ( \20325 , \20318 , \20324 );
not \U$19949 ( \20326 , \2534 );
not \U$19950 ( \20327 , \19315 );
or \U$19951 ( \20328 , \20326 , \20327 );
and \U$19952 ( \20329 , RIc226d40_19, \13465 );
not \U$19953 ( \20330 , RIc226d40_19);
and \U$19954 ( \20331 , \20330 , \9051 );
or \U$19955 ( \20332 , \20329 , \20331 );
nand \U$19956 ( \20333 , \20332 , \2518 );
nand \U$19957 ( \20334 , \20328 , \20333 );
xor \U$19958 ( \20335 , \20325 , \20334 );
not \U$19959 ( \20336 , \4383 );
not \U$19960 ( \20337 , \19931 );
or \U$19961 ( \20338 , \20336 , \20337 );
not \U$19962 ( \20339 , RIc2265c0_35);
not \U$19963 ( \20340 , \4122 );
or \U$19964 ( \20341 , \20339 , \20340 );
nand \U$19965 ( \20342 , \5569 , \16314 );
nand \U$19966 ( \20343 , \20341 , \20342 );
nand \U$19967 ( \20344 , \20343 , \4381 );
nand \U$19968 ( \20345 , \20338 , \20344 );
and \U$19969 ( \20346 , \20335 , \20345 );
and \U$19970 ( \20347 , \20325 , \20334 );
or \U$19971 ( \20348 , \20346 , \20347 );
not \U$19972 ( \20349 , \20348 );
not \U$19973 ( \20350 , \5215 );
not \U$19974 ( \20351 , \5179 );
and \U$19975 ( \20352 , \20350 , \20351 );
and \U$19976 ( \20353 , \13515 , \2692 );
nor \U$19977 ( \20354 , \20352 , \20353 );
not \U$19978 ( \20355 , \20354 );
not \U$19979 ( \20356 , \5185 );
and \U$19980 ( \20357 , \20355 , \20356 );
and \U$19981 ( \20358 , \19341 , \3631 );
nor \U$19982 ( \20359 , \20357 , \20358 );
not \U$19983 ( \20360 , \19365 );
not \U$19984 ( \20361 , \20360 );
not \U$19985 ( \20362 , \7038 );
and \U$19986 ( \20363 , \20361 , \20362 );
not \U$19987 ( \20364 , RIc226b60_23);
not \U$19988 ( \20365 , \11565 );
or \U$19989 ( \20366 , \20364 , \20365 );
not \U$19990 ( \20367 , \8951 );
not \U$19991 ( \20368 , \20367 );
nand \U$19992 ( \20369 , \20368 , \1911 );
nand \U$19993 ( \20370 , \20366 , \20369 );
and \U$19994 ( \20371 , \20370 , \10214 );
nor \U$19995 ( \20372 , \20363 , \20371 );
nand \U$19996 ( \20373 , \20359 , \20372 );
not \U$19997 ( \20374 , \2138 );
not \U$19998 ( \20375 , RIc226980_27);
not \U$19999 ( \20376 , \17579 );
or \U$20000 ( \20377 , \20375 , \20376 );
nand \U$20001 ( \20378 , \16532 , \2133 );
nand \U$20002 ( \20379 , \20377 , \20378 );
not \U$20003 ( \20380 , \20379 );
or \U$20004 ( \20381 , \20374 , \20380 );
nand \U$20005 ( \20382 , \19384 , \2154 );
nand \U$20006 ( \20383 , \20381 , \20382 );
and \U$20007 ( \20384 , \20373 , \20383 );
nor \U$20008 ( \20385 , \20359 , \20372 );
nor \U$20009 ( \20386 , \20384 , \20385 );
nand \U$20010 ( \20387 , \20349 , \20386 );
not \U$20011 ( \20388 , \20387 );
xor \U$20012 ( \20389 , \19806 , \19814 );
not \U$20013 ( \20390 , \19742 );
nand \U$20014 ( \20391 , \20390 , \1120 );
not \U$20015 ( \20392 , \13487 );
not \U$20016 ( \20393 , \20392 );
and \U$20017 ( \20394 , \1139 , \20393 );
not \U$20018 ( \20395 , \1139 );
and \U$20019 ( \20396 , \20395 , \15623 );
nor \U$20020 ( \20397 , \20394 , \20396 );
not \U$20021 ( \20398 , \20397 );
nand \U$20022 ( \20399 , \20398 , \1118 );
nand \U$20023 ( \20400 , \20391 , \20399 );
xor \U$20024 ( \20401 , \20389 , \20400 );
not \U$20025 ( \20402 , \1306 );
not \U$20026 ( \20403 , RIc227100_11);
not \U$20027 ( \20404 , \17625 );
or \U$20028 ( \20405 , \20403 , \20404 );
not \U$20029 ( \20406 , \16492 );
nand \U$20030 ( \20407 , \20406 , \1685 );
nand \U$20031 ( \20408 , \20405 , \20407 );
not \U$20032 ( \20409 , \20408 );
or \U$20033 ( \20410 , \20402 , \20409 );
nand \U$20034 ( \20411 , \19834 , \1311 );
nand \U$20035 ( \20412 , \20410 , \20411 );
and \U$20036 ( \20413 , \20401 , \20412 );
and \U$20037 ( \20414 , \20389 , \20400 );
or \U$20038 ( \20415 , \20413 , \20414 );
not \U$20039 ( \20416 , \2697 );
not \U$20040 ( \20417 , RIc2267a0_31);
not \U$20041 ( \20418 , \17549 );
or \U$20042 ( \20419 , \20417 , \20418 );
nand \U$20043 ( \20420 , \6071 , \3648 );
nand \U$20044 ( \20421 , \20419 , \20420 );
not \U$20045 ( \20422 , \20421 );
or \U$20046 ( \20423 , \20416 , \20422 );
nand \U$20047 ( \20424 , \19861 , \2710 );
nand \U$20048 ( \20425 , \20423 , \20424 );
xor \U$20049 ( \20426 , \20415 , \20425 );
not \U$20050 ( \20427 , \9740 );
not \U$20051 ( \20428 , \19846 );
and \U$20052 ( \20429 , \20427 , \20428 );
and \U$20053 ( \20430 , \6720 , \9144 );
nor \U$20054 ( \20431 , \20429 , \20430 );
not \U$20055 ( \20432 , \20431 );
nand \U$20056 ( \20433 , \20432 , \2078 );
not \U$20057 ( \20434 , \19848 );
nand \U$20058 ( \20435 , \20434 , \9142 );
nand \U$20059 ( \20436 , \20433 , \20435 );
and \U$20060 ( \20437 , \20426 , \20436 );
and \U$20061 ( \20438 , \20415 , \20425 );
or \U$20062 ( \20439 , \20437 , \20438 );
not \U$20063 ( \20440 , \20439 );
or \U$20064 ( \20441 , \20388 , \20440 );
not \U$20065 ( \20442 , \20386 );
nand \U$20066 ( \20443 , \20442 , \20348 );
nand \U$20067 ( \20444 , \20441 , \20443 );
nand \U$20068 ( \20445 , \20315 , \20444 );
not \U$20069 ( \20446 , \20264 );
not \U$20070 ( \20447 , \20313 );
nand \U$20071 ( \20448 , \20446 , \20447 );
nand \U$20072 ( \20449 , \20445 , \20448 );
not \U$20073 ( \20450 , \20449 );
xor \U$20074 ( \20451 , \19302 , \19305 );
xnor \U$20075 ( \20452 , \20451 , \19392 );
nand \U$20076 ( \20453 , \20450 , \20452 );
not \U$20077 ( \20454 , \20453 );
or \U$20078 ( \20455 , \20254 , \20454 );
not \U$20079 ( \20456 , \20452 );
nand \U$20080 ( \20457 , \20456 , \20449 );
nand \U$20081 ( \20458 , \20455 , \20457 );
not \U$20082 ( \20459 , \20458 );
or \U$20083 ( \20460 , \20063 , \20459 );
not \U$20084 ( \20461 , \20459 );
not \U$20085 ( \20462 , \20063 );
or \U$20086 ( \20463 , \20461 , \20462 );
xnor \U$20087 ( \20464 , \19871 , \19663 );
xor \U$20088 ( \20465 , \20464 , \19874 );
not \U$20089 ( \20466 , \20465 );
xor \U$20090 ( \20467 , \19509 , \19507 );
xnor \U$20091 ( \20468 , \20467 , \19578 );
not \U$20092 ( \20469 , \20468 );
not \U$20093 ( \20470 , \20469 );
or \U$20094 ( \20471 , \20466 , \20470 );
or \U$20095 ( \20472 , \20469 , \20465 );
xor \U$20096 ( \20473 , \19669 , \19671 );
xor \U$20097 ( \20474 , \20473 , \19709 );
xor \U$20098 ( \20475 , \19641 , \19653 );
buf \U$20099 ( \20476 , \19629 );
and \U$20100 ( \20477 , \20475 , \20476 );
not \U$20101 ( \20478 , \20475 );
not \U$20102 ( \20479 , \20476 );
and \U$20103 ( \20480 , \20478 , \20479 );
nor \U$20104 ( \20481 , \20477 , \20480 );
buf \U$20105 ( \20482 , \20481 );
not \U$20106 ( \20483 , \20482 );
xor \U$20107 ( \20484 , \19682 , \19694 );
xor \U$20108 ( \20485 , \20484 , \19707 );
not \U$20109 ( \20486 , \20485 );
or \U$20110 ( \20487 , \20483 , \20486 );
or \U$20111 ( \20488 , \20485 , \20482 );
xor \U$20112 ( \20489 , \19553 , \19562 );
xor \U$20113 ( \20490 , \20489 , \19573 );
nand \U$20114 ( \20491 , \20488 , \20490 );
nand \U$20115 ( \20492 , \20487 , \20491 );
xor \U$20116 ( \20493 , \20474 , \20492 );
xor \U$20117 ( \20494 , \19548 , \19512 );
xor \U$20118 ( \20495 , \20494 , \19576 );
and \U$20119 ( \20496 , \20493 , \20495 );
and \U$20120 ( \20497 , \20474 , \20492 );
or \U$20121 ( \20498 , \20496 , \20497 );
nand \U$20122 ( \20499 , \20472 , \20498 );
nand \U$20123 ( \20500 , \20471 , \20499 );
nand \U$20124 ( \20501 , \20463 , \20500 );
nand \U$20125 ( \20502 , \20460 , \20501 );
xor \U$20126 ( \20503 , \19878 , \19880 );
xor \U$20127 ( \20504 , \20503 , \19983 );
xor \U$20128 ( \20505 , \20502 , \20504 );
xor \U$20129 ( \20506 , \19465 , \19467 );
xor \U$20130 ( \20507 , \20506 , \19470 );
xor \U$20131 ( \20508 , \19916 , \19918 );
xor \U$20132 ( \20509 , \20508 , \19971 );
or \U$20133 ( \20510 , \20507 , \20509 );
xor \U$20134 ( \20511 , \19655 , \19659 );
xor \U$20135 ( \20512 , \20511 , \19619 );
not \U$20136 ( \20513 , \20512 );
not \U$20137 ( \20514 , \20513 );
not \U$20138 ( \20515 , \1339 );
not \U$20139 ( \20516 , \19821 );
or \U$20140 ( \20517 , \20515 , \20516 );
not \U$20141 ( \20518 , RIc2271f0_9);
not \U$20142 ( \20519 , \19721 );
not \U$20143 ( \20520 , \20519 );
or \U$20144 ( \20521 , \20518 , \20520 );
nand \U$20145 ( \20522 , \19721 , \1351 );
nand \U$20146 ( \20523 , \20521 , \20522 );
nand \U$20147 ( \20524 , \20523 , \1363 );
nand \U$20148 ( \20525 , \20517 , \20524 );
and \U$20149 ( \20526 , \16248 , \954 );
not \U$20150 ( \20527 , RIc2272e0_7);
not \U$20151 ( \20528 , \16482 );
not \U$20152 ( \20529 , \20528 );
or \U$20153 ( \20530 , \20527 , \20529 );
nand \U$20154 ( \20531 , \16256 , \1139 );
nand \U$20155 ( \20532 , \20530 , \20531 );
not \U$20156 ( \20533 , \20532 );
not \U$20157 ( \20534 , \1118 );
or \U$20158 ( \20535 , \20533 , \20534 );
or \U$20159 ( \20536 , \20397 , \1119 );
nand \U$20160 ( \20537 , \20535 , \20536 );
xor \U$20161 ( \20538 , \20526 , \20537 );
not \U$20162 ( \20539 , \1363 );
not \U$20163 ( \20540 , RIc2271f0_9);
not \U$20164 ( \20541 , \12846 );
or \U$20165 ( \20542 , \20540 , \20541 );
nand \U$20166 ( \20543 , \12845 , \1351 );
nand \U$20167 ( \20544 , \20542 , \20543 );
not \U$20168 ( \20545 , \20544 );
or \U$20169 ( \20546 , \20539 , \20545 );
nand \U$20170 ( \20547 , \20523 , \1339 );
nand \U$20171 ( \20548 , \20546 , \20547 );
and \U$20172 ( \20549 , \20538 , \20548 );
and \U$20173 ( \20550 , \20526 , \20537 );
or \U$20174 ( \20551 , \20549 , \20550 );
xor \U$20175 ( \20552 , \20525 , \20551 );
not \U$20176 ( \20553 , \1945 );
not \U$20177 ( \20554 , RIc226e30_17);
not \U$20178 ( \20555 , \17015 );
or \U$20179 ( \20556 , \20554 , \20555 );
nand \U$20180 ( \20557 , \10986 , \1935 );
nand \U$20181 ( \20558 , \20556 , \20557 );
not \U$20182 ( \20559 , \20558 );
or \U$20183 ( \20560 , \20553 , \20559 );
nand \U$20184 ( \20561 , \19955 , \1963 );
nand \U$20185 ( \20562 , \20560 , \20561 );
and \U$20186 ( \20563 , \20552 , \20562 );
and \U$20187 ( \20564 , \20525 , \20551 );
or \U$20188 ( \20565 , \20563 , \20564 );
not \U$20189 ( \20566 , \15164 );
and \U$20190 ( \20567 , RIc225a80_59, \3580 );
not \U$20191 ( \20568 , RIc225a80_59);
and \U$20192 ( \20569 , \20568 , \3579 );
or \U$20193 ( \20570 , \20567 , \20569 );
not \U$20194 ( \20571 , \20570 );
or \U$20195 ( \20572 , \20566 , \20571 );
nand \U$20196 ( \20573 , \19680 , \12670 );
nand \U$20197 ( \20574 , \20572 , \20573 );
xor \U$20198 ( \20575 , \20565 , \20574 );
not \U$20199 ( \20576 , \9444 );
not \U$20200 ( \20577 , \19541 );
or \U$20201 ( \20578 , \20576 , \20577 );
not \U$20202 ( \20579 , RIc225e40_51);
not \U$20203 ( \20580 , \2234 );
or \U$20204 ( \20581 , \20579 , \20580 );
nand \U$20205 ( \20582 , \18087 , \12423 );
nand \U$20206 ( \20583 , \20581 , \20582 );
nand \U$20207 ( \20584 , \20583 , \9459 );
nand \U$20208 ( \20585 , \20578 , \20584 );
and \U$20209 ( \20586 , \20575 , \20585 );
and \U$20210 ( \20587 , \20565 , \20574 );
or \U$20211 ( \20588 , \20586 , \20587 );
xor \U$20212 ( \20589 , \19523 , \19534 );
xor \U$20213 ( \20590 , \20589 , \19545 );
xor \U$20214 ( \20591 , \20588 , \20590 );
xor \U$20215 ( \20592 , \19617 , \19597 );
xor \U$20216 ( \20593 , \20592 , \19608 );
and \U$20217 ( \20594 , \20591 , \20593 );
and \U$20218 ( \20595 , \20588 , \20590 );
or \U$20219 ( \20596 , \20594 , \20595 );
not \U$20220 ( \20597 , \20596 );
or \U$20221 ( \20598 , \20514 , \20597 );
not \U$20222 ( \20599 , \20512 );
not \U$20223 ( \20600 , \20596 );
not \U$20224 ( \20601 , \20600 );
or \U$20225 ( \20602 , \20599 , \20601 );
xor \U$20226 ( \20603 , \19921 , \19933 );
xor \U$20227 ( \20604 , \20603 , \19960 );
not \U$20228 ( \20605 , \1682 );
not \U$20229 ( \20606 , \20323 );
or \U$20230 ( \20607 , \20605 , \20606 );
and \U$20231 ( \20608 , \1296 , \10086 );
not \U$20232 ( \20609 , \1296 );
buf \U$20233 ( \20610 , \10360 );
and \U$20234 ( \20611 , \20609 , \20610 );
nor \U$20235 ( \20612 , \20608 , \20611 );
not \U$20236 ( \20613 , \20612 );
nand \U$20237 ( \20614 , \20613 , \1678 );
nand \U$20238 ( \20615 , \20607 , \20614 );
not \U$20239 ( \20616 , \2358 );
not \U$20240 ( \20617 , \19942 );
or \U$20241 ( \20618 , \20616 , \20617 );
not \U$20242 ( \20619 , RIc226f20_15);
not \U$20243 ( \20620 , \10263 );
or \U$20244 ( \20621 , \20619 , \20620 );
nand \U$20245 ( \20622 , \9299 , \1674 );
nand \U$20246 ( \20623 , \20621 , \20622 );
nand \U$20247 ( \20624 , \20623 , \2320 );
nand \U$20248 ( \20625 , \20618 , \20624 );
xor \U$20249 ( \20626 , \20615 , \20625 );
not \U$20250 ( \20627 , \2518 );
not \U$20251 ( \20628 , RIc226d40_19);
not \U$20252 ( \20629 , \11394 );
or \U$20253 ( \20630 , \20628 , \20629 );
nand \U$20254 ( \20631 , \10653 , \2523 );
nand \U$20255 ( \20632 , \20630 , \20631 );
not \U$20256 ( \20633 , \20632 );
or \U$20257 ( \20634 , \20627 , \20633 );
nand \U$20258 ( \20635 , \20332 , \2534 );
nand \U$20259 ( \20636 , \20634 , \20635 );
and \U$20260 ( \20637 , \20626 , \20636 );
and \U$20261 ( \20638 , \20615 , \20625 );
or \U$20262 ( \20639 , \20637 , \20638 );
not \U$20263 ( \20640 , \20431 );
not \U$20264 ( \20641 , \2086 );
not \U$20265 ( \20642 , \20641 );
and \U$20266 ( \20643 , \20640 , \20642 );
and \U$20267 ( \20644 , RIc226890_29, \15699 );
not \U$20268 ( \20645 , RIc226890_29);
not \U$20269 ( \20646 , \10609 );
and \U$20270 ( \20647 , \20645 , \20646 );
or \U$20271 ( \20648 , \20644 , \20647 );
and \U$20272 ( \20649 , \20648 , \2784 );
nor \U$20273 ( \20650 , \20643 , \20649 );
not \U$20274 ( \20651 , \20650 );
not \U$20275 ( \20652 , \20651 );
not \U$20276 ( \20653 , \3629 );
not \U$20277 ( \20654 , RIc2266b0_33);
buf \U$20278 ( \20655 , \5663 );
not \U$20279 ( \20656 , \20655 );
not \U$20280 ( \20657 , \20656 );
or \U$20281 ( \20658 , \20654 , \20657 );
nand \U$20282 ( \20659 , \6726 , \9425 );
nand \U$20283 ( \20660 , \20658 , \20659 );
not \U$20284 ( \20661 , \20660 );
or \U$20285 ( \20662 , \20653 , \20661 );
not \U$20286 ( \20663 , \20354 );
nand \U$20287 ( \20664 , \20663 , \3631 );
nand \U$20288 ( \20665 , \20662 , \20664 );
not \U$20289 ( \20666 , \20665 );
or \U$20290 ( \20667 , \20652 , \20666 );
not \U$20291 ( \20668 , \20665 );
not \U$20292 ( \20669 , \20668 );
not \U$20293 ( \20670 , \20650 );
or \U$20294 ( \20671 , \20669 , \20670 );
not \U$20295 ( \20672 , \2138 );
not \U$20296 ( \20673 , RIc226980_27);
not \U$20297 ( \20674 , \12727 );
not \U$20298 ( \20675 , \20674 );
or \U$20299 ( \20676 , \20673 , \20675 );
nand \U$20300 ( \20677 , \12727 , \2799 );
nand \U$20301 ( \20678 , \20676 , \20677 );
not \U$20302 ( \20679 , \20678 );
or \U$20303 ( \20680 , \20672 , \20679 );
nand \U$20304 ( \20681 , \20379 , \2154 );
nand \U$20305 ( \20682 , \20680 , \20681 );
nand \U$20306 ( \20683 , \20671 , \20682 );
nand \U$20307 ( \20684 , \20667 , \20683 );
xor \U$20308 ( \20685 , \20639 , \20684 );
not \U$20309 ( \20686 , \1311 );
not \U$20310 ( \20687 , \20408 );
or \U$20311 ( \20688 , \20686 , \20687 );
not \U$20312 ( \20689 , RIc227100_11);
not \U$20313 ( \20690 , \12756 );
not \U$20314 ( \20691 , \20690 );
or \U$20315 ( \20692 , \20689 , \20691 );
not \U$20316 ( \20693 , \12755 );
not \U$20317 ( \20694 , \20693 );
nand \U$20318 ( \20695 , \20694 , \1302 );
nand \U$20319 ( \20696 , \20692 , \20695 );
nand \U$20320 ( \20697 , \20696 , \1306 );
nand \U$20321 ( \20698 , \20688 , \20697 );
not \U$20322 ( \20699 , \20698 );
not \U$20323 ( \20700 , RIc227010_13);
not \U$20324 ( \20701 , \13211 );
not \U$20325 ( \20702 , \20701 );
not \U$20326 ( \20703 , \20702 );
or \U$20327 ( \20704 , \20700 , \20703 );
nand \U$20328 ( \20705 , \20701 , \3841 );
nand \U$20329 ( \20706 , \20704 , \20705 );
not \U$20330 ( \20707 , \20706 );
not \U$20331 ( \20708 , \1678 );
or \U$20332 ( \20709 , \20707 , \20708 );
or \U$20333 ( \20710 , \20612 , \1757 );
nand \U$20334 ( \20711 , \20709 , \20710 );
not \U$20335 ( \20712 , \20711 );
or \U$20336 ( \20713 , \20699 , \20712 );
or \U$20337 ( \20714 , \20711 , \20698 );
or \U$20338 ( \20715 , RIc227268_8, RIc2271f0_9);
nand \U$20339 ( \20716 , \20715 , \18182 );
and \U$20340 ( \20717 , RIc227268_8, RIc2271f0_9);
nor \U$20341 ( \20718 , \20717 , \1139 );
and \U$20342 ( \20719 , \20716 , \20718 );
not \U$20343 ( \20720 , \1120 );
not \U$20344 ( \20721 , \20532 );
or \U$20345 ( \20722 , \20720 , \20721 );
and \U$20346 ( \20723 , \18356 , RIc2272e0_7);
and \U$20347 ( \20724 , \18367 , \1139 );
nor \U$20348 ( \20725 , \20723 , \20724 );
or \U$20349 ( \20726 , \20725 , \1117 );
nand \U$20350 ( \20727 , \20722 , \20726 );
and \U$20351 ( \20728 , \20719 , \20727 );
nand \U$20352 ( \20729 , \20714 , \20728 );
nand \U$20353 ( \20730 , \20713 , \20729 );
not \U$20354 ( \20731 , \2710 );
not \U$20355 ( \20732 , \20421 );
or \U$20356 ( \20733 , \20731 , \20732 );
not \U$20357 ( \20734 , RIc2267a0_31);
not \U$20358 ( \20735 , \14192 );
or \U$20359 ( \20736 , \20734 , \20735 );
nand \U$20360 ( \20737 , \6492 , \3648 );
nand \U$20361 ( \20738 , \20736 , \20737 );
nand \U$20362 ( \20739 , \20738 , \2697 );
nand \U$20363 ( \20740 , \20733 , \20739 );
xor \U$20364 ( \20741 , \20730 , \20740 );
not \U$20365 ( \20742 , \4381 );
not \U$20366 ( \20743 , RIc2265c0_35);
not \U$20367 ( \20744 , \18450 );
or \U$20368 ( \20745 , \20743 , \20744 );
nand \U$20369 ( \20746 , \4407 , \3620 );
nand \U$20370 ( \20747 , \20745 , \20746 );
not \U$20371 ( \20748 , \20747 );
or \U$20372 ( \20749 , \20742 , \20748 );
nand \U$20373 ( \20750 , \20343 , \5135 );
nand \U$20374 ( \20751 , \20749 , \20750 );
and \U$20375 ( \20752 , \20741 , \20751 );
and \U$20376 ( \20753 , \20730 , \20740 );
or \U$20377 ( \20754 , \20752 , \20753 );
and \U$20378 ( \20755 , \20685 , \20754 );
and \U$20379 ( \20756 , \20639 , \20684 );
or \U$20380 ( \20757 , \20755 , \20756 );
xor \U$20381 ( \20758 , \20604 , \20757 );
xor \U$20382 ( \20759 , \19936 , \19946 );
xor \U$20383 ( \20760 , \20759 , \19957 );
xor \U$20384 ( \20761 , \20325 , \20334 );
xor \U$20385 ( \20762 , \20761 , \20345 );
xor \U$20386 ( \20763 , \20760 , \20762 );
not \U$20387 ( \20764 , \1930 );
not \U$20388 ( \20765 , \20370 );
or \U$20389 ( \20766 , \20764 , \20765 );
not \U$20390 ( \20767 , RIc226b60_23);
not \U$20391 ( \20768 , \8975 );
or \U$20392 ( \20769 , \20767 , \20768 );
nand \U$20393 ( \20770 , \8974 , \2111 );
nand \U$20394 ( \20771 , \20769 , \20770 );
nand \U$20395 ( \20772 , \20771 , \10214 );
nand \U$20396 ( \20773 , \20766 , \20772 );
not \U$20397 ( \20774 , \2367 );
not \U$20398 ( \20775 , \20232 );
or \U$20399 ( \20776 , \20774 , \20775 );
not \U$20400 ( \20777 , RIc226c50_21);
not \U$20401 ( \20778 , \9212 );
or \U$20402 ( \20779 , \20777 , \20778 );
nand \U$20403 ( \20780 , \9211 , \2370 );
nand \U$20404 ( \20781 , \20779 , \20780 );
nand \U$20405 ( \20782 , \20781 , \2392 );
nand \U$20406 ( \20783 , \20776 , \20782 );
xor \U$20407 ( \20784 , \20773 , \20783 );
not \U$20408 ( \20785 , \2860 );
not \U$20409 ( \20786 , RIc226a70_25);
not \U$20410 ( \20787 , \8810 );
or \U$20411 ( \20788 , \20786 , \20787 );
nand \U$20412 ( \20789 , \10859 , \1905 );
nand \U$20413 ( \20790 , \20788 , \20789 );
not \U$20414 ( \20791 , \20790 );
or \U$20415 ( \20792 , \20785 , \20791 );
nand \U$20416 ( \20793 , \20221 , \2173 );
nand \U$20417 ( \20794 , \20792 , \20793 );
and \U$20418 ( \20795 , \20784 , \20794 );
and \U$20419 ( \20796 , \20773 , \20783 );
or \U$20420 ( \20797 , \20795 , \20796 );
and \U$20421 ( \20798 , \20763 , \20797 );
and \U$20422 ( \20799 , \20760 , \20762 );
or \U$20423 ( \20800 , \20798 , \20799 );
and \U$20424 ( \20801 , \20758 , \20800 );
and \U$20425 ( \20802 , \20604 , \20757 );
or \U$20426 ( \20803 , \20801 , \20802 );
nand \U$20427 ( \20804 , \20602 , \20803 );
nand \U$20428 ( \20805 , \20598 , \20804 );
nand \U$20429 ( \20806 , \20510 , \20805 );
nand \U$20430 ( \20807 , \20507 , \20509 );
and \U$20431 ( \20808 , \20806 , \20807 );
not \U$20432 ( \20809 , \20808 );
not \U$20433 ( \20810 , \20809 );
xor \U$20434 ( \20811 , \19891 , \19975 );
xor \U$20435 ( \20812 , \20811 , \19979 );
not \U$20436 ( \20813 , \20812 );
not \U$20437 ( \20814 , \20813 );
or \U$20438 ( \20815 , \20810 , \20814 );
not \U$20439 ( \20816 , \20812 );
not \U$20440 ( \20817 , \20808 );
or \U$20441 ( \20818 , \20816 , \20817 );
xor \U$20442 ( \20819 , \19456 , \19473 );
xor \U$20443 ( \20820 , \20819 , \19476 );
nand \U$20444 ( \20821 , \20818 , \20820 );
nand \U$20445 ( \20822 , \20815 , \20821 );
and \U$20446 ( \20823 , \20505 , \20822 );
and \U$20447 ( \20824 , \20502 , \20504 );
or \U$20448 ( \20825 , \20823 , \20824 );
buf \U$20449 ( \20826 , \20825 );
and \U$20450 ( \20827 , \20054 , \20826 );
not \U$20451 ( \20828 , \20040 );
nor \U$20452 ( \20829 , \20828 , \20053 );
nor \U$20453 ( \20830 , \20827 , \20829 );
nand \U$20454 ( \20831 , \20038 , \20830 );
not \U$20455 ( \20832 , \20831 );
not \U$20456 ( \20833 , \20813 );
not \U$20457 ( \20834 , \20808 );
or \U$20458 ( \20835 , \20833 , \20834 );
nand \U$20459 ( \20836 , \20809 , \20812 );
nand \U$20460 ( \20837 , \20835 , \20836 );
and \U$20461 ( \20838 , \20837 , \20820 );
not \U$20462 ( \20839 , \20837 );
not \U$20463 ( \20840 , \20820 );
and \U$20464 ( \20841 , \20839 , \20840 );
nor \U$20465 ( \20842 , \20838 , \20841 );
xor \U$20466 ( \20843 , \20604 , \20757 );
xor \U$20467 ( \20844 , \20843 , \20800 );
xor \U$20468 ( \20845 , \20639 , \20684 );
xor \U$20469 ( \20846 , \20845 , \20754 );
xor \U$20470 ( \20847 , \20415 , \20425 );
xor \U$20471 ( \20848 , \20847 , \20436 );
xor \U$20472 ( \20849 , \20565 , \20574 );
xor \U$20473 ( \20850 , \20849 , \20585 );
xor \U$20474 ( \20851 , \20848 , \20850 );
xor \U$20475 ( \20852 , \20389 , \20400 );
xor \U$20476 ( \20853 , \20852 , \20412 );
not \U$20477 ( \20854 , \15719 );
not \U$20478 ( \20855 , RIc225990_61);
not \U$20479 ( \20856 , \1393 );
or \U$20480 ( \20857 , \20855 , \20856 );
nand \U$20481 ( \20858 , \5247 , \10338 );
nand \U$20482 ( \20859 , \20857 , \20858 );
not \U$20483 ( \20860 , \20859 );
or \U$20484 ( \20861 , \20854 , \20860 );
buf \U$20485 ( \20862 , \15729 );
nand \U$20486 ( \20863 , \20092 , \20862 );
nand \U$20487 ( \20864 , \20861 , \20863 );
xor \U$20488 ( \20865 , \20853 , \20864 );
not \U$20489 ( \20866 , \10445 );
not \U$20490 ( \20867 , RIc225f30_49);
not \U$20491 ( \20868 , \2015 );
or \U$20492 ( \20869 , \20867 , \20868 );
nand \U$20493 ( \20870 , \3508 , \9541 );
nand \U$20494 ( \20871 , \20869 , \20870 );
not \U$20495 ( \20872 , \20871 );
or \U$20496 ( \20873 , \20866 , \20872 );
nand \U$20497 ( \20874 , \20210 , \9552 );
nand \U$20498 ( \20875 , \20873 , \20874 );
and \U$20499 ( \20876 , \20865 , \20875 );
and \U$20500 ( \20877 , \20853 , \20864 );
or \U$20501 ( \20878 , \20876 , \20877 );
xor \U$20502 ( \20879 , \20851 , \20878 );
xor \U$20503 ( \20880 , \20846 , \20879 );
not \U$20504 ( \20881 , \20665 );
not \U$20505 ( \20882 , \20650 );
or \U$20506 ( \20883 , \20881 , \20882 );
nand \U$20507 ( \20884 , \20668 , \20651 );
nand \U$20508 ( \20885 , \20883 , \20884 );
xor \U$20509 ( \20886 , \20885 , \20682 );
not \U$20510 ( \20887 , \11965 );
not \U$20511 ( \20888 , RIc225b70_57);
not \U$20512 ( \20889 , \12382 );
or \U$20513 ( \20890 , \20888 , \20889 );
nand \U$20514 ( \20891 , \4474 , \15262 );
nand \U$20515 ( \20892 , \20890 , \20891 );
not \U$20516 ( \20893 , \20892 );
or \U$20517 ( \20894 , \20887 , \20893 );
not \U$20518 ( \20895 , RIc225b70_57);
not \U$20519 ( \20896 , \4178 );
or \U$20520 ( \20897 , \20895 , \20896 );
nand \U$20521 ( \20898 , \1730 , \11033 );
nand \U$20522 ( \20899 , \20897 , \20898 );
nand \U$20523 ( \20900 , \20899 , \11974 );
nand \U$20524 ( \20901 , \20894 , \20900 );
not \U$20525 ( \20902 , \9552 );
not \U$20526 ( \20903 , \20871 );
or \U$20527 ( \20904 , \20902 , \20903 );
and \U$20528 ( \20905 , \2592 , RIc225f30_49);
not \U$20529 ( \20906 , \2592 );
and \U$20530 ( \20907 , \20906 , \9541 );
or \U$20531 ( \20908 , \20905 , \20907 );
nand \U$20532 ( \20909 , \20908 , \10445 );
nand \U$20533 ( \20910 , \20904 , \20909 );
xor \U$20534 ( \20911 , \20901 , \20910 );
not \U$20535 ( \20912 , \9619 );
not \U$20536 ( \20913 , RIc226020_47);
not \U$20537 ( \20914 , \2556 );
or \U$20538 ( \20915 , \20913 , \20914 );
nand \U$20539 ( \20916 , \3450 , \9624 );
nand \U$20540 ( \20917 , \20915 , \20916 );
not \U$20541 ( \20918 , \20917 );
or \U$20542 ( \20919 , \20912 , \20918 );
not \U$20543 ( \20920 , RIc226020_47);
not \U$20544 ( \20921 , \5819 );
or \U$20545 ( \20922 , \20920 , \20921 );
nand \U$20546 ( \20923 , \2480 , \9624 );
nand \U$20547 ( \20924 , \20922 , \20923 );
nand \U$20548 ( \20925 , \20924 , \9641 );
nand \U$20549 ( \20926 , \20919 , \20925 );
and \U$20550 ( \20927 , \20911 , \20926 );
and \U$20551 ( \20928 , \20901 , \20910 );
or \U$20552 ( \20929 , \20927 , \20928 );
xor \U$20553 ( \20930 , \20886 , \20929 );
not \U$20554 ( \20931 , \9398 );
not \U$20555 ( \20932 , \20116 );
or \U$20556 ( \20933 , \20931 , \20932 );
not \U$20557 ( \20934 , RIc226110_45);
not \U$20558 ( \20935 , \3021 );
or \U$20559 ( \20936 , \20934 , \20935 );
nand \U$20560 ( \20937 , \2498 , \14390 );
nand \U$20561 ( \20938 , \20936 , \20937 );
nand \U$20562 ( \20939 , \20938 , \9384 );
nand \U$20563 ( \20940 , \20933 , \20939 );
not \U$20564 ( \20941 , \9641 );
not \U$20565 ( \20942 , \20917 );
or \U$20566 ( \20943 , \20941 , \20942 );
nand \U$20567 ( \20944 , \20101 , \9619 );
nand \U$20568 ( \20945 , \20943 , \20944 );
xor \U$20569 ( \20946 , \20940 , \20945 );
not \U$20570 ( \20947 , \11965 );
not \U$20571 ( \20948 , \20899 );
or \U$20572 ( \20949 , \20947 , \20948 );
nand \U$20573 ( \20950 , \20080 , \11974 );
nand \U$20574 ( \20951 , \20949 , \20950 );
xor \U$20575 ( \20952 , \20946 , \20951 );
and \U$20576 ( \20953 , \20930 , \20952 );
and \U$20577 ( \20954 , \20886 , \20929 );
or \U$20578 ( \20955 , \20953 , \20954 );
and \U$20579 ( \20956 , \20880 , \20955 );
and \U$20580 ( \20957 , \20846 , \20879 );
or \U$20581 ( \20958 , \20956 , \20957 );
xor \U$20582 ( \20959 , \20844 , \20958 );
xor \U$20583 ( \20960 , \20372 , \20383 );
xor \U$20584 ( \20961 , \20960 , \20359 );
xor \U$20585 ( \20962 , \20225 , \20237 );
xor \U$20586 ( \20963 , \20962 , \20212 );
xor \U$20587 ( \20964 , \20961 , \20963 );
not \U$20588 ( \20965 , \9705 );
not \U$20589 ( \20966 , \20185 );
or \U$20590 ( \20967 , \20965 , \20966 );
and \U$20591 ( \20968 , \6303 , \2634 );
not \U$20592 ( \20969 , \6303 );
and \U$20593 ( \20970 , \20969 , \4227 );
nor \U$20594 ( \20971 , \20968 , \20970 );
not \U$20595 ( \20972 , \20971 );
nand \U$20596 ( \20973 , \20972 , \9690 );
nand \U$20597 ( \20974 , \20967 , \20973 );
not \U$20598 ( \20975 , \6307 );
not \U$20599 ( \20976 , \20274 );
or \U$20600 ( \20977 , \20975 , \20976 );
not \U$20601 ( \20978 , RIc2263e0_39);
not \U$20602 ( \20979 , \11321 );
or \U$20603 ( \20980 , \20978 , \20979 );
not \U$20604 ( \20981 , RIc2263e0_39);
nand \U$20605 ( \20982 , \20981 , \11324 );
nand \U$20606 ( \20983 , \20980 , \20982 );
nand \U$20607 ( \20984 , \20983 , \6688 );
nand \U$20608 ( \20985 , \20977 , \20984 );
nor \U$20609 ( \20986 , \20974 , \20985 );
not \U$20610 ( \20987 , \12945 );
not \U$20611 ( \20988 , \20169 );
or \U$20612 ( \20989 , \20987 , \20988 );
not \U$20613 ( \20990 , RIc225d50_53);
not \U$20614 ( \20991 , \9570 );
or \U$20615 ( \20992 , \20990 , \20991 );
nand \U$20616 ( \20993 , \2443 , \11585 );
nand \U$20617 ( \20994 , \20992 , \20993 );
nand \U$20618 ( \20995 , \20994 , \8777 );
nand \U$20619 ( \20996 , \20989 , \20995 );
not \U$20620 ( \20997 , \20996 );
or \U$20621 ( \20998 , \20986 , \20997 );
nand \U$20622 ( \20999 , \20974 , \20985 );
nand \U$20623 ( \21000 , \20998 , \20999 );
xnor \U$20624 ( \21001 , \20964 , \21000 );
not \U$20625 ( \21002 , \9129 );
not \U$20626 ( \21003 , \20129 );
or \U$20627 ( \21004 , \21002 , \21003 );
not \U$20628 ( \21005 , RIc226200_43);
not \U$20629 ( \21006 , \2063 );
or \U$20630 ( \21007 , \21005 , \21006 );
nand \U$20631 ( \21008 , \3008 , \13805 );
nand \U$20632 ( \21009 , \21007 , \21008 );
nand \U$20633 ( \21010 , \21009 , \9110 );
nand \U$20634 ( \21011 , \21004 , \21010 );
not \U$20635 ( \21012 , \11117 );
not \U$20636 ( \21013 , RIc225c60_55);
not \U$20637 ( \21014 , \3092 );
or \U$20638 ( \21015 , \21013 , \21014 );
nand \U$20639 ( \21016 , \8989 , \11108 );
nand \U$20640 ( \21017 , \21015 , \21016 );
not \U$20641 ( \21018 , \21017 );
or \U$20642 ( \21019 , \21012 , \21018 );
nand \U$20643 ( \21020 , \20140 , \11038 );
nand \U$20644 ( \21021 , \21019 , \21020 );
xor \U$20645 ( \21022 , \21011 , \21021 );
not \U$20646 ( \21023 , \16891 );
not \U$20647 ( \21024 , RIc2258a0_63);
not \U$20648 ( \21025 , \3993 );
or \U$20649 ( \21026 , \21024 , \21025 );
nand \U$20650 ( \21027 , \1403 , \16880 );
nand \U$20651 ( \21028 , \21026 , \21027 );
not \U$20652 ( \21029 , \21028 );
or \U$20653 ( \21030 , \21023 , \21029 );
nand \U$20654 ( \21031 , \20158 , RIc225828_64);
nand \U$20655 ( \21032 , \21030 , \21031 );
and \U$20656 ( \21033 , \21022 , \21032 );
and \U$20657 ( \21034 , \21011 , \21021 );
or \U$20658 ( \21035 , \21033 , \21034 );
not \U$20659 ( \21036 , \20951 );
not \U$20660 ( \21037 , \20940 );
or \U$20661 ( \21038 , \21036 , \21037 );
or \U$20662 ( \21039 , \20940 , \20951 );
nand \U$20663 ( \21040 , \21039 , \20945 );
nand \U$20664 ( \21041 , \21038 , \21040 );
xor \U$20665 ( \21042 , \21035 , \21041 );
not \U$20666 ( \21043 , \9459 );
not \U$20667 ( \21044 , RIc225e40_51);
not \U$20668 ( \21045 , \4009 );
or \U$20669 ( \21046 , \21044 , \21045 );
nand \U$20670 ( \21047 , \4008 , \9450 );
nand \U$20671 ( \21048 , \21046 , \21047 );
not \U$20672 ( \21049 , \21048 );
or \U$20673 ( \21050 , \21043 , \21049 );
nand \U$20674 ( \21051 , \20583 , \9444 );
nand \U$20675 ( \21052 , \21050 , \21051 );
not \U$20676 ( \21053 , \21052 );
not \U$20677 ( \21054 , \15164 );
and \U$20678 ( \21055 , RIc225a80_59, \1949 );
not \U$20679 ( \21056 , RIc225a80_59);
and \U$20680 ( \21057 , \21056 , \3918 );
or \U$20681 ( \21058 , \21055 , \21057 );
not \U$20682 ( \21059 , \21058 );
or \U$20683 ( \21060 , \21054 , \21059 );
nand \U$20684 ( \21061 , \20570 , \12670 );
nand \U$20685 ( \21062 , \21060 , \21061 );
not \U$20686 ( \21063 , \21062 );
or \U$20687 ( \21064 , \21053 , \21063 );
or \U$20688 ( \21065 , \21062 , \21052 );
not \U$20689 ( \21066 , \5519 );
not \U$20690 ( \21067 , \20283 );
or \U$20691 ( \21068 , \21066 , \21067 );
not \U$20692 ( \21069 , RIc2264d0_37);
not \U$20693 ( \21070 , \19926 );
or \U$20694 ( \21071 , \21069 , \21070 );
nand \U$20695 ( \21072 , \3641 , \4371 );
nand \U$20696 ( \21073 , \21071 , \21072 );
nand \U$20697 ( \21074 , \21073 , \5509 );
nand \U$20698 ( \21075 , \21068 , \21074 );
nand \U$20699 ( \21076 , \21065 , \21075 );
nand \U$20700 ( \21077 , \21064 , \21076 );
xor \U$20701 ( \21078 , \21042 , \21077 );
xor \U$20702 ( \21079 , \21001 , \21078 );
not \U$20703 ( \21080 , \1682 );
not \U$20704 ( \21081 , \20706 );
or \U$20705 ( \21082 , \21080 , \21081 );
not \U$20706 ( \21083 , RIc227010_13);
not \U$20707 ( \21084 , \10356 );
not \U$20708 ( \21085 , \21084 );
or \U$20709 ( \21086 , \21083 , \21085 );
nand \U$20710 ( \21087 , \13497 , \1758 );
nand \U$20711 ( \21088 , \21086 , \21087 );
nand \U$20712 ( \21089 , \21088 , \1678 );
nand \U$20713 ( \21090 , \21082 , \21089 );
and \U$20714 ( \21091 , \18182 , \1120 );
not \U$20715 ( \21092 , \1339 );
not \U$20716 ( \21093 , RIc2271f0_9);
not \U$20717 ( \21094 , \13487 );
not \U$20718 ( \21095 , \21094 );
or \U$20719 ( \21096 , \21093 , \21095 );
not \U$20720 ( \21097 , \21094 );
nand \U$20721 ( \21098 , \21097 , \1342 );
nand \U$20722 ( \21099 , \21096 , \21098 );
not \U$20723 ( \21100 , \21099 );
or \U$20724 ( \21101 , \21092 , \21100 );
not \U$20725 ( \21102 , \16256 );
and \U$20726 ( \21103 , \1342 , \21102 );
not \U$20727 ( \21104 , \1342 );
and \U$20728 ( \21105 , \21104 , \16482 );
nor \U$20729 ( \21106 , \21103 , \21105 );
nand \U$20730 ( \21107 , \21106 , \1362 );
nand \U$20731 ( \21108 , \21101 , \21107 );
xor \U$20732 ( \21109 , \21091 , \21108 );
not \U$20733 ( \21110 , \1306 );
not \U$20734 ( \21111 , RIc227100_11);
not \U$20735 ( \21112 , \18158 );
or \U$20736 ( \21113 , \21111 , \21112 );
nand \U$20737 ( \21114 , \18161 , \3351 );
nand \U$20738 ( \21115 , \21113 , \21114 );
not \U$20739 ( \21116 , \21115 );
or \U$20740 ( \21117 , \21110 , \21116 );
not \U$20741 ( \21118 , RIc227100_11);
not \U$20742 ( \21119 , \15444 );
or \U$20743 ( \21120 , \21118 , \21119 );
nand \U$20744 ( \21121 , \15443 , \1685 );
nand \U$20745 ( \21122 , \21120 , \21121 );
nand \U$20746 ( \21123 , \21122 , \1310 );
nand \U$20747 ( \21124 , \21117 , \21123 );
and \U$20748 ( \21125 , \21109 , \21124 );
and \U$20749 ( \21126 , \21091 , \21108 );
or \U$20750 ( \21127 , \21125 , \21126 );
xor \U$20751 ( \21128 , \21090 , \21127 );
not \U$20752 ( \21129 , \2518 );
and \U$20753 ( \21130 , \2523 , \9250 );
not \U$20754 ( \21131 , \2523 );
and \U$20755 ( \21132 , \21131 , \17014 );
nor \U$20756 ( \21133 , \21130 , \21132 );
not \U$20757 ( \21134 , \21133 );
or \U$20758 ( \21135 , \21129 , \21134 );
not \U$20759 ( \21136 , RIc226d40_19);
not \U$20760 ( \21137 , \10814 );
or \U$20761 ( \21138 , \21136 , \21137 );
nand \U$20762 ( \21139 , \10110 , \3338 );
nand \U$20763 ( \21140 , \21138 , \21139 );
nand \U$20764 ( \21141 , \21140 , \2534 );
nand \U$20765 ( \21142 , \21135 , \21141 );
and \U$20766 ( \21143 , \21128 , \21142 );
and \U$20767 ( \21144 , \21090 , \21127 );
or \U$20768 ( \21145 , \21143 , \21144 );
not \U$20769 ( \21146 , \1945 );
not \U$20770 ( \21147 , RIc226e30_17);
not \U$20771 ( \21148 , \10263 );
or \U$20772 ( \21149 , \21147 , \21148 );
not \U$20773 ( \21150 , \9297 );
nand \U$20774 ( \21151 , \21150 , \1935 );
nand \U$20775 ( \21152 , \21149 , \21151 );
not \U$20776 ( \21153 , \21152 );
or \U$20777 ( \21154 , \21146 , \21153 );
not \U$20778 ( \21155 , RIc226e30_17);
not \U$20779 ( \21156 , \9275 );
not \U$20780 ( \21157 , \21156 );
or \U$20781 ( \21158 , \21155 , \21157 );
nand \U$20782 ( \21159 , \9275 , \1952 );
nand \U$20783 ( \21160 , \21158 , \21159 );
nand \U$20784 ( \21161 , \21160 , \1963 );
nand \U$20785 ( \21162 , \21154 , \21161 );
not \U$20786 ( \21163 , \2358 );
not \U$20787 ( \21164 , RIc226f20_15);
not \U$20788 ( \21165 , \13442 );
or \U$20789 ( \21166 , \21164 , \21165 );
nand \U$20790 ( \21167 , \9320 , \2301 );
nand \U$20791 ( \21168 , \21166 , \21167 );
not \U$20792 ( \21169 , \21168 );
or \U$20793 ( \21170 , \21163 , \21169 );
not \U$20794 ( \21171 , RIc226f20_15);
not \U$20795 ( \21172 , \10086 );
not \U$20796 ( \21173 , \21172 );
or \U$20797 ( \21174 , \21171 , \21173 );
not \U$20798 ( \21175 , \16945 );
nand \U$20799 ( \21176 , \21175 , \2301 );
nand \U$20800 ( \21177 , \21174 , \21176 );
nand \U$20801 ( \21178 , \21177 , \2320 );
nand \U$20802 ( \21179 , \21170 , \21178 );
xor \U$20803 ( \21180 , \21162 , \21179 );
not \U$20804 ( \21181 , \2367 );
not \U$20805 ( \21182 , RIc226c50_21);
not \U$20806 ( \21183 , \9051 );
not \U$20807 ( \21184 , \21183 );
or \U$20808 ( \21185 , \21182 , \21184 );
not \U$20809 ( \21186 , \13465 );
nand \U$20810 ( \21187 , \21186 , \2370 );
nand \U$20811 ( \21188 , \21185 , \21187 );
not \U$20812 ( \21189 , \21188 );
or \U$20813 ( \21190 , \21181 , \21189 );
not \U$20814 ( \21191 , RIc226c50_21);
not \U$20815 ( \21192 , \19789 );
or \U$20816 ( \21193 , \21191 , \21192 );
nand \U$20817 ( \21194 , \19790 , \2370 );
nand \U$20818 ( \21195 , \21193 , \21194 );
nand \U$20819 ( \21196 , \21195 , \2392 );
nand \U$20820 ( \21197 , \21190 , \21196 );
and \U$20821 ( \21198 , \21180 , \21197 );
and \U$20822 ( \21199 , \21162 , \21179 );
or \U$20823 ( \21200 , \21198 , \21199 );
xor \U$20824 ( \21201 , \21145 , \21200 );
not \U$20825 ( \21202 , \18037 );
not \U$20826 ( \21203 , \21058 );
or \U$20827 ( \21204 , \21202 , \21203 );
and \U$20828 ( \21205 , RIc225a80_59, \1487 );
not \U$20829 ( \21206 , RIc225a80_59);
and \U$20830 ( \21207 , \21206 , \3043 );
or \U$20831 ( \21208 , \21205 , \21207 );
nand \U$20832 ( \21209 , \21208 , \15164 );
nand \U$20833 ( \21210 , \21204 , \21209 );
and \U$20834 ( \21211 , \21201 , \21210 );
and \U$20835 ( \21212 , \21145 , \21200 );
or \U$20836 ( \21213 , \21211 , \21212 );
xor \U$20837 ( \21214 , \20853 , \20864 );
xor \U$20838 ( \21215 , \21214 , \20875 );
xor \U$20839 ( \21216 , \21213 , \21215 );
xor \U$20840 ( \21217 , \21052 , \21062 );
xor \U$20841 ( \21218 , \21217 , \21075 );
and \U$20842 ( \21219 , \21216 , \21218 );
and \U$20843 ( \21220 , \21213 , \21215 );
or \U$20844 ( \21221 , \21219 , \21220 );
and \U$20845 ( \21222 , \21079 , \21221 );
and \U$20846 ( \21223 , \21001 , \21078 );
or \U$20847 ( \21224 , \21222 , \21223 );
and \U$20848 ( \21225 , \20959 , \21224 );
and \U$20849 ( \21226 , \20844 , \20958 );
or \U$20850 ( \21227 , \21225 , \21226 );
not \U$20851 ( \21228 , \21227 );
not \U$20852 ( \21229 , \19903 );
not \U$20853 ( \21230 , \19911 );
or \U$20854 ( \21231 , \21229 , \21230 );
not \U$20855 ( \21232 , \19903 );
nand \U$20856 ( \21233 , \21232 , \19910 );
nand \U$20857 ( \21234 , \21231 , \21233 );
buf \U$20858 ( \21235 , \19906 );
not \U$20859 ( \21236 , \21235 );
and \U$20860 ( \21237 , \21234 , \21236 );
not \U$20861 ( \21238 , \21234 );
and \U$20862 ( \21239 , \21238 , \21235 );
nor \U$20863 ( \21240 , \21237 , \21239 );
xor \U$20864 ( \21241 , \19963 , \19965 );
xor \U$20865 ( \21242 , \21241 , \19968 );
xor \U$20866 ( \21243 , \21240 , \21242 );
not \U$20867 ( \21244 , \20264 );
not \U$20868 ( \21245 , \20444 );
or \U$20869 ( \21246 , \21244 , \21245 );
or \U$20870 ( \21247 , \20444 , \20264 );
nand \U$20871 ( \21248 , \21246 , \21247 );
and \U$20872 ( \21249 , \21248 , \20447 );
not \U$20873 ( \21250 , \21248 );
and \U$20874 ( \21251 , \21250 , \20313 );
nor \U$20875 ( \21252 , \21249 , \21251 );
xor \U$20876 ( \21253 , \21243 , \21252 );
not \U$20877 ( \21254 , \21253 );
xor \U$20878 ( \21255 , \20588 , \20590 );
xor \U$20879 ( \21256 , \21255 , \20593 );
not \U$20880 ( \21257 , \21256 );
xor \U$20881 ( \21258 , \20760 , \20762 );
xor \U$20882 ( \21259 , \21258 , \20797 );
not \U$20883 ( \21260 , \21259 );
xor \U$20884 ( \21261 , \20773 , \20783 );
xor \U$20885 ( \21262 , \21261 , \20794 );
not \U$20886 ( \21263 , \21262 );
not \U$20887 ( \21264 , \6307 );
not \U$20888 ( \21265 , \20983 );
or \U$20889 ( \21266 , \21264 , \21265 );
not \U$20890 ( \21267 , RIc2263e0_39);
not \U$20891 ( \21268 , \11672 );
or \U$20892 ( \21269 , \21267 , \21268 );
nand \U$20893 ( \21270 , \2980 , \5498 );
nand \U$20894 ( \21271 , \21269 , \21270 );
nand \U$20895 ( \21272 , \21271 , \6689 );
nand \U$20896 ( \21273 , \21266 , \21272 );
not \U$20897 ( \21274 , \21273 );
not \U$20898 ( \21275 , \20971 );
not \U$20899 ( \21276 , \9705 );
not \U$20900 ( \21277 , \21276 );
and \U$20901 ( \21278 , \21275 , \21277 );
not \U$20902 ( \21279 , RIc2262f0_41);
not \U$20903 ( \21280 , \3715 );
or \U$20904 ( \21281 , \21279 , \21280 );
nand \U$20905 ( \21282 , \15217 , \9822 );
nand \U$20906 ( \21283 , \21281 , \21282 );
and \U$20907 ( \21284 , \21283 , \9690 );
nor \U$20908 ( \21285 , \21278 , \21284 );
not \U$20909 ( \21286 , \21285 );
not \U$20910 ( \21287 , \21286 );
or \U$20911 ( \21288 , \21274 , \21287 );
not \U$20912 ( \21289 , \21273 );
not \U$20913 ( \21290 , \21289 );
not \U$20914 ( \21291 , \21285 );
or \U$20915 ( \21292 , \21290 , \21291 );
not \U$20916 ( \21293 , \8777 );
and \U$20917 ( \21294 , RIc225d50_53, \18086 );
not \U$20918 ( \21295 , RIc225d50_53);
and \U$20919 ( \21296 , \21295 , \11648 );
or \U$20920 ( \21297 , \21294 , \21296 );
not \U$20921 ( \21298 , \21297 );
or \U$20922 ( \21299 , \21293 , \21298 );
nand \U$20923 ( \21300 , \20994 , \9555 );
nand \U$20924 ( \21301 , \21299 , \21300 );
nand \U$20925 ( \21302 , \21292 , \21301 );
nand \U$20926 ( \21303 , \21288 , \21302 );
not \U$20927 ( \21304 , \21303 );
or \U$20928 ( \21305 , \21263 , \21304 );
or \U$20929 ( \21306 , \21303 , \21262 );
not \U$20930 ( \21307 , RIc225828_64);
not \U$20931 ( \21308 , \21028 );
or \U$20932 ( \21309 , \21307 , \21308 );
not \U$20933 ( \21310 , RIc2258a0_63);
not \U$20934 ( \21311 , \3670 );
or \U$20935 ( \21312 , \21310 , \21311 );
nand \U$20936 ( \21313 , \1371 , \16880 );
nand \U$20937 ( \21314 , \21312 , \21313 );
nand \U$20938 ( \21315 , \21314 , \20159 );
nand \U$20939 ( \21316 , \21309 , \21315 );
not \U$20940 ( \21317 , \21316 );
not \U$20941 ( \21318 , \11708 );
not \U$20942 ( \21319 , \21048 );
or \U$20943 ( \21320 , \21318 , \21319 );
not \U$20944 ( \21321 , RIc225e40_51);
not \U$20945 ( \21322 , \5767 );
or \U$20946 ( \21323 , \21321 , \21322 );
nand \U$20947 ( \21324 , \3834 , \9450 );
nand \U$20948 ( \21325 , \21323 , \21324 );
nand \U$20949 ( \21326 , \21325 , \9459 );
nand \U$20950 ( \21327 , \21320 , \21326 );
not \U$20951 ( \21328 , \21327 );
or \U$20952 ( \21329 , \21317 , \21328 );
or \U$20953 ( \21330 , \21316 , \21327 );
xor \U$20954 ( \21331 , \20728 , \20698 );
xnor \U$20955 ( \21332 , \21331 , \20711 );
not \U$20956 ( \21333 , \21332 );
nand \U$20957 ( \21334 , \21330 , \21333 );
nand \U$20958 ( \21335 , \21329 , \21334 );
nand \U$20959 ( \21336 , \21306 , \21335 );
nand \U$20960 ( \21337 , \21305 , \21336 );
not \U$20961 ( \21338 , \21337 );
or \U$20962 ( \21339 , \21260 , \21338 );
or \U$20963 ( \21340 , \21337 , \21259 );
not \U$20964 ( \21341 , \15719 );
and \U$20965 ( \21342 , RIc225990_61, \1531 );
not \U$20966 ( \21343 , RIc225990_61);
and \U$20967 ( \21344 , \21343 , \3581 );
or \U$20968 ( \21345 , \21342 , \21344 );
not \U$20969 ( \21346 , \21345 );
or \U$20970 ( \21347 , \21341 , \21346 );
nand \U$20971 ( \21348 , \20859 , \15729 );
nand \U$20972 ( \21349 , \21347 , \21348 );
not \U$20973 ( \21350 , \21349 );
not \U$20974 ( \21351 , \2860 );
not \U$20975 ( \21352 , RIc226a70_25);
not \U$20976 ( \21353 , \20367 );
or \U$20977 ( \21354 , \21352 , \21353 );
nand \U$20978 ( \21355 , \8952 , \6107 );
nand \U$20979 ( \21356 , \21354 , \21355 );
not \U$20980 ( \21357 , \21356 );
or \U$20981 ( \21358 , \21351 , \21357 );
nand \U$20982 ( \21359 , \20790 , \2173 );
nand \U$20983 ( \21360 , \21358 , \21359 );
not \U$20984 ( \21361 , \21360 );
nand \U$20985 ( \21362 , \21350 , \21361 );
not \U$20986 ( \21363 , \4383 );
not \U$20987 ( \21364 , \20747 );
or \U$20988 ( \21365 , \21363 , \21364 );
not \U$20989 ( \21366 , RIc2265c0_35);
not \U$20990 ( \21367 , \5216 );
or \U$20991 ( \21368 , \21366 , \21367 );
not \U$20992 ( \21369 , \13512 );
nand \U$20993 ( \21370 , \21369 , \9587 );
nand \U$20994 ( \21371 , \21368 , \21370 );
nand \U$20995 ( \21372 , \21371 , \4381 );
nand \U$20996 ( \21373 , \21365 , \21372 );
and \U$20997 ( \21374 , \21362 , \21373 );
nor \U$20998 ( \21375 , \21350 , \21361 );
nor \U$20999 ( \21376 , \21374 , \21375 );
not \U$21000 ( \21377 , \21376 );
not \U$21001 ( \21378 , \21377 );
not \U$21002 ( \21379 , \9934 );
not \U$21003 ( \21380 , RIc226110_45);
not \U$21004 ( \21381 , \12548 );
or \U$21005 ( \21382 , \21380 , \21381 );
nand \U$21006 ( \21383 , \2720 , \9100 );
nand \U$21007 ( \21384 , \21382 , \21383 );
not \U$21008 ( \21385 , \21384 );
or \U$21009 ( \21386 , \21379 , \21385 );
nand \U$21010 ( \21387 , \20938 , \11825 );
nand \U$21011 ( \21388 , \21386 , \21387 );
not \U$21012 ( \21389 , \11697 );
not \U$21013 ( \21390 , RIc225c60_55);
not \U$21014 ( \21391 , \3686 );
or \U$21015 ( \21392 , \21390 , \21391 );
nand \U$21016 ( \21393 , \2422 , \11041 );
nand \U$21017 ( \21394 , \21392 , \21393 );
not \U$21018 ( \21395 , \21394 );
or \U$21019 ( \21396 , \21389 , \21395 );
nand \U$21020 ( \21397 , \21017 , \13025 );
nand \U$21021 ( \21398 , \21396 , \21397 );
xor \U$21022 ( \21399 , \21388 , \21398 );
not \U$21023 ( \21400 , \9110 );
not \U$21024 ( \21401 , RIc226200_43);
not \U$21025 ( \21402 , \12310 );
or \U$21026 ( \21403 , \21401 , \21402 );
nand \U$21027 ( \21404 , \11515 , \9106 );
nand \U$21028 ( \21405 , \21403 , \21404 );
not \U$21029 ( \21406 , \21405 );
or \U$21030 ( \21407 , \21400 , \21406 );
nand \U$21031 ( \21408 , \21009 , \9205 );
nand \U$21032 ( \21409 , \21407 , \21408 );
and \U$21033 ( \21410 , \21399 , \21409 );
and \U$21034 ( \21411 , \21388 , \21398 );
or \U$21035 ( \21412 , \21410 , \21411 );
not \U$21036 ( \21413 , \21412 );
or \U$21037 ( \21414 , \21378 , \21413 );
not \U$21038 ( \21415 , \21412 );
not \U$21039 ( \21416 , \21415 );
not \U$21040 ( \21417 , \21376 );
or \U$21041 ( \21418 , \21416 , \21417 );
xor \U$21042 ( \21419 , \20730 , \20740 );
xor \U$21043 ( \21420 , \21419 , \20751 );
nand \U$21044 ( \21421 , \21418 , \21420 );
nand \U$21045 ( \21422 , \21414 , \21421 );
nand \U$21046 ( \21423 , \21340 , \21422 );
nand \U$21047 ( \21424 , \21339 , \21423 );
not \U$21048 ( \21425 , \21424 );
or \U$21049 ( \21426 , \21257 , \21425 );
or \U$21050 ( \21427 , \21424 , \21256 );
xor \U$21051 ( \21428 , \20525 , \20551 );
xor \U$21052 ( \21429 , \21428 , \20562 );
not \U$21053 ( \21430 , \2358 );
not \U$21054 ( \21431 , \20623 );
or \U$21055 ( \21432 , \21430 , \21431 );
nand \U$21056 ( \21433 , \21168 , \2320 );
nand \U$21057 ( \21434 , \21432 , \21433 );
not \U$21058 ( \21435 , \21434 );
not \U$21059 ( \21436 , \2697 );
not \U$21060 ( \21437 , RIc2267a0_31);
not \U$21061 ( \21438 , \9740 );
not \U$21062 ( \21439 , \21438 );
or \U$21063 ( \21440 , \21437 , \21439 );
nand \U$21064 ( \21441 , \9740 , \2705 );
nand \U$21065 ( \21442 , \21440 , \21441 );
not \U$21066 ( \21443 , \21442 );
or \U$21067 ( \21444 , \21436 , \21443 );
nand \U$21068 ( \21445 , \20738 , \2710 );
nand \U$21069 ( \21446 , \21444 , \21445 );
not \U$21070 ( \21447 , \21446 );
or \U$21071 ( \21448 , \21435 , \21447 );
or \U$21072 ( \21449 , \21446 , \21434 );
not \U$21073 ( \21450 , \1945 );
not \U$21074 ( \21451 , \21160 );
or \U$21075 ( \21452 , \21450 , \21451 );
nand \U$21076 ( \21453 , \20558 , \1963 );
nand \U$21077 ( \21454 , \21452 , \21453 );
nand \U$21078 ( \21455 , \21449 , \21454 );
nand \U$21079 ( \21456 , \21448 , \21455 );
xor \U$21080 ( \21457 , \21429 , \21456 );
xor \U$21081 ( \21458 , \20526 , \20537 );
xor \U$21082 ( \21459 , \21458 , \20548 );
not \U$21083 ( \21460 , \2534 );
not \U$21084 ( \21461 , \20632 );
or \U$21085 ( \21462 , \21460 , \21461 );
nand \U$21086 ( \21463 , \21140 , \2518 );
nand \U$21087 ( \21464 , \21462 , \21463 );
xor \U$21088 ( \21465 , \21459 , \21464 );
not \U$21089 ( \21466 , \2367 );
not \U$21090 ( \21467 , \20781 );
or \U$21091 ( \21468 , \21466 , \21467 );
nand \U$21092 ( \21469 , \21188 , \2392 );
nand \U$21093 ( \21470 , \21468 , \21469 );
and \U$21094 ( \21471 , \21465 , \21470 );
and \U$21095 ( \21472 , \21459 , \21464 );
or \U$21096 ( \21473 , \21471 , \21472 );
and \U$21097 ( \21474 , \21457 , \21473 );
and \U$21098 ( \21475 , \21429 , \21456 );
or \U$21099 ( \21476 , \21474 , \21475 );
not \U$21100 ( \21477 , \21476 );
xor \U$21101 ( \21478 , \20131 , \20120 );
xnor \U$21102 ( \21479 , \21478 , \20144 );
nand \U$21103 ( \21480 , \21477 , \21479 );
not \U$21104 ( \21481 , \21480 );
xor \U$21105 ( \21482 , \20615 , \20625 );
xor \U$21106 ( \21483 , \21482 , \20636 );
not \U$21107 ( \21484 , \10214 );
not \U$21108 ( \21485 , RIc226b60_23);
not \U$21109 ( \21486 , \8910 );
or \U$21110 ( \21487 , \21485 , \21486 );
nand \U$21111 ( \21488 , \12406 , \5637 );
nand \U$21112 ( \21489 , \21487 , \21488 );
not \U$21113 ( \21490 , \21489 );
or \U$21114 ( \21491 , \21484 , \21490 );
nand \U$21115 ( \21492 , \20771 , \5365 );
nand \U$21116 ( \21493 , \21491 , \21492 );
not \U$21117 ( \21494 , \21493 );
not \U$21118 ( \21495 , \3631 );
not \U$21119 ( \21496 , \20660 );
or \U$21120 ( \21497 , \21495 , \21496 );
not \U$21121 ( \21498 , RIc2266b0_33);
not \U$21122 ( \21499 , \17549 );
or \U$21123 ( \21500 , \21498 , \21499 );
nand \U$21124 ( \21501 , \9875 , \5179 );
nand \U$21125 ( \21502 , \21500 , \21501 );
nand \U$21126 ( \21503 , \21502 , \3629 );
nand \U$21127 ( \21504 , \21497 , \21503 );
not \U$21128 ( \21505 , \21504 );
or \U$21129 ( \21506 , \21494 , \21505 );
or \U$21130 ( \21507 , \21504 , \21493 );
not \U$21131 ( \21508 , \5519 );
not \U$21132 ( \21509 , \21073 );
or \U$21133 ( \21510 , \21508 , \21509 );
not \U$21134 ( \21511 , RIc2264d0_37);
not \U$21135 ( \21512 , \16519 );
not \U$21136 ( \21513 , \21512 );
or \U$21137 ( \21514 , \21511 , \21513 );
nand \U$21138 ( \21515 , \4418 , \4371 );
nand \U$21139 ( \21516 , \21514 , \21515 );
nand \U$21140 ( \21517 , \21516 , \5509 );
nand \U$21141 ( \21518 , \21510 , \21517 );
nand \U$21142 ( \21519 , \21507 , \21518 );
nand \U$21143 ( \21520 , \21506 , \21519 );
xor \U$21144 ( \21521 , \21483 , \21520 );
not \U$21145 ( \21522 , \1339 );
not \U$21146 ( \21523 , \20544 );
or \U$21147 ( \21524 , \21522 , \21523 );
nand \U$21148 ( \21525 , \21099 , \1363 );
nand \U$21149 ( \21526 , \21524 , \21525 );
xor \U$21150 ( \21527 , \20719 , \20727 );
xor \U$21151 ( \21528 , \21526 , \21527 );
not \U$21152 ( \21529 , \1311 );
not \U$21153 ( \21530 , \20696 );
or \U$21154 ( \21531 , \21529 , \21530 );
nand \U$21155 ( \21532 , \21122 , \1306 );
nand \U$21156 ( \21533 , \21531 , \21532 );
and \U$21157 ( \21534 , \21528 , \21533 );
and \U$21158 ( \21535 , \21526 , \21527 );
or \U$21159 ( \21536 , \21534 , \21535 );
not \U$21160 ( \21537 , \9142 );
not \U$21161 ( \21538 , \20648 );
or \U$21162 ( \21539 , \21537 , \21538 );
and \U$21163 ( \21540 , RIc226890_29, \16531 );
not \U$21164 ( \21541 , RIc226890_29);
and \U$21165 ( \21542 , \21541 , \8886 );
or \U$21166 ( \21543 , \21540 , \21542 );
nand \U$21167 ( \21544 , \21543 , \2784 );
nand \U$21168 ( \21545 , \21539 , \21544 );
xor \U$21169 ( \21546 , \21536 , \21545 );
not \U$21170 ( \21547 , \2154 );
not \U$21171 ( \21548 , \20678 );
or \U$21172 ( \21549 , \21547 , \21548 );
not \U$21173 ( \21550 , RIc226980_27);
not \U$21174 ( \21551 , \9897 );
or \U$21175 ( \21552 , \21550 , \21551 );
nand \U$21176 ( \21553 , \20216 , \2799 );
nand \U$21177 ( \21554 , \21552 , \21553 );
nand \U$21178 ( \21555 , \21554 , \2138 );
nand \U$21179 ( \21556 , \21549 , \21555 );
and \U$21180 ( \21557 , \21546 , \21556 );
and \U$21181 ( \21558 , \21536 , \21545 );
or \U$21182 ( \21559 , \21557 , \21558 );
and \U$21183 ( \21560 , \21521 , \21559 );
and \U$21184 ( \21561 , \21483 , \21520 );
or \U$21185 ( \21562 , \21560 , \21561 );
not \U$21186 ( \21563 , \21562 );
or \U$21187 ( \21564 , \21481 , \21563 );
not \U$21188 ( \21565 , \21479 );
nand \U$21189 ( \21566 , \21565 , \21476 );
nand \U$21190 ( \21567 , \21564 , \21566 );
nand \U$21191 ( \21568 , \21427 , \21567 );
nand \U$21192 ( \21569 , \21426 , \21568 );
not \U$21193 ( \21570 , \21569 );
nand \U$21194 ( \21571 , \21254 , \21570 );
not \U$21195 ( \21572 , \21571 );
or \U$21196 ( \21573 , \21228 , \21572 );
nand \U$21197 ( \21574 , \21569 , \21253 );
nand \U$21198 ( \21575 , \21573 , \21574 );
not \U$21199 ( \21576 , \21575 );
xor \U$21200 ( \21577 , \21240 , \21242 );
and \U$21201 ( \21578 , \21577 , \21252 );
and \U$21202 ( \21579 , \21240 , \21242 );
or \U$21203 ( \21580 , \21578 , \21579 );
xor \U$21204 ( \21581 , \20449 , \20452 );
xor \U$21205 ( \21582 , \21581 , \20253 );
xor \U$21206 ( \21583 , \21580 , \21582 );
xor \U$21207 ( \21584 , \20298 , \20308 );
xnor \U$21208 ( \21585 , \21584 , \20296 );
not \U$21209 ( \21586 , \20249 );
not \U$21210 ( \21587 , \20243 );
or \U$21211 ( \21588 , \21586 , \21587 );
nand \U$21212 ( \21589 , \20242 , \20201 );
nand \U$21213 ( \21590 , \21588 , \21589 );
and \U$21214 ( \21591 , \21590 , \20247 );
not \U$21215 ( \21592 , \21590 );
not \U$21216 ( \21593 , \20247 );
and \U$21217 ( \21594 , \21592 , \21593 );
nor \U$21218 ( \21595 , \21591 , \21594 );
xor \U$21219 ( \21596 , \21585 , \21595 );
and \U$21220 ( \21597 , \20187 , \20161 );
not \U$21221 ( \21598 , \20187 );
and \U$21222 ( \21599 , \21598 , \20162 );
or \U$21223 ( \21600 , \21597 , \21599 );
xor \U$21224 ( \21601 , \21600 , \20172 );
xor \U$21225 ( \21602 , \20084 , \20094 );
xor \U$21226 ( \21603 , \21602 , \20105 );
or \U$21227 ( \21604 , \21601 , \21603 );
xor \U$21228 ( \21605 , \20294 , \20287 );
xnor \U$21229 ( \21606 , \21605 , \20277 );
not \U$21230 ( \21607 , \21606 );
nand \U$21231 ( \21608 , \21604 , \21607 );
nand \U$21232 ( \21609 , \21601 , \21603 );
nand \U$21233 ( \21610 , \21608 , \21609 );
and \U$21234 ( \21611 , \21596 , \21610 );
and \U$21235 ( \21612 , \21585 , \21595 );
or \U$21236 ( \21613 , \21611 , \21612 );
not \U$21237 ( \21614 , \21613 );
not \U$21238 ( \21615 , \20074 );
not \U$21239 ( \21616 , \20251 );
not \U$21240 ( \21617 , \21616 );
or \U$21241 ( \21618 , \21615 , \21617 );
not \U$21242 ( \21619 , \20248 );
not \U$21243 ( \21620 , \20250 );
or \U$21244 ( \21621 , \21619 , \21620 );
nand \U$21245 ( \21622 , \21621 , \20073 );
nand \U$21246 ( \21623 , \21618 , \21622 );
not \U$21247 ( \21624 , \20194 );
and \U$21248 ( \21625 , \21623 , \21624 );
not \U$21249 ( \21626 , \21623 );
and \U$21250 ( \21627 , \21626 , \20194 );
nor \U$21251 ( \21628 , \21625 , \21627 );
not \U$21252 ( \21629 , \21628 );
not \U$21253 ( \21630 , \21629 );
or \U$21254 ( \21631 , \21614 , \21630 );
or \U$21255 ( \21632 , \21629 , \21613 );
not \U$21256 ( \21633 , \20961 );
not \U$21257 ( \21634 , \21000 );
or \U$21258 ( \21635 , \21633 , \21634 );
or \U$21259 ( \21636 , \21000 , \20961 );
not \U$21260 ( \21637 , \20963 );
nand \U$21261 ( \21638 , \21636 , \21637 );
nand \U$21262 ( \21639 , \21635 , \21638 );
not \U$21263 ( \21640 , \21041 );
not \U$21264 ( \21641 , \21035 );
or \U$21265 ( \21642 , \21640 , \21641 );
or \U$21266 ( \21643 , \21035 , \21041 );
nand \U$21267 ( \21644 , \21643 , \21077 );
nand \U$21268 ( \21645 , \21642 , \21644 );
or \U$21269 ( \21646 , \21639 , \21645 );
xor \U$21270 ( \21647 , \20348 , \20442 );
xor \U$21271 ( \21648 , \21647 , \20439 );
nand \U$21272 ( \21649 , \21646 , \21648 );
nand \U$21273 ( \21650 , \21645 , \21639 );
nand \U$21274 ( \21651 , \21649 , \21650 );
nand \U$21275 ( \21652 , \21632 , \21651 );
nand \U$21276 ( \21653 , \21631 , \21652 );
xor \U$21277 ( \21654 , \21583 , \21653 );
not \U$21278 ( \21655 , \21654 );
not \U$21279 ( \21656 , \21655 );
or \U$21280 ( \21657 , \21576 , \21656 );
not \U$21281 ( \21658 , \21654 );
not \U$21282 ( \21659 , \21575 );
not \U$21283 ( \21660 , \21659 );
or \U$21284 ( \21661 , \21658 , \21660 );
xor \U$21285 ( \21662 , \21648 , \21645 );
xor \U$21286 ( \21663 , \21662 , \21639 );
xor \U$21287 ( \21664 , \21585 , \21595 );
xor \U$21288 ( \21665 , \21664 , \21610 );
or \U$21289 ( \21666 , \21663 , \21665 );
xor \U$21290 ( \21667 , \20848 , \20850 );
and \U$21291 ( \21668 , \21667 , \20878 );
and \U$21292 ( \21669 , \20848 , \20850 );
or \U$21293 ( \21670 , \21668 , \21669 );
not \U$21294 ( \21671 , \20147 );
not \U$21295 ( \21672 , \20189 );
or \U$21296 ( \21673 , \21671 , \21672 );
or \U$21297 ( \21674 , \20147 , \20189 );
nand \U$21298 ( \21675 , \21673 , \21674 );
buf \U$21299 ( \21676 , \20108 );
and \U$21300 ( \21677 , \21675 , \21676 );
not \U$21301 ( \21678 , \21675 );
not \U$21302 ( \21679 , \21676 );
and \U$21303 ( \21680 , \21678 , \21679 );
nor \U$21304 ( \21681 , \21677 , \21680 );
not \U$21305 ( \21682 , \21681 );
and \U$21306 ( \21683 , \21670 , \21682 );
not \U$21307 ( \21684 , \21670 );
and \U$21308 ( \21685 , \21684 , \21681 );
or \U$21309 ( \21686 , \21683 , \21685 );
xor \U$21310 ( \21687 , \20481 , \20490 );
xnor \U$21311 ( \21688 , \21687 , \20485 );
buf \U$21312 ( \21689 , \21688 );
not \U$21313 ( \21690 , \21689 );
and \U$21314 ( \21691 , \21686 , \21690 );
not \U$21315 ( \21692 , \21686 );
and \U$21316 ( \21693 , \21692 , \21689 );
nor \U$21317 ( \21694 , \21691 , \21693 );
nand \U$21318 ( \21695 , \21666 , \21694 );
nand \U$21319 ( \21696 , \21663 , \21665 );
nand \U$21320 ( \21697 , \21695 , \21696 );
not \U$21321 ( \21698 , \21613 );
not \U$21322 ( \21699 , \21628 );
not \U$21323 ( \21700 , \21651 );
and \U$21324 ( \21701 , \21699 , \21700 );
and \U$21325 ( \21702 , \21651 , \21628 );
nor \U$21326 ( \21703 , \21701 , \21702 );
not \U$21327 ( \21704 , \21703 );
or \U$21328 ( \21705 , \21698 , \21704 );
or \U$21329 ( \21706 , \21703 , \21613 );
nand \U$21330 ( \21707 , \21705 , \21706 );
xor \U$21331 ( \21708 , \21697 , \21707 );
not \U$21332 ( \21709 , \21688 );
not \U$21333 ( \21710 , \21709 );
not \U$21334 ( \21711 , \21681 );
or \U$21335 ( \21712 , \21710 , \21711 );
not \U$21336 ( \21713 , \21682 );
not \U$21337 ( \21714 , \21688 );
or \U$21338 ( \21715 , \21713 , \21714 );
nand \U$21339 ( \21716 , \21715 , \21670 );
nand \U$21340 ( \21717 , \21712 , \21716 );
not \U$21341 ( \21718 , \21717 );
xor \U$21342 ( \21719 , \20474 , \20492 );
xor \U$21343 ( \21720 , \21719 , \20495 );
not \U$21344 ( \21721 , \21720 );
and \U$21345 ( \21722 , \21718 , \21721 );
not \U$21346 ( \21723 , \21718 );
and \U$21347 ( \21724 , \21723 , \21720 );
nor \U$21348 ( \21725 , \21722 , \21724 );
xor \U$21349 ( \21726 , \20512 , \20596 );
xor \U$21350 ( \21727 , \21726 , \20803 );
not \U$21351 ( \21728 , \21727 );
and \U$21352 ( \21729 , \21725 , \21728 );
not \U$21353 ( \21730 , \21725 );
and \U$21354 ( \21731 , \21730 , \21727 );
nor \U$21355 ( \21732 , \21729 , \21731 );
and \U$21356 ( \21733 , \21708 , \21732 );
and \U$21357 ( \21734 , \21697 , \21707 );
or \U$21358 ( \21735 , \21733 , \21734 );
nand \U$21359 ( \21736 , \21661 , \21735 );
nand \U$21360 ( \21737 , \21657 , \21736 );
xor \U$21361 ( \21738 , \20842 , \21737 );
not \U$21362 ( \21739 , \21582 );
not \U$21363 ( \21740 , \21739 );
not \U$21364 ( \21741 , \21653 );
or \U$21365 ( \21742 , \21740 , \21741 );
or \U$21366 ( \21743 , \21739 , \21653 );
buf \U$21367 ( \21744 , \21580 );
nand \U$21368 ( \21745 , \21743 , \21744 );
nand \U$21369 ( \21746 , \21742 , \21745 );
not \U$21370 ( \21747 , \21746 );
not \U$21371 ( \21748 , \20458 );
not \U$21372 ( \21749 , \20063 );
or \U$21373 ( \21750 , \21748 , \21749 );
or \U$21374 ( \21751 , \20458 , \20063 );
nand \U$21375 ( \21752 , \21750 , \21751 );
not \U$21376 ( \21753 , \20500 );
and \U$21377 ( \21754 , \21752 , \21753 );
not \U$21378 ( \21755 , \21752 );
and \U$21379 ( \21756 , \21755 , \20500 );
nor \U$21380 ( \21757 , \21754 , \21756 );
and \U$21381 ( \21758 , \21747 , \21757 );
not \U$21382 ( \21759 , \21747 );
not \U$21383 ( \21760 , \21757 );
and \U$21384 ( \21761 , \21759 , \21760 );
nor \U$21385 ( \21762 , \21758 , \21761 );
not \U$21386 ( \21763 , \20465 );
not \U$21387 ( \21764 , \21763 );
not \U$21388 ( \21765 , \20469 );
or \U$21389 ( \21766 , \21764 , \21765 );
nand \U$21390 ( \21767 , \20468 , \20465 );
nand \U$21391 ( \21768 , \21766 , \21767 );
not \U$21392 ( \21769 , \20498 );
and \U$21393 ( \21770 , \21768 , \21769 );
not \U$21394 ( \21771 , \21768 );
and \U$21395 ( \21772 , \21771 , \20498 );
nor \U$21396 ( \21773 , \21770 , \21772 );
not \U$21397 ( \21774 , \21773 );
not \U$21398 ( \21775 , \21774 );
nand \U$21399 ( \21776 , \21727 , \21718 );
not \U$21400 ( \21777 , \21721 );
and \U$21401 ( \21778 , \21776 , \21777 );
nor \U$21402 ( \21779 , \21727 , \21718 );
nor \U$21403 ( \21780 , \21778 , \21779 );
not \U$21404 ( \21781 , \21780 );
not \U$21405 ( \21782 , \21781 );
or \U$21406 ( \21783 , \21775 , \21782 );
xor \U$21407 ( \21784 , \20805 , \20509 );
xor \U$21408 ( \21785 , \21784 , \20507 );
nand \U$21409 ( \21786 , \21773 , \21780 );
nand \U$21410 ( \21787 , \21785 , \21786 );
nand \U$21411 ( \21788 , \21783 , \21787 );
and \U$21412 ( \21789 , \21762 , \21788 );
not \U$21413 ( \21790 , \21762 );
not \U$21414 ( \21791 , \21788 );
and \U$21415 ( \21792 , \21790 , \21791 );
nor \U$21416 ( \21793 , \21789 , \21792 );
and \U$21417 ( \21794 , \21738 , \21793 );
and \U$21418 ( \21795 , \20842 , \21737 );
or \U$21419 ( \21796 , \21794 , \21795 );
not \U$21420 ( \21797 , \21796 );
xor \U$21421 ( \21798 , \19440 , \19479 );
xor \U$21422 ( \21799 , \21798 , \19482 );
not \U$21423 ( \21800 , \21760 );
not \U$21424 ( \21801 , \21746 );
or \U$21425 ( \21802 , \21800 , \21801 );
not \U$21426 ( \21803 , \21747 );
not \U$21427 ( \21804 , \21757 );
or \U$21428 ( \21805 , \21803 , \21804 );
nand \U$21429 ( \21806 , \21805 , \21788 );
nand \U$21430 ( \21807 , \21802 , \21806 );
xor \U$21431 ( \21808 , \21799 , \21807 );
xor \U$21432 ( \21809 , \20502 , \20504 );
xor \U$21433 ( \21810 , \21809 , \20822 );
xor \U$21434 ( \21811 , \21808 , \21810 );
not \U$21435 ( \21812 , \21811 );
or \U$21436 ( \21813 , \21797 , \21812 );
xor \U$21437 ( \21814 , \20842 , \21737 );
xor \U$21438 ( \21815 , \21814 , \21793 );
and \U$21439 ( \21816 , \21781 , \21774 );
not \U$21440 ( \21817 , \21781 );
and \U$21441 ( \21818 , \21817 , \21773 );
nor \U$21442 ( \21819 , \21816 , \21818 );
and \U$21443 ( \21820 , \21819 , \21785 );
not \U$21444 ( \21821 , \21819 );
not \U$21445 ( \21822 , \21785 );
and \U$21446 ( \21823 , \21821 , \21822 );
nor \U$21447 ( \21824 , \21820 , \21823 );
buf \U$21448 ( \21825 , \21824 );
not \U$21449 ( \21826 , \21659 );
not \U$21450 ( \21827 , \21655 );
or \U$21451 ( \21828 , \21826 , \21827 );
nand \U$21452 ( \21829 , \21654 , \21575 );
nand \U$21453 ( \21830 , \21828 , \21829 );
and \U$21454 ( \21831 , \21830 , \21735 );
not \U$21455 ( \21832 , \21830 );
not \U$21456 ( \21833 , \21735 );
and \U$21457 ( \21834 , \21832 , \21833 );
nor \U$21458 ( \21835 , \21831 , \21834 );
or \U$21459 ( \21836 , \21825 , \21835 );
xor \U$21460 ( \21837 , \21011 , \21021 );
xor \U$21461 ( \21838 , \21837 , \21032 );
xor \U$21462 ( \21839 , \21429 , \21456 );
xor \U$21463 ( \21840 , \21839 , \21473 );
xor \U$21464 ( \21841 , \21838 , \21840 );
and \U$21465 ( \21842 , \20985 , \20997 );
not \U$21466 ( \21843 , \20985 );
and \U$21467 ( \21844 , \21843 , \20996 );
or \U$21468 ( \21845 , \21842 , \21844 );
and \U$21469 ( \21846 , \21845 , \20974 );
not \U$21470 ( \21847 , \21845 );
not \U$21471 ( \21848 , \20974 );
and \U$21472 ( \21849 , \21847 , \21848 );
nor \U$21473 ( \21850 , \21846 , \21849 );
and \U$21474 ( \21851 , \21841 , \21850 );
and \U$21475 ( \21852 , \21838 , \21840 );
or \U$21476 ( \21853 , \21851 , \21852 );
not \U$21477 ( \21854 , \21607 );
not \U$21478 ( \21855 , \21603 );
not \U$21479 ( \21856 , \21855 );
or \U$21480 ( \21857 , \21854 , \21856 );
nand \U$21481 ( \21858 , \21603 , \21606 );
nand \U$21482 ( \21859 , \21857 , \21858 );
xor \U$21483 ( \21860 , \21859 , \21601 );
xor \U$21484 ( \21861 , \21853 , \21860 );
not \U$21485 ( \21862 , \2860 );
not \U$21486 ( \21863 , RIc226a70_25);
not \U$21487 ( \21864 , \11094 );
or \U$21488 ( \21865 , \21863 , \21864 );
buf \U$21489 ( \21866 , \8973 );
not \U$21490 ( \21867 , \21866 );
nand \U$21491 ( \21868 , \21867 , \1905 );
nand \U$21492 ( \21869 , \21865 , \21868 );
not \U$21493 ( \21870 , \21869 );
or \U$21494 ( \21871 , \21862 , \21870 );
nand \U$21495 ( \21872 , \21356 , \2173 );
nand \U$21496 ( \21873 , \21871 , \21872 );
not \U$21497 ( \21874 , \21873 );
not \U$21498 ( \21875 , \3631 );
not \U$21499 ( \21876 , \21502 );
or \U$21500 ( \21877 , \21875 , \21876 );
not \U$21501 ( \21878 , RIc2266b0_33);
not \U$21502 ( \21879 , \12698 );
or \U$21503 ( \21880 , \21878 , \21879 );
nand \U$21504 ( \21881 , \6492 , \6890 );
nand \U$21505 ( \21882 , \21880 , \21881 );
nand \U$21506 ( \21883 , \21882 , \3629 );
nand \U$21507 ( \21884 , \21877 , \21883 );
not \U$21508 ( \21885 , \21884 );
nand \U$21509 ( \21886 , \21874 , \21885 );
not \U$21510 ( \21887 , \4381 );
not \U$21511 ( \21888 , RIc2265c0_35);
not \U$21512 ( \21889 , \5664 );
or \U$21513 ( \21890 , \21888 , \21889 );
nand \U$21514 ( \21891 , \6726 , \4376 );
nand \U$21515 ( \21892 , \21890 , \21891 );
not \U$21516 ( \21893 , \21892 );
or \U$21517 ( \21894 , \21887 , \21893 );
nand \U$21518 ( \21895 , \21371 , \4383 );
nand \U$21519 ( \21896 , \21894 , \21895 );
and \U$21520 ( \21897 , \21886 , \21896 );
nor \U$21521 ( \21898 , \21874 , \21885 );
nor \U$21522 ( \21899 , \21897 , \21898 );
not \U$21523 ( \21900 , \21899 );
not \U$21524 ( \21901 , \21900 );
not \U$21525 ( \21902 , \2138 );
not \U$21526 ( \21903 , RIc226980_27);
not \U$21527 ( \21904 , \8807 );
or \U$21528 ( \21905 , \21903 , \21904 );
nand \U$21529 ( \21906 , \10859 , \16510 );
nand \U$21530 ( \21907 , \21905 , \21906 );
not \U$21531 ( \21908 , \21907 );
or \U$21532 ( \21909 , \21902 , \21908 );
nand \U$21533 ( \21910 , \21554 , \2154 );
nand \U$21534 ( \21911 , \21909 , \21910 );
not \U$21535 ( \21912 , \21911 );
and \U$21536 ( \21913 , \21489 , \1930 );
and \U$21537 ( \21914 , RIc226b60_23, \13129 );
not \U$21538 ( \21915 , RIc226b60_23);
and \U$21539 ( \21916 , \21915 , \8924 );
or \U$21540 ( \21917 , \21914 , \21916 );
and \U$21541 ( \21918 , \21917 , \1915 );
nor \U$21542 ( \21919 , \21913 , \21918 );
not \U$21543 ( \21920 , \21919 );
not \U$21544 ( \21921 , \21920 );
or \U$21545 ( \21922 , \21912 , \21921 );
not \U$21546 ( \21923 , \21919 );
not \U$21547 ( \21924 , \21911 );
not \U$21548 ( \21925 , \21924 );
or \U$21549 ( \21926 , \21923 , \21925 );
not \U$21550 ( \21927 , \5519 );
not \U$21551 ( \21928 , \21516 );
or \U$21552 ( \21929 , \21927 , \21928 );
not \U$21553 ( \21930 , RIc2264d0_37);
not \U$21554 ( \21931 , \10220 );
or \U$21555 ( \21932 , \21930 , \21931 );
nand \U$21556 ( \21933 , \4406 , \4371 );
nand \U$21557 ( \21934 , \21932 , \21933 );
nand \U$21558 ( \21935 , \21934 , \5509 );
nand \U$21559 ( \21936 , \21929 , \21935 );
nand \U$21560 ( \21937 , \21926 , \21936 );
nand \U$21561 ( \21938 , \21922 , \21937 );
not \U$21562 ( \21939 , \21938 );
or \U$21563 ( \21940 , \21901 , \21939 );
not \U$21564 ( \21941 , \21938 );
not \U$21565 ( \21942 , \21941 );
not \U$21566 ( \21943 , \21899 );
or \U$21567 ( \21944 , \21942 , \21943 );
or \U$21568 ( \21945 , RIc227178_10, RIc227100_11);
nand \U$21569 ( \21946 , \21945 , \16248 );
and \U$21570 ( \21947 , RIc227178_10, RIc227100_11);
nor \U$21571 ( \21948 , \21947 , \1351 );
and \U$21572 ( \21949 , \21946 , \21948 );
not \U$21573 ( \21950 , \1339 );
not \U$21574 ( \21951 , \21106 );
or \U$21575 ( \21952 , \21950 , \21951 );
or \U$21576 ( \21953 , \18367 , \1342 );
not \U$21577 ( \21954 , \16248 );
or \U$21578 ( \21955 , \21954 , RIc2271f0_9);
nand \U$21579 ( \21956 , \21953 , \21955 );
nand \U$21580 ( \21957 , \21956 , \1362 );
nand \U$21581 ( \21958 , \21952 , \21957 );
and \U$21582 ( \21959 , \21949 , \21958 );
not \U$21583 ( \21960 , \1678 );
and \U$21584 ( \21961 , RIc227010_13, \13198 );
not \U$21585 ( \21962 , RIc227010_13);
and \U$21586 ( \21963 , \21962 , \12755 );
or \U$21587 ( \21964 , \21961 , \21963 );
not \U$21588 ( \21965 , \21964 );
or \U$21589 ( \21966 , \21960 , \21965 );
nand \U$21590 ( \21967 , \21088 , \1682 );
nand \U$21591 ( \21968 , \21966 , \21967 );
xor \U$21592 ( \21969 , \21959 , \21968 );
not \U$21593 ( \21970 , \2318 );
not \U$21594 ( \21971 , \21177 );
or \U$21595 ( \21972 , \21970 , \21971 );
not \U$21596 ( \21973 , RIc226f20_15);
not \U$21597 ( \21974 , \10198 );
or \U$21598 ( \21975 , \21973 , \21974 );
not \U$21599 ( \21976 , \10198 );
nand \U$21600 ( \21977 , \21976 , \2301 );
nand \U$21601 ( \21978 , \21975 , \21977 );
nand \U$21602 ( \21979 , \21978 , \2320 );
nand \U$21603 ( \21980 , \21972 , \21979 );
and \U$21604 ( \21981 , \21969 , \21980 );
and \U$21605 ( \21982 , \21959 , \21968 );
or \U$21606 ( \21983 , \21981 , \21982 );
not \U$21607 ( \21984 , \2697 );
not \U$21608 ( \21985 , RIc2267a0_31);
not \U$21609 ( \21986 , \10142 );
or \U$21610 ( \21987 , \21985 , \21986 );
nand \U$21611 ( \21988 , \10310 , \2705 );
nand \U$21612 ( \21989 , \21987 , \21988 );
not \U$21613 ( \21990 , \21989 );
or \U$21614 ( \21991 , \21984 , \21990 );
nand \U$21615 ( \21992 , \21442 , \2710 );
nand \U$21616 ( \21993 , \21991 , \21992 );
xor \U$21617 ( \21994 , \21983 , \21993 );
not \U$21618 ( \21995 , \2784 );
and \U$21619 ( \21996 , RIc226890_29, \12724 );
not \U$21620 ( \21997 , RIc226890_29);
and \U$21621 ( \21998 , \21997 , \12727 );
or \U$21622 ( \21999 , \21996 , \21998 );
not \U$21623 ( \22000 , \21999 );
or \U$21624 ( \22001 , \21995 , \22000 );
nand \U$21625 ( \22002 , \21543 , \9142 );
nand \U$21626 ( \22003 , \22001 , \22002 );
and \U$21627 ( \22004 , \21994 , \22003 );
and \U$21628 ( \22005 , \21983 , \21993 );
or \U$21629 ( \22006 , \22004 , \22005 );
nand \U$21630 ( \22007 , \21944 , \22006 );
nand \U$21631 ( \22008 , \21940 , \22007 );
not \U$21632 ( \22009 , \22008 );
xor \U$21633 ( \22010 , \21483 , \21520 );
xor \U$21634 ( \22011 , \22010 , \21559 );
not \U$21635 ( \22012 , \22011 );
or \U$21636 ( \22013 , \22009 , \22012 );
not \U$21637 ( \22014 , \22008 );
not \U$21638 ( \22015 , \22014 );
not \U$21639 ( \22016 , \22011 );
not \U$21640 ( \22017 , \22016 );
or \U$21641 ( \22018 , \22015 , \22017 );
xor \U$21642 ( \22019 , \21536 , \21545 );
xor \U$21643 ( \22020 , \22019 , \21556 );
xor \U$21644 ( \22021 , \21493 , \21504 );
xor \U$21645 ( \22022 , \22021 , \21518 );
xor \U$21646 ( \22023 , \22020 , \22022 );
not \U$21647 ( \22024 , \9934 );
not \U$21648 ( \22025 , RIc226110_45);
not \U$21649 ( \22026 , \11841 );
or \U$21650 ( \22027 , \22025 , \22026 );
nand \U$21651 ( \22028 , \2064 , \9100 );
nand \U$21652 ( \22029 , \22027 , \22028 );
not \U$21653 ( \22030 , \22029 );
or \U$21654 ( \22031 , \22024 , \22030 );
nand \U$21655 ( \22032 , \21384 , \9398 );
nand \U$21656 ( \22033 , \22031 , \22032 );
not \U$21657 ( \22034 , \22033 );
not \U$21658 ( \22035 , \22034 );
not \U$21659 ( \22036 , \11974 );
not \U$21660 ( \22037 , \20892 );
or \U$21661 ( \22038 , \22036 , \22037 );
not \U$21662 ( \22039 , RIc225b70_57);
not \U$21663 ( \22040 , \10930 );
or \U$21664 ( \22041 , \22039 , \22040 );
nand \U$21665 ( \22042 , \8989 , \10074 );
nand \U$21666 ( \22043 , \22041 , \22042 );
nand \U$21667 ( \22044 , \22043 , \11965 );
nand \U$21668 ( \22045 , \22038 , \22044 );
not \U$21669 ( \22046 , \22045 );
not \U$21670 ( \22047 , \22046 );
or \U$21671 ( \22048 , \22035 , \22047 );
not \U$21672 ( \22049 , \9619 );
not \U$21673 ( \22050 , \20924 );
or \U$21674 ( \22051 , \22049 , \22050 );
and \U$21675 ( \22052 , RIc226020_47, \11854 );
not \U$21676 ( \22053 , RIc226020_47);
and \U$21677 ( \22054 , \22053 , \2498 );
or \U$21678 ( \22055 , \22052 , \22054 );
nand \U$21679 ( \22056 , \22055 , \10001 );
nand \U$21680 ( \22057 , \22051 , \22056 );
nand \U$21681 ( \22058 , \22048 , \22057 );
nand \U$21682 ( \22059 , \22033 , \22045 );
nand \U$21683 ( \22060 , \22058 , \22059 );
and \U$21684 ( \22061 , \22023 , \22060 );
and \U$21685 ( \22062 , \22020 , \22022 );
or \U$21686 ( \22063 , \22061 , \22062 );
nand \U$21687 ( \22064 , \22018 , \22063 );
nand \U$21688 ( \22065 , \22013 , \22064 );
and \U$21689 ( \22066 , \21861 , \22065 );
and \U$21690 ( \22067 , \21853 , \21860 );
or \U$21691 ( \22068 , \22066 , \22067 );
not \U$21692 ( \22069 , \22068 );
xor \U$21693 ( \22070 , \21256 , \21567 );
not \U$21694 ( \22071 , \21424 );
and \U$21695 ( \22072 , \22070 , \22071 );
not \U$21696 ( \22073 , \22070 );
and \U$21697 ( \22074 , \22073 , \21424 );
nor \U$21698 ( \22075 , \22072 , \22074 );
not \U$21699 ( \22076 , \22075 );
not \U$21700 ( \22077 , \22076 );
or \U$21701 ( \22078 , \22069 , \22077 );
not \U$21702 ( \22079 , \22068 );
not \U$21703 ( \22080 , \22079 );
not \U$21704 ( \22081 , \22075 );
or \U$21705 ( \22082 , \22080 , \22081 );
xor \U$21706 ( \22083 , \21476 , \21565 );
xnor \U$21707 ( \22084 , \22083 , \21562 );
not \U$21708 ( \22085 , \22084 );
xor \U$21709 ( \22086 , \21259 , \21337 );
xnor \U$21710 ( \22087 , \22086 , \21422 );
not \U$21711 ( \22088 , \22087 );
or \U$21712 ( \22089 , \22085 , \22088 );
xor \U$21713 ( \22090 , \21526 , \21527 );
xor \U$21714 ( \22091 , \22090 , \21533 );
not \U$21715 ( \22092 , \9552 );
not \U$21716 ( \22093 , \20908 );
or \U$21717 ( \22094 , \22092 , \22093 );
not \U$21718 ( \22095 , RIc225f30_49);
not \U$21719 ( \22096 , \9361 );
or \U$21720 ( \22097 , \22095 , \22096 );
nand \U$21721 ( \22098 , \10899 , \11289 );
nand \U$21722 ( \22099 , \22097 , \22098 );
nand \U$21723 ( \22100 , \22099 , \10445 );
nand \U$21724 ( \22101 , \22094 , \22100 );
xor \U$21725 ( \22102 , \22091 , \22101 );
not \U$21726 ( \22103 , \15719 );
not \U$21727 ( \22104 , RIc225990_61);
not \U$21728 ( \22105 , \1949 );
or \U$21729 ( \22106 , \22104 , \22105 );
nand \U$21730 ( \22107 , \3439 , \12806 );
nand \U$21731 ( \22108 , \22106 , \22107 );
not \U$21732 ( \22109 , \22108 );
or \U$21733 ( \22110 , \22103 , \22109 );
nand \U$21734 ( \22111 , \21345 , \20862 );
nand \U$21735 ( \22112 , \22110 , \22111 );
and \U$21736 ( \22113 , \22102 , \22112 );
and \U$21737 ( \22114 , \22091 , \22101 );
or \U$21738 ( \22115 , \22113 , \22114 );
xor \U$21739 ( \22116 , \21459 , \21464 );
xor \U$21740 ( \22117 , \22116 , \21470 );
not \U$21741 ( \22118 , \22117 );
xor \U$21742 ( \22119 , \21434 , \21454 );
xnor \U$21743 ( \22120 , \21446 , \22119 );
nand \U$21744 ( \22121 , \22118 , \22120 );
nand \U$21745 ( \22122 , \22115 , \22121 );
not \U$21746 ( \22123 , \22120 );
nand \U$21747 ( \22124 , \22123 , \22117 );
nand \U$21748 ( \22125 , \22122 , \22124 );
not \U$21749 ( \22126 , \6307 );
not \U$21750 ( \22127 , \21271 );
or \U$21751 ( \22128 , \22126 , \22127 );
not \U$21752 ( \22129 , RIc2263e0_39);
not \U$21753 ( \22130 , \14299 );
or \U$21754 ( \22131 , \22129 , \22130 );
nand \U$21755 ( \22132 , \3640 , \5498 );
nand \U$21756 ( \22133 , \22131 , \22132 );
nand \U$21757 ( \22134 , \22133 , \6689 );
nand \U$21758 ( \22135 , \22128 , \22134 );
not \U$21759 ( \22136 , \9459 );
not \U$21760 ( \22137 , RIc225e40_51);
not \U$21761 ( \22138 , \3509 );
or \U$21762 ( \22139 , \22137 , \22138 );
not \U$21763 ( \22140 , RIc225e40_51);
nand \U$21764 ( \22141 , \9434 , \22140 );
nand \U$21765 ( \22142 , \22139 , \22141 );
not \U$21766 ( \22143 , \22142 );
or \U$21767 ( \22144 , \22136 , \22143 );
nand \U$21768 ( \22145 , \21325 , \9444 );
nand \U$21769 ( \22146 , \22144 , \22145 );
xor \U$21770 ( \22147 , \22135 , \22146 );
not \U$21771 ( \22148 , \9488 );
not \U$21772 ( \22149 , RIc225d50_53);
not \U$21773 ( \22150 , \2257 );
or \U$21774 ( \22151 , \22149 , \22150 );
nand \U$21775 ( \22152 , \9608 , \8772 );
nand \U$21776 ( \22153 , \22151 , \22152 );
not \U$21777 ( \22154 , \22153 );
or \U$21778 ( \22155 , \22148 , \22154 );
nand \U$21779 ( \22156 , \21297 , \12945 );
nand \U$21780 ( \22157 , \22155 , \22156 );
and \U$21781 ( \22158 , \22147 , \22157 );
and \U$21782 ( \22159 , \22135 , \22146 );
or \U$21783 ( \22160 , \22158 , \22159 );
not \U$21784 ( \22161 , \21373 );
not \U$21785 ( \22162 , \21361 );
or \U$21786 ( \22163 , \22161 , \22162 );
or \U$21787 ( \22164 , \21361 , \21373 );
nand \U$21788 ( \22165 , \22163 , \22164 );
and \U$21789 ( \22166 , \22165 , \21349 );
not \U$21790 ( \22167 , \22165 );
and \U$21791 ( \22168 , \22167 , \21350 );
nor \U$21792 ( \22169 , \22166 , \22168 );
xor \U$21793 ( \22170 , \22160 , \22169 );
not \U$21794 ( \22171 , \11118 );
not \U$21795 ( \22172 , RIc225c60_55);
not \U$21796 ( \22173 , \2834 );
or \U$21797 ( \22174 , \22172 , \22173 );
nand \U$21798 ( \22175 , \5269 , \11108 );
nand \U$21799 ( \22176 , \22174 , \22175 );
not \U$21800 ( \22177 , \22176 );
or \U$21801 ( \22178 , \22171 , \22177 );
nand \U$21802 ( \22179 , \21394 , \13025 );
nand \U$21803 ( \22180 , \22178 , \22179 );
not \U$21804 ( \22181 , \9705 );
not \U$21805 ( \22182 , \21283 );
or \U$21806 ( \22183 , \22181 , \22182 );
and \U$21807 ( \22184 , RIc2262f0_41, \11321 );
not \U$21808 ( \22185 , RIc2262f0_41);
and \U$21809 ( \22186 , \22185 , \11324 );
or \U$21810 ( \22187 , \22184 , \22186 );
nand \U$21811 ( \22188 , \22187 , \9690 );
nand \U$21812 ( \22189 , \22183 , \22188 );
xor \U$21813 ( \22190 , \22180 , \22189 );
not \U$21814 ( \22191 , \9205 );
not \U$21815 ( \22192 , \21405 );
or \U$21816 ( \22193 , \22191 , \22192 );
not \U$21817 ( \22194 , RIc226200_43);
not \U$21818 ( \22195 , \4228 );
or \U$21819 ( \22196 , \22194 , \22195 );
not \U$21820 ( \22197 , \2635 );
nand \U$21821 ( \22198 , \22197 , \9106 );
nand \U$21822 ( \22199 , \22196 , \22198 );
nand \U$21823 ( \22200 , \22199 , \9110 );
nand \U$21824 ( \22201 , \22193 , \22200 );
and \U$21825 ( \22202 , \22190 , \22201 );
and \U$21826 ( \22203 , \22180 , \22189 );
or \U$21827 ( \22204 , \22202 , \22203 );
and \U$21828 ( \22205 , \22170 , \22204 );
and \U$21829 ( \22206 , \22160 , \22169 );
or \U$21830 ( \22207 , \22205 , \22206 );
xor \U$21831 ( \22208 , \22125 , \22207 );
xor \U$21832 ( \22209 , \20886 , \20929 );
xor \U$21833 ( \22210 , \22209 , \20952 );
and \U$21834 ( \22211 , \22208 , \22210 );
and \U$21835 ( \22212 , \22125 , \22207 );
or \U$21836 ( \22213 , \22211 , \22212 );
nand \U$21837 ( \22214 , \22089 , \22213 );
not \U$21838 ( \22215 , \22084 );
not \U$21839 ( \22216 , \22087 );
nand \U$21840 ( \22217 , \22215 , \22216 );
nand \U$21841 ( \22218 , \22214 , \22217 );
nand \U$21842 ( \22219 , \22082 , \22218 );
nand \U$21843 ( \22220 , \22078 , \22219 );
not \U$21844 ( \22221 , \22220 );
and \U$21845 ( \22222 , \21253 , \21569 );
not \U$21846 ( \22223 , \21253 );
and \U$21847 ( \22224 , \22223 , \21570 );
nor \U$21848 ( \22225 , \22222 , \22224 );
xnor \U$21849 ( \22226 , \22225 , \21227 );
nand \U$21850 ( \22227 , \22221 , \22226 );
not \U$21851 ( \22228 , \22227 );
xor \U$21852 ( \22229 , \21697 , \21707 );
xor \U$21853 ( \22230 , \22229 , \21732 );
not \U$21854 ( \22231 , \22230 );
or \U$21855 ( \22232 , \22228 , \22231 );
not \U$21856 ( \22233 , \22226 );
nand \U$21857 ( \22234 , \22233 , \22220 );
nand \U$21858 ( \22235 , \22232 , \22234 );
nand \U$21859 ( \22236 , \21836 , \22235 );
nand \U$21860 ( \22237 , \21835 , \21825 );
nand \U$21861 ( \22238 , \22236 , \22237 );
nand \U$21862 ( \22239 , \21815 , \22238 );
nand \U$21863 ( \22240 , \21813 , \22239 );
not \U$21864 ( \22241 , \21811 );
not \U$21865 ( \22242 , \21796 );
nand \U$21866 ( \22243 , \22241 , \22242 );
nand \U$21867 ( \22244 , \22240 , \22243 );
not \U$21868 ( \22245 , \20825 );
xor \U$21869 ( \22246 , \20040 , \22245 );
xnor \U$21870 ( \22247 , \22246 , \20052 );
xor \U$21871 ( \22248 , \21799 , \21807 );
and \U$21872 ( \22249 , \22248 , \21810 );
and \U$21873 ( \22250 , \21799 , \21807 );
or \U$21874 ( \22251 , \22249 , \22250 );
nor \U$21875 ( \22252 , \22247 , \22251 );
or \U$21876 ( \22253 , \22244 , \22252 );
nand \U$21877 ( \22254 , \22247 , \22251 );
nand \U$21878 ( \22255 , \22253 , \22254 );
not \U$21879 ( \22256 , \22255 );
or \U$21880 ( \22257 , \20832 , \22256 );
not \U$21881 ( \22258 , \20038 );
not \U$21882 ( \22259 , \20830 );
nand \U$21883 ( \22260 , \22258 , \22259 );
nand \U$21884 ( \22261 , \22257 , \22260 );
buf \U$21885 ( \22262 , \20004 );
nand \U$21886 ( \22263 , \19435 , \19995 );
and \U$21887 ( \22264 , \22262 , \22263 , \20023 , \18889 );
nand \U$21888 ( \22265 , \22261 , \22264 );
nand \U$21889 ( \22266 , \20027 , \22265 );
not \U$21890 ( \22267 , \22266 );
or \U$21891 ( \22268 , \17459 , \22267 );
not \U$21892 ( \22269 , \15100 );
not \U$21893 ( \22270 , \17456 );
not \U$21894 ( \22271 , \16737 );
not \U$21895 ( \22272 , \16197 );
or \U$21896 ( \22273 , \22271 , \22272 );
nand \U$21897 ( \22274 , \16742 , \17444 );
nand \U$21898 ( \22275 , \22273 , \22274 );
nand \U$21899 ( \22276 , \22275 , \16739 );
or \U$21900 ( \22277 , \22276 , \16194 );
nand \U$21901 ( \22278 , \15572 , \16193 );
nand \U$21902 ( \22279 , \22277 , \22278 );
not \U$21903 ( \22280 , \22279 );
or \U$21904 ( \22281 , \22270 , \22280 );
not \U$21905 ( \22282 , \17455 );
not \U$21906 ( \22283 , \17453 );
nand \U$21907 ( \22284 , \22282 , \22283 );
nand \U$21908 ( \22285 , \22281 , \22284 );
not \U$21909 ( \22286 , \22285 );
or \U$21910 ( \22287 , \22269 , \22286 );
not \U$21911 ( \22288 , \15098 );
not \U$21912 ( \22289 , \14092 );
nand \U$21913 ( \22290 , \12921 , \13559 );
or \U$21914 ( \22291 , \22289 , \22290 );
not \U$21915 ( \22292 , \14091 );
buf \U$21916 ( \22293 , \14085 );
nand \U$21917 ( \22294 , \22292 , \22293 );
nand \U$21918 ( \22295 , \22291 , \22294 );
not \U$21919 ( \22296 , \22295 );
or \U$21920 ( \22297 , \22288 , \22296 );
not \U$21921 ( \22298 , \15097 );
nand \U$21922 ( \22299 , \22298 , \15094 );
nand \U$21923 ( \22300 , \22297 , \22299 );
buf \U$21924 ( \22301 , \15090 );
and \U$21925 ( \22302 , \22300 , \22301 );
nor \U$21926 ( \22303 , \14583 , \15089 );
nor \U$21927 ( \22304 , \22302 , \22303 );
nand \U$21928 ( \22305 , \22287 , \22304 );
not \U$21929 ( \22306 , \22305 );
nand \U$21930 ( \22307 , \22268 , \22306 );
not \U$21931 ( \22308 , \5509 );
not \U$21932 ( \22309 , RIc2264d0_37);
not \U$21933 ( \22310 , \1530 );
or \U$21934 ( \22311 , \22309 , \22310 );
nand \U$21935 ( \22312 , \3579 , \12522 );
nand \U$21936 ( \22313 , \22311 , \22312 );
not \U$21937 ( \22314 , \22313 );
or \U$21938 ( \22315 , \22308 , \22314 );
not \U$21939 ( \22316 , RIc2264d0_37);
not \U$21940 ( \22317 , \3496 );
or \U$21941 ( \22318 , \22316 , \22317 );
not \U$21942 ( \22319 , \2380 );
nand \U$21943 ( \22320 , \22319 , \4371 );
nand \U$21944 ( \22321 , \22318 , \22320 );
nand \U$21945 ( \22322 , \22321 , \5519 );
nand \U$21946 ( \22323 , \22315 , \22322 );
not \U$21947 ( \22324 , \22323 );
not \U$21948 ( \22325 , \2860 );
not \U$21949 ( \22326 , RIc226a70_25);
not \U$21950 ( \22327 , \2592 );
or \U$21951 ( \22328 , \22326 , \22327 );
not \U$21952 ( \22329 , \2591 );
nand \U$21953 ( \22330 , \22329 , \1905 );
nand \U$21954 ( \22331 , \22328 , \22330 );
not \U$21955 ( \22332 , \22331 );
or \U$21956 ( \22333 , \22325 , \22332 );
not \U$21957 ( \22334 , RIc226a70_25);
not \U$21958 ( \22335 , \2015 );
or \U$21959 ( \22336 , \22334 , \22335 );
nand \U$21960 ( \22337 , \3508 , \13838 );
nand \U$21961 ( \22338 , \22336 , \22337 );
nand \U$21962 ( \22339 , \22338 , \2173 );
nand \U$21963 ( \22340 , \22333 , \22339 );
not \U$21964 ( \22341 , \22340 );
not \U$21965 ( \22342 , \22341 );
or \U$21966 ( \22343 , \22324 , \22342 );
not \U$21967 ( \22344 , \22323 );
nand \U$21968 ( \22345 , \22344 , \22340 );
nand \U$21969 ( \22346 , \22343 , \22345 );
not \U$21970 ( \22347 , \9110 );
not \U$21971 ( \22348 , RIc226200_43);
not \U$21972 ( \22349 , \10450 );
or \U$21973 ( \22350 , \22348 , \22349 );
nand \U$21974 ( \22351 , \840 , \9125 );
nand \U$21975 ( \22352 , \22350 , \22351 );
not \U$21976 ( \22353 , \22352 );
or \U$21977 ( \22354 , \22347 , \22353 );
not \U$21978 ( \22355 , RIc226200_43);
not \U$21979 ( \22356 , \13077 );
or \U$21980 ( \22357 , \22355 , \22356 );
nand \U$21981 ( \22358 , \888 , \9117 );
nand \U$21982 ( \22359 , \22357 , \22358 );
nand \U$21983 ( \22360 , \22359 , \9205 );
nand \U$21984 ( \22361 , \22354 , \22360 );
not \U$21985 ( \22362 , \22361 );
and \U$21986 ( \22363 , \22346 , \22362 );
not \U$21987 ( \22364 , \22346 );
and \U$21988 ( \22365 , \22364 , \22361 );
nor \U$21989 ( \22366 , \22363 , \22365 );
not \U$21990 ( \22367 , \22366 );
not \U$21991 ( \22368 , \22367 );
not \U$21992 ( \22369 , \4383 );
not \U$21993 ( \22370 , RIc2265c0_35);
not \U$21994 ( \22371 , \3438 );
or \U$21995 ( \22372 , \22370 , \22371 );
nand \U$21996 ( \22373 , \3439 , \4376 );
nand \U$21997 ( \22374 , \22372 , \22373 );
not \U$21998 ( \22375 , \22374 );
or \U$21999 ( \22376 , \22369 , \22375 );
and \U$22000 ( \22377 , \1485 , \3620 );
not \U$22001 ( \22378 , \1485 );
and \U$22002 ( \22379 , \22378 , RIc2265c0_35);
or \U$22003 ( \22380 , \22377 , \22379 );
nand \U$22004 ( \22381 , \22380 , \4381 );
nand \U$22005 ( \22382 , \22376 , \22381 );
not \U$22006 ( \22383 , \1930 );
not \U$22007 ( \22384 , RIc226b60_23);
not \U$22008 ( \22385 , \9361 );
or \U$22009 ( \22386 , \22384 , \22385 );
not \U$22010 ( \22387 , RIc226b60_23);
not \U$22011 ( \22388 , \15908 );
nand \U$22012 ( \22389 , \22387 , \22388 );
nand \U$22013 ( \22390 , \22386 , \22389 );
not \U$22014 ( \22391 , \22390 );
or \U$22015 ( \22392 , \22383 , \22391 );
not \U$22016 ( \22393 , RIc226b60_23);
not \U$22017 ( \22394 , \2476 );
or \U$22018 ( \22395 , \22393 , \22394 );
nand \U$22019 ( \22396 , \3036 , \1927 );
nand \U$22020 ( \22397 , \22395 , \22396 );
nand \U$22021 ( \22398 , \22397 , \1915 );
nand \U$22022 ( \22399 , \22392 , \22398 );
not \U$22023 ( \22400 , \22399 );
and \U$22024 ( \22401 , \22382 , \22400 );
not \U$22025 ( \22402 , \22382 );
and \U$22026 ( \22403 , \22402 , \22399 );
or \U$22027 ( \22404 , \22401 , \22403 );
not \U$22028 ( \22405 , RIc226c50_21);
not \U$22029 ( \22406 , \3022 );
or \U$22030 ( \22407 , \22405 , \22406 );
not \U$22031 ( \22408 , \11854 );
nand \U$22032 ( \22409 , \22408 , \2383 );
nand \U$22033 ( \22410 , \22407 , \22409 );
and \U$22034 ( \22411 , \22410 , \2367 );
not \U$22035 ( \22412 , RIc226c50_21);
not \U$22036 ( \22413 , \2670 );
or \U$22037 ( \22414 , \22412 , \22413 );
nand \U$22038 ( \22415 , \4564 , \2370 );
nand \U$22039 ( \22416 , \22414 , \22415 );
and \U$22040 ( \22417 , \22416 , \2392 );
nor \U$22041 ( \22418 , \22411 , \22417 );
buf \U$22042 ( \22419 , \22418 );
and \U$22043 ( \22420 , \22404 , \22419 );
not \U$22044 ( \22421 , \22404 );
not \U$22045 ( \22422 , \22419 );
and \U$22046 ( \22423 , \22421 , \22422 );
nor \U$22047 ( \22424 , \22420 , \22423 );
not \U$22048 ( \22425 , \22424 );
not \U$22049 ( \22426 , \22425 );
or \U$22050 ( \22427 , \22368 , \22426 );
not \U$22051 ( \22428 , \22424 );
not \U$22052 ( \22429 , \22366 );
or \U$22053 ( \22430 , \22428 , \22429 );
and \U$22054 ( \22431 , RIc226890_29, \2225 );
not \U$22055 ( \22432 , RIc226890_29);
and \U$22056 ( \22433 , \22432 , \2233 );
or \U$22057 ( \22434 , \22431 , \22433 );
not \U$22058 ( \22435 , \22434 );
not \U$22059 ( \22436 , \9142 );
not \U$22060 ( \22437 , \22436 );
and \U$22061 ( \22438 , \22435 , \22437 );
and \U$22062 ( \22439 , RIc226890_29, \4009 );
not \U$22063 ( \22440 , RIc226890_29);
and \U$22064 ( \22441 , \22440 , \4008 );
or \U$22065 ( \22442 , \22439 , \22441 );
and \U$22066 ( \22443 , \22442 , \2784 );
nor \U$22067 ( \22444 , \22438 , \22443 );
not \U$22068 ( \22445 , \22444 );
not \U$22069 ( \22446 , \22445 );
not \U$22070 ( \22447 , \2697 );
not \U$22071 ( \22448 , RIc2267a0_31);
not \U$22072 ( \22449 , \9570 );
or \U$22073 ( \22450 , \22448 , \22449 );
nand \U$22074 ( \22451 , \5269 , \2705 );
nand \U$22075 ( \22452 , \22450 , \22451 );
not \U$22076 ( \22453 , \22452 );
or \U$22077 ( \22454 , \22447 , \22453 );
not \U$22078 ( \22455 , RIc2267a0_31);
not \U$22079 ( \22456 , \9479 );
or \U$22080 ( \22457 , \22455 , \22456 );
nand \U$22081 ( \22458 , \2422 , \2705 );
nand \U$22082 ( \22459 , \22457 , \22458 );
nand \U$22083 ( \22460 , \2711 , \22459 );
nand \U$22084 ( \22461 , \22454 , \22460 );
not \U$22085 ( \22462 , \22461 );
or \U$22086 ( \22463 , \22446 , \22462 );
or \U$22087 ( \22464 , \22461 , \22445 );
not \U$22088 ( \22465 , \9705 );
not \U$22089 ( \22466 , \11715 );
not \U$22090 ( \22467 , \9822 );
or \U$22091 ( \22468 , \22466 , \22467 );
not \U$22092 ( \22469 , \1020 );
nand \U$22093 ( \22470 , \22469 , RIc2262f0_41);
nand \U$22094 ( \22471 , \22468 , \22470 );
not \U$22095 ( \22472 , \22471 );
or \U$22096 ( \22473 , \22465 , \22472 );
not \U$22097 ( \22474 , RIc2262f0_41);
not \U$22098 ( \22475 , \11260 );
or \U$22099 ( \22476 , \22474 , \22475 );
nand \U$22100 ( \22477 , \9540 , \6303 );
nand \U$22101 ( \22478 , \22476 , \22477 );
nand \U$22102 ( \22479 , \22478 , \9690 );
nand \U$22103 ( \22480 , \22473 , \22479 );
nand \U$22104 ( \22481 , \22464 , \22480 );
nand \U$22105 ( \22482 , \22463 , \22481 );
nand \U$22106 ( \22483 , \22430 , \22482 );
nand \U$22107 ( \22484 , \22427 , \22483 );
not \U$22108 ( \22485 , \22484 );
not \U$22109 ( \22486 , \9934 );
not \U$22110 ( \22487 , RIc226110_45);
not \U$22111 ( \22488 , \11112 );
or \U$22112 ( \22489 , \22487 , \22488 );
nand \U$22113 ( \22490 , \3957 , \9379 );
nand \U$22114 ( \22491 , \22489 , \22490 );
not \U$22115 ( \22492 , \22491 );
or \U$22116 ( \22493 , \22486 , \22492 );
nand \U$22117 ( \22494 , \11825 , RIc226110_45);
nand \U$22118 ( \22495 , \22493 , \22494 );
not \U$22119 ( \22496 , \1082 );
not \U$22120 ( \22497 , \1078 );
not \U$22121 ( \22498 , \16532 );
or \U$22122 ( \22499 , \22497 , \22498 );
not \U$22123 ( \22500 , \16532 );
nand \U$22124 ( \22501 , \22500 , RIc2274c0_3);
nand \U$22125 ( \22502 , \22499 , \22501 );
not \U$22126 ( \22503 , \22502 );
or \U$22127 ( \22504 , \22496 , \22503 );
and \U$22128 ( \22505 , \12727 , \1027 );
not \U$22129 ( \22506 , \12727 );
and \U$22130 ( \22507 , \22506 , RIc2274c0_3);
or \U$22131 ( \22508 , \22505 , \22507 );
nand \U$22132 ( \22509 , \22508 , \1040 );
nand \U$22133 ( \22510 , \22504 , \22509 );
xor \U$22134 ( \22511 , \22495 , \22510 );
and \U$22135 ( \22512 , RIc2275b0_1, \8807 );
not \U$22136 ( \22513 , RIc2275b0_1);
and \U$22137 ( \22514 , \22513 , \8811 );
nor \U$22138 ( \22515 , \22512 , \22514 );
or \U$22139 ( \22516 , \22515 , \855 );
xor \U$22140 ( \22517 , RIc2275b0_1, \20216 );
not \U$22141 ( \22518 , \22517 );
or \U$22142 ( \22519 , \22518 , \899 );
nand \U$22143 ( \22520 , \22516 , \22519 );
xor \U$22144 ( \22521 , \22511 , \22520 );
not \U$22145 ( \22522 , \3629 );
not \U$22146 ( \22523 , RIc2266b0_33);
not \U$22147 ( \22524 , \9700 );
or \U$22148 ( \22525 , \22523 , \22524 );
nand \U$22149 ( \22526 , \2346 , \6355 );
nand \U$22150 ( \22527 , \22525 , \22526 );
not \U$22151 ( \22528 , \22527 );
or \U$22152 ( \22529 , \22522 , \22528 );
not \U$22153 ( \22530 , RIc2266b0_33);
not \U$22154 ( \22531 , \4182 );
or \U$22155 ( \22532 , \22530 , \22531 );
nand \U$22156 ( \22533 , \9196 , \5179 );
nand \U$22157 ( \22534 , \22532 , \22533 );
nand \U$22158 ( \22535 , \22534 , \3631 );
nand \U$22159 ( \22536 , \22529 , \22535 );
not \U$22160 ( \22537 , \22536 );
not \U$22161 ( \22538 , \1963 );
not \U$22162 ( \22539 , RIc226e30_17);
not \U$22163 ( \22540 , \4228 );
or \U$22164 ( \22541 , \22539 , \22540 );
not \U$22165 ( \22542 , \9188 );
nand \U$22166 ( \22543 , \22542 , \1935 );
nand \U$22167 ( \22544 , \22541 , \22543 );
not \U$22168 ( \22545 , \22544 );
or \U$22169 ( \22546 , \22538 , \22545 );
not \U$22170 ( \22547 , RIc226e30_17);
not \U$22171 ( \22548 , \2104 );
or \U$22172 ( \22549 , \22547 , \22548 );
nand \U$22173 ( \22550 , \9654 , \1952 );
nand \U$22174 ( \22551 , \22549 , \22550 );
nand \U$22175 ( \22552 , \22551 , \1945 );
nand \U$22176 ( \22553 , \22546 , \22552 );
not \U$22177 ( \22554 , \22553 );
or \U$22178 ( \22555 , \22537 , \22554 );
or \U$22179 ( \22556 , \22536 , \22553 );
not \U$22180 ( \22557 , \2358 );
not \U$22181 ( \22558 , RIc226f20_15);
not \U$22182 ( \22559 , \3116 );
or \U$22183 ( \22560 , \22558 , \22559 );
not \U$22184 ( \22561 , \3116 );
nand \U$22185 ( \22562 , \22561 , \2301 );
nand \U$22186 ( \22563 , \22560 , \22562 );
not \U$22187 ( \22564 , \22563 );
or \U$22188 ( \22565 , \22557 , \22564 );
not \U$22189 ( \22566 , RIc226f20_15);
not \U$22190 ( \22567 , \6439 );
or \U$22191 ( \22568 , \22566 , \22567 );
nand \U$22192 ( \22569 , \2981 , \2301 );
nand \U$22193 ( \22570 , \22568 , \22569 );
nand \U$22194 ( \22571 , \22570 , \2320 );
nand \U$22195 ( \22572 , \22565 , \22571 );
nand \U$22196 ( \22573 , \22556 , \22572 );
nand \U$22197 ( \22574 , \22555 , \22573 );
xor \U$22198 ( \22575 , \22521 , \22574 );
not \U$22199 ( \22576 , \6307 );
not \U$22200 ( \22577 , RIc2263e0_39);
not \U$22201 ( \22578 , \3993 );
or \U$22202 ( \22579 , \22577 , \22578 );
nand \U$22203 ( \22580 , \9540 , \8990 );
nand \U$22204 ( \22581 , \22579 , \22580 );
not \U$22205 ( \22582 , \22581 );
or \U$22206 ( \22583 , \22576 , \22582 );
not \U$22207 ( \22584 , RIc2263e0_39);
not \U$22208 ( \22585 , \1372 );
or \U$22209 ( \22586 , \22584 , \22585 );
nand \U$22210 ( \22587 , \1371 , \5498 );
nand \U$22211 ( \22588 , \22586 , \22587 );
nand \U$22212 ( \22589 , \22588 , \6689 );
nand \U$22213 ( \22590 , \22583 , \22589 );
not \U$22214 ( \22591 , \2086 );
and \U$22215 ( \22592 , RIc226890_29, \2833 );
not \U$22216 ( \22593 , RIc226890_29);
and \U$22217 ( \22594 , \22593 , \2443 );
or \U$22218 ( \22595 , \22592 , \22594 );
not \U$22219 ( \22596 , \22595 );
or \U$22220 ( \22597 , \22591 , \22596 );
not \U$22221 ( \22598 , \22434 );
nand \U$22222 ( \22599 , \22598 , \2784 );
nand \U$22223 ( \22600 , \22597 , \22599 );
xor \U$22224 ( \22601 , \22590 , \22600 );
not \U$22225 ( \22602 , \2138 );
not \U$22226 ( \22603 , RIc226980_27);
not \U$22227 ( \22604 , \3835 );
or \U$22228 ( \22605 , \22603 , \22604 );
nand \U$22229 ( \22606 , \3834 , \2150 );
nand \U$22230 ( \22607 , \22605 , \22606 );
not \U$22231 ( \22608 , \22607 );
or \U$22232 ( \22609 , \22602 , \22608 );
not \U$22233 ( \22610 , RIc226980_27);
not \U$22234 ( \22611 , \4009 );
or \U$22235 ( \22612 , \22610 , \22611 );
nand \U$22236 ( \22613 , \4008 , \2799 );
nand \U$22237 ( \22614 , \22612 , \22613 );
nand \U$22238 ( \22615 , \22614 , \2154 );
nand \U$22239 ( \22616 , \22609 , \22615 );
and \U$22240 ( \22617 , \22601 , \22616 );
and \U$22241 ( \22618 , \22590 , \22600 );
or \U$22242 ( \22619 , \22617 , \22618 );
xor \U$22243 ( \22620 , \22575 , \22619 );
not \U$22244 ( \22621 , \22620 );
not \U$22245 ( \22622 , \22621 );
or \U$22246 ( \22623 , \22485 , \22622 );
not \U$22247 ( \22624 , \22484 );
nand \U$22248 ( \22625 , \22624 , \22620 );
nand \U$22249 ( \22626 , \22623 , \22625 );
not \U$22250 ( \22627 , RIc226110_45);
not \U$22251 ( \22628 , \3071 );
or \U$22252 ( \22629 , \22627 , \22628 );
nand \U$22253 ( \22630 , \1072 , \9100 );
nand \U$22254 ( \22631 , \22629 , \22630 );
and \U$22255 ( \22632 , \22631 , \9934 );
and \U$22256 ( \22633 , \22491 , \9398 );
nor \U$22257 ( \22634 , \22632 , \22633 );
not \U$22258 ( \22635 , \22634 );
not \U$22259 ( \22636 , \22635 );
not \U$22260 ( \22637 , \9705 );
not \U$22261 ( \22638 , RIc2262f0_41);
not \U$22262 ( \22639 , \1558 );
or \U$22263 ( \22640 , \22638 , \22639 );
not \U$22264 ( \22641 , \1558 );
nand \U$22265 ( \22642 , \22641 , \6303 );
nand \U$22266 ( \22643 , \22640 , \22642 );
not \U$22267 ( \22644 , \22643 );
or \U$22268 ( \22645 , \22637 , \22644 );
nand \U$22269 ( \22646 , \22471 , \9690 );
nand \U$22270 ( \22647 , \22645 , \22646 );
not \U$22271 ( \22648 , \22647 );
not \U$22272 ( \22649 , \22648 );
or \U$22273 ( \22650 , \22636 , \22649 );
nand \U$22274 ( \22651 , \22647 , \22634 );
nand \U$22275 ( \22652 , \22650 , \22651 );
not \U$22276 ( \22653 , \2711 );
not \U$22277 ( \22654 , RIc2267a0_31);
not \U$22278 ( \22655 , \10936 );
or \U$22279 ( \22656 , \22654 , \22655 );
nand \U$22280 ( \22657 , \2305 , \3648 );
nand \U$22281 ( \22658 , \22656 , \22657 );
not \U$22282 ( \22659 , \22658 );
or \U$22283 ( \22660 , \22653 , \22659 );
nand \U$22284 ( \22661 , \2697 , \22459 );
nand \U$22285 ( \22662 , \22660 , \22661 );
not \U$22286 ( \22663 , \22662 );
and \U$22287 ( \22664 , \22652 , \22663 );
not \U$22288 ( \22665 , \22652 );
and \U$22289 ( \22666 , \22665 , \22662 );
nor \U$22290 ( \22667 , \22664 , \22666 );
not \U$22291 ( \22668 , \22667 );
not \U$22292 ( \22669 , \22668 );
xor \U$22293 ( \22670 , \22590 , \22600 );
xor \U$22294 ( \22671 , \22670 , \22616 );
not \U$22295 ( \22672 , \22671 );
or \U$22296 ( \22673 , \22669 , \22672 );
or \U$22297 ( \22674 , \22671 , \22668 );
xor \U$22298 ( \22675 , \22553 , \22572 );
xor \U$22299 ( \22676 , \22675 , \22536 );
nand \U$22300 ( \22677 , \22674 , \22676 );
nand \U$22301 ( \22678 , \22673 , \22677 );
and \U$22302 ( \22679 , \22626 , \22678 );
not \U$22303 ( \22680 , \22626 );
not \U$22304 ( \22681 , \22678 );
and \U$22305 ( \22682 , \22680 , \22681 );
nor \U$22306 ( \22683 , \22679 , \22682 );
not \U$22307 ( \22684 , \2173 );
not \U$22308 ( \22685 , \22331 );
or \U$22309 ( \22686 , \22684 , \22685 );
not \U$22310 ( \22687 , RIc226a70_25);
not \U$22311 ( \22688 , \4802 );
or \U$22312 ( \22689 , \22687 , \22688 );
nand \U$22313 ( \22690 , \9942 , \2190 );
nand \U$22314 ( \22691 , \22689 , \22690 );
nand \U$22315 ( \22692 , \22691 , \2195 );
nand \U$22316 ( \22693 , \22686 , \22692 );
not \U$22317 ( \22694 , \5519 );
not \U$22318 ( \22695 , \22313 );
or \U$22319 ( \22696 , \22694 , \22695 );
not \U$22320 ( \22697 , RIc2264d0_37);
not \U$22321 ( \22698 , \1948 );
or \U$22322 ( \22699 , \22697 , \22698 );
nand \U$22323 ( \22700 , \1332 , \12522 );
nand \U$22324 ( \22701 , \22699 , \22700 );
nand \U$22325 ( \22702 , \22701 , \5509 );
nand \U$22326 ( \22703 , \22696 , \22702 );
xor \U$22327 ( \22704 , \22693 , \22703 );
not \U$22328 ( \22705 , \1915 );
not \U$22329 ( \22706 , RIc226b60_23);
not \U$22330 ( \22707 , \12989 );
or \U$22331 ( \22708 , \22706 , \22707 );
nand \U$22332 ( \22709 , \2895 , \1927 );
nand \U$22333 ( \22710 , \22708 , \22709 );
not \U$22334 ( \22711 , \22710 );
or \U$22335 ( \22712 , \22705 , \22711 );
nand \U$22336 ( \22713 , \22397 , \1930 );
nand \U$22337 ( \22714 , \22712 , \22713 );
xor \U$22338 ( \22715 , \22704 , \22714 );
not \U$22339 ( \22716 , \22715 );
not \U$22340 ( \22717 , \9129 );
not \U$22341 ( \22718 , \22352 );
or \U$22342 ( \22719 , \22717 , \22718 );
not \U$22343 ( \22720 , RIc226200_43);
not \U$22344 ( \22721 , \982 );
or \U$22345 ( \22722 , \22720 , \22721 );
nand \U$22346 ( \22723 , \3464 , \9125 );
nand \U$22347 ( \22724 , \22722 , \22723 );
nand \U$22348 ( \22725 , \22724 , \9110 );
nand \U$22349 ( \22726 , \22719 , \22725 );
not \U$22350 ( \22727 , \6307 );
not \U$22351 ( \22728 , \22588 );
or \U$22352 ( \22729 , \22727 , \22728 );
not \U$22353 ( \22730 , RIc2263e0_39);
not \U$22354 ( \22731 , \2380 );
or \U$22355 ( \22732 , \22730 , \22731 );
not \U$22356 ( \22733 , \19678 );
nand \U$22357 ( \22734 , \22733 , \5498 );
nand \U$22358 ( \22735 , \22732 , \22734 );
nand \U$22359 ( \22736 , \22735 , \6688 );
nand \U$22360 ( \22737 , \22729 , \22736 );
xor \U$22361 ( \22738 , \22726 , \22737 );
not \U$22362 ( \22739 , \2154 );
not \U$22363 ( \22740 , \22607 );
or \U$22364 ( \22741 , \22739 , \22740 );
not \U$22365 ( \22742 , RIc226980_27);
not \U$22366 ( \22743 , \11890 );
or \U$22367 ( \22744 , \22742 , \22743 );
nand \U$22368 ( \22745 , \3508 , \2799 );
nand \U$22369 ( \22746 , \22744 , \22745 );
nand \U$22370 ( \22747 , \22746 , \2138 );
nand \U$22371 ( \22748 , \22741 , \22747 );
xnor \U$22372 ( \22749 , \22738 , \22748 );
nand \U$22373 ( \22750 , \22716 , \22749 );
not \U$22374 ( \22751 , \9639 );
not \U$22375 ( \22752 , \14672 );
or \U$22376 ( \22753 , \22751 , \22752 );
not \U$22377 ( \22754 , RIc226020_47);
not \U$22378 ( \22755 , \2700 );
or \U$22379 ( \22756 , \22754 , \22755 );
not \U$22380 ( \22757 , \11112 );
nand \U$22381 ( \22758 , \22757 , \9624 );
nand \U$22382 ( \22759 , \22756 , \22758 );
nand \U$22383 ( \22760 , \22759 , \12304 );
nand \U$22384 ( \22761 , \22753 , \22760 );
not \U$22385 ( \22762 , \3629 );
not \U$22386 ( \22763 , \14693 );
or \U$22387 ( \22764 , \22762 , \22763 );
not \U$22388 ( \22765 , RIc2266b0_33);
not \U$22389 ( \22766 , \3092 );
or \U$22390 ( \22767 , \22765 , \22766 );
nand \U$22391 ( \22768 , \2297 , \6355 );
nand \U$22392 ( \22769 , \22767 , \22768 );
nand \U$22393 ( \22770 , \22769 , \3631 );
nand \U$22394 ( \22771 , \22764 , \22770 );
xor \U$22395 ( \22772 , \22761 , \22771 );
not \U$22396 ( \22773 , \1945 );
not \U$22397 ( \22774 , \14750 );
or \U$22398 ( \22775 , \22773 , \22774 );
not \U$22399 ( \22776 , RIc226e30_17);
not \U$22400 ( \22777 , \9513 );
or \U$22401 ( \22778 , \22776 , \22777 );
nand \U$22402 ( \22779 , \5160 , \1952 );
nand \U$22403 ( \22780 , \22778 , \22779 );
nand \U$22404 ( \22781 , \22780 , \1963 );
nand \U$22405 ( \22782 , \22775 , \22781 );
and \U$22406 ( \22783 , \22772 , \22782 );
and \U$22407 ( \22784 , \22761 , \22771 );
or \U$22408 ( \22785 , \22783 , \22784 );
and \U$22409 ( \22786 , \22750 , \22785 );
nor \U$22410 ( \22787 , \22716 , \22749 );
nor \U$22411 ( \22788 , \22786 , \22787 );
not \U$22412 ( \22789 , \22788 );
not \U$22413 ( \22790 , \22789 );
not \U$22414 ( \22791 , \9398 );
not \U$22415 ( \22792 , \22631 );
or \U$22416 ( \22793 , \22791 , \22792 );
not \U$22417 ( \22794 , \888 );
not \U$22418 ( \22795 , RIc226110_45);
not \U$22419 ( \22796 , \22795 );
and \U$22420 ( \22797 , \22794 , \22796 );
not \U$22421 ( \22798 , \17294 );
and \U$22422 ( \22799 , \22798 , \9379 );
nor \U$22423 ( \22800 , \22797 , \22799 );
not \U$22424 ( \22801 , \22800 );
nand \U$22425 ( \22802 , \22801 , \9384 );
nand \U$22426 ( \22803 , \22793 , \22802 );
not \U$22427 ( \22804 , \1963 );
not \U$22428 ( \22805 , \22551 );
or \U$22429 ( \22806 , \22804 , \22805 );
nand \U$22430 ( \22807 , \22780 , \1945 );
nand \U$22431 ( \22808 , \22806 , \22807 );
xor \U$22432 ( \22809 , \22803 , \22808 );
not \U$22433 ( \22810 , \2358 );
not \U$22434 ( \22811 , \22570 );
or \U$22435 ( \22812 , \22810 , \22811 );
and \U$22436 ( \22813 , RIc226f20_15, \4049 );
not \U$22437 ( \22814 , RIc226f20_15);
and \U$22438 ( \22815 , \22814 , \3641 );
or \U$22439 ( \22816 , \22813 , \22815 );
nand \U$22440 ( \22817 , \22816 , \2320 );
nand \U$22441 ( \22818 , \22812 , \22817 );
xnor \U$22442 ( \22819 , \22809 , \22818 );
xor \U$22443 ( \22820 , \22480 , \22444 );
xor \U$22444 ( \22821 , \22820 , \22461 );
nand \U$22445 ( \22822 , \22819 , \22821 );
not \U$22446 ( \22823 , \4381 );
and \U$22447 ( \22824 , RIc2265c0_35, \13235 );
not \U$22448 ( \22825 , RIc2265c0_35);
and \U$22449 ( \22826 , \22825 , \17977 );
or \U$22450 ( \22827 , \22824 , \22826 );
not \U$22451 ( \22828 , \22827 );
or \U$22452 ( \22829 , \22823 , \22828 );
nand \U$22453 ( \22830 , \22380 , \4383 );
nand \U$22454 ( \22831 , \22829 , \22830 );
not \U$22455 ( \22832 , \2392 );
not \U$22456 ( \22833 , RIc226c50_21);
not \U$22457 ( \22834 , \11841 );
or \U$22458 ( \22835 , \22833 , \22834 );
nand \U$22459 ( \22836 , \2064 , \2383 );
nand \U$22460 ( \22837 , \22835 , \22836 );
not \U$22461 ( \22838 , \22837 );
or \U$22462 ( \22839 , \22832 , \22838 );
nand \U$22463 ( \22840 , \22416 , \2367 );
nand \U$22464 ( \22841 , \22839 , \22840 );
xor \U$22465 ( \22842 , \22831 , \22841 );
not \U$22466 ( \22843 , \2518 );
not \U$22467 ( \22844 , RIc226d40_19);
not \U$22468 ( \22845 , \9188 );
or \U$22469 ( \22846 , \22844 , \22845 );
nand \U$22470 ( \22847 , \9805 , \1941 );
nand \U$22471 ( \22848 , \22846 , \22847 );
not \U$22472 ( \22849 , \22848 );
or \U$22473 ( \22850 , \22843 , \22849 );
not \U$22474 ( \22851 , RIc226d40_19);
not \U$22475 ( \22852 , \2043 );
or \U$22476 ( \22853 , \22851 , \22852 );
nand \U$22477 ( \22854 , \11515 , \3338 );
nand \U$22478 ( \22855 , \22853 , \22854 );
nand \U$22479 ( \22856 , \22855 , \2534 );
nand \U$22480 ( \22857 , \22850 , \22856 );
xor \U$22481 ( \22858 , \22842 , \22857 );
and \U$22482 ( \22859 , \22822 , \22858 );
nor \U$22483 ( \22860 , \22819 , \22821 );
nor \U$22484 ( \22861 , \22859 , \22860 );
not \U$22485 ( \22862 , \22861 );
not \U$22486 ( \22863 , \22862 );
or \U$22487 ( \22864 , \22790 , \22863 );
not \U$22488 ( \22865 , \22861 );
not \U$22489 ( \22866 , \22788 );
or \U$22490 ( \22867 , \22865 , \22866 );
not \U$22491 ( \22868 , \3629 );
not \U$22492 ( \22869 , \22769 );
or \U$22493 ( \22870 , \22868 , \22869 );
nand \U$22494 ( \22871 , \22527 , \3631 );
nand \U$22495 ( \22872 , \22870 , \22871 );
not \U$22496 ( \22873 , \22872 );
not \U$22497 ( \22874 , \1579 );
not \U$22498 ( \22875 , \11566 );
xor \U$22499 ( \22876 , RIc2275b0_1, \22875 );
not \U$22500 ( \22877 , \22876 );
or \U$22501 ( \22878 , \22874 , \22877 );
xor \U$22502 ( \22879 , RIc2275b0_1, \11994 );
nand \U$22503 ( \22880 , \22879 , \854 );
nand \U$22504 ( \22881 , \22878 , \22880 );
not \U$22505 ( \22882 , RIc2275b0_1);
nor \U$22506 ( \22883 , \22882 , \8910 );
or \U$22507 ( \22884 , \22881 , \22883 );
not \U$22508 ( \22885 , \22884 );
or \U$22509 ( \22886 , \22873 , \22885 );
nand \U$22510 ( \22887 , \22881 , \22883 );
nand \U$22511 ( \22888 , \22886 , \22887 );
not \U$22512 ( \22889 , \1340 );
not \U$22513 ( \22890 , RIc2271f0_9);
not \U$22514 ( \22891 , \5665 );
or \U$22515 ( \22892 , \22890 , \22891 );
buf \U$22516 ( \22893 , \5663 );
nand \U$22517 ( \22894 , \22893 , \1342 );
nand \U$22518 ( \22895 , \22892 , \22894 );
not \U$22519 ( \22896 , \22895 );
or \U$22520 ( \22897 , \22889 , \22896 );
not \U$22521 ( \22898 , \1351 );
not \U$22522 ( \22899 , \6071 );
or \U$22523 ( \22900 , \22898 , \22899 );
not \U$22524 ( \22901 , \9769 );
nand \U$22525 ( \22902 , \22901 , RIc2271f0_9);
nand \U$22526 ( \22903 , \22900 , \22902 );
nand \U$22527 ( \22904 , \22903 , \1363 );
nand \U$22528 ( \22905 , \22897 , \22904 );
not \U$22529 ( \22906 , \22905 );
not \U$22530 ( \22907 , \22906 );
not \U$22531 ( \22908 , \951 );
not \U$22532 ( \22909 , RIc2273d0_5);
not \U$22533 ( \22910 , \16531 );
or \U$22534 ( \22911 , \22909 , \22910 );
nand \U$22535 ( \22912 , \8886 , \946 );
nand \U$22536 ( \22913 , \22911 , \22912 );
not \U$22537 ( \22914 , \22913 );
or \U$22538 ( \22915 , \22908 , \22914 );
not \U$22539 ( \22916 , RIc2273d0_5);
not \U$22540 ( \22917 , \10142 );
or \U$22541 ( \22918 , \22916 , \22917 );
nand \U$22542 ( \22919 , \10310 , \946 );
nand \U$22543 ( \22920 , \22918 , \22919 );
nand \U$22544 ( \22921 , \22920 , \954 );
nand \U$22545 ( \22922 , \22915 , \22921 );
not \U$22546 ( \22923 , \22922 );
not \U$22547 ( \22924 , \1121 );
not \U$22548 ( \22925 , RIc2272e0_7);
not \U$22549 ( \22926 , \10125 );
or \U$22550 ( \22927 , \22925 , \22926 );
not \U$22551 ( \22928 , \6492 );
not \U$22552 ( \22929 , \22928 );
nand \U$22553 ( \22930 , \22929 , \4241 );
nand \U$22554 ( \22931 , \22927 , \22930 );
not \U$22555 ( \22932 , \22931 );
or \U$22556 ( \22933 , \22924 , \22932 );
not \U$22557 ( \22934 , RIc2272e0_7);
not \U$22558 ( \22935 , \18410 );
or \U$22559 ( \22936 , \22934 , \22935 );
nand \U$22560 ( \22937 , \9740 , \1139 );
nand \U$22561 ( \22938 , \22936 , \22937 );
nand \U$22562 ( \22939 , \22938 , \1118 );
nand \U$22563 ( \22940 , \22933 , \22939 );
not \U$22564 ( \22941 , \22940 );
not \U$22565 ( \22942 , \22941 );
or \U$22566 ( \22943 , \22923 , \22942 );
or \U$22567 ( \22944 , \22922 , \22941 );
nand \U$22568 ( \22945 , \22943 , \22944 );
not \U$22569 ( \22946 , \22945 );
or \U$22570 ( \22947 , \22907 , \22946 );
or \U$22571 ( \22948 , \22945 , \22906 );
nand \U$22572 ( \22949 , \22947 , \22948 );
xor \U$22573 ( \22950 , \22888 , \22949 );
not \U$22574 ( \22951 , \22803 );
not \U$22575 ( \22952 , \22818 );
or \U$22576 ( \22953 , \22951 , \22952 );
or \U$22577 ( \22954 , \22818 , \22803 );
nand \U$22578 ( \22955 , \22954 , \22808 );
nand \U$22579 ( \22956 , \22953 , \22955 );
xor \U$22580 ( \22957 , \22950 , \22956 );
nand \U$22581 ( \22958 , \22867 , \22957 );
nand \U$22582 ( \22959 , \22864 , \22958 );
not \U$22583 ( \22960 , \22959 );
not \U$22584 ( \22961 , \22960 );
and \U$22585 ( \22962 , RIc2275b0_1, \11994 );
not \U$22586 ( \22963 , \1082 );
not \U$22587 ( \22964 , \22508 );
or \U$22588 ( \22965 , \22963 , \22964 );
not \U$22589 ( \22966 , RIc2274c0_3);
not \U$22590 ( \22967 , \20217 );
or \U$22591 ( \22968 , \22966 , \22967 );
not \U$22592 ( \22969 , \9900 );
nand \U$22593 ( \22970 , \22969 , \2896 );
nand \U$22594 ( \22971 , \22968 , \22970 );
nand \U$22595 ( \22972 , \22971 , \1040 );
nand \U$22596 ( \22973 , \22965 , \22972 );
xor \U$22597 ( \22974 , \22962 , \22973 );
not \U$22598 ( \22975 , \854 );
not \U$22599 ( \22976 , \22876 );
or \U$22600 ( \22977 , \22975 , \22976 );
not \U$22601 ( \22978 , \22515 );
nand \U$22602 ( \22979 , \22978 , \1579 );
nand \U$22603 ( \22980 , \22977 , \22979 );
xnor \U$22604 ( \22981 , \22974 , \22980 );
not \U$22605 ( \22982 , \22981 );
not \U$22606 ( \22983 , \22982 );
not \U$22607 ( \22984 , \9619 );
not \U$22608 ( \22985 , \22984 );
not \U$22609 ( \22986 , \9640 );
or \U$22610 ( \22987 , \22985 , \22986 );
nand \U$22611 ( \22988 , \22987 , RIc226020_47);
not \U$22612 ( \22989 , \1311 );
not \U$22613 ( \22990 , \1302 );
not \U$22614 ( \22991 , \18450 );
not \U$22615 ( \22992 , \22991 );
or \U$22616 ( \22993 , \22990 , \22992 );
not \U$22617 ( \22994 , \4407 );
nand \U$22618 ( \22995 , \22994 , RIc227100_11);
nand \U$22619 ( \22996 , \22993 , \22995 );
not \U$22620 ( \22997 , \22996 );
or \U$22621 ( \22998 , \22989 , \22997 );
not \U$22622 ( \22999 , RIc227100_11);
not \U$22623 ( \23000 , \9850 );
or \U$22624 ( \23001 , \22999 , \23000 );
nand \U$22625 ( \23002 , \13515 , \1302 );
nand \U$22626 ( \23003 , \23001 , \23002 );
nand \U$22627 ( \23004 , \23003 , \1307 );
nand \U$22628 ( \23005 , \22998 , \23004 );
xor \U$22629 ( \23006 , \22988 , \23005 );
not \U$22630 ( \23007 , \1682 );
not \U$22631 ( \23008 , RIc227010_13);
not \U$22632 ( \23009 , \4049 );
or \U$22633 ( \23010 , \23008 , \23009 );
nand \U$22634 ( \23011 , \15768 , \2427 );
nand \U$22635 ( \23012 , \23010 , \23011 );
not \U$22636 ( \23013 , \23012 );
or \U$22637 ( \23014 , \23007 , \23013 );
xnor \U$22638 ( \23015 , RIc227010_13, \4414 );
nand \U$22639 ( \23016 , \23015 , \1680 );
nand \U$22640 ( \23017 , \23014 , \23016 );
xnor \U$22641 ( \23018 , \23006 , \23017 );
not \U$22642 ( \23019 , \23018 );
not \U$22643 ( \23020 , \23019 );
or \U$22644 ( \23021 , \22983 , \23020 );
not \U$22645 ( \23022 , \23018 );
not \U$22646 ( \23023 , \22981 );
or \U$22647 ( \23024 , \23022 , \23023 );
xor \U$22648 ( \23025 , \22831 , \22841 );
and \U$22649 ( \23026 , \23025 , \22857 );
and \U$22650 ( \23027 , \22831 , \22841 );
or \U$22651 ( \23028 , \23026 , \23027 );
nand \U$22652 ( \23029 , \23024 , \23028 );
nand \U$22653 ( \23030 , \23021 , \23029 );
xor \U$22654 ( \23031 , \22888 , \22949 );
and \U$22655 ( \23032 , \23031 , \22956 );
and \U$22656 ( \23033 , \22888 , \22949 );
or \U$22657 ( \23034 , \23032 , \23033 );
xor \U$22658 ( \23035 , \23030 , \23034 );
not \U$22659 ( \23036 , \1082 );
not \U$22660 ( \23037 , \22971 );
or \U$22661 ( \23038 , \23036 , \23037 );
not \U$22662 ( \23039 , RIc2274c0_3);
not \U$22663 ( \23040 , \10858 );
or \U$22664 ( \23041 , \23039 , \23040 );
not \U$22665 ( \23042 , \10295 );
nand \U$22666 ( \23043 , \23042 , \2896 );
nand \U$22667 ( \23044 , \23041 , \23043 );
nand \U$22668 ( \23045 , \23044 , \1040 );
nand \U$22669 ( \23046 , \23038 , \23045 );
not \U$22670 ( \23047 , \10001 );
not \U$22671 ( \23048 , \22759 );
or \U$22672 ( \23049 , \23047 , \23048 );
nand \U$22673 ( \23050 , \9619 , RIc226020_47);
nand \U$22674 ( \23051 , \23049 , \23050 );
xor \U$22675 ( \23052 , \23046 , \23051 );
not \U$22676 ( \23053 , \954 );
not \U$22677 ( \23054 , \22913 );
or \U$22678 ( \23055 , \23053 , \23054 );
not \U$22679 ( \23056 , RIc2273d0_5);
not \U$22680 ( \23057 , \8857 );
or \U$22681 ( \23058 , \23056 , \23057 );
not \U$22682 ( \23059 , \12724 );
nand \U$22683 ( \23060 , \23059 , \946 );
nand \U$22684 ( \23061 , \23058 , \23060 );
nand \U$22685 ( \23062 , \23061 , \951 );
nand \U$22686 ( \23063 , \23055 , \23062 );
and \U$22687 ( \23064 , \23052 , \23063 );
and \U$22688 ( \23065 , \23046 , \23051 );
or \U$22689 ( \23066 , \23064 , \23065 );
xor \U$22690 ( \23067 , \22693 , \22703 );
and \U$22691 ( \23068 , \23067 , \22714 );
and \U$22692 ( \23069 , \22693 , \22703 );
or \U$22693 ( \23070 , \23068 , \23069 );
xor \U$22694 ( \23071 , \23066 , \23070 );
xor \U$22695 ( \23072 , \22726 , \22737 );
and \U$22696 ( \23073 , \23072 , \22748 );
and \U$22697 ( \23074 , \22726 , \22737 );
or \U$22698 ( \23075 , \23073 , \23074 );
and \U$22699 ( \23076 , \23071 , \23075 );
and \U$22700 ( \23077 , \23066 , \23070 );
or \U$22701 ( \23078 , \23076 , \23077 );
xor \U$22702 ( \23079 , \23035 , \23078 );
not \U$22703 ( \23080 , \23079 );
or \U$22704 ( \23081 , \22961 , \23080 );
or \U$22705 ( \23082 , \23079 , \22960 );
nand \U$22706 ( \23083 , \23081 , \23082 );
xnor \U$22707 ( \23084 , \22683 , \23083 );
not \U$22708 ( \23085 , \23084 );
not \U$22709 ( \23086 , \23085 );
not \U$22710 ( \23087 , \1363 );
not \U$22711 ( \23088 , \14923 );
or \U$22712 ( \23089 , \23087 , \23088 );
not \U$22713 ( \23090 , RIc2271f0_9);
not \U$22714 ( \23091 , \12698 );
or \U$22715 ( \23092 , \23090 , \23091 );
nand \U$22716 ( \23093 , \6492 , \1351 );
nand \U$22717 ( \23094 , \23092 , \23093 );
nand \U$22718 ( \23095 , \23094 , \1339 );
nand \U$22719 ( \23096 , \23089 , \23095 );
not \U$22720 ( \23097 , \1311 );
not \U$22721 ( \23098 , RIc227100_11);
not \U$22722 ( \23099 , \15603 );
or \U$22723 ( \23100 , \23098 , \23099 );
nand \U$22724 ( \23101 , \12791 , \3351 );
nand \U$22725 ( \23102 , \23100 , \23101 );
not \U$22726 ( \23103 , \23102 );
or \U$22727 ( \23104 , \23097 , \23103 );
nand \U$22728 ( \23105 , \15000 , \1307 );
nand \U$22729 ( \23106 , \23104 , \23105 );
not \U$22730 ( \23107 , \23106 );
xor \U$22731 ( \23108 , \23096 , \23107 );
not \U$22732 ( \23109 , \1682 );
and \U$22733 ( \23110 , RIc227010_13, \18450 );
not \U$22734 ( \23111 , RIc227010_13);
and \U$22735 ( \23112 , \23111 , \4407 );
or \U$22736 ( \23113 , \23110 , \23112 );
not \U$22737 ( \23114 , \23113 );
or \U$22738 ( \23115 , \23109 , \23114 );
nand \U$22739 ( \23116 , \15009 , \3250 );
nand \U$22740 ( \23117 , \23115 , \23116 );
xor \U$22741 ( \23118 , \23108 , \23117 );
not \U$22742 ( \23119 , \23118 );
or \U$22743 ( \23120 , \14676 , \14686 );
and \U$22744 ( \23121 , \23120 , \14697 );
and \U$22745 ( \23122 , \14676 , \14686 );
nor \U$22746 ( \23123 , \23121 , \23122 );
not \U$22747 ( \23124 , \23123 );
or \U$22748 ( \23125 , \23119 , \23124 );
xor \U$22749 ( \23126 , \14609 , \14618 );
and \U$22750 ( \23127 , \23126 , \14629 );
and \U$22751 ( \23128 , \14609 , \14618 );
or \U$22752 ( \23129 , \23127 , \23128 );
nand \U$22753 ( \23130 , \23125 , \23129 );
not \U$22754 ( \23131 , \23118 );
not \U$22755 ( \23132 , \23123 );
nand \U$22756 ( \23133 , \23131 , \23132 );
nand \U$22757 ( \23134 , \23130 , \23133 );
not \U$22758 ( \23135 , \23134 );
not \U$22759 ( \23136 , \23135 );
not \U$22760 ( \23137 , \1118 );
not \U$22761 ( \23138 , \14907 );
or \U$22762 ( \23139 , \23137 , \23138 );
not \U$22763 ( \23140 , RIc2272e0_7);
not \U$22764 ( \23141 , \10609 );
or \U$22765 ( \23142 , \23140 , \23141 );
nand \U$22766 ( \23143 , \10141 , \1139 );
nand \U$22767 ( \23144 , \23142 , \23143 );
nand \U$22768 ( \23145 , \23144 , \1120 );
nand \U$22769 ( \23146 , \23139 , \23145 );
not \U$22770 ( \23147 , \954 );
not \U$22771 ( \23148 , \23061 );
or \U$22772 ( \23149 , \23147 , \23148 );
not \U$22773 ( \23150 , \14911 );
nand \U$22774 ( \23151 , \23150 , \951 );
nand \U$22775 ( \23152 , \23149 , \23151 );
xor \U$22776 ( \23153 , \23146 , \23152 );
not \U$22777 ( \23154 , \1040 );
not \U$22778 ( \23155 , \14986 );
or \U$22779 ( \23156 , \23154 , \23155 );
nand \U$22780 ( \23157 , \23044 , \1082 );
nand \U$22781 ( \23158 , \23156 , \23157 );
and \U$22782 ( \23159 , \23153 , \23158 );
and \U$22783 ( \23160 , \23146 , \23152 );
or \U$22784 ( \23161 , \23159 , \23160 );
not \U$22785 ( \23162 , \14609 );
not \U$22786 ( \23163 , \2173 );
not \U$22787 ( \23164 , \22691 );
or \U$22788 ( \23165 , \23163 , \23164 );
nand \U$22789 ( \23166 , \14935 , \2860 );
nand \U$22790 ( \23167 , \23165 , \23166 );
xor \U$22791 ( \23168 , \23162 , \23167 );
not \U$22792 ( \23169 , \6307 );
not \U$22793 ( \23170 , \22735 );
or \U$22794 ( \23171 , \23169 , \23170 );
nand \U$22795 ( \23172 , \14945 , \6689 );
nand \U$22796 ( \23173 , \23171 , \23172 );
and \U$22797 ( \23174 , \23168 , \23173 );
and \U$22798 ( \23175 , \23162 , \23167 );
or \U$22799 ( \23176 , \23174 , \23175 );
xor \U$22800 ( \23177 , \23161 , \23176 );
not \U$22801 ( \23178 , \9110 );
not \U$22802 ( \23179 , \14684 );
or \U$22803 ( \23180 , \23178 , \23179 );
nand \U$22804 ( \23181 , \22724 , \9129 );
nand \U$22805 ( \23182 , \23180 , \23181 );
not \U$22806 ( \23183 , \9816 );
not \U$22807 ( \23184 , \22478 );
or \U$22808 ( \23185 , \23183 , \23184 );
nand \U$22809 ( \23186 , \14627 , \9690 );
nand \U$22810 ( \23187 , \23185 , \23186 );
xor \U$22811 ( \23188 , \23182 , \23187 );
not \U$22812 ( \23189 , \3653 );
not \U$22813 ( \23190 , \22452 );
or \U$22814 ( \23191 , \23189 , \23190 );
nand \U$22815 ( \23192 , \14616 , \2697 );
nand \U$22816 ( \23193 , \23191 , \23192 );
and \U$22817 ( \23194 , \23188 , \23193 );
and \U$22818 ( \23195 , \23182 , \23187 );
or \U$22819 ( \23196 , \23194 , \23195 );
xor \U$22820 ( \23197 , \23177 , \23196 );
not \U$22821 ( \23198 , \23197 );
not \U$22822 ( \23199 , \23198 );
or \U$22823 ( \23200 , \23136 , \23199 );
xor \U$22824 ( \23201 , \23162 , \23167 );
xor \U$22825 ( \23202 , \23201 , \23173 );
xor \U$22826 ( \23203 , \22761 , \22771 );
xor \U$22827 ( \23204 , \23203 , \22782 );
xor \U$22828 ( \23205 , \23202 , \23204 );
not \U$22829 ( \23206 , \2086 );
not \U$22830 ( \23207 , \22442 );
or \U$22831 ( \23208 , \23206 , \23207 );
nand \U$22832 ( \23209 , \14640 , \2078 );
nand \U$22833 ( \23210 , \23208 , \23209 );
not \U$22834 ( \23211 , \22800 );
not \U$22835 ( \23212 , \9398 );
not \U$22836 ( \23213 , \23212 );
and \U$22837 ( \23214 , \23211 , \23213 );
and \U$22838 ( \23215 , \14662 , \9934 );
nor \U$22839 ( \23216 , \23214 , \23215 );
not \U$22840 ( \23217 , \23216 );
xor \U$22841 ( \23218 , \23210 , \23217 );
not \U$22842 ( \23219 , \2154 );
not \U$22843 ( \23220 , \22746 );
or \U$22844 ( \23221 , \23219 , \23220 );
nand \U$22845 ( \23222 , \2138 , \14649 );
nand \U$22846 ( \23223 , \23221 , \23222 );
xor \U$22847 ( \23224 , \23218 , \23223 );
and \U$22848 ( \23225 , \23205 , \23224 );
and \U$22849 ( \23226 , \23202 , \23204 );
or \U$22850 ( \23227 , \23225 , \23226 );
nand \U$22851 ( \23228 , \23200 , \23227 );
not \U$22852 ( \23229 , \23135 );
nand \U$22853 ( \23230 , \23229 , \23197 );
nand \U$22854 ( \23231 , \23228 , \23230 );
not \U$22855 ( \23232 , \1363 );
not \U$22856 ( \23233 , \23094 );
or \U$22857 ( \23234 , \23232 , \23233 );
nand \U$22858 ( \23235 , \22903 , \1339 );
nand \U$22859 ( \23236 , \23234 , \23235 );
not \U$22860 ( \23237 , \1120 );
not \U$22861 ( \23238 , \22938 );
or \U$22862 ( \23239 , \23237 , \23238 );
nand \U$22863 ( \23240 , \23144 , \1118 );
nand \U$22864 ( \23241 , \23239 , \23240 );
not \U$22865 ( \23242 , \23241 );
xor \U$22866 ( \23243 , \23236 , \23242 );
not \U$22867 ( \23244 , \1311 );
not \U$22868 ( \23245 , \23003 );
or \U$22869 ( \23246 , \23244 , \23245 );
nand \U$22870 ( \23247 , \23102 , \1307 );
nand \U$22871 ( \23248 , \23246 , \23247 );
xor \U$22872 ( \23249 , \23243 , \23248 );
not \U$22873 ( \23250 , \23249 );
xor \U$22874 ( \23251 , \22883 , \22881 );
xnor \U$22875 ( \23252 , \23251 , \22872 );
not \U$22876 ( \23253 , \23252 );
or \U$22877 ( \23254 , \23250 , \23253 );
not \U$22878 ( \23255 , \23210 );
not \U$22879 ( \23256 , \23217 );
or \U$22880 ( \23257 , \23255 , \23256 );
not \U$22881 ( \23258 , \23210 );
not \U$22882 ( \23259 , \23258 );
not \U$22883 ( \23260 , \23216 );
or \U$22884 ( \23261 , \23259 , \23260 );
nand \U$22885 ( \23262 , \23261 , \23223 );
nand \U$22886 ( \23263 , \23257 , \23262 );
nand \U$22887 ( \23264 , \23254 , \23263 );
not \U$22888 ( \23265 , \23249 );
not \U$22889 ( \23266 , \23252 );
nand \U$22890 ( \23267 , \23265 , \23266 );
nand \U$22891 ( \23268 , \23264 , \23267 );
not \U$22892 ( \23269 , \2367 );
not \U$22893 ( \23270 , \22837 );
or \U$22894 ( \23271 , \23269 , \23270 );
nand \U$22895 ( \23272 , \14730 , \2392 );
nand \U$22896 ( \23273 , \23271 , \23272 );
not \U$22897 ( \23274 , \5509 );
not \U$22898 ( \23275 , \14958 );
or \U$22899 ( \23276 , \23274 , \23275 );
nand \U$22900 ( \23277 , \22701 , \5519 );
nand \U$22901 ( \23278 , \23276 , \23277 );
xor \U$22902 ( \23279 , \23273 , \23278 );
not \U$22903 ( \23280 , \1930 );
not \U$22904 ( \23281 , \22710 );
or \U$22905 ( \23282 , \23280 , \23281 );
nand \U$22906 ( \23283 , \14719 , \1915 );
nand \U$22907 ( \23284 , \23282 , \23283 );
and \U$22908 ( \23285 , \23279 , \23284 );
and \U$22909 ( \23286 , \23273 , \23278 );
or \U$22910 ( \23287 , \23285 , \23286 );
xor \U$22911 ( \23288 , \23046 , \23051 );
xor \U$22912 ( \23289 , \23288 , \23063 );
nor \U$22913 ( \23290 , \23287 , \23289 );
not \U$22914 ( \23291 , \1579 );
not \U$22915 ( \23292 , \22879 );
or \U$22916 ( \23293 , \23291 , \23292 );
nand \U$22917 ( \23294 , \14970 , \854 );
nand \U$22918 ( \23295 , \23293 , \23294 );
not \U$22919 ( \23296 , \5741 );
not \U$22920 ( \23297 , \14742 );
or \U$22921 ( \23298 , \23296 , \23297 );
nand \U$22922 ( \23299 , \22827 , \5135 );
nand \U$22923 ( \23300 , \23298 , \23299 );
xor \U$22924 ( \23301 , \23295 , \23300 );
not \U$22925 ( \23302 , \2534 );
not \U$22926 ( \23303 , \22848 );
or \U$22927 ( \23304 , \23302 , \23303 );
nand \U$22928 ( \23305 , \14761 , \2518 );
nand \U$22929 ( \23306 , \23304 , \23305 );
and \U$22930 ( \23307 , \23301 , \23306 );
and \U$22931 ( \23308 , \23295 , \23300 );
or \U$22932 ( \23309 , \23307 , \23308 );
not \U$22933 ( \23310 , \23309 );
or \U$22934 ( \23311 , \23290 , \23310 );
nand \U$22935 ( \23312 , \23287 , \23289 );
nand \U$22936 ( \23313 , \23311 , \23312 );
xor \U$22937 ( \23314 , \23268 , \23313 );
xor \U$22938 ( \23315 , \23066 , \23070 );
xor \U$22939 ( \23316 , \23315 , \23075 );
xor \U$22940 ( \23317 , \23314 , \23316 );
xor \U$22941 ( \23318 , \23231 , \23317 );
xor \U$22942 ( \23319 , \22957 , \22862 );
xor \U$22943 ( \23320 , \23319 , \22789 );
and \U$22944 ( \23321 , \23318 , \23320 );
and \U$22945 ( \23322 , \23231 , \23317 );
or \U$22946 ( \23323 , \23321 , \23322 );
not \U$22947 ( \23324 , \1682 );
not \U$22948 ( \23325 , \23015 );
or \U$22949 ( \23326 , \23324 , \23325 );
nand \U$22950 ( \23327 , \23113 , \1680 );
nand \U$22951 ( \23328 , \23326 , \23327 );
not \U$22952 ( \23329 , \23328 );
not \U$22953 ( \23330 , \2534 );
not \U$22954 ( \23331 , \3010 );
not \U$22955 ( \23332 , \23331 );
not \U$22956 ( \23333 , \2523 );
or \U$22957 ( \23334 , \23332 , \23333 );
not \U$22958 ( \23335 , \4240 );
nand \U$22959 ( \23336 , \23335 , RIc226d40_19);
nand \U$22960 ( \23337 , \23334 , \23336 );
not \U$22961 ( \23338 , \23337 );
or \U$22962 ( \23339 , \23330 , \23338 );
nand \U$22963 ( \23340 , \22855 , \2518 );
nand \U$22964 ( \23341 , \23339 , \23340 );
not \U$22965 ( \23342 , \23341 );
not \U$22966 ( \23343 , \23342 );
not \U$22967 ( \23344 , \23343 );
or \U$22968 ( \23345 , \23329 , \23344 );
not \U$22969 ( \23346 , \23328 );
nand \U$22970 ( \23347 , \23342 , \23346 );
not \U$22971 ( \23348 , \23236 );
not \U$22972 ( \23349 , \23348 );
not \U$22973 ( \23350 , \23242 );
or \U$22974 ( \23351 , \23349 , \23350 );
nand \U$22975 ( \23352 , \23351 , \23248 );
nand \U$22976 ( \23353 , \23241 , \23236 );
nand \U$22977 ( \23354 , \23352 , \23353 );
nand \U$22978 ( \23355 , \23347 , \23354 );
nand \U$22979 ( \23356 , \23345 , \23355 );
not \U$22980 ( \23357 , \22534 );
not \U$22981 ( \23358 , \3629 );
or \U$22982 ( \23359 , \23357 , \23358 );
not \U$22983 ( \23360 , RIc2266b0_33);
not \U$22984 ( \23361 , \3044 );
or \U$22985 ( \23362 , \23360 , \23361 );
nand \U$22986 ( \23363 , \9116 , \12551 );
nand \U$22987 ( \23364 , \23362 , \23363 );
nand \U$22988 ( \23365 , \23364 , \3631 );
nand \U$22989 ( \23366 , \23359 , \23365 );
not \U$22990 ( \23367 , \5135 );
not \U$22991 ( \23368 , RIc2265c0_35);
not \U$22992 ( \23369 , \1531 );
or \U$22993 ( \23370 , \23368 , \23369 );
nand \U$22994 ( \23371 , \3581 , \3620 );
nand \U$22995 ( \23372 , \23370 , \23371 );
not \U$22996 ( \23373 , \23372 );
or \U$22997 ( \23374 , \23367 , \23373 );
nand \U$22998 ( \23375 , \22374 , \5741 );
nand \U$22999 ( \23376 , \23374 , \23375 );
xor \U$23000 ( \23377 , \23366 , \23376 );
not \U$23001 ( \23378 , \2392 );
not \U$23002 ( \23379 , \22410 );
or \U$23003 ( \23380 , \23378 , \23379 );
not \U$23004 ( \23381 , RIc226c50_21);
not \U$23005 ( \23382 , \2476 );
or \U$23006 ( \23383 , \23381 , \23382 );
nand \U$23007 ( \23384 , \20114 , \3204 );
nand \U$23008 ( \23385 , \23383 , \23384 );
nand \U$23009 ( \23386 , \23385 , \2367 );
nand \U$23010 ( \23387 , \23380 , \23386 );
xor \U$23011 ( \23388 , \23377 , \23387 );
not \U$23012 ( \23389 , \23388 );
and \U$23013 ( \23390 , \23356 , \23389 );
not \U$23014 ( \23391 , \23356 );
and \U$23015 ( \23392 , \23391 , \23388 );
nor \U$23016 ( \23393 , \23390 , \23392 );
not \U$23017 ( \23394 , \23393 );
nor \U$23018 ( \23395 , \22922 , \22905 );
or \U$23019 ( \23396 , \23395 , \22941 );
nand \U$23020 ( \23397 , \22922 , \22905 );
nand \U$23021 ( \23398 , \23396 , \23397 );
or \U$23022 ( \23399 , \22973 , \22962 );
nand \U$23023 ( \23400 , \23399 , \22980 );
nand \U$23024 ( \23401 , \22973 , \22962 );
nand \U$23025 ( \23402 , \23400 , \23401 );
xor \U$23026 ( \23403 , \23398 , \23402 );
not \U$23027 ( \23404 , \22988 );
not \U$23028 ( \23405 , \23017 );
or \U$23029 ( \23406 , \23404 , \23405 );
or \U$23030 ( \23407 , \23017 , \22988 );
nand \U$23031 ( \23408 , \23407 , \23005 );
nand \U$23032 ( \23409 , \23406 , \23408 );
xor \U$23033 ( \23410 , \23403 , \23409 );
not \U$23034 ( \23411 , \23410 );
and \U$23035 ( \23412 , \23394 , \23411 );
and \U$23036 ( \23413 , \23393 , \23410 );
nor \U$23037 ( \23414 , \23412 , \23413 );
not \U$23038 ( \23415 , \9552 );
not \U$23039 ( \23416 , \23415 );
not \U$23040 ( \23417 , \9533 );
or \U$23041 ( \23418 , \23416 , \23417 );
nand \U$23042 ( \23419 , \23418 , RIc225f30_49);
not \U$23043 ( \23420 , \23419 );
not \U$23044 ( \23421 , \9212 );
nand \U$23045 ( \23422 , \23421 , RIc2275b0_1);
nand \U$23046 ( \23423 , \23420 , \23422 );
not \U$23047 ( \23424 , \23423 );
not \U$23048 ( \23425 , \2358 );
not \U$23049 ( \23426 , \22816 );
or \U$23050 ( \23427 , \23425 , \23426 );
nand \U$23051 ( \23428 , \15020 , \2320 );
nand \U$23052 ( \23429 , \23427 , \23428 );
not \U$23053 ( \23430 , \23429 );
or \U$23054 ( \23431 , \23424 , \23430 );
not \U$23055 ( \23432 , \23422 );
nand \U$23056 ( \23433 , \23432 , \23419 );
nand \U$23057 ( \23434 , \23431 , \23433 );
xor \U$23058 ( \23435 , \23346 , \23434 );
nor \U$23059 ( \23436 , \23117 , \23096 );
or \U$23060 ( \23437 , \23436 , \23107 );
nand \U$23061 ( \23438 , \23117 , \23096 );
nand \U$23062 ( \23439 , \23437 , \23438 );
and \U$23063 ( \23440 , \23435 , \23439 );
and \U$23064 ( \23441 , \23346 , \23434 );
or \U$23065 ( \23442 , \23440 , \23441 );
not \U$23066 ( \23443 , \23442 );
not \U$23067 ( \23444 , \23443 );
not \U$23068 ( \23445 , \23328 );
not \U$23069 ( \23446 , \23341 );
not \U$23070 ( \23447 , \23446 );
or \U$23071 ( \23448 , \23445 , \23447 );
nand \U$23072 ( \23449 , \23341 , \23346 );
nand \U$23073 ( \23450 , \23448 , \23449 );
not \U$23074 ( \23451 , \23354 );
and \U$23075 ( \23452 , \23450 , \23451 );
not \U$23076 ( \23453 , \23450 );
and \U$23077 ( \23454 , \23453 , \23354 );
nor \U$23078 ( \23455 , \23452 , \23454 );
not \U$23079 ( \23456 , \23455 );
or \U$23080 ( \23457 , \23444 , \23456 );
xor \U$23081 ( \23458 , \23161 , \23176 );
and \U$23082 ( \23459 , \23458 , \23196 );
and \U$23083 ( \23460 , \23161 , \23176 );
or \U$23084 ( \23461 , \23459 , \23460 );
nand \U$23085 ( \23462 , \23457 , \23461 );
not \U$23086 ( \23463 , \23455 );
nand \U$23087 ( \23464 , \23463 , \23442 );
and \U$23088 ( \23465 , \23462 , \23464 );
xor \U$23089 ( \23466 , \23414 , \23465 );
xor \U$23090 ( \23467 , \23268 , \23313 );
and \U$23091 ( \23468 , \23467 , \23316 );
and \U$23092 ( \23469 , \23268 , \23313 );
or \U$23093 ( \23470 , \23468 , \23469 );
xnor \U$23094 ( \23471 , \23466 , \23470 );
xor \U$23095 ( \23472 , \23323 , \23471 );
not \U$23096 ( \23473 , \23472 );
or \U$23097 ( \23474 , \23086 , \23473 );
not \U$23098 ( \23475 , \23472 );
not \U$23099 ( \23476 , \23085 );
nand \U$23100 ( \23477 , \23475 , \23476 );
nand \U$23101 ( \23478 , \23474 , \23477 );
xnor \U$23102 ( \23479 , \23249 , \23263 );
and \U$23103 ( \23480 , \23479 , \23266 );
not \U$23104 ( \23481 , \23479 );
and \U$23105 ( \23482 , \23481 , \23252 );
nor \U$23106 ( \23483 , \23480 , \23482 );
xor \U$23107 ( \23484 , \22726 , \22737 );
xor \U$23108 ( \23485 , \23484 , \22748 );
xor \U$23109 ( \23486 , \22785 , \23485 );
xor \U$23110 ( \23487 , \23486 , \22715 );
xor \U$23111 ( \23488 , \23483 , \23487 );
xor \U$23112 ( \23489 , \22858 , \22821 );
xor \U$23113 ( \23490 , \23489 , \22819 );
and \U$23114 ( \23491 , \23488 , \23490 );
and \U$23115 ( \23492 , \23483 , \23487 );
or \U$23116 ( \23493 , \23491 , \23492 );
and \U$23117 ( \23494 , \23028 , \22981 );
not \U$23118 ( \23495 , \23028 );
and \U$23119 ( \23496 , \23495 , \22982 );
or \U$23120 ( \23497 , \23494 , \23496 );
xor \U$23121 ( \23498 , \23497 , \23019 );
xor \U$23122 ( \23499 , \22482 , \22425 );
xor \U$23123 ( \23500 , \23499 , \22367 );
xor \U$23124 ( \23501 , \23498 , \23500 );
xor \U$23125 ( \23502 , \22667 , \22671 );
xor \U$23126 ( \23503 , \23502 , \22676 );
xnor \U$23127 ( \23504 , \23501 , \23503 );
xor \U$23128 ( \23505 , \23493 , \23504 );
not \U$23129 ( \23506 , \23429 );
not \U$23130 ( \23507 , \23422 );
not \U$23131 ( \23508 , \23419 );
and \U$23132 ( \23509 , \23507 , \23508 );
and \U$23133 ( \23510 , \23422 , \23419 );
nor \U$23134 ( \23511 , \23509 , \23510 );
not \U$23135 ( \23512 , \23511 );
or \U$23136 ( \23513 , \23506 , \23512 );
or \U$23137 ( \23514 , \23429 , \23511 );
nand \U$23138 ( \23515 , \23513 , \23514 );
not \U$23139 ( \23516 , \14916 );
not \U$23140 ( \23517 , \23516 );
not \U$23141 ( \23518 , \14927 );
or \U$23142 ( \23519 , \23517 , \23518 );
or \U$23143 ( \23520 , \23516 , \14927 );
nand \U$23144 ( \23521 , \23520 , \14909 );
nand \U$23145 ( \23522 , \23519 , \23521 );
xor \U$23146 ( \23523 , \23515 , \23522 );
xor \U$23147 ( \23524 , \15002 , \15013 );
and \U$23148 ( \23525 , \23524 , \15024 );
and \U$23149 ( \23526 , \15002 , \15013 );
or \U$23150 ( \23527 , \23525 , \23526 );
and \U$23151 ( \23528 , \23523 , \23527 );
and \U$23152 ( \23529 , \23515 , \23522 );
or \U$23153 ( \23530 , \23528 , \23529 );
xor \U$23154 ( \23531 , \23346 , \23434 );
xor \U$23155 ( \23532 , \23531 , \23439 );
xor \U$23156 ( \23533 , \23530 , \23532 );
xor \U$23157 ( \23534 , \14974 , \14979 );
and \U$23158 ( \23535 , \23534 , \14990 );
and \U$23159 ( \23536 , \14974 , \14979 );
or \U$23160 ( \23537 , \23535 , \23536 );
xor \U$23161 ( \23538 , \23146 , \23152 );
xor \U$23162 ( \23539 , \23538 , \23158 );
xor \U$23163 ( \23540 , \23537 , \23539 );
xor \U$23164 ( \23541 , \14642 , \14651 );
and \U$23165 ( \23542 , \23541 , \14664 );
and \U$23166 ( \23543 , \14642 , \14651 );
or \U$23167 ( \23544 , \23542 , \23543 );
and \U$23168 ( \23545 , \23540 , \23544 );
and \U$23169 ( \23546 , \23537 , \23539 );
or \U$23170 ( \23547 , \23545 , \23546 );
and \U$23171 ( \23548 , \23533 , \23547 );
and \U$23172 ( \23549 , \23530 , \23532 );
or \U$23173 ( \23550 , \23548 , \23549 );
not \U$23174 ( \23551 , \23463 );
not \U$23175 ( \23552 , \23443 );
or \U$23176 ( \23553 , \23551 , \23552 );
nand \U$23177 ( \23554 , \23455 , \23442 );
nand \U$23178 ( \23555 , \23553 , \23554 );
xor \U$23179 ( \23556 , \23555 , \23461 );
xor \U$23180 ( \23557 , \23550 , \23556 );
xor \U$23181 ( \23558 , \14939 , \14949 );
and \U$23182 ( \23559 , \23558 , \14960 );
and \U$23183 ( \23560 , \14939 , \14949 );
or \U$23184 ( \23561 , \23559 , \23560 );
xor \U$23185 ( \23562 , \14711 , \14721 );
and \U$23186 ( \23563 , \23562 , \14732 );
and \U$23187 ( \23564 , \14711 , \14721 );
or \U$23188 ( \23565 , \23563 , \23564 );
xor \U$23189 ( \23566 , \23561 , \23565 );
xor \U$23190 ( \23567 , \14744 , \14754 );
and \U$23191 ( \23568 , \23567 , \14765 );
and \U$23192 ( \23569 , \14744 , \14754 );
or \U$23193 ( \23570 , \23568 , \23569 );
and \U$23194 ( \23571 , \23566 , \23570 );
and \U$23195 ( \23572 , \23561 , \23565 );
or \U$23196 ( \23573 , \23571 , \23572 );
xor \U$23197 ( \23574 , \23295 , \23300 );
xor \U$23198 ( \23575 , \23574 , \23306 );
xor \U$23199 ( \23576 , \23182 , \23187 );
xor \U$23200 ( \23577 , \23576 , \23193 );
xor \U$23201 ( \23578 , \23575 , \23577 );
xor \U$23202 ( \23579 , \23273 , \23278 );
xor \U$23203 ( \23580 , \23579 , \23284 );
and \U$23204 ( \23581 , \23578 , \23580 );
and \U$23205 ( \23582 , \23575 , \23577 );
or \U$23206 ( \23583 , \23581 , \23582 );
xor \U$23207 ( \23584 , \23573 , \23583 );
xor \U$23208 ( \23585 , \23289 , \23287 );
xor \U$23209 ( \23586 , \23585 , \23309 );
and \U$23210 ( \23587 , \23584 , \23586 );
and \U$23211 ( \23588 , \23573 , \23583 );
or \U$23212 ( \23589 , \23587 , \23588 );
xor \U$23213 ( \23590 , \23557 , \23589 );
xor \U$23214 ( \23591 , \23505 , \23590 );
buf \U$23215 ( \23592 , \23591 );
not \U$23216 ( \23593 , \23592 );
xor \U$23217 ( \23594 , \23530 , \23532 );
xor \U$23218 ( \23595 , \23594 , \23547 );
not \U$23219 ( \23596 , \23595 );
xor \U$23220 ( \23597 , \23561 , \23565 );
xor \U$23221 ( \23598 , \23597 , \23570 );
not \U$23222 ( \23599 , \23598 );
xor \U$23223 ( \23600 , \23537 , \23539 );
xor \U$23224 ( \23601 , \23600 , \23544 );
not \U$23225 ( \23602 , \23601 );
or \U$23226 ( \23603 , \23599 , \23602 );
or \U$23227 ( \23604 , \23598 , \23601 );
not \U$23228 ( \23605 , \14849 );
nand \U$23229 ( \23606 , \23605 , \14840 );
not \U$23230 ( \23607 , \23606 );
not \U$23231 ( \23608 , \14832 );
or \U$23232 ( \23609 , \23607 , \23608 );
nand \U$23233 ( \23610 , \14839 , \14849 );
nand \U$23234 ( \23611 , \23609 , \23610 );
nand \U$23235 ( \23612 , \23604 , \23611 );
nand \U$23236 ( \23613 , \23603 , \23612 );
not \U$23237 ( \23614 , \23613 );
or \U$23238 ( \23615 , \23596 , \23614 );
or \U$23239 ( \23616 , \23613 , \23595 );
xor \U$23240 ( \23617 , \23515 , \23522 );
xor \U$23241 ( \23618 , \23617 , \23527 );
not \U$23242 ( \23619 , \23618 );
not \U$23243 ( \23620 , \23619 );
xor \U$23244 ( \23621 , \14991 , \15025 );
and \U$23245 ( \23622 , \23621 , \15035 );
and \U$23246 ( \23623 , \14991 , \15025 );
or \U$23247 ( \23624 , \23622 , \23623 );
not \U$23248 ( \23625 , \23624 );
not \U$23249 ( \23626 , \23625 );
or \U$23250 ( \23627 , \23620 , \23626 );
xor \U$23251 ( \23628 , \15048 , \15052 );
and \U$23252 ( \23629 , \23628 , \15060 );
and \U$23253 ( \23630 , \15048 , \15052 );
or \U$23254 ( \23631 , \23629 , \23630 );
nand \U$23255 ( \23632 , \23627 , \23631 );
nand \U$23256 ( \23633 , \23624 , \23618 );
nand \U$23257 ( \23634 , \23632 , \23633 );
nand \U$23258 ( \23635 , \23616 , \23634 );
nand \U$23259 ( \23636 , \23615 , \23635 );
xor \U$23260 ( \23637 , \23573 , \23583 );
xor \U$23261 ( \23638 , \23637 , \23586 );
not \U$23262 ( \23639 , \23638 );
buf \U$23263 ( \23640 , \14707 );
or \U$23264 ( \23641 , \14766 , \23640 );
nand \U$23265 ( \23642 , \23641 , \14733 );
nand \U$23266 ( \23643 , \14766 , \23640 );
nand \U$23267 ( \23644 , \23642 , \23643 );
xor \U$23268 ( \23645 , \23575 , \23577 );
xor \U$23269 ( \23646 , \23645 , \23580 );
xor \U$23270 ( \23647 , \23644 , \23646 );
xor \U$23271 ( \23648 , \23202 , \23204 );
xor \U$23272 ( \23649 , \23648 , \23224 );
and \U$23273 ( \23650 , \23647 , \23649 );
and \U$23274 ( \23651 , \23644 , \23646 );
or \U$23275 ( \23652 , \23650 , \23651 );
not \U$23276 ( \23653 , \23652 );
or \U$23277 ( \23654 , \23639 , \23653 );
or \U$23278 ( \23655 , \23638 , \23652 );
not \U$23279 ( \23656 , \14928 );
not \U$23280 ( \23657 , \14899 );
not \U$23281 ( \23658 , \23657 );
or \U$23282 ( \23659 , \23656 , \23658 );
nand \U$23283 ( \23660 , \23659 , \14961 );
or \U$23284 ( \23661 , \23657 , \14928 );
nand \U$23285 ( \23662 , \23660 , \23661 );
not \U$23286 ( \23663 , \23662 );
xor \U$23287 ( \23664 , \23118 , \23129 );
and \U$23288 ( \23665 , \23664 , \23132 );
not \U$23289 ( \23666 , \23664 );
and \U$23290 ( \23667 , \23666 , \23123 );
nor \U$23291 ( \23668 , \23665 , \23667 );
not \U$23292 ( \23669 , \23668 );
not \U$23293 ( \23670 , \23669 );
or \U$23294 ( \23671 , \23663 , \23670 );
or \U$23295 ( \23672 , \23669 , \23662 );
xor \U$23296 ( \23673 , \14630 , \14665 );
and \U$23297 ( \23674 , \23673 , \14698 );
and \U$23298 ( \23675 , \14630 , \14665 );
or \U$23299 ( \23676 , \23674 , \23675 );
nand \U$23300 ( \23677 , \23672 , \23676 );
nand \U$23301 ( \23678 , \23671 , \23677 );
nand \U$23302 ( \23679 , \23655 , \23678 );
nand \U$23303 ( \23680 , \23654 , \23679 );
xor \U$23304 ( \23681 , \23636 , \23680 );
xor \U$23305 ( \23682 , \23231 , \23317 );
xor \U$23306 ( \23683 , \23682 , \23320 );
xor \U$23307 ( \23684 , \23681 , \23683 );
not \U$23308 ( \23685 , \23684 );
or \U$23309 ( \23686 , \23593 , \23685 );
or \U$23310 ( \23687 , \23592 , \23684 );
not \U$23311 ( \23688 , \23134 );
not \U$23312 ( \23689 , \23198 );
or \U$23313 ( \23690 , \23688 , \23689 );
nand \U$23314 ( \23691 , \23197 , \23135 );
nand \U$23315 ( \23692 , \23690 , \23691 );
not \U$23316 ( \23693 , \23227 );
xor \U$23317 ( \23694 , \23692 , \23693 );
not \U$23318 ( \23695 , \23694 );
not \U$23319 ( \23696 , \23695 );
xor \U$23320 ( \23697 , \23483 , \23487 );
xor \U$23321 ( \23698 , \23697 , \23490 );
not \U$23322 ( \23699 , \23698 );
not \U$23323 ( \23700 , \23699 );
not \U$23324 ( \23701 , \23700 );
or \U$23325 ( \23702 , \23696 , \23701 );
not \U$23326 ( \23703 , \23694 );
not \U$23327 ( \23704 , \23699 );
or \U$23328 ( \23705 , \23703 , \23704 );
and \U$23329 ( \23706 , \23631 , \23618 );
not \U$23330 ( \23707 , \23631 );
and \U$23331 ( \23708 , \23707 , \23619 );
nor \U$23332 ( \23709 , \23706 , \23708 );
and \U$23333 ( \23710 , \23709 , \23625 );
not \U$23334 ( \23711 , \23709 );
and \U$23335 ( \23712 , \23711 , \23624 );
nor \U$23336 ( \23713 , \23710 , \23712 );
not \U$23337 ( \23714 , \14868 );
not \U$23338 ( \23715 , \14859 );
or \U$23339 ( \23716 , \23714 , \23715 );
or \U$23340 ( \23717 , \14868 , \14859 );
nand \U$23341 ( \23718 , \23717 , \14873 );
nand \U$23342 ( \23719 , \23716 , \23718 );
not \U$23343 ( \23720 , \23719 );
nand \U$23344 ( \23721 , \23713 , \23720 );
not \U$23345 ( \23722 , \15061 );
not \U$23346 ( \23723 , \15043 );
or \U$23347 ( \23724 , \23722 , \23723 );
or \U$23348 ( \23725 , \15061 , \15043 );
nand \U$23349 ( \23726 , \23725 , \15036 );
nand \U$23350 ( \23727 , \23724 , \23726 );
and \U$23351 ( \23728 , \23721 , \23727 );
nor \U$23352 ( \23729 , \23713 , \23720 );
nor \U$23353 ( \23730 , \23728 , \23729 );
not \U$23354 ( \23731 , \23730 );
nand \U$23355 ( \23732 , \23705 , \23731 );
nand \U$23356 ( \23733 , \23702 , \23732 );
nand \U$23357 ( \23734 , \23687 , \23733 );
nand \U$23358 ( \23735 , \23686 , \23734 );
xor \U$23359 ( \23736 , \23478 , \23735 );
xor \U$23360 ( \23737 , \23550 , \23556 );
and \U$23361 ( \23738 , \23737 , \23589 );
and \U$23362 ( \23739 , \23550 , \23556 );
or \U$23363 ( \23740 , \23738 , \23739 );
not \U$23364 ( \23741 , \23498 );
nand \U$23365 ( \23742 , \23741 , \23503 );
and \U$23366 ( \23743 , \23742 , \23500 );
not \U$23367 ( \23744 , \23498 );
nor \U$23368 ( \23745 , \23744 , \23503 );
nor \U$23369 ( \23746 , \23743 , \23745 );
not \U$23370 ( \23747 , \23746 );
not \U$23371 ( \23748 , \22399 );
not \U$23372 ( \23749 , \22418 );
not \U$23373 ( \23750 , \23749 );
or \U$23374 ( \23751 , \23748 , \23750 );
not \U$23375 ( \23752 , \22418 );
not \U$23376 ( \23753 , \22400 );
or \U$23377 ( \23754 , \23752 , \23753 );
nand \U$23378 ( \23755 , \23754 , \22382 );
nand \U$23379 ( \23756 , \23751 , \23755 );
not \U$23380 ( \23757 , \23756 );
not \U$23381 ( \23758 , \6718 );
and \U$23382 ( \23759 , \946 , \23758 );
not \U$23383 ( \23760 , \946 );
and \U$23384 ( \23761 , \23760 , \9740 );
or \U$23385 ( \23762 , \23759 , \23761 );
not \U$23386 ( \23763 , \23762 );
not \U$23387 ( \23764 , \955 );
and \U$23388 ( \23765 , \23763 , \23764 );
and \U$23389 ( \23766 , \22920 , \950 );
nor \U$23390 ( \23767 , \23765 , \23766 );
not \U$23391 ( \23768 , \1118 );
not \U$23392 ( \23769 , \22931 );
or \U$23393 ( \23770 , \23768 , \23769 );
not \U$23394 ( \23771 , RIc2272e0_7);
not \U$23395 ( \23772 , \13687 );
not \U$23396 ( \23773 , \23772 );
not \U$23397 ( \23774 , \23773 );
or \U$23398 ( \23775 , \23771 , \23774 );
buf \U$23399 ( \23776 , \14998 );
nand \U$23400 ( \23777 , \23776 , \940 );
nand \U$23401 ( \23778 , \23775 , \23777 );
nand \U$23402 ( \23779 , \23778 , \1121 );
nand \U$23403 ( \23780 , \23770 , \23779 );
xor \U$23404 ( \23781 , \23767 , \23780 );
not \U$23405 ( \23782 , \1363 );
not \U$23406 ( \23783 , \22895 );
or \U$23407 ( \23784 , \23782 , \23783 );
and \U$23408 ( \23785 , \5216 , RIc2271f0_9);
not \U$23409 ( \23786 , \5216 );
and \U$23410 ( \23787 , \23786 , \1351 );
or \U$23411 ( \23788 , \23785 , \23787 );
nand \U$23412 ( \23789 , \23788 , \1340 );
nand \U$23413 ( \23790 , \23784 , \23789 );
xor \U$23414 ( \23791 , \23781 , \23790 );
not \U$23415 ( \23792 , \23791 );
and \U$23416 ( \23793 , \23757 , \23792 );
and \U$23417 ( \23794 , \23756 , \23791 );
nor \U$23418 ( \23795 , \23793 , \23794 );
not \U$23419 ( \23796 , \22361 );
not \U$23420 ( \23797 , \22340 );
or \U$23421 ( \23798 , \23796 , \23797 );
not \U$23422 ( \23799 , \22362 );
not \U$23423 ( \23800 , \22341 );
or \U$23424 ( \23801 , \23799 , \23800 );
nand \U$23425 ( \23802 , \23801 , \22323 );
nand \U$23426 ( \23803 , \23798 , \23802 );
and \U$23427 ( \23804 , \23795 , \23803 );
not \U$23428 ( \23805 , \23795 );
not \U$23429 ( \23806 , \23803 );
and \U$23430 ( \23807 , \23805 , \23806 );
nor \U$23431 ( \23808 , \23804 , \23807 );
not \U$23432 ( \23809 , \23808 );
not \U$23433 ( \23810 , \2784 );
not \U$23434 ( \23811 , \22595 );
or \U$23435 ( \23812 , \23810 , \23811 );
xor \U$23436 ( \23813 , RIc226890_29, \2421 );
nand \U$23437 ( \23814 , \23813 , \9142 );
nand \U$23438 ( \23815 , \23812 , \23814 );
not \U$23439 ( \23816 , \9129 );
not \U$23440 ( \23817 , RIc226200_43);
not \U$23441 ( \23818 , \3071 );
or \U$23442 ( \23819 , \23817 , \23818 );
nand \U$23443 ( \23820 , \1072 , \9117 );
nand \U$23444 ( \23821 , \23819 , \23820 );
not \U$23445 ( \23822 , \23821 );
or \U$23446 ( \23823 , \23816 , \23822 );
nand \U$23447 ( \23824 , \22359 , \9110 );
nand \U$23448 ( \23825 , \23823 , \23824 );
xor \U$23449 ( \23826 , \23815 , \23825 );
not \U$23450 ( \23827 , \1682 );
not \U$23451 ( \23828 , RIc227010_13);
not \U$23452 ( \23829 , \12493 );
or \U$23453 ( \23830 , \23828 , \23829 );
nand \U$23454 ( \23831 , \2980 , \1296 );
nand \U$23455 ( \23832 , \23830 , \23831 );
not \U$23456 ( \23833 , \23832 );
or \U$23457 ( \23834 , \23827 , \23833 );
nand \U$23458 ( \23835 , \23012 , \3250 );
nand \U$23459 ( \23836 , \23834 , \23835 );
and \U$23460 ( \23837 , \23826 , \23836 );
not \U$23461 ( \23838 , \23826 );
not \U$23462 ( \23839 , \23836 );
and \U$23463 ( \23840 , \23838 , \23839 );
nor \U$23464 ( \23841 , \23837 , \23840 );
not \U$23465 ( \23842 , \5365 );
not \U$23466 ( \23843 , RIc226b60_23);
not \U$23467 ( \23844 , \9422 );
or \U$23468 ( \23845 , \23843 , \23844 );
nand \U$23469 ( \23846 , \3291 , \1927 );
nand \U$23470 ( \23847 , \23845 , \23846 );
not \U$23471 ( \23848 , \23847 );
or \U$23472 ( \23849 , \23842 , \23848 );
nand \U$23473 ( \23850 , \22390 , \1915 );
nand \U$23474 ( \23851 , \23849 , \23850 );
not \U$23475 ( \23852 , \9690 );
not \U$23476 ( \23853 , \22643 );
or \U$23477 ( \23854 , \23852 , \23853 );
not \U$23478 ( \23855 , RIc2262f0_41);
not \U$23479 ( \23856 , \4608 );
or \U$23480 ( \23857 , \23855 , \23856 );
not \U$23481 ( \23858 , \10450 );
nand \U$23482 ( \23859 , \23858 , \10679 );
nand \U$23483 ( \23860 , \23857 , \23859 );
nand \U$23484 ( \23861 , \23860 , \9816 );
nand \U$23485 ( \23862 , \23854 , \23861 );
xor \U$23486 ( \23863 , \23851 , \23862 );
not \U$23487 ( \23864 , \2860 );
not \U$23488 ( \23865 , \22338 );
or \U$23489 ( \23866 , \23864 , \23865 );
and \U$23490 ( \23867 , RIc226a70_25, \9408 );
not \U$23491 ( \23868 , RIc226a70_25);
and \U$23492 ( \23869 , \23868 , \12509 );
or \U$23493 ( \23870 , \23867 , \23869 );
nand \U$23494 ( \23871 , \23870 , \2173 );
nand \U$23495 ( \23872 , \23866 , \23871 );
xor \U$23496 ( \23873 , \23863 , \23872 );
xor \U$23497 ( \23874 , \23841 , \23873 );
and \U$23498 ( \23875 , RIc2275b0_1, \22875 );
not \U$23499 ( \23876 , \2697 );
not \U$23500 ( \23877 , \22658 );
or \U$23501 ( \23878 , \23876 , \23877 );
not \U$23502 ( \23879 , RIc2267a0_31);
not \U$23503 ( \23880 , \12382 );
or \U$23504 ( \23881 , \23879 , \23880 );
not \U$23505 ( \23882 , \18961 );
nand \U$23506 ( \23883 , \23882 , \2072 );
nand \U$23507 ( \23884 , \23881 , \23883 );
nand \U$23508 ( \23885 , \23884 , \2710 );
nand \U$23509 ( \23886 , \23878 , \23885 );
xor \U$23510 ( \23887 , \23875 , \23886 );
not \U$23511 ( \23888 , \2358 );
buf \U$23512 ( \23889 , \10532 );
and \U$23513 ( \23890 , \23889 , RIc226f20_15);
not \U$23514 ( \23891 , \23889 );
and \U$23515 ( \23892 , \23891 , \2301 );
or \U$23516 ( \23893 , \23890 , \23892 );
not \U$23517 ( \23894 , \23893 );
or \U$23518 ( \23895 , \23888 , \23894 );
nand \U$23519 ( \23896 , \22563 , \2320 );
nand \U$23520 ( \23897 , \23895 , \23896 );
xor \U$23521 ( \23898 , \23887 , \23897 );
xor \U$23522 ( \23899 , \23874 , \23898 );
not \U$23523 ( \23900 , \23899 );
or \U$23524 ( \23901 , \23809 , \23900 );
or \U$23525 ( \23902 , \23808 , \23899 );
nand \U$23526 ( \23903 , \23901 , \23902 );
nor \U$23527 ( \23904 , \22662 , \22635 );
or \U$23528 ( \23905 , \23904 , \22648 );
nand \U$23529 ( \23906 , \22662 , \22635 );
nand \U$23530 ( \23907 , \23905 , \23906 );
and \U$23531 ( \23908 , \22996 , \9904 );
not \U$23532 ( \23909 , \1291 );
not \U$23533 ( \23910 , \13525 );
not \U$23534 ( \23911 , \23910 );
or \U$23535 ( \23912 , \23909 , \23911 );
not \U$23536 ( \23913 , \4418 );
nand \U$23537 ( \23914 , \23913 , RIc227100_11);
nand \U$23538 ( \23915 , \23912 , \23914 );
and \U$23539 ( \23916 , \23915 , \1311 );
nor \U$23540 ( \23917 , \23908 , \23916 );
not \U$23541 ( \23918 , \1945 );
not \U$23542 ( \23919 , \22544 );
or \U$23543 ( \23920 , \23918 , \23919 );
not \U$23544 ( \23921 , RIc226e30_17);
not \U$23545 ( \23922 , \2043 );
or \U$23546 ( \23923 , \23921 , \23922 );
nand \U$23547 ( \23924 , \20183 , \1935 );
nand \U$23548 ( \23925 , \23923 , \23924 );
nand \U$23549 ( \23926 , \23925 , \1963 );
nand \U$23550 ( \23927 , \23920 , \23926 );
xor \U$23551 ( \23928 , \23917 , \23927 );
not \U$23552 ( \23929 , \2518 );
not \U$23553 ( \23930 , \23337 );
or \U$23554 ( \23931 , \23929 , \23930 );
not \U$23555 ( \23932 , RIc226d40_19);
not \U$23556 ( \23933 , \2671 );
or \U$23557 ( \23934 , \23932 , \23933 );
nand \U$23558 ( \23935 , \17831 , \3338 );
nand \U$23559 ( \23936 , \23934 , \23935 );
nand \U$23560 ( \23937 , \23936 , \2534 );
nand \U$23561 ( \23938 , \23931 , \23937 );
xor \U$23562 ( \23939 , \23928 , \23938 );
xor \U$23563 ( \23940 , \23907 , \23939 );
not \U$23564 ( \23941 , \2138 );
not \U$23565 ( \23942 , \22614 );
or \U$23566 ( \23943 , \23941 , \23942 );
not \U$23567 ( \23944 , RIc226980_27);
not \U$23568 ( \23945 , \18086 );
or \U$23569 ( \23946 , \23944 , \23945 );
not \U$23570 ( \23947 , \19226 );
nand \U$23571 ( \23948 , \23947 , \2133 );
nand \U$23572 ( \23949 , \23946 , \23948 );
nand \U$23573 ( \23950 , \23949 , \2154 );
nand \U$23574 ( \23951 , \23943 , \23950 );
not \U$23575 ( \23952 , \6307 );
not \U$23576 ( \23953 , RIc2263e0_39);
not \U$23577 ( \23954 , \11714 );
or \U$23578 ( \23955 , \23953 , \23954 );
nand \U$23579 ( \23956 , \2119 , \8990 );
nand \U$23580 ( \23957 , \23955 , \23956 );
not \U$23581 ( \23958 , \23957 );
or \U$23582 ( \23959 , \23952 , \23958 );
nand \U$23583 ( \23960 , \22581 , \6689 );
nand \U$23584 ( \23961 , \23959 , \23960 );
not \U$23585 ( \23962 , \23961 );
xor \U$23586 ( \23963 , \23951 , \23962 );
not \U$23587 ( \23964 , \5519 );
not \U$23588 ( \23965 , RIc2264d0_37);
not \U$23589 ( \23966 , \1440 );
or \U$23590 ( \23967 , \23965 , \23966 );
nand \U$23591 ( \23968 , \1371 , \5504 );
nand \U$23592 ( \23969 , \23967 , \23968 );
not \U$23593 ( \23970 , \23969 );
or \U$23594 ( \23971 , \23964 , \23970 );
nand \U$23595 ( \23972 , \22321 , \5509 );
nand \U$23596 ( \23973 , \23971 , \23972 );
xnor \U$23597 ( \23974 , \23963 , \23973 );
xor \U$23598 ( \23975 , \23940 , \23974 );
and \U$23599 ( \23976 , \23903 , \23975 );
not \U$23600 ( \23977 , \23903 );
not \U$23601 ( \23978 , \23975 );
and \U$23602 ( \23979 , \23977 , \23978 );
nor \U$23603 ( \23980 , \23976 , \23979 );
not \U$23604 ( \23981 , \23980 );
or \U$23605 ( \23982 , \23747 , \23981 );
or \U$23606 ( \23983 , \23746 , \23980 );
nand \U$23607 ( \23984 , \23982 , \23983 );
xor \U$23608 ( \23985 , \23740 , \23984 );
xor \U$23609 ( \23986 , \23493 , \23504 );
and \U$23610 ( \23987 , \23986 , \23590 );
and \U$23611 ( \23988 , \23493 , \23504 );
or \U$23612 ( \23989 , \23987 , \23988 );
xor \U$23613 ( \23990 , \23985 , \23989 );
xor \U$23614 ( \23991 , \23636 , \23680 );
and \U$23615 ( \23992 , \23991 , \23683 );
and \U$23616 ( \23993 , \23636 , \23680 );
or \U$23617 ( \23994 , \23992 , \23993 );
xor \U$23618 ( \23995 , \23990 , \23994 );
xnor \U$23619 ( \23996 , \23736 , \23995 );
xor \U$23620 ( \23997 , \23595 , \23634 );
xnor \U$23621 ( \23998 , \23997 , \23613 );
xor \U$23622 ( \23999 , \23678 , \23638 );
xnor \U$23623 ( \24000 , \23999 , \23652 );
xor \U$23624 ( \24001 , \23998 , \24000 );
xor \U$23625 ( \24002 , \14882 , \14891 );
and \U$23626 ( \24003 , \24002 , \14962 );
and \U$23627 ( \24004 , \14882 , \14891 );
or \U$23628 ( \24005 , \24003 , \24004 );
xor \U$23629 ( \24006 , \23611 , \23601 );
xnor \U$23630 ( \24007 , \24006 , \23598 );
xor \U$23631 ( \24008 , \24005 , \24007 );
xor \U$23632 ( \24009 , \23662 , \23676 );
xor \U$23633 ( \24010 , \24009 , \23668 );
and \U$23634 ( \24011 , \24008 , \24010 );
and \U$23635 ( \24012 , \24005 , \24007 );
or \U$23636 ( \24013 , \24011 , \24012 );
and \U$23637 ( \24014 , \24001 , \24013 );
and \U$23638 ( \24015 , \23998 , \24000 );
or \U$23639 ( \24016 , \24014 , \24015 );
xor \U$23640 ( \24017 , \23644 , \23646 );
xor \U$23641 ( \24018 , \24017 , \23649 );
buf \U$23642 ( \24019 , \14699 );
not \U$23643 ( \24020 , \24019 );
buf \U$23644 ( \24021 , \14768 );
not \U$23645 ( \24022 , \24021 );
or \U$23646 ( \24023 , \24020 , \24022 );
or \U$23647 ( \24024 , \24021 , \24019 );
nand \U$23648 ( \24025 , \24024 , \14778 );
nand \U$23649 ( \24026 , \24023 , \24025 );
or \U$23650 ( \24027 , \24018 , \24026 );
not \U$23651 ( \24028 , \14817 );
not \U$23652 ( \24029 , \14810 );
or \U$23653 ( \24030 , \24028 , \24029 );
not \U$23654 ( \24031 , \14816 );
not \U$23655 ( \24032 , \14810 );
not \U$23656 ( \24033 , \24032 );
or \U$23657 ( \24034 , \24031 , \24033 );
nand \U$23658 ( \24035 , \24034 , \14827 );
nand \U$23659 ( \24036 , \24030 , \24035 );
and \U$23660 ( \24037 , \24027 , \24036 );
and \U$23661 ( \24038 , \24026 , \24018 );
nor \U$23662 ( \24039 , \24037 , \24038 );
xor \U$23663 ( \24040 , \23694 , \23698 );
xnor \U$23664 ( \24041 , \24040 , \23730 );
xor \U$23665 ( \24042 , \24039 , \24041 );
and \U$23666 ( \24043 , \23727 , \23719 );
not \U$23667 ( \24044 , \23727 );
and \U$23668 ( \24045 , \24044 , \23720 );
nor \U$23669 ( \24046 , \24043 , \24045 );
xnor \U$23670 ( \24047 , \24046 , \23713 );
not \U$23671 ( \24048 , \24047 );
xor \U$23672 ( \24049 , \24005 , \24007 );
xor \U$23673 ( \24050 , \24049 , \24010 );
nand \U$23674 ( \24051 , \24048 , \24050 );
nand \U$23675 ( \24052 , \14963 , \14878 );
and \U$23676 ( \24053 , \24052 , \15063 );
nor \U$23677 ( \24054 , \14878 , \14963 );
nor \U$23678 ( \24055 , \24053 , \24054 );
not \U$23679 ( \24056 , \24055 );
and \U$23680 ( \24057 , \24051 , \24056 );
not \U$23681 ( \24058 , \24047 );
nor \U$23682 ( \24059 , \24058 , \24050 );
nor \U$23683 ( \24060 , \24057 , \24059 );
and \U$23684 ( \24061 , \24042 , \24060 );
and \U$23685 ( \24062 , \24039 , \24041 );
or \U$23686 ( \24063 , \24061 , \24062 );
xor \U$23687 ( \24064 , \24016 , \24063 );
xor \U$23688 ( \24065 , \23733 , \23591 );
xnor \U$23689 ( \24066 , \24065 , \23684 );
and \U$23690 ( \24067 , \24064 , \24066 );
and \U$23691 ( \24068 , \24016 , \24063 );
or \U$23692 ( \24069 , \24067 , \24068 );
nand \U$23693 ( \24070 , \23996 , \24069 );
xor \U$23694 ( \24071 , \23998 , \24000 );
xor \U$23695 ( \24072 , \24071 , \24013 );
xor \U$23696 ( \24073 , \24039 , \24041 );
xor \U$23697 ( \24074 , \24073 , \24060 );
xor \U$23698 ( \24075 , \24072 , \24074 );
not \U$23699 ( \24076 , \14607 );
not \U$23700 ( \24077 , \24076 );
not \U$23701 ( \24078 , \24077 );
not \U$23702 ( \24079 , \14782 );
or \U$23703 ( \24080 , \24078 , \24079 );
not \U$23704 ( \24081 , \14779 );
not \U$23705 ( \24082 , \24076 );
or \U$23706 ( \24083 , \24081 , \24082 );
nand \U$23707 ( \24084 , \24083 , \14791 );
nand \U$23708 ( \24085 , \24080 , \24084 );
not \U$23709 ( \24086 , \24085 );
xor \U$23710 ( \24087 , \24026 , \24018 );
not \U$23711 ( \24088 , \24036 );
and \U$23712 ( \24089 , \24087 , \24088 );
not \U$23713 ( \24090 , \24087 );
and \U$23714 ( \24091 , \24090 , \24036 );
nor \U$23715 ( \24092 , \24089 , \24091 );
buf \U$23716 ( \24093 , \24092 );
nand \U$23717 ( \24094 , \24086 , \24093 );
xor \U$23718 ( \24095 , \24055 , \24047 );
xor \U$23719 ( \24096 , \24095 , \24050 );
and \U$23720 ( \24097 , \24094 , \24096 );
not \U$23721 ( \24098 , \24085 );
nor \U$23722 ( \24099 , \24098 , \24093 );
nor \U$23723 ( \24100 , \24097 , \24099 );
xor \U$23724 ( \24101 , \24075 , \24100 );
not \U$23725 ( \24102 , \15074 );
not \U$23726 ( \24103 , \14828 );
nand \U$23727 ( \24104 , \15068 , \24103 );
not \U$23728 ( \24105 , \24104 );
or \U$23729 ( \24106 , \24102 , \24105 );
nand \U$23730 ( \24107 , \15069 , \14828 );
nand \U$23731 ( \24108 , \24106 , \24107 );
not \U$23732 ( \24109 , \24108 );
xnor \U$23733 ( \24110 , \24092 , \24085 );
xor \U$23734 ( \24111 , \24110 , \24096 );
not \U$23735 ( \24112 , \24111 );
nand \U$23736 ( \24113 , \24109 , \24112 );
not \U$23737 ( \24114 , \14599 );
nand \U$23738 ( \24115 , \24114 , \14792 );
not \U$23739 ( \24116 , \24115 );
not \U$23740 ( \24117 , \14589 );
or \U$23741 ( \24118 , \24116 , \24117 );
not \U$23742 ( \24119 , \14792 );
nand \U$23743 ( \24120 , \24119 , \14795 );
nand \U$23744 ( \24121 , \24118 , \24120 );
buf \U$23745 ( \24122 , \24121 );
and \U$23746 ( \24123 , \24113 , \24122 );
not \U$23747 ( \24124 , \24108 );
nor \U$23748 ( \24125 , \24124 , \24112 );
nor \U$23749 ( \24126 , \24123 , \24125 );
nand \U$23750 ( \24127 , \24101 , \24126 );
buf \U$23751 ( \24128 , \24127 );
xor \U$23752 ( \24129 , \24016 , \24063 );
xor \U$23753 ( \24130 , \24129 , \24066 );
xor \U$23754 ( \24131 , \24072 , \24074 );
and \U$23755 ( \24132 , \24131 , \24100 );
and \U$23756 ( \24133 , \24072 , \24074 );
or \U$23757 ( \24134 , \24132 , \24133 );
nand \U$23758 ( \24135 , \24130 , \24134 );
not \U$23759 ( \24136 , \14801 );
not \U$23760 ( \24137 , \15075 );
or \U$23761 ( \24138 , \24136 , \24137 );
or \U$23762 ( \24139 , \14801 , \15075 );
nand \U$23763 ( \24140 , \24139 , \15087 );
nand \U$23764 ( \24141 , \24138 , \24140 );
not \U$23765 ( \24142 , \24141 );
not \U$23766 ( \24143 , \15074 );
not \U$23767 ( \24144 , \24104 );
or \U$23768 ( \24145 , \24143 , \24144 );
nand \U$23769 ( \24146 , \24145 , \24107 );
not \U$23770 ( \24147 , \24121 );
xor \U$23771 ( \24148 , \24146 , \24147 );
xnor \U$23772 ( \24149 , \24148 , \24111 );
buf \U$23773 ( \24150 , \24149 );
not \U$23774 ( \24151 , \24150 );
nand \U$23775 ( \24152 , \24142 , \24151 );
and \U$23776 ( \24153 , \24070 , \24128 , \24135 , \24152 );
not \U$23777 ( \24154 , \23746 );
not \U$23778 ( \24155 , \24154 );
not \U$23779 ( \24156 , \23980 );
or \U$23780 ( \24157 , \24155 , \24156 );
not \U$23781 ( \24158 , \23746 );
not \U$23782 ( \24159 , \23980 );
not \U$23783 ( \24160 , \24159 );
or \U$23784 ( \24161 , \24158 , \24160 );
nand \U$23785 ( \24162 , \24161 , \23740 );
nand \U$23786 ( \24163 , \24157 , \24162 );
buf \U$23787 ( \24164 , \24163 );
not \U$23788 ( \24165 , \24164 );
not \U$23789 ( \24166 , \23808 );
not \U$23790 ( \24167 , \24166 );
not \U$23791 ( \24168 , \23899 );
or \U$23792 ( \24169 , \24167 , \24168 );
or \U$23793 ( \24170 , \24166 , \23899 );
nand \U$23794 ( \24171 , \24170 , \23975 );
nand \U$23795 ( \24172 , \24169 , \24171 );
not \U$23796 ( \24173 , \24172 );
not \U$23797 ( \24174 , \24173 );
not \U$23798 ( \24175 , \954 );
not \U$23799 ( \24176 , RIc2273d0_5);
not \U$23800 ( \24177 , \22928 );
or \U$23801 ( \24178 , \24176 , \24177 );
nand \U$23802 ( \24179 , \6494 , \946 );
nand \U$23803 ( \24180 , \24178 , \24179 );
not \U$23804 ( \24181 , \24180 );
or \U$23805 ( \24182 , \24175 , \24181 );
not \U$23806 ( \24183 , \23762 );
nand \U$23807 ( \24184 , \24183 , \950 );
nand \U$23808 ( \24185 , \24182 , \24184 );
not \U$23809 ( \24186 , \1121 );
not \U$23810 ( \24187 , RIc2272e0_7);
not \U$23811 ( \24188 , \5665 );
or \U$23812 ( \24189 , \24187 , \24188 );
nand \U$23813 ( \24190 , \6726 , \1139 );
nand \U$23814 ( \24191 , \24189 , \24190 );
not \U$23815 ( \24192 , \24191 );
or \U$23816 ( \24193 , \24186 , \24192 );
nand \U$23817 ( \24194 , \23778 , \1118 );
nand \U$23818 ( \24195 , \24193 , \24194 );
xor \U$23819 ( \24196 , \24185 , \24195 );
not \U$23820 ( \24197 , \1040 );
not \U$23821 ( \24198 , \22502 );
or \U$23822 ( \24199 , \24197 , \24198 );
not \U$23823 ( \24200 , RIc2274c0_3);
not \U$23824 ( \24201 , \15699 );
or \U$23825 ( \24202 , \24200 , \24201 );
nand \U$23826 ( \24203 , \10141 , \1078 );
nand \U$23827 ( \24204 , \24202 , \24203 );
nand \U$23828 ( \24205 , \24204 , \1082 );
nand \U$23829 ( \24206 , \24199 , \24205 );
xor \U$23830 ( \24207 , \24196 , \24206 );
and \U$23831 ( \24208 , \8811 , RIc2275b0_1);
not \U$23832 ( \24209 , \1579 );
and \U$23833 ( \24210 , RIc2275b0_1, \20674 );
not \U$23834 ( \24211 , RIc2275b0_1);
and \U$23835 ( \24212 , \24211 , \12727 );
or \U$23836 ( \24213 , \24210 , \24212 );
not \U$23837 ( \24214 , \24213 );
or \U$23838 ( \24215 , \24209 , \24214 );
nand \U$23839 ( \24216 , \22517 , \854 );
nand \U$23840 ( \24217 , \24215 , \24216 );
xor \U$23841 ( \24218 , \24208 , \24217 );
not \U$23842 ( \24219 , \2710 );
not \U$23843 ( \24220 , RIc2267a0_31);
not \U$23844 ( \24221 , \9197 );
or \U$23845 ( \24222 , \24220 , \24221 );
not \U$23846 ( \24223 , \13235 );
nand \U$23847 ( \24224 , \24223 , \6902 );
nand \U$23848 ( \24225 , \24222 , \24224 );
not \U$23849 ( \24226 , \24225 );
or \U$23850 ( \24227 , \24219 , \24226 );
nand \U$23851 ( \24228 , \23884 , \2697 );
nand \U$23852 ( \24229 , \24227 , \24228 );
xor \U$23853 ( \24230 , \24218 , \24229 );
xor \U$23854 ( \24231 , \24207 , \24230 );
xor \U$23855 ( \24232 , \23366 , \23376 );
and \U$23856 ( \24233 , \24232 , \23387 );
and \U$23857 ( \24234 , \23366 , \23376 );
or \U$23858 ( \24235 , \24233 , \24234 );
xor \U$23859 ( \24236 , \24231 , \24235 );
not \U$23860 ( \24237 , \24236 );
xor \U$23861 ( \24238 , \23917 , \23927 );
and \U$23862 ( \24239 , \24238 , \23938 );
and \U$23863 ( \24240 , \23917 , \23927 );
or \U$23864 ( \24241 , \24239 , \24240 );
not \U$23865 ( \24242 , \23825 );
not \U$23866 ( \24243 , \23815 );
or \U$23867 ( \24244 , \24242 , \24243 );
or \U$23868 ( \24245 , \23815 , \23825 );
nand \U$23869 ( \24246 , \24245 , \23836 );
nand \U$23870 ( \24247 , \24244 , \24246 );
not \U$23871 ( \24248 , \24247 );
nor \U$23872 ( \24249 , \23973 , \23951 );
or \U$23873 ( \24250 , \24249 , \23962 );
nand \U$23874 ( \24251 , \23973 , \23951 );
nand \U$23875 ( \24252 , \24250 , \24251 );
not \U$23876 ( \24253 , \24252 );
not \U$23877 ( \24254 , \24253 );
or \U$23878 ( \24255 , \24248 , \24254 );
not \U$23879 ( \24256 , \24247 );
nand \U$23880 ( \24257 , \24256 , \24252 );
nand \U$23881 ( \24258 , \24255 , \24257 );
xnor \U$23882 ( \24259 , \24241 , \24258 );
not \U$23883 ( \24260 , \24259 );
or \U$23884 ( \24261 , \24237 , \24260 );
or \U$23885 ( \24262 , \24236 , \24259 );
nand \U$23886 ( \24263 , \24261 , \24262 );
not \U$23887 ( \24264 , \3631 );
not \U$23888 ( \24265 , RIc2266b0_33);
not \U$23889 ( \24266 , \3438 );
or \U$23890 ( \24267 , \24265 , \24266 );
nand \U$23891 ( \24268 , \3439 , \5179 );
nand \U$23892 ( \24269 , \24267 , \24268 );
not \U$23893 ( \24270 , \24269 );
or \U$23894 ( \24271 , \24264 , \24270 );
nand \U$23895 ( \24272 , \23364 , \3629 );
nand \U$23896 ( \24273 , \24271 , \24272 );
not \U$23897 ( \24274 , \2518 );
not \U$23898 ( \24275 , \23936 );
or \U$23899 ( \24276 , \24274 , \24275 );
not \U$23900 ( \24277 , RIc226d40_19);
not \U$23901 ( \24278 , \3022 );
or \U$23902 ( \24279 , \24277 , \24278 );
nand \U$23903 ( \24280 , \2500 , \1941 );
nand \U$23904 ( \24281 , \24279 , \24280 );
nand \U$23905 ( \24282 , \24281 , \2534 );
nand \U$23906 ( \24283 , \24276 , \24282 );
xor \U$23907 ( \24284 , \24273 , \24283 );
not \U$23908 ( \24285 , \1963 );
not \U$23909 ( \24286 , RIc226e30_17);
not \U$23910 ( \24287 , \3010 );
or \U$23911 ( \24288 , \24286 , \24287 );
nand \U$23912 ( \24289 , \23331 , \1935 );
nand \U$23913 ( \24290 , \24288 , \24289 );
not \U$23914 ( \24291 , \24290 );
or \U$23915 ( \24292 , \24285 , \24291 );
nand \U$23916 ( \24293 , \23925 , \1945 );
nand \U$23917 ( \24294 , \24292 , \24293 );
and \U$23918 ( \24295 , \24284 , \24294 );
not \U$23919 ( \24296 , \24284 );
not \U$23920 ( \24297 , \24294 );
and \U$23921 ( \24298 , \24296 , \24297 );
nor \U$23922 ( \24299 , \24295 , \24298 );
not \U$23923 ( \24300 , \1930 );
not \U$23924 ( \24301 , RIc226b60_23);
not \U$23925 ( \24302 , \2014 );
not \U$23926 ( \24303 , \24302 );
or \U$23927 ( \24304 , \24301 , \24303 );
nand \U$23928 ( \24305 , \2014 , \2111 );
nand \U$23929 ( \24306 , \24304 , \24305 );
not \U$23930 ( \24307 , \24306 );
or \U$23931 ( \24308 , \24300 , \24307 );
nand \U$23932 ( \24309 , \23847 , \1915 );
nand \U$23933 ( \24310 , \24308 , \24309 );
not \U$23934 ( \24311 , \2392 );
not \U$23935 ( \24312 , \23385 );
or \U$23936 ( \24313 , \24311 , \24312 );
not \U$23937 ( \24314 , RIc226c50_21);
not \U$23938 ( \24315 , \2556 );
or \U$23939 ( \24316 , \24314 , \24315 );
not \U$23940 ( \24317 , \9361 );
nand \U$23941 ( \24318 , \24317 , \2383 );
nand \U$23942 ( \24319 , \24316 , \24318 );
nand \U$23943 ( \24320 , \24319 , \2367 );
nand \U$23944 ( \24321 , \24313 , \24320 );
xor \U$23945 ( \24322 , \24310 , \24321 );
not \U$23946 ( \24323 , \5135 );
not \U$23947 ( \24324 , RIc2265c0_35);
not \U$23948 ( \24325 , \1393 );
or \U$23949 ( \24326 , \24324 , \24325 );
nand \U$23950 ( \24327 , \5247 , \3620 );
nand \U$23951 ( \24328 , \24326 , \24327 );
not \U$23952 ( \24329 , \24328 );
or \U$23953 ( \24330 , \24323 , \24329 );
nand \U$23954 ( \24331 , \23372 , \4381 );
nand \U$23955 ( \24332 , \24330 , \24331 );
xor \U$23956 ( \24333 , \24322 , \24332 );
not \U$23957 ( \24334 , \24333 );
and \U$23958 ( \24335 , \24299 , \24334 );
not \U$23959 ( \24336 , \24299 );
and \U$23960 ( \24337 , \24336 , \24333 );
nor \U$23961 ( \24338 , \24335 , \24337 );
not \U$23962 ( \24339 , \6689 );
not \U$23963 ( \24340 , \23957 );
or \U$23964 ( \24341 , \24339 , \24340 );
not \U$23965 ( \24342 , RIc2263e0_39);
not \U$23966 ( \24343 , \1558 );
or \U$23967 ( \24344 , \24342 , \24343 );
nand \U$23968 ( \24345 , \22641 , \5498 );
nand \U$23969 ( \24346 , \24344 , \24345 );
nand \U$23970 ( \24347 , \24346 , \6307 );
nand \U$23971 ( \24348 , \24341 , \24347 );
not \U$23972 ( \24349 , \2154 );
not \U$23973 ( \24350 , RIc226980_27);
not \U$23974 ( \24351 , \2833 );
or \U$23975 ( \24352 , \24350 , \24351 );
nand \U$23976 ( \24353 , \5949 , \16510 );
nand \U$23977 ( \24354 , \24352 , \24353 );
not \U$23978 ( \24355 , \24354 );
or \U$23979 ( \24356 , \24349 , \24355 );
nand \U$23980 ( \24357 , \23949 , \2138 );
nand \U$23981 ( \24358 , \24356 , \24357 );
xor \U$23982 ( \24359 , \24348 , \24358 );
not \U$23983 ( \24360 , \2784 );
not \U$23984 ( \24361 , \23813 );
or \U$23985 ( \24362 , \24360 , \24361 );
not \U$23986 ( \24363 , RIc226890_29);
not \U$23987 ( \24364 , \2304 );
or \U$23988 ( \24365 , \24363 , \24364 );
not \U$23989 ( \24366 , \3092 );
nand \U$23990 ( \24367 , \24366 , \9144 );
nand \U$23991 ( \24368 , \24365 , \24367 );
nand \U$23992 ( \24369 , \24368 , \2086 );
nand \U$23993 ( \24370 , \24362 , \24369 );
and \U$23994 ( \24371 , \24359 , \24370 );
not \U$23995 ( \24372 , \24359 );
not \U$23996 ( \24373 , \24370 );
and \U$23997 ( \24374 , \24372 , \24373 );
nor \U$23998 ( \24375 , \24371 , \24374 );
xor \U$23999 ( \24376 , \24338 , \24375 );
and \U$24000 ( \24377 , \24263 , \24376 );
not \U$24001 ( \24378 , \24263 );
not \U$24002 ( \24379 , \24376 );
and \U$24003 ( \24380 , \24378 , \24379 );
nor \U$24004 ( \24381 , \24377 , \24380 );
not \U$24005 ( \24382 , \24381 );
not \U$24006 ( \24383 , \24382 );
or \U$24007 ( \24384 , \24174 , \24383 );
nand \U$24008 ( \24385 , \24381 , \24172 );
nand \U$24009 ( \24386 , \24384 , \24385 );
nand \U$24010 ( \24387 , \23414 , \23465 );
and \U$24011 ( \24388 , \24387 , \23470 );
nor \U$24012 ( \24389 , \23465 , \23414 );
nor \U$24013 ( \24390 , \24388 , \24389 );
and \U$24014 ( \24391 , \24386 , \24390 );
not \U$24015 ( \24392 , \24386 );
not \U$24016 ( \24393 , \24390 );
and \U$24017 ( \24394 , \24392 , \24393 );
nor \U$24018 ( \24395 , \24391 , \24394 );
buf \U$24019 ( \24396 , \24395 );
nand \U$24020 ( \24397 , \24165 , \24396 );
not \U$24021 ( \24398 , \24397 );
not \U$24022 ( \24399 , \23471 );
not \U$24023 ( \24400 , \23084 );
or \U$24024 ( \24401 , \24399 , \24400 );
nand \U$24025 ( \24402 , \24401 , \23323 );
not \U$24026 ( \24403 , \23471 );
nand \U$24027 ( \24404 , \24403 , \23085 );
nand \U$24028 ( \24405 , \24402 , \24404 );
not \U$24029 ( \24406 , \24405 );
or \U$24030 ( \24407 , \24398 , \24406 );
not \U$24031 ( \24408 , \24396 );
nand \U$24032 ( \24409 , \24408 , \24164 );
nand \U$24033 ( \24410 , \24407 , \24409 );
not \U$24034 ( \24411 , \9110 );
not \U$24035 ( \24412 , \23821 );
or \U$24036 ( \24413 , \24411 , \24412 );
not \U$24037 ( \24414 , RIc226200_43);
not \U$24038 ( \24415 , \2701 );
or \U$24039 ( \24416 , \24414 , \24415 );
nand \U$24040 ( \24417 , \931 , \9117 );
nand \U$24041 ( \24418 , \24416 , \24417 );
nand \U$24042 ( \24419 , \24418 , \9205 );
nand \U$24043 ( \24420 , \24413 , \24419 );
not \U$24044 ( \24421 , \1682 );
not \U$24045 ( \24422 , RIc227010_13);
not \U$24046 ( \24423 , \9513 );
or \U$24047 ( \24424 , \24422 , \24423 );
nand \U$24048 ( \24425 , \5160 , \2427 );
nand \U$24049 ( \24426 , \24424 , \24425 );
not \U$24050 ( \24427 , \24426 );
or \U$24051 ( \24428 , \24421 , \24427 );
nand \U$24052 ( \24429 , \23832 , \1680 );
nand \U$24053 ( \24430 , \24428 , \24429 );
xor \U$24054 ( \24431 , \24420 , \24430 );
not \U$24055 ( \24432 , \2320 );
not \U$24056 ( \24433 , \23893 );
or \U$24057 ( \24434 , \24432 , \24433 );
not \U$24058 ( \24435 , RIc226f20_15);
not \U$24059 ( \24436 , \4228 );
or \U$24060 ( \24437 , \24435 , \24436 );
nand \U$24061 ( \24438 , \2636 , \1674 );
nand \U$24062 ( \24439 , \24437 , \24438 );
nand \U$24063 ( \24440 , \2358 , \24439 );
nand \U$24064 ( \24441 , \24434 , \24440 );
xnor \U$24065 ( \24442 , \24431 , \24441 );
not \U$24066 ( \24443 , \5509 );
not \U$24067 ( \24444 , \23969 );
or \U$24068 ( \24445 , \24443 , \24444 );
not \U$24069 ( \24446 , RIc2264d0_37);
not \U$24070 ( \24447 , \17161 );
or \U$24071 ( \24448 , \24446 , \24447 );
not \U$24072 ( \24449 , \9539 );
nand \U$24073 ( \24450 , \24449 , \5514 );
nand \U$24074 ( \24451 , \24448 , \24450 );
nand \U$24075 ( \24452 , \24451 , \5519 );
nand \U$24076 ( \24453 , \24445 , \24452 );
not \U$24077 ( \24454 , \24453 );
not \U$24078 ( \24455 , \24454 );
not \U$24079 ( \24456 , \2860 );
not \U$24080 ( \24457 , \23870 );
or \U$24081 ( \24458 , \24456 , \24457 );
not \U$24082 ( \24459 , RIc226a70_25);
not \U$24083 ( \24460 , \2258 );
or \U$24084 ( \24461 , \24459 , \24460 );
nand \U$24085 ( \24462 , \4008 , \1905 );
nand \U$24086 ( \24463 , \24461 , \24462 );
nand \U$24087 ( \24464 , \24463 , \2173 );
nand \U$24088 ( \24465 , \24458 , \24464 );
not \U$24089 ( \24466 , \9690 );
not \U$24090 ( \24467 , \23860 );
or \U$24091 ( \24468 , \24466 , \24467 );
not \U$24092 ( \24469 , RIc2262f0_41);
not \U$24093 ( \24470 , \4024 );
or \U$24094 ( \24471 , \24469 , \24470 );
nand \U$24095 ( \24472 , \888 , \6303 );
nand \U$24096 ( \24473 , \24471 , \24472 );
nand \U$24097 ( \24474 , \24473 , \9816 );
nand \U$24098 ( \24475 , \24468 , \24474 );
xor \U$24099 ( \24476 , \24465 , \24475 );
not \U$24100 ( \24477 , \24476 );
or \U$24101 ( \24478 , \24455 , \24477 );
or \U$24102 ( \24479 , \24476 , \24454 );
nand \U$24103 ( \24480 , \24478 , \24479 );
and \U$24104 ( \24481 , \24442 , \24480 );
not \U$24105 ( \24482 , \24442 );
not \U$24106 ( \24483 , \24480 );
and \U$24107 ( \24484 , \24482 , \24483 );
or \U$24108 ( \24485 , \24481 , \24484 );
xor \U$24109 ( \24486 , \23398 , \23402 );
and \U$24110 ( \24487 , \24486 , \23409 );
and \U$24111 ( \24488 , \23398 , \23402 );
or \U$24112 ( \24489 , \24487 , \24488 );
xor \U$24113 ( \24490 , \24485 , \24489 );
not \U$24114 ( \24491 , \23388 );
not \U$24115 ( \24492 , \23410 );
or \U$24116 ( \24493 , \24491 , \24492 );
or \U$24117 ( \24494 , \23410 , \23388 );
nand \U$24118 ( \24495 , \24494 , \23356 );
nand \U$24119 ( \24496 , \24493 , \24495 );
xor \U$24120 ( \24497 , \24490 , \24496 );
xor \U$24121 ( \24498 , \23030 , \23034 );
and \U$24122 ( \24499 , \24498 , \23078 );
and \U$24123 ( \24500 , \23030 , \23034 );
or \U$24124 ( \24501 , \24499 , \24500 );
and \U$24125 ( \24502 , \24497 , \24501 );
and \U$24126 ( \24503 , \24490 , \24496 );
or \U$24127 ( \24504 , \24502 , \24503 );
not \U$24128 ( \24505 , \23917 );
xor \U$24129 ( \24506 , \22495 , \22510 );
and \U$24130 ( \24507 , \24506 , \22520 );
and \U$24131 ( \24508 , \22495 , \22510 );
or \U$24132 ( \24509 , \24507 , \24508 );
xor \U$24133 ( \24510 , \24505 , \24509 );
not \U$24134 ( \24511 , \23790 );
not \U$24135 ( \24512 , \23767 );
not \U$24136 ( \24513 , \24512 );
or \U$24137 ( \24514 , \24511 , \24513 );
or \U$24138 ( \24515 , \24512 , \23790 );
nand \U$24139 ( \24516 , \24515 , \23780 );
nand \U$24140 ( \24517 , \24514 , \24516 );
xor \U$24141 ( \24518 , \24510 , \24517 );
not \U$24142 ( \24519 , \23803 );
not \U$24143 ( \24520 , \23756 );
or \U$24144 ( \24521 , \24519 , \24520 );
or \U$24145 ( \24522 , \23803 , \23756 );
not \U$24146 ( \24523 , \23791 );
nand \U$24147 ( \24524 , \24522 , \24523 );
nand \U$24148 ( \24525 , \24521 , \24524 );
xor \U$24149 ( \24526 , \24518 , \24525 );
xor \U$24150 ( \24527 , \22521 , \22574 );
and \U$24151 ( \24528 , \24527 , \22619 );
and \U$24152 ( \24529 , \22521 , \22574 );
or \U$24153 ( \24530 , \24528 , \24529 );
xor \U$24154 ( \24531 , \24526 , \24530 );
not \U$24155 ( \24532 , \22678 );
not \U$24156 ( \24533 , \22620 );
or \U$24157 ( \24534 , \24532 , \24533 );
or \U$24158 ( \24535 , \22620 , \22678 );
nand \U$24159 ( \24536 , \24535 , \22484 );
nand \U$24160 ( \24537 , \24534 , \24536 );
xor \U$24161 ( \24538 , \24531 , \24537 );
not \U$24162 ( \24539 , \23974 );
not \U$24163 ( \24540 , \23907 );
or \U$24164 ( \24541 , \24539 , \24540 );
or \U$24165 ( \24542 , \23974 , \23907 );
nand \U$24166 ( \24543 , \24542 , \23939 );
nand \U$24167 ( \24544 , \24541 , \24543 );
or \U$24168 ( \24545 , \9934 , \11825 );
nand \U$24169 ( \24546 , \24545 , RIc226110_45);
not \U$24170 ( \24547 , \1340 );
not \U$24171 ( \24548 , RIc2271f0_9);
not \U$24172 ( \24549 , \4407 );
not \U$24173 ( \24550 , \24549 );
or \U$24174 ( \24551 , \24548 , \24550 );
nand \U$24175 ( \24552 , \6079 , \1351 );
nand \U$24176 ( \24553 , \24551 , \24552 );
not \U$24177 ( \24554 , \24553 );
or \U$24178 ( \24555 , \24547 , \24554 );
nand \U$24179 ( \24556 , \23788 , \1363 );
nand \U$24180 ( \24557 , \24555 , \24556 );
xor \U$24181 ( \24558 , \24546 , \24557 );
not \U$24182 ( \24559 , \1311 );
not \U$24183 ( \24560 , RIc227100_11);
not \U$24184 ( \24561 , \19926 );
or \U$24185 ( \24562 , \24560 , \24561 );
nand \U$24186 ( \24563 , \15768 , \3351 );
nand \U$24187 ( \24564 , \24562 , \24563 );
not \U$24188 ( \24565 , \24564 );
or \U$24189 ( \24566 , \24559 , \24565 );
nand \U$24190 ( \24567 , \23915 , \1307 );
nand \U$24191 ( \24568 , \24566 , \24567 );
xor \U$24192 ( \24569 , \24558 , \24568 );
xor \U$24193 ( \24570 , \23875 , \23886 );
and \U$24194 ( \24571 , \24570 , \23897 );
and \U$24195 ( \24572 , \23875 , \23886 );
or \U$24196 ( \24573 , \24571 , \24572 );
xor \U$24197 ( \24574 , \24569 , \24573 );
xor \U$24198 ( \24575 , \23851 , \23862 );
and \U$24199 ( \24576 , \24575 , \23872 );
and \U$24200 ( \24577 , \23851 , \23862 );
or \U$24201 ( \24578 , \24576 , \24577 );
xor \U$24202 ( \24579 , \24574 , \24578 );
xor \U$24203 ( \24580 , \24544 , \24579 );
xor \U$24204 ( \24581 , \23841 , \23873 );
and \U$24205 ( \24582 , \24581 , \23898 );
and \U$24206 ( \24583 , \23841 , \23873 );
or \U$24207 ( \24584 , \24582 , \24583 );
xor \U$24208 ( \24585 , \24580 , \24584 );
and \U$24209 ( \24586 , \24538 , \24585 );
and \U$24210 ( \24587 , \24531 , \24537 );
or \U$24211 ( \24588 , \24586 , \24587 );
xor \U$24212 ( \24589 , \24504 , \24588 );
not \U$24213 ( \24590 , \1363 );
not \U$24214 ( \24591 , \24553 );
or \U$24215 ( \24592 , \24590 , \24591 );
not \U$24216 ( \24593 , RIc2271f0_9);
not \U$24217 ( \24594 , \4123 );
or \U$24218 ( \24595 , \24593 , \24594 );
nand \U$24219 ( \24596 , \5569 , \1342 );
nand \U$24220 ( \24597 , \24595 , \24596 );
nand \U$24221 ( \24598 , \24597 , \1340 );
nand \U$24222 ( \24599 , \24592 , \24598 );
not \U$24223 ( \24600 , \24599 );
not \U$24224 ( \24601 , \2358 );
not \U$24225 ( \24602 , RIc226f20_15);
not \U$24226 ( \24603 , \2043 );
or \U$24227 ( \24604 , \24602 , \24603 );
nand \U$24228 ( \24605 , \5528 , \2301 );
nand \U$24229 ( \24606 , \24604 , \24605 );
not \U$24230 ( \24607 , \24606 );
or \U$24231 ( \24608 , \24601 , \24607 );
nand \U$24232 ( \24609 , \24439 , \2320 );
nand \U$24233 ( \24610 , \24608 , \24609 );
xor \U$24234 ( \24611 , \24600 , \24610 );
xor \U$24235 ( \24612 , \24546 , \24557 );
and \U$24236 ( \24613 , \24612 , \24568 );
and \U$24237 ( \24614 , \24546 , \24557 );
or \U$24238 ( \24615 , \24613 , \24614 );
xor \U$24239 ( \24616 , \24611 , \24615 );
xor \U$24240 ( \24617 , \24207 , \24230 );
and \U$24241 ( \24618 , \24617 , \24235 );
and \U$24242 ( \24619 , \24207 , \24230 );
or \U$24243 ( \24620 , \24618 , \24619 );
xor \U$24244 ( \24621 , \24616 , \24620 );
xor \U$24245 ( \24622 , \24569 , \24573 );
and \U$24246 ( \24623 , \24622 , \24578 );
and \U$24247 ( \24624 , \24569 , \24573 );
or \U$24248 ( \24625 , \24623 , \24624 );
xor \U$24249 ( \24626 , \24621 , \24625 );
not \U$24250 ( \24627 , \24626 );
xor \U$24251 ( \24628 , \24544 , \24579 );
and \U$24252 ( \24629 , \24628 , \24584 );
and \U$24253 ( \24630 , \24544 , \24579 );
or \U$24254 ( \24631 , \24629 , \24630 );
not \U$24255 ( \24632 , \24631 );
not \U$24256 ( \24633 , \24632 );
or \U$24257 ( \24634 , \24627 , \24633 );
not \U$24258 ( \24635 , \24626 );
nand \U$24259 ( \24636 , \24635 , \24631 );
nand \U$24260 ( \24637 , \24634 , \24636 );
not \U$24261 ( \24638 , \24376 );
not \U$24262 ( \24639 , \24259 );
or \U$24263 ( \24640 , \24638 , \24639 );
nand \U$24264 ( \24641 , \24640 , \24236 );
not \U$24265 ( \24642 , \24259 );
nand \U$24266 ( \24643 , \24642 , \24379 );
nand \U$24267 ( \24644 , \24641 , \24643 );
not \U$24268 ( \24645 , \24644 );
and \U$24269 ( \24646 , \24637 , \24645 );
not \U$24270 ( \24647 , \24637 );
and \U$24271 ( \24648 , \24647 , \24644 );
nor \U$24272 ( \24649 , \24646 , \24648 );
xnor \U$24273 ( \24650 , \24589 , \24649 );
not \U$24274 ( \24651 , \24173 );
not \U$24275 ( \24652 , \24390 );
or \U$24276 ( \24653 , \24651 , \24652 );
nand \U$24277 ( \24654 , \24653 , \24382 );
not \U$24278 ( \24655 , \24173 );
nand \U$24279 ( \24656 , \24655 , \24393 );
nand \U$24280 ( \24657 , \24654 , \24656 );
not \U$24281 ( \24658 , \24657 );
xor \U$24282 ( \24659 , \24208 , \24217 );
and \U$24283 ( \24660 , \24659 , \24229 );
and \U$24284 ( \24661 , \24208 , \24217 );
or \U$24285 ( \24662 , \24660 , \24661 );
not \U$24286 ( \24663 , \951 );
not \U$24287 ( \24664 , \24180 );
or \U$24288 ( \24665 , \24663 , \24664 );
not \U$24289 ( \24666 , RIc2273d0_5);
not \U$24290 ( \24667 , \17549 );
or \U$24291 ( \24668 , \24666 , \24667 );
nand \U$24292 ( \24669 , \23772 , \946 );
nand \U$24293 ( \24670 , \24668 , \24669 );
nand \U$24294 ( \24671 , \24670 , \954 );
nand \U$24295 ( \24672 , \24665 , \24671 );
not \U$24296 ( \24673 , \1082 );
and \U$24297 ( \24674 , \9859 , RIc2274c0_3);
not \U$24298 ( \24675 , \9859 );
and \U$24299 ( \24676 , \24675 , \2896 );
or \U$24300 ( \24677 , \24674 , \24676 );
not \U$24301 ( \24678 , \24677 );
or \U$24302 ( \24679 , \24673 , \24678 );
nand \U$24303 ( \24680 , \24204 , \1040 );
nand \U$24304 ( \24681 , \24679 , \24680 );
xor \U$24305 ( \24682 , \24672 , \24681 );
not \U$24306 ( \24683 , \1118 );
not \U$24307 ( \24684 , \24191 );
or \U$24308 ( \24685 , \24683 , \24684 );
not \U$24309 ( \24686 , RIc2272e0_7);
not \U$24310 ( \24687 , \5216 );
or \U$24311 ( \24688 , \24686 , \24687 );
nand \U$24312 ( \24689 , \5217 , \1139 );
nand \U$24313 ( \24690 , \24688 , \24689 );
nand \U$24314 ( \24691 , \24690 , \1121 );
nand \U$24315 ( \24692 , \24685 , \24691 );
xor \U$24316 ( \24693 , \24682 , \24692 );
xor \U$24317 ( \24694 , \24662 , \24693 );
xor \U$24318 ( \24695 , \24310 , \24321 );
and \U$24319 ( \24696 , \24695 , \24332 );
and \U$24320 ( \24697 , \24310 , \24321 );
or \U$24321 ( \24698 , \24696 , \24697 );
xor \U$24322 ( \24699 , \24694 , \24698 );
not \U$24323 ( \24700 , \24299 );
not \U$24324 ( \24701 , \24333 );
or \U$24325 ( \24702 , \24700 , \24701 );
or \U$24326 ( \24703 , \24333 , \24299 );
nand \U$24327 ( \24704 , \24703 , \24375 );
nand \U$24328 ( \24705 , \24702 , \24704 );
xor \U$24329 ( \24706 , \24699 , \24705 );
not \U$24330 ( \24707 , \9705 );
not \U$24331 ( \24708 , RIc2262f0_41);
not \U$24332 ( \24709 , \9491 );
or \U$24333 ( \24710 , \24708 , \24709 );
nand \U$24334 ( \24711 , \1072 , \6303 );
nand \U$24335 ( \24712 , \24710 , \24711 );
not \U$24336 ( \24713 , \24712 );
or \U$24337 ( \24714 , \24707 , \24713 );
nand \U$24338 ( \24715 , \24473 , \9690 );
nand \U$24339 ( \24716 , \24714 , \24715 );
not \U$24340 ( \24717 , \5519 );
not \U$24341 ( \24718 , RIc2264d0_37);
not \U$24342 ( \24719 , \11714 );
or \U$24343 ( \24720 , \24718 , \24719 );
nand \U$24344 ( \24721 , \1454 , \4371 );
nand \U$24345 ( \24722 , \24720 , \24721 );
not \U$24346 ( \24723 , \24722 );
or \U$24347 ( \24724 , \24717 , \24723 );
nand \U$24348 ( \24725 , \24451 , \5509 );
nand \U$24349 ( \24726 , \24724 , \24725 );
xor \U$24350 ( \24727 , \24716 , \24726 );
not \U$24351 ( \24728 , \2154 );
not \U$24352 ( \24729 , RIc226980_27);
not \U$24353 ( \24730 , \3686 );
or \U$24354 ( \24731 , \24729 , \24730 );
nand \U$24355 ( \24732 , \2423 , \16510 );
nand \U$24356 ( \24733 , \24731 , \24732 );
not \U$24357 ( \24734 , \24733 );
or \U$24358 ( \24735 , \24728 , \24734 );
nand \U$24359 ( \24736 , \24354 , \2138 );
nand \U$24360 ( \24737 , \24735 , \24736 );
xor \U$24361 ( \24738 , \24727 , \24737 );
not \U$24362 ( \24739 , \3631 );
not \U$24363 ( \24740 , RIc2266b0_33);
not \U$24364 ( \24741 , \1530 );
or \U$24365 ( \24742 , \24740 , \24741 );
nand \U$24366 ( \24743 , \3579 , \2692 );
nand \U$24367 ( \24744 , \24742 , \24743 );
not \U$24368 ( \24745 , \24744 );
or \U$24369 ( \24746 , \24739 , \24745 );
nand \U$24370 ( \24747 , \24269 , \3629 );
nand \U$24371 ( \24748 , \24746 , \24747 );
not \U$24372 ( \24749 , \6689 );
not \U$24373 ( \24750 , \24346 );
or \U$24374 ( \24751 , \24749 , \24750 );
not \U$24375 ( \24752 , RIc2263e0_39);
not \U$24376 ( \24753 , \2178 );
or \U$24377 ( \24754 , \24752 , \24753 );
nand \U$24378 ( \24755 , \840 , \8998 );
nand \U$24379 ( \24756 , \24754 , \24755 );
nand \U$24380 ( \24757 , \24756 , \6307 );
nand \U$24381 ( \24758 , \24751 , \24757 );
xor \U$24382 ( \24759 , \24748 , \24758 );
not \U$24383 ( \24760 , \2367 );
not \U$24384 ( \24761 , RIc226c50_21);
not \U$24385 ( \24762 , \3292 );
or \U$24386 ( \24763 , \24761 , \24762 );
nand \U$24387 ( \24764 , \2593 , \3204 );
nand \U$24388 ( \24765 , \24763 , \24764 );
not \U$24389 ( \24766 , \24765 );
or \U$24390 ( \24767 , \24760 , \24766 );
nand \U$24391 ( \24768 , \24319 , \2392 );
nand \U$24392 ( \24769 , \24767 , \24768 );
xor \U$24393 ( \24770 , \24759 , \24769 );
xor \U$24394 ( \24771 , \24738 , \24770 );
not \U$24395 ( \24772 , \2711 );
and \U$24396 ( \24773 , \3044 , RIc2267a0_31);
not \U$24397 ( \24774 , \3044 );
and \U$24398 ( \24775 , \24774 , \2705 );
or \U$24399 ( \24776 , \24773 , \24775 );
not \U$24400 ( \24777 , \24776 );
or \U$24401 ( \24778 , \24772 , \24777 );
nand \U$24402 ( \24779 , \24225 , \2697 );
nand \U$24403 ( \24780 , \24778 , \24779 );
not \U$24404 ( \24781 , \1945 );
not \U$24405 ( \24782 , \24290 );
or \U$24406 ( \24783 , \24781 , \24782 );
not \U$24407 ( \24784 , RIc226e30_17);
not \U$24408 ( \24785 , \3810 );
or \U$24409 ( \24786 , \24784 , \24785 );
nand \U$24410 ( \24787 , \2720 , \1960 );
nand \U$24411 ( \24788 , \24786 , \24787 );
nand \U$24412 ( \24789 , \24788 , \1963 );
nand \U$24413 ( \24790 , \24783 , \24789 );
xor \U$24414 ( \24791 , \24780 , \24790 );
not \U$24415 ( \24792 , \2534 );
and \U$24416 ( \24793 , RIc226d40_19, \5819 );
not \U$24417 ( \24794 , RIc226d40_19);
and \U$24418 ( \24795 , \24794 , \2480 );
or \U$24419 ( \24796 , \24793 , \24795 );
not \U$24420 ( \24797 , \24796 );
or \U$24421 ( \24798 , \24792 , \24797 );
nand \U$24422 ( \24799 , \24281 , \2518 );
nand \U$24423 ( \24800 , \24798 , \24799 );
xor \U$24424 ( \24801 , \24791 , \24800 );
xor \U$24425 ( \24802 , \24771 , \24801 );
xor \U$24426 ( \24803 , \24706 , \24802 );
not \U$24427 ( \24804 , \24247 );
not \U$24428 ( \24805 , \24241 );
or \U$24429 ( \24806 , \24804 , \24805 );
or \U$24430 ( \24807 , \24241 , \24247 );
nand \U$24431 ( \24808 , \24807 , \24252 );
nand \U$24432 ( \24809 , \24806 , \24808 );
not \U$24433 ( \24810 , \24809 );
not \U$24434 ( \24811 , \24475 );
not \U$24435 ( \24812 , \24465 );
or \U$24436 ( \24813 , \24811 , \24812 );
or \U$24437 ( \24814 , \24465 , \24475 );
nand \U$24438 ( \24815 , \24814 , \24453 );
nand \U$24439 ( \24816 , \24813 , \24815 );
not \U$24440 ( \24817 , \24370 );
not \U$24441 ( \24818 , \24358 );
or \U$24442 ( \24819 , \24817 , \24818 );
or \U$24443 ( \24820 , \24358 , \24370 );
nand \U$24444 ( \24821 , \24820 , \24348 );
nand \U$24445 ( \24822 , \24819 , \24821 );
xor \U$24446 ( \24823 , \24816 , \24822 );
not \U$24447 ( \24824 , \24420 );
not \U$24448 ( \24825 , \24430 );
or \U$24449 ( \24826 , \24824 , \24825 );
or \U$24450 ( \24827 , \24430 , \24420 );
nand \U$24451 ( \24828 , \24827 , \24441 );
nand \U$24452 ( \24829 , \24826 , \24828 );
xnor \U$24453 ( \24830 , \24823 , \24829 );
not \U$24454 ( \24831 , \24830 );
or \U$24455 ( \24832 , \24810 , \24831 );
or \U$24456 ( \24833 , \24809 , \24830 );
nand \U$24457 ( \24834 , \24832 , \24833 );
xor \U$24458 ( \24835 , \24185 , \24195 );
and \U$24459 ( \24836 , \24835 , \24206 );
and \U$24460 ( \24837 , \24185 , \24195 );
or \U$24461 ( \24838 , \24836 , \24837 );
and \U$24462 ( \24839 , RIc2275b0_1, \20216 );
and \U$24463 ( \24840 , \24418 , \9110 );
not \U$24464 ( \24841 , \9129 );
nor \U$24465 ( \24842 , \24841 , \9106 );
nor \U$24466 ( \24843 , \24840 , \24842 );
not \U$24467 ( \24844 , \24843 );
xor \U$24468 ( \24845 , \24839 , \24844 );
not \U$24469 ( \24846 , \1579 );
xor \U$24470 ( \24847 , RIc2275b0_1, \8886 );
not \U$24471 ( \24848 , \24847 );
or \U$24472 ( \24849 , \24846 , \24848 );
nand \U$24473 ( \24850 , \24213 , \854 );
nand \U$24474 ( \24851 , \24849 , \24850 );
xnor \U$24475 ( \24852 , \24845 , \24851 );
xor \U$24476 ( \24853 , \24838 , \24852 );
or \U$24477 ( \24854 , \24294 , \24273 );
nand \U$24478 ( \24855 , \24854 , \24283 );
nand \U$24479 ( \24856 , \24294 , \24273 );
and \U$24480 ( \24857 , \24855 , \24856 );
xnor \U$24481 ( \24858 , \24853 , \24857 );
and \U$24482 ( \24859 , \24834 , \24858 );
not \U$24483 ( \24860 , \24834 );
not \U$24484 ( \24861 , \24858 );
and \U$24485 ( \24862 , \24860 , \24861 );
nor \U$24486 ( \24863 , \24859 , \24862 );
and \U$24487 ( \24864 , \24803 , \24863 );
not \U$24488 ( \24865 , \24803 );
not \U$24489 ( \24866 , \24863 );
and \U$24490 ( \24867 , \24865 , \24866 );
or \U$24491 ( \24868 , \24864 , \24867 );
not \U$24492 ( \24869 , \2086 );
xnor \U$24493 ( \24870 , RIc226890_29, \9700 );
not \U$24494 ( \24871 , \24870 );
or \U$24495 ( \24872 , \24869 , \24871 );
nand \U$24496 ( \24873 , \24368 , \2784 );
nand \U$24497 ( \24874 , \24872 , \24873 );
not \U$24498 ( \24875 , \1311 );
not \U$24499 ( \24876 , RIc227100_11);
not \U$24500 ( \24877 , \11672 );
or \U$24501 ( \24878 , \24876 , \24877 );
nand \U$24502 ( \24879 , \2981 , \1291 );
nand \U$24503 ( \24880 , \24878 , \24879 );
not \U$24504 ( \24881 , \24880 );
or \U$24505 ( \24882 , \24875 , \24881 );
nand \U$24506 ( \24883 , \24564 , \1307 );
nand \U$24507 ( \24884 , \24882 , \24883 );
xor \U$24508 ( \24885 , \24874 , \24884 );
not \U$24509 ( \24886 , \1682 );
not \U$24510 ( \24887 , RIc227010_13);
not \U$24511 ( \24888 , \23889 );
or \U$24512 ( \24889 , \24887 , \24888 );
nand \U$24513 ( \24890 , \4501 , \1296 );
nand \U$24514 ( \24891 , \24889 , \24890 );
not \U$24515 ( \24892 , \24891 );
or \U$24516 ( \24893 , \24886 , \24892 );
nand \U$24517 ( \24894 , \24426 , \3250 );
nand \U$24518 ( \24895 , \24893 , \24894 );
xor \U$24519 ( \24896 , \24885 , \24895 );
not \U$24520 ( \24897 , \2172 );
not \U$24521 ( \24898 , RIc226a70_25);
not \U$24522 ( \24899 , \2234 );
or \U$24523 ( \24900 , \24898 , \24899 );
nand \U$24524 ( \24901 , \18087 , \3982 );
nand \U$24525 ( \24902 , \24900 , \24901 );
not \U$24526 ( \24903 , \24902 );
or \U$24527 ( \24904 , \24897 , \24903 );
nand \U$24528 ( \24905 , \24463 , \2860 );
nand \U$24529 ( \24906 , \24904 , \24905 );
not \U$24530 ( \24907 , \5135 );
not \U$24531 ( \24908 , RIc2265c0_35);
not \U$24532 ( \24909 , \1372 );
or \U$24533 ( \24910 , \24908 , \24909 );
nand \U$24534 ( \24911 , \2373 , \3620 );
nand \U$24535 ( \24912 , \24910 , \24911 );
not \U$24536 ( \24913 , \24912 );
or \U$24537 ( \24914 , \24907 , \24913 );
nand \U$24538 ( \24915 , \24328 , \5741 );
nand \U$24539 ( \24916 , \24914 , \24915 );
xor \U$24540 ( \24917 , \24906 , \24916 );
not \U$24541 ( \24918 , \1930 );
not \U$24542 ( \24919 , RIc226b60_23);
not \U$24543 ( \24920 , \5768 );
or \U$24544 ( \24921 , \24919 , \24920 );
nand \U$24545 ( \24922 , \3840 , \2111 );
nand \U$24546 ( \24923 , \24921 , \24922 );
not \U$24547 ( \24924 , \24923 );
or \U$24548 ( \24925 , \24918 , \24924 );
nand \U$24549 ( \24926 , \24306 , \1915 );
nand \U$24550 ( \24927 , \24925 , \24926 );
xor \U$24551 ( \24928 , \24917 , \24927 );
xor \U$24552 ( \24929 , \24896 , \24928 );
xor \U$24553 ( \24930 , \24505 , \24509 );
and \U$24554 ( \24931 , \24930 , \24517 );
and \U$24555 ( \24932 , \24505 , \24509 );
or \U$24556 ( \24933 , \24931 , \24932 );
xor \U$24557 ( \24934 , \24929 , \24933 );
not \U$24558 ( \24935 , \24934 );
not \U$24559 ( \24936 , \24480 );
nand \U$24560 ( \24937 , \24936 , \24442 );
and \U$24561 ( \24938 , \24937 , \24489 );
nor \U$24562 ( \24939 , \24442 , \24483 );
nor \U$24563 ( \24940 , \24938 , \24939 );
not \U$24564 ( \24941 , \24940 );
and \U$24565 ( \24942 , \24935 , \24941 );
and \U$24566 ( \24943 , \24934 , \24940 );
nor \U$24567 ( \24944 , \24942 , \24943 );
xor \U$24568 ( \24945 , \24518 , \24525 );
and \U$24569 ( \24946 , \24945 , \24530 );
and \U$24570 ( \24947 , \24518 , \24525 );
or \U$24571 ( \24948 , \24946 , \24947 );
and \U$24572 ( \24949 , \24944 , \24948 );
not \U$24573 ( \24950 , \24944 );
not \U$24574 ( \24951 , \24948 );
and \U$24575 ( \24952 , \24950 , \24951 );
nor \U$24576 ( \24953 , \24949 , \24952 );
and \U$24577 ( \24954 , \24868 , \24953 );
not \U$24578 ( \24955 , \24868 );
not \U$24579 ( \24956 , \24953 );
and \U$24580 ( \24957 , \24955 , \24956 );
nor \U$24581 ( \24958 , \24954 , \24957 );
not \U$24582 ( \24959 , \24958 );
or \U$24583 ( \24960 , \24658 , \24959 );
or \U$24584 ( \24961 , \24657 , \24958 );
nand \U$24585 ( \24962 , \24960 , \24961 );
xor \U$24586 ( \24963 , \24490 , \24496 );
xor \U$24587 ( \24964 , \24963 , \24501 );
not \U$24588 ( \24965 , \24964 );
xor \U$24589 ( \24966 , \24531 , \24537 );
xor \U$24590 ( \24967 , \24966 , \24585 );
not \U$24591 ( \24968 , \24967 );
or \U$24592 ( \24969 , \24965 , \24968 );
or \U$24593 ( \24970 , \24967 , \24964 );
buf \U$24594 ( \24971 , \23079 );
not \U$24595 ( \24972 , \24971 );
not \U$24596 ( \24973 , \22683 );
or \U$24597 ( \24974 , \24972 , \24973 );
or \U$24598 ( \24975 , \24971 , \22683 );
not \U$24599 ( \24976 , \22960 );
nand \U$24600 ( \24977 , \24975 , \24976 );
nand \U$24601 ( \24978 , \24974 , \24977 );
nand \U$24602 ( \24979 , \24970 , \24978 );
nand \U$24603 ( \24980 , \24969 , \24979 );
and \U$24604 ( \24981 , \24962 , \24980 );
not \U$24605 ( \24982 , \24962 );
not \U$24606 ( \24983 , \24980 );
and \U$24607 ( \24984 , \24982 , \24983 );
nor \U$24608 ( \24985 , \24981 , \24984 );
xor \U$24609 ( \24986 , \24650 , \24985 );
xor \U$24610 ( \24987 , \24410 , \24986 );
xnor \U$24611 ( \24988 , \24978 , \24964 );
xnor \U$24612 ( \24989 , \24988 , \24967 );
not \U$24613 ( \24990 , \24405 );
xor \U$24614 ( \24991 , \24163 , \24395 );
not \U$24615 ( \24992 , \24991 );
or \U$24616 ( \24993 , \24990 , \24992 );
or \U$24617 ( \24994 , \24991 , \24405 );
nand \U$24618 ( \24995 , \24993 , \24994 );
xor \U$24619 ( \24996 , \24989 , \24995 );
xor \U$24620 ( \24997 , \23985 , \23989 );
and \U$24621 ( \24998 , \24997 , \23994 );
and \U$24622 ( \24999 , \23985 , \23989 );
or \U$24623 ( \25000 , \24998 , \24999 );
and \U$24624 ( \25001 , \24996 , \25000 );
and \U$24625 ( \25002 , \24989 , \24995 );
or \U$24626 ( \25003 , \25001 , \25002 );
or \U$24627 ( \25004 , \24987 , \25003 );
xor \U$24628 ( \25005 , \24989 , \24995 );
xor \U$24629 ( \25006 , \25005 , \25000 );
not \U$24630 ( \25007 , \25006 );
or \U$24631 ( \25008 , \23995 , \23478 );
nand \U$24632 ( \25009 , \25008 , \23735 );
nand \U$24633 ( \25010 , \23995 , \23478 );
nand \U$24634 ( \25011 , \25009 , \25010 );
not \U$24635 ( \25012 , \25011 );
nand \U$24636 ( \25013 , \25007 , \25012 );
nand \U$24637 ( \25014 , \25004 , \25013 );
not \U$24638 ( \25015 , \24934 );
nand \U$24639 ( \25016 , \25015 , \24940 );
not \U$24640 ( \25017 , \25016 );
not \U$24641 ( \25018 , \24948 );
or \U$24642 ( \25019 , \25017 , \25018 );
not \U$24643 ( \25020 , \24940 );
nand \U$24644 ( \25021 , \25020 , \24934 );
nand \U$24645 ( \25022 , \25019 , \25021 );
not \U$24646 ( \25023 , \24626 );
not \U$24647 ( \25024 , \24631 );
or \U$24648 ( \25025 , \25023 , \25024 );
not \U$24649 ( \25026 , \24626 );
nand \U$24650 ( \25027 , \25026 , \24632 );
nand \U$24651 ( \25028 , \24644 , \25027 );
nand \U$24652 ( \25029 , \25025 , \25028 );
xor \U$24653 ( \25030 , \25022 , \25029 );
not \U$24654 ( \25031 , \24861 );
buf \U$24655 ( \25032 , \24830 );
not \U$24656 ( \25033 , \25032 );
not \U$24657 ( \25034 , \25033 );
or \U$24658 ( \25035 , \25031 , \25034 );
not \U$24659 ( \25036 , \24858 );
not \U$24660 ( \25037 , \25032 );
or \U$24661 ( \25038 , \25036 , \25037 );
nand \U$24662 ( \25039 , \25038 , \24809 );
nand \U$24663 ( \25040 , \25035 , \25039 );
not \U$24664 ( \25041 , \24839 );
nand \U$24665 ( \25042 , \25041 , \24843 );
not \U$24666 ( \25043 , \25042 );
not \U$24667 ( \25044 , \24851 );
or \U$24668 ( \25045 , \25043 , \25044 );
nand \U$24669 ( \25046 , \24844 , \24839 );
nand \U$24670 ( \25047 , \25045 , \25046 );
xor \U$24671 ( \25048 , \24672 , \24681 );
and \U$24672 ( \25049 , \25048 , \24692 );
and \U$24673 ( \25050 , \24672 , \24681 );
or \U$24674 ( \25051 , \25049 , \25050 );
xor \U$24675 ( \25052 , \25047 , \25051 );
not \U$24676 ( \25053 , \1082 );
and \U$24677 ( \25054 , \6493 , RIc2274c0_3);
not \U$24678 ( \25055 , \6493 );
and \U$24679 ( \25056 , \25055 , \1032 );
or \U$24680 ( \25057 , \25054 , \25056 );
not \U$24681 ( \25058 , \25057 );
or \U$24682 ( \25059 , \25053 , \25058 );
nand \U$24683 ( \25060 , \24677 , \1040 );
nand \U$24684 ( \25061 , \25059 , \25060 );
not \U$24685 ( \25062 , \954 );
not \U$24686 ( \25063 , RIc2273d0_5);
not \U$24687 ( \25064 , \5665 );
or \U$24688 ( \25065 , \25063 , \25064 );
nand \U$24689 ( \25066 , \19859 , \946 );
nand \U$24690 ( \25067 , \25065 , \25066 );
not \U$24691 ( \25068 , \25067 );
or \U$24692 ( \25069 , \25062 , \25068 );
nand \U$24693 ( \25070 , \24670 , \951 );
nand \U$24694 ( \25071 , \25069 , \25070 );
xor \U$24695 ( \25072 , \25061 , \25071 );
not \U$24696 ( \25073 , \854 );
not \U$24697 ( \25074 , \24847 );
or \U$24698 ( \25075 , \25073 , \25074 );
and \U$24699 ( \25076 , RIc2275b0_1, \15699 );
not \U$24700 ( \25077 , RIc2275b0_1);
and \U$24701 ( \25078 , \25077 , \20646 );
or \U$24702 ( \25079 , \25076 , \25078 );
nand \U$24703 ( \25080 , \25079 , \1579 );
nand \U$24704 ( \25081 , \25075 , \25080 );
xor \U$24705 ( \25082 , \25072 , \25081 );
xor \U$24706 ( \25083 , \25052 , \25082 );
buf \U$24707 ( \25084 , \24816 );
not \U$24708 ( \25085 , \25084 );
not \U$24709 ( \25086 , \24829 );
or \U$24710 ( \25087 , \25085 , \25086 );
or \U$24711 ( \25088 , \24829 , \25084 );
nand \U$24712 ( \25089 , \25088 , \24822 );
nand \U$24713 ( \25090 , \25087 , \25089 );
xor \U$24714 ( \25091 , \25083 , \25090 );
xor \U$24715 ( \25092 , \24738 , \24770 );
and \U$24716 ( \25093 , \25092 , \24801 );
and \U$24717 ( \25094 , \24738 , \24770 );
or \U$24718 ( \25095 , \25093 , \25094 );
xor \U$24719 ( \25096 , \25091 , \25095 );
not \U$24720 ( \25097 , \25096 );
and \U$24721 ( \25098 , \25040 , \25097 );
not \U$24722 ( \25099 , \25040 );
and \U$24723 ( \25100 , \25099 , \25096 );
or \U$24724 ( \25101 , \25098 , \25100 );
xor \U$24725 ( \25102 , \24600 , \24610 );
and \U$24726 ( \25103 , \25102 , \24615 );
and \U$24727 ( \25104 , \24600 , \24610 );
or \U$24728 ( \25105 , \25103 , \25104 );
not \U$24729 ( \25106 , \24838 );
nand \U$24730 ( \25107 , \25106 , \24852 );
not \U$24731 ( \25108 , \25107 );
not \U$24732 ( \25109 , \24857 );
not \U$24733 ( \25110 , \25109 );
or \U$24734 ( \25111 , \25108 , \25110 );
not \U$24735 ( \25112 , \24852 );
nand \U$24736 ( \25113 , \25112 , \24838 );
nand \U$24737 ( \25114 , \25111 , \25113 );
xor \U$24738 ( \25115 , \25105 , \25114 );
xor \U$24739 ( \25116 , \24662 , \24693 );
and \U$24740 ( \25117 , \25116 , \24698 );
and \U$24741 ( \25118 , \24662 , \24693 );
or \U$24742 ( \25119 , \25117 , \25118 );
xnor \U$24743 ( \25120 , \25115 , \25119 );
and \U$24744 ( \25121 , \25101 , \25120 );
not \U$24745 ( \25122 , \25101 );
not \U$24746 ( \25123 , \25120 );
and \U$24747 ( \25124 , \25122 , \25123 );
nor \U$24748 ( \25125 , \25121 , \25124 );
not \U$24749 ( \25126 , \25125 );
xnor \U$24750 ( \25127 , \25030 , \25126 );
not \U$24751 ( \25128 , \24866 );
not \U$24752 ( \25129 , \24803 );
not \U$24753 ( \25130 , \25129 );
not \U$24754 ( \25131 , \25130 );
or \U$24755 ( \25132 , \25128 , \25131 );
not \U$24756 ( \25133 , \25129 );
not \U$24757 ( \25134 , \24863 );
or \U$24758 ( \25135 , \25133 , \25134 );
nand \U$24759 ( \25136 , \25135 , \24956 );
nand \U$24760 ( \25137 , \25132 , \25136 );
not \U$24761 ( \25138 , \25137 );
not \U$24762 ( \25139 , \25138 );
xor \U$24763 ( \25140 , \24699 , \24705 );
and \U$24764 ( \25141 , \25140 , \24802 );
and \U$24765 ( \25142 , \24699 , \24705 );
or \U$24766 ( \25143 , \25141 , \25142 );
or \U$24767 ( \25144 , \9110 , \9129 );
nand \U$24768 ( \25145 , \25144 , RIc226200_43);
not \U$24769 ( \25146 , \1121 );
not \U$24770 ( \25147 , RIc2272e0_7);
not \U$24771 ( \25148 , \18450 );
or \U$24772 ( \25149 , \25147 , \25148 );
nand \U$24773 ( \25150 , \22991 , \940 );
nand \U$24774 ( \25151 , \25149 , \25150 );
not \U$24775 ( \25152 , \25151 );
or \U$24776 ( \25153 , \25146 , \25152 );
nand \U$24777 ( \25154 , \24690 , \1118 );
nand \U$24778 ( \25155 , \25153 , \25154 );
xor \U$24779 ( \25156 , \25145 , \25155 );
not \U$24780 ( \25157 , \1340 );
not \U$24781 ( \25158 , RIc2271f0_9);
not \U$24782 ( \25159 , \19926 );
or \U$24783 ( \25160 , \25158 , \25159 );
nand \U$24784 ( \25161 , \3641 , \1351 );
nand \U$24785 ( \25162 , \25160 , \25161 );
not \U$24786 ( \25163 , \25162 );
or \U$24787 ( \25164 , \25157 , \25163 );
nand \U$24788 ( \25165 , \24597 , \1597 );
nand \U$24789 ( \25166 , \25164 , \25165 );
xor \U$24790 ( \25167 , \25156 , \25166 );
xor \U$24791 ( \25168 , \24874 , \24884 );
and \U$24792 ( \25169 , \25168 , \24895 );
and \U$24793 ( \25170 , \24874 , \24884 );
or \U$24794 ( \25171 , \25169 , \25170 );
xor \U$24795 ( \25172 , \25167 , \25171 );
xor \U$24796 ( \25173 , \24780 , \24790 );
and \U$24797 ( \25174 , \25173 , \24800 );
and \U$24798 ( \25175 , \24780 , \24790 );
or \U$24799 ( \25176 , \25174 , \25175 );
xor \U$24800 ( \25177 , \25172 , \25176 );
xor \U$24801 ( \25178 , \24748 , \24758 );
and \U$24802 ( \25179 , \25178 , \24769 );
and \U$24803 ( \25180 , \24748 , \24758 );
or \U$24804 ( \25181 , \25179 , \25180 );
xor \U$24805 ( \25182 , \24906 , \24916 );
and \U$24806 ( \25183 , \25182 , \24927 );
and \U$24807 ( \25184 , \24906 , \24916 );
or \U$24808 ( \25185 , \25183 , \25184 );
not \U$24809 ( \25186 , \25185 );
and \U$24810 ( \25187 , \25181 , \25186 );
not \U$24811 ( \25188 , \25181 );
and \U$24812 ( \25189 , \25188 , \25185 );
or \U$24813 ( \25190 , \25187 , \25189 );
or \U$24814 ( \25191 , \24726 , \24716 );
and \U$24815 ( \25192 , \25191 , \24737 );
and \U$24816 ( \25193 , \24716 , \24726 );
nor \U$24817 ( \25194 , \25192 , \25193 );
not \U$24818 ( \25195 , \25194 );
and \U$24819 ( \25196 , \25190 , \25195 );
not \U$24820 ( \25197 , \25190 );
and \U$24821 ( \25198 , \25197 , \25194 );
nor \U$24822 ( \25199 , \25196 , \25198 );
xor \U$24823 ( \25200 , \25177 , \25199 );
xor \U$24824 ( \25201 , \24896 , \24928 );
and \U$24825 ( \25202 , \25201 , \24933 );
and \U$24826 ( \25203 , \24896 , \24928 );
or \U$24827 ( \25204 , \25202 , \25203 );
and \U$24828 ( \25205 , \25200 , \25204 );
not \U$24829 ( \25206 , \25200 );
not \U$24830 ( \25207 , \25204 );
and \U$24831 ( \25208 , \25206 , \25207 );
nor \U$24832 ( \25209 , \25205 , \25208 );
xor \U$24833 ( \25210 , \25143 , \25209 );
not \U$24834 ( \25211 , \1963 );
not \U$24835 ( \25212 , RIc226e30_17);
not \U$24836 ( \25213 , \12989 );
or \U$24837 ( \25214 , \25212 , \25213 );
not \U$24838 ( \25215 , \4195 );
nand \U$24839 ( \25216 , \25215 , \1952 );
nand \U$24840 ( \25217 , \25214 , \25216 );
not \U$24841 ( \25218 , \25217 );
or \U$24842 ( \25219 , \25211 , \25218 );
nand \U$24843 ( \25220 , \24788 , \1945 );
nand \U$24844 ( \25221 , \25219 , \25220 );
xor \U$24845 ( \25222 , \24599 , \25221 );
not \U$24846 ( \25223 , \2320 );
not \U$24847 ( \25224 , \24606 );
or \U$24848 ( \25225 , \25223 , \25224 );
not \U$24849 ( \25226 , RIc226f20_15);
not \U$24850 ( \25227 , \4240 );
not \U$24851 ( \25228 , \25227 );
or \U$24852 ( \25229 , \25226 , \25228 );
nand \U$24853 ( \25230 , \23331 , \2301 );
nand \U$24854 ( \25231 , \25229 , \25230 );
nand \U$24855 ( \25232 , \25231 , \2358 );
nand \U$24856 ( \25233 , \25225 , \25232 );
xor \U$24857 ( \25234 , \25222 , \25233 );
not \U$24858 ( \25235 , RIc2275b0_1);
nor \U$24859 ( \25236 , \25235 , \12724 );
not \U$24860 ( \25237 , \2086 );
and \U$24861 ( \25238 , RIc226890_29, \2615 );
not \U$24862 ( \25239 , RIc226890_29);
and \U$24863 ( \25240 , \25239 , \1730 );
or \U$24864 ( \25241 , \25238 , \25240 );
not \U$24865 ( \25242 , \25241 );
or \U$24866 ( \25243 , \25237 , \25242 );
nand \U$24867 ( \25244 , \24870 , \2078 );
nand \U$24868 ( \25245 , \25243 , \25244 );
xor \U$24869 ( \25246 , \25236 , \25245 );
not \U$24870 ( \25247 , \3250 );
not \U$24871 ( \25248 , \24891 );
or \U$24872 ( \25249 , \25247 , \25248 );
not \U$24873 ( \25250 , RIc227010_13);
not \U$24874 ( \25251 , \3564 );
or \U$24875 ( \25252 , \25250 , \25251 );
nand \U$24876 ( \25253 , \2636 , \2427 );
nand \U$24877 ( \25254 , \25252 , \25253 );
nand \U$24878 ( \25255 , \25254 , \1682 );
nand \U$24879 ( \25256 , \25249 , \25255 );
xor \U$24880 ( \25257 , \25246 , \25256 );
xor \U$24881 ( \25258 , \25234 , \25257 );
not \U$24882 ( \25259 , \5135 );
and \U$24883 ( \25260 , \1404 , RIc2265c0_35);
not \U$24884 ( \25261 , \1404 );
and \U$24885 ( \25262 , \25261 , \16314 );
or \U$24886 ( \25263 , \25260 , \25262 );
not \U$24887 ( \25264 , \25263 );
or \U$24888 ( \25265 , \25259 , \25264 );
nand \U$24889 ( \25266 , \24912 , \5741 );
nand \U$24890 ( \25267 , \25265 , \25266 );
not \U$24891 ( \25268 , \5509 );
not \U$24892 ( \25269 , \24722 );
or \U$24893 ( \25270 , \25268 , \25269 );
not \U$24894 ( \25271 , RIc2264d0_37);
not \U$24895 ( \25272 , \1559 );
or \U$24896 ( \25273 , \25271 , \25272 );
nand \U$24897 ( \25274 , \984 , \12522 );
nand \U$24898 ( \25275 , \25273 , \25274 );
nand \U$24899 ( \25276 , \25275 , \5519 );
nand \U$24900 ( \25277 , \25270 , \25276 );
xor \U$24901 ( \25278 , \25267 , \25277 );
not \U$24902 ( \25279 , \2173 );
not \U$24903 ( \25280 , RIc226a70_25);
not \U$24904 ( \25281 , \2834 );
or \U$24905 ( \25282 , \25280 , \25281 );
not \U$24906 ( \25283 , \5270 );
nand \U$24907 ( \25284 , \25283 , \1905 );
nand \U$24908 ( \25285 , \25282 , \25284 );
not \U$24909 ( \25286 , \25285 );
or \U$24910 ( \25287 , \25279 , \25286 );
nand \U$24911 ( \25288 , \24902 , \2195 );
nand \U$24912 ( \25289 , \25287 , \25288 );
xor \U$24913 ( \25290 , \25278 , \25289 );
xor \U$24914 ( \25291 , \25258 , \25290 );
and \U$24915 ( \25292 , \9573 , \891 );
not \U$24916 ( \25293 , \9573 );
and \U$24917 ( \25294 , \25293 , \2865 );
nor \U$24918 ( \25295 , \25292 , \25294 );
not \U$24919 ( \25296 , \25295 );
not \U$24920 ( \25297 , \6308 );
and \U$24921 ( \25298 , \25296 , \25297 );
not \U$24922 ( \25299 , \24756 );
nor \U$24923 ( \25300 , \25299 , \17125 );
nor \U$24924 ( \25301 , \25298 , \25300 );
not \U$24925 ( \25302 , RIc226b60_23);
not \U$24926 ( \25303 , \2258 );
or \U$24927 ( \25304 , \25302 , \25303 );
nand \U$24928 ( \25305 , \2261 , \1919 );
nand \U$24929 ( \25306 , \25304 , \25305 );
and \U$24930 ( \25307 , \1930 , \25306 );
and \U$24931 ( \25308 , \24923 , \1915 );
nor \U$24932 ( \25309 , \25307 , \25308 );
xor \U$24933 ( \25310 , \25301 , \25309 );
not \U$24934 ( \25311 , \24744 );
nor \U$24935 ( \25312 , \25311 , \5185 );
and \U$24936 ( \25313 , \9943 , \22319 );
not \U$24937 ( \25314 , \9943 );
and \U$24938 ( \25315 , \25314 , \1393 );
nor \U$24939 ( \25316 , \25313 , \25315 );
nor \U$24940 ( \25317 , \25316 , \4440 );
nor \U$24941 ( \25318 , \25312 , \25317 );
xor \U$24942 ( \25319 , \25310 , \25318 );
not \U$24943 ( \25320 , \2711 );
not \U$24944 ( \25321 , RIc2267a0_31);
not \U$24945 ( \25322 , \1333 );
or \U$24946 ( \25323 , \25321 , \25322 );
nand \U$24947 ( \25324 , \3918 , \6902 );
nand \U$24948 ( \25325 , \25323 , \25324 );
not \U$24949 ( \25326 , \25325 );
or \U$24950 ( \25327 , \25320 , \25326 );
nand \U$24951 ( \25328 , \24776 , \2697 );
nand \U$24952 ( \25329 , \25327 , \25328 );
not \U$24953 ( \25330 , \2367 );
not \U$24954 ( \25331 , RIc226c50_21);
not \U$24955 ( \25332 , \2015 );
or \U$24956 ( \25333 , \25331 , \25332 );
nand \U$24957 ( \25334 , \3508 , \2370 );
nand \U$24958 ( \25335 , \25333 , \25334 );
not \U$24959 ( \25336 , \25335 );
or \U$24960 ( \25337 , \25330 , \25336 );
nand \U$24961 ( \25338 , \24765 , \2392 );
nand \U$24962 ( \25339 , \25337 , \25338 );
xor \U$24963 ( \25340 , \25329 , \25339 );
not \U$24964 ( \25341 , \2534 );
not \U$24965 ( \25342 , RIc226d40_19);
not \U$24966 ( \25343 , \3447 );
or \U$24967 ( \25344 , \25342 , \25343 );
nand \U$24968 ( \25345 , \3450 , \1941 );
nand \U$24969 ( \25346 , \25344 , \25345 );
not \U$24970 ( \25347 , \25346 );
or \U$24971 ( \25348 , \25341 , \25347 );
nand \U$24972 ( \25349 , \24796 , \2518 );
nand \U$24973 ( \25350 , \25348 , \25349 );
xor \U$24974 ( \25351 , \25340 , \25350 );
xor \U$24975 ( \25352 , \25319 , \25351 );
not \U$24976 ( \25353 , RIc2262f0_41);
not \U$24977 ( \25354 , \932 );
or \U$24978 ( \25355 , \25353 , \25354 );
not \U$24979 ( \25356 , \2701 );
nand \U$24980 ( \25357 , \25356 , \6303 );
nand \U$24981 ( \25358 , \25355 , \25357 );
not \U$24982 ( \25359 , \25358 );
not \U$24983 ( \25360 , \9816 );
or \U$24984 ( \25361 , \25359 , \25360 );
not \U$24985 ( \25362 , \24712 );
or \U$24986 ( \25363 , \25362 , \16459 );
nand \U$24987 ( \25364 , \25361 , \25363 );
not \U$24988 ( \25365 , \2138 );
not \U$24989 ( \25366 , \24733 );
or \U$24990 ( \25367 , \25365 , \25366 );
not \U$24991 ( \25368 , RIc226980_27);
not \U$24992 ( \25369 , \10936 );
or \U$24993 ( \25370 , \25368 , \25369 );
nand \U$24994 ( \25371 , \2305 , \2133 );
nand \U$24995 ( \25372 , \25370 , \25371 );
nand \U$24996 ( \25373 , \25372 , \2154 );
nand \U$24997 ( \25374 , \25367 , \25373 );
xor \U$24998 ( \25375 , \25364 , \25374 );
not \U$24999 ( \25376 , \1311 );
not \U$25000 ( \25377 , RIc227100_11);
not \U$25001 ( \25378 , \3121 );
or \U$25002 ( \25379 , \25377 , \25378 );
nand \U$25003 ( \25380 , \3122 , \1302 );
nand \U$25004 ( \25381 , \25379 , \25380 );
not \U$25005 ( \25382 , \25381 );
or \U$25006 ( \25383 , \25376 , \25382 );
nand \U$25007 ( \25384 , \24880 , \1307 );
nand \U$25008 ( \25385 , \25383 , \25384 );
xor \U$25009 ( \25386 , \25375 , \25385 );
xnor \U$25010 ( \25387 , \25352 , \25386 );
xor \U$25011 ( \25388 , \25291 , \25387 );
xor \U$25012 ( \25389 , \24616 , \24620 );
and \U$25013 ( \25390 , \25389 , \24625 );
and \U$25014 ( \25391 , \24616 , \24620 );
or \U$25015 ( \25392 , \25390 , \25391 );
xor \U$25016 ( \25393 , \25388 , \25392 );
xnor \U$25017 ( \25394 , \25210 , \25393 );
not \U$25018 ( \25395 , \25394 );
not \U$25019 ( \25396 , \25395 );
or \U$25020 ( \25397 , \25139 , \25396 );
nand \U$25021 ( \25398 , \25394 , \25137 );
nand \U$25022 ( \25399 , \25397 , \25398 );
not \U$25023 ( \25400 , \25399 );
not \U$25024 ( \25401 , \24504 );
not \U$25025 ( \25402 , \24649 );
not \U$25026 ( \25403 , \25402 );
or \U$25027 ( \25404 , \25401 , \25403 );
not \U$25028 ( \25405 , \24504 );
not \U$25029 ( \25406 , \25405 );
not \U$25030 ( \25407 , \24649 );
or \U$25031 ( \25408 , \25406 , \25407 );
nand \U$25032 ( \25409 , \25408 , \24588 );
nand \U$25033 ( \25410 , \25404 , \25409 );
not \U$25034 ( \25411 , \25410 );
not \U$25035 ( \25412 , \25411 );
and \U$25036 ( \25413 , \25400 , \25412 );
and \U$25037 ( \25414 , \25399 , \25411 );
nor \U$25038 ( \25415 , \25413 , \25414 );
xor \U$25039 ( \25416 , \25127 , \25415 );
not \U$25040 ( \25417 , \24983 );
buf \U$25041 ( \25418 , \24958 );
not \U$25042 ( \25419 , \25418 );
or \U$25043 ( \25420 , \25417 , \25419 );
nand \U$25044 ( \25421 , \25420 , \24657 );
not \U$25045 ( \25422 , \25418 );
nand \U$25046 ( \25423 , \25422 , \24980 );
and \U$25047 ( \25424 , \25421 , \25423 );
xor \U$25048 ( \25425 , \25416 , \25424 );
or \U$25049 ( \25426 , \24650 , \24985 );
and \U$25050 ( \25427 , \25426 , \24410 );
and \U$25051 ( \25428 , \24650 , \24985 );
nor \U$25052 ( \25429 , \25427 , \25428 );
nand \U$25053 ( \25430 , \25425 , \25429 );
xor \U$25054 ( \25431 , \25329 , \25339 );
and \U$25055 ( \25432 , \25431 , \25350 );
and \U$25056 ( \25433 , \25329 , \25339 );
or \U$25057 ( \25434 , \25432 , \25433 );
not \U$25058 ( \25435 , \2367 );
not \U$25059 ( \25436 , RIc226c50_21);
not \U$25060 ( \25437 , \1990 );
or \U$25061 ( \25438 , \25436 , \25437 );
not \U$25062 ( \25439 , \3835 );
nand \U$25063 ( \25440 , \25439 , \4475 );
nand \U$25064 ( \25441 , \25438 , \25440 );
not \U$25065 ( \25442 , \25441 );
or \U$25066 ( \25443 , \25435 , \25442 );
nand \U$25067 ( \25444 , \25335 , \2392 );
nand \U$25068 ( \25445 , \25443 , \25444 );
not \U$25069 ( \25446 , \5509 );
not \U$25070 ( \25447 , \25275 );
or \U$25071 ( \25448 , \25446 , \25447 );
not \U$25072 ( \25449 , RIc2264d0_37);
not \U$25073 ( \25450 , \2178 );
or \U$25074 ( \25451 , \25449 , \25450 );
nand \U$25075 ( \25452 , \841 , \4371 );
nand \U$25076 ( \25453 , \25451 , \25452 );
nand \U$25077 ( \25454 , \25453 , \5519 );
nand \U$25078 ( \25455 , \25448 , \25454 );
xor \U$25079 ( \25456 , \25445 , \25455 );
not \U$25080 ( \25457 , \3631 );
not \U$25081 ( \25458 , RIc2266b0_33);
not \U$25082 ( \25459 , \1372 );
or \U$25083 ( \25460 , \25458 , \25459 );
nand \U$25084 ( \25461 , \1223 , \9425 );
nand \U$25085 ( \25462 , \25460 , \25461 );
not \U$25086 ( \25463 , \25462 );
or \U$25087 ( \25464 , \25457 , \25463 );
not \U$25088 ( \25465 , \25316 );
nand \U$25089 ( \25466 , \25465 , \3629 );
nand \U$25090 ( \25467 , \25464 , \25466 );
xor \U$25091 ( \25468 , \25456 , \25467 );
xor \U$25092 ( \25469 , \25434 , \25468 );
not \U$25093 ( \25470 , \1340 );
not \U$25094 ( \25471 , RIc2271f0_9);
not \U$25095 ( \25472 , \17703 );
or \U$25096 ( \25473 , \25471 , \25472 );
nand \U$25097 ( \25474 , \3732 , \1342 );
nand \U$25098 ( \25475 , \25473 , \25474 );
not \U$25099 ( \25476 , \25475 );
or \U$25100 ( \25477 , \25470 , \25476 );
nand \U$25101 ( \25478 , \1597 , \25162 );
nand \U$25102 ( \25479 , \25477 , \25478 );
not \U$25103 ( \25480 , RIc2263e0_39);
not \U$25104 ( \25481 , \1074 );
or \U$25105 ( \25482 , \25480 , \25481 );
not \U$25106 ( \25483 , RIc2263e0_39);
nand \U$25107 ( \25484 , \1073 , \25483 );
nand \U$25108 ( \25485 , \25482 , \25484 );
not \U$25109 ( \25486 , \25485 );
not \U$25110 ( \25487 , \6307 );
or \U$25111 ( \25488 , \25486 , \25487 );
not \U$25112 ( \25489 , \25295 );
nand \U$25113 ( \25490 , \25489 , \6689 );
nand \U$25114 ( \25491 , \25488 , \25490 );
xor \U$25115 ( \25492 , \25479 , \25491 );
not \U$25116 ( \25493 , \1311 );
not \U$25117 ( \25494 , RIc227100_11);
not \U$25118 ( \25495 , \6425 );
or \U$25119 ( \25496 , \25494 , \25495 );
nand \U$25120 ( \25497 , \4501 , \3351 );
nand \U$25121 ( \25498 , \25496 , \25497 );
not \U$25122 ( \25499 , \25498 );
or \U$25123 ( \25500 , \25493 , \25499 );
nand \U$25124 ( \25501 , \25381 , \1307 );
nand \U$25125 ( \25502 , \25500 , \25501 );
xor \U$25126 ( \25503 , \25492 , \25502 );
xor \U$25127 ( \25504 , \25469 , \25503 );
xor \U$25128 ( \25505 , \24599 , \25221 );
and \U$25129 ( \25506 , \25505 , \25233 );
and \U$25130 ( \25507 , \24599 , \25221 );
or \U$25131 ( \25508 , \25506 , \25507 );
not \U$25132 ( \25509 , \25508 );
not \U$25133 ( \25510 , \2518 );
not \U$25134 ( \25511 , \25346 );
or \U$25135 ( \25512 , \25510 , \25511 );
not \U$25136 ( \25513 , RIc226d40_19);
not \U$25137 ( \25514 , \2592 );
or \U$25138 ( \25515 , \25513 , \25514 );
nand \U$25139 ( \25516 , \3183 , \2523 );
nand \U$25140 ( \25517 , \25515 , \25516 );
nand \U$25141 ( \25518 , \25517 , \2534 );
nand \U$25142 ( \25519 , \25512 , \25518 );
not \U$25143 ( \25520 , \1963 );
not \U$25144 ( \25521 , RIc226e30_17);
not \U$25145 ( \25522 , \2476 );
or \U$25146 ( \25523 , \25521 , \25522 );
nand \U$25147 ( \25524 , \20114 , \1952 );
nand \U$25148 ( \25525 , \25523 , \25524 );
not \U$25149 ( \25526 , \25525 );
or \U$25150 ( \25527 , \25520 , \25526 );
nand \U$25151 ( \25528 , \25217 , \1945 );
nand \U$25152 ( \25529 , \25527 , \25528 );
xor \U$25153 ( \25530 , \25519 , \25529 );
not \U$25154 ( \25531 , \3653 );
not \U$25155 ( \25532 , RIc2267a0_31);
not \U$25156 ( \25533 , \1531 );
or \U$25157 ( \25534 , \25532 , \25533 );
nand \U$25158 ( \25535 , \1532 , \2072 );
nand \U$25159 ( \25536 , \25534 , \25535 );
not \U$25160 ( \25537 , \25536 );
or \U$25161 ( \25538 , \25531 , \25537 );
nand \U$25162 ( \25539 , \25325 , \2697 );
nand \U$25163 ( \25540 , \25538 , \25539 );
xor \U$25164 ( \25541 , \25530 , \25540 );
xor \U$25165 ( \25542 , \25509 , \25541 );
not \U$25166 ( \25543 , RIc226a70_25);
not \U$25167 ( \25544 , \2424 );
or \U$25168 ( \25545 , \25543 , \25544 );
nand \U$25169 ( \25546 , \4457 , \1905 );
nand \U$25170 ( \25547 , \25545 , \25546 );
and \U$25171 ( \25548 , \25547 , \2173 );
and \U$25172 ( \25549 , \25285 , \2195 );
nor \U$25173 ( \25550 , \25548 , \25549 );
not \U$25174 ( \25551 , RIc2265c0_35);
not \U$25175 ( \25552 , \2120 );
or \U$25176 ( \25553 , \25551 , \25552 );
nand \U$25177 ( \25554 , \1455 , \4376 );
nand \U$25178 ( \25555 , \25553 , \25554 );
and \U$25179 ( \25556 , \25555 , \5135 );
and \U$25180 ( \25557 , \25263 , \5741 );
nor \U$25181 ( \25558 , \25556 , \25557 );
xor \U$25182 ( \25559 , \25550 , \25558 );
not \U$25183 ( \25560 , \1930 );
not \U$25184 ( \25561 , \2229 );
not \U$25185 ( \25562 , \1911 );
and \U$25186 ( \25563 , \25561 , \25562 );
and \U$25187 ( \25564 , \5697 , \1911 );
nor \U$25188 ( \25565 , \25563 , \25564 );
nor \U$25189 ( \25566 , \25560 , \25565 );
not \U$25190 ( \25567 , \25306 );
nor \U$25191 ( \25568 , \25567 , \5643 );
nor \U$25192 ( \25569 , \25566 , \25568 );
xor \U$25193 ( \25570 , \25559 , \25569 );
xor \U$25194 ( \25571 , \25542 , \25570 );
xor \U$25195 ( \25572 , \25504 , \25571 );
or \U$25196 ( \25573 , \25114 , \25105 );
nand \U$25197 ( \25574 , \25573 , \25119 );
nand \U$25198 ( \25575 , \25114 , \25105 );
nand \U$25199 ( \25576 , \25574 , \25575 );
xnor \U$25200 ( \25577 , \25572 , \25576 );
not \U$25201 ( \25578 , \25120 );
not \U$25202 ( \25579 , \25097 );
or \U$25203 ( \25580 , \25578 , \25579 );
nand \U$25204 ( \25581 , \25580 , \25040 );
nand \U$25205 ( \25582 , \25096 , \25123 );
and \U$25206 ( \25583 , \25581 , \25582 );
xor \U$25207 ( \25584 , \25577 , \25583 );
not \U$25208 ( \25585 , \25194 );
not \U$25209 ( \25586 , \25186 );
or \U$25210 ( \25587 , \25585 , \25586 );
nand \U$25211 ( \25588 , \25587 , \25181 );
nand \U$25212 ( \25589 , \25185 , \25195 );
and \U$25213 ( \25590 , \25588 , \25589 );
not \U$25214 ( \25591 , \25590 );
xor \U$25215 ( \25592 , \25047 , \25051 );
and \U$25216 ( \25593 , \25592 , \25082 );
and \U$25217 ( \25594 , \25047 , \25051 );
or \U$25218 ( \25595 , \25593 , \25594 );
not \U$25219 ( \25596 , \25595 );
and \U$25220 ( \25597 , \25591 , \25596 );
and \U$25221 ( \25598 , \25590 , \25595 );
nor \U$25222 ( \25599 , \25597 , \25598 );
xor \U$25223 ( \25600 , \25301 , \25309 );
and \U$25224 ( \25601 , \25600 , \25318 );
and \U$25225 ( \25602 , \25301 , \25309 );
or \U$25226 ( \25603 , \25601 , \25602 );
not \U$25227 ( \25604 , \25603 );
not \U$25228 ( \25605 , \25604 );
or \U$25229 ( \25606 , \25374 , \25364 );
and \U$25230 ( \25607 , \25606 , \25385 );
and \U$25231 ( \25608 , \25364 , \25374 );
nor \U$25232 ( \25609 , \25607 , \25608 );
not \U$25233 ( \25610 , \25609 );
or \U$25234 ( \25611 , \25605 , \25610 );
not \U$25235 ( \25612 , \25609 );
nand \U$25236 ( \25613 , \25612 , \25603 );
nand \U$25237 ( \25614 , \25611 , \25613 );
xor \U$25238 ( \25615 , \25267 , \25277 );
and \U$25239 ( \25616 , \25615 , \25289 );
and \U$25240 ( \25617 , \25267 , \25277 );
or \U$25241 ( \25618 , \25616 , \25617 );
xnor \U$25242 ( \25619 , \25614 , \25618 );
xor \U$25243 ( \25620 , \25599 , \25619 );
or \U$25244 ( \25621 , \25083 , \25090 );
and \U$25245 ( \25622 , \25621 , \25095 );
and \U$25246 ( \25623 , \25083 , \25090 );
nor \U$25247 ( \25624 , \25622 , \25623 );
not \U$25248 ( \25625 , \25624 );
and \U$25249 ( \25626 , \25620 , \25625 );
not \U$25250 ( \25627 , \25620 );
and \U$25251 ( \25628 , \25627 , \25624 );
nor \U$25252 ( \25629 , \25626 , \25628 );
not \U$25253 ( \25630 , \2320 );
not \U$25254 ( \25631 , \25231 );
or \U$25255 ( \25632 , \25630 , \25631 );
not \U$25256 ( \25633 , RIc226f20_15);
not \U$25257 ( \25634 , \2671 );
or \U$25258 ( \25635 , \25633 , \25634 );
nand \U$25259 ( \25636 , \2720 , \1674 );
nand \U$25260 ( \25637 , \25635 , \25636 );
nand \U$25261 ( \25638 , \25637 , \2358 );
nand \U$25262 ( \25639 , \25632 , \25638 );
not \U$25263 ( \25640 , \2078 );
not \U$25264 ( \25641 , \25241 );
or \U$25265 ( \25642 , \25640 , \25641 );
and \U$25266 ( \25643 , RIc226890_29, \1487 );
not \U$25267 ( \25644 , RIc226890_29);
and \U$25268 ( \25645 , \25644 , \1486 );
or \U$25269 ( \25646 , \25643 , \25645 );
nand \U$25270 ( \25647 , \25646 , \2086 );
nand \U$25271 ( \25648 , \25642 , \25647 );
xor \U$25272 ( \25649 , \25639 , \25648 );
not \U$25273 ( \25650 , \1682 );
not \U$25274 ( \25651 , RIc227010_13);
not \U$25275 ( \25652 , \5527 );
or \U$25276 ( \25653 , \25651 , \25652 );
nand \U$25277 ( \25654 , \3800 , \1296 );
nand \U$25278 ( \25655 , \25653 , \25654 );
not \U$25279 ( \25656 , \25655 );
or \U$25280 ( \25657 , \25650 , \25656 );
nand \U$25281 ( \25658 , \25254 , \3250 );
nand \U$25282 ( \25659 , \25657 , \25658 );
buf \U$25283 ( \25660 , \25659 );
xor \U$25284 ( \25661 , \25649 , \25660 );
not \U$25285 ( \25662 , \9817 );
not \U$25286 ( \25663 , \6303 );
and \U$25287 ( \25664 , \25662 , \25663 );
and \U$25288 ( \25665 , \25358 , \9690 );
nor \U$25289 ( \25666 , \25664 , \25665 );
xor \U$25290 ( \25667 , \25145 , \25155 );
and \U$25291 ( \25668 , \25667 , \25166 );
and \U$25292 ( \25669 , \25145 , \25155 );
or \U$25293 ( \25670 , \25668 , \25669 );
xor \U$25294 ( \25671 , \25666 , \25670 );
xor \U$25295 ( \25672 , \25061 , \25071 );
and \U$25296 ( \25673 , \25672 , \25081 );
and \U$25297 ( \25674 , \25061 , \25071 );
or \U$25298 ( \25675 , \25673 , \25674 );
xor \U$25299 ( \25676 , \25671 , \25675 );
xor \U$25300 ( \25677 , \25661 , \25676 );
xor \U$25301 ( \25678 , \25167 , \25171 );
and \U$25302 ( \25679 , \25678 , \25176 );
and \U$25303 ( \25680 , \25167 , \25171 );
or \U$25304 ( \25681 , \25679 , \25680 );
xnor \U$25305 ( \25682 , \25677 , \25681 );
and \U$25306 ( \25683 , \25629 , \25682 );
not \U$25307 ( \25684 , \25629 );
not \U$25308 ( \25685 , \25682 );
and \U$25309 ( \25686 , \25684 , \25685 );
nor \U$25310 ( \25687 , \25683 , \25686 );
xor \U$25311 ( \25688 , \25584 , \25687 );
nand \U$25312 ( \25689 , \25394 , \25138 );
not \U$25313 ( \25690 , \25689 );
not \U$25314 ( \25691 , \25410 );
or \U$25315 ( \25692 , \25690 , \25691 );
nand \U$25316 ( \25693 , \25395 , \25137 );
nand \U$25317 ( \25694 , \25692 , \25693 );
not \U$25318 ( \25695 , \25694 );
xor \U$25319 ( \25696 , \25688 , \25695 );
or \U$25320 ( \25697 , \25199 , \25177 );
and \U$25321 ( \25698 , \25697 , \25204 );
and \U$25322 ( \25699 , \25177 , \25199 );
nor \U$25323 ( \25700 , \25698 , \25699 );
and \U$25324 ( \25701 , RIc2275b0_1, \8886 );
not \U$25325 ( \25702 , \1082 );
not \U$25326 ( \25703 , RIc2274c0_3);
not \U$25327 ( \25704 , \23776 );
not \U$25328 ( \25705 , \25704 );
or \U$25329 ( \25706 , \25703 , \25705 );
not \U$25330 ( \25707 , \16555 );
nand \U$25331 ( \25708 , \25707 , \1027 );
nand \U$25332 ( \25709 , \25706 , \25708 );
not \U$25333 ( \25710 , \25709 );
or \U$25334 ( \25711 , \25702 , \25710 );
nand \U$25335 ( \25712 , \25057 , \1040 );
nand \U$25336 ( \25713 , \25711 , \25712 );
xor \U$25337 ( \25714 , \25701 , \25713 );
not \U$25338 ( \25715 , \2154 );
not \U$25339 ( \25716 , RIc226980_27);
not \U$25340 ( \25717 , \2347 );
or \U$25341 ( \25718 , \25716 , \25717 );
nand \U$25342 ( \25719 , \2354 , \2133 );
nand \U$25343 ( \25720 , \25718 , \25719 );
not \U$25344 ( \25721 , \25720 );
or \U$25345 ( \25722 , \25715 , \25721 );
nand \U$25346 ( \25723 , \25372 , \2138 );
nand \U$25347 ( \25724 , \25722 , \25723 );
xor \U$25348 ( \25725 , \25714 , \25724 );
not \U$25349 ( \25726 , \25725 );
not \U$25350 ( \25727 , \854 );
not \U$25351 ( \25728 , \25079 );
or \U$25352 ( \25729 , \25727 , \25728 );
and \U$25353 ( \25730 , RIc2275b0_1, \6719 );
not \U$25354 ( \25731 , RIc2275b0_1);
and \U$25355 ( \25732 , \25731 , \6720 );
or \U$25356 ( \25733 , \25730 , \25732 );
nand \U$25357 ( \25734 , \25733 , \1579 );
nand \U$25358 ( \25735 , \25729 , \25734 );
not \U$25359 ( \25736 , \1118 );
not \U$25360 ( \25737 , \25151 );
or \U$25361 ( \25738 , \25736 , \25737 );
not \U$25362 ( \25739 , RIc2272e0_7);
not \U$25363 ( \25740 , \4123 );
or \U$25364 ( \25741 , \25739 , \25740 );
nand \U$25365 ( \25742 , \16519 , \1139 );
nand \U$25366 ( \25743 , \25741 , \25742 );
nand \U$25367 ( \25744 , \25743 , \1121 );
nand \U$25368 ( \25745 , \25738 , \25744 );
xor \U$25369 ( \25746 , \25735 , \25745 );
not \U$25370 ( \25747 , \951 );
not \U$25371 ( \25748 , \25067 );
or \U$25372 ( \25749 , \25747 , \25748 );
not \U$25373 ( \25750 , RIc2273d0_5);
not \U$25374 ( \25751 , \5216 );
or \U$25375 ( \25752 , \25750 , \25751 );
nand \U$25376 ( \25753 , \5217 , \946 );
nand \U$25377 ( \25754 , \25752 , \25753 );
nand \U$25378 ( \25755 , \25754 , \954 );
nand \U$25379 ( \25756 , \25749 , \25755 );
xnor \U$25380 ( \25757 , \25746 , \25756 );
not \U$25381 ( \25758 , \25757 );
or \U$25382 ( \25759 , \25726 , \25758 );
or \U$25383 ( \25760 , \25725 , \25757 );
nand \U$25384 ( \25761 , \25759 , \25760 );
xor \U$25385 ( \25762 , \25236 , \25245 );
and \U$25386 ( \25763 , \25762 , \25256 );
and \U$25387 ( \25764 , \25236 , \25245 );
or \U$25388 ( \25765 , \25763 , \25764 );
and \U$25389 ( \25766 , \25761 , \25765 );
not \U$25390 ( \25767 , \25761 );
not \U$25391 ( \25768 , \25765 );
and \U$25392 ( \25769 , \25767 , \25768 );
nor \U$25393 ( \25770 , \25766 , \25769 );
not \U$25394 ( \25771 , \25386 );
not \U$25395 ( \25772 , \25351 );
or \U$25396 ( \25773 , \25771 , \25772 );
or \U$25397 ( \25774 , \25351 , \25386 );
not \U$25398 ( \25775 , \25319 );
nand \U$25399 ( \25776 , \25774 , \25775 );
nand \U$25400 ( \25777 , \25773 , \25776 );
xor \U$25401 ( \25778 , \25770 , \25777 );
xor \U$25402 ( \25779 , \25234 , \25257 );
and \U$25403 ( \25780 , \25779 , \25290 );
and \U$25404 ( \25781 , \25234 , \25257 );
or \U$25405 ( \25782 , \25780 , \25781 );
xor \U$25406 ( \25783 , \25778 , \25782 );
xor \U$25407 ( \25784 , \25700 , \25783 );
xor \U$25408 ( \25785 , \25291 , \25387 );
and \U$25409 ( \25786 , \25785 , \25392 );
and \U$25410 ( \25787 , \25291 , \25387 );
or \U$25411 ( \25788 , \25786 , \25787 );
xnor \U$25412 ( \25789 , \25784 , \25788 );
not \U$25413 ( \25790 , \25393 );
buf \U$25414 ( \25791 , \25209 );
not \U$25415 ( \25792 , \25791 );
or \U$25416 ( \25793 , \25790 , \25792 );
or \U$25417 ( \25794 , \25791 , \25393 );
nand \U$25418 ( \25795 , \25794 , \25143 );
nand \U$25419 ( \25796 , \25793 , \25795 );
and \U$25420 ( \25797 , \25789 , \25796 );
not \U$25421 ( \25798 , \25789 );
not \U$25422 ( \25799 , \25796 );
and \U$25423 ( \25800 , \25798 , \25799 );
nor \U$25424 ( \25801 , \25797 , \25800 );
not \U$25425 ( \25802 , \25126 );
not \U$25426 ( \25803 , \25022 );
or \U$25427 ( \25804 , \25802 , \25803 );
not \U$25428 ( \25805 , \25022 );
not \U$25429 ( \25806 , \25805 );
not \U$25430 ( \25807 , \25125 );
or \U$25431 ( \25808 , \25806 , \25807 );
nand \U$25432 ( \25809 , \25808 , \25029 );
nand \U$25433 ( \25810 , \25804 , \25809 );
not \U$25434 ( \25811 , \25810 );
and \U$25435 ( \25812 , \25801 , \25811 );
not \U$25436 ( \25813 , \25801 );
and \U$25437 ( \25814 , \25813 , \25810 );
nor \U$25438 ( \25815 , \25812 , \25814 );
xor \U$25439 ( \25816 , \25696 , \25815 );
xor \U$25440 ( \25817 , \25127 , \25415 );
and \U$25441 ( \25818 , \25817 , \25424 );
and \U$25442 ( \25819 , \25127 , \25415 );
or \U$25443 ( \25820 , \25818 , \25819 );
nand \U$25444 ( \25821 , \25816 , \25820 );
nand \U$25445 ( \25822 , \25430 , \25821 );
nor \U$25446 ( \25823 , \25014 , \25822 );
and \U$25447 ( \25824 , \24153 , \25823 );
xor \U$25448 ( \25825 , \25701 , \25713 );
and \U$25449 ( \25826 , \25825 , \25724 );
and \U$25450 ( \25827 , \25701 , \25713 );
or \U$25451 ( \25828 , \25826 , \25827 );
nand \U$25452 ( \25829 , \20646 , RIc2275b0_1);
and \U$25453 ( \25830 , \6730 , \1082 );
and \U$25454 ( \25831 , \25709 , \1040 );
nor \U$25455 ( \25832 , \25830 , \25831 );
xor \U$25456 ( \25833 , \25829 , \25832 );
not \U$25457 ( \25834 , \25733 );
nor \U$25458 ( \25835 , \25834 , \855 );
xnor \U$25459 ( \25836 , \6494 , RIc2275b0_1);
nor \U$25460 ( \25837 , \25836 , \899 );
nor \U$25461 ( \25838 , \25835 , \25837 );
xor \U$25462 ( \25839 , \25833 , \25838 );
and \U$25463 ( \25840 , \25828 , \25839 );
not \U$25464 ( \25841 , \25828 );
not \U$25465 ( \25842 , \25839 );
and \U$25466 ( \25843 , \25841 , \25842 );
or \U$25467 ( \25844 , \25840 , \25843 );
and \U$25468 ( \25845 , \16459 , \9817 );
nor \U$25469 ( \25846 , \25845 , \12937 );
not \U$25470 ( \25847 , \25754 );
not \U$25471 ( \25848 , \25847 );
not \U$25472 ( \25849 , \952 );
and \U$25473 ( \25850 , \25848 , \25849 );
and \U$25474 ( \25851 , \6742 , \954 );
nor \U$25475 ( \25852 , \25850 , \25851 );
xor \U$25476 ( \25853 , \25846 , \25852 );
not \U$25477 ( \25854 , \25743 );
not \U$25478 ( \25855 , \25854 );
not \U$25479 ( \25856 , \1117 );
and \U$25480 ( \25857 , \25855 , \25856 );
and \U$25481 ( \25858 , \6826 , \1121 );
nor \U$25482 ( \25859 , \25857 , \25858 );
xor \U$25483 ( \25860 , \25853 , \25859 );
and \U$25484 ( \25861 , \25844 , \25860 );
not \U$25485 ( \25862 , \25844 );
not \U$25486 ( \25863 , \25860 );
and \U$25487 ( \25864 , \25862 , \25863 );
nor \U$25488 ( \25865 , \25861 , \25864 );
not \U$25489 ( \25866 , \2697 );
not \U$25490 ( \25867 , \25536 );
or \U$25491 ( \25868 , \25866 , \25867 );
nand \U$25492 ( \25869 , \6904 , \2711 );
nand \U$25493 ( \25870 , \25868 , \25869 );
not \U$25494 ( \25871 , \5509 );
not \U$25495 ( \25872 , \25453 );
or \U$25496 ( \25873 , \25871 , \25872 );
nand \U$25497 ( \25874 , \6801 , \5519 );
nand \U$25498 ( \25875 , \25873 , \25874 );
xor \U$25499 ( \25876 , \25870 , \25875 );
not \U$25500 ( \25877 , \2518 );
not \U$25501 ( \25878 , \25517 );
or \U$25502 ( \25879 , \25877 , \25878 );
nand \U$25503 ( \25880 , \6773 , \2534 );
nand \U$25504 ( \25881 , \25879 , \25880 );
xor \U$25505 ( \25882 , \25876 , \25881 );
not \U$25506 ( \25883 , \25565 );
not \U$25507 ( \25884 , \5643 );
and \U$25508 ( \25885 , \25883 , \25884 );
and \U$25509 ( \25886 , \6813 , \1930 );
nor \U$25510 ( \25887 , \25885 , \25886 );
not \U$25511 ( \25888 , \3629 );
not \U$25512 ( \25889 , \25462 );
or \U$25513 ( \25890 , \25888 , \25889 );
nand \U$25514 ( \25891 , \6892 , \3631 );
nand \U$25515 ( \25892 , \25890 , \25891 );
xor \U$25516 ( \25893 , \25887 , \25892 );
not \U$25517 ( \25894 , \2392 );
not \U$25518 ( \25895 , \25441 );
or \U$25519 ( \25896 , \25894 , \25895 );
nand \U$25520 ( \25897 , \6881 , \2367 );
nand \U$25521 ( \25898 , \25896 , \25897 );
not \U$25522 ( \25899 , \25898 );
xor \U$25523 ( \25900 , \25893 , \25899 );
xor \U$25524 ( \25901 , \25882 , \25900 );
not \U$25525 ( \25902 , \6689 );
not \U$25526 ( \25903 , \25485 );
or \U$25527 ( \25904 , \25902 , \25903 );
nand \U$25528 ( \25905 , \6696 , \6307 );
nand \U$25529 ( \25906 , \25904 , \25905 );
not \U$25530 ( \25907 , \5741 );
not \U$25531 ( \25908 , \25555 );
or \U$25532 ( \25909 , \25907 , \25908 );
nand \U$25533 ( \25910 , \6786 , \5135 );
nand \U$25534 ( \25911 , \25909 , \25910 );
xor \U$25535 ( \25912 , \25906 , \25911 );
not \U$25536 ( \25913 , \2195 );
not \U$25537 ( \25914 , \25547 );
or \U$25538 ( \25915 , \25913 , \25914 );
and \U$25539 ( \25916 , \2306 , \1905 );
not \U$25540 ( \25917 , \2306 );
and \U$25541 ( \25918 , \25917 , RIc226a70_25);
or \U$25542 ( \25919 , \25916 , \25918 );
nand \U$25543 ( \25920 , \25919 , \2173 );
nand \U$25544 ( \25921 , \25915 , \25920 );
xor \U$25545 ( \25922 , \25912 , \25921 );
not \U$25546 ( \25923 , \25922 );
and \U$25547 ( \25924 , \25901 , \25923 );
not \U$25548 ( \25925 , \25901 );
and \U$25549 ( \25926 , \25925 , \25922 );
nor \U$25550 ( \25927 , \25924 , \25926 );
xor \U$25551 ( \25928 , \25865 , \25927 );
or \U$25552 ( \25929 , \25676 , \25661 );
nand \U$25553 ( \25930 , \25929 , \25681 );
nand \U$25554 ( \25931 , \25676 , \25661 );
and \U$25555 ( \25932 , \25930 , \25931 );
and \U$25556 ( \25933 , \25928 , \25932 );
and \U$25557 ( \25934 , \25865 , \25927 );
or \U$25558 ( \25935 , \25933 , \25934 );
xor \U$25559 ( \25936 , \6764 , \6775 );
xnor \U$25560 ( \25937 , \25936 , \6788 );
xor \U$25561 ( \25938 , \6883 , \6894 );
xor \U$25562 ( \25939 , \25938 , \6906 );
xor \U$25563 ( \25940 , \25937 , \25939 );
and \U$25564 ( \25941 , \1340 , \6429 );
not \U$25565 ( \25942 , RIc2271f0_9);
not \U$25566 ( \25943 , \3116 );
or \U$25567 ( \25944 , \25942 , \25943 );
nand \U$25568 ( \25945 , \3120 , \1351 );
nand \U$25569 ( \25946 , \25944 , \25945 );
and \U$25570 ( \25947 , \25946 , \1363 );
nor \U$25571 ( \25948 , \25941 , \25947 );
not \U$25572 ( \25949 , \1579 );
not \U$25573 ( \25950 , \6496 );
or \U$25574 ( \25951 , \25949 , \25950 );
not \U$25575 ( \25952 , \25836 );
nand \U$25576 ( \25953 , \25952 , \854 );
nand \U$25577 ( \25954 , \25951 , \25953 );
not \U$25578 ( \25955 , \25919 );
not \U$25579 ( \25956 , \2195 );
or \U$25580 ( \25957 , \25955 , \25956 );
not \U$25581 ( \25958 , \6508 );
nand \U$25582 ( \25959 , \25958 , \2173 );
nand \U$25583 ( \25960 , \25957 , \25959 );
xor \U$25584 ( \25961 , \25954 , \25960 );
xnor \U$25585 ( \25962 , \25948 , \25961 );
xor \U$25586 ( \25963 , \25940 , \25962 );
nand \U$25587 ( \25964 , \25768 , \25757 );
and \U$25588 ( \25965 , \25964 , \25725 );
nor \U$25589 ( \25966 , \25768 , \25757 );
nor \U$25590 ( \25967 , \25965 , \25966 );
not \U$25591 ( \25968 , \25603 );
not \U$25592 ( \25969 , \25609 );
or \U$25593 ( \25970 , \25968 , \25969 );
nand \U$25594 ( \25971 , \25970 , \25618 );
nand \U$25595 ( \25972 , \25612 , \25604 );
and \U$25596 ( \25973 , \25971 , \25972 );
xor \U$25597 ( \25974 , \25967 , \25973 );
nand \U$25598 ( \25975 , \25570 , \25509 );
and \U$25599 ( \25976 , \25975 , \25541 );
nor \U$25600 ( \25977 , \25570 , \25509 );
nor \U$25601 ( \25978 , \25976 , \25977 );
and \U$25602 ( \25979 , \25974 , \25978 );
and \U$25603 ( \25980 , \25967 , \25973 );
or \U$25604 ( \25981 , \25979 , \25980 );
xor \U$25605 ( \25982 , \25963 , \25981 );
not \U$25606 ( \25983 , \25860 );
not \U$25607 ( \25984 , \25839 );
or \U$25608 ( \25985 , \25983 , \25984 );
nand \U$25609 ( \25986 , \25985 , \25828 );
nand \U$25610 ( \25987 , \25842 , \25863 );
and \U$25611 ( \25988 , \25986 , \25987 );
xor \U$25612 ( \25989 , \25829 , \25832 );
and \U$25613 ( \25990 , \25989 , \25838 );
and \U$25614 ( \25991 , \25829 , \25832 );
or \U$25615 ( \25992 , \25990 , \25991 );
xor \U$25616 ( \25993 , \25846 , \25852 );
and \U$25617 ( \25994 , \25993 , \25859 );
and \U$25618 ( \25995 , \25846 , \25852 );
or \U$25619 ( \25996 , \25994 , \25995 );
xor \U$25620 ( \25997 , \25992 , \25996 );
xor \U$25621 ( \25998 , \6721 , \6732 );
xnor \U$25622 ( \25999 , \25998 , \6746 );
xor \U$25623 ( \26000 , \25997 , \25999 );
not \U$25624 ( \26001 , \26000 );
xor \U$25625 ( \26002 , \25988 , \26001 );
not \U$25626 ( \26003 , \25455 );
not \U$25627 ( \26004 , \25445 );
or \U$25628 ( \26005 , \26003 , \26004 );
or \U$25629 ( \26006 , \25445 , \25455 );
nand \U$25630 ( \26007 , \26006 , \25467 );
nand \U$25631 ( \26008 , \26005 , \26007 );
not \U$25632 ( \26009 , \26008 );
xor \U$25633 ( \26010 , \25550 , \25558 );
and \U$25634 ( \26011 , \26010 , \25569 );
and \U$25635 ( \26012 , \25550 , \25558 );
or \U$25636 ( \26013 , \26011 , \26012 );
not \U$25637 ( \26014 , \26013 );
not \U$25638 ( \26015 , \26014 );
or \U$25639 ( \26016 , \26009 , \26015 );
not \U$25640 ( \26017 , \26008 );
not \U$25641 ( \26018 , \26017 );
not \U$25642 ( \26019 , \26013 );
or \U$25643 ( \26020 , \26018 , \26019 );
not \U$25644 ( \26021 , \25491 );
not \U$25645 ( \26022 , \25479 );
or \U$25646 ( \26023 , \26021 , \26022 );
or \U$25647 ( \26024 , \25479 , \25491 );
nand \U$25648 ( \26025 , \26024 , \25502 );
nand \U$25649 ( \26026 , \26023 , \26025 );
nand \U$25650 ( \26027 , \26020 , \26026 );
nand \U$25651 ( \26028 , \26016 , \26027 );
xor \U$25652 ( \26029 , \26002 , \26028 );
xor \U$25653 ( \26030 , \25982 , \26029 );
xor \U$25654 ( \26031 , \25935 , \26030 );
not \U$25655 ( \26032 , \1963 );
not \U$25656 ( \26033 , \6838 );
or \U$25657 ( \26034 , \26032 , \26033 );
not \U$25658 ( \26035 , \7140 );
nand \U$25659 ( \26036 , \26035 , \25525 );
nand \U$25660 ( \26037 , \26034 , \26036 );
not \U$25661 ( \26038 , \2358 );
not \U$25662 ( \26039 , \6864 );
or \U$25663 ( \26040 , \26038 , \26039 );
nand \U$25664 ( \26041 , \25637 , \2320 );
nand \U$25665 ( \26042 , \26040 , \26041 );
xor \U$25666 ( \26043 , \26037 , \26042 );
not \U$25667 ( \26044 , \2078 );
not \U$25668 ( \26045 , \25646 );
or \U$25669 ( \26046 , \26044 , \26045 );
nand \U$25670 ( \26047 , \6762 , \2086 );
nand \U$25671 ( \26048 , \26046 , \26047 );
xnor \U$25672 ( \26049 , \26043 , \26048 );
not \U$25673 ( \26050 , \1682 );
not \U$25674 ( \26051 , RIc227010_13);
not \U$25675 ( \26052 , \3011 );
or \U$25676 ( \26053 , \26051 , \26052 );
nand \U$25677 ( \26054 , \4240 , \2427 );
nand \U$25678 ( \26055 , \26053 , \26054 );
not \U$25679 ( \26056 , \26055 );
or \U$25680 ( \26057 , \26050 , \26056 );
nand \U$25681 ( \26058 , \25655 , \1680 );
nand \U$25682 ( \26059 , \26057 , \26058 );
not \U$25683 ( \26060 , \26059 );
xor \U$25684 ( \26061 , \25666 , \26060 );
not \U$25685 ( \26062 , \25735 );
not \U$25686 ( \26063 , \25756 );
or \U$25687 ( \26064 , \26062 , \26063 );
or \U$25688 ( \26065 , \25756 , \25735 );
nand \U$25689 ( \26066 , \26065 , \25745 );
nand \U$25690 ( \26067 , \26064 , \26066 );
xnor \U$25691 ( \26068 , \26061 , \26067 );
xor \U$25692 ( \26069 , \26049 , \26068 );
xor \U$25693 ( \26070 , \25666 , \25670 );
and \U$25694 ( \26071 , \26070 , \25675 );
and \U$25695 ( \26072 , \25666 , \25670 );
or \U$25696 ( \26073 , \26071 , \26072 );
xnor \U$25697 ( \26074 , \26069 , \26073 );
xor \U$25698 ( \26075 , \25967 , \25973 );
xor \U$25699 ( \26076 , \26075 , \25978 );
xor \U$25700 ( \26077 , \26074 , \26076 );
nand \U$25701 ( \26078 , \25619 , \25590 );
and \U$25702 ( \26079 , \26078 , \25595 );
nor \U$25703 ( \26080 , \25619 , \25590 );
nor \U$25704 ( \26081 , \26079 , \26080 );
and \U$25705 ( \26082 , \26077 , \26081 );
and \U$25706 ( \26083 , \26074 , \26076 );
or \U$25707 ( \26084 , \26082 , \26083 );
xor \U$25708 ( \26085 , \26031 , \26084 );
not \U$25709 ( \26086 , \25783 );
buf \U$25710 ( \26087 , \25700 );
nand \U$25711 ( \26088 , \26086 , \26087 );
and \U$25712 ( \26089 , \26088 , \25788 );
nor \U$25713 ( \26090 , \26086 , \26087 );
nor \U$25714 ( \26091 , \26089 , \26090 );
or \U$25715 ( \26092 , \25782 , \25770 );
nand \U$25716 ( \26093 , \26092 , \25777 );
nand \U$25717 ( \26094 , \25782 , \25770 );
and \U$25718 ( \26095 , \26093 , \26094 );
not \U$25719 ( \26096 , \25540 );
not \U$25720 ( \26097 , \25529 );
or \U$25721 ( \26098 , \26096 , \26097 );
or \U$25722 ( \26099 , \25540 , \25529 );
nand \U$25723 ( \26100 , \26099 , \25519 );
nand \U$25724 ( \26101 , \26098 , \26100 );
not \U$25725 ( \26102 , \25648 );
not \U$25726 ( \26103 , \25639 );
or \U$25727 ( \26104 , \26102 , \26103 );
or \U$25728 ( \26105 , \25639 , \25648 );
nand \U$25729 ( \26106 , \26105 , \25659 );
nand \U$25730 ( \26107 , \26104 , \26106 );
not \U$25731 ( \26108 , \26107 );
xor \U$25732 ( \26109 , \26101 , \26108 );
not \U$25733 ( \26110 , \1340 );
not \U$25734 ( \26111 , \25946 );
or \U$25735 ( \26112 , \26110 , \26111 );
nand \U$25736 ( \26113 , \25475 , \1363 );
nand \U$25737 ( \26114 , \26112 , \26113 );
not \U$25738 ( \26115 , \6850 );
not \U$25739 ( \26116 , \2155 );
and \U$25740 ( \26117 , \26115 , \26116 );
and \U$25741 ( \26118 , \25720 , \2138 );
nor \U$25742 ( \26119 , \26117 , \26118 );
xor \U$25743 ( \26120 , \26114 , \26119 );
not \U$25744 ( \26121 , \1307 );
not \U$25745 ( \26122 , \25498 );
or \U$25746 ( \26123 , \26121 , \26122 );
not \U$25747 ( \26124 , RIc227100_11);
not \U$25748 ( \26125 , \3564 );
or \U$25749 ( \26126 , \26124 , \26125 );
nand \U$25750 ( \26127 , \2636 , \1685 );
nand \U$25751 ( \26128 , \26126 , \26127 );
nand \U$25752 ( \26129 , \26128 , \1311 );
nand \U$25753 ( \26130 , \26123 , \26129 );
xor \U$25754 ( \26131 , \26120 , \26130 );
xnor \U$25755 ( \26132 , \26109 , \26131 );
not \U$25756 ( \26133 , \26026 );
not \U$25757 ( \26134 , \26017 );
or \U$25758 ( \26135 , \26133 , \26134 );
or \U$25759 ( \26136 , \26017 , \26026 );
nand \U$25760 ( \26137 , \26135 , \26136 );
and \U$25761 ( \26138 , \26137 , \26013 );
not \U$25762 ( \26139 , \26137 );
and \U$25763 ( \26140 , \26139 , \26014 );
nor \U$25764 ( \26141 , \26138 , \26140 );
xor \U$25765 ( \26142 , \26132 , \26141 );
xor \U$25766 ( \26143 , \25434 , \25468 );
and \U$25767 ( \26144 , \26143 , \25503 );
and \U$25768 ( \26145 , \25434 , \25468 );
or \U$25769 ( \26146 , \26144 , \26145 );
xnor \U$25770 ( \26147 , \26142 , \26146 );
xor \U$25771 ( \26148 , \26095 , \26147 );
xor \U$25772 ( \26149 , \25865 , \25927 );
xor \U$25773 ( \26150 , \26149 , \25932 );
xor \U$25774 ( \26151 , \26148 , \26150 );
xor \U$25775 ( \26152 , \26091 , \26151 );
or \U$25776 ( \26153 , \25571 , \25504 );
and \U$25777 ( \26154 , \26153 , \25576 );
and \U$25778 ( \26155 , \25504 , \25571 );
nor \U$25779 ( \26156 , \26154 , \26155 );
not \U$25780 ( \26157 , \25682 );
not \U$25781 ( \26158 , \25624 );
or \U$25782 ( \26159 , \26157 , \26158 );
nand \U$25783 ( \26160 , \26159 , \25620 );
nand \U$25784 ( \26161 , \25625 , \25685 );
and \U$25785 ( \26162 , \26160 , \26161 );
xor \U$25786 ( \26163 , \26156 , \26162 );
xor \U$25787 ( \26164 , \26074 , \26076 );
xor \U$25788 ( \26165 , \26164 , \26081 );
xor \U$25789 ( \26166 , \26163 , \26165 );
and \U$25790 ( \26167 , \26152 , \26166 );
and \U$25791 ( \26168 , \26091 , \26151 );
or \U$25792 ( \26169 , \26167 , \26168 );
xor \U$25793 ( \26170 , \26085 , \26169 );
nand \U$25794 ( \26171 , \26132 , \26141 );
and \U$25795 ( \26172 , \26171 , \26146 );
nor \U$25796 ( \26173 , \26141 , \26132 );
nor \U$25797 ( \26174 , \26172 , \26173 );
nand \U$25798 ( \26175 , \26131 , \26108 );
and \U$25799 ( \26176 , \26175 , \26101 );
nor \U$25800 ( \26177 , \26131 , \26108 );
nor \U$25801 ( \26178 , \26176 , \26177 );
not \U$25802 ( \26179 , \26048 );
not \U$25803 ( \26180 , \26042 );
or \U$25804 ( \26181 , \26179 , \26180 );
or \U$25805 ( \26182 , \26042 , \26048 );
nand \U$25806 ( \26183 , \26182 , \26037 );
nand \U$25807 ( \26184 , \26181 , \26183 );
xor \U$25808 ( \26185 , \25870 , \25875 );
and \U$25809 ( \26186 , \26185 , \25881 );
and \U$25810 ( \26187 , \25870 , \25875 );
or \U$25811 ( \26188 , \26186 , \26187 );
xor \U$25812 ( \26189 , \26184 , \26188 );
not \U$25813 ( \26190 , \1311 );
not \U$25814 ( \26191 , \6570 );
or \U$25815 ( \26192 , \26190 , \26191 );
nand \U$25816 ( \26193 , \26128 , \1307 );
nand \U$25817 ( \26194 , \26192 , \26193 );
xor \U$25818 ( \26195 , \6700 , \26194 );
not \U$25819 ( \26196 , \3250 );
not \U$25820 ( \26197 , \26055 );
or \U$25821 ( \26198 , \26196 , \26197 );
nand \U$25822 ( \26199 , \6591 , \1682 );
nand \U$25823 ( \26200 , \26198 , \26199 );
xnor \U$25824 ( \26201 , \26195 , \26200 );
xnor \U$25825 ( \26202 , \26189 , \26201 );
xor \U$25826 ( \26203 , \26178 , \26202 );
or \U$25827 ( \26204 , \25900 , \25882 );
and \U$25828 ( \26205 , \26204 , \25922 );
and \U$25829 ( \26206 , \25882 , \25900 );
nor \U$25830 ( \26207 , \26205 , \26206 );
xor \U$25831 ( \26208 , \26203 , \26207 );
xor \U$25832 ( \26209 , \26174 , \26208 );
nand \U$25833 ( \26210 , \26068 , \26049 );
and \U$25834 ( \26211 , \26210 , \26073 );
nor \U$25835 ( \26212 , \26068 , \26049 );
nor \U$25836 ( \26213 , \26211 , \26212 );
not \U$25837 ( \26214 , \6803 );
not \U$25838 ( \26215 , \6816 );
or \U$25839 ( \26216 , \26214 , \26215 );
nand \U$25840 ( \26217 , \6815 , \6804 );
nand \U$25841 ( \26218 , \26216 , \26217 );
not \U$25842 ( \26219 , \6828 );
and \U$25843 ( \26220 , \26218 , \26219 );
not \U$25844 ( \26221 , \26218 );
and \U$25845 ( \26222 , \26221 , \6828 );
nor \U$25846 ( \26223 , \26220 , \26222 );
not \U$25847 ( \26224 , \26060 );
not \U$25848 ( \26225 , \25666 );
or \U$25849 ( \26226 , \26224 , \26225 );
nand \U$25850 ( \26227 , \26226 , \26067 );
not \U$25851 ( \26228 , \25666 );
nand \U$25852 ( \26229 , \26228 , \26059 );
and \U$25853 ( \26230 , \26227 , \26229 );
xor \U$25854 ( \26231 , \26223 , \26230 );
xor \U$25855 ( \26232 , \6842 , \6854 );
xor \U$25856 ( \26233 , \26232 , \6866 );
xor \U$25857 ( \26234 , \26231 , \26233 );
xor \U$25858 ( \26235 , \26213 , \26234 );
not \U$25859 ( \26236 , \25899 );
not \U$25860 ( \26237 , \25887 );
or \U$25861 ( \26238 , \26236 , \26237 );
nand \U$25862 ( \26239 , \26238 , \25892 );
not \U$25863 ( \26240 , \25887 );
nand \U$25864 ( \26241 , \26240 , \25898 );
nand \U$25865 ( \26242 , \26239 , \26241 );
not \U$25866 ( \26243 , \26242 );
or \U$25867 ( \26244 , \25911 , \25921 );
nand \U$25868 ( \26245 , \26244 , \25906 );
nand \U$25869 ( \26246 , \25921 , \25911 );
and \U$25870 ( \26247 , \26245 , \26246 );
not \U$25871 ( \26248 , \26247 );
or \U$25872 ( \26249 , \26243 , \26248 );
or \U$25873 ( \26250 , \26247 , \26242 );
nand \U$25874 ( \26251 , \26249 , \26250 );
not \U$25875 ( \26252 , \26119 );
not \U$25876 ( \26253 , \26252 );
not \U$25877 ( \26254 , \26114 );
or \U$25878 ( \26255 , \26253 , \26254 );
or \U$25879 ( \26256 , \26114 , \26252 );
nand \U$25880 ( \26257 , \26256 , \26130 );
nand \U$25881 ( \26258 , \26255 , \26257 );
not \U$25882 ( \26259 , \26258 );
and \U$25883 ( \26260 , \26251 , \26259 );
not \U$25884 ( \26261 , \26251 );
and \U$25885 ( \26262 , \26261 , \26258 );
nor \U$25886 ( \26263 , \26260 , \26262 );
xor \U$25887 ( \26264 , \26235 , \26263 );
xor \U$25888 ( \26265 , \26209 , \26264 );
xor \U$25889 ( \26266 , \26095 , \26147 );
and \U$25890 ( \26267 , \26266 , \26150 );
and \U$25891 ( \26268 , \26095 , \26147 );
or \U$25892 ( \26269 , \26267 , \26268 );
xor \U$25893 ( \26270 , \26265 , \26269 );
xor \U$25894 ( \26271 , \26156 , \26162 );
and \U$25895 ( \26272 , \26271 , \26165 );
and \U$25896 ( \26273 , \26156 , \26162 );
or \U$25897 ( \26274 , \26272 , \26273 );
xor \U$25898 ( \26275 , \26270 , \26274 );
xor \U$25899 ( \26276 , \26170 , \26275 );
xor \U$25900 ( \26277 , \25577 , \25583 );
and \U$25901 ( \26278 , \26277 , \25687 );
and \U$25902 ( \26279 , \25577 , \25583 );
or \U$25903 ( \26280 , \26278 , \26279 );
not \U$25904 ( \26281 , \25810 );
not \U$25905 ( \26282 , \25789 );
nand \U$25906 ( \26283 , \26282 , \25799 );
not \U$25907 ( \26284 , \26283 );
or \U$25908 ( \26285 , \26281 , \26284 );
not \U$25909 ( \26286 , \26282 );
nand \U$25910 ( \26287 , \26286 , \25796 );
nand \U$25911 ( \26288 , \26285 , \26287 );
not \U$25912 ( \26289 , \26288 );
xor \U$25913 ( \26290 , \26280 , \26289 );
xor \U$25914 ( \26291 , \26091 , \26151 );
xor \U$25915 ( \26292 , \26291 , \26166 );
and \U$25916 ( \26293 , \26290 , \26292 );
and \U$25917 ( \26294 , \26280 , \26289 );
or \U$25918 ( \26295 , \26293 , \26294 );
nand \U$25919 ( \26296 , \26276 , \26295 );
xor \U$25920 ( \26297 , \26280 , \26289 );
xor \U$25921 ( \26298 , \26297 , \26292 );
xor \U$25922 ( \26299 , \25688 , \25695 );
and \U$25923 ( \26300 , \26299 , \25815 );
and \U$25924 ( \26301 , \25688 , \25695 );
or \U$25925 ( \26302 , \26300 , \26301 );
nand \U$25926 ( \26303 , \26298 , \26302 );
and \U$25927 ( \26304 , \26296 , \26303 );
xor \U$25928 ( \26305 , \25935 , \26030 );
and \U$25929 ( \26306 , \26305 , \26084 );
and \U$25930 ( \26307 , \25935 , \26030 );
or \U$25931 ( \26308 , \26306 , \26307 );
xor \U$25932 ( \26309 , \26178 , \26202 );
and \U$25933 ( \26310 , \26309 , \26207 );
and \U$25934 ( \26311 , \26178 , \26202 );
or \U$25935 ( \26312 , \26310 , \26311 );
xor \U$25936 ( \26313 , \6316 , \6299 );
xnor \U$25937 ( \26314 , \26313 , \6289 );
xor \U$25938 ( \26315 , \6495 , \6502 );
xor \U$25939 ( \26316 , \26315 , \6514 );
xor \U$25940 ( \26317 , \26314 , \26316 );
not \U$25941 ( \26318 , \25960 );
nand \U$25942 ( \26319 , \26318 , \25948 );
and \U$25943 ( \26320 , \26319 , \25954 );
nor \U$25944 ( \26321 , \26318 , \25948 );
nor \U$25945 ( \26322 , \26320 , \26321 );
xor \U$25946 ( \26323 , \26317 , \26322 );
or \U$25947 ( \26324 , \26184 , \26201 );
nand \U$25948 ( \26325 , \26324 , \26188 );
nand \U$25949 ( \26326 , \26201 , \26184 );
and \U$25950 ( \26327 , \26325 , \26326 );
xor \U$25951 ( \26328 , \26323 , \26327 );
xor \U$25952 ( \26329 , \6831 , \6870 );
xnor \U$25953 ( \26330 , \26329 , \6909 );
xor \U$25954 ( \26331 , \26328 , \26330 );
xor \U$25955 ( \26332 , \26312 , \26331 );
xor \U$25956 ( \26333 , \26213 , \26234 );
and \U$25957 ( \26334 , \26333 , \26263 );
and \U$25958 ( \26335 , \26213 , \26234 );
or \U$25959 ( \26336 , \26334 , \26335 );
xor \U$25960 ( \26337 , \26332 , \26336 );
xor \U$25961 ( \26338 , \26174 , \26208 );
and \U$25962 ( \26339 , \26338 , \26264 );
and \U$25963 ( \26340 , \26174 , \26208 );
or \U$25964 ( \26341 , \26339 , \26340 );
xor \U$25965 ( \26342 , \26337 , \26341 );
not \U$25966 ( \26343 , \25939 );
nand \U$25967 ( \26344 , \26343 , \25937 );
and \U$25968 ( \26345 , \26344 , \25962 );
nor \U$25969 ( \26346 , \26343 , \25937 );
nor \U$25970 ( \26347 , \26345 , \26346 );
xor \U$25971 ( \26348 , \26223 , \26230 );
and \U$25972 ( \26349 , \26348 , \26233 );
and \U$25973 ( \26350 , \26223 , \26230 );
or \U$25974 ( \26351 , \26349 , \26350 );
xor \U$25975 ( \26352 , \26347 , \26351 );
not \U$25976 ( \26353 , \26194 );
not \U$25977 ( \26354 , \26200 );
nand \U$25978 ( \26355 , \26353 , \26354 );
and \U$25979 ( \26356 , \26355 , \6751 );
not \U$25980 ( \26357 , \26194 );
nor \U$25981 ( \26358 , \26357 , \26354 );
nor \U$25982 ( \26359 , \26356 , \26358 );
xor \U$25983 ( \26360 , \6538 , \6547 );
xor \U$25984 ( \26361 , \26360 , \6527 );
xor \U$25985 ( \26362 , \26359 , \26361 );
xor \U$25986 ( \26363 , \6419 , \6445 );
xnor \U$25987 ( \26364 , \26363 , \6431 );
xor \U$25988 ( \26365 , \26362 , \26364 );
xor \U$25989 ( \26366 , \26352 , \26365 );
not \U$25990 ( \26367 , \6361 );
not \U$25991 ( \26368 , \6348 );
or \U$25992 ( \26369 , \26367 , \26368 );
or \U$25993 ( \26370 , \6348 , \6361 );
nand \U$25994 ( \26371 , \26369 , \26370 );
and \U$25995 ( \26372 , \26371 , \6336 );
not \U$25996 ( \26373 , \26371 );
and \U$25997 ( \26374 , \26373 , \6335 );
nor \U$25998 ( \26375 , \26372 , \26374 );
xor \U$25999 ( \26376 , \6404 , \6391 );
xnor \U$26000 ( \26377 , \26376 , \6389 );
xor \U$26001 ( \26378 , \26375 , \26377 );
xor \U$26002 ( \26379 , \6572 , \6582 );
xnor \U$26003 ( \26380 , \26379 , \6593 );
xor \U$26004 ( \26381 , \26378 , \26380 );
nand \U$26005 ( \26382 , \26000 , \25988 );
and \U$26006 ( \26383 , \26028 , \26382 );
not \U$26007 ( \26384 , \26001 );
nor \U$26008 ( \26385 , \26384 , \25988 );
nor \U$26009 ( \26386 , \26383 , \26385 );
xor \U$26010 ( \26387 , \26381 , \26386 );
xor \U$26011 ( \26388 , \25992 , \25996 );
and \U$26012 ( \26389 , \26388 , \25999 );
and \U$26013 ( \26390 , \25992 , \25996 );
or \U$26014 ( \26391 , \26389 , \26390 );
xor \U$26015 ( \26392 , \6748 , \6751 );
xor \U$26016 ( \26393 , \26392 , \6790 );
xor \U$26017 ( \26394 , \26391 , \26393 );
or \U$26018 ( \26395 , \26258 , \26242 );
not \U$26019 ( \26396 , \26247 );
nand \U$26020 ( \26397 , \26395 , \26396 );
nand \U$26021 ( \26398 , \26242 , \26258 );
and \U$26022 ( \26399 , \26397 , \26398 );
xor \U$26023 ( \26400 , \26394 , \26399 );
xor \U$26024 ( \26401 , \26387 , \26400 );
xor \U$26025 ( \26402 , \26366 , \26401 );
xor \U$26026 ( \26403 , \25963 , \25981 );
and \U$26027 ( \26404 , \26403 , \26029 );
and \U$26028 ( \26405 , \25963 , \25981 );
or \U$26029 ( \26406 , \26404 , \26405 );
xor \U$26030 ( \26407 , \26402 , \26406 );
xor \U$26031 ( \26408 , \26342 , \26407 );
xor \U$26032 ( \26409 , \26308 , \26408 );
xor \U$26033 ( \26410 , \26265 , \26269 );
and \U$26034 ( \26411 , \26410 , \26274 );
and \U$26035 ( \26412 , \26265 , \26269 );
or \U$26036 ( \26413 , \26411 , \26412 );
xor \U$26037 ( \26414 , \26409 , \26413 );
xor \U$26038 ( \26415 , \26085 , \26169 );
and \U$26039 ( \26416 , \26415 , \26275 );
and \U$26040 ( \26417 , \26085 , \26169 );
or \U$26041 ( \26418 , \26416 , \26417 );
nand \U$26042 ( \26419 , \26414 , \26418 );
xor \U$26043 ( \26420 , \26308 , \26408 );
and \U$26044 ( \26421 , \26420 , \26413 );
and \U$26045 ( \26422 , \26308 , \26408 );
or \U$26046 ( \26423 , \26421 , \26422 );
xor \U$26047 ( \26424 , \26314 , \26316 );
and \U$26048 ( \26425 , \26424 , \26322 );
and \U$26049 ( \26426 , \26314 , \26316 );
or \U$26050 ( \26427 , \26425 , \26426 );
xor \U$26051 ( \26428 , \26359 , \26361 );
and \U$26052 ( \26429 , \26428 , \26364 );
and \U$26053 ( \26430 , \26359 , \26361 );
or \U$26054 ( \26431 , \26429 , \26430 );
xor \U$26055 ( \26432 , \26427 , \26431 );
xor \U$26056 ( \26433 , \26375 , \26377 );
and \U$26057 ( \26434 , \26433 , \26380 );
and \U$26058 ( \26435 , \26375 , \26377 );
or \U$26059 ( \26436 , \26434 , \26435 );
xor \U$26060 ( \26437 , \26432 , \26436 );
xor \U$26061 ( \26438 , \26381 , \26386 );
and \U$26062 ( \26439 , \26438 , \26400 );
and \U$26063 ( \26440 , \26381 , \26386 );
or \U$26064 ( \26441 , \26439 , \26440 );
xor \U$26065 ( \26442 , \26437 , \26441 );
xor \U$26066 ( \26443 , \6596 , \6602 );
xor \U$26067 ( \26444 , \26443 , \6606 );
xor \U$26068 ( \26445 , \6687 , \6792 );
xnor \U$26069 ( \26446 , \26445 , \6911 );
xor \U$26070 ( \26447 , \26444 , \26446 );
xor \U$26071 ( \26448 , \26391 , \26393 );
and \U$26072 ( \26449 , \26448 , \26399 );
and \U$26073 ( \26450 , \26391 , \26393 );
or \U$26074 ( \26451 , \26449 , \26450 );
xor \U$26075 ( \26452 , \26447 , \26451 );
xor \U$26076 ( \26453 , \26442 , \26452 );
xor \U$26077 ( \26454 , \26312 , \26331 );
and \U$26078 ( \26455 , \26454 , \26336 );
and \U$26079 ( \26456 , \26312 , \26331 );
or \U$26080 ( \26457 , \26455 , \26456 );
xor \U$26081 ( \26458 , \26347 , \26351 );
and \U$26082 ( \26459 , \26458 , \26365 );
and \U$26083 ( \26460 , \26347 , \26351 );
or \U$26084 ( \26461 , \26459 , \26460 );
xor \U$26085 ( \26462 , \26323 , \26327 );
and \U$26086 ( \26463 , \26462 , \26330 );
and \U$26087 ( \26464 , \26323 , \26327 );
or \U$26088 ( \26465 , \26463 , \26464 );
xor \U$26089 ( \26466 , \26461 , \26465 );
not \U$26090 ( \26467 , \6556 );
not \U$26091 ( \26468 , \6517 );
or \U$26092 ( \26469 , \26467 , \26468 );
nand \U$26093 ( \26470 , \6559 , \6555 );
nand \U$26094 ( \26471 , \26469 , \26470 );
and \U$26095 ( \26472 , \26471 , \6551 );
not \U$26096 ( \26473 , \26471 );
and \U$26097 ( \26474 , \26473 , \6558 );
nor \U$26098 ( \26475 , \26472 , \26474 );
xor \U$26099 ( \26476 , \6447 , \6406 );
xnor \U$26100 ( \26477 , \26476 , \6364 );
xor \U$26101 ( \26478 , \26475 , \26477 );
xor \U$26102 ( \26479 , \6469 , \6467 );
xnor \U$26103 ( \26480 , \26479 , \6472 );
xor \U$26104 ( \26481 , \26478 , \26480 );
xor \U$26105 ( \26482 , \26466 , \26481 );
xor \U$26106 ( \26483 , \26457 , \26482 );
xor \U$26107 ( \26484 , \26366 , \26401 );
and \U$26108 ( \26485 , \26484 , \26406 );
and \U$26109 ( \26486 , \26366 , \26401 );
or \U$26110 ( \26487 , \26485 , \26486 );
xor \U$26111 ( \26488 , \26483 , \26487 );
xor \U$26112 ( \26489 , \26453 , \26488 );
xor \U$26113 ( \26490 , \26337 , \26341 );
and \U$26114 ( \26491 , \26490 , \26407 );
and \U$26115 ( \26492 , \26337 , \26341 );
or \U$26116 ( \26493 , \26491 , \26492 );
xor \U$26117 ( \26494 , \26489 , \26493 );
nand \U$26118 ( \26495 , \26423 , \26494 );
and \U$26119 ( \26496 , \26304 , \26419 , \26495 );
xor \U$26120 ( \26497 , \6648 , \6645 );
and \U$26121 ( \26498 , \26497 , \6641 );
not \U$26122 ( \26499 , \26497 );
and \U$26123 ( \26500 , \26499 , \6647 );
nor \U$26124 ( \26501 , \26498 , \26500 );
xor \U$26125 ( \26502 , \6682 , \6679 );
xnor \U$26126 ( \26503 , \26502 , \6914 );
xor \U$26127 ( \26504 , \26501 , \26503 );
xor \U$26128 ( \26505 , \26444 , \26446 );
and \U$26129 ( \26506 , \26505 , \26451 );
and \U$26130 ( \26507 , \26444 , \26446 );
or \U$26131 ( \26508 , \26506 , \26507 );
xor \U$26132 ( \26509 , \26504 , \26508 );
xor \U$26133 ( \26510 , \26461 , \26465 );
and \U$26134 ( \26511 , \26510 , \26481 );
and \U$26135 ( \26512 , \26461 , \26465 );
or \U$26136 ( \26513 , \26511 , \26512 );
xor \U$26137 ( \26514 , \26427 , \26431 );
and \U$26138 ( \26515 , \26514 , \26436 );
and \U$26139 ( \26516 , \26427 , \26431 );
or \U$26140 ( \26517 , \26515 , \26516 );
not \U$26141 ( \26518 , \6611 );
not \U$26142 ( \26519 , \6561 );
and \U$26143 ( \26520 , \26518 , \26519 );
and \U$26144 ( \26521 , \6611 , \6561 );
nor \U$26145 ( \26522 , \26520 , \26521 );
not \U$26146 ( \26523 , \26522 );
not \U$26147 ( \26524 , \6475 );
not \U$26148 ( \26525 , \26524 );
and \U$26149 ( \26526 , \26523 , \26525 );
and \U$26150 ( \26527 , \26522 , \26524 );
nor \U$26151 ( \26528 , \26526 , \26527 );
xor \U$26152 ( \26529 , \26517 , \26528 );
xor \U$26153 ( \26530 , \26475 , \26477 );
and \U$26154 ( \26531 , \26530 , \26480 );
and \U$26155 ( \26532 , \26475 , \26477 );
or \U$26156 ( \26533 , \26531 , \26532 );
xor \U$26157 ( \26534 , \26529 , \26533 );
xor \U$26158 ( \26535 , \26513 , \26534 );
xor \U$26159 ( \26536 , \26437 , \26441 );
and \U$26160 ( \26537 , \26536 , \26452 );
and \U$26161 ( \26538 , \26437 , \26441 );
or \U$26162 ( \26539 , \26537 , \26538 );
xor \U$26163 ( \26540 , \26535 , \26539 );
xor \U$26164 ( \26541 , \26509 , \26540 );
xor \U$26165 ( \26542 , \26457 , \26482 );
and \U$26166 ( \26543 , \26542 , \26487 );
and \U$26167 ( \26544 , \26457 , \26482 );
or \U$26168 ( \26545 , \26543 , \26544 );
xor \U$26169 ( \26546 , \26541 , \26545 );
xor \U$26170 ( \26547 , \26453 , \26488 );
and \U$26171 ( \26548 , \26547 , \26493 );
and \U$26172 ( \26549 , \26453 , \26488 );
or \U$26173 ( \26550 , \26548 , \26549 );
nand \U$26174 ( \26551 , \26546 , \26550 );
xor \U$26175 ( \26552 , \26501 , \26503 );
and \U$26176 ( \26553 , \26552 , \26508 );
and \U$26177 ( \26554 , \26501 , \26503 );
or \U$26178 ( \26555 , \26553 , \26554 );
not \U$26179 ( \26556 , \6614 );
not \U$26180 ( \26557 , \6652 );
or \U$26181 ( \26558 , \26556 , \26557 );
nand \U$26182 ( \26559 , \6626 , \6653 );
nand \U$26183 ( \26560 , \26558 , \26559 );
not \U$26184 ( \26561 , \6650 );
and \U$26185 ( \26562 , \26560 , \26561 );
not \U$26186 ( \26563 , \26560 );
and \U$26187 ( \26564 , \26563 , \6650 );
nor \U$26188 ( \26565 , \26562 , \26564 );
xor \U$26189 ( \26566 , \26517 , \26528 );
and \U$26190 ( \26567 , \26566 , \26533 );
and \U$26191 ( \26568 , \26517 , \26528 );
or \U$26192 ( \26569 , \26567 , \26568 );
xor \U$26193 ( \26570 , \26565 , \26569 );
xnor \U$26194 ( \26571 , \6668 , \6916 );
and \U$26195 ( \26572 , \26571 , \6671 );
not \U$26196 ( \26573 , \26571 );
and \U$26197 ( \26574 , \26573 , \6919 );
nor \U$26198 ( \26575 , \26572 , \26574 );
xor \U$26199 ( \26576 , \26570 , \26575 );
xor \U$26200 ( \26577 , \26555 , \26576 );
xor \U$26201 ( \26578 , \26513 , \26534 );
and \U$26202 ( \26579 , \26578 , \26539 );
and \U$26203 ( \26580 , \26513 , \26534 );
or \U$26204 ( \26581 , \26579 , \26580 );
xor \U$26205 ( \26582 , \26577 , \26581 );
xor \U$26206 ( \26583 , \26509 , \26540 );
and \U$26207 ( \26584 , \26583 , \26545 );
and \U$26208 ( \26585 , \26509 , \26540 );
or \U$26209 ( \26586 , \26584 , \26585 );
nand \U$26210 ( \26587 , \26582 , \26586 );
xor \U$26211 ( \26588 , \6456 , \6458 );
xnor \U$26212 ( \26589 , \26588 , \6461 );
xor \U$26213 ( \26590 , \26565 , \26569 );
and \U$26214 ( \26591 , \26590 , \26575 );
and \U$26215 ( \26592 , \26565 , \26569 );
or \U$26216 ( \26593 , \26591 , \26592 );
xor \U$26217 ( \26594 , \26589 , \26593 );
xor \U$26218 ( \26595 , \6665 , \6655 );
xnor \U$26219 ( \26596 , \26595 , \6921 );
xor \U$26220 ( \26597 , \26594 , \26596 );
xor \U$26221 ( \26598 , \26555 , \26576 );
and \U$26222 ( \26599 , \26598 , \26581 );
and \U$26223 ( \26600 , \26555 , \26576 );
or \U$26224 ( \26601 , \26599 , \26600 );
nand \U$26225 ( \26602 , \26597 , \26601 );
xor \U$26226 ( \26603 , \6464 , \6925 );
xnor \U$26227 ( \26604 , \26603 , \6933 );
xor \U$26228 ( \26605 , \26589 , \26593 );
and \U$26229 ( \26606 , \26605 , \26596 );
and \U$26230 ( \26607 , \26589 , \26593 );
or \U$26231 ( \26608 , \26606 , \26607 );
nand \U$26232 ( \26609 , \26604 , \26608 );
and \U$26233 ( \26610 , \26551 , \26587 , \26602 , \26609 );
nand \U$26234 ( \26611 , \25824 , \26496 , \26610 );
not \U$26235 ( \26612 , \26611 );
nand \U$26236 ( \26613 , \22307 , \26612 );
not \U$26237 ( \26614 , \26496 );
not \U$26238 ( \26615 , \25823 );
not \U$26239 ( \26616 , \24070 );
not \U$26240 ( \26617 , \24135 );
nand \U$26241 ( \26618 , \24149 , \24141 );
not \U$26242 ( \26619 , \26618 );
nand \U$26243 ( \26620 , \26619 , \24127 );
not \U$26244 ( \26621 , \24101 );
not \U$26245 ( \26622 , \24126 );
nand \U$26246 ( \26623 , \26621 , \26622 );
nand \U$26247 ( \26624 , \26620 , \26623 );
not \U$26248 ( \26625 , \26624 );
or \U$26249 ( \26626 , \26617 , \26625 );
or \U$26250 ( \26627 , \24130 , \24134 );
nand \U$26251 ( \26628 , \26626 , \26627 );
not \U$26252 ( \26629 , \26628 );
or \U$26253 ( \26630 , \26616 , \26629 );
or \U$26254 ( \26631 , \23996 , \24069 );
nand \U$26255 ( \26632 , \26630 , \26631 );
not \U$26256 ( \26633 , \26632 );
or \U$26257 ( \26634 , \26615 , \26633 );
not \U$26258 ( \26635 , \25430 );
xor \U$26259 ( \26636 , \24410 , \24986 );
nor \U$26260 ( \26637 , \25003 , \26636 );
nand \U$26261 ( \26638 , \25006 , \25011 );
or \U$26262 ( \26639 , \26637 , \26638 );
xor \U$26263 ( \26640 , \24986 , \24410 );
nand \U$26264 ( \26641 , \26640 , \25003 );
nand \U$26265 ( \26642 , \26639 , \26641 );
not \U$26266 ( \26643 , \26642 );
or \U$26267 ( \26644 , \26635 , \26643 );
or \U$26268 ( \26645 , \25425 , \25429 );
nand \U$26269 ( \26646 , \26644 , \26645 );
buf \U$26270 ( \26647 , \25821 );
and \U$26271 ( \26648 , \26646 , \26647 );
nor \U$26272 ( \26649 , \25820 , \25816 );
nor \U$26273 ( \26650 , \26648 , \26649 );
nand \U$26274 ( \26651 , \26634 , \26650 );
not \U$26275 ( \26652 , \26651 );
or \U$26276 ( \26653 , \26614 , \26652 );
not \U$26277 ( \26654 , \26419 );
not \U$26278 ( \26655 , \26296 );
nor \U$26279 ( \26656 , \26298 , \26302 );
not \U$26280 ( \26657 , \26656 );
or \U$26281 ( \26658 , \26655 , \26657 );
or \U$26282 ( \26659 , \26276 , \26295 );
nand \U$26283 ( \26660 , \26658 , \26659 );
not \U$26284 ( \26661 , \26660 );
or \U$26285 ( \26662 , \26654 , \26661 );
or \U$26286 ( \26663 , \26414 , \26418 );
nand \U$26287 ( \26664 , \26662 , \26663 );
buf \U$26288 ( \26665 , \26495 );
and \U$26289 ( \26666 , \26664 , \26665 );
nor \U$26290 ( \26667 , \26423 , \26494 );
nor \U$26291 ( \26668 , \26666 , \26667 );
nand \U$26292 ( \26669 , \26653 , \26668 );
nand \U$26293 ( \26670 , \26669 , \26610 );
nand \U$26294 ( \26671 , \26613 , \26670 );
not \U$26295 ( \26672 , \5509 );
not \U$26296 ( \26673 , RIc2264d0_37);
not \U$26297 ( \26674 , \23758 );
or \U$26298 ( \26675 , \26673 , \26674 );
not \U$26299 ( \26676 , RIc2264d0_37);
nand \U$26300 ( \26677 , \26676 , \6718 );
nand \U$26301 ( \26678 , \26675 , \26677 );
not \U$26302 ( \26679 , \26678 );
or \U$26303 ( \26680 , \26672 , \26679 );
not \U$26304 ( \26681 , \6492 );
xor \U$26305 ( \26682 , \4371 , \26681 );
nand \U$26306 ( \26683 , \26682 , \5519 );
nand \U$26307 ( \26684 , \26680 , \26683 );
not \U$26308 ( \26685 , \6688 );
not \U$26309 ( \26686 , RIc2263e0_39);
not \U$26310 ( \26687 , \13687 );
or \U$26311 ( \26688 , \26686 , \26687 );
nand \U$26312 ( \26689 , \9769 , \6694 );
nand \U$26313 ( \26690 , \26688 , \26689 );
not \U$26314 ( \26691 , \26690 );
or \U$26315 ( \26692 , \26685 , \26691 );
not \U$26316 ( \26693 , RIc2263e0_39);
not \U$26317 ( \26694 , \5664 );
or \U$26318 ( \26695 , \26693 , \26694 );
nand \U$26319 ( \26696 , \5663 , \25483 );
nand \U$26320 ( \26697 , \26695 , \26696 );
nand \U$26321 ( \26698 , \26697 , \6307 );
nand \U$26322 ( \26699 , \26692 , \26698 );
xor \U$26323 ( \26700 , \26684 , \26699 );
not \U$26324 ( \26701 , \9690 );
not \U$26325 ( \26702 , RIc2262f0_41);
not \U$26326 ( \26703 , \5216 );
or \U$26327 ( \26704 , \26702 , \26703 );
nand \U$26328 ( \26705 , \15007 , \17820 );
nand \U$26329 ( \26706 , \26704 , \26705 );
not \U$26330 ( \26707 , \26706 );
or \U$26331 ( \26708 , \26701 , \26707 );
not \U$26332 ( \26709 , RIc2262f0_41);
not \U$26333 ( \26710 , \6076 );
or \U$26334 ( \26711 , \26709 , \26710 );
nand \U$26335 ( \26712 , \4406 , \6303 );
nand \U$26336 ( \26713 , \26711 , \26712 );
nand \U$26337 ( \26714 , \26713 , \9816 );
nand \U$26338 ( \26715 , \26708 , \26714 );
xnor \U$26339 ( \26716 , \26700 , \26715 );
not \U$26340 ( \26717 , \26716 );
not \U$26341 ( \26718 , \2697 );
xor \U$26342 ( \26719 , RIc2267a0_31, \8951 );
not \U$26343 ( \26720 , \26719 );
or \U$26344 ( \26721 , \26718 , \26720 );
and \U$26345 ( \26722 , RIc2267a0_31, \10295 );
not \U$26346 ( \26723 , RIc2267a0_31);
and \U$26347 ( \26724 , \26723 , \8806 );
or \U$26348 ( \26725 , \26722 , \26724 );
nand \U$26349 ( \26726 , \26725 , \2710 );
nand \U$26350 ( \26727 , \26721 , \26726 );
not \U$26351 ( \26728 , \2784 );
and \U$26352 ( \26729 , RIc226890_29, \8910 );
not \U$26353 ( \26730 , RIc226890_29);
and \U$26354 ( \26731 , \26730 , \14968 );
or \U$26355 ( \26732 , \26729 , \26731 );
not \U$26356 ( \26733 , \26732 );
or \U$26357 ( \26734 , \26728 , \26733 );
and \U$26358 ( \26735 , RIc226890_29, \8978 );
not \U$26359 ( \26736 , RIc226890_29);
and \U$26360 ( \26737 , \26736 , \10748 );
nor \U$26361 ( \26738 , \26735 , \26737 );
not \U$26362 ( \26739 , \26738 );
nand \U$26363 ( \26740 , \26739 , \9142 );
nand \U$26364 ( \26741 , \26734 , \26740 );
xor \U$26365 ( \26742 , \26727 , \26741 );
not \U$26366 ( \26743 , \9205 );
not \U$26367 ( \26744 , RIc226200_43);
not \U$26368 ( \26745 , \4049 );
or \U$26369 ( \26746 , \26744 , \26745 );
nand \U$26370 ( \26747 , \3640 , \13805 );
nand \U$26371 ( \26748 , \26746 , \26747 );
not \U$26372 ( \26749 , \26748 );
or \U$26373 ( \26750 , \26743 , \26749 );
not \U$26374 ( \26751 , RIc226200_43);
not \U$26375 ( \26752 , \4417 );
or \U$26376 ( \26753 , \26751 , \26752 );
nand \U$26377 ( \26754 , \16519 , \9117 );
nand \U$26378 ( \26755 , \26753 , \26754 );
nand \U$26379 ( \26756 , \26755 , \9110 );
nand \U$26380 ( \26757 , \26750 , \26756 );
xor \U$26381 ( \26758 , \26742 , \26757 );
not \U$26382 ( \26759 , \26758 );
not \U$26383 ( \26760 , \26759 );
or \U$26384 ( \26761 , \26717 , \26760 );
not \U$26385 ( \26762 , \1963 );
not \U$26386 ( \26763 , RIc226e30_17);
not \U$26387 ( \26764 , \20693 );
or \U$26388 ( \26765 , \26763 , \26764 );
nand \U$26389 ( \26766 , \12755 , \1960 );
nand \U$26390 ( \26767 , \26765 , \26766 );
not \U$26391 ( \26768 , \26767 );
or \U$26392 ( \26769 , \26762 , \26768 );
not \U$26393 ( \26770 , RIc226e30_17);
not \U$26394 ( \26771 , \15444 );
or \U$26395 ( \26772 , \26770 , \26771 );
nand \U$26396 ( \26773 , \12825 , \1960 );
nand \U$26397 ( \26774 , \26772 , \26773 );
nand \U$26398 ( \26775 , \26774 , \1945 );
nand \U$26399 ( \26776 , \26769 , \26775 );
and \U$26400 ( \26777 , \16248 , \1681 );
not \U$26401 ( \26778 , \26777 );
not \U$26402 ( \26779 , \2318 );
and \U$26403 ( \26780 , \13487 , \2351 );
not \U$26404 ( \26781 , \13487 );
and \U$26405 ( \26782 , \26781 , RIc226f20_15);
or \U$26406 ( \26783 , \26780 , \26782 );
not \U$26407 ( \26784 , \26783 );
or \U$26408 ( \26785 , \26779 , \26784 );
not \U$26409 ( \26786 , RIc226f20_15);
not \U$26410 ( \26787 , \16259 );
or \U$26411 ( \26788 , \26786 , \26787 );
nand \U$26412 ( \26789 , \16482 , \1674 );
nand \U$26413 ( \26790 , \26788 , \26789 );
nand \U$26414 ( \26791 , \26790 , \2319 );
nand \U$26415 ( \26792 , \26785 , \26791 );
not \U$26416 ( \26793 , \26792 );
nand \U$26417 ( \26794 , \26778 , \26793 );
not \U$26418 ( \26795 , \26794 );
not \U$26419 ( \26796 , \1945 );
not \U$26420 ( \26797 , RIc226e30_17);
not \U$26421 ( \26798 , \18158 );
or \U$26422 ( \26799 , \26797 , \26798 );
nand \U$26423 ( \26800 , \18161 , \1960 );
nand \U$26424 ( \26801 , \26799 , \26800 );
not \U$26425 ( \26802 , \26801 );
or \U$26426 ( \26803 , \26796 , \26802 );
nand \U$26427 ( \26804 , \26774 , \1963 );
nand \U$26428 ( \26805 , \26803 , \26804 );
not \U$26429 ( \26806 , \26805 );
or \U$26430 ( \26807 , \26795 , \26806 );
nand \U$26431 ( \26808 , \26792 , \26777 );
nand \U$26432 ( \26809 , \26807 , \26808 );
xor \U$26433 ( \26810 , \26776 , \26809 );
not \U$26434 ( \26811 , \2154 );
and \U$26435 ( \26812 , RIc226980_27, \9224 );
not \U$26436 ( \26813 , RIc226980_27);
and \U$26437 ( \26814 , \26813 , \9050 );
or \U$26438 ( \26815 , \26812 , \26814 );
not \U$26439 ( \26816 , \26815 );
or \U$26440 ( \26817 , \26811 , \26816 );
not \U$26441 ( \26818 , RIc226980_27);
not \U$26442 ( \26819 , \10652 );
or \U$26443 ( \26820 , \26818 , \26819 );
nand \U$26444 ( \26821 , \9072 , \2150 );
nand \U$26445 ( \26822 , \26820 , \26821 );
nand \U$26446 ( \26823 , \26822 , \2138 );
nand \U$26447 ( \26824 , \26817 , \26823 );
xor \U$26448 ( \26825 , \26810 , \26824 );
not \U$26449 ( \26826 , \9459 );
not \U$26450 ( \26827 , RIc225e40_51);
not \U$26451 ( \26828 , \12977 );
or \U$26452 ( \26829 , \26827 , \26828 );
nand \U$26453 ( \26830 , \3008 , \11795 );
nand \U$26454 ( \26831 , \26829 , \26830 );
not \U$26455 ( \26832 , \26831 );
or \U$26456 ( \26833 , \26826 , \26832 );
not \U$26457 ( \26834 , RIc225e40_51);
not \U$26458 ( \26835 , \2670 );
or \U$26459 ( \26836 , \26834 , \26835 );
nand \U$26460 ( \26837 , \16642 , \9450 );
nand \U$26461 ( \26838 , \26836 , \26837 );
nand \U$26462 ( \26839 , \26838 , \9444 );
nand \U$26463 ( \26840 , \26833 , \26839 );
xor \U$26464 ( \26841 , \26825 , \26840 );
not \U$26465 ( \26842 , \15164 );
and \U$26466 ( \26843 , RIc225a80_59, \4009 );
not \U$26467 ( \26844 , RIc225a80_59);
and \U$26468 ( \26845 , \26844 , \9608 );
or \U$26469 ( \26846 , \26843 , \26845 );
not \U$26470 ( \26847 , \26846 );
or \U$26471 ( \26848 , \26842 , \26847 );
and \U$26472 ( \26849 , RIc225a80_59, \16762 );
not \U$26473 ( \26850 , RIc225a80_59);
and \U$26474 ( \26851 , \26850 , \9600 );
or \U$26475 ( \26852 , \26849 , \26851 );
nand \U$26476 ( \26853 , \26852 , \12670 );
nand \U$26477 ( \26854 , \26848 , \26853 );
and \U$26478 ( \26855 , \26841 , \26854 );
and \U$26479 ( \26856 , \26825 , \26840 );
or \U$26480 ( \26857 , \26855 , \26856 );
nand \U$26481 ( \26858 , \26761 , \26857 );
not \U$26482 ( \26859 , \26716 );
nand \U$26483 ( \26860 , \26859 , \26758 );
nand \U$26484 ( \26861 , \26858 , \26860 );
or \U$26485 ( \26862 , RIc227088_12, RIc227010_13);
nand \U$26486 ( \26863 , \26862 , \18357 );
and \U$26487 ( \26864 , RIc227088_12, RIc227010_13);
nor \U$26488 ( \26865 , \26864 , \1291 );
and \U$26489 ( \26866 , \26863 , \26865 );
not \U$26490 ( \26867 , \1310 );
not \U$26491 ( \26868 , RIc227100_11);
not \U$26492 ( \26869 , \21102 );
or \U$26493 ( \26870 , \26868 , \26869 );
nand \U$26494 ( \26871 , \16482 , \1685 );
nand \U$26495 ( \26872 , \26870 , \26871 );
not \U$26496 ( \26873 , \26872 );
or \U$26497 ( \26874 , \26867 , \26873 );
or \U$26498 ( \26875 , \16248 , \3351 );
or \U$26499 ( \26876 , \18181 , RIc227100_11);
nand \U$26500 ( \26877 , \26875 , \26876 );
nand \U$26501 ( \26878 , \26877 , \1306 );
nand \U$26502 ( \26879 , \26874 , \26878 );
xor \U$26503 ( \26880 , \26866 , \26879 );
not \U$26504 ( \26881 , \1682 );
not \U$26505 ( \26882 , RIc227010_13);
not \U$26506 ( \26883 , \18158 );
or \U$26507 ( \26884 , \26882 , \26883 );
nand \U$26508 ( \26885 , \18161 , \2427 );
nand \U$26509 ( \26886 , \26884 , \26885 );
not \U$26510 ( \26887 , \26886 );
or \U$26511 ( \26888 , \26881 , \26887 );
not \U$26512 ( \26889 , RIc227010_13);
not \U$26513 ( \26890 , \20392 );
or \U$26514 ( \26891 , \26889 , \26890 );
nand \U$26515 ( \26892 , \13487 , \1758 );
nand \U$26516 ( \26893 , \26891 , \26892 );
nand \U$26517 ( \26894 , \26893 , \1678 );
nand \U$26518 ( \26895 , \26888 , \26894 );
xor \U$26519 ( \26896 , \26880 , \26895 );
not \U$26520 ( \26897 , \1963 );
not \U$26521 ( \26898 , RIc226e30_17);
not \U$26522 ( \26899 , \10198 );
or \U$26523 ( \26900 , \26898 , \26899 );
nand \U$26524 ( \26901 , \10197 , \1960 );
nand \U$26525 ( \26902 , \26900 , \26901 );
not \U$26526 ( \26903 , \26902 );
or \U$26527 ( \26904 , \26897 , \26903 );
not \U$26528 ( \26905 , RIc226e30_17);
not \U$26529 ( \26906 , \21084 );
or \U$26530 ( \26907 , \26905 , \26906 );
nand \U$26531 ( \26908 , \13497 , \1960 );
nand \U$26532 ( \26909 , \26907 , \26908 );
nand \U$26533 ( \26910 , \26909 , \1945 );
nand \U$26534 ( \26911 , \26904 , \26910 );
xor \U$26535 ( \26912 , \26896 , \26911 );
not \U$26536 ( \26913 , \5519 );
not \U$26537 ( \26914 , RIc2264d0_37);
not \U$26538 ( \26915 , \16555 );
or \U$26539 ( \26916 , \26914 , \26915 );
nand \U$26540 ( \26917 , \6071 , \5504 );
nand \U$26541 ( \26918 , \26916 , \26917 );
not \U$26542 ( \26919 , \26918 );
or \U$26543 ( \26920 , \26913 , \26919 );
nand \U$26544 ( \26921 , \26682 , \5509 );
nand \U$26545 ( \26922 , \26920 , \26921 );
xor \U$26546 ( \26923 , \26912 , \26922 );
not \U$26547 ( \26924 , \4383 );
not \U$26548 ( \26925 , RIc2265c0_35);
not \U$26549 ( \26926 , \9859 );
or \U$26550 ( \26927 , \26925 , \26926 );
not \U$26551 ( \26928 , \23758 );
nand \U$26552 ( \26929 , \26928 , \4376 );
nand \U$26553 ( \26930 , \26927 , \26929 );
not \U$26554 ( \26931 , \26930 );
or \U$26555 ( \26932 , \26924 , \26931 );
and \U$26556 ( \26933 , \3620 , \10609 );
not \U$26557 ( \26934 , \3620 );
and \U$26558 ( \26935 , \26934 , \10141 );
nor \U$26559 ( \26936 , \26933 , \26935 );
nand \U$26560 ( \26937 , \26936 , \4381 );
nand \U$26561 ( \26938 , \26932 , \26937 );
xor \U$26562 ( \26939 , \26923 , \26938 );
not \U$26563 ( \26940 , \2154 );
not \U$26564 ( \26941 , RIc226980_27);
not \U$26565 ( \26942 , \8910 );
or \U$26566 ( \26943 , \26941 , \26942 );
nand \U$26567 ( \26944 , \12406 , \2150 );
nand \U$26568 ( \26945 , \26943 , \26944 );
not \U$26569 ( \26946 , \26945 );
or \U$26570 ( \26947 , \26940 , \26946 );
not \U$26571 ( \26948 , RIc226980_27);
not \U$26572 ( \26949 , \9215 );
or \U$26573 ( \26950 , \26948 , \26949 );
nand \U$26574 ( \26951 , \9211 , \2150 );
nand \U$26575 ( \26952 , \26950 , \26951 );
nand \U$26576 ( \26953 , \26952 , \2138 );
nand \U$26577 ( \26954 , \26947 , \26953 );
not \U$26578 ( \26955 , \2710 );
not \U$26579 ( \26956 , RIc2267a0_31);
not \U$26580 ( \26957 , \9897 );
or \U$26581 ( \26958 , \26956 , \26957 );
nand \U$26582 ( \26959 , \8829 , \3648 );
nand \U$26583 ( \26960 , \26958 , \26959 );
not \U$26584 ( \26961 , \26960 );
or \U$26585 ( \26962 , \26955 , \26961 );
nand \U$26586 ( \26963 , \26725 , \2697 );
nand \U$26587 ( \26964 , \26962 , \26963 );
not \U$26588 ( \26965 , \26964 );
and \U$26589 ( \26966 , \26954 , \26965 );
not \U$26590 ( \26967 , \26954 );
not \U$26591 ( \26968 , \2710 );
not \U$26592 ( \26969 , \26960 );
or \U$26593 ( \26970 , \26968 , \26969 );
nand \U$26594 ( \26971 , \26970 , \26963 );
and \U$26595 ( \26972 , \26967 , \26971 );
or \U$26596 ( \26973 , \26966 , \26972 );
not \U$26597 ( \26974 , \26738 );
not \U$26598 ( \26975 , \2077 );
and \U$26599 ( \26976 , \26974 , \26975 );
and \U$26600 ( \26977 , RIc226890_29, \20367 );
not \U$26601 ( \26978 , RIc226890_29);
and \U$26602 ( \26979 , \26978 , \8951 );
or \U$26603 ( \26980 , \26977 , \26979 );
and \U$26604 ( \26981 , \26980 , \9142 );
nor \U$26605 ( \26982 , \26976 , \26981 );
buf \U$26606 ( \26983 , \26982 );
not \U$26607 ( \26984 , \26983 );
and \U$26608 ( \26985 , \26973 , \26984 );
not \U$26609 ( \26986 , \26973 );
and \U$26610 ( \26987 , \26986 , \26983 );
nor \U$26611 ( \26988 , \26985 , \26987 );
xor \U$26612 ( \26989 , \26939 , \26988 );
not \U$26613 ( \26990 , \9690 );
not \U$26614 ( \26991 , \26713 );
or \U$26615 ( \26992 , \26990 , \26991 );
not \U$26616 ( \26993 , \9822 );
not \U$26617 ( \26994 , \10209 );
or \U$26618 ( \26995 , \26993 , \26994 );
not \U$26619 ( \26996 , \16519 );
nand \U$26620 ( \26997 , \26996 , RIc2262f0_41);
nand \U$26621 ( \26998 , \26995 , \26997 );
nand \U$26622 ( \26999 , \26998 , \9705 );
nand \U$26623 ( \27000 , \26992 , \26999 );
not \U$26624 ( \27001 , \3631 );
not \U$26625 ( \27002 , RIc2266b0_33);
not \U$26626 ( \27003 , \8887 );
or \U$26627 ( \27004 , \27002 , \27003 );
nand \U$26628 ( \27005 , \8886 , \5179 );
nand \U$26629 ( \27006 , \27004 , \27005 );
not \U$26630 ( \27007 , \27006 );
or \U$26631 ( \27008 , \27001 , \27007 );
not \U$26632 ( \27009 , RIc2266b0_33);
not \U$26633 ( \27010 , \12724 );
or \U$26634 ( \27011 , \27009 , \27010 );
nand \U$26635 ( \27012 , \12727 , \9425 );
nand \U$26636 ( \27013 , \27011 , \27012 );
nand \U$26637 ( \27014 , \27013 , \3629 );
nand \U$26638 ( \27015 , \27008 , \27014 );
xor \U$26639 ( \27016 , \27000 , \27015 );
not \U$26640 ( \27017 , \26697 );
not \U$26641 ( \27018 , \27017 );
not \U$26642 ( \27019 , \6313 );
and \U$26643 ( \27020 , \27018 , \27019 );
not \U$26644 ( \27021 , \5498 );
not \U$26645 ( \27022 , \18459 );
or \U$26646 ( \27023 , \27021 , \27022 );
not \U$26647 ( \27024 , \10231 );
nand \U$26648 ( \27025 , \27024 , RIc2263e0_39);
nand \U$26649 ( \27026 , \27023 , \27025 );
and \U$26650 ( \27027 , \27026 , \6307 );
nor \U$26651 ( \27028 , \27020 , \27027 );
xnor \U$26652 ( \27029 , \27016 , \27028 );
xor \U$26653 ( \27030 , \26989 , \27029 );
xor \U$26654 ( \27031 , \26861 , \27030 );
not \U$26655 ( \27032 , \9552 );
not \U$26656 ( \27033 , RIc225f30_49);
not \U$26657 ( \27034 , \3009 );
or \U$26658 ( \27035 , \27033 , \27034 );
nand \U$26659 ( \27036 , \11844 , \9549 );
nand \U$26660 ( \27037 , \27035 , \27036 );
not \U$26661 ( \27038 , \27037 );
or \U$26662 ( \27039 , \27032 , \27038 );
not \U$26663 ( \27040 , RIc225f30_49);
not \U$26664 ( \27041 , \5526 );
or \U$26665 ( \27042 , \27040 , \27041 );
nand \U$26666 ( \27043 , \2042 , \9541 );
nand \U$26667 ( \27044 , \27042 , \27043 );
nand \U$26668 ( \27045 , \27044 , \10445 );
nand \U$26669 ( \27046 , \27039 , \27045 );
not \U$26670 ( \27047 , \11974 );
and \U$26671 ( \27048 , RIc225b70_57, \2258 );
not \U$26672 ( \27049 , RIc225b70_57);
and \U$26673 ( \27050 , \27049 , \9608 );
or \U$26674 ( \27051 , \27048 , \27050 );
not \U$26675 ( \27052 , \27051 );
or \U$26676 ( \27053 , \27047 , \27052 );
not \U$26677 ( \27054 , RIc225b70_57);
not \U$26678 ( \27055 , \12508 );
or \U$26679 ( \27056 , \27054 , \27055 );
nand \U$26680 ( \27057 , \1988 , \11033 );
nand \U$26681 ( \27058 , \27056 , \27057 );
nand \U$26682 ( \27059 , \27058 , \11965 );
nand \U$26683 ( \27060 , \27053 , \27059 );
and \U$26684 ( \27061 , \27046 , \27060 );
not \U$26685 ( \27062 , \27046 );
not \U$26686 ( \27063 , \27060 );
and \U$26687 ( \27064 , \27062 , \27063 );
nor \U$26688 ( \27065 , \27061 , \27064 );
not \U$26689 ( \27066 , \12304 );
not \U$26690 ( \27067 , RIc226020_47);
not \U$26691 ( \27068 , \9804 );
or \U$26692 ( \27069 , \27067 , \27068 );
nand \U$26693 ( \27070 , \9805 , \9373 );
nand \U$26694 ( \27071 , \27069 , \27070 );
not \U$26695 ( \27072 , \27071 );
or \U$26696 ( \27073 , \27066 , \27072 );
and \U$26697 ( \27074 , RIc226020_47, \10532 );
not \U$26698 ( \27075 , RIc226020_47);
and \U$26699 ( \27076 , \27075 , \9654 );
or \U$26700 ( \27077 , \27074 , \27076 );
nand \U$26701 ( \27078 , \27077 , \9641 );
nand \U$26702 ( \27079 , \27073 , \27078 );
and \U$26703 ( \27080 , \27065 , \27079 );
not \U$26704 ( \27081 , \27065 );
not \U$26705 ( \27082 , \27079 );
and \U$26706 ( \27083 , \27081 , \27082 );
or \U$26707 ( \27084 , \27080 , \27083 );
not \U$26708 ( \27085 , \27084 );
and \U$26709 ( \27086 , \2421 , \12806 );
not \U$26710 ( \27087 , \2421 );
and \U$26711 ( \27088 , \27087 , RIc225990_61);
or \U$26712 ( \27089 , \27086 , \27088 );
and \U$26713 ( \27090 , \27089 , \15719 );
and \U$26714 ( \27091 , \10933 , \12806 );
not \U$26715 ( \27092 , \10933 );
and \U$26716 ( \27093 , \27092 , RIc225990_61);
or \U$26717 ( \27094 , \27091 , \27093 );
and \U$26718 ( \27095 , \27094 , \15729 );
nor \U$26719 ( \27096 , \27090 , \27095 );
not \U$26720 ( \27097 , \3115 );
not \U$26721 ( \27098 , \22795 );
and \U$26722 ( \27099 , \27097 , \27098 );
and \U$26723 ( \27100 , \3115 , \22795 );
nor \U$26724 ( \27101 , \27099 , \27100 );
not \U$26725 ( \27102 , \27101 );
not \U$26726 ( \27103 , \23212 );
and \U$26727 ( \27104 , \27102 , \27103 );
not \U$26728 ( \27105 , RIc226110_45);
not \U$26729 ( \27106 , \10496 );
or \U$26730 ( \27107 , \27105 , \27106 );
nand \U$26731 ( \27108 , \3725 , \14660 );
nand \U$26732 ( \27109 , \27107 , \27108 );
and \U$26733 ( \27110 , \27109 , \9384 );
nor \U$26734 ( \27111 , \27104 , \27110 );
xor \U$26735 ( \27112 , \27096 , \27111 );
not \U$26736 ( \27113 , RIc225c60_55);
not \U$26737 ( \27114 , \11890 );
or \U$26738 ( \27115 , \27113 , \27114 );
nand \U$26739 ( \27116 , \2014 , \8767 );
nand \U$26740 ( \27117 , \27115 , \27116 );
and \U$26741 ( \27118 , \27117 , \13025 );
and \U$26742 ( \27119 , \2585 , \11108 );
not \U$26743 ( \27120 , \2585 );
and \U$26744 ( \27121 , \27120 , RIc225c60_55);
or \U$26745 ( \27122 , \27119 , \27121 );
and \U$26746 ( \27123 , \27122 , \11697 );
nor \U$26747 ( \27124 , \27118 , \27123 );
xor \U$26748 ( \27125 , \27112 , \27124 );
not \U$26749 ( \27126 , \27125 );
or \U$26750 ( \27127 , \27085 , \27126 );
or \U$26751 ( \27128 , RIc226f98_14, RIc226f20_15);
nand \U$26752 ( \27129 , \27128 , \16248 );
and \U$26753 ( \27130 , RIc226f98_14, RIc226f20_15);
nor \U$26754 ( \27131 , \27130 , \1758 );
and \U$26755 ( \27132 , \27129 , \27131 );
not \U$26756 ( \27133 , \1682 );
not \U$26757 ( \27134 , RIc227010_13);
not \U$26758 ( \27135 , \21102 );
or \U$26759 ( \27136 , \27134 , \27135 );
nand \U$26760 ( \27137 , \16482 , \1758 );
nand \U$26761 ( \27138 , \27136 , \27137 );
not \U$26762 ( \27139 , \27138 );
or \U$26763 ( \27140 , \27133 , \27139 );
or \U$26764 ( \27141 , \16248 , \1758 );
or \U$26765 ( \27142 , \21954 , RIc227010_13);
nand \U$26766 ( \27143 , \27141 , \27142 );
nand \U$26767 ( \27144 , \27143 , \1677 );
nand \U$26768 ( \27145 , \27140 , \27144 );
and \U$26769 ( \27146 , \27132 , \27145 );
not \U$26770 ( \27147 , \1945 );
not \U$26771 ( \27148 , \26767 );
or \U$26772 ( \27149 , \27147 , \27148 );
nand \U$26773 ( \27150 , \26909 , \1963 );
nand \U$26774 ( \27151 , \27149 , \27150 );
xor \U$26775 ( \27152 , \27146 , \27151 );
not \U$26776 ( \27153 , \2534 );
not \U$26777 ( \27154 , RIc226d40_19);
not \U$26778 ( \27155 , \10360 );
or \U$26779 ( \27156 , \27154 , \27155 );
nand \U$26780 ( \27157 , \10086 , \1941 );
nand \U$26781 ( \27158 , \27156 , \27157 );
not \U$26782 ( \27159 , \27158 );
or \U$26783 ( \27160 , \27153 , \27159 );
not \U$26784 ( \27161 , RIc226d40_19);
not \U$26785 ( \27162 , \10369 );
or \U$26786 ( \27163 , \27161 , \27162 );
nand \U$26787 ( \27164 , \10370 , \3338 );
nand \U$26788 ( \27165 , \27163 , \27164 );
nand \U$26789 ( \27166 , \27165 , \2518 );
nand \U$26790 ( \27167 , \27160 , \27166 );
xor \U$26791 ( \27168 , \27152 , \27167 );
not \U$26792 ( \27169 , \9555 );
and \U$26793 ( \27170 , RIc225d50_53, \2555 );
not \U$26794 ( \27171 , RIc225d50_53);
and \U$26795 ( \27172 , \27171 , \9942 );
or \U$26796 ( \27173 , \27170 , \27172 );
not \U$26797 ( \27174 , \27173 );
or \U$26798 ( \27175 , \27169 , \27174 );
not \U$26799 ( \27176 , RIc225d50_53);
not \U$26800 ( \27177 , \15382 );
or \U$26801 ( \27178 , \27176 , \27177 );
nand \U$26802 ( \27179 , \2475 , \8772 );
nand \U$26803 ( \27180 , \27178 , \27179 );
nand \U$26804 ( \27181 , \27180 , \8777 );
nand \U$26805 ( \27182 , \27175 , \27181 );
xor \U$26806 ( \27183 , \27168 , \27182 );
not \U$26807 ( \27184 , \15164 );
not \U$26808 ( \27185 , \26852 );
or \U$26809 ( \27186 , \27184 , \27185 );
and \U$26810 ( \27187 , RIc225a80_59, \9570 );
not \U$26811 ( \27188 , RIc225a80_59);
and \U$26812 ( \27189 , \27188 , \2443 );
or \U$26813 ( \27190 , \27187 , \27189 );
nand \U$26814 ( \27191 , \27190 , \12670 );
nand \U$26815 ( \27192 , \27186 , \27191 );
xor \U$26816 ( \27193 , \27183 , \27192 );
nand \U$26817 ( \27194 , \27127 , \27193 );
not \U$26818 ( \27195 , \27125 );
not \U$26819 ( \27196 , \27084 );
nand \U$26820 ( \27197 , \27195 , \27196 );
nand \U$26821 ( \27198 , \27194 , \27197 );
and \U$26822 ( \27199 , \27031 , \27198 );
and \U$26823 ( \27200 , \26861 , \27030 );
or \U$26824 ( \27201 , \27199 , \27200 );
and \U$26825 ( \27202 , \18357 , \1310 );
not \U$26826 ( \27203 , \1682 );
not \U$26827 ( \27204 , \26893 );
or \U$26828 ( \27205 , \27203 , \27204 );
nand \U$26829 ( \27206 , \27138 , \1678 );
nand \U$26830 ( \27207 , \27205 , \27206 );
xor \U$26831 ( \27208 , \27202 , \27207 );
and \U$26832 ( \27209 , RIc226f20_15, \15444 );
not \U$26833 ( \27210 , RIc226f20_15);
and \U$26834 ( \27211 , \27210 , \19721 );
nor \U$26835 ( \27212 , \27209 , \27211 );
not \U$26836 ( \27213 , \2318 );
or \U$26837 ( \27214 , \27212 , \27213 );
not \U$26838 ( \27215 , RIc226f20_15);
not \U$26839 ( \27216 , \18158 );
or \U$26840 ( \27217 , \27215 , \27216 );
nand \U$26841 ( \27218 , \18161 , \2301 );
nand \U$26842 ( \27219 , \27217 , \27218 );
nand \U$26843 ( \27220 , \27219 , \2320 );
nand \U$26844 ( \27221 , \27214 , \27220 );
and \U$26845 ( \27222 , \27208 , \27221 );
and \U$26846 ( \27223 , \27202 , \27207 );
or \U$26847 ( \27224 , \27222 , \27223 );
not \U$26848 ( \27225 , \2358 );
and \U$26849 ( \27226 , RIc226f20_15, \16042 );
not \U$26850 ( \27227 , RIc226f20_15);
and \U$26851 ( \27228 , \27227 , \12755 );
or \U$26852 ( \27229 , \27226 , \27228 );
not \U$26853 ( \27230 , \27229 );
or \U$26854 ( \27231 , \27225 , \27230 );
or \U$26855 ( \27232 , \27212 , \2321 );
nand \U$26856 ( \27233 , \27231 , \27232 );
xor \U$26857 ( \27234 , \27224 , \27233 );
not \U$26858 ( \27235 , \10214 );
not \U$26859 ( \27236 , RIc226b60_23);
not \U$26860 ( \27237 , \9251 );
or \U$26861 ( \27238 , \27236 , \27237 );
buf \U$26862 ( \27239 , \17014 );
nand \U$26863 ( \27240 , \27239 , \1911 );
nand \U$26864 ( \27241 , \27238 , \27240 );
not \U$26865 ( \27242 , \27241 );
or \U$26866 ( \27243 , \27235 , \27242 );
not \U$26867 ( \27244 , RIc226b60_23);
not \U$26868 ( \27245 , \10814 );
or \U$26869 ( \27246 , \27244 , \27245 );
nand \U$26870 ( \27247 , \10110 , \2111 );
nand \U$26871 ( \27248 , \27246 , \27247 );
nand \U$26872 ( \27249 , \27248 , \1930 );
nand \U$26873 ( \27250 , \27243 , \27249 );
and \U$26874 ( \27251 , \27234 , \27250 );
and \U$26875 ( \27252 , \27224 , \27233 );
or \U$26876 ( \27253 , \27251 , \27252 );
nand \U$26877 ( \27254 , \26982 , \26965 );
and \U$26878 ( \27255 , \27254 , \26954 );
nor \U$26879 ( \27256 , \26982 , \26965 );
nor \U$26880 ( \27257 , \27255 , \27256 );
xor \U$26881 ( \27258 , \27253 , \27257 );
not \U$26882 ( \27259 , \27000 );
nand \U$26883 ( \27260 , \27259 , \27028 );
and \U$26884 ( \27261 , \27260 , \27015 );
not \U$26885 ( \27262 , \27000 );
nor \U$26886 ( \27263 , \27262 , \27028 );
nor \U$26887 ( \27264 , \27261 , \27263 );
xor \U$26888 ( \27265 , \27258 , \27264 );
not \U$26889 ( \27266 , \2195 );
not \U$26890 ( \27267 , RIc226a70_25);
not \U$26891 ( \27268 , \9073 );
or \U$26892 ( \27269 , \27267 , \27268 );
nand \U$26893 ( \27270 , \9072 , \1905 );
nand \U$26894 ( \27271 , \27269 , \27270 );
not \U$26895 ( \27272 , \27271 );
or \U$26896 ( \27273 , \27266 , \27272 );
not \U$26897 ( \27274 , RIc226a70_25);
not \U$26898 ( \27275 , \9046 );
or \U$26899 ( \27276 , \27274 , \27275 );
nand \U$26900 ( \27277 , \10644 , \2187 );
nand \U$26901 ( \27278 , \27276 , \27277 );
nand \U$26902 ( \27279 , \27278 , \2173 );
nand \U$26903 ( \27280 , \27273 , \27279 );
not \U$26904 ( \27281 , \2392 );
not \U$26905 ( \27282 , RIc226c50_21);
not \U$26906 ( \27283 , \9300 );
or \U$26907 ( \27284 , \27282 , \27283 );
nand \U$26908 ( \27285 , \21150 , \10834 );
nand \U$26909 ( \27286 , \27284 , \27285 );
not \U$26910 ( \27287 , \27286 );
or \U$26911 ( \27288 , \27281 , \27287 );
not \U$26912 ( \27289 , RIc226c50_21);
not \U$26913 ( \27290 , \10800 );
or \U$26914 ( \27291 , \27289 , \27290 );
nand \U$26915 ( \27292 , \9275 , \2370 );
nand \U$26916 ( \27293 , \27291 , \27292 );
nand \U$26917 ( \27294 , \27293 , \2367 );
nand \U$26918 ( \27295 , \27288 , \27294 );
not \U$26919 ( \27296 , \2534 );
not \U$26920 ( \27297 , RIc226d40_19);
not \U$26921 ( \27298 , \12100 );
or \U$26922 ( \27299 , \27297 , \27298 );
nand \U$26923 ( \27300 , \9320 , \2523 );
nand \U$26924 ( \27301 , \27299 , \27300 );
not \U$26925 ( \27302 , \27301 );
or \U$26926 ( \27303 , \27296 , \27302 );
nand \U$26927 ( \27304 , \27158 , \2518 );
nand \U$26928 ( \27305 , \27303 , \27304 );
xor \U$26929 ( \27306 , \27295 , \27305 );
xor \U$26930 ( \27307 , \27280 , \27306 );
xor \U$26931 ( \27308 , \26684 , \26715 );
and \U$26932 ( \27309 , \27308 , \26699 );
and \U$26933 ( \27310 , \26684 , \26715 );
or \U$26934 ( \27311 , \27309 , \27310 );
xor \U$26935 ( \27312 , \27307 , \27311 );
xor \U$26936 ( \27313 , \26727 , \26741 );
and \U$26937 ( \27314 , \27313 , \26757 );
and \U$26938 ( \27315 , \26727 , \26741 );
or \U$26939 ( \27316 , \27314 , \27315 );
and \U$26940 ( \27317 , \27312 , \27316 );
and \U$26941 ( \27318 , \27307 , \27311 );
or \U$26942 ( \27319 , \27317 , \27318 );
xor \U$26943 ( \27320 , \27265 , \27319 );
xor \U$26944 ( \27321 , \26939 , \26988 );
and \U$26945 ( \27322 , \27321 , \27029 );
and \U$26946 ( \27323 , \26939 , \26988 );
or \U$26947 ( \27324 , \27322 , \27323 );
xor \U$26948 ( \27325 , \27320 , \27324 );
xor \U$26949 ( \27326 , \27201 , \27325 );
xor \U$26950 ( \27327 , \27202 , \27207 );
xor \U$26951 ( \27328 , \27327 , \27221 );
not \U$26952 ( \27329 , \2173 );
not \U$26953 ( \27330 , \27271 );
or \U$26954 ( \27331 , \27329 , \27330 );
not \U$26955 ( \27332 , RIc226a70_25);
not \U$26956 ( \27333 , \13223 );
or \U$26957 ( \27334 , \27332 , \27333 );
nand \U$26958 ( \27335 , \10110 , \1905 );
nand \U$26959 ( \27336 , \27334 , \27335 );
nand \U$26960 ( \27337 , \27336 , \2195 );
nand \U$26961 ( \27338 , \27331 , \27337 );
xor \U$26962 ( \27339 , \27328 , \27338 );
not \U$26963 ( \27340 , \2154 );
not \U$26964 ( \27341 , \26952 );
or \U$26965 ( \27342 , \27340 , \27341 );
nand \U$26966 ( \27343 , \26815 , \2138 );
nand \U$26967 ( \27344 , \27342 , \27343 );
xor \U$26968 ( \27345 , \27339 , \27344 );
not \U$26969 ( \27346 , \2367 );
not \U$26970 ( \27347 , \27286 );
or \U$26971 ( \27348 , \27346 , \27347 );
not \U$26972 ( \27349 , RIc226c50_21);
not \U$26973 ( \27350 , \13442 );
or \U$26974 ( \27351 , \27349 , \27350 );
nand \U$26975 ( \27352 , \9324 , \3204 );
nand \U$26976 ( \27353 , \27351 , \27352 );
nand \U$26977 ( \27354 , \27353 , \2392 );
nand \U$26978 ( \27355 , \27348 , \27354 );
not \U$26979 ( \27356 , \1930 );
not \U$26980 ( \27357 , \27241 );
or \U$26981 ( \27358 , \27356 , \27357 );
and \U$26982 ( \27359 , \9274 , \5637 );
not \U$26983 ( \27360 , \9274 );
and \U$26984 ( \27361 , \27360 , RIc226b60_23);
or \U$26985 ( \27362 , \27359 , \27361 );
nand \U$26986 ( \27363 , \27362 , \10214 );
nand \U$26987 ( \27364 , \27358 , \27363 );
xor \U$26988 ( \27365 , \27355 , \27364 );
not \U$26989 ( \27366 , \3631 );
not \U$26990 ( \27367 , \27013 );
or \U$26991 ( \27368 , \27366 , \27367 );
not \U$26992 ( \27369 , RIc2266b0_33);
not \U$26993 ( \27370 , \8830 );
or \U$26994 ( \27371 , \27369 , \27370 );
nand \U$26995 ( \27372 , \20216 , \5179 );
nand \U$26996 ( \27373 , \27371 , \27372 );
nand \U$26997 ( \27374 , \27373 , \3629 );
nand \U$26998 ( \27375 , \27368 , \27374 );
xor \U$26999 ( \27376 , \27365 , \27375 );
xor \U$27000 ( \27377 , \27345 , \27376 );
not \U$27001 ( \27378 , \5135 );
not \U$27002 ( \27379 , RIc2265c0_35);
not \U$27003 ( \27380 , \16531 );
or \U$27004 ( \27381 , \27379 , \27380 );
nand \U$27005 ( \27382 , \8886 , \3620 );
nand \U$27006 ( \27383 , \27381 , \27382 );
not \U$27007 ( \27384 , \27383 );
or \U$27008 ( \27385 , \27378 , \27384 );
not \U$27009 ( \27386 , RIc2265c0_35);
not \U$27010 ( \27387 , \8857 );
or \U$27011 ( \27388 , \27386 , \27387 );
nand \U$27012 ( \27389 , \8856 , \4376 );
nand \U$27013 ( \27390 , \27388 , \27389 );
nand \U$27014 ( \27391 , \27390 , \4381 );
nand \U$27015 ( \27392 , \27385 , \27391 );
not \U$27016 ( \27393 , \16891 );
not \U$27017 ( \27394 , RIc2258a0_63);
not \U$27018 ( \27395 , \3091 );
or \U$27019 ( \27396 , \27394 , \27395 );
nand \U$27020 ( \27397 , \10933 , \16880 );
nand \U$27021 ( \27398 , \27396 , \27397 );
not \U$27022 ( \27399 , \27398 );
or \U$27023 ( \27400 , \27393 , \27399 );
and \U$27024 ( \27401 , \2353 , \16880 );
not \U$27025 ( \27402 , \2353 );
and \U$27026 ( \27403 , \27402 , RIc2258a0_63);
or \U$27027 ( \27404 , \27401 , \27403 );
nand \U$27028 ( \27405 , \27404 , RIc225828_64);
nand \U$27029 ( \27406 , \27400 , \27405 );
or \U$27030 ( \27407 , \27392 , \27406 );
not \U$27031 ( \27408 , \10445 );
not \U$27032 ( \27409 , RIc225f30_49);
not \U$27033 ( \27410 , \4227 );
or \U$27034 ( \27411 , \27409 , \27410 );
nand \U$27035 ( \27412 , \2634 , \11289 );
nand \U$27036 ( \27413 , \27411 , \27412 );
not \U$27037 ( \27414 , \27413 );
or \U$27038 ( \27415 , \27408 , \27414 );
nand \U$27039 ( \27416 , \27044 , \9552 );
nand \U$27040 ( \27417 , \27415 , \27416 );
nand \U$27041 ( \27418 , \27407 , \27417 );
nand \U$27042 ( \27419 , \27406 , \27392 );
nand \U$27043 ( \27420 , \27418 , \27419 );
and \U$27044 ( \27421 , \27377 , \27420 );
and \U$27045 ( \27422 , \27345 , \27376 );
or \U$27046 ( \27423 , \27421 , \27422 );
not \U$27047 ( \27424 , \2318 );
not \U$27048 ( \27425 , \27219 );
or \U$27049 ( \27426 , \27424 , \27425 );
nand \U$27050 ( \27427 , \26783 , \2320 );
nand \U$27051 ( \27428 , \27426 , \27427 );
xor \U$27052 ( \27429 , \27132 , \27145 );
xor \U$27053 ( \27430 , \27428 , \27429 );
not \U$27054 ( \27431 , \2534 );
not \U$27055 ( \27432 , \27165 );
or \U$27056 ( \27433 , \27431 , \27432 );
not \U$27057 ( \27434 , RIc226d40_19);
not \U$27058 ( \27435 , \16492 );
or \U$27059 ( \27436 , \27434 , \27435 );
nand \U$27060 ( \27437 , \3338 , \13497 );
nand \U$27061 ( \27438 , \27436 , \27437 );
nand \U$27062 ( \27439 , \27438 , \2518 );
nand \U$27063 ( \27440 , \27433 , \27439 );
and \U$27064 ( \27441 , \27430 , \27440 );
and \U$27065 ( \27442 , \27428 , \27429 );
or \U$27066 ( \27443 , \27441 , \27442 );
not \U$27067 ( \27444 , \4381 );
not \U$27068 ( \27445 , \27383 );
or \U$27069 ( \27446 , \27444 , \27445 );
nand \U$27070 ( \27447 , \26936 , \4383 );
nand \U$27071 ( \27448 , \27446 , \27447 );
xor \U$27072 ( \27449 , \27443 , \27448 );
not \U$27073 ( \27450 , RIc225828_64);
not \U$27074 ( \27451 , RIc2258a0_63);
not \U$27075 ( \27452 , \4181 );
or \U$27076 ( \27453 , \27451 , \27452 );
nand \U$27077 ( \27454 , \17977 , \16880 );
nand \U$27078 ( \27455 , \27453 , \27454 );
not \U$27079 ( \27456 , \27455 );
or \U$27080 ( \27457 , \27450 , \27456 );
not \U$27081 ( \27458 , RIc2258a0_63);
not \U$27082 ( \27459 , \2347 );
or \U$27083 ( \27460 , \27458 , \27459 );
nand \U$27084 ( \27461 , \2346 , \16880 );
nand \U$27085 ( \27462 , \27460 , \27461 );
nand \U$27086 ( \27463 , \27462 , \16891 );
nand \U$27087 ( \27464 , \27457 , \27463 );
xor \U$27088 ( \27465 , \27449 , \27464 );
not \U$27089 ( \27466 , \11117 );
not \U$27090 ( \27467 , RIc225c60_55);
not \U$27091 ( \27468 , \10896 );
or \U$27092 ( \27469 , \27467 , \27468 );
nand \U$27093 ( \27470 , \3446 , \11108 );
nand \U$27094 ( \27471 , \27469 , \27470 );
not \U$27095 ( \27472 , \27471 );
or \U$27096 ( \27473 , \27466 , \27472 );
nand \U$27097 ( \27474 , \27122 , \13024 );
nand \U$27098 ( \27475 , \27473 , \27474 );
buf \U$27099 ( \27476 , \27475 );
not \U$27100 ( \27477 , \27476 );
not \U$27101 ( \27478 , \15729 );
not \U$27102 ( \27479 , \27089 );
or \U$27103 ( \27480 , \27478 , \27479 );
and \U$27104 ( \27481 , RIc225990_61, \9570 );
not \U$27105 ( \27482 , RIc225990_61);
and \U$27106 ( \27483 , \27482 , \2443 );
or \U$27107 ( \27484 , \27481 , \27483 );
nand \U$27108 ( \27485 , \27484 , \15719 );
nand \U$27109 ( \27486 , \27480 , \27485 );
not \U$27110 ( \27487 , \27486 );
or \U$27111 ( \27488 , \27477 , \27487 );
or \U$27112 ( \27489 , \27486 , \27476 );
not \U$27113 ( \27490 , \8777 );
not \U$27114 ( \27491 , RIc225d50_53);
not \U$27115 ( \27492 , \4195 );
or \U$27116 ( \27493 , \27491 , \27492 );
nand \U$27117 ( \27494 , \2498 , \8772 );
nand \U$27118 ( \27495 , \27493 , \27494 );
not \U$27119 ( \27496 , \27495 );
or \U$27120 ( \27497 , \27490 , \27496 );
nand \U$27121 ( \27498 , \27180 , \9555 );
nand \U$27122 ( \27499 , \27497 , \27498 );
nand \U$27123 ( \27500 , \27489 , \27499 );
nand \U$27124 ( \27501 , \27488 , \27500 );
xor \U$27125 ( \27502 , \27465 , \27501 );
not \U$27126 ( \27503 , \11965 );
and \U$27127 ( \27504 , RIc225b70_57, \9433 );
not \U$27128 ( \27505 , RIc225b70_57);
and \U$27129 ( \27506 , \27505 , \2013 );
or \U$27130 ( \27507 , \27504 , \27506 );
not \U$27131 ( \27508 , \27507 );
or \U$27132 ( \27509 , \27503 , \27508 );
nand \U$27133 ( \27510 , \27058 , \15267 );
nand \U$27134 ( \27511 , \27509 , \27510 );
not \U$27135 ( \27512 , \9398 );
not \U$27136 ( \27513 , \27109 );
or \U$27137 ( \27514 , \27512 , \27513 );
not \U$27138 ( \27515 , RIc226110_45);
not \U$27139 ( \27516 , \9674 );
or \U$27140 ( \27517 , \27515 , \27516 );
nand \U$27141 ( \27518 , \3640 , \9379 );
nand \U$27142 ( \27519 , \27517 , \27518 );
nand \U$27143 ( \27520 , \27519 , \9934 );
nand \U$27144 ( \27521 , \27514 , \27520 );
xor \U$27145 ( \27522 , \27511 , \27521 );
not \U$27146 ( \27523 , \10953 );
not \U$27147 ( \27524 , \27077 );
or \U$27148 ( \27525 , \27523 , \27524 );
not \U$27149 ( \27526 , RIc226020_47);
not \U$27150 ( \27527 , \9513 );
or \U$27151 ( \27528 , \27526 , \27527 );
not \U$27152 ( \27529 , RIc226020_47);
nand \U$27153 ( \27530 , \27529 , \11324 );
nand \U$27154 ( \27531 , \27528 , \27530 );
nand \U$27155 ( \27532 , \27531 , \10001 );
nand \U$27156 ( \27533 , \27525 , \27532 );
and \U$27157 ( \27534 , \27522 , \27533 );
and \U$27158 ( \27535 , \27511 , \27521 );
or \U$27159 ( \27536 , \27534 , \27535 );
and \U$27160 ( \27537 , \27502 , \27536 );
and \U$27161 ( \27538 , \27465 , \27501 );
or \U$27162 ( \27539 , \27537 , \27538 );
xor \U$27163 ( \27540 , \27423 , \27539 );
not \U$27164 ( \27541 , \27063 );
not \U$27165 ( \27542 , \27082 );
or \U$27166 ( \27543 , \27541 , \27542 );
nand \U$27167 ( \27544 , \27543 , \27046 );
not \U$27168 ( \27545 , \27063 );
nand \U$27169 ( \27546 , \27545 , \27079 );
nand \U$27170 ( \27547 , \27544 , \27546 );
buf \U$27171 ( \27548 , \27547 );
xor \U$27172 ( \27549 , \27168 , \27182 );
and \U$27173 ( \27550 , \27549 , \27192 );
and \U$27174 ( \27551 , \27168 , \27182 );
or \U$27175 ( \27552 , \27550 , \27551 );
xor \U$27176 ( \27553 , \27096 , \27111 );
and \U$27177 ( \27554 , \27553 , \27124 );
and \U$27178 ( \27555 , \27096 , \27111 );
or \U$27179 ( \27556 , \27554 , \27555 );
and \U$27180 ( \27557 , \27552 , \27556 );
not \U$27181 ( \27558 , \27552 );
not \U$27182 ( \27559 , \27556 );
and \U$27183 ( \27560 , \27558 , \27559 );
or \U$27184 ( \27561 , \27557 , \27560 );
xor \U$27185 ( \27562 , \27548 , \27561 );
and \U$27186 ( \27563 , \27540 , \27562 );
and \U$27187 ( \27564 , \27423 , \27539 );
or \U$27188 ( \27565 , \27563 , \27564 );
xor \U$27189 ( \27566 , \27326 , \27565 );
not \U$27190 ( \27567 , \27566 );
and \U$27191 ( \27568 , \16248 , \1338 );
not \U$27192 ( \27569 , \1310 );
and \U$27193 ( \27570 , \13487 , \1302 );
not \U$27194 ( \27571 , \13487 );
and \U$27195 ( \27572 , \27571 , RIc227100_11);
or \U$27196 ( \27573 , \27570 , \27572 );
not \U$27197 ( \27574 , \27573 );
or \U$27198 ( \27575 , \27569 , \27574 );
nand \U$27199 ( \27576 , \26872 , \1306 );
nand \U$27200 ( \27577 , \27575 , \27576 );
xor \U$27201 ( \27578 , \27568 , \27577 );
not \U$27202 ( \27579 , \1682 );
not \U$27203 ( \27580 , RIc227010_13);
not \U$27204 ( \27581 , \18167 );
or \U$27205 ( \27582 , \27580 , \27581 );
nand \U$27206 ( \27583 , \12825 , \1758 );
nand \U$27207 ( \27584 , \27582 , \27583 );
not \U$27208 ( \27585 , \27584 );
or \U$27209 ( \27586 , \27579 , \27585 );
nand \U$27210 ( \27587 , \26886 , \1678 );
nand \U$27211 ( \27588 , \27586 , \27587 );
xor \U$27212 ( \27589 , \27578 , \27588 );
not \U$27213 ( \27590 , \1914 );
not \U$27214 ( \27591 , \27248 );
or \U$27215 ( \27592 , \27590 , \27591 );
not \U$27216 ( \27593 , RIc226b60_23);
not \U$27217 ( \27594 , \9076 );
or \U$27218 ( \27595 , \27593 , \27594 );
nand \U$27219 ( \27596 , \9071 , \1911 );
nand \U$27220 ( \27597 , \27595 , \27596 );
nand \U$27221 ( \27598 , \27597 , \1930 );
nand \U$27222 ( \27599 , \27592 , \27598 );
xor \U$27223 ( \27600 , \27589 , \27599 );
not \U$27224 ( \27601 , \2392 );
not \U$27225 ( \27602 , \27293 );
or \U$27226 ( \27603 , \27601 , \27602 );
not \U$27227 ( \27604 , RIc226c50_21);
not \U$27228 ( \27605 , \9255 );
or \U$27229 ( \27606 , \27604 , \27605 );
nand \U$27230 ( \27607 , \10986 , \2383 );
nand \U$27231 ( \27608 , \27606 , \27607 );
nand \U$27232 ( \27609 , \27608 , \2367 );
nand \U$27233 ( \27610 , \27603 , \27609 );
xor \U$27234 ( \27611 , \27600 , \27610 );
not \U$27235 ( \27612 , \2518 );
not \U$27236 ( \27613 , \27301 );
or \U$27237 ( \27614 , \27612 , \27613 );
not \U$27238 ( \27615 , RIc226d40_19);
not \U$27239 ( \27616 , \9297 );
or \U$27240 ( \27617 , \27615 , \27616 );
nand \U$27241 ( \27618 , \9298 , \2523 );
nand \U$27242 ( \27619 , \27617 , \27618 );
nand \U$27243 ( \27620 , \27619 , \2533 );
nand \U$27244 ( \27621 , \27614 , \27620 );
not \U$27245 ( \27622 , \2172 );
not \U$27246 ( \27623 , RIc226a70_25);
not \U$27247 ( \27624 , \11405 );
or \U$27248 ( \27625 , \27623 , \27624 );
nand \U$27249 ( \27626 , \8924 , \2190 );
nand \U$27250 ( \27627 , \27625 , \27626 );
not \U$27251 ( \27628 , \27627 );
or \U$27252 ( \27629 , \27622 , \27628 );
nand \U$27253 ( \27630 , \27278 , \2195 );
nand \U$27254 ( \27631 , \27629 , \27630 );
xor \U$27255 ( \27632 , \27621 , \27631 );
not \U$27256 ( \27633 , \2710 );
and \U$27257 ( \27634 , \8856 , \6902 );
not \U$27258 ( \27635 , \8856 );
and \U$27259 ( \27636 , \27635 , RIc2267a0_31);
or \U$27260 ( \27637 , \27634 , \27636 );
not \U$27261 ( \27638 , \27637 );
or \U$27262 ( \27639 , \27633 , \27638 );
nand \U$27263 ( \27640 , \26960 , \2697 );
nand \U$27264 ( \27641 , \27639 , \27640 );
xor \U$27265 ( \27642 , \27632 , \27641 );
xor \U$27266 ( \27643 , \27611 , \27642 );
xor \U$27267 ( \27644 , \26912 , \26922 );
and \U$27268 ( \27645 , \27644 , \26938 );
and \U$27269 ( \27646 , \26912 , \26922 );
or \U$27270 ( \27647 , \27645 , \27646 );
xor \U$27271 ( \27648 , \27643 , \27647 );
not \U$27272 ( \27649 , \27559 );
not \U$27273 ( \27650 , \27547 );
or \U$27274 ( \27651 , \27649 , \27650 );
not \U$27275 ( \27652 , \27547 );
not \U$27276 ( \27653 , \27652 );
not \U$27277 ( \27654 , \27556 );
or \U$27278 ( \27655 , \27653 , \27654 );
nand \U$27279 ( \27656 , \27655 , \27552 );
nand \U$27280 ( \27657 , \27651 , \27656 );
xor \U$27281 ( \27658 , \27648 , \27657 );
not \U$27282 ( \27659 , \10214 );
not \U$27283 ( \27660 , RIc226b60_23);
not \U$27284 ( \27661 , \10263 );
or \U$27285 ( \27662 , \27660 , \27661 );
nand \U$27286 ( \27663 , \9298 , \1927 );
nand \U$27287 ( \27664 , \27662 , \27663 );
not \U$27288 ( \27665 , \27664 );
or \U$27289 ( \27666 , \27659 , \27665 );
nand \U$27290 ( \27667 , \27362 , \1930 );
nand \U$27291 ( \27668 , \27666 , \27667 );
not \U$27292 ( \27669 , \2367 );
not \U$27293 ( \27670 , \27353 );
or \U$27294 ( \27671 , \27669 , \27670 );
not \U$27295 ( \27672 , RIc226c50_21);
not \U$27296 ( \27673 , \12862 );
or \U$27297 ( \27674 , \27672 , \27673 );
nand \U$27298 ( \27675 , \10086 , \2383 );
nand \U$27299 ( \27676 , \27674 , \27675 );
nand \U$27300 ( \27677 , \27676 , \2391 );
nand \U$27301 ( \27678 , \27671 , \27677 );
xor \U$27302 ( \27679 , \27668 , \27678 );
not \U$27303 ( \27680 , \2195 );
not \U$27304 ( \27681 , RIc226a70_25);
not \U$27305 ( \27682 , \11488 );
or \U$27306 ( \27683 , \27681 , \27682 );
nand \U$27307 ( \27684 , \10986 , \2190 );
nand \U$27308 ( \27685 , \27683 , \27684 );
not \U$27309 ( \27686 , \27685 );
or \U$27310 ( \27687 , \27680 , \27686 );
nand \U$27311 ( \27688 , \27336 , \2173 );
nand \U$27312 ( \27689 , \27687 , \27688 );
and \U$27313 ( \27690 , \27679 , \27689 );
and \U$27314 ( \27691 , \27668 , \27678 );
or \U$27315 ( \27692 , \27690 , \27691 );
not \U$27316 ( \27693 , \27692 );
not \U$27317 ( \27694 , \9444 );
not \U$27318 ( \27695 , RIc225e40_51);
not \U$27319 ( \27696 , \2894 );
or \U$27320 ( \27697 , \27695 , \27696 );
nand \U$27321 ( \27698 , \2500 , \22140 );
nand \U$27322 ( \27699 , \27697 , \27698 );
not \U$27323 ( \27700 , \27699 );
or \U$27324 ( \27701 , \27694 , \27700 );
nand \U$27325 ( \27702 , \26838 , \9459 );
nand \U$27326 ( \27703 , \27701 , \27702 );
not \U$27327 ( \27704 , \27703 );
or \U$27328 ( \27705 , \27693 , \27704 );
or \U$27329 ( \27706 , \27703 , \27692 );
xor \U$27330 ( \27707 , \26776 , \26809 );
and \U$27331 ( \27708 , \27707 , \26824 );
and \U$27332 ( \27709 , \26776 , \26809 );
or \U$27333 ( \27710 , \27708 , \27709 );
nand \U$27334 ( \27711 , \27706 , \27710 );
nand \U$27335 ( \27712 , \27705 , \27711 );
not \U$27336 ( \27713 , \9129 );
not \U$27337 ( \27714 , RIc226200_43);
not \U$27338 ( \27715 , \17703 );
or \U$27339 ( \27716 , \27714 , \27715 );
nand \U$27340 ( \27717 , \2980 , \9106 );
nand \U$27341 ( \27718 , \27716 , \27717 );
not \U$27342 ( \27719 , \27718 );
or \U$27343 ( \27720 , \27713 , \27719 );
nand \U$27344 ( \27721 , \26748 , \9110 );
nand \U$27345 ( \27722 , \27720 , \27721 );
not \U$27346 ( \27723 , \11118 );
not \U$27347 ( \27724 , \27117 );
or \U$27348 ( \27725 , \27723 , \27724 );
not \U$27349 ( \27726 , RIc225c60_55);
not \U$27350 ( \27727 , \9408 );
or \U$27351 ( \27728 , \27726 , \27727 );
nand \U$27352 ( \27729 , \3834 , \16788 );
nand \U$27353 ( \27730 , \27728 , \27729 );
nand \U$27354 ( \27731 , \27730 , \12532 );
nand \U$27355 ( \27732 , \27725 , \27731 );
xor \U$27356 ( \27733 , \27722 , \27732 );
not \U$27357 ( \27734 , \11577 );
not \U$27358 ( \27735 , RIc225d50_53);
not \U$27359 ( \27736 , \2586 );
or \U$27360 ( \27737 , \27735 , \27736 );
nand \U$27361 ( \27738 , \3183 , \8782 );
nand \U$27362 ( \27739 , \27737 , \27738 );
not \U$27363 ( \27740 , \27739 );
or \U$27364 ( \27741 , \27734 , \27740 );
nand \U$27365 ( \27742 , \27173 , \9488 );
nand \U$27366 ( \27743 , \27741 , \27742 );
xor \U$27367 ( \27744 , \27733 , \27743 );
xor \U$27368 ( \27745 , \27712 , \27744 );
not \U$27369 ( \27746 , \9458 );
not \U$27370 ( \27747 , \27699 );
or \U$27371 ( \27748 , \27746 , \27747 );
not \U$27372 ( \27749 , RIc225e40_51);
not \U$27373 ( \27750 , \5819 );
or \U$27374 ( \27751 , \27749 , \27750 );
nand \U$27375 ( \27752 , \2480 , \11795 );
nand \U$27376 ( \27753 , \27751 , \27752 );
nand \U$27377 ( \27754 , \27753 , \11708 );
nand \U$27378 ( \27755 , \27748 , \27754 );
not \U$27379 ( \27756 , \15164 );
not \U$27380 ( \27757 , \27190 );
or \U$27381 ( \27758 , \27756 , \27757 );
and \U$27382 ( \27759 , RIc225a80_59, \3686 );
not \U$27383 ( \27760 , RIc225a80_59);
not \U$27384 ( \27761 , \13914 );
and \U$27385 ( \27762 , \27760 , \27761 );
or \U$27386 ( \27763 , \27759 , \27762 );
nand \U$27387 ( \27764 , \27763 , \12670 );
nand \U$27388 ( \27765 , \27758 , \27764 );
not \U$27389 ( \27766 , \27765 );
and \U$27390 ( \27767 , \27755 , \27766 );
not \U$27391 ( \27768 , \27755 );
and \U$27392 ( \27769 , \27768 , \27765 );
or \U$27393 ( \27770 , \27767 , \27769 );
not \U$27394 ( \27771 , \20159 );
not \U$27395 ( \27772 , \27455 );
or \U$27396 ( \27773 , \27771 , \27772 );
not \U$27397 ( \27774 , RIc2258a0_63);
not \U$27398 ( \27775 , \3783 );
or \U$27399 ( \27776 , \27774 , \27775 );
nand \U$27400 ( \27777 , \3043 , \16880 );
nand \U$27401 ( \27778 , \27776 , \27777 );
nand \U$27402 ( \27779 , \27778 , RIc225828_64);
nand \U$27403 ( \27780 , \27773 , \27779 );
and \U$27404 ( \27781 , \27770 , \27780 );
not \U$27405 ( \27782 , \27770 );
not \U$27406 ( \27783 , \27780 );
and \U$27407 ( \27784 , \27782 , \27783 );
nor \U$27408 ( \27785 , \27781 , \27784 );
and \U$27409 ( \27786 , \27745 , \27785 );
and \U$27410 ( \27787 , \27712 , \27744 );
or \U$27411 ( \27788 , \27786 , \27787 );
xor \U$27412 ( \27789 , \27658 , \27788 );
xor \U$27413 ( \27790 , \26880 , \26895 );
and \U$27414 ( \27791 , \27790 , \26911 );
and \U$27415 ( \27792 , \26880 , \26895 );
or \U$27416 ( \27793 , \27791 , \27792 );
not \U$27417 ( \27794 , \5135 );
not \U$27418 ( \27795 , RIc2265c0_35);
not \U$27419 ( \27796 , \6493 );
or \U$27420 ( \27797 , \27795 , \27796 );
buf \U$27421 ( \27798 , \6492 );
nand \U$27422 ( \27799 , \27798 , \3620 );
nand \U$27423 ( \27800 , \27797 , \27799 );
not \U$27424 ( \27801 , \27800 );
or \U$27425 ( \27802 , \27794 , \27801 );
nand \U$27426 ( \27803 , \26930 , \5741 );
nand \U$27427 ( \27804 , \27802 , \27803 );
xor \U$27428 ( \27805 , \27793 , \27804 );
not \U$27429 ( \27806 , \15719 );
not \U$27430 ( \27807 , RIc225990_61);
not \U$27431 ( \27808 , \12382 );
or \U$27432 ( \27809 , \27807 , \27808 );
nand \U$27433 ( \27810 , \2353 , \10338 );
nand \U$27434 ( \27811 , \27809 , \27810 );
not \U$27435 ( \27812 , \27811 );
or \U$27436 ( \27813 , \27806 , \27812 );
not \U$27437 ( \27814 , RIc225990_61);
not \U$27438 ( \27815 , \4181 );
or \U$27439 ( \27816 , \27814 , \27815 );
nand \U$27440 ( \27817 , \9196 , \12806 );
nand \U$27441 ( \27818 , \27816 , \27817 );
nand \U$27442 ( \27819 , \27818 , \15729 );
nand \U$27443 ( \27820 , \27813 , \27819 );
xor \U$27444 ( \27821 , \27805 , \27820 );
not \U$27445 ( \27822 , \5519 );
not \U$27446 ( \27823 , RIc2264d0_37);
not \U$27447 ( \27824 , \15603 );
or \U$27448 ( \27825 , \27823 , \27824 );
nand \U$27449 ( \27826 , \20655 , \5504 );
nand \U$27450 ( \27827 , \27825 , \27826 );
not \U$27451 ( \27828 , \27827 );
or \U$27452 ( \27829 , \27822 , \27828 );
nand \U$27453 ( \27830 , \26918 , \5509 );
nand \U$27454 ( \27831 , \27829 , \27830 );
not \U$27455 ( \27832 , \6307 );
not \U$27456 ( \27833 , RIc2263e0_39);
not \U$27457 ( \27834 , \10220 );
or \U$27458 ( \27835 , \27833 , \27834 );
nand \U$27459 ( \27836 , \4407 , \25483 );
nand \U$27460 ( \27837 , \27835 , \27836 );
not \U$27461 ( \27838 , \27837 );
or \U$27462 ( \27839 , \27832 , \27838 );
nand \U$27463 ( \27840 , \27026 , \6689 );
nand \U$27464 ( \27841 , \27839 , \27840 );
xor \U$27465 ( \27842 , \27831 , \27841 );
not \U$27466 ( \27843 , \9705 );
not \U$27467 ( \27844 , RIc2262f0_41);
not \U$27468 ( \27845 , \4049 );
or \U$27469 ( \27846 , \27844 , \27845 );
nand \U$27470 ( \27847 , \15768 , \6303 );
nand \U$27471 ( \27848 , \27846 , \27847 );
not \U$27472 ( \27849 , \27848 );
or \U$27473 ( \27850 , \27843 , \27849 );
nand \U$27474 ( \27851 , \26998 , \9690 );
nand \U$27475 ( \27852 , \27850 , \27851 );
xor \U$27476 ( \27853 , \27842 , \27852 );
xor \U$27477 ( \27854 , \27821 , \27853 );
not \U$27478 ( \27855 , \27780 );
not \U$27479 ( \27856 , \27765 );
or \U$27480 ( \27857 , \27855 , \27856 );
not \U$27481 ( \27858 , \27766 );
not \U$27482 ( \27859 , \27783 );
or \U$27483 ( \27860 , \27858 , \27859 );
nand \U$27484 ( \27861 , \27860 , \27755 );
nand \U$27485 ( \27862 , \27857 , \27861 );
xor \U$27486 ( \27863 , \27854 , \27862 );
xor \U$27487 ( \27864 , \27443 , \27448 );
and \U$27488 ( \27865 , \27864 , \27464 );
and \U$27489 ( \27866 , \27443 , \27448 );
or \U$27490 ( \27867 , \27865 , \27866 );
xor \U$27491 ( \27868 , \27146 , \27151 );
and \U$27492 ( \27869 , \27868 , \27167 );
and \U$27493 ( \27870 , \27146 , \27151 );
or \U$27494 ( \27871 , \27869 , \27870 );
not \U$27495 ( \27872 , \20862 );
not \U$27496 ( \27873 , \27811 );
or \U$27497 ( \27874 , \27872 , \27873 );
nand \U$27498 ( \27875 , \27094 , \15719 );
nand \U$27499 ( \27876 , \27874 , \27875 );
xor \U$27500 ( \27877 , \27871 , \27876 );
not \U$27501 ( \27878 , \10445 );
not \U$27502 ( \27879 , \27037 );
or \U$27503 ( \27880 , \27878 , \27879 );
not \U$27504 ( \27881 , RIc225f30_49);
not \U$27505 ( \27882 , \2670 );
or \U$27506 ( \27883 , \27881 , \27882 );
nand \U$27507 ( \27884 , \17831 , \9549 );
nand \U$27508 ( \27885 , \27883 , \27884 );
nand \U$27509 ( \27886 , \27885 , \9552 );
nand \U$27510 ( \27887 , \27880 , \27886 );
xor \U$27511 ( \27888 , \27877 , \27887 );
xor \U$27512 ( \27889 , \27867 , \27888 );
not \U$27513 ( \27890 , \9619 );
not \U$27514 ( \27891 , RIc226020_47);
not \U$27515 ( \27892 , \11068 );
or \U$27516 ( \27893 , \27891 , \27892 );
nand \U$27517 ( \27894 , \11515 , \9373 );
nand \U$27518 ( \27895 , \27893 , \27894 );
not \U$27519 ( \27896 , \27895 );
or \U$27520 ( \27897 , \27890 , \27896 );
nand \U$27521 ( \27898 , \27071 , \10001 );
nand \U$27522 ( \27899 , \27897 , \27898 );
not \U$27523 ( \27900 , \11965 );
not \U$27524 ( \27901 , \27051 );
or \U$27525 ( \27902 , \27900 , \27901 );
not \U$27526 ( \27903 , RIc225b70_57);
not \U$27527 ( \27904 , \2233 );
or \U$27528 ( \27905 , \27903 , \27904 );
not \U$27529 ( \27906 , \9599 );
nand \U$27530 ( \27907 , \27906 , \15262 );
nand \U$27531 ( \27908 , \27905 , \27907 );
nand \U$27532 ( \27909 , \27908 , \11974 );
nand \U$27533 ( \27910 , \27902 , \27909 );
not \U$27534 ( \27911 , \27910 );
and \U$27535 ( \27912 , \27899 , \27911 );
not \U$27536 ( \27913 , \27899 );
and \U$27537 ( \27914 , \27913 , \27910 );
or \U$27538 ( \27915 , \27912 , \27914 );
not \U$27539 ( \27916 , \4500 );
not \U$27540 ( \27917 , \9100 );
and \U$27541 ( \27918 , \27916 , \27917 );
and \U$27542 ( \27919 , \15217 , \9100 );
nor \U$27543 ( \27920 , \27918 , \27919 );
not \U$27544 ( \27921 , \27920 );
not \U$27545 ( \27922 , \23212 );
and \U$27546 ( \27923 , \27921 , \27922 );
not \U$27547 ( \27924 , \27101 );
and \U$27548 ( \27925 , \27924 , \9934 );
nor \U$27549 ( \27926 , \27923 , \27925 );
buf \U$27550 ( \27927 , \27926 );
xnor \U$27551 ( \27928 , \27915 , \27927 );
and \U$27552 ( \27929 , \27889 , \27928 );
and \U$27553 ( \27930 , \27867 , \27888 );
or \U$27554 ( \27931 , \27929 , \27930 );
xor \U$27555 ( \27932 , \27863 , \27931 );
nand \U$27556 ( \27933 , \27911 , \27926 );
and \U$27557 ( \27934 , \27933 , \27899 );
nor \U$27558 ( \27935 , \27911 , \27926 );
nor \U$27559 ( \27936 , \27934 , \27935 );
not \U$27560 ( \27937 , \27936 );
xor \U$27561 ( \27938 , \27871 , \27876 );
and \U$27562 ( \27939 , \27938 , \27887 );
and \U$27563 ( \27940 , \27871 , \27876 );
or \U$27564 ( \27941 , \27939 , \27940 );
xor \U$27565 ( \27942 , \27937 , \27941 );
not \U$27566 ( \27943 , \27743 );
not \U$27567 ( \27944 , \27722 );
nand \U$27568 ( \27945 , \27943 , \27944 );
and \U$27569 ( \27946 , \27945 , \27732 );
not \U$27570 ( \27947 , \27743 );
nor \U$27571 ( \27948 , \27947 , \27944 );
nor \U$27572 ( \27949 , \27946 , \27948 );
not \U$27573 ( \27950 , \27949 );
xor \U$27574 ( \27951 , \27942 , \27950 );
xor \U$27575 ( \27952 , \27932 , \27951 );
xor \U$27576 ( \27953 , \27789 , \27952 );
xor \U$27577 ( \27954 , \27867 , \27888 );
xor \U$27578 ( \27955 , \27954 , \27928 );
xor \U$27579 ( \27956 , \27712 , \27744 );
xor \U$27580 ( \27957 , \27956 , \27785 );
xor \U$27581 ( \27958 , \27955 , \27957 );
xor \U$27582 ( \27959 , \27428 , \27429 );
xor \U$27583 ( \27960 , \27959 , \27440 );
or \U$27584 ( \27961 , RIc226ea8_16, RIc226e30_17);
nand \U$27585 ( \27962 , \27961 , \16248 );
and \U$27586 ( \27963 , RIc226ea8_16, RIc226e30_17);
nor \U$27587 ( \27964 , \27963 , \1674 );
and \U$27588 ( \27965 , \27962 , \27964 );
not \U$27589 ( \27966 , \2318 );
not \U$27590 ( \27967 , \26790 );
or \U$27591 ( \27968 , \27966 , \27967 );
or \U$27592 ( \27969 , \18357 , \2351 );
or \U$27593 ( \27970 , \18356 , RIc226f20_15);
nand \U$27594 ( \27971 , \27969 , \27970 );
nand \U$27595 ( \27972 , \27971 , \2319 );
nand \U$27596 ( \27973 , \27968 , \27972 );
and \U$27597 ( \27974 , \27965 , \27973 );
not \U$27598 ( \27975 , \2518 );
not \U$27599 ( \27976 , RIc226d40_19);
not \U$27600 ( \27977 , \13198 );
or \U$27601 ( \27978 , \27976 , \27977 );
nand \U$27602 ( \27979 , \12755 , \1941 );
nand \U$27603 ( \27980 , \27978 , \27979 );
not \U$27604 ( \27981 , \27980 );
or \U$27605 ( \27982 , \27975 , \27981 );
nand \U$27606 ( \27983 , \27438 , \2533 );
nand \U$27607 ( \27984 , \27982 , \27983 );
xor \U$27608 ( \27985 , \27974 , \27984 );
not \U$27609 ( \27986 , \2367 );
not \U$27610 ( \27987 , \27676 );
or \U$27611 ( \27988 , \27986 , \27987 );
not \U$27612 ( \27989 , RIc226c50_21);
not \U$27613 ( \27990 , \10370 );
not \U$27614 ( \27991 , \27990 );
or \U$27615 ( \27992 , \27989 , \27991 );
nand \U$27616 ( \27993 , \21976 , \3204 );
nand \U$27617 ( \27994 , \27992 , \27993 );
nand \U$27618 ( \27995 , \27994 , \2391 );
nand \U$27619 ( \27996 , \27988 , \27995 );
and \U$27620 ( \27997 , \27985 , \27996 );
and \U$27621 ( \27998 , \27974 , \27984 );
or \U$27622 ( \27999 , \27997 , \27998 );
xor \U$27623 ( \28000 , \27960 , \27999 );
not \U$27624 ( \28001 , \5509 );
and \U$27625 ( \28002 , \9728 , RIc2264d0_37);
not \U$27626 ( \28003 , \9728 );
and \U$27627 ( \28004 , \28003 , \4371 );
or \U$27628 ( \28005 , \28002 , \28004 );
not \U$27629 ( \28006 , \28005 );
or \U$27630 ( \28007 , \28001 , \28006 );
nand \U$27631 ( \28008 , \26678 , \5519 );
nand \U$27632 ( \28009 , \28007 , \28008 );
and \U$27633 ( \28010 , \28000 , \28009 );
and \U$27634 ( \28011 , \27960 , \27999 );
or \U$27635 ( \28012 , \28010 , \28011 );
not \U$27636 ( \28013 , \2710 );
not \U$27637 ( \28014 , \26719 );
or \U$27638 ( \28015 , \28013 , \28014 );
not \U$27639 ( \28016 , RIc2267a0_31);
not \U$27640 ( \28017 , \8978 );
or \U$27641 ( \28018 , \28016 , \28017 );
nand \U$27642 ( \28019 , \8979 , \2705 );
nand \U$27643 ( \28020 , \28018 , \28019 );
nand \U$27644 ( \28021 , \28020 , \2697 );
nand \U$27645 ( \28022 , \28015 , \28021 );
not \U$27646 ( \28023 , \2086 );
not \U$27647 ( \28024 , \26732 );
or \U$27648 ( \28025 , \28023 , \28024 );
not \U$27649 ( \28026 , \8924 );
and \U$27650 ( \28027 , RIc226890_29, \28026 );
not \U$27651 ( \28028 , RIc226890_29);
and \U$27652 ( \28029 , \28028 , \8924 );
or \U$27653 ( \28030 , \28027 , \28029 );
nand \U$27654 ( \28031 , \28030 , \2784 );
nand \U$27655 ( \28032 , \28025 , \28031 );
xor \U$27656 ( \28033 , \28022 , \28032 );
not \U$27657 ( \28034 , \3629 );
not \U$27658 ( \28035 , RIc2266b0_33);
not \U$27659 ( \28036 , \8810 );
or \U$27660 ( \28037 , \28035 , \28036 );
nand \U$27661 ( \28038 , \8806 , \6890 );
nand \U$27662 ( \28039 , \28037 , \28038 );
not \U$27663 ( \28040 , \28039 );
or \U$27664 ( \28041 , \28034 , \28040 );
nand \U$27665 ( \28042 , \27373 , \3631 );
nand \U$27666 ( \28043 , \28041 , \28042 );
and \U$27667 ( \28044 , \28033 , \28043 );
and \U$27668 ( \28045 , \28022 , \28032 );
or \U$27669 ( \28046 , \28044 , \28045 );
xor \U$27670 ( \28047 , \28012 , \28046 );
not \U$27671 ( \28048 , \6307 );
not \U$27672 ( \28049 , \26690 );
or \U$27673 ( \28050 , \28048 , \28049 );
and \U$27674 ( \28051 , \9573 , \9775 );
not \U$27675 ( \28052 , \9573 );
and \U$27676 ( \28053 , \28052 , \6492 );
nor \U$27677 ( \28054 , \28051 , \28053 );
nand \U$27678 ( \28055 , \28054 , \6688 );
nand \U$27679 ( \28056 , \28050 , \28055 );
not \U$27680 ( \28057 , \9129 );
not \U$27681 ( \28058 , \26755 );
or \U$27682 ( \28059 , \28057 , \28058 );
not \U$27683 ( \28060 , RIc226200_43);
not \U$27684 ( \28061 , \10277 );
or \U$27685 ( \28062 , \28060 , \28061 );
nand \U$27686 ( \28063 , \4406 , \13805 );
nand \U$27687 ( \28064 , \28062 , \28063 );
nand \U$27688 ( \28065 , \28064 , \9110 );
nand \U$27689 ( \28066 , \28059 , \28065 );
xor \U$27690 ( \28067 , \28056 , \28066 );
not \U$27691 ( \28068 , \9816 );
not \U$27692 ( \28069 , \26706 );
or \U$27693 ( \28070 , \28068 , \28069 );
not \U$27694 ( \28071 , RIc2262f0_41);
not \U$27695 ( \28072 , \15603 );
or \U$27696 ( \28073 , \28071 , \28072 );
nand \U$27697 ( \28074 , \12791 , \9822 );
nand \U$27698 ( \28075 , \28073 , \28074 );
nand \U$27699 ( \28076 , \28075 , \9690 );
nand \U$27700 ( \28077 , \28070 , \28076 );
and \U$27701 ( \28078 , \28067 , \28077 );
and \U$27702 ( \28079 , \28056 , \28066 );
or \U$27703 ( \28080 , \28078 , \28079 );
xor \U$27704 ( \28081 , \28047 , \28080 );
xor \U$27705 ( \28082 , \27668 , \27678 );
xor \U$27706 ( \28083 , \28082 , \27689 );
not \U$27707 ( \28084 , \28083 );
not \U$27708 ( \28085 , \2195 );
not \U$27709 ( \28086 , RIc226a70_25);
not \U$27710 ( \28087 , \10800 );
or \U$27711 ( \28088 , \28086 , \28087 );
nand \U$27712 ( \28089 , \9275 , \9662 );
nand \U$27713 ( \28090 , \28088 , \28089 );
not \U$27714 ( \28091 , \28090 );
or \U$27715 ( \28092 , \28085 , \28091 );
nand \U$27716 ( \28093 , \27685 , \2172 );
nand \U$27717 ( \28094 , \28092 , \28093 );
not \U$27718 ( \28095 , \2138 );
not \U$27719 ( \28096 , RIc226980_27);
not \U$27720 ( \28097 , \13223 );
or \U$27721 ( \28098 , \28096 , \28097 );
nand \U$27722 ( \28099 , \10110 , \2799 );
nand \U$27723 ( \28100 , \28098 , \28099 );
not \U$27724 ( \28101 , \28100 );
or \U$27725 ( \28102 , \28095 , \28101 );
nand \U$27726 ( \28103 , \26822 , \2154 );
nand \U$27727 ( \28104 , \28102 , \28103 );
xor \U$27728 ( \28105 , \28094 , \28104 );
not \U$27729 ( \28106 , \9398 );
not \U$27730 ( \28107 , \27519 );
or \U$27731 ( \28108 , \28106 , \28107 );
not \U$27732 ( \28109 , RIc226110_45);
not \U$27733 ( \28110 , \4122 );
or \U$27734 ( \28111 , \28109 , \28110 );
nand \U$27735 ( \28112 , \4121 , \9379 );
nand \U$27736 ( \28113 , \28111 , \28112 );
nand \U$27737 ( \28114 , \28113 , \9382 );
nand \U$27738 ( \28115 , \28108 , \28114 );
and \U$27739 ( \28116 , \28105 , \28115 );
and \U$27740 ( \28117 , \28094 , \28104 );
or \U$27741 ( \28118 , \28116 , \28117 );
not \U$27742 ( \28119 , \28118 );
nand \U$27743 ( \28120 , \28084 , \28119 );
not \U$27744 ( \28121 , \28120 );
xor \U$27745 ( \28122 , \27965 , \27973 );
not \U$27746 ( \28123 , \1963 );
not \U$27747 ( \28124 , \26801 );
or \U$27748 ( \28125 , \28123 , \28124 );
not \U$27749 ( \28126 , RIc226e30_17);
not \U$27750 ( \28127 , \20392 );
or \U$27751 ( \28128 , \28126 , \28127 );
nand \U$27752 ( \28129 , \13487 , \1960 );
nand \U$27753 ( \28130 , \28128 , \28129 );
nand \U$27754 ( \28131 , \28130 , \1945 );
nand \U$27755 ( \28132 , \28125 , \28131 );
xor \U$27756 ( \28133 , \28122 , \28132 );
not \U$27757 ( \28134 , \2533 );
not \U$27758 ( \28135 , \27980 );
or \U$27759 ( \28136 , \28134 , \28135 );
not \U$27760 ( \28137 , RIc226d40_19);
not \U$27761 ( \28138 , \15444 );
or \U$27762 ( \28139 , \28137 , \28138 );
nand \U$27763 ( \28140 , \12825 , \1941 );
nand \U$27764 ( \28141 , \28139 , \28140 );
nand \U$27765 ( \28142 , \28141 , \2518 );
nand \U$27766 ( \28143 , \28136 , \28142 );
and \U$27767 ( \28144 , \28133 , \28143 );
and \U$27768 ( \28145 , \28122 , \28132 );
or \U$27769 ( \28146 , \28144 , \28145 );
not \U$27770 ( \28147 , \4381 );
not \U$27771 ( \28148 , RIc2265c0_35);
buf \U$27772 ( \28149 , \9900 );
not \U$27773 ( \28150 , \28149 );
or \U$27774 ( \28151 , \28148 , \28150 );
nand \U$27775 ( \28152 , \22969 , \3620 );
nand \U$27776 ( \28153 , \28151 , \28152 );
not \U$27777 ( \28154 , \28153 );
or \U$27778 ( \28155 , \28147 , \28154 );
nand \U$27779 ( \28156 , \27390 , \4383 );
nand \U$27780 ( \28157 , \28155 , \28156 );
xor \U$27781 ( \28158 , \28146 , \28157 );
not \U$27782 ( \28159 , \9534 );
not \U$27783 ( \28160 , RIc225f30_49);
not \U$27784 ( \28161 , \2104 );
or \U$27785 ( \28162 , \28160 , \28161 );
not \U$27786 ( \28163 , RIc225f30_49);
nand \U$27787 ( \28164 , \4500 , \28163 );
nand \U$27788 ( \28165 , \28162 , \28164 );
not \U$27789 ( \28166 , \28165 );
or \U$27790 ( \28167 , \28159 , \28166 );
nand \U$27791 ( \28168 , \27413 , \9552 );
nand \U$27792 ( \28169 , \28167 , \28168 );
and \U$27793 ( \28170 , \28158 , \28169 );
and \U$27794 ( \28171 , \28146 , \28157 );
or \U$27795 ( \28172 , \28170 , \28171 );
not \U$27796 ( \28173 , \28172 );
or \U$27797 ( \28174 , \28121 , \28173 );
nand \U$27798 ( \28175 , \28118 , \28083 );
nand \U$27799 ( \28176 , \28174 , \28175 );
xor \U$27800 ( \28177 , \28081 , \28176 );
xor \U$27801 ( \28178 , \27345 , \27376 );
xor \U$27802 ( \28179 , \28178 , \27420 );
and \U$27803 ( \28180 , \28177 , \28179 );
and \U$27804 ( \28181 , \28081 , \28176 );
or \U$27805 ( \28182 , \28180 , \28181 );
and \U$27806 ( \28183 , \27958 , \28182 );
and \U$27807 ( \28184 , \27955 , \27957 );
or \U$27808 ( \28185 , \28183 , \28184 );
xor \U$27809 ( \28186 , \27953 , \28185 );
not \U$27810 ( \28187 , \28186 );
or \U$27811 ( \28188 , \27567 , \28187 );
or \U$27812 ( \28189 , \27566 , \28186 );
not \U$27813 ( \28190 , \2086 );
not \U$27814 ( \28191 , \28030 );
or \U$27815 ( \28192 , \28190 , \28191 );
and \U$27816 ( \28193 , RIc226890_29, \9049 );
not \U$27817 ( \28194 , RIc226890_29);
and \U$27818 ( \28195 , \28194 , \10644 );
or \U$27819 ( \28196 , \28193 , \28195 );
nand \U$27820 ( \28197 , \28196 , \2078 );
nand \U$27821 ( \28198 , \28192 , \28197 );
not \U$27822 ( \28199 , \28198 );
not \U$27823 ( \28200 , RIc226b60_23);
not \U$27824 ( \28201 , \9321 );
or \U$27825 ( \28202 , \28200 , \28201 );
nand \U$27826 ( \28203 , \9320 , \5637 );
nand \U$27827 ( \28204 , \28202 , \28203 );
not \U$27828 ( \28205 , \28204 );
not \U$27829 ( \28206 , \1914 );
or \U$27830 ( \28207 , \28205 , \28206 );
nand \U$27831 ( \28208 , \27664 , \1930 );
nand \U$27832 ( \28209 , \28207 , \28208 );
not \U$27833 ( \28210 , \28209 );
and \U$27834 ( \28211 , \28199 , \28210 );
xor \U$27835 ( \28212 , \26793 , \26777 );
xor \U$27836 ( \28213 , \28212 , \26805 );
nor \U$27837 ( \28214 , \28211 , \28213 );
and \U$27838 ( \28215 , \28198 , \28209 );
nor \U$27839 ( \28216 , \28214 , \28215 );
not \U$27840 ( \28217 , \6688 );
and \U$27841 ( \28218 , RIc2263e0_39, \6718 );
not \U$27842 ( \28219 , RIc2263e0_39);
and \U$27843 ( \28220 , \28219 , \18410 );
nor \U$27844 ( \28221 , \28218 , \28220 );
not \U$27845 ( \28222 , \28221 );
or \U$27846 ( \28223 , \28217 , \28222 );
nand \U$27847 ( \28224 , \28054 , \6307 );
nand \U$27848 ( \28225 , \28223 , \28224 );
not \U$27849 ( \28226 , \28225 );
not \U$27850 ( \28227 , \5509 );
not \U$27851 ( \28228 , RIc2264d0_37);
not \U$27852 ( \28229 , \12228 );
or \U$27853 ( \28230 , \28228 , \28229 );
not \U$27854 ( \28231 , RIc2264d0_37);
nand \U$27855 ( \28232 , \28231 , \8885 );
nand \U$27856 ( \28233 , \28230 , \28232 );
not \U$27857 ( \28234 , \28233 );
or \U$27858 ( \28235 , \28227 , \28234 );
nand \U$27859 ( \28236 , \28005 , \5519 );
nand \U$27860 ( \28237 , \28235 , \28236 );
not \U$27861 ( \28238 , \28237 );
nand \U$27862 ( \28239 , \28226 , \28238 );
not \U$27863 ( \28240 , \28239 );
not \U$27864 ( \28241 , \9690 );
not \U$27865 ( \28242 , RIc2262f0_41);
not \U$27866 ( \28243 , \17549 );
or \U$27867 ( \28244 , \28242 , \28243 );
nand \U$27868 ( \28245 , \14998 , \12937 );
nand \U$27869 ( \28246 , \28244 , \28245 );
not \U$27870 ( \28247 , \28246 );
or \U$27871 ( \28248 , \28241 , \28247 );
nand \U$27872 ( \28249 , \28075 , \9816 );
nand \U$27873 ( \28250 , \28248 , \28249 );
not \U$27874 ( \28251 , \28250 );
or \U$27875 ( \28252 , \28240 , \28251 );
nand \U$27876 ( \28253 , \28225 , \28237 );
nand \U$27877 ( \28254 , \28252 , \28253 );
not \U$27878 ( \28255 , \28254 );
xor \U$27879 ( \28256 , \28216 , \28255 );
not \U$27880 ( \28257 , RIc226200_43);
not \U$27881 ( \28258 , \9850 );
or \U$27882 ( \28259 , \28257 , \28258 );
nand \U$27883 ( \28260 , \5215 , \9117 );
nand \U$27884 ( \28261 , \28259 , \28260 );
and \U$27885 ( \28262 , \9110 , \28261 );
and \U$27886 ( \28263 , \28064 , \9205 );
nor \U$27887 ( \28264 , \28262 , \28263 );
not \U$27888 ( \28265 , \28020 );
not \U$27889 ( \28266 , \28265 );
not \U$27890 ( \28267 , \18740 );
and \U$27891 ( \28268 , \28266 , \28267 );
and \U$27892 ( \28269 , \8910 , RIc2267a0_31);
not \U$27893 ( \28270 , \8910 );
and \U$27894 ( \28271 , \28270 , \2705 );
or \U$27895 ( \28272 , \28269 , \28271 );
and \U$27896 ( \28273 , \28272 , \2697 );
nor \U$27897 ( \28274 , \28268 , \28273 );
nand \U$27898 ( \28275 , \28264 , \28274 );
not \U$27899 ( \28276 , \3631 );
not \U$27900 ( \28277 , \28039 );
or \U$27901 ( \28278 , \28276 , \28277 );
not \U$27902 ( \28279 , RIc2266b0_33);
not \U$27903 ( \28280 , \9915 );
or \U$27904 ( \28281 , \28279 , \28280 );
nand \U$27905 ( \28282 , \8951 , \5179 );
nand \U$27906 ( \28283 , \28281 , \28282 );
nand \U$27907 ( \28284 , \28283 , \3629 );
nand \U$27908 ( \28285 , \28278 , \28284 );
and \U$27909 ( \28286 , \28275 , \28285 );
nor \U$27910 ( \28287 , \28264 , \28274 );
nor \U$27911 ( \28288 , \28286 , \28287 );
and \U$27912 ( \28289 , \28256 , \28288 );
and \U$27913 ( \28290 , \28216 , \28255 );
or \U$27914 ( \28291 , \28289 , \28290 );
xor \U$27915 ( \28292 , \27710 , \27692 );
xnor \U$27916 ( \28293 , \28292 , \27703 );
and \U$27917 ( \28294 , \28291 , \28293 );
not \U$27918 ( \28295 , \28291 );
not \U$27919 ( \28296 , \28293 );
and \U$27920 ( \28297 , \28295 , \28296 );
nor \U$27921 ( \28298 , \28294 , \28297 );
not \U$27922 ( \28299 , \28298 );
not \U$27923 ( \28300 , \28299 );
not \U$27924 ( \28301 , \12670 );
not \U$27925 ( \28302 , \26846 );
or \U$27926 ( \28303 , \28301 , \28302 );
not \U$27927 ( \28304 , RIc225a80_59);
not \U$27928 ( \28305 , \12508 );
or \U$27929 ( \28306 , \28304 , \28305 );
not \U$27930 ( \28307 , RIc225a80_59);
nand \U$27931 ( \28308 , \28307 , \1988 );
nand \U$27932 ( \28309 , \28306 , \28308 );
nand \U$27933 ( \28310 , \28309 , \15164 );
nand \U$27934 ( \28311 , \28303 , \28310 );
not \U$27935 ( \28312 , \28311 );
not \U$27936 ( \28313 , \11708 );
not \U$27937 ( \28314 , \26831 );
or \U$27938 ( \28315 , \28313 , \28314 );
not \U$27939 ( \28316 , RIc225e40_51);
not \U$27940 ( \28317 , \5526 );
or \U$27941 ( \28318 , \28316 , \28317 );
nand \U$27942 ( \28319 , \2042 , \9450 );
nand \U$27943 ( \28320 , \28318 , \28319 );
nand \U$27944 ( \28321 , \28320 , \9459 );
nand \U$27945 ( \28322 , \28315 , \28321 );
not \U$27946 ( \28323 , \28322 );
nand \U$27947 ( \28324 , \28312 , \28323 );
xor \U$27948 ( \28325 , \27974 , \27984 );
xor \U$27949 ( \28326 , \28325 , \27996 );
and \U$27950 ( \28327 , \28324 , \28326 );
nor \U$27951 ( \28328 , \28312 , \28323 );
nor \U$27952 ( \28329 , \28327 , \28328 );
not \U$27953 ( \28330 , \28329 );
not \U$27954 ( \28331 , RIc2258a0_63);
not \U$27955 ( \28332 , \13914 );
or \U$27956 ( \28333 , \28331 , \28332 );
not \U$27957 ( \28334 , RIc2258a0_63);
nand \U$27958 ( \28335 , \28334 , \2421 );
nand \U$27959 ( \28336 , \28333 , \28335 );
and \U$27960 ( \28337 , \28336 , \16891 );
and \U$27961 ( \28338 , \27398 , RIc225828_64);
nor \U$27962 ( \28339 , \28337 , \28338 );
not \U$27963 ( \28340 , \28339 );
not \U$27964 ( \28341 , \28340 );
and \U$27965 ( \28342 , RIc225990_61, \2225 );
not \U$27966 ( \28343 , RIc225990_61);
and \U$27967 ( \28344 , \28343 , \9599 );
nor \U$27968 ( \28345 , \28342 , \28344 );
and \U$27969 ( \28346 , \28345 , \15719 );
and \U$27970 ( \28347 , \27484 , \15729 );
nor \U$27971 ( \28348 , \28346 , \28347 );
not \U$27972 ( \28349 , \28348 );
not \U$27973 ( \28350 , \28349 );
or \U$27974 ( \28351 , \28341 , \28350 );
not \U$27975 ( \28352 , \28339 );
not \U$27976 ( \28353 , \28348 );
or \U$27977 ( \28354 , \28352 , \28353 );
not \U$27978 ( \28355 , \11118 );
and \U$27979 ( \28356 , RIc225c60_55, \2476 );
not \U$27980 ( \28357 , RIc225c60_55);
and \U$27981 ( \28358 , \28357 , \3036 );
or \U$27982 ( \28359 , \28356 , \28358 );
not \U$27983 ( \28360 , \28359 );
or \U$27984 ( \28361 , \28355 , \28360 );
nand \U$27985 ( \28362 , \27471 , \12532 );
nand \U$27986 ( \28363 , \28361 , \28362 );
nand \U$27987 ( \28364 , \28354 , \28363 );
nand \U$27988 ( \28365 , \28351 , \28364 );
not \U$27989 ( \28366 , \28365 );
not \U$27990 ( \28367 , \28366 );
or \U$27991 ( \28368 , \28330 , \28367 );
xor \U$27992 ( \28369 , \27960 , \27999 );
xor \U$27993 ( \28370 , \28369 , \28009 );
nand \U$27994 ( \28371 , \28368 , \28370 );
not \U$27995 ( \28372 , \28329 );
nand \U$27996 ( \28373 , \28372 , \28365 );
and \U$27997 ( \28374 , \28371 , \28373 );
not \U$27998 ( \28375 , \28374 );
not \U$27999 ( \28376 , \28375 );
or \U$28000 ( \28377 , \28300 , \28376 );
nand \U$28001 ( \28378 , \28374 , \28298 );
nand \U$28002 ( \28379 , \28377 , \28378 );
buf \U$28003 ( \28380 , \28379 );
not \U$28004 ( \28381 , \28380 );
xor \U$28005 ( \28382 , \28081 , \28176 );
xor \U$28006 ( \28383 , \28382 , \28179 );
not \U$28007 ( \28384 , \28383 );
or \U$28008 ( \28385 , \28381 , \28384 );
or \U$28009 ( \28386 , \28380 , \28383 );
and \U$28010 ( \28387 , \28083 , \28118 );
not \U$28011 ( \28388 , \28083 );
and \U$28012 ( \28389 , \28388 , \28119 );
nor \U$28013 ( \28390 , \28387 , \28389 );
not \U$28014 ( \28391 , \28390 );
and \U$28015 ( \28392 , \28172 , \28391 );
not \U$28016 ( \28393 , \28172 );
and \U$28017 ( \28394 , \28393 , \28390 );
nor \U$28018 ( \28395 , \28392 , \28394 );
not \U$28019 ( \28396 , \28395 );
not \U$28020 ( \28397 , \28396 );
xor \U$28021 ( \28398 , \28225 , \28237 );
xnor \U$28022 ( \28399 , \28398 , \28250 );
not \U$28023 ( \28400 , \28399 );
not \U$28024 ( \28401 , \28400 );
not \U$28025 ( \28402 , \28285 );
not \U$28026 ( \28403 , \28264 );
or \U$28027 ( \28404 , \28402 , \28403 );
or \U$28028 ( \28405 , \28285 , \28264 );
nand \U$28029 ( \28406 , \28404 , \28405 );
not \U$28030 ( \28407 , \28274 );
and \U$28031 ( \28408 , \28406 , \28407 );
not \U$28032 ( \28409 , \28406 );
and \U$28033 ( \28410 , \28409 , \28274 );
nor \U$28034 ( \28411 , \28408 , \28410 );
not \U$28035 ( \28412 , \28411 );
or \U$28036 ( \28413 , \28401 , \28412 );
not \U$28037 ( \28414 , \28399 );
not \U$28038 ( \28415 , \28411 );
not \U$28039 ( \28416 , \28415 );
or \U$28040 ( \28417 , \28414 , \28416 );
not \U$28041 ( \28418 , \16891 );
not \U$28042 ( \28419 , RIc2258a0_63);
not \U$28043 ( \28420 , \2444 );
or \U$28044 ( \28421 , \28419 , \28420 );
nand \U$28045 ( \28422 , \2443 , \16880 );
nand \U$28046 ( \28423 , \28421 , \28422 );
not \U$28047 ( \28424 , \28423 );
or \U$28048 ( \28425 , \28418 , \28424 );
nand \U$28049 ( \28426 , \28336 , RIc225828_64);
nand \U$28050 ( \28427 , \28425 , \28426 );
not \U$28051 ( \28428 , \28427 );
not \U$28052 ( \28429 , \28428 );
not \U$28053 ( \28430 , RIc226020_47);
not \U$28054 ( \28431 , \9674 );
or \U$28055 ( \28432 , \28430 , \28431 );
nand \U$28056 ( \28433 , \3640 , \9624 );
nand \U$28057 ( \28434 , \28432 , \28433 );
not \U$28058 ( \28435 , \28434 );
not \U$28059 ( \28436 , \28435 );
not \U$28060 ( \28437 , \9640 );
and \U$28061 ( \28438 , \28436 , \28437 );
not \U$28062 ( \28439 , RIc226020_47);
not \U$28063 ( \28440 , \12493 );
or \U$28064 ( \28441 , \28439 , \28440 );
nand \U$28065 ( \28442 , \2980 , \9624 );
nand \U$28066 ( \28443 , \28441 , \28442 );
and \U$28067 ( \28444 , \28443 , \10953 );
nor \U$28068 ( \28445 , \28438 , \28444 );
not \U$28069 ( \28446 , \28445 );
or \U$28070 ( \28447 , \28429 , \28446 );
not \U$28071 ( \28448 , \11118 );
not \U$28072 ( \28449 , RIc225c60_55);
not \U$28073 ( \28450 , \2894 );
or \U$28074 ( \28451 , \28449 , \28450 );
nand \U$28075 ( \28452 , \4196 , \8767 );
nand \U$28076 ( \28453 , \28451 , \28452 );
not \U$28077 ( \28454 , \28453 );
or \U$28078 ( \28455 , \28448 , \28454 );
nand \U$28079 ( \28456 , \28359 , \11038 );
nand \U$28080 ( \28457 , \28455 , \28456 );
nand \U$28081 ( \28458 , \28447 , \28457 );
not \U$28082 ( \28459 , \28445 );
nand \U$28083 ( \28460 , \28459 , \28427 );
nand \U$28084 ( \28461 , \28458 , \28460 );
nand \U$28085 ( \28462 , \28417 , \28461 );
nand \U$28086 ( \28463 , \28413 , \28462 );
not \U$28087 ( \28464 , \28463 );
or \U$28088 ( \28465 , \28397 , \28464 );
not \U$28089 ( \28466 , \28395 );
not \U$28090 ( \28467 , \28463 );
not \U$28091 ( \28468 , \28467 );
or \U$28092 ( \28469 , \28466 , \28468 );
not \U$28093 ( \28470 , \9205 );
not \U$28094 ( \28471 , \28261 );
or \U$28095 ( \28472 , \28470 , \28471 );
not \U$28096 ( \28473 , RIc226200_43);
not \U$28097 ( \28474 , \5664 );
or \U$28098 ( \28475 , \28473 , \28474 );
nand \U$28099 ( \28476 , \5663 , \9117 );
nand \U$28100 ( \28477 , \28475 , \28476 );
nand \U$28101 ( \28478 , \28477 , \9110 );
nand \U$28102 ( \28479 , \28472 , \28478 );
not \U$28103 ( \28480 , \2710 );
not \U$28104 ( \28481 , \28272 );
or \U$28105 ( \28482 , \28480 , \28481 );
and \U$28106 ( \28483 , RIc2267a0_31, \28026 );
not \U$28107 ( \28484 , RIc2267a0_31);
and \U$28108 ( \28485 , \28484 , \8924 );
or \U$28109 ( \28486 , \28483 , \28485 );
nand \U$28110 ( \28487 , \28486 , \2697 );
nand \U$28111 ( \28488 , \28482 , \28487 );
xor \U$28112 ( \28489 , \28479 , \28488 );
not \U$28113 ( \28490 , \9398 );
not \U$28114 ( \28491 , \28113 );
or \U$28115 ( \28492 , \28490 , \28491 );
not \U$28116 ( \28493 , RIc226110_45);
not \U$28117 ( \28494 , \9842 );
or \U$28118 ( \28495 , \28493 , \28494 );
nand \U$28119 ( \28496 , \4406 , \9100 );
nand \U$28120 ( \28497 , \28495 , \28496 );
nand \U$28121 ( \28498 , \28497 , \9934 );
nand \U$28122 ( \28499 , \28492 , \28498 );
and \U$28123 ( \28500 , \28489 , \28499 );
and \U$28124 ( \28501 , \28479 , \28488 );
or \U$28125 ( \28502 , \28500 , \28501 );
not \U$28126 ( \28503 , \15719 );
and \U$28127 ( \28504 , RIc225990_61, \2257 );
not \U$28128 ( \28505 , RIc225990_61);
and \U$28129 ( \28506 , \28505 , \4008 );
or \U$28130 ( \28507 , \28504 , \28506 );
not \U$28131 ( \28508 , \28507 );
or \U$28132 ( \28509 , \28503 , \28508 );
nand \U$28133 ( \28510 , \28345 , \15729 );
nand \U$28134 ( \28511 , \28509 , \28510 );
not \U$28135 ( \28512 , \9555 );
and \U$28136 ( \28513 , RIc225d50_53, \3810 );
not \U$28137 ( \28514 , RIc225d50_53);
and \U$28138 ( \28515 , \28514 , \2720 );
or \U$28139 ( \28516 , \28513 , \28515 );
not \U$28140 ( \28517 , \28516 );
or \U$28141 ( \28518 , \28512 , \28517 );
and \U$28142 ( \28519 , RIc225d50_53, \2063 );
not \U$28143 ( \28520 , RIc225d50_53);
and \U$28144 ( \28521 , \28520 , \3008 );
or \U$28145 ( \28522 , \28519 , \28521 );
nand \U$28146 ( \28523 , \28522 , \9488 );
nand \U$28147 ( \28524 , \28518 , \28523 );
xor \U$28148 ( \28525 , \28511 , \28524 );
not \U$28149 ( \28526 , \15164 );
and \U$28150 ( \28527 , RIc225a80_59, \9433 );
not \U$28151 ( \28528 , RIc225a80_59);
and \U$28152 ( \28529 , \28528 , \2014 );
or \U$28153 ( \28530 , \28527 , \28529 );
not \U$28154 ( \28531 , \28530 );
or \U$28155 ( \28532 , \28526 , \28531 );
nand \U$28156 ( \28533 , \28309 , \12670 );
nand \U$28157 ( \28534 , \28532 , \28533 );
and \U$28158 ( \28535 , \28525 , \28534 );
and \U$28159 ( \28536 , \28511 , \28524 );
or \U$28160 ( \28537 , \28535 , \28536 );
xor \U$28161 ( \28538 , \28502 , \28537 );
xor \U$28162 ( \28539 , \28146 , \28157 );
xor \U$28163 ( \28540 , \28539 , \28169 );
and \U$28164 ( \28541 , \28538 , \28540 );
and \U$28165 ( \28542 , \28502 , \28537 );
or \U$28166 ( \28543 , \28541 , \28542 );
nand \U$28167 ( \28544 , \28469 , \28543 );
nand \U$28168 ( \28545 , \28465 , \28544 );
nand \U$28169 ( \28546 , \28386 , \28545 );
nand \U$28170 ( \28547 , \28385 , \28546 );
not \U$28171 ( \28548 , \28547 );
xor \U$28172 ( \28549 , \27955 , \27957 );
xor \U$28173 ( \28550 , \28549 , \28182 );
not \U$28174 ( \28551 , \28550 );
nand \U$28175 ( \28552 , \28548 , \28551 );
not \U$28176 ( \28553 , \28552 );
nand \U$28177 ( \28554 , \28291 , \28293 );
not \U$28178 ( \28555 , \28554 );
not \U$28179 ( \28556 , \28375 );
or \U$28180 ( \28557 , \28555 , \28556 );
not \U$28181 ( \28558 , \28291 );
nand \U$28182 ( \28559 , \28558 , \28296 );
nand \U$28183 ( \28560 , \28557 , \28559 );
xor \U$28184 ( \28561 , \27224 , \27233 );
xor \U$28185 ( \28562 , \28561 , \27250 );
xor \U$28186 ( \28563 , \27328 , \27338 );
and \U$28187 ( \28564 , \28563 , \27344 );
and \U$28188 ( \28565 , \27328 , \27338 );
or \U$28189 ( \28566 , \28564 , \28565 );
xor \U$28190 ( \28567 , \28562 , \28566 );
xor \U$28191 ( \28568 , \27355 , \27364 );
and \U$28192 ( \28569 , \28568 , \27375 );
and \U$28193 ( \28570 , \27355 , \27364 );
or \U$28194 ( \28571 , \28569 , \28570 );
xor \U$28195 ( \28572 , \28567 , \28571 );
xor \U$28196 ( \28573 , \28012 , \28046 );
and \U$28197 ( \28574 , \28573 , \28080 );
and \U$28198 ( \28575 , \28012 , \28046 );
or \U$28199 ( \28576 , \28574 , \28575 );
xor \U$28200 ( \28577 , \28572 , \28576 );
xor \U$28201 ( \28578 , \27307 , \27311 );
xor \U$28202 ( \28579 , \28578 , \27316 );
xor \U$28203 ( \28580 , \28577 , \28579 );
xor \U$28204 ( \28581 , \28560 , \28580 );
xor \U$28205 ( \28582 , \27423 , \27539 );
xor \U$28206 ( \28583 , \28582 , \27562 );
xor \U$28207 ( \28584 , \28581 , \28583 );
not \U$28208 ( \28585 , \28584 );
or \U$28209 ( \28586 , \28553 , \28585 );
nand \U$28210 ( \28587 , \28547 , \28550 );
nand \U$28211 ( \28588 , \28586 , \28587 );
nand \U$28212 ( \28589 , \28189 , \28588 );
nand \U$28213 ( \28590 , \28188 , \28589 );
not \U$28214 ( \28591 , \28590 );
not \U$28215 ( \28592 , \9458 );
not \U$28216 ( \28593 , RIc225e40_51);
not \U$28217 ( \28594 , \2554 );
or \U$28218 ( \28595 , \28593 , \28594 );
nand \U$28219 ( \28596 , \3446 , \9450 );
nand \U$28220 ( \28597 , \28595 , \28596 );
not \U$28221 ( \28598 , \28597 );
or \U$28222 ( \28599 , \28592 , \28598 );
not \U$28223 ( \28600 , RIc225e40_51);
not \U$28224 ( \28601 , \12519 );
or \U$28225 ( \28602 , \28600 , \28601 );
nand \U$28226 ( \28603 , \2590 , \12423 );
nand \U$28227 ( \28604 , \28602 , \28603 );
nand \U$28228 ( \28605 , \28604 , \9444 );
nand \U$28229 ( \28606 , \28599 , \28605 );
not \U$28230 ( \28607 , \15164 );
and \U$28231 ( \28608 , RIc225a80_59, \3092 );
not \U$28232 ( \28609 , RIc225a80_59);
and \U$28233 ( \28610 , \28609 , \8989 );
or \U$28234 ( \28611 , \28608 , \28610 );
not \U$28235 ( \28612 , \28611 );
or \U$28236 ( \28613 , \28607 , \28612 );
and \U$28237 ( \28614 , RIc225a80_59, \4473 );
not \U$28238 ( \28615 , RIc225a80_59);
and \U$28239 ( \28616 , \28615 , \2353 );
or \U$28240 ( \28617 , \28614 , \28616 );
nand \U$28241 ( \28618 , \28617 , \12670 );
nand \U$28242 ( \28619 , \28613 , \28618 );
xor \U$28243 ( \28620 , \28606 , \28619 );
not \U$28244 ( \28621 , \8777 );
and \U$28245 ( \28622 , \9433 , RIc225d50_53);
not \U$28246 ( \28623 , \9433 );
and \U$28247 ( \28624 , \28623 , \8772 );
or \U$28248 ( \28625 , \28622 , \28624 );
not \U$28249 ( \28626 , \28625 );
or \U$28250 ( \28627 , \28621 , \28626 );
not \U$28251 ( \28628 , RIc225d50_53);
not \U$28252 ( \28629 , \12508 );
or \U$28253 ( \28630 , \28628 , \28629 );
nand \U$28254 ( \28631 , \1988 , \11585 );
nand \U$28255 ( \28632 , \28630 , \28631 );
nand \U$28256 ( \28633 , \28632 , \9555 );
nand \U$28257 ( \28634 , \28627 , \28633 );
xor \U$28258 ( \28635 , \28620 , \28634 );
not \U$28259 ( \28636 , \27280 );
not \U$28260 ( \28637 , \27295 );
or \U$28261 ( \28638 , \28636 , \28637 );
or \U$28262 ( \28639 , \27280 , \27295 );
nand \U$28263 ( \28640 , \28639 , \27305 );
nand \U$28264 ( \28641 , \28638 , \28640 );
not \U$28265 ( \28642 , \12670 );
not \U$28266 ( \28643 , \28611 );
or \U$28267 ( \28644 , \28642 , \28643 );
nand \U$28268 ( \28645 , \27763 , \15164 );
nand \U$28269 ( \28646 , \28644 , \28645 );
xor \U$28270 ( \28647 , \28641 , \28646 );
not \U$28271 ( \28648 , \9459 );
not \U$28272 ( \28649 , \27753 );
or \U$28273 ( \28650 , \28648 , \28649 );
nand \U$28274 ( \28651 , \28597 , \9444 );
nand \U$28275 ( \28652 , \28650 , \28651 );
and \U$28276 ( \28653 , \28647 , \28652 );
and \U$28277 ( \28654 , \28641 , \28646 );
or \U$28278 ( \28655 , \28653 , \28654 );
and \U$28279 ( \28656 , \28635 , \28655 );
not \U$28280 ( \28657 , \28635 );
not \U$28281 ( \28658 , \28655 );
and \U$28282 ( \28659 , \28657 , \28658 );
nor \U$28283 ( \28660 , \28656 , \28659 );
and \U$28284 ( \28661 , \26866 , \26879 );
not \U$28285 ( \28662 , \2320 );
not \U$28286 ( \28663 , \27229 );
or \U$28287 ( \28664 , \28662 , \28663 );
not \U$28288 ( \28665 , RIc226f20_15);
not \U$28289 ( \28666 , \16492 );
or \U$28290 ( \28667 , \28665 , \28666 );
nand \U$28291 ( \28668 , \13497 , \2351 );
nand \U$28292 ( \28669 , \28667 , \28668 );
nand \U$28293 ( \28670 , \28669 , \2318 );
nand \U$28294 ( \28671 , \28664 , \28670 );
xor \U$28295 ( \28672 , \28661 , \28671 );
not \U$28296 ( \28673 , \1963 );
not \U$28297 ( \28674 , RIc226e30_17);
not \U$28298 ( \28675 , \12862 );
or \U$28299 ( \28676 , \28674 , \28675 );
nand \U$28300 ( \28677 , \10086 , \1960 );
nand \U$28301 ( \28678 , \28676 , \28677 );
not \U$28302 ( \28679 , \28678 );
or \U$28303 ( \28680 , \28673 , \28679 );
nand \U$28304 ( \28681 , \26902 , \1945 );
nand \U$28305 ( \28682 , \28680 , \28681 );
and \U$28306 ( \28683 , \28672 , \28682 );
and \U$28307 ( \28684 , \28661 , \28671 );
or \U$28308 ( \28685 , \28683 , \28684 );
not \U$28309 ( \28686 , \15719 );
not \U$28310 ( \28687 , \27818 );
or \U$28311 ( \28688 , \28686 , \28687 );
not \U$28312 ( \28689 , RIc225990_61);
not \U$28313 ( \28690 , \9115 );
or \U$28314 ( \28691 , \28689 , \28690 );
nand \U$28315 ( \28692 , \3043 , \12806 );
nand \U$28316 ( \28693 , \28691 , \28692 );
nand \U$28317 ( \28694 , \28693 , \15729 );
nand \U$28318 ( \28695 , \28688 , \28694 );
xor \U$28319 ( \28696 , \28685 , \28695 );
not \U$28320 ( \28697 , \10445 );
not \U$28321 ( \28698 , RIc225f30_49);
not \U$28322 ( \28699 , \12989 );
or \U$28323 ( \28700 , \28698 , \28699 );
nand \U$28324 ( \28701 , \2500 , \9549 );
nand \U$28325 ( \28702 , \28700 , \28701 );
not \U$28326 ( \28703 , \28702 );
or \U$28327 ( \28704 , \28697 , \28703 );
not \U$28328 ( \28705 , RIc225f30_49);
not \U$28329 ( \28706 , \2475 );
not \U$28330 ( \28707 , \28706 );
or \U$28331 ( \28708 , \28705 , \28707 );
not \U$28332 ( \28709 , RIc225f30_49);
nand \U$28333 ( \28710 , \28709 , \3036 );
nand \U$28334 ( \28711 , \28708 , \28710 );
nand \U$28335 ( \28712 , \28711 , \9552 );
nand \U$28336 ( \28713 , \28704 , \28712 );
xor \U$28337 ( \28714 , \28696 , \28713 );
and \U$28338 ( \28715 , \28660 , \28714 );
not \U$28339 ( \28716 , \28660 );
not \U$28340 ( \28717 , \28714 );
and \U$28341 ( \28718 , \28716 , \28717 );
nor \U$28342 ( \28719 , \28715 , \28718 );
xor \U$28343 ( \28720 , \27568 , \27577 );
and \U$28344 ( \28721 , \28720 , \27588 );
and \U$28345 ( \28722 , \27568 , \27577 );
or \U$28346 ( \28723 , \28721 , \28722 );
not \U$28347 ( \28724 , \2320 );
not \U$28348 ( \28725 , \28669 );
or \U$28349 ( \28726 , \28724 , \28725 );
nand \U$28350 ( \28727 , \21978 , \2318 );
nand \U$28351 ( \28728 , \28726 , \28727 );
xor \U$28352 ( \28729 , \28723 , \28728 );
not \U$28353 ( \28730 , \2391 );
not \U$28354 ( \28731 , \27608 );
or \U$28355 ( \28732 , \28730 , \28731 );
not \U$28356 ( \28733 , RIc226c50_21);
not \U$28357 ( \28734 , \13223 );
or \U$28358 ( \28735 , \28733 , \28734 );
nand \U$28359 ( \28736 , \10110 , \2370 );
nand \U$28360 ( \28737 , \28735 , \28736 );
nand \U$28361 ( \28738 , \28737 , \2367 );
nand \U$28362 ( \28739 , \28732 , \28738 );
xor \U$28363 ( \28740 , \28729 , \28739 );
xor \U$28364 ( \28741 , \27589 , \27599 );
and \U$28365 ( \28742 , \28741 , \27610 );
and \U$28366 ( \28743 , \27589 , \27599 );
or \U$28367 ( \28744 , \28742 , \28743 );
xor \U$28368 ( \28745 , \28740 , \28744 );
not \U$28369 ( \28746 , \16891 );
not \U$28370 ( \28747 , RIc2258a0_63);
not \U$28371 ( \28748 , \3438 );
or \U$28372 ( \28749 , \28747 , \28748 );
not \U$28373 ( \28750 , RIc2258a0_63);
nand \U$28374 ( \28751 , \1332 , \28750 );
nand \U$28375 ( \28752 , \28749 , \28751 );
not \U$28376 ( \28753 , \28752 );
or \U$28377 ( \28754 , \28746 , \28753 );
not \U$28378 ( \28755 , RIc2258a0_63);
not \U$28379 ( \28756 , \4590 );
or \U$28380 ( \28757 , \28755 , \28756 );
nand \U$28381 ( \28758 , \1529 , \16880 );
nand \U$28382 ( \28759 , \28757 , \28758 );
nand \U$28383 ( \28760 , \28759 , RIc225828_64);
nand \U$28384 ( \28761 , \28754 , \28760 );
xor \U$28385 ( \28762 , \28745 , \28761 );
xor \U$28386 ( \28763 , \27611 , \27642 );
and \U$28387 ( \28764 , \28763 , \27647 );
and \U$28388 ( \28765 , \27611 , \27642 );
or \U$28389 ( \28766 , \28764 , \28765 );
xor \U$28390 ( \28767 , \28762 , \28766 );
not \U$28391 ( \28768 , RIc226200_43);
not \U$28392 ( \28769 , \3119 );
or \U$28393 ( \28770 , \28768 , \28769 );
nand \U$28394 ( \28771 , \3115 , \9125 );
nand \U$28395 ( \28772 , \28770 , \28771 );
not \U$28396 ( \28773 , \28772 );
not \U$28397 ( \28774 , \28773 );
not \U$28398 ( \28775 , \9109 );
and \U$28399 ( \28776 , \28774 , \28775 );
not \U$28400 ( \28777 , RIc226200_43);
not \U$28401 ( \28778 , \2104 );
or \U$28402 ( \28779 , \28777 , \28778 );
not \U$28403 ( \28780 , \3715 );
nand \U$28404 ( \28781 , \28780 , \13805 );
nand \U$28405 ( \28782 , \28779 , \28781 );
and \U$28406 ( \28783 , \28782 , \9205 );
nor \U$28407 ( \28784 , \28776 , \28783 );
not \U$28408 ( \28785 , \28784 );
not \U$28409 ( \28786 , \9705 );
xor \U$28410 ( \28787 , RIc2262f0_41, \3725 );
not \U$28411 ( \28788 , \28787 );
or \U$28412 ( \28789 , \28786 , \28788 );
nand \U$28413 ( \28790 , \27848 , \9690 );
nand \U$28414 ( \28791 , \28789 , \28790 );
not \U$28415 ( \28792 , \28791 );
not \U$28416 ( \28793 , \11117 );
not \U$28417 ( \28794 , RIc225c60_55);
not \U$28418 ( \28795 , \4009 );
or \U$28419 ( \28796 , \28794 , \28795 );
nand \U$28420 ( \28797 , \4008 , \11041 );
nand \U$28421 ( \28798 , \28796 , \28797 );
not \U$28422 ( \28799 , \28798 );
or \U$28423 ( \28800 , \28793 , \28799 );
not \U$28424 ( \28801 , RIc225c60_55);
not \U$28425 ( \28802 , \16762 );
or \U$28426 ( \28803 , \28801 , \28802 );
nand \U$28427 ( \28804 , \18087 , \11108 );
nand \U$28428 ( \28805 , \28803 , \28804 );
nand \U$28429 ( \28806 , \28805 , \12532 );
nand \U$28430 ( \28807 , \28800 , \28806 );
not \U$28431 ( \28808 , \28807 );
not \U$28432 ( \28809 , \28808 );
or \U$28433 ( \28810 , \28792 , \28809 );
or \U$28434 ( \28811 , \28808 , \28791 );
nand \U$28435 ( \28812 , \28810 , \28811 );
xor \U$28436 ( \28813 , \28785 , \28812 );
xor \U$28437 ( \28814 , \28767 , \28813 );
xor \U$28438 ( \28815 , \28719 , \28814 );
xor \U$28439 ( \28816 , \27265 , \27319 );
and \U$28440 ( \28817 , \28816 , \27324 );
and \U$28441 ( \28818 , \27265 , \27319 );
or \U$28442 ( \28819 , \28817 , \28818 );
xor \U$28443 ( \28820 , \28815 , \28819 );
not \U$28444 ( \28821 , \28820 );
not \U$28445 ( \28822 , \28821 );
not \U$28446 ( \28823 , \27257 );
not \U$28447 ( \28824 , \27264 );
or \U$28448 ( \28825 , \28823 , \28824 );
nand \U$28449 ( \28826 , \28825 , \27253 );
not \U$28450 ( \28827 , \27264 );
not \U$28451 ( \28828 , \27257 );
nand \U$28452 ( \28829 , \28827 , \28828 );
and \U$28453 ( \28830 , \28826 , \28829 );
not \U$28454 ( \28831 , \2518 );
not \U$28455 ( \28832 , \27619 );
or \U$28456 ( \28833 , \28831 , \28832 );
not \U$28457 ( \28834 , RIc226d40_19);
not \U$28458 ( \28835 , \10800 );
or \U$28459 ( \28836 , \28834 , \28835 );
nand \U$28460 ( \28837 , \9274 , \2523 );
nand \U$28461 ( \28838 , \28836 , \28837 );
nand \U$28462 ( \28839 , \28838 , \2533 );
nand \U$28463 ( \28840 , \28833 , \28839 );
not \U$28464 ( \28841 , RIc226b60_23);
not \U$28465 ( \28842 , \9049 );
or \U$28466 ( \28843 , \28841 , \28842 );
nand \U$28467 ( \28844 , \9045 , \1927 );
nand \U$28468 ( \28845 , \28843 , \28844 );
not \U$28469 ( \28846 , \28845 );
not \U$28470 ( \28847 , \1930 );
or \U$28471 ( \28848 , \28846 , \28847 );
nand \U$28472 ( \28849 , \27597 , \1914 );
nand \U$28473 ( \28850 , \28848 , \28849 );
xor \U$28474 ( \28851 , \28840 , \28850 );
not \U$28475 ( \28852 , \1963 );
not \U$28476 ( \28853 , RIc226e30_17);
not \U$28477 ( \28854 , \9321 );
or \U$28478 ( \28855 , \28853 , \28854 );
nand \U$28479 ( \28856 , \9324 , \1960 );
nand \U$28480 ( \28857 , \28855 , \28856 );
not \U$28481 ( \28858 , \28857 );
or \U$28482 ( \28859 , \28852 , \28858 );
nand \U$28483 ( \28860 , \28678 , \1945 );
nand \U$28484 ( \28861 , \28859 , \28860 );
xor \U$28485 ( \28862 , \28851 , \28861 );
xor \U$28486 ( \28863 , \27621 , \27631 );
and \U$28487 ( \28864 , \28863 , \27641 );
and \U$28488 ( \28865 , \27621 , \27631 );
or \U$28489 ( \28866 , \28864 , \28865 );
xor \U$28490 ( \28867 , \28862 , \28866 );
not \U$28491 ( \28868 , \2086 );
and \U$28492 ( \28869 , RIc226890_29, \8807 );
not \U$28493 ( \28870 , RIc226890_29);
and \U$28494 ( \28871 , \28870 , \8806 );
or \U$28495 ( \28872 , \28869 , \28871 );
not \U$28496 ( \28873 , \28872 );
or \U$28497 ( \28874 , \28868 , \28873 );
nand \U$28498 ( \28875 , \26980 , \2784 );
nand \U$28499 ( \28876 , \28874 , \28875 );
not \U$28500 ( \28877 , \3629 );
not \U$28501 ( \28878 , \27006 );
or \U$28502 ( \28879 , \28877 , \28878 );
not \U$28503 ( \28880 , RIc2266b0_33);
not \U$28504 ( \28881 , \15699 );
or \U$28505 ( \28882 , \28880 , \28881 );
nand \U$28506 ( \28883 , \10141 , \12551 );
nand \U$28507 ( \28884 , \28882 , \28883 );
nand \U$28508 ( \28885 , \28884 , \3631 );
nand \U$28509 ( \28886 , \28879 , \28885 );
nor \U$28510 ( \28887 , \28876 , \28886 );
not \U$28511 ( \28888 , RIc226980_27);
not \U$28512 ( \28889 , \21866 );
or \U$28513 ( \28890 , \28888 , \28889 );
nand \U$28514 ( \28891 , \8974 , \4528 );
nand \U$28515 ( \28892 , \28890 , \28891 );
and \U$28516 ( \28893 , \28892 , \2154 );
and \U$28517 ( \28894 , \26945 , \2138 );
nor \U$28518 ( \28895 , \28893 , \28894 );
or \U$28519 ( \28896 , \28887 , \28895 );
nand \U$28520 ( \28897 , \28886 , \28876 );
nand \U$28521 ( \28898 , \28896 , \28897 );
xor \U$28522 ( \28899 , \28867 , \28898 );
and \U$28523 ( \28900 , \28830 , \28899 );
not \U$28524 ( \28901 , \28830 );
not \U$28525 ( \28902 , \28899 );
and \U$28526 ( \28903 , \28901 , \28902 );
or \U$28527 ( \28904 , \28900 , \28903 );
not \U$28528 ( \28905 , \27937 );
not \U$28529 ( \28906 , \27950 );
or \U$28530 ( \28907 , \28905 , \28906 );
not \U$28531 ( \28908 , \27949 );
not \U$28532 ( \28909 , \27936 );
or \U$28533 ( \28910 , \28908 , \28909 );
nand \U$28534 ( \28911 , \28910 , \27941 );
nand \U$28535 ( \28912 , \28907 , \28911 );
xor \U$28536 ( \28913 , \28904 , \28912 );
xor \U$28537 ( \28914 , \27648 , \27657 );
and \U$28538 ( \28915 , \28914 , \27788 );
and \U$28539 ( \28916 , \27648 , \27657 );
or \U$28540 ( \28917 , \28915 , \28916 );
xor \U$28541 ( \28918 , \28913 , \28917 );
xor \U$28542 ( \28919 , \27863 , \27931 );
and \U$28543 ( \28920 , \28919 , \27951 );
and \U$28544 ( \28921 , \27863 , \27931 );
or \U$28545 ( \28922 , \28920 , \28921 );
xnor \U$28546 ( \28923 , \28918 , \28922 );
not \U$28547 ( \28924 , \28923 );
not \U$28548 ( \28925 , \28924 );
or \U$28549 ( \28926 , \28822 , \28925 );
nand \U$28550 ( \28927 , \28923 , \28820 );
nand \U$28551 ( \28928 , \28926 , \28927 );
or \U$28552 ( \28929 , \27201 , \27325 );
and \U$28553 ( \28930 , \27565 , \28929 );
and \U$28554 ( \28931 , \27201 , \27325 );
nor \U$28555 ( \28932 , \28930 , \28931 );
and \U$28556 ( \28933 , \28928 , \28932 );
not \U$28557 ( \28934 , \28928 );
not \U$28558 ( \28935 , \28932 );
and \U$28559 ( \28936 , \28934 , \28935 );
nor \U$28560 ( \28937 , \28933 , \28936 );
not \U$28561 ( \28938 , \28937 );
and \U$28562 ( \28939 , \28591 , \28938 );
and \U$28563 ( \28940 , \28590 , \28937 );
nor \U$28564 ( \28941 , \28939 , \28940 );
buf \U$28565 ( \28942 , \27789 );
not \U$28566 ( \28943 , \28942 );
not \U$28567 ( \28944 , \27952 );
nand \U$28568 ( \28945 , \28943 , \28944 );
and \U$28569 ( \28946 , \28945 , \28185 );
not \U$28570 ( \28947 , \28942 );
nor \U$28571 ( \28948 , \28947 , \28944 );
nor \U$28572 ( \28949 , \28946 , \28948 );
not \U$28573 ( \28950 , \28949 );
xor \U$28574 ( \28951 , \28661 , \28671 );
xor \U$28575 ( \28952 , \28951 , \28682 );
not \U$28576 ( \28953 , RIc225828_64);
not \U$28577 ( \28954 , \28752 );
or \U$28578 ( \28955 , \28953 , \28954 );
nand \U$28579 ( \28956 , \16891 , \27778 );
nand \U$28580 ( \28957 , \28955 , \28956 );
xor \U$28581 ( \28958 , \28952 , \28957 );
not \U$28582 ( \28959 , \8788 );
not \U$28583 ( \28960 , \28625 );
or \U$28584 ( \28961 , \28959 , \28960 );
nand \U$28585 ( \28962 , \27739 , \9488 );
nand \U$28586 ( \28963 , \28961 , \28962 );
xnor \U$28587 ( \28964 , \28958 , \28963 );
not \U$28588 ( \28965 , \28964 );
not \U$28589 ( \28966 , \28965 );
not \U$28590 ( \28967 , \9129 );
not \U$28591 ( \28968 , \28772 );
or \U$28592 ( \28969 , \28967 , \28968 );
nand \U$28593 ( \28970 , \27718 , \9110 );
nand \U$28594 ( \28971 , \28969 , \28970 );
not \U$28595 ( \28972 , \28971 );
not \U$28596 ( \28973 , \28972 );
not \U$28597 ( \28974 , \13025 );
not \U$28598 ( \28975 , \28798 );
or \U$28599 ( \28976 , \28974 , \28975 );
nand \U$28600 ( \28977 , \27730 , \11697 );
nand \U$28601 ( \28978 , \28976 , \28977 );
not \U$28602 ( \28979 , \28978 );
and \U$28603 ( \28980 , \28973 , \28979 );
and \U$28604 ( \28981 , \28972 , \28978 );
nor \U$28605 ( \28982 , \28980 , \28981 );
not \U$28606 ( \28983 , \27920 );
not \U$28607 ( \28984 , \9934 );
not \U$28608 ( \28985 , \28984 );
and \U$28609 ( \28986 , \28983 , \28985 );
not \U$28610 ( \28987 , RIc226110_45);
not \U$28611 ( \28988 , \14476 );
or \U$28612 ( \28989 , \28987 , \28988 );
nand \U$28613 ( \28990 , \18240 , \14390 );
nand \U$28614 ( \28991 , \28989 , \28990 );
and \U$28615 ( \28992 , \28991 , \9398 );
nor \U$28616 ( \28993 , \28986 , \28992 );
and \U$28617 ( \28994 , \28982 , \28993 );
not \U$28618 ( \28995 , \28982 );
not \U$28619 ( \28996 , \28993 );
and \U$28620 ( \28997 , \28995 , \28996 );
nor \U$28621 ( \28998 , \28994 , \28997 );
not \U$28622 ( \28999 , \28998 );
not \U$28623 ( \29000 , \28999 );
or \U$28624 ( \29001 , \28966 , \29000 );
nand \U$28625 ( \29002 , \28998 , \28964 );
nand \U$28626 ( \29003 , \29001 , \29002 );
xor \U$28627 ( \29004 , \28562 , \28566 );
and \U$28628 ( \29005 , \29004 , \28571 );
and \U$28629 ( \29006 , \28562 , \28566 );
or \U$28630 ( \29007 , \29005 , \29006 );
not \U$28631 ( \29008 , \29007 );
and \U$28632 ( \29009 , \29003 , \29008 );
not \U$28633 ( \29010 , \29003 );
and \U$28634 ( \29011 , \29010 , \29007 );
nor \U$28635 ( \29012 , \29009 , \29011 );
not \U$28636 ( \29013 , \29012 );
not \U$28637 ( \29014 , \29013 );
xor \U$28638 ( \29015 , \28886 , \28876 );
not \U$28639 ( \29016 , \28895 );
xor \U$28640 ( \29017 , \29015 , \29016 );
xor \U$28641 ( \29018 , \28641 , \28646 );
xor \U$28642 ( \29019 , \29018 , \28652 );
xor \U$28643 ( \29020 , \29017 , \29019 );
not \U$28644 ( \29021 , \12304 );
not \U$28645 ( \29022 , RIc226020_47);
not \U$28646 ( \29023 , \12977 );
or \U$28647 ( \29024 , \29022 , \29023 );
nand \U$28648 ( \29025 , \11844 , \9373 );
nand \U$28649 ( \29026 , \29024 , \29025 );
not \U$28650 ( \29027 , \29026 );
or \U$28651 ( \29028 , \29021 , \29027 );
nand \U$28652 ( \29029 , \27895 , \10001 );
nand \U$28653 ( \29030 , \29028 , \29029 );
not \U$28654 ( \29031 , \29030 );
not \U$28655 ( \29032 , \9552 );
not \U$28656 ( \29033 , \28702 );
or \U$28657 ( \29034 , \29032 , \29033 );
nand \U$28658 ( \29035 , \27885 , \9534 );
nand \U$28659 ( \29036 , \29034 , \29035 );
not \U$28660 ( \29037 , \29036 );
not \U$28661 ( \29038 , \29037 );
or \U$28662 ( \29039 , \29031 , \29038 );
or \U$28663 ( \29040 , \29030 , \29037 );
nand \U$28664 ( \29041 , \29039 , \29040 );
not \U$28665 ( \29042 , \27908 );
not \U$28666 ( \29043 , \29042 );
not \U$28667 ( \29044 , \11965 );
not \U$28668 ( \29045 , \29044 );
and \U$28669 ( \29046 , \29043 , \29045 );
not \U$28670 ( \29047 , RIc225b70_57);
not \U$28671 ( \29048 , \2444 );
or \U$28672 ( \29049 , \29047 , \29048 );
nand \U$28673 ( \29050 , \5949 , \10074 );
nand \U$28674 ( \29051 , \29049 , \29050 );
and \U$28675 ( \29052 , \29051 , \11974 );
nor \U$28676 ( \29053 , \29046 , \29052 );
and \U$28677 ( \29054 , \29041 , \29053 );
not \U$28678 ( \29055 , \29041 );
not \U$28679 ( \29056 , \29053 );
and \U$28680 ( \29057 , \29055 , \29056 );
nor \U$28681 ( \29058 , \29054 , \29057 );
xor \U$28682 ( \29059 , \29020 , \29058 );
not \U$28683 ( \29060 , \29059 );
not \U$28684 ( \29061 , \29060 );
or \U$28685 ( \29062 , \29014 , \29061 );
not \U$28686 ( \29063 , \29059 );
not \U$28687 ( \29064 , \29012 );
or \U$28688 ( \29065 , \29063 , \29064 );
xor \U$28689 ( \29066 , \28572 , \28576 );
and \U$28690 ( \29067 , \29066 , \28579 );
and \U$28691 ( \29068 , \28572 , \28576 );
or \U$28692 ( \29069 , \29067 , \29068 );
nand \U$28693 ( \29070 , \29065 , \29069 );
nand \U$28694 ( \29071 , \29062 , \29070 );
xor \U$28695 ( \29072 , \27831 , \27841 );
and \U$28696 ( \29073 , \29072 , \27852 );
and \U$28697 ( \29074 , \27831 , \27841 );
or \U$28698 ( \29075 , \29073 , \29074 );
xor \U$28699 ( \29076 , \27793 , \27804 );
and \U$28700 ( \29077 , \29076 , \27820 );
and \U$28701 ( \29078 , \27793 , \27804 );
or \U$28702 ( \29079 , \29077 , \29078 );
xor \U$28703 ( \29080 , \29075 , \29079 );
not \U$28704 ( \29081 , \29037 );
not \U$28705 ( \29082 , \29053 );
or \U$28706 ( \29083 , \29081 , \29082 );
nand \U$28707 ( \29084 , \29083 , \29030 );
nand \U$28708 ( \29085 , \29056 , \29036 );
nand \U$28709 ( \29086 , \29084 , \29085 );
xor \U$28710 ( \29087 , \29080 , \29086 );
not \U$28711 ( \29088 , \29087 );
not \U$28712 ( \29089 , \29088 );
not \U$28713 ( \29090 , \29017 );
nand \U$28714 ( \29091 , \29058 , \29090 );
and \U$28715 ( \29092 , \29091 , \29019 );
nor \U$28716 ( \29093 , \29058 , \29090 );
nor \U$28717 ( \29094 , \29092 , \29093 );
not \U$28718 ( \29095 , \29094 );
not \U$28719 ( \29096 , \29095 );
or \U$28720 ( \29097 , \29089 , \29096 );
nand \U$28721 ( \29098 , \29094 , \29087 );
nand \U$28722 ( \29099 , \29097 , \29098 );
not \U$28723 ( \29100 , \28965 );
buf \U$28724 ( \29101 , \28998 );
not \U$28725 ( \29102 , \29101 );
or \U$28726 ( \29103 , \29100 , \29102 );
or \U$28727 ( \29104 , \29101 , \28965 );
nand \U$28728 ( \29105 , \29104 , \29007 );
nand \U$28729 ( \29106 , \29103 , \29105 );
and \U$28730 ( \29107 , \29099 , \29106 );
not \U$28731 ( \29108 , \29099 );
not \U$28732 ( \29109 , \29106 );
and \U$28733 ( \29110 , \29108 , \29109 );
nor \U$28734 ( \29111 , \29107 , \29110 );
xor \U$28735 ( \29112 , \29071 , \29111 );
not \U$28736 ( \29113 , \6689 );
not \U$28737 ( \29114 , \27837 );
or \U$28738 ( \29115 , \29113 , \29114 );
not \U$28739 ( \29116 , RIc2263e0_39);
not \U$28740 ( \29117 , \4414 );
or \U$28741 ( \29118 , \29116 , \29117 );
nand \U$28742 ( \29119 , \16519 , \5498 );
nand \U$28743 ( \29120 , \29118 , \29119 );
nand \U$28744 ( \29121 , \29120 , \6307 );
nand \U$28745 ( \29122 , \29115 , \29121 );
not \U$28746 ( \29123 , RIc226a70_25);
not \U$28747 ( \29124 , \8910 );
or \U$28748 ( \29125 , \29123 , \29124 );
not \U$28749 ( \29126 , \12403 );
nand \U$28750 ( \29127 , \29126 , \1905 );
nand \U$28751 ( \29128 , \29125 , \29127 );
and \U$28752 ( \29129 , \29128 , \2172 );
and \U$28753 ( \29130 , \27627 , \2195 );
nor \U$28754 ( \29131 , \29129 , \29130 );
xor \U$28755 ( \29132 , \29122 , \29131 );
not \U$28756 ( \29133 , \3629 );
not \U$28757 ( \29134 , \28884 );
or \U$28758 ( \29135 , \29133 , \29134 );
not \U$28759 ( \29136 , RIc2266b0_33);
not \U$28760 ( \29137 , \23758 );
or \U$28761 ( \29138 , \29136 , \29137 );
nand \U$28762 ( \29139 , \6718 , \2692 );
nand \U$28763 ( \29140 , \29138 , \29139 );
nand \U$28764 ( \29141 , \29140 , \3631 );
nand \U$28765 ( \29142 , \29135 , \29141 );
not \U$28766 ( \29143 , \29142 );
and \U$28767 ( \29144 , \29132 , \29143 );
not \U$28768 ( \29145 , \29132 );
and \U$28769 ( \29146 , \29145 , \29142 );
nor \U$28770 ( \29147 , \29144 , \29146 );
not \U$28771 ( \29148 , \29147 );
not \U$28772 ( \29149 , \29148 );
not \U$28773 ( \29150 , \2154 );
not \U$28774 ( \29151 , RIc226980_27);
not \U$28775 ( \29152 , \20367 );
or \U$28776 ( \29153 , \29151 , \29152 );
nand \U$28777 ( \29154 , \9916 , \2799 );
nand \U$28778 ( \29155 , \29153 , \29154 );
not \U$28779 ( \29156 , \29155 );
or \U$28780 ( \29157 , \29150 , \29156 );
nand \U$28781 ( \29158 , \28892 , \2138 );
nand \U$28782 ( \29159 , \29157 , \29158 );
not \U$28783 ( \29160 , \2784 );
not \U$28784 ( \29161 , \28872 );
or \U$28785 ( \29162 , \29160 , \29161 );
and \U$28786 ( \29163 , RIc226890_29, \20217 );
not \U$28787 ( \29164 , RIc226890_29);
and \U$28788 ( \29165 , \29164 , \20216 );
or \U$28789 ( \29166 , \29163 , \29165 );
nand \U$28790 ( \29167 , \29166 , \9142 );
nand \U$28791 ( \29168 , \29162 , \29167 );
xor \U$28792 ( \29169 , \29159 , \29168 );
not \U$28793 ( \29170 , \2710 );
not \U$28794 ( \29171 , RIc2267a0_31);
not \U$28795 ( \29172 , \9884 );
or \U$28796 ( \29173 , \29171 , \29172 );
nand \U$28797 ( \29174 , \8886 , \3648 );
nand \U$28798 ( \29175 , \29173 , \29174 );
not \U$28799 ( \29176 , \29175 );
or \U$28800 ( \29177 , \29170 , \29176 );
nand \U$28801 ( \29178 , \27637 , \2697 );
nand \U$28802 ( \29179 , \29177 , \29178 );
xnor \U$28803 ( \29180 , \29169 , \29179 );
not \U$28804 ( \29181 , \29180 );
not \U$28805 ( \29182 , \29181 );
or \U$28806 ( \29183 , \29149 , \29182 );
nand \U$28807 ( \29184 , \29180 , \29147 );
nand \U$28808 ( \29185 , \29183 , \29184 );
not \U$28809 ( \29186 , \9934 );
not \U$28810 ( \29187 , \28991 );
or \U$28811 ( \29188 , \29186 , \29187 );
not \U$28812 ( \29189 , RIc226110_45);
not \U$28813 ( \29190 , \3798 );
or \U$28814 ( \29191 , \29189 , \29190 );
nand \U$28815 ( \29192 , \2730 , \22795 );
nand \U$28816 ( \29193 , \29191 , \29192 );
nand \U$28817 ( \29194 , \29193 , \9398 );
nand \U$28818 ( \29195 , \29188 , \29194 );
not \U$28819 ( \29196 , \9619 );
not \U$28820 ( \29197 , RIc226020_47);
not \U$28821 ( \29198 , \3810 );
or \U$28822 ( \29199 , \29197 , \29198 );
nand \U$28823 ( \29200 , \9139 , \11607 );
nand \U$28824 ( \29201 , \29199 , \29200 );
not \U$28825 ( \29202 , \29201 );
or \U$28826 ( \29203 , \29196 , \29202 );
nand \U$28827 ( \29204 , \29026 , \10001 );
nand \U$28828 ( \29205 , \29203 , \29204 );
xor \U$28829 ( \29206 , \29195 , \29205 );
not \U$28830 ( \29207 , \11965 );
not \U$28831 ( \29208 , \29051 );
or \U$28832 ( \29209 , \29207 , \29208 );
not \U$28833 ( \29210 , RIc225b70_57);
not \U$28834 ( \29211 , \9479 );
or \U$28835 ( \29212 , \29210 , \29211 );
nand \U$28836 ( \29213 , \27761 , \15262 );
nand \U$28837 ( \29214 , \29212 , \29213 );
nand \U$28838 ( \29215 , \29214 , \15267 );
nand \U$28839 ( \29216 , \29209 , \29215 );
xor \U$28840 ( \29217 , \29206 , \29216 );
xor \U$28841 ( \29218 , \29185 , \29217 );
xor \U$28842 ( \29219 , \27821 , \27853 );
and \U$28843 ( \29220 , \29219 , \27862 );
and \U$28844 ( \29221 , \27821 , \27853 );
or \U$28845 ( \29222 , \29220 , \29221 );
not \U$28846 ( \29223 , \29222 );
xor \U$28847 ( \29224 , \29218 , \29223 );
xor \U$28848 ( \29225 , \21949 , \21958 );
not \U$28849 ( \29226 , \1310 );
not \U$28850 ( \29227 , \21115 );
or \U$28851 ( \29228 , \29226 , \29227 );
nand \U$28852 ( \29229 , \27573 , \1306 );
nand \U$28853 ( \29230 , \29228 , \29229 );
xor \U$28854 ( \29231 , \29225 , \29230 );
not \U$28855 ( \29232 , \1682 );
not \U$28856 ( \29233 , \21964 );
or \U$28857 ( \29234 , \29232 , \29233 );
nand \U$28858 ( \29235 , \27584 , \1678 );
nand \U$28859 ( \29236 , \29234 , \29235 );
xor \U$28860 ( \29237 , \29231 , \29236 );
not \U$28861 ( \29238 , \4381 );
not \U$28862 ( \29239 , \27800 );
or \U$28863 ( \29240 , \29238 , \29239 );
not \U$28864 ( \29241 , RIc2265c0_35);
not \U$28865 ( \29242 , \9765 );
or \U$28866 ( \29243 , \29241 , \29242 );
nand \U$28867 ( \29244 , \9770 , \3620 );
nand \U$28868 ( \29245 , \29243 , \29244 );
nand \U$28869 ( \29246 , \29245 , \4383 );
nand \U$28870 ( \29247 , \29240 , \29246 );
xor \U$28871 ( \29248 , \29237 , \29247 );
not \U$28872 ( \29249 , \5509 );
not \U$28873 ( \29250 , \27827 );
or \U$28874 ( \29251 , \29249 , \29250 );
not \U$28875 ( \29252 , RIc2264d0_37);
not \U$28876 ( \29253 , \10230 );
or \U$28877 ( \29254 , \29252 , \29253 );
nand \U$28878 ( \29255 , \10231 , \5514 );
nand \U$28879 ( \29256 , \29254 , \29255 );
nand \U$28880 ( \29257 , \29256 , \5519 );
nand \U$28881 ( \29258 , \29251 , \29257 );
xor \U$28882 ( \29259 , \29248 , \29258 );
not \U$28883 ( \29260 , \28996 );
not \U$28884 ( \29261 , \28971 );
or \U$28885 ( \29262 , \29260 , \29261 );
not \U$28886 ( \29263 , \28972 );
not \U$28887 ( \29264 , \28993 );
or \U$28888 ( \29265 , \29263 , \29264 );
nand \U$28889 ( \29266 , \29265 , \28978 );
nand \U$28890 ( \29267 , \29262 , \29266 );
xor \U$28891 ( \29268 , \29259 , \29267 );
not \U$28892 ( \29269 , \28957 );
not \U$28893 ( \29270 , \28963 );
or \U$28894 ( \29271 , \29269 , \29270 );
or \U$28895 ( \29272 , \28963 , \28957 );
nand \U$28896 ( \29273 , \29272 , \28952 );
nand \U$28897 ( \29274 , \29271 , \29273 );
xor \U$28898 ( \29275 , \29268 , \29274 );
not \U$28899 ( \29276 , \29275 );
and \U$28900 ( \29277 , \29224 , \29276 );
not \U$28901 ( \29278 , \29224 );
and \U$28902 ( \29279 , \29278 , \29275 );
nor \U$28903 ( \29280 , \29277 , \29279 );
xor \U$28904 ( \29281 , \29112 , \29280 );
not \U$28905 ( \29282 , \29281 );
or \U$28906 ( \29283 , \28950 , \29282 );
or \U$28907 ( \29284 , \28949 , \29281 );
nand \U$28908 ( \29285 , \29283 , \29284 );
not \U$28909 ( \29286 , \29059 );
not \U$28910 ( \29287 , \29013 );
or \U$28911 ( \29288 , \29286 , \29287 );
nand \U$28912 ( \29289 , \29060 , \29012 );
nand \U$28913 ( \29290 , \29288 , \29289 );
xor \U$28914 ( \29291 , \29290 , \29069 );
not \U$28915 ( \29292 , \29291 );
not \U$28916 ( \29293 , \26759 );
not \U$28917 ( \29294 , \26859 );
or \U$28918 ( \29295 , \29293 , \29294 );
nand \U$28919 ( \29296 , \26758 , \26716 );
nand \U$28920 ( \29297 , \29295 , \29296 );
xor \U$28921 ( \29298 , \29297 , \26857 );
xor \U$28922 ( \29299 , \28022 , \28032 );
xor \U$28923 ( \29300 , \29299 , \28043 );
xor \U$28924 ( \29301 , \28056 , \28066 );
xor \U$28925 ( \29302 , \29301 , \28077 );
xor \U$28926 ( \29303 , \29300 , \29302 );
not \U$28927 ( \29304 , \11965 );
not \U$28928 ( \29305 , RIc225b70_57);
not \U$28929 ( \29306 , \9422 );
or \U$28930 ( \29307 , \29305 , \29306 );
nand \U$28931 ( \29308 , \2590 , \10074 );
nand \U$28932 ( \29309 , \29307 , \29308 );
not \U$28933 ( \29310 , \29309 );
or \U$28934 ( \29311 , \29304 , \29310 );
nand \U$28935 ( \29312 , \27507 , \11974 );
nand \U$28936 ( \29313 , \29311 , \29312 );
not \U$28937 ( \29314 , \8777 );
not \U$28938 ( \29315 , \28516 );
or \U$28939 ( \29316 , \29314 , \29315 );
nand \U$28940 ( \29317 , \27495 , \9555 );
nand \U$28941 ( \29318 , \29316 , \29317 );
or \U$28942 ( \29319 , \29313 , \29318 );
not \U$28943 ( \29320 , \9641 );
not \U$28944 ( \29321 , \28443 );
or \U$28945 ( \29322 , \29320 , \29321 );
nand \U$28946 ( \29323 , \27531 , \12304 );
nand \U$28947 ( \29324 , \29322 , \29323 );
nand \U$28948 ( \29325 , \29319 , \29324 );
nand \U$28949 ( \29326 , \29313 , \29318 );
nand \U$28950 ( \29327 , \29325 , \29326 );
and \U$28951 ( \29328 , \29303 , \29327 );
and \U$28952 ( \29329 , \29300 , \29302 );
or \U$28953 ( \29330 , \29328 , \29329 );
or \U$28954 ( \29331 , \29298 , \29330 );
xor \U$28955 ( \29332 , \27475 , \27499 );
not \U$28956 ( \29333 , \27486 );
and \U$28957 ( \29334 , \29332 , \29333 );
not \U$28958 ( \29335 , \29332 );
and \U$28959 ( \29336 , \29335 , \27486 );
nor \U$28960 ( \29337 , \29334 , \29336 );
not \U$28961 ( \29338 , \29337 );
not \U$28962 ( \29339 , \29338 );
xor \U$28963 ( \29340 , \27511 , \27521 );
xor \U$28964 ( \29341 , \29340 , \27533 );
not \U$28965 ( \29342 , \29341 );
or \U$28966 ( \29343 , \29339 , \29342 );
or \U$28967 ( \29344 , \29341 , \29338 );
xor \U$28968 ( \29345 , \27392 , \27406 );
xnor \U$28969 ( \29346 , \29345 , \27417 );
not \U$28970 ( \29347 , \29346 );
nand \U$28971 ( \29348 , \29344 , \29347 );
nand \U$28972 ( \29349 , \29343 , \29348 );
nand \U$28973 ( \29350 , \29331 , \29349 );
nand \U$28974 ( \29351 , \29298 , \29330 );
nand \U$28975 ( \29352 , \29350 , \29351 );
xor \U$28976 ( \29353 , \26861 , \27030 );
xor \U$28977 ( \29354 , \29353 , \27198 );
xor \U$28978 ( \29355 , \29352 , \29354 );
not \U$28979 ( \29356 , \27193 );
not \U$28980 ( \29357 , \27125 );
or \U$28981 ( \29358 , \29356 , \29357 );
or \U$28982 ( \29359 , \27125 , \27193 );
nand \U$28983 ( \29360 , \29358 , \29359 );
and \U$28984 ( \29361 , \29360 , \27196 );
not \U$28985 ( \29362 , \29360 );
and \U$28986 ( \29363 , \29362 , \27084 );
nor \U$28987 ( \29364 , \29361 , \29363 );
xor \U$28988 ( \29365 , \27465 , \27501 );
xor \U$28989 ( \29366 , \29365 , \27536 );
or \U$28990 ( \29367 , \29364 , \29366 );
xor \U$28991 ( \29368 , \26825 , \26840 );
xor \U$28992 ( \29369 , \29368 , \26854 );
not \U$28993 ( \29370 , \29369 );
xor \U$28994 ( \29371 , \28094 , \28104 );
xor \U$28995 ( \29372 , \29371 , \28115 );
xor \U$28996 ( \29373 , \28213 , \28209 );
xnor \U$28997 ( \29374 , \29373 , \28198 );
or \U$28998 ( \29375 , \29372 , \29374 );
or \U$28999 ( \29376 , RIc226db8_18, RIc226d40_19);
nand \U$29000 ( \29377 , \29376 , \18182 );
and \U$29001 ( \29378 , RIc226db8_18, RIc226d40_19);
nor \U$29002 ( \29379 , \29378 , \1960 );
and \U$29003 ( \29380 , \29377 , \29379 );
not \U$29004 ( \29381 , \1963 );
not \U$29005 ( \29382 , RIc226e30_17);
not \U$29006 ( \29383 , \21102 );
or \U$29007 ( \29384 , \29382 , \29383 );
not \U$29008 ( \29385 , \16259 );
nand \U$29009 ( \29386 , \29385 , \1952 );
nand \U$29010 ( \29387 , \29384 , \29386 );
not \U$29011 ( \29388 , \29387 );
or \U$29012 ( \29389 , \29381 , \29388 );
or \U$29013 ( \29390 , \16248 , \1935 );
or \U$29014 ( \29391 , \18181 , RIc226e30_17);
nand \U$29015 ( \29392 , \29390 , \29391 );
nand \U$29016 ( \29393 , \29392 , \1944 );
nand \U$29017 ( \29394 , \29389 , \29393 );
and \U$29018 ( \29395 , \29380 , \29394 );
not \U$29019 ( \29396 , \2391 );
not \U$29020 ( \29397 , RIc226c50_21);
not \U$29021 ( \29398 , \13198 );
or \U$29022 ( \29399 , \29397 , \29398 );
nand \U$29023 ( \29400 , \12755 , \2370 );
nand \U$29024 ( \29401 , \29399 , \29400 );
not \U$29025 ( \29402 , \29401 );
or \U$29026 ( \29403 , \29396 , \29402 );
not \U$29027 ( \29404 , RIc226c50_21);
not \U$29028 ( \29405 , \21084 );
or \U$29029 ( \29406 , \29404 , \29405 );
nand \U$29030 ( \29407 , \13497 , \10834 );
nand \U$29031 ( \29408 , \29406 , \29407 );
nand \U$29032 ( \29409 , \29408 , \2367 );
nand \U$29033 ( \29410 , \29403 , \29409 );
xor \U$29034 ( \29411 , \29395 , \29410 );
not \U$29035 ( \29412 , \1930 );
not \U$29036 ( \29413 , RIc226b60_23);
not \U$29037 ( \29414 , \21172 );
or \U$29038 ( \29415 , \29413 , \29414 );
nand \U$29039 ( \29416 , \10086 , \2111 );
nand \U$29040 ( \29417 , \29415 , \29416 );
not \U$29041 ( \29418 , \29417 );
or \U$29042 ( \29419 , \29412 , \29418 );
not \U$29043 ( \29420 , RIc226b60_23);
not \U$29044 ( \29421 , \10198 );
or \U$29045 ( \29422 , \29420 , \29421 );
not \U$29046 ( \29423 , \13211 );
nand \U$29047 ( \29424 , \29423 , \2111 );
nand \U$29048 ( \29425 , \29422 , \29424 );
nand \U$29049 ( \29426 , \29425 , \1914 );
nand \U$29050 ( \29427 , \29419 , \29426 );
and \U$29051 ( \29428 , \29411 , \29427 );
and \U$29052 ( \29429 , \29395 , \29410 );
or \U$29053 ( \29430 , \29428 , \29429 );
not \U$29054 ( \29431 , \5509 );
not \U$29055 ( \29432 , RIc2264d0_37);
not \U$29056 ( \29433 , \10322 );
or \U$29057 ( \29434 , \29432 , \29433 );
nand \U$29058 ( \29435 , \8856 , \4371 );
nand \U$29059 ( \29436 , \29434 , \29435 );
not \U$29060 ( \29437 , \29436 );
or \U$29061 ( \29438 , \29431 , \29437 );
nand \U$29062 ( \29439 , \28233 , \5519 );
nand \U$29063 ( \29440 , \29438 , \29439 );
xor \U$29064 ( \29441 , \29430 , \29440 );
not \U$29065 ( \29442 , \6689 );
not \U$29066 ( \29443 , RIc2263e0_39);
not \U$29067 ( \29444 , \15699 );
or \U$29068 ( \29445 , \29443 , \29444 );
not \U$29069 ( \29446 , \10307 );
nand \U$29070 ( \29447 , \29446 , \6694 );
nand \U$29071 ( \29448 , \29445 , \29447 );
not \U$29072 ( \29449 , \29448 );
or \U$29073 ( \29450 , \29442 , \29449 );
nand \U$29074 ( \29451 , \28221 , \6307 );
nand \U$29075 ( \29452 , \29450 , \29451 );
and \U$29076 ( \29453 , \29441 , \29452 );
and \U$29077 ( \29454 , \29430 , \29440 );
or \U$29078 ( \29455 , \29453 , \29454 );
and \U$29079 ( \29456 , \29375 , \29455 );
and \U$29080 ( \29457 , \29372 , \29374 );
nor \U$29081 ( \29458 , \29456 , \29457 );
not \U$29082 ( \29459 , \29458 );
not \U$29083 ( \29460 , \29459 );
or \U$29084 ( \29461 , \29370 , \29460 );
not \U$29085 ( \29462 , \29369 );
not \U$29086 ( \29463 , \29462 );
not \U$29087 ( \29464 , \29458 );
or \U$29088 ( \29465 , \29463 , \29464 );
not \U$29089 ( \29466 , \2195 );
not \U$29090 ( \29467 , RIc226a70_25);
not \U$29091 ( \29468 , \9297 );
or \U$29092 ( \29469 , \29467 , \29468 );
nand \U$29093 ( \29470 , \9299 , \2187 );
nand \U$29094 ( \29471 , \29469 , \29470 );
not \U$29095 ( \29472 , \29471 );
or \U$29096 ( \29473 , \29466 , \29472 );
nand \U$29097 ( \29474 , \28090 , \2173 );
nand \U$29098 ( \29475 , \29473 , \29474 );
not \U$29099 ( \29476 , \29475 );
and \U$29100 ( \29477 , \28204 , \1930 );
and \U$29101 ( \29478 , \29417 , \1914 );
nor \U$29102 ( \29479 , \29477 , \29478 );
not \U$29103 ( \29480 , \29479 );
not \U$29104 ( \29481 , \29480 );
or \U$29105 ( \29482 , \29476 , \29481 );
or \U$29106 ( \29483 , \29480 , \29475 );
not \U$29107 ( \29484 , \2138 );
not \U$29108 ( \29485 , RIc226980_27);
not \U$29109 ( \29486 , \11488 );
or \U$29110 ( \29487 , \29485 , \29486 );
nand \U$29111 ( \29488 , \9256 , \2150 );
nand \U$29112 ( \29489 , \29487 , \29488 );
not \U$29113 ( \29490 , \29489 );
or \U$29114 ( \29491 , \29484 , \29490 );
nand \U$29115 ( \29492 , \28100 , \2154 );
nand \U$29116 ( \29493 , \29491 , \29492 );
nand \U$29117 ( \29494 , \29483 , \29493 );
nand \U$29118 ( \29495 , \29482 , \29494 );
not \U$29119 ( \29496 , \29495 );
and \U$29120 ( \29497 , \16248 , \2318 );
not \U$29121 ( \29498 , \1963 );
not \U$29122 ( \29499 , \28130 );
or \U$29123 ( \29500 , \29498 , \29499 );
nand \U$29124 ( \29501 , \1944 , \29387 );
nand \U$29125 ( \29502 , \29500 , \29501 );
xor \U$29126 ( \29503 , \29497 , \29502 );
not \U$29127 ( \29504 , \2517 );
not \U$29128 ( \29505 , RIc226d40_19);
not \U$29129 ( \29506 , \15629 );
or \U$29130 ( \29507 , \29505 , \29506 );
nand \U$29131 ( \29508 , \18161 , \1941 );
nand \U$29132 ( \29509 , \29507 , \29508 );
not \U$29133 ( \29510 , \29509 );
or \U$29134 ( \29511 , \29504 , \29510 );
nand \U$29135 ( \29512 , \28141 , \2533 );
nand \U$29136 ( \29513 , \29511 , \29512 );
and \U$29137 ( \29514 , \29503 , \29513 );
and \U$29138 ( \29515 , \29497 , \29502 );
or \U$29139 ( \29516 , \29514 , \29515 );
not \U$29140 ( \29517 , \2391 );
not \U$29141 ( \29518 , \29408 );
or \U$29142 ( \29519 , \29517 , \29518 );
nand \U$29143 ( \29520 , \27994 , \2367 );
nand \U$29144 ( \29521 , \29519 , \29520 );
xor \U$29145 ( \29522 , \29516 , \29521 );
not \U$29146 ( \29523 , \2078 );
and \U$29147 ( \29524 , RIc226890_29, \10652 );
not \U$29148 ( \29525 , RIc226890_29);
and \U$29149 ( \29526 , \29525 , \9072 );
or \U$29150 ( \29527 , \29524 , \29526 );
not \U$29151 ( \29528 , \29527 );
or \U$29152 ( \29529 , \29523 , \29528 );
nand \U$29153 ( \29530 , \28196 , \2086 );
nand \U$29154 ( \29531 , \29529 , \29530 );
and \U$29155 ( \29532 , \29522 , \29531 );
and \U$29156 ( \29533 , \29516 , \29521 );
or \U$29157 ( \29534 , \29532 , \29533 );
not \U$29158 ( \29535 , \29534 );
nand \U$29159 ( \29536 , \29496 , \29535 );
not \U$29160 ( \29537 , \29536 );
xor \U$29161 ( \29538 , \28122 , \28132 );
xor \U$29162 ( \29539 , \29538 , \28143 );
not \U$29163 ( \29540 , \3629 );
not \U$29164 ( \29541 , RIc2266b0_33);
not \U$29165 ( \29542 , \11094 );
or \U$29166 ( \29543 , \29541 , \29542 );
nand \U$29167 ( \29544 , \8974 , \6890 );
nand \U$29168 ( \29545 , \29543 , \29544 );
not \U$29169 ( \29546 , \29545 );
or \U$29170 ( \29547 , \29540 , \29546 );
nand \U$29171 ( \29548 , \28283 , \3631 );
nand \U$29172 ( \29549 , \29547 , \29548 );
xor \U$29173 ( \29550 , \29539 , \29549 );
not \U$29174 ( \29551 , \9690 );
not \U$29175 ( \29552 , RIc2262f0_41);
not \U$29176 ( \29553 , \22928 );
or \U$29177 ( \29554 , \29552 , \29553 );
not \U$29178 ( \29555 , \9775 );
nand \U$29179 ( \29556 , \29555 , \12937 );
nand \U$29180 ( \29557 , \29554 , \29556 );
not \U$29181 ( \29558 , \29557 );
or \U$29182 ( \29559 , \29551 , \29558 );
nand \U$29183 ( \29560 , \28246 , \9816 );
nand \U$29184 ( \29561 , \29559 , \29560 );
and \U$29185 ( \29562 , \29550 , \29561 );
and \U$29186 ( \29563 , \29539 , \29549 );
or \U$29187 ( \29564 , \29562 , \29563 );
not \U$29188 ( \29565 , \29564 );
or \U$29189 ( \29566 , \29537 , \29565 );
nand \U$29190 ( \29567 , \29495 , \29534 );
nand \U$29191 ( \29568 , \29566 , \29567 );
nand \U$29192 ( \29569 , \29465 , \29568 );
nand \U$29193 ( \29570 , \29461 , \29569 );
nand \U$29194 ( \29571 , \29367 , \29570 );
nand \U$29195 ( \29572 , \29364 , \29366 );
nand \U$29196 ( \29573 , \29571 , \29572 );
and \U$29197 ( \29574 , \29355 , \29573 );
and \U$29198 ( \29575 , \29352 , \29354 );
or \U$29199 ( \29576 , \29574 , \29575 );
not \U$29200 ( \29577 , \29576 );
or \U$29201 ( \29578 , \29292 , \29577 );
or \U$29202 ( \29579 , \29576 , \29291 );
not \U$29203 ( \29580 , \28583 );
or \U$29204 ( \29581 , \28560 , \28580 );
not \U$29205 ( \29582 , \29581 );
or \U$29206 ( \29583 , \29580 , \29582 );
nand \U$29207 ( \29584 , \28560 , \28580 );
nand \U$29208 ( \29585 , \29583 , \29584 );
nand \U$29209 ( \29586 , \29579 , \29585 );
nand \U$29210 ( \29587 , \29578 , \29586 );
not \U$29211 ( \29588 , \29587 );
and \U$29212 ( \29589 , \29285 , \29588 );
not \U$29213 ( \29590 , \29285 );
and \U$29214 ( \29591 , \29590 , \29587 );
nor \U$29215 ( \29592 , \29589 , \29591 );
not \U$29216 ( \29593 , \29592 );
and \U$29217 ( \29594 , \28941 , \29593 );
not \U$29218 ( \29595 , \28941 );
and \U$29219 ( \29596 , \29595 , \29592 );
nor \U$29220 ( \29597 , \29594 , \29596 );
xor \U$29221 ( \29598 , \29291 , \29585 );
xnor \U$29222 ( \29599 , \29598 , \29576 );
xor \U$29223 ( \29600 , \29300 , \29302 );
xor \U$29224 ( \29601 , \29600 , \29327 );
not \U$29225 ( \29602 , \29601 );
xor \U$29226 ( \29603 , \28216 , \28255 );
xor \U$29227 ( \29604 , \29603 , \28288 );
nand \U$29228 ( \29605 , \29602 , \29604 );
xor \U$29229 ( \29606 , \28370 , \28365 );
xnor \U$29230 ( \29607 , \29606 , \28329 );
and \U$29231 ( \29608 , \29605 , \29607 );
nor \U$29232 ( \29609 , \29602 , \29604 );
nor \U$29233 ( \29610 , \29608 , \29609 );
xor \U$29234 ( \29611 , \29330 , \29349 );
xnor \U$29235 ( \29612 , \29611 , \29298 );
xor \U$29236 ( \29613 , \29610 , \29612 );
not \U$29237 ( \29614 , \29337 );
not \U$29238 ( \29615 , \29614 );
not \U$29239 ( \29616 , \29346 );
or \U$29240 ( \29617 , \29615 , \29616 );
or \U$29241 ( \29618 , \29338 , \29346 );
nand \U$29242 ( \29619 , \29617 , \29618 );
not \U$29243 ( \29620 , \29341 );
and \U$29244 ( \29621 , \29619 , \29620 );
not \U$29245 ( \29622 , \29619 );
and \U$29246 ( \29623 , \29622 , \29341 );
nor \U$29247 ( \29624 , \29621 , \29623 );
not \U$29248 ( \29625 , \29624 );
not \U$29249 ( \29626 , \5135 );
not \U$29250 ( \29627 , \28153 );
or \U$29251 ( \29628 , \29626 , \29627 );
not \U$29252 ( \29629 , RIc2265c0_35);
not \U$29253 ( \29630 , \15684 );
or \U$29254 ( \29631 , \29629 , \29630 );
nand \U$29255 ( \29632 , \8806 , \16314 );
nand \U$29256 ( \29633 , \29631 , \29632 );
nand \U$29257 ( \29634 , \29633 , \4381 );
nand \U$29258 ( \29635 , \29628 , \29634 );
not \U$29259 ( \29636 , \11965 );
not \U$29260 ( \29637 , RIc225b70_57);
not \U$29261 ( \29638 , \4803 );
or \U$29262 ( \29639 , \29637 , \29638 );
nand \U$29263 ( \29640 , \9364 , \12475 );
nand \U$29264 ( \29641 , \29639 , \29640 );
not \U$29265 ( \29642 , \29641 );
or \U$29266 ( \29643 , \29636 , \29642 );
nand \U$29267 ( \29644 , \29309 , \11974 );
nand \U$29268 ( \29645 , \29643 , \29644 );
xor \U$29269 ( \29646 , \29635 , \29645 );
not \U$29270 ( \29647 , \9534 );
not \U$29271 ( \29648 , RIc225f30_49);
not \U$29272 ( \29649 , \9513 );
or \U$29273 ( \29650 , \29648 , \29649 );
nand \U$29274 ( \29651 , \11324 , \9549 );
nand \U$29275 ( \29652 , \29650 , \29651 );
not \U$29276 ( \29653 , \29652 );
or \U$29277 ( \29654 , \29647 , \29653 );
nand \U$29278 ( \29655 , \28165 , \9552 );
nand \U$29279 ( \29656 , \29654 , \29655 );
and \U$29280 ( \29657 , \29646 , \29656 );
and \U$29281 ( \29658 , \29635 , \29645 );
or \U$29282 ( \29659 , \29657 , \29658 );
not \U$29283 ( \29660 , \29659 );
and \U$29284 ( \29661 , \28363 , \28348 );
not \U$29285 ( \29662 , \28363 );
and \U$29286 ( \29663 , \29662 , \28349 );
or \U$29287 ( \29664 , \29661 , \29663 );
and \U$29288 ( \29665 , \29664 , \28339 );
not \U$29289 ( \29666 , \29664 );
and \U$29290 ( \29667 , \29666 , \28340 );
nor \U$29291 ( \29668 , \29665 , \29667 );
nand \U$29292 ( \29669 , \29660 , \29668 );
xor \U$29293 ( \29670 , \29516 , \29521 );
xor \U$29294 ( \29671 , \29670 , \29531 );
xor \U$29295 ( \29672 , \29497 , \29502 );
xor \U$29296 ( \29673 , \29672 , \29513 );
not \U$29297 ( \29674 , \2173 );
not \U$29298 ( \29675 , \29471 );
or \U$29299 ( \29676 , \29674 , \29675 );
not \U$29300 ( \29677 , RIc226a70_25);
not \U$29301 ( \29678 , \12100 );
or \U$29302 ( \29679 , \29677 , \29678 );
nand \U$29303 ( \29680 , \9324 , \2190 );
nand \U$29304 ( \29681 , \29679 , \29680 );
nand \U$29305 ( \29682 , \29681 , \2195 );
nand \U$29306 ( \29683 , \29676 , \29682 );
xor \U$29307 ( \29684 , \29673 , \29683 );
not \U$29308 ( \29685 , \2154 );
not \U$29309 ( \29686 , \29489 );
or \U$29310 ( \29687 , \29685 , \29686 );
not \U$29311 ( \29688 , RIc226980_27);
not \U$29312 ( \29689 , \9274 );
not \U$29313 ( \29690 , \29689 );
or \U$29314 ( \29691 , \29688 , \29690 );
nand \U$29315 ( \29692 , \10976 , \4528 );
nand \U$29316 ( \29693 , \29691 , \29692 );
nand \U$29317 ( \29694 , \29693 , \2138 );
nand \U$29318 ( \29695 , \29687 , \29694 );
and \U$29319 ( \29696 , \29684 , \29695 );
and \U$29320 ( \29697 , \29673 , \29683 );
or \U$29321 ( \29698 , \29696 , \29697 );
xor \U$29322 ( \29699 , \29671 , \29698 );
not \U$29323 ( \29700 , \9459 );
not \U$29324 ( \29701 , RIc225e40_51);
not \U$29325 ( \29702 , \9188 );
or \U$29326 ( \29703 , \29701 , \29702 );
nand \U$29327 ( \29704 , \9805 , \12423 );
nand \U$29328 ( \29705 , \29703 , \29704 );
not \U$29329 ( \29706 , \29705 );
or \U$29330 ( \29707 , \29700 , \29706 );
nand \U$29331 ( \29708 , \28320 , \9444 );
nand \U$29332 ( \29709 , \29707 , \29708 );
and \U$29333 ( \29710 , \29699 , \29709 );
and \U$29334 ( \29711 , \29671 , \29698 );
or \U$29335 ( \29712 , \29710 , \29711 );
and \U$29336 ( \29713 , \29669 , \29712 );
not \U$29337 ( \29714 , \29659 );
nor \U$29338 ( \29715 , \29714 , \29668 );
nor \U$29339 ( \29716 , \29713 , \29715 );
not \U$29340 ( \29717 , \29716 );
or \U$29341 ( \29718 , \29625 , \29717 );
xor \U$29342 ( \29719 , \28326 , \28322 );
xnor \U$29343 ( \29720 , \29719 , \28312 );
xor \U$29344 ( \29721 , \29318 , \29313 );
xor \U$29345 ( \29722 , \29721 , \29324 );
xor \U$29346 ( \29723 , \29720 , \29722 );
and \U$29347 ( \29724 , \29493 , \29479 );
not \U$29348 ( \29725 , \29493 );
and \U$29349 ( \29726 , \29725 , \29480 );
nor \U$29350 ( \29727 , \29724 , \29726 );
xor \U$29351 ( \29728 , \29727 , \29475 );
not \U$29352 ( \29729 , \6071 );
not \U$29353 ( \29730 , \12456 );
and \U$29354 ( \29731 , \29729 , \29730 );
and \U$29355 ( \29732 , \23772 , \9125 );
nor \U$29356 ( \29733 , \29731 , \29732 );
not \U$29357 ( \29734 , \29733 );
not \U$29358 ( \29735 , \9109 );
and \U$29359 ( \29736 , \29734 , \29735 );
and \U$29360 ( \29737 , \28477 , \9129 );
nor \U$29361 ( \29738 , \29736 , \29737 );
not \U$29362 ( \29739 , \9382 );
not \U$29363 ( \29740 , RIc226110_45);
not \U$29364 ( \29741 , \9754 );
or \U$29365 ( \29742 , \29740 , \29741 );
nand \U$29366 ( \29743 , \5215 , \9379 );
nand \U$29367 ( \29744 , \29742 , \29743 );
not \U$29368 ( \29745 , \29744 );
or \U$29369 ( \29746 , \29739 , \29745 );
nand \U$29370 ( \29747 , \28497 , \11825 );
nand \U$29371 ( \29748 , \29746 , \29747 );
not \U$29372 ( \29749 , \29748 );
nand \U$29373 ( \29750 , \29738 , \29749 );
not \U$29374 ( \29751 , \9639 );
not \U$29375 ( \29752 , RIc226020_47);
not \U$29376 ( \29753 , \4414 );
or \U$29377 ( \29754 , \29752 , \29753 );
nand \U$29378 ( \29755 , \16519 , \11607 );
nand \U$29379 ( \29756 , \29754 , \29755 );
not \U$29380 ( \29757 , \29756 );
or \U$29381 ( \29758 , \29751 , \29757 );
nand \U$29382 ( \29759 , \28434 , \9619 );
nand \U$29383 ( \29760 , \29758 , \29759 );
and \U$29384 ( \29761 , \29750 , \29760 );
nor \U$29385 ( \29762 , \29738 , \29749 );
nor \U$29386 ( \29763 , \29761 , \29762 );
or \U$29387 ( \29764 , \29728 , \29763 );
not \U$29388 ( \29765 , \29728 );
not \U$29389 ( \29766 , \29763 );
or \U$29390 ( \29767 , \29765 , \29766 );
xor \U$29391 ( \29768 , \29380 , \29394 );
not \U$29392 ( \29769 , \2533 );
not \U$29393 ( \29770 , \29509 );
or \U$29394 ( \29771 , \29769 , \29770 );
not \U$29395 ( \29772 , RIc226d40_19);
not \U$29396 ( \29773 , \21094 );
or \U$29397 ( \29774 , \29772 , \29773 );
nand \U$29398 ( \29775 , \13487 , \1941 );
nand \U$29399 ( \29776 , \29774 , \29775 );
nand \U$29400 ( \29777 , \29776 , \2518 );
nand \U$29401 ( \29778 , \29771 , \29777 );
xor \U$29402 ( \29779 , \29768 , \29778 );
not \U$29403 ( \29780 , \1930 );
not \U$29404 ( \29781 , \29425 );
or \U$29405 ( \29782 , \29780 , \29781 );
not \U$29406 ( \29783 , RIc226b60_23);
not \U$29407 ( \29784 , \17625 );
or \U$29408 ( \29785 , \29783 , \29784 );
nand \U$29409 ( \29786 , \10356 , \1927 );
nand \U$29410 ( \29787 , \29785 , \29786 );
nand \U$29411 ( \29788 , \29787 , \1914 );
nand \U$29412 ( \29789 , \29782 , \29788 );
and \U$29413 ( \29790 , \29779 , \29789 );
and \U$29414 ( \29791 , \29768 , \29778 );
or \U$29415 ( \29792 , \29790 , \29791 );
not \U$29416 ( \29793 , \6307 );
not \U$29417 ( \29794 , \29448 );
or \U$29418 ( \29795 , \29793 , \29794 );
not \U$29419 ( \29796 , RIc2263e0_39);
not \U$29420 ( \29797 , \17579 );
or \U$29421 ( \29798 , \29796 , \29797 );
nand \U$29422 ( \29799 , \8886 , \8998 );
nand \U$29423 ( \29800 , \29798 , \29799 );
nand \U$29424 ( \29801 , \29800 , \6688 );
nand \U$29425 ( \29802 , \29795 , \29801 );
xor \U$29426 ( \29803 , \29792 , \29802 );
not \U$29427 ( \29804 , \9690 );
not \U$29428 ( \29805 , RIc2262f0_41);
not \U$29429 ( \29806 , \21438 );
or \U$29430 ( \29807 , \29805 , \29806 );
nand \U$29431 ( \29808 , \6720 , \12937 );
nand \U$29432 ( \29809 , \29807 , \29808 );
not \U$29433 ( \29810 , \29809 );
or \U$29434 ( \29811 , \29804 , \29810 );
nand \U$29435 ( \29812 , \29557 , \9816 );
nand \U$29436 ( \29813 , \29811 , \29812 );
and \U$29437 ( \29814 , \29803 , \29813 );
and \U$29438 ( \29815 , \29792 , \29802 );
or \U$29439 ( \29816 , \29814 , \29815 );
nand \U$29440 ( \29817 , \29767 , \29816 );
nand \U$29441 ( \29818 , \29764 , \29817 );
and \U$29442 ( \29819 , \29723 , \29818 );
and \U$29443 ( \29820 , \29720 , \29722 );
or \U$29444 ( \29821 , \29819 , \29820 );
nand \U$29445 ( \29822 , \29718 , \29821 );
not \U$29446 ( \29823 , \29716 );
not \U$29447 ( \29824 , \29624 );
nand \U$29448 ( \29825 , \29823 , \29824 );
and \U$29449 ( \29826 , \29822 , \29825 );
and \U$29450 ( \29827 , \29613 , \29826 );
and \U$29451 ( \29828 , \29610 , \29612 );
or \U$29452 ( \29829 , \29827 , \29828 );
not \U$29453 ( \29830 , \29829 );
xor \U$29454 ( \29831 , \29352 , \29354 );
xor \U$29455 ( \29832 , \29831 , \29573 );
nor \U$29456 ( \29833 , \29830 , \29832 );
xor \U$29457 ( \29834 , \28545 , \28379 );
not \U$29458 ( \29835 , \28383 );
and \U$29459 ( \29836 , \29834 , \29835 );
not \U$29460 ( \29837 , \29834 );
and \U$29461 ( \29838 , \29837 , \28383 );
nor \U$29462 ( \29839 , \29836 , \29838 );
xor \U$29463 ( \29840 , \29570 , \29366 );
not \U$29464 ( \29841 , \29364 );
and \U$29465 ( \29842 , \29840 , \29841 );
not \U$29466 ( \29843 , \29840 );
and \U$29467 ( \29844 , \29843 , \29364 );
nor \U$29468 ( \29845 , \29842 , \29844 );
nand \U$29469 ( \29846 , \29839 , \29845 );
and \U$29470 ( \29847 , \29568 , \29462 );
not \U$29471 ( \29848 , \29568 );
and \U$29472 ( \29849 , \29848 , \29369 );
nor \U$29473 ( \29850 , \29847 , \29849 );
xor \U$29474 ( \29851 , \29850 , \29459 );
not \U$29475 ( \29852 , \29851 );
not \U$29476 ( \29853 , \29852 );
xor \U$29477 ( \29854 , \29495 , \29535 );
xnor \U$29478 ( \29855 , \29854 , \29564 );
xor \U$29479 ( \29856 , \29374 , \29372 );
xor \U$29480 ( \29857 , \29856 , \29455 );
xor \U$29481 ( \29858 , \29855 , \29857 );
xor \U$29482 ( \29859 , \29430 , \29440 );
xor \U$29483 ( \29860 , \29859 , \29452 );
xor \U$29484 ( \29861 , \29539 , \29549 );
xor \U$29485 ( \29862 , \29861 , \29561 );
xor \U$29486 ( \29863 , \29860 , \29862 );
not \U$29487 ( \29864 , \28507 );
not \U$29488 ( \29865 , \29864 );
not \U$29489 ( \29866 , \20862 );
not \U$29490 ( \29867 , \29866 );
and \U$29491 ( \29868 , \29865 , \29867 );
and \U$29492 ( \29869 , \12806 , \1989 );
not \U$29493 ( \29870 , \12806 );
and \U$29494 ( \29871 , \29870 , \3838 );
or \U$29495 ( \29872 , \29869 , \29871 );
not \U$29496 ( \29873 , \29872 );
and \U$29497 ( \29874 , \29873 , \15719 );
nor \U$29498 ( \29875 , \29868 , \29874 );
not \U$29499 ( \29876 , \29875 );
not \U$29500 ( \29877 , \11974 );
not \U$29501 ( \29878 , \29641 );
or \U$29502 ( \29879 , \29877 , \29878 );
not \U$29503 ( \29880 , RIc225b70_57);
not \U$29504 ( \29881 , \28706 );
or \U$29505 ( \29882 , \29880 , \29881 );
nand \U$29506 ( \29883 , \17819 , \10074 );
nand \U$29507 ( \29884 , \29882 , \29883 );
nand \U$29508 ( \29885 , \29884 , \11965 );
nand \U$29509 ( \29886 , \29879 , \29885 );
not \U$29510 ( \29887 , \29886 );
not \U$29511 ( \29888 , \29887 );
or \U$29512 ( \29889 , \29876 , \29888 );
not \U$29513 ( \29890 , \12532 );
not \U$29514 ( \29891 , \28453 );
or \U$29515 ( \29892 , \29890 , \29891 );
not \U$29516 ( \29893 , RIc225c60_55);
not \U$29517 ( \29894 , \2670 );
or \U$29518 ( \29895 , \29893 , \29894 );
nand \U$29519 ( \29896 , \16642 , \11108 );
nand \U$29520 ( \29897 , \29895 , \29896 );
nand \U$29521 ( \29898 , \29897 , \11117 );
nand \U$29522 ( \29899 , \29892 , \29898 );
nand \U$29523 ( \29900 , \29889 , \29899 );
not \U$29524 ( \29901 , \29875 );
nand \U$29525 ( \29902 , \29901 , \29886 );
nand \U$29526 ( \29903 , \29900 , \29902 );
and \U$29527 ( \29904 , \29863 , \29903 );
and \U$29528 ( \29905 , \29860 , \29862 );
or \U$29529 ( \29906 , \29904 , \29905 );
and \U$29530 ( \29907 , \29858 , \29906 );
and \U$29531 ( \29908 , \29855 , \29857 );
or \U$29532 ( \29909 , \29907 , \29908 );
not \U$29533 ( \29910 , \29909 );
or \U$29534 ( \29911 , \29853 , \29910 );
not \U$29535 ( \29912 , \29851 );
not \U$29536 ( \29913 , \29909 );
not \U$29537 ( \29914 , \29913 );
or \U$29538 ( \29915 , \29912 , \29914 );
not \U$29539 ( \29916 , \2078 );
and \U$29540 ( \29917 , RIc226890_29, \10111 );
not \U$29541 ( \29918 , RIc226890_29);
and \U$29542 ( \29919 , \29918 , \10110 );
or \U$29543 ( \29920 , \29917 , \29919 );
not \U$29544 ( \29921 , \29920 );
or \U$29545 ( \29922 , \29916 , \29921 );
nand \U$29546 ( \29923 , \29527 , \9142 );
nand \U$29547 ( \29924 , \29922 , \29923 );
not \U$29548 ( \29925 , \2710 );
not \U$29549 ( \29926 , \28486 );
or \U$29550 ( \29927 , \29925 , \29926 );
not \U$29551 ( \29928 , RIc2267a0_31);
not \U$29552 ( \29929 , \10645 );
or \U$29553 ( \29930 , \29928 , \29929 );
nand \U$29554 ( \29931 , \9225 , \3648 );
nand \U$29555 ( \29932 , \29930 , \29931 );
nand \U$29556 ( \29933 , \29932 , \2697 );
nand \U$29557 ( \29934 , \29927 , \29933 );
xor \U$29558 ( \29935 , \29924 , \29934 );
not \U$29559 ( \29936 , \3631 );
not \U$29560 ( \29937 , \29545 );
or \U$29561 ( \29938 , \29936 , \29937 );
not \U$29562 ( \29939 , \2692 );
not \U$29563 ( \29940 , \14968 );
or \U$29564 ( \29941 , \29939 , \29940 );
not \U$29565 ( \29942 , \8913 );
nand \U$29566 ( \29943 , \29942 , RIc2266b0_33);
nand \U$29567 ( \29944 , \29941 , \29943 );
nand \U$29568 ( \29945 , \29944 , \3629 );
nand \U$29569 ( \29946 , \29938 , \29945 );
and \U$29570 ( \29947 , \29935 , \29946 );
and \U$29571 ( \29948 , \29924 , \29934 );
or \U$29572 ( \29949 , \29947 , \29948 );
not \U$29573 ( \29950 , \29949 );
not \U$29574 ( \29951 , \4381 );
not \U$29575 ( \29952 , RIc2265c0_35);
not \U$29576 ( \29953 , \9915 );
or \U$29577 ( \29954 , \29952 , \29953 );
nand \U$29578 ( \29955 , \8951 , \3620 );
nand \U$29579 ( \29956 , \29954 , \29955 );
not \U$29580 ( \29957 , \29956 );
or \U$29581 ( \29958 , \29951 , \29957 );
nand \U$29582 ( \29959 , \29633 , \4383 );
nand \U$29583 ( \29960 , \29958 , \29959 );
not \U$29584 ( \29961 , \29960 );
not \U$29585 ( \29962 , \5509 );
not \U$29586 ( \29963 , RIc2264d0_37);
not \U$29587 ( \29964 , \9897 );
or \U$29588 ( \29965 , \29963 , \29964 );
nand \U$29589 ( \29966 , \8831 , \4371 );
nand \U$29590 ( \29967 , \29965 , \29966 );
not \U$29591 ( \29968 , \29967 );
or \U$29592 ( \29969 , \29962 , \29968 );
nand \U$29593 ( \29970 , \29436 , \5519 );
nand \U$29594 ( \29971 , \29969 , \29970 );
not \U$29595 ( \29972 , \29971 );
nand \U$29596 ( \29973 , \29961 , \29972 );
not \U$29597 ( \29974 , \29973 );
not \U$29598 ( \29975 , \9552 );
not \U$29599 ( \29976 , \29652 );
or \U$29600 ( \29977 , \29975 , \29976 );
not \U$29601 ( \29978 , RIc225f30_49);
not \U$29602 ( \29979 , \3726 );
or \U$29603 ( \29980 , \29978 , \29979 );
nand \U$29604 ( \29981 , \2980 , \9541 );
nand \U$29605 ( \29982 , \29980 , \29981 );
nand \U$29606 ( \29983 , \29982 , \9532 );
nand \U$29607 ( \29984 , \29977 , \29983 );
not \U$29608 ( \29985 , \29984 );
or \U$29609 ( \29986 , \29974 , \29985 );
nand \U$29610 ( \29987 , \29971 , \29960 );
nand \U$29611 ( \29988 , \29986 , \29987 );
not \U$29612 ( \29989 , \29988 );
or \U$29613 ( \29990 , \29950 , \29989 );
or \U$29614 ( \29991 , \29988 , \29949 );
not \U$29615 ( \29992 , \8777 );
not \U$29616 ( \29993 , RIc225d50_53);
not \U$29617 ( \29994 , \3798 );
or \U$29618 ( \29995 , \29993 , \29994 );
nand \U$29619 ( \29996 , \2042 , \11391 );
nand \U$29620 ( \29997 , \29995 , \29996 );
not \U$29621 ( \29998 , \29997 );
or \U$29622 ( \29999 , \29992 , \29998 );
nand \U$29623 ( \30000 , \28522 , \9555 );
nand \U$29624 ( \30001 , \29999 , \30000 );
not \U$29625 ( \30002 , \30001 );
not \U$29626 ( \30003 , RIc225828_64);
not \U$29627 ( \30004 , \28423 );
or \U$29628 ( \30005 , \30003 , \30004 );
not \U$29629 ( \30006 , RIc2258a0_63);
not \U$29630 ( \30007 , \19226 );
or \U$29631 ( \30008 , \30006 , \30007 );
nand \U$29632 ( \30009 , \11648 , \15620 );
nand \U$29633 ( \30010 , \30008 , \30009 );
nand \U$29634 ( \30011 , \30010 , \16891 );
nand \U$29635 ( \30012 , \30005 , \30011 );
not \U$29636 ( \30013 , \30012 );
or \U$29637 ( \30014 , \30002 , \30013 );
or \U$29638 ( \30015 , \30012 , \30001 );
xor \U$29639 ( \30016 , \29395 , \29410 );
xor \U$29640 ( \30017 , \30016 , \29427 );
nand \U$29641 ( \30018 , \30015 , \30017 );
nand \U$29642 ( \30019 , \30014 , \30018 );
nand \U$29643 ( \30020 , \29991 , \30019 );
nand \U$29644 ( \30021 , \29990 , \30020 );
not \U$29645 ( \30022 , \30021 );
xor \U$29646 ( \30023 , \28479 , \28488 );
xor \U$29647 ( \30024 , \30023 , \28499 );
not \U$29648 ( \30025 , \30024 );
xor \U$29649 ( \30026 , \28511 , \28524 );
xor \U$29650 ( \30027 , \30026 , \28534 );
not \U$29651 ( \30028 , \30027 );
or \U$29652 ( \30029 , \30025 , \30028 );
or \U$29653 ( \30030 , \30027 , \30024 );
not \U$29654 ( \30031 , \2367 );
not \U$29655 ( \30032 , \29401 );
or \U$29656 ( \30033 , \30031 , \30032 );
not \U$29657 ( \30034 , RIc226c50_21);
not \U$29658 ( \30035 , \18167 );
or \U$29659 ( \30036 , \30034 , \30035 );
nand \U$29660 ( \30037 , \19721 , \3204 );
nand \U$29661 ( \30038 , \30036 , \30037 );
nand \U$29662 ( \30039 , \30038 , \2392 );
nand \U$29663 ( \30040 , \30033 , \30039 );
and \U$29664 ( \30041 , \16248 , \1963 );
not \U$29665 ( \30042 , \2533 );
not \U$29666 ( \30043 , \29776 );
or \U$29667 ( \30044 , \30042 , \30043 );
not \U$29668 ( \30045 , RIc226d40_19);
not \U$29669 ( \30046 , \20528 );
or \U$29670 ( \30047 , \30045 , \30046 );
nand \U$29671 ( \30048 , \16482 , \1941 );
nand \U$29672 ( \30049 , \30047 , \30048 );
nand \U$29673 ( \30050 , \30049 , \2517 );
nand \U$29674 ( \30051 , \30044 , \30050 );
xor \U$29675 ( \30052 , \30041 , \30051 );
not \U$29676 ( \30053 , \2391 );
not \U$29677 ( \30054 , RIc226c50_21);
not \U$29678 ( \30055 , \15630 );
or \U$29679 ( \30056 , \30054 , \30055 );
nand \U$29680 ( \30057 , \12845 , \10834 );
nand \U$29681 ( \30058 , \30056 , \30057 );
not \U$29682 ( \30059 , \30058 );
or \U$29683 ( \30060 , \30053 , \30059 );
nand \U$29684 ( \30061 , \30038 , \2367 );
nand \U$29685 ( \30062 , \30060 , \30061 );
and \U$29686 ( \30063 , \30052 , \30062 );
and \U$29687 ( \30064 , \30041 , \30051 );
or \U$29688 ( \30065 , \30063 , \30064 );
xor \U$29689 ( \30066 , \30040 , \30065 );
not \U$29690 ( \30067 , \2138 );
not \U$29691 ( \30068 , RIc226980_27);
buf \U$29692 ( \30069 , \10263 );
not \U$29693 ( \30070 , \30069 );
or \U$29694 ( \30071 , \30068 , \30070 );
nand \U$29695 ( \30072 , \9299 , \2150 );
nand \U$29696 ( \30073 , \30071 , \30072 );
not \U$29697 ( \30074 , \30073 );
or \U$29698 ( \30075 , \30067 , \30074 );
nand \U$29699 ( \30076 , \29693 , \2154 );
nand \U$29700 ( \30077 , \30075 , \30076 );
and \U$29701 ( \30078 , \30066 , \30077 );
and \U$29702 ( \30079 , \30040 , \30065 );
or \U$29703 ( \30080 , \30078 , \30079 );
not \U$29704 ( \30081 , \12670 );
not \U$29705 ( \30082 , \28530 );
or \U$29706 ( \30083 , \30081 , \30082 );
not \U$29707 ( \30084 , RIc225a80_59);
not \U$29708 ( \30085 , \2592 );
or \U$29709 ( \30086 , \30084 , \30085 );
not \U$29710 ( \30087 , RIc225a80_59);
nand \U$29711 ( \30088 , \30087 , \3291 );
nand \U$29712 ( \30089 , \30086 , \30088 );
nand \U$29713 ( \30090 , \30089 , \15164 );
nand \U$29714 ( \30091 , \30083 , \30090 );
xor \U$29715 ( \30092 , \30080 , \30091 );
not \U$29716 ( \30093 , \9459 );
not \U$29717 ( \30094 , RIc225e40_51);
not \U$29718 ( \30095 , \2104 );
or \U$29719 ( \30096 , \30094 , \30095 );
nand \U$29720 ( \30097 , \4501 , \9450 );
nand \U$29721 ( \30098 , \30096 , \30097 );
not \U$29722 ( \30099 , \30098 );
or \U$29723 ( \30100 , \30093 , \30099 );
nand \U$29724 ( \30101 , \29705 , \9445 );
nand \U$29725 ( \30102 , \30100 , \30101 );
and \U$29726 ( \30103 , \30092 , \30102 );
and \U$29727 ( \30104 , \30080 , \30091 );
or \U$29728 ( \30105 , \30103 , \30104 );
nand \U$29729 ( \30106 , \30030 , \30105 );
nand \U$29730 ( \30107 , \30029 , \30106 );
not \U$29731 ( \30108 , \30107 );
or \U$29732 ( \30109 , \30022 , \30108 );
or \U$29733 ( \30110 , \30107 , \30021 );
not \U$29734 ( \30111 , \28400 );
not \U$29735 ( \30112 , \28415 );
or \U$29736 ( \30113 , \30111 , \30112 );
nand \U$29737 ( \30114 , \28411 , \28399 );
nand \U$29738 ( \30115 , \30113 , \30114 );
and \U$29739 ( \30116 , \30115 , \28461 );
not \U$29740 ( \30117 , \30115 );
not \U$29741 ( \30118 , \28461 );
and \U$29742 ( \30119 , \30117 , \30118 );
nor \U$29743 ( \30120 , \30116 , \30119 );
nand \U$29744 ( \30121 , \30110 , \30120 );
nand \U$29745 ( \30122 , \30109 , \30121 );
nand \U$29746 ( \30123 , \29915 , \30122 );
nand \U$29747 ( \30124 , \29911 , \30123 );
and \U$29748 ( \30125 , \29846 , \30124 );
nor \U$29749 ( \30126 , \29839 , \29845 );
nor \U$29750 ( \30127 , \30125 , \30126 );
or \U$29751 ( \30128 , \29833 , \30127 );
not \U$29752 ( \30129 , \29829 );
nand \U$29753 ( \30130 , \30129 , \29832 );
nand \U$29754 ( \30131 , \30128 , \30130 );
not \U$29755 ( \30132 , \30131 );
xor \U$29756 ( \30133 , \29599 , \30132 );
xor \U$29757 ( \30134 , \27566 , \28186 );
xnor \U$29758 ( \30135 , \30134 , \28588 );
and \U$29759 ( \30136 , \30133 , \30135 );
and \U$29760 ( \30137 , \29599 , \30132 );
or \U$29761 ( \30138 , \30136 , \30137 );
nand \U$29762 ( \30139 , \29597 , \30138 );
buf \U$29763 ( \30140 , \30139 );
not \U$29764 ( \30141 , \30140 );
xor \U$29765 ( \30142 , \29599 , \30132 );
xor \U$29766 ( \30143 , \30142 , \30135 );
and \U$29767 ( \30144 , \28547 , \28550 );
not \U$29768 ( \30145 , \28547 );
and \U$29769 ( \30146 , \30145 , \28551 );
nor \U$29770 ( \30147 , \30144 , \30146 );
xnor \U$29771 ( \30148 , \30147 , \28584 );
xor \U$29772 ( \30149 , \29610 , \29612 );
xor \U$29773 ( \30150 , \30149 , \29826 );
xor \U$29774 ( \30151 , \29604 , \29601 );
xnor \U$29775 ( \30152 , \30151 , \29607 );
not \U$29776 ( \30153 , \28396 );
not \U$29777 ( \30154 , \28467 );
or \U$29778 ( \30155 , \30153 , \30154 );
nand \U$29779 ( \30156 , \28463 , \28395 );
nand \U$29780 ( \30157 , \30155 , \30156 );
and \U$29781 ( \30158 , \30157 , \28543 );
not \U$29782 ( \30159 , \30157 );
not \U$29783 ( \30160 , \28543 );
and \U$29784 ( \30161 , \30159 , \30160 );
nor \U$29785 ( \30162 , \30158 , \30161 );
xor \U$29786 ( \30163 , \30152 , \30162 );
xor \U$29787 ( \30164 , \28502 , \28537 );
xor \U$29788 ( \30165 , \30164 , \28540 );
xor \U$29789 ( \30166 , \29635 , \29645 );
xor \U$29790 ( \30167 , \30166 , \29656 );
not \U$29791 ( \30168 , \30167 );
not \U$29792 ( \30169 , \28459 );
not \U$29793 ( \30170 , \28457 );
not \U$29794 ( \30171 , \30170 );
or \U$29795 ( \30172 , \30169 , \30171 );
nand \U$29796 ( \30173 , \28457 , \28445 );
nand \U$29797 ( \30174 , \30172 , \30173 );
and \U$29798 ( \30175 , \30174 , \28428 );
not \U$29799 ( \30176 , \30174 );
and \U$29800 ( \30177 , \30176 , \28427 );
nor \U$29801 ( \30178 , \30175 , \30177 );
not \U$29802 ( \30179 , \30178 );
not \U$29803 ( \30180 , \30179 );
or \U$29804 ( \30181 , \30168 , \30180 );
not \U$29805 ( \30182 , \30167 );
not \U$29806 ( \30183 , \30182 );
not \U$29807 ( \30184 , \30178 );
or \U$29808 ( \30185 , \30183 , \30184 );
xor \U$29809 ( \30186 , \29671 , \29698 );
xor \U$29810 ( \30187 , \30186 , \29709 );
nand \U$29811 ( \30188 , \30185 , \30187 );
nand \U$29812 ( \30189 , \30181 , \30188 );
xor \U$29813 ( \30190 , \30165 , \30189 );
xor \U$29814 ( \30191 , \29720 , \29722 );
xor \U$29815 ( \30192 , \30191 , \29818 );
and \U$29816 ( \30193 , \30190 , \30192 );
and \U$29817 ( \30194 , \30165 , \30189 );
or \U$29818 ( \30195 , \30193 , \30194 );
and \U$29819 ( \30196 , \30163 , \30195 );
and \U$29820 ( \30197 , \30152 , \30162 );
or \U$29821 ( \30198 , \30196 , \30197 );
not \U$29822 ( \30199 , \30198 );
nand \U$29823 ( \30200 , \30150 , \30199 );
not \U$29824 ( \30201 , \30200 );
xor \U$29825 ( \30202 , \29851 , \30122 );
xor \U$29826 ( \30203 , \30202 , \29909 );
not \U$29827 ( \30204 , \30203 );
not \U$29828 ( \30205 , \30204 );
xor \U$29829 ( \30206 , \29716 , \29821 );
buf \U$29830 ( \30207 , \29624 );
xnor \U$29831 ( \30208 , \30206 , \30207 );
not \U$29832 ( \30209 , \30208 );
not \U$29833 ( \30210 , \30209 );
or \U$29834 ( \30211 , \30205 , \30210 );
not \U$29835 ( \30212 , \30208 );
not \U$29836 ( \30213 , \30203 );
or \U$29837 ( \30214 , \30212 , \30213 );
xor \U$29838 ( \30215 , \29712 , \29659 );
xnor \U$29839 ( \30216 , \30215 , \29668 );
not \U$29840 ( \30217 , \30216 );
not \U$29841 ( \30218 , RIc225828_64);
not \U$29842 ( \30219 , \30010 );
or \U$29843 ( \30220 , \30218 , \30219 );
not \U$29844 ( \30221 , RIc2258a0_63);
not \U$29845 ( \30222 , \4009 );
or \U$29846 ( \30223 , \30221 , \30222 );
nand \U$29847 ( \30224 , \9608 , \28750 );
nand \U$29848 ( \30225 , \30223 , \30224 );
nand \U$29849 ( \30226 , \30225 , \16891 );
nand \U$29850 ( \30227 , \30220 , \30226 );
not \U$29851 ( \30228 , \30227 );
not \U$29852 ( \30229 , \11974 );
not \U$29853 ( \30230 , \29884 );
or \U$29854 ( \30231 , \30229 , \30230 );
not \U$29855 ( \30232 , RIc225b70_57);
not \U$29856 ( \30233 , \11854 );
or \U$29857 ( \30234 , \30232 , \30233 );
nand \U$29858 ( \30235 , \12990 , \10074 );
nand \U$29859 ( \30236 , \30234 , \30235 );
nand \U$29860 ( \30237 , \30236 , \11965 );
nand \U$29861 ( \30238 , \30231 , \30237 );
not \U$29862 ( \30239 , \30238 );
or \U$29863 ( \30240 , \30228 , \30239 );
or \U$29864 ( \30241 , \30238 , \30227 );
not \U$29865 ( \30242 , \11038 );
not \U$29866 ( \30243 , \29897 );
or \U$29867 ( \30244 , \30242 , \30243 );
not \U$29868 ( \30245 , RIc225c60_55);
not \U$29869 ( \30246 , \12977 );
or \U$29870 ( \30247 , \30245 , \30246 );
nand \U$29871 ( \30248 , \11844 , \11108 );
nand \U$29872 ( \30249 , \30247 , \30248 );
nand \U$29873 ( \30250 , \30249 , \11117 );
nand \U$29874 ( \30251 , \30244 , \30250 );
nand \U$29875 ( \30252 , \30241 , \30251 );
nand \U$29876 ( \30253 , \30240 , \30252 );
not \U$29877 ( \30254 , \30253 );
not \U$29878 ( \30255 , \30254 );
and \U$29879 ( \30256 , \11585 , \2634 );
not \U$29880 ( \30257 , \11585 );
and \U$29881 ( \30258 , \30257 , \14476 );
nor \U$29882 ( \30259 , \30256 , \30258 );
not \U$29883 ( \30260 , \30259 );
not \U$29884 ( \30261 , \8776 );
and \U$29885 ( \30262 , \30260 , \30261 );
and \U$29886 ( \30263 , \29997 , \11577 );
nor \U$29887 ( \30264 , \30262 , \30263 );
not \U$29888 ( \30265 , \30264 );
and \U$29889 ( \30266 , \30089 , \18037 );
not \U$29890 ( \30267 , RIc225a80_59);
not \U$29891 ( \30268 , \4802 );
or \U$29892 ( \30269 , \30267 , \30268 );
nand \U$29893 ( \30270 , \9360 , \17064 );
nand \U$29894 ( \30271 , \30269 , \30270 );
and \U$29895 ( \30272 , \30271 , \15164 );
nor \U$29896 ( \30273 , \30266 , \30272 );
not \U$29897 ( \30274 , \30273 );
or \U$29898 ( \30275 , \30265 , \30274 );
not \U$29899 ( \30276 , \9458 );
not \U$29900 ( \30277 , RIc225e40_51);
not \U$29901 ( \30278 , \3116 );
or \U$29902 ( \30279 , \30277 , \30278 );
not \U$29903 ( \30280 , \15755 );
nand \U$29904 ( \30281 , \30280 , \22140 );
nand \U$29905 ( \30282 , \30279 , \30281 );
not \U$29906 ( \30283 , \30282 );
or \U$29907 ( \30284 , \30276 , \30283 );
nand \U$29908 ( \30285 , \30098 , \9445 );
nand \U$29909 ( \30286 , \30284 , \30285 );
nand \U$29910 ( \30287 , \30275 , \30286 );
not \U$29911 ( \30288 , \30273 );
not \U$29912 ( \30289 , \30264 );
nand \U$29913 ( \30290 , \30288 , \30289 );
nand \U$29914 ( \30291 , \30287 , \30290 );
not \U$29915 ( \30292 , \30291 );
not \U$29916 ( \30293 , \30292 );
or \U$29917 ( \30294 , \30255 , \30293 );
not \U$29918 ( \30295 , \4381 );
not \U$29919 ( \30296 , RIc2265c0_35);
not \U$29920 ( \30297 , \8978 );
or \U$29921 ( \30298 , \30296 , \30297 );
nand \U$29922 ( \30299 , \8974 , \3620 );
nand \U$29923 ( \30300 , \30298 , \30299 );
not \U$29924 ( \30301 , \30300 );
or \U$29925 ( \30302 , \30295 , \30301 );
nand \U$29926 ( \30303 , \29956 , \5135 );
nand \U$29927 ( \30304 , \30302 , \30303 );
not \U$29928 ( \30305 , \9552 );
not \U$29929 ( \30306 , \29982 );
or \U$29930 ( \30307 , \30305 , \30306 );
not \U$29931 ( \30308 , RIc225f30_49);
not \U$29932 ( \30309 , \19926 );
or \U$29933 ( \30310 , \30308 , \30309 );
nand \U$29934 ( \30311 , \3641 , \28163 );
nand \U$29935 ( \30312 , \30310 , \30311 );
nand \U$29936 ( \30313 , \30312 , \9534 );
nand \U$29937 ( \30314 , \30307 , \30313 );
xor \U$29938 ( \30315 , \30304 , \30314 );
or \U$29939 ( \30316 , \29872 , \29866 );
not \U$29940 ( \30317 , RIc225990_61);
not \U$29941 ( \30318 , \9433 );
or \U$29942 ( \30319 , \30317 , \30318 );
nand \U$29943 ( \30320 , \9434 , \12806 );
nand \U$29944 ( \30321 , \30319 , \30320 );
nand \U$29945 ( \30322 , \30321 , \15719 );
nand \U$29946 ( \30323 , \30316 , \30322 );
and \U$29947 ( \30324 , \30315 , \30323 );
and \U$29948 ( \30325 , \30304 , \30314 );
or \U$29949 ( \30326 , \30324 , \30325 );
nand \U$29950 ( \30327 , \30294 , \30326 );
not \U$29951 ( \30328 , \30254 );
nand \U$29952 ( \30329 , \30328 , \30291 );
nand \U$29953 ( \30330 , \30327 , \30329 );
not \U$29954 ( \30331 , \30330 );
not \U$29955 ( \30332 , \2172 );
not \U$29956 ( \30333 , \29681 );
or \U$29957 ( \30334 , \30332 , \30333 );
not \U$29958 ( \30335 , RIc226a70_25);
not \U$29959 ( \30336 , \12862 );
or \U$29960 ( \30337 , \30335 , \30336 );
nand \U$29961 ( \30338 , \21175 , \6107 );
nand \U$29962 ( \30339 , \30337 , \30338 );
nand \U$29963 ( \30340 , \30339 , \2195 );
nand \U$29964 ( \30341 , \30334 , \30340 );
not \U$29965 ( \30342 , \30341 );
not \U$29966 ( \30343 , \30342 );
not \U$29967 ( \30344 , \2086 );
not \U$29968 ( \30345 , \29920 );
or \U$29969 ( \30346 , \30344 , \30345 );
and \U$29970 ( \30347 , RIc226890_29, \9250 );
not \U$29971 ( \30348 , RIc226890_29);
and \U$29972 ( \30349 , \30348 , \9254 );
or \U$29973 ( \30350 , \30347 , \30349 );
nand \U$29974 ( \30351 , \30350 , \2078 );
nand \U$29975 ( \30352 , \30346 , \30351 );
not \U$29976 ( \30353 , \30352 );
not \U$29977 ( \30354 , \30353 );
or \U$29978 ( \30355 , \30343 , \30354 );
not \U$29979 ( \30356 , \2710 );
not \U$29980 ( \30357 , \29932 );
or \U$29981 ( \30358 , \30356 , \30357 );
not \U$29982 ( \30359 , RIc2267a0_31);
not \U$29983 ( \30360 , \11478 );
or \U$29984 ( \30361 , \30359 , \30360 );
nand \U$29985 ( \30362 , \9077 , \3648 );
nand \U$29986 ( \30363 , \30361 , \30362 );
nand \U$29987 ( \30364 , \30363 , \2697 );
nand \U$29988 ( \30365 , \30358 , \30364 );
nand \U$29989 ( \30366 , \30355 , \30365 );
nand \U$29990 ( \30367 , \30352 , \30341 );
nand \U$29991 ( \30368 , \30366 , \30367 );
xor \U$29992 ( \30369 , \29924 , \29934 );
xor \U$29993 ( \30370 , \30369 , \29946 );
xor \U$29994 ( \30371 , \30368 , \30370 );
xor \U$29995 ( \30372 , \1911 , \12755 );
not \U$29996 ( \30373 , \30372 );
not \U$29997 ( \30374 , \10213 );
and \U$29998 ( \30375 , \30373 , \30374 );
and \U$29999 ( \30376 , \29787 , \1930 );
nor \U$30000 ( \30377 , \30375 , \30376 );
not \U$30001 ( \30378 , \30377 );
and \U$30002 ( \30379 , \30339 , \2172 );
not \U$30003 ( \30380 , \2194 );
and \U$30004 ( \30381 , \3982 , \10197 );
not \U$30005 ( \30382 , \3982 );
and \U$30006 ( \30383 , \30382 , \10198 );
nor \U$30007 ( \30384 , \30381 , \30383 );
nor \U$30008 ( \30385 , \30380 , \30384 );
nor \U$30009 ( \30386 , \30379 , \30385 );
not \U$30010 ( \30387 , \30386 );
or \U$30011 ( \30388 , \30378 , \30387 );
or \U$30012 ( \30389 , RIc226cc8_20, RIc226c50_21);
nand \U$30013 ( \30390 , \30389 , \18367 );
and \U$30014 ( \30391 , RIc226cc8_20, RIc226c50_21);
nor \U$30015 ( \30392 , \30391 , \1941 );
and \U$30016 ( \30393 , \30390 , \30392 );
not \U$30017 ( \30394 , \2533 );
not \U$30018 ( \30395 , \30049 );
or \U$30019 ( \30396 , \30394 , \30395 );
or \U$30020 ( \30397 , \18357 , \1941 );
or \U$30021 ( \30398 , \18181 , RIc226d40_19);
nand \U$30022 ( \30399 , \30397 , \30398 );
nand \U$30023 ( \30400 , \30399 , \2517 );
nand \U$30024 ( \30401 , \30396 , \30400 );
and \U$30025 ( \30402 , \30393 , \30401 );
nand \U$30026 ( \30403 , \30388 , \30402 );
not \U$30027 ( \30404 , \30386 );
not \U$30028 ( \30405 , \30377 );
nand \U$30029 ( \30406 , \30404 , \30405 );
nand \U$30030 ( \30407 , \30403 , \30406 );
not \U$30031 ( \30408 , \5509 );
not \U$30032 ( \30409 , RIc2264d0_37);
not \U$30033 ( \30410 , \8810 );
or \U$30034 ( \30411 , \30409 , \30410 );
nand \U$30035 ( \30412 , \8811 , \4371 );
nand \U$30036 ( \30413 , \30411 , \30412 );
not \U$30037 ( \30414 , \30413 );
or \U$30038 ( \30415 , \30408 , \30414 );
nand \U$30039 ( \30416 , \29967 , \5519 );
nand \U$30040 ( \30417 , \30415 , \30416 );
xor \U$30041 ( \30418 , \30407 , \30417 );
not \U$30042 ( \30419 , \6689 );
not \U$30043 ( \30420 , RIc2263e0_39);
not \U$30044 ( \30421 , \20674 );
or \U$30045 ( \30422 , \30420 , \30421 );
nand \U$30046 ( \30423 , \12727 , \8998 );
nand \U$30047 ( \30424 , \30422 , \30423 );
not \U$30048 ( \30425 , \30424 );
or \U$30049 ( \30426 , \30419 , \30425 );
nand \U$30050 ( \30427 , \29800 , \6307 );
nand \U$30051 ( \30428 , \30426 , \30427 );
and \U$30052 ( \30429 , \30418 , \30428 );
and \U$30053 ( \30430 , \30407 , \30417 );
or \U$30054 ( \30431 , \30429 , \30430 );
and \U$30055 ( \30432 , \30371 , \30431 );
and \U$30056 ( \30433 , \30368 , \30370 );
or \U$30057 ( \30434 , \30432 , \30433 );
not \U$30058 ( \30435 , \30434 );
nand \U$30059 ( \30436 , \30331 , \30435 );
xor \U$30060 ( \30437 , \29673 , \29683 );
xor \U$30061 ( \30438 , \30437 , \29695 );
and \U$30062 ( \30439 , RIc2266b0_33, \13129 );
not \U$30063 ( \30440 , RIc2266b0_33);
and \U$30064 ( \30441 , \30440 , \8924 );
nor \U$30065 ( \30442 , \30439 , \30441 );
not \U$30066 ( \30443 , \30442 );
not \U$30067 ( \30444 , \5185 );
and \U$30068 ( \30445 , \30443 , \30444 );
and \U$30069 ( \30446 , \29944 , \3631 );
nor \U$30070 ( \30447 , \30445 , \30446 );
not \U$30071 ( \30448 , \30447 );
and \U$30072 ( \30449 , \29744 , \9398 );
not \U$30073 ( \30450 , RIc226110_45);
not \U$30074 ( \30451 , \5664 );
or \U$30075 ( \30452 , \30450 , \30451 );
nand \U$30076 ( \30453 , \5663 , \10429 );
nand \U$30077 ( \30454 , \30452 , \30453 );
and \U$30078 ( \30455 , \30454 , \9934 );
nor \U$30079 ( \30456 , \30449 , \30455 );
not \U$30080 ( \30457 , \30456 );
or \U$30081 ( \30458 , \30448 , \30457 );
not \U$30082 ( \30459 , \10001 );
not \U$30083 ( \30460 , RIc226020_47);
not \U$30084 ( \30461 , \6076 );
or \U$30085 ( \30462 , \30460 , \30461 );
nand \U$30086 ( \30463 , \4406 , \11607 );
nand \U$30087 ( \30464 , \30462 , \30463 );
not \U$30088 ( \30465 , \30464 );
or \U$30089 ( \30466 , \30459 , \30465 );
nand \U$30090 ( \30467 , \29756 , \9619 );
nand \U$30091 ( \30468 , \30466 , \30467 );
nand \U$30092 ( \30469 , \30458 , \30468 );
not \U$30093 ( \30470 , \30447 );
not \U$30094 ( \30471 , \30456 );
nand \U$30095 ( \30472 , \30470 , \30471 );
nand \U$30096 ( \30473 , \30469 , \30472 );
xor \U$30097 ( \30474 , \30438 , \30473 );
xor \U$30098 ( \30475 , \29768 , \29778 );
xor \U$30099 ( \30476 , \30475 , \29789 );
not \U$30100 ( \30477 , \9110 );
not \U$30101 ( \30478 , RIc226200_43);
not \U$30102 ( \30479 , \9775 );
or \U$30103 ( \30480 , \30478 , \30479 );
nand \U$30104 ( \30481 , \13805 , \6492 );
nand \U$30105 ( \30482 , \30480 , \30481 );
not \U$30106 ( \30483 , \30482 );
or \U$30107 ( \30484 , \30477 , \30483 );
not \U$30108 ( \30485 , \9205 );
or \U$30109 ( \30486 , \29733 , \30485 );
nand \U$30110 ( \30487 , \30484 , \30486 );
xor \U$30111 ( \30488 , \30476 , \30487 );
not \U$30112 ( \30489 , \9816 );
not \U$30113 ( \30490 , \29809 );
or \U$30114 ( \30491 , \30489 , \30490 );
not \U$30115 ( \30492 , RIc2262f0_41);
not \U$30116 ( \30493 , \10142 );
or \U$30117 ( \30494 , \30492 , \30493 );
nand \U$30118 ( \30495 , \20646 , \6303 );
nand \U$30119 ( \30496 , \30494 , \30495 );
nand \U$30120 ( \30497 , \30496 , \9690 );
nand \U$30121 ( \30498 , \30491 , \30497 );
and \U$30122 ( \30499 , \30488 , \30498 );
and \U$30123 ( \30500 , \30476 , \30487 );
or \U$30124 ( \30501 , \30499 , \30500 );
and \U$30125 ( \30502 , \30474 , \30501 );
and \U$30126 ( \30503 , \30438 , \30473 );
or \U$30127 ( \30504 , \30502 , \30503 );
and \U$30128 ( \30505 , \30436 , \30504 );
nor \U$30129 ( \30506 , \30331 , \30435 );
nor \U$30130 ( \30507 , \30505 , \30506 );
not \U$30131 ( \30508 , \30507 );
not \U$30132 ( \30509 , \30508 );
or \U$30133 ( \30510 , \30217 , \30509 );
not \U$30134 ( \30511 , \30216 );
not \U$30135 ( \30512 , \30511 );
not \U$30136 ( \30513 , \30507 );
or \U$30137 ( \30514 , \30512 , \30513 );
xor \U$30138 ( \30515 , \29855 , \29857 );
xor \U$30139 ( \30516 , \30515 , \29906 );
nand \U$30140 ( \30517 , \30514 , \30516 );
nand \U$30141 ( \30518 , \30510 , \30517 );
nand \U$30142 ( \30519 , \30214 , \30518 );
nand \U$30143 ( \30520 , \30211 , \30519 );
not \U$30144 ( \30521 , \30520 );
or \U$30145 ( \30522 , \30201 , \30521 );
not \U$30146 ( \30523 , \30150 );
nand \U$30147 ( \30524 , \30523 , \30198 );
nand \U$30148 ( \30525 , \30522 , \30524 );
not \U$30149 ( \30526 , \30525 );
xor \U$30150 ( \30527 , \30148 , \30526 );
not \U$30151 ( \30528 , \29829 );
not \U$30152 ( \30529 , \29832 );
or \U$30153 ( \30530 , \30528 , \30529 );
or \U$30154 ( \30531 , \29832 , \29829 );
nand \U$30155 ( \30532 , \30530 , \30531 );
xor \U$30156 ( \30533 , \30127 , \30532 );
and \U$30157 ( \30534 , \30527 , \30533 );
and \U$30158 ( \30535 , \30148 , \30526 );
or \U$30159 ( \30536 , \30534 , \30535 );
nand \U$30160 ( \30537 , \30143 , \30536 );
not \U$30161 ( \30538 , \30537 );
not \U$30162 ( \30539 , \30124 );
not \U$30163 ( \30540 , \29845 );
and \U$30164 ( \30541 , \30539 , \30540 );
and \U$30165 ( \30542 , \29845 , \30124 );
nor \U$30166 ( \30543 , \30541 , \30542 );
not \U$30167 ( \30544 , \29839 );
and \U$30168 ( \30545 , \30543 , \30544 );
not \U$30169 ( \30546 , \30543 );
and \U$30170 ( \30547 , \30546 , \29839 );
nor \U$30171 ( \30548 , \30545 , \30547 );
xor \U$30172 ( \30549 , \30165 , \30189 );
xor \U$30173 ( \30550 , \30549 , \30192 );
not \U$30174 ( \30551 , \30550 );
xor \U$30175 ( \30552 , \30027 , \30024 );
buf \U$30176 ( \30553 , \30105 );
xor \U$30177 ( \30554 , \30552 , \30553 );
xor \U$30178 ( \30555 , \30040 , \30065 );
xor \U$30179 ( \30556 , \30555 , \30077 );
xor \U$30180 ( \30557 , \30041 , \30051 );
xor \U$30181 ( \30558 , \30557 , \30062 );
and \U$30182 ( \30559 , RIc226890_29, \10975 );
not \U$30183 ( \30560 , RIc226890_29);
and \U$30184 ( \30561 , \30560 , \9275 );
or \U$30185 ( \30562 , \30559 , \30561 );
not \U$30186 ( \30563 , \30562 );
or \U$30187 ( \30564 , \30563 , \3930 );
not \U$30188 ( \30565 , \30350 );
or \U$30189 ( \30566 , \30565 , \20641 );
nand \U$30190 ( \30567 , \30564 , \30566 );
xor \U$30191 ( \30568 , \30558 , \30567 );
not \U$30192 ( \30569 , \2154 );
not \U$30193 ( \30570 , \30073 );
or \U$30194 ( \30571 , \30569 , \30570 );
not \U$30195 ( \30572 , RIc226980_27);
buf \U$30196 ( \30573 , \9320 );
not \U$30197 ( \30574 , \30573 );
not \U$30198 ( \30575 , \30574 );
or \U$30199 ( \30576 , \30572 , \30575 );
nand \U$30200 ( \30577 , \30573 , \2150 );
nand \U$30201 ( \30578 , \30576 , \30577 );
nand \U$30202 ( \30579 , \30578 , \2138 );
nand \U$30203 ( \30580 , \30571 , \30579 );
and \U$30204 ( \30581 , \30568 , \30580 );
and \U$30205 ( \30582 , \30558 , \30567 );
or \U$30206 ( \30583 , \30581 , \30582 );
xor \U$30207 ( \30584 , \30556 , \30583 );
not \U$30208 ( \30585 , \30341 );
not \U$30209 ( \30586 , \30353 );
or \U$30210 ( \30587 , \30585 , \30586 );
or \U$30211 ( \30588 , \30353 , \30341 );
nand \U$30212 ( \30589 , \30587 , \30588 );
xor \U$30213 ( \30590 , \30365 , \30589 );
and \U$30214 ( \30591 , \30584 , \30590 );
and \U$30215 ( \30592 , \30556 , \30583 );
or \U$30216 ( \30593 , \30591 , \30592 );
not \U$30217 ( \30594 , \2710 );
not \U$30218 ( \30595 , \30363 );
or \U$30219 ( \30596 , \30594 , \30595 );
not \U$30220 ( \30597 , RIc2267a0_31);
not \U$30221 ( \30598 , \13223 );
or \U$30222 ( \30599 , \30597 , \30598 );
nand \U$30223 ( \30600 , \10110 , \2705 );
nand \U$30224 ( \30601 , \30599 , \30600 );
nand \U$30225 ( \30602 , \30601 , \2697 );
nand \U$30226 ( \30603 , \30596 , \30602 );
not \U$30227 ( \30604 , RIc2266b0_33);
not \U$30228 ( \30605 , \13465 );
or \U$30229 ( \30606 , \30604 , \30605 );
nand \U$30230 ( \30607 , \9225 , \9943 );
nand \U$30231 ( \30608 , \30606 , \30607 );
not \U$30232 ( \30609 , \30608 );
not \U$30233 ( \30610 , \3629 );
or \U$30234 ( \30611 , \30609 , \30610 );
not \U$30235 ( \30612 , \30442 );
nand \U$30236 ( \30613 , \30612 , \3631 );
nand \U$30237 ( \30614 , \30611 , \30613 );
xor \U$30238 ( \30615 , \30603 , \30614 );
not \U$30239 ( \30616 , \12304 );
not \U$30240 ( \30617 , \30464 );
or \U$30241 ( \30618 , \30616 , \30617 );
not \U$30242 ( \30619 , \13515 );
and \U$30243 ( \30620 , RIc226020_47, \30619 );
not \U$30244 ( \30621 , RIc226020_47);
and \U$30245 ( \30622 , \30621 , \5217 );
nor \U$30246 ( \30623 , \30620 , \30622 );
or \U$30247 ( \30624 , \30623 , \9640 );
nand \U$30248 ( \30625 , \30618 , \30624 );
and \U$30249 ( \30626 , \30615 , \30625 );
and \U$30250 ( \30627 , \30603 , \30614 );
or \U$30251 ( \30628 , \30626 , \30627 );
not \U$30252 ( \30629 , \30628 );
not \U$30253 ( \30630 , \9110 );
not \U$30254 ( \30631 , RIc226200_43);
not \U$30255 ( \30632 , \23758 );
or \U$30256 ( \30633 , \30631 , \30632 );
not \U$30257 ( \30634 , \18410 );
nand \U$30258 ( \30635 , \30634 , \13805 );
nand \U$30259 ( \30636 , \30633 , \30635 );
not \U$30260 ( \30637 , \30636 );
or \U$30261 ( \30638 , \30630 , \30637 );
nand \U$30262 ( \30639 , \30482 , \9129 );
nand \U$30263 ( \30640 , \30638 , \30639 );
not \U$30264 ( \30641 , \9398 );
not \U$30265 ( \30642 , \30454 );
or \U$30266 ( \30643 , \30641 , \30642 );
not \U$30267 ( \30644 , RIc226110_45);
not \U$30268 ( \30645 , \9765 );
or \U$30269 ( \30646 , \30644 , \30645 );
nand \U$30270 ( \30647 , \6071 , \9379 );
nand \U$30271 ( \30648 , \30646 , \30647 );
nand \U$30272 ( \30649 , \30648 , \9934 );
nand \U$30273 ( \30650 , \30643 , \30649 );
nor \U$30274 ( \30651 , \30640 , \30650 );
not \U$30275 ( \30652 , \9552 );
not \U$30276 ( \30653 , \30312 );
or \U$30277 ( \30654 , \30652 , \30653 );
not \U$30278 ( \30655 , RIc225f30_49);
not \U$30279 ( \30656 , \4414 );
or \U$30280 ( \30657 , \30655 , \30656 );
not \U$30281 ( \30658 , \4122 );
nand \U$30282 ( \30659 , \30658 , \9549 );
nand \U$30283 ( \30660 , \30657 , \30659 );
nand \U$30284 ( \30661 , \30660 , \10445 );
nand \U$30285 ( \30662 , \30654 , \30661 );
not \U$30286 ( \30663 , \30662 );
or \U$30287 ( \30664 , \30651 , \30663 );
nand \U$30288 ( \30665 , \30640 , \30650 );
nand \U$30289 ( \30666 , \30664 , \30665 );
not \U$30290 ( \30667 , \30666 );
or \U$30291 ( \30668 , \30629 , \30667 );
not \U$30292 ( \30669 , \30628 );
not \U$30293 ( \30670 , \30669 );
not \U$30294 ( \30671 , \30666 );
not \U$30295 ( \30672 , \30671 );
or \U$30296 ( \30673 , \30670 , \30672 );
xor \U$30297 ( \30674 , \30393 , \30401 );
not \U$30298 ( \30675 , \2367 );
not \U$30299 ( \30676 , \30058 );
or \U$30300 ( \30677 , \30675 , \30676 );
not \U$30301 ( \30678 , RIc226c50_21);
not \U$30302 ( \30679 , \13487 );
not \U$30303 ( \30680 , \30679 );
or \U$30304 ( \30681 , \30678 , \30680 );
nand \U$30305 ( \30682 , \13488 , \3204 );
nand \U$30306 ( \30683 , \30681 , \30682 );
nand \U$30307 ( \30684 , \30683 , \2391 );
nand \U$30308 ( \30685 , \30677 , \30684 );
xor \U$30309 ( \30686 , \30674 , \30685 );
not \U$30310 ( \30687 , \2195 );
not \U$30311 ( \30688 , RIc226a70_25);
not \U$30312 ( \30689 , \17625 );
or \U$30313 ( \30690 , \30688 , \30689 );
nand \U$30314 ( \30691 , \20406 , \3982 );
nand \U$30315 ( \30692 , \30690 , \30691 );
not \U$30316 ( \30693 , \30692 );
or \U$30317 ( \30694 , \30687 , \30693 );
not \U$30318 ( \30695 , \30384 );
nand \U$30319 ( \30696 , \30695 , \2172 );
nand \U$30320 ( \30697 , \30694 , \30696 );
and \U$30321 ( \30698 , \30686 , \30697 );
and \U$30322 ( \30699 , \30674 , \30685 );
or \U$30323 ( \30700 , \30698 , \30699 );
not \U$30324 ( \30701 , \6688 );
not \U$30325 ( \30702 , RIc2263e0_39);
not \U$30326 ( \30703 , \9900 );
or \U$30327 ( \30704 , \30702 , \30703 );
nand \U$30328 ( \30705 , \10289 , \8990 );
nand \U$30329 ( \30706 , \30704 , \30705 );
not \U$30330 ( \30707 , \30706 );
or \U$30331 ( \30708 , \30701 , \30707 );
nand \U$30332 ( \30709 , \30424 , \6307 );
nand \U$30333 ( \30710 , \30708 , \30709 );
xor \U$30334 ( \30711 , \30700 , \30710 );
not \U$30335 ( \30712 , \9690 );
and \U$30336 ( \30713 , \8886 , \12937 );
not \U$30337 ( \30714 , \8886 );
and \U$30338 ( \30715 , \30714 , RIc2262f0_41);
or \U$30339 ( \30716 , \30713 , \30715 );
not \U$30340 ( \30717 , \30716 );
or \U$30341 ( \30718 , \30712 , \30717 );
nand \U$30342 ( \30719 , \30496 , \9705 );
nand \U$30343 ( \30720 , \30718 , \30719 );
and \U$30344 ( \30721 , \30711 , \30720 );
and \U$30345 ( \30722 , \30700 , \30710 );
or \U$30346 ( \30723 , \30721 , \30722 );
nand \U$30347 ( \30724 , \30673 , \30723 );
nand \U$30348 ( \30725 , \30668 , \30724 );
xor \U$30349 ( \30726 , \30593 , \30725 );
xor \U$30350 ( \30727 , \30407 , \30417 );
xor \U$30351 ( \30728 , \30727 , \30428 );
not \U$30352 ( \30729 , \30468 );
not \U$30353 ( \30730 , \30447 );
and \U$30354 ( \30731 , \30729 , \30730 );
and \U$30355 ( \30732 , \30468 , \30447 );
nor \U$30356 ( \30733 , \30731 , \30732 );
and \U$30357 ( \30734 , \30733 , \30471 );
not \U$30358 ( \30735 , \30733 );
and \U$30359 ( \30736 , \30735 , \30456 );
or \U$30360 ( \30737 , \30734 , \30736 );
or \U$30361 ( \30738 , \30728 , \30737 );
xor \U$30362 ( \30739 , \30476 , \30487 );
xor \U$30363 ( \30740 , \30739 , \30498 );
nand \U$30364 ( \30741 , \30738 , \30740 );
nand \U$30365 ( \30742 , \30737 , \30728 );
nand \U$30366 ( \30743 , \30741 , \30742 );
and \U$30367 ( \30744 , \30726 , \30743 );
and \U$30368 ( \30745 , \30593 , \30725 );
or \U$30369 ( \30746 , \30744 , \30745 );
xor \U$30370 ( \30747 , \30554 , \30746 );
and \U$30371 ( \30748 , \30504 , \30434 );
not \U$30372 ( \30749 , \30504 );
and \U$30373 ( \30750 , \30749 , \30435 );
nor \U$30374 ( \30751 , \30748 , \30750 );
and \U$30375 ( \30752 , \30751 , \30330 );
not \U$30376 ( \30753 , \30751 );
and \U$30377 ( \30754 , \30753 , \30331 );
nor \U$30378 ( \30755 , \30752 , \30754 );
and \U$30379 ( \30756 , \30747 , \30755 );
and \U$30380 ( \30757 , \30554 , \30746 );
or \U$30381 ( \30758 , \30756 , \30757 );
not \U$30382 ( \30759 , \30758 );
or \U$30383 ( \30760 , \30551 , \30759 );
or \U$30384 ( \30761 , \30550 , \30758 );
and \U$30385 ( \30762 , \29760 , \29748 );
not \U$30386 ( \30763 , \29760 );
and \U$30387 ( \30764 , \30763 , \29749 );
nor \U$30388 ( \30765 , \30762 , \30764 );
not \U$30389 ( \30766 , \29738 );
and \U$30390 ( \30767 , \30765 , \30766 );
not \U$30391 ( \30768 , \30765 );
and \U$30392 ( \30769 , \30768 , \29738 );
nor \U$30393 ( \30770 , \30767 , \30769 );
not \U$30394 ( \30771 , \30770 );
not \U$30395 ( \30772 , \30771 );
not \U$30396 ( \30773 , \29984 );
not \U$30397 ( \30774 , \29972 );
not \U$30398 ( \30775 , \29960 );
and \U$30399 ( \30776 , \30774 , \30775 );
and \U$30400 ( \30777 , \29960 , \29972 );
nor \U$30401 ( \30778 , \30776 , \30777 );
not \U$30402 ( \30779 , \30778 );
or \U$30403 ( \30780 , \30773 , \30779 );
or \U$30404 ( \30781 , \29984 , \30778 );
nand \U$30405 ( \30782 , \30780 , \30781 );
not \U$30406 ( \30783 , \30782 );
or \U$30407 ( \30784 , \30772 , \30783 );
not \U$30408 ( \30785 , \30782 );
nand \U$30409 ( \30786 , \30785 , \30770 );
nand \U$30410 ( \30787 , \30784 , \30786 );
xor \U$30411 ( \30788 , \29792 , \29802 );
xor \U$30412 ( \30789 , \30788 , \29813 );
not \U$30413 ( \30790 , \30789 );
and \U$30414 ( \30791 , \30787 , \30790 );
not \U$30415 ( \30792 , \30787 );
and \U$30416 ( \30793 , \30792 , \30789 );
nor \U$30417 ( \30794 , \30791 , \30793 );
not \U$30418 ( \30795 , \30794 );
not \U$30419 ( \30796 , \30795 );
not \U$30420 ( \30797 , \30253 );
not \U$30421 ( \30798 , \30326 );
not \U$30422 ( \30799 , \30798 );
or \U$30423 ( \30800 , \30797 , \30799 );
nand \U$30424 ( \30801 , \30254 , \30326 );
nand \U$30425 ( \30802 , \30800 , \30801 );
and \U$30426 ( \30803 , \30802 , \30292 );
not \U$30427 ( \30804 , \30802 );
and \U$30428 ( \30805 , \30804 , \30291 );
nor \U$30429 ( \30806 , \30803 , \30805 );
not \U$30430 ( \30807 , \30806 );
not \U$30431 ( \30808 , \30807 );
or \U$30432 ( \30809 , \30796 , \30808 );
xor \U$30433 ( \30810 , \30304 , \30314 );
xor \U$30434 ( \30811 , \30810 , \30323 );
not \U$30435 ( \30812 , \30372 );
nand \U$30436 ( \30813 , \30812 , \1930 );
not \U$30437 ( \30814 , RIc226b60_23);
not \U$30438 ( \30815 , \19721 );
not \U$30439 ( \30816 , \30815 );
or \U$30440 ( \30817 , \30814 , \30816 );
nand \U$30441 ( \30818 , \19721 , \1927 );
nand \U$30442 ( \30819 , \30817 , \30818 );
nand \U$30443 ( \30820 , \30819 , \1914 );
nand \U$30444 ( \30821 , \30813 , \30820 );
and \U$30445 ( \30822 , \16248 , \2533 );
not \U$30446 ( \30823 , \2367 );
not \U$30447 ( \30824 , \30683 );
or \U$30448 ( \30825 , \30823 , \30824 );
not \U$30449 ( \30826 , RIc226c50_21);
not \U$30450 ( \30827 , \16256 );
not \U$30451 ( \30828 , \30827 );
or \U$30452 ( \30829 , \30826 , \30828 );
nand \U$30453 ( \30830 , \16256 , \2383 );
nand \U$30454 ( \30831 , \30829 , \30830 );
nand \U$30455 ( \30832 , \30831 , \2391 );
nand \U$30456 ( \30833 , \30825 , \30832 );
xor \U$30457 ( \30834 , \30822 , \30833 );
not \U$30458 ( \30835 , \1914 );
not \U$30459 ( \30836 , RIc226b60_23);
not \U$30460 ( \30837 , \12846 );
or \U$30461 ( \30838 , \30836 , \30837 );
nand \U$30462 ( \30839 , \18161 , \5637 );
nand \U$30463 ( \30840 , \30838 , \30839 );
not \U$30464 ( \30841 , \30840 );
or \U$30465 ( \30842 , \30835 , \30841 );
nand \U$30466 ( \30843 , \30819 , \1930 );
nand \U$30467 ( \30844 , \30842 , \30843 );
and \U$30468 ( \30845 , \30834 , \30844 );
and \U$30469 ( \30846 , \30822 , \30833 );
or \U$30470 ( \30847 , \30845 , \30846 );
xor \U$30471 ( \30848 , \30821 , \30847 );
not \U$30472 ( \30849 , \2784 );
and \U$30473 ( \30850 , RIc226890_29, \10263 );
not \U$30474 ( \30851 , RIc226890_29);
not \U$30475 ( \30852 , \30069 );
and \U$30476 ( \30853 , \30851 , \30852 );
or \U$30477 ( \30854 , \30850 , \30853 );
not \U$30478 ( \30855 , \30854 );
or \U$30479 ( \30856 , \30849 , \30855 );
nand \U$30480 ( \30857 , \30562 , \2086 );
nand \U$30481 ( \30858 , \30856 , \30857 );
and \U$30482 ( \30859 , \30848 , \30858 );
and \U$30483 ( \30860 , \30821 , \30847 );
or \U$30484 ( \30861 , \30859 , \30860 );
not \U$30485 ( \30862 , \2154 );
not \U$30486 ( \30863 , \30578 );
or \U$30487 ( \30864 , \30862 , \30863 );
not \U$30488 ( \30865 , RIc226980_27);
not \U$30489 ( \30866 , \16945 );
or \U$30490 ( \30867 , \30865 , \30866 );
nand \U$30491 ( \30868 , \10086 , \2150 );
nand \U$30492 ( \30869 , \30867 , \30868 );
nand \U$30493 ( \30870 , \30869 , \2138 );
nand \U$30494 ( \30871 , \30864 , \30870 );
not \U$30495 ( \30872 , \30871 );
not \U$30496 ( \30873 , \2697 );
not \U$30497 ( \30874 , RIc2267a0_31);
buf \U$30498 ( \30875 , \9255 );
not \U$30499 ( \30876 , \30875 );
or \U$30500 ( \30877 , \30874 , \30876 );
not \U$30501 ( \30878 , \11488 );
nand \U$30502 ( \30879 , \30878 , \2705 );
nand \U$30503 ( \30880 , \30877 , \30879 );
not \U$30504 ( \30881 , \30880 );
or \U$30505 ( \30882 , \30873 , \30881 );
nand \U$30506 ( \30883 , \30601 , \2710 );
nand \U$30507 ( \30884 , \30882 , \30883 );
not \U$30508 ( \30885 , \30884 );
or \U$30509 ( \30886 , \30872 , \30885 );
or \U$30510 ( \30887 , \30884 , \30871 );
not \U$30511 ( \30888 , \3631 );
not \U$30512 ( \30889 , \30608 );
or \U$30513 ( \30890 , \30888 , \30889 );
not \U$30514 ( \30891 , RIc2266b0_33);
not \U$30515 ( \30892 , \10652 );
or \U$30516 ( \30893 , \30891 , \30892 );
nand \U$30517 ( \30894 , \10653 , \5179 );
nand \U$30518 ( \30895 , \30893 , \30894 );
nand \U$30519 ( \30896 , \30895 , \3629 );
nand \U$30520 ( \30897 , \30890 , \30896 );
nand \U$30521 ( \30898 , \30887 , \30897 );
nand \U$30522 ( \30899 , \30886 , \30898 );
xor \U$30523 ( \30900 , \30861 , \30899 );
not \U$30524 ( \30901 , \9459 );
not \U$30525 ( \30902 , RIc225e40_51);
not \U$30526 ( \30903 , \6439 );
or \U$30527 ( \30904 , \30902 , \30903 );
nand \U$30528 ( \30905 , \3728 , \22140 );
nand \U$30529 ( \30906 , \30904 , \30905 );
not \U$30530 ( \30907 , \30906 );
or \U$30531 ( \30908 , \30901 , \30907 );
nand \U$30532 ( \30909 , \30282 , \9444 );
nand \U$30533 ( \30910 , \30908 , \30909 );
and \U$30534 ( \30911 , \30900 , \30910 );
and \U$30535 ( \30912 , \30861 , \30899 );
or \U$30536 ( \30913 , \30911 , \30912 );
xor \U$30537 ( \30914 , \30811 , \30913 );
not \U$30538 ( \30915 , \30289 );
and \U$30539 ( \30916 , \30273 , \30915 );
not \U$30540 ( \30917 , \30273 );
not \U$30541 ( \30918 , \30264 );
and \U$30542 ( \30919 , \30917 , \30918 );
or \U$30543 ( \30920 , \30916 , \30919 );
and \U$30544 ( \30921 , \30286 , \30920 );
not \U$30545 ( \30922 , \30286 );
not \U$30546 ( \30923 , \30289 );
and \U$30547 ( \30924 , \30288 , \30923 );
not \U$30548 ( \30925 , \30288 );
not \U$30549 ( \30926 , \30264 );
and \U$30550 ( \30927 , \30925 , \30926 );
or \U$30551 ( \30928 , \30924 , \30927 );
and \U$30552 ( \30929 , \30922 , \30928 );
or \U$30553 ( \30930 , \30921 , \30929 );
and \U$30554 ( \30931 , \30914 , \30930 );
and \U$30555 ( \30932 , \30811 , \30913 );
or \U$30556 ( \30933 , \30931 , \30932 );
nand \U$30557 ( \30934 , \30806 , \30794 );
nand \U$30558 ( \30935 , \30933 , \30934 );
nand \U$30559 ( \30936 , \30809 , \30935 );
not \U$30560 ( \30937 , \30936 );
xor \U$30561 ( \30938 , \29728 , \29816 );
xnor \U$30562 ( \30939 , \30938 , \29763 );
not \U$30563 ( \30940 , \30770 );
not \U$30564 ( \30941 , \30782 );
or \U$30565 ( \30942 , \30940 , \30941 );
not \U$30566 ( \30943 , \30785 );
not \U$30567 ( \30944 , \30771 );
or \U$30568 ( \30945 , \30943 , \30944 );
nand \U$30569 ( \30946 , \30945 , \30789 );
nand \U$30570 ( \30947 , \30942 , \30946 );
and \U$30571 ( \30948 , \30939 , \30947 );
not \U$30572 ( \30949 , \30939 );
not \U$30573 ( \30950 , \30947 );
and \U$30574 ( \30951 , \30949 , \30950 );
or \U$30575 ( \30952 , \30948 , \30951 );
not \U$30576 ( \30953 , \29949 );
and \U$30577 ( \30954 , \30019 , \30953 );
not \U$30578 ( \30955 , \30019 );
and \U$30579 ( \30956 , \30955 , \29949 );
nor \U$30580 ( \30957 , \30954 , \30956 );
and \U$30581 ( \30958 , \30957 , \29988 );
not \U$30582 ( \30959 , \30957 );
not \U$30583 ( \30960 , \29988 );
and \U$30584 ( \30961 , \30959 , \30960 );
nor \U$30585 ( \30962 , \30958 , \30961 );
not \U$30586 ( \30963 , \30962 );
and \U$30587 ( \30964 , \30952 , \30963 );
not \U$30588 ( \30965 , \30952 );
not \U$30589 ( \30966 , \30963 );
and \U$30590 ( \30967 , \30965 , \30966 );
nor \U$30591 ( \30968 , \30964 , \30967 );
not \U$30592 ( \30969 , \30968 );
or \U$30593 ( \30970 , \30937 , \30969 );
or \U$30594 ( \30971 , \30936 , \30968 );
xor \U$30595 ( \30972 , \30368 , \30370 );
xor \U$30596 ( \30973 , \30972 , \30431 );
xor \U$30597 ( \30974 , \30438 , \30473 );
xor \U$30598 ( \30975 , \30974 , \30501 );
xor \U$30599 ( \30976 , \30973 , \30975 );
not \U$30600 ( \30977 , \5741 );
not \U$30601 ( \30978 , RIc2265c0_35);
not \U$30602 ( \30979 , \9787 );
or \U$30603 ( \30980 , \30978 , \30979 );
nand \U$30604 ( \30981 , \12406 , \4376 );
nand \U$30605 ( \30982 , \30980 , \30981 );
not \U$30606 ( \30983 , \30982 );
or \U$30607 ( \30984 , \30977 , \30983 );
nand \U$30608 ( \30985 , \30300 , \4383 );
nand \U$30609 ( \30986 , \30984 , \30985 );
not \U$30610 ( \30987 , \5509 );
not \U$30611 ( \30988 , RIc2264d0_37);
not \U$30612 ( \30989 , \13370 );
or \U$30613 ( \30990 , \30988 , \30989 );
nand \U$30614 ( \30991 , \20368 , \4371 );
nand \U$30615 ( \30992 , \30990 , \30991 );
not \U$30616 ( \30993 , \30992 );
or \U$30617 ( \30994 , \30987 , \30993 );
nand \U$30618 ( \30995 , \30413 , \5519 );
nand \U$30619 ( \30996 , \30994 , \30995 );
xor \U$30620 ( \30997 , \30986 , \30996 );
not \U$30621 ( \30998 , \11965 );
not \U$30622 ( \30999 , RIc225b70_57);
not \U$30623 ( \31000 , \2670 );
or \U$30624 ( \31001 , \30999 , \31000 );
nand \U$30625 ( \31002 , \17831 , \11033 );
nand \U$30626 ( \31003 , \31001 , \31002 );
not \U$30627 ( \31004 , \31003 );
or \U$30628 ( \31005 , \30998 , \31004 );
nand \U$30629 ( \31006 , \30236 , \15267 );
nand \U$30630 ( \31007 , \31005 , \31006 );
and \U$30631 ( \31008 , \30997 , \31007 );
and \U$30632 ( \31009 , \30986 , \30996 );
or \U$30633 ( \31010 , \31008 , \31009 );
not \U$30634 ( \31011 , RIc225828_64);
not \U$30635 ( \31012 , \30225 );
or \U$30636 ( \31013 , \31011 , \31012 );
not \U$30637 ( \31014 , RIc2258a0_63);
not \U$30638 ( \31015 , \3839 );
or \U$30639 ( \31016 , \31014 , \31015 );
nand \U$30640 ( \31017 , \3834 , \16880 );
nand \U$30641 ( \31018 , \31016 , \31017 );
nand \U$30642 ( \31019 , \31018 , \16891 );
nand \U$30643 ( \31020 , \31013 , \31019 );
not \U$30644 ( \31021 , \31020 );
not \U$30645 ( \31022 , \15729 );
not \U$30646 ( \31023 , \30321 );
or \U$30647 ( \31024 , \31022 , \31023 );
not \U$30648 ( \31025 , RIc225990_61);
not \U$30649 ( \31026 , \2586 );
or \U$30650 ( \31027 , \31025 , \31026 );
nand \U$30651 ( \31028 , \3183 , \12806 );
nand \U$30652 ( \31029 , \31027 , \31028 );
nand \U$30653 ( \31030 , \31029 , \15719 );
nand \U$30654 ( \31031 , \31024 , \31030 );
not \U$30655 ( \31032 , \31031 );
or \U$30656 ( \31033 , \31021 , \31032 );
or \U$30657 ( \31034 , \31031 , \31020 );
not \U$30658 ( \31035 , \11038 );
not \U$30659 ( \31036 , \30249 );
or \U$30660 ( \31037 , \31035 , \31036 );
not \U$30661 ( \31038 , RIc225c60_55);
not \U$30662 ( \31039 , \5526 );
or \U$30663 ( \31040 , \31038 , \31039 );
nand \U$30664 ( \31041 , \2730 , \11108 );
nand \U$30665 ( \31042 , \31040 , \31041 );
nand \U$30666 ( \31043 , \31042 , \11118 );
nand \U$30667 ( \31044 , \31037 , \31043 );
nand \U$30668 ( \31045 , \31034 , \31044 );
nand \U$30669 ( \31046 , \31033 , \31045 );
xor \U$30670 ( \31047 , \31010 , \31046 );
not \U$30671 ( \31048 , \12670 );
not \U$30672 ( \31049 , \30271 );
or \U$30673 ( \31050 , \31048 , \31049 );
not \U$30674 ( \31051 , RIc225a80_59);
not \U$30675 ( \31052 , \2476 );
or \U$30676 ( \31053 , \31051 , \31052 );
not \U$30677 ( \31054 , \28706 );
nand \U$30678 ( \31055 , \31054 , \17064 );
nand \U$30679 ( \31056 , \31053 , \31055 );
nand \U$30680 ( \31057 , \31056 , \15164 );
nand \U$30681 ( \31058 , \31050 , \31057 );
not \U$30682 ( \31059 , \31058 );
not \U$30683 ( \31060 , \8777 );
and \U$30684 ( \31061 , RIc225d50_53, \9651 );
not \U$30685 ( \31062 , RIc225d50_53);
and \U$30686 ( \31063 , \31062 , \10533 );
or \U$30687 ( \31064 , \31061 , \31063 );
not \U$30688 ( \31065 , \31064 );
or \U$30689 ( \31066 , \31060 , \31065 );
not \U$30690 ( \31067 , \30259 );
nand \U$30691 ( \31068 , \31067 , \12945 );
nand \U$30692 ( \31069 , \31066 , \31068 );
not \U$30693 ( \31070 , \31069 );
or \U$30694 ( \31071 , \31059 , \31070 );
or \U$30695 ( \31072 , \31069 , \31058 );
xor \U$30696 ( \31073 , \30402 , \30405 );
xnor \U$30697 ( \31074 , \31073 , \30404 );
not \U$30698 ( \31075 , \31074 );
nand \U$30699 ( \31076 , \31072 , \31075 );
nand \U$30700 ( \31077 , \31071 , \31076 );
and \U$30701 ( \31078 , \31047 , \31077 );
and \U$30702 ( \31079 , \31010 , \31046 );
or \U$30703 ( \31080 , \31078 , \31079 );
and \U$30704 ( \31081 , \30976 , \31080 );
and \U$30705 ( \31082 , \30973 , \30975 );
or \U$30706 ( \31083 , \31081 , \31082 );
nand \U$30707 ( \31084 , \30971 , \31083 );
nand \U$30708 ( \31085 , \30970 , \31084 );
nand \U$30709 ( \31086 , \30761 , \31085 );
nand \U$30710 ( \31087 , \30760 , \31086 );
not \U$30711 ( \31088 , \31087 );
xor \U$30712 ( \31089 , \30152 , \30162 );
xor \U$30713 ( \31090 , \31089 , \30195 );
not \U$30714 ( \31091 , \31090 );
not \U$30715 ( \31092 , \30963 );
not \U$30716 ( \31093 , \30947 );
or \U$30717 ( \31094 , \31092 , \31093 );
not \U$30718 ( \31095 , \30950 );
not \U$30719 ( \31096 , \30962 );
or \U$30720 ( \31097 , \31095 , \31096 );
not \U$30721 ( \31098 , \30939 );
nand \U$30722 ( \31099 , \31097 , \31098 );
nand \U$30723 ( \31100 , \31094 , \31099 );
and \U$30724 ( \31101 , \30107 , \30021 );
not \U$30725 ( \31102 , \30107 );
not \U$30726 ( \31103 , \30021 );
and \U$30727 ( \31104 , \31102 , \31103 );
nor \U$30728 ( \31105 , \31101 , \31104 );
xor \U$30729 ( \31106 , \31105 , \30120 );
xor \U$30730 ( \31107 , \31100 , \31106 );
xor \U$30731 ( \31108 , \30187 , \30167 );
xor \U$30732 ( \31109 , \31108 , \30178 );
not \U$30733 ( \31110 , \31109 );
not \U$30734 ( \31111 , \31110 );
xor \U$30735 ( \31112 , \29860 , \29862 );
xor \U$30736 ( \31113 , \31112 , \29903 );
not \U$30737 ( \31114 , \31113 );
or \U$30738 ( \31115 , \31111 , \31114 );
not \U$30739 ( \31116 , \31113 );
not \U$30740 ( \31117 , \31116 );
not \U$30741 ( \31118 , \31109 );
or \U$30742 ( \31119 , \31117 , \31118 );
not \U$30743 ( \31120 , \30012 );
not \U$30744 ( \31121 , \30001 );
not \U$30745 ( \31122 , \30017 );
not \U$30746 ( \31123 , \31122 );
and \U$30747 ( \31124 , \31121 , \31123 );
and \U$30748 ( \31125 , \30001 , \31122 );
nor \U$30749 ( \31126 , \31124 , \31125 );
not \U$30750 ( \31127 , \31126 );
or \U$30751 ( \31128 , \31120 , \31127 );
or \U$30752 ( \31129 , \31126 , \30012 );
nand \U$30753 ( \31130 , \31128 , \31129 );
xnor \U$30754 ( \31131 , \29899 , \29887 );
xnor \U$30755 ( \31132 , \29875 , \31131 );
xor \U$30756 ( \31133 , \31130 , \31132 );
xor \U$30757 ( \31134 , \30080 , \30091 );
xor \U$30758 ( \31135 , \31134 , \30102 );
and \U$30759 ( \31136 , \31133 , \31135 );
and \U$30760 ( \31137 , \31130 , \31132 );
or \U$30761 ( \31138 , \31136 , \31137 );
nand \U$30762 ( \31139 , \31119 , \31138 );
nand \U$30763 ( \31140 , \31115 , \31139 );
and \U$30764 ( \31141 , \31107 , \31140 );
and \U$30765 ( \31142 , \31100 , \31106 );
or \U$30766 ( \31143 , \31141 , \31142 );
not \U$30767 ( \31144 , \31143 );
nand \U$30768 ( \31145 , \31091 , \31144 );
not \U$30769 ( \31146 , \31145 );
or \U$30770 ( \31147 , \31088 , \31146 );
not \U$30771 ( \31148 , \31144 );
nand \U$30772 ( \31149 , \31148 , \31090 );
nand \U$30773 ( \31150 , \31147 , \31149 );
not \U$30774 ( \31151 , \31150 );
xor \U$30775 ( \31152 , \30548 , \31151 );
not \U$30776 ( \31153 , \30199 );
not \U$30777 ( \31154 , \30523 );
or \U$30778 ( \31155 , \31153 , \31154 );
nand \U$30779 ( \31156 , \30150 , \30198 );
nand \U$30780 ( \31157 , \31155 , \31156 );
not \U$30781 ( \31158 , \30520 );
and \U$30782 ( \31159 , \31157 , \31158 );
not \U$30783 ( \31160 , \31157 );
and \U$30784 ( \31161 , \31160 , \30520 );
nor \U$30785 ( \31162 , \31159 , \31161 );
xor \U$30786 ( \31163 , \31152 , \31162 );
xor \U$30787 ( \31164 , \31143 , \31090 );
xnor \U$30788 ( \31165 , \31164 , \31087 );
xor \U$30789 ( \31166 , \30518 , \30208 );
xor \U$30790 ( \31167 , \31166 , \30203 );
not \U$30791 ( \31168 , \31167 );
nand \U$30792 ( \31169 , \31165 , \31168 );
xor \U$30793 ( \31170 , \31100 , \31106 );
xor \U$30794 ( \31171 , \31170 , \31140 );
not \U$30795 ( \31172 , \31171 );
xor \U$30796 ( \31173 , \30216 , \30516 );
xnor \U$30797 ( \31174 , \31173 , \30508 );
nand \U$30798 ( \31175 , \31172 , \31174 );
not \U$30799 ( \31176 , \31175 );
xor \U$30800 ( \31177 , \30550 , \30758 );
xor \U$30801 ( \31178 , \31177 , \31085 );
not \U$30802 ( \31179 , \31178 );
or \U$30803 ( \31180 , \31176 , \31179 );
or \U$30804 ( \31181 , \31172 , \31174 );
nand \U$30805 ( \31182 , \31180 , \31181 );
and \U$30806 ( \31183 , \31169 , \31182 );
nor \U$30807 ( \31184 , \31165 , \31168 );
nor \U$30808 ( \31185 , \31183 , \31184 );
nor \U$30809 ( \31186 , \31163 , \31185 );
xor \U$30810 ( \31187 , \30148 , \30526 );
xor \U$30811 ( \31188 , \31187 , \30533 );
xor \U$30812 ( \31189 , \30548 , \31151 );
and \U$30813 ( \31190 , \31189 , \31162 );
and \U$30814 ( \31191 , \30548 , \31151 );
or \U$30815 ( \31192 , \31190 , \31191 );
nand \U$30816 ( \31193 , \31188 , \31192 );
nand \U$30817 ( \31194 , \31186 , \31193 );
or \U$30818 ( \31195 , \31188 , \31192 );
nand \U$30819 ( \31196 , \31194 , \31195 );
not \U$30820 ( \31197 , \31196 );
or \U$30821 ( \31198 , \30538 , \31197 );
not \U$30822 ( \31199 , \30143 );
not \U$30823 ( \31200 , \30536 );
nand \U$30824 ( \31201 , \31199 , \31200 );
nand \U$30825 ( \31202 , \31198 , \31201 );
not \U$30826 ( \31203 , \31202 );
or \U$30827 ( \31204 , \30141 , \31203 );
or \U$30828 ( \31205 , \29597 , \30138 );
nand \U$30829 ( \31206 , \31204 , \31205 );
not \U$30830 ( \31207 , \31206 );
not \U$30831 ( \31208 , \30806 );
not \U$30832 ( \31209 , \30795 );
or \U$30833 ( \31210 , \31208 , \31209 );
nand \U$30834 ( \31211 , \30807 , \30794 );
nand \U$30835 ( \31212 , \31210 , \31211 );
and \U$30836 ( \31213 , \31212 , \30933 );
not \U$30837 ( \31214 , \31212 );
not \U$30838 ( \31215 , \30933 );
and \U$30839 ( \31216 , \31214 , \31215 );
nor \U$30840 ( \31217 , \31213 , \31216 );
not \U$30841 ( \31218 , \2784 );
and \U$30842 ( \31219 , RIc226890_29, \9321 );
not \U$30843 ( \31220 , RIc226890_29);
and \U$30844 ( \31221 , \31220 , \30573 );
or \U$30845 ( \31222 , \31219 , \31221 );
not \U$30846 ( \31223 , \31222 );
or \U$30847 ( \31224 , \31218 , \31223 );
nand \U$30848 ( \31225 , \30854 , \9142 );
nand \U$30849 ( \31226 , \31224 , \31225 );
not \U$30850 ( \31227 , \4383 );
not \U$30851 ( \31228 , RIc2265c0_35);
not \U$30852 ( \31229 , \28026 );
or \U$30853 ( \31230 , \31228 , \31229 );
nand \U$30854 ( \31231 , \9211 , \3620 );
nand \U$30855 ( \31232 , \31230 , \31231 );
not \U$30856 ( \31233 , \31232 );
or \U$30857 ( \31234 , \31227 , \31233 );
not \U$30858 ( \31235 , RIc2265c0_35);
not \U$30859 ( \31236 , \9046 );
or \U$30860 ( \31237 , \31235 , \31236 );
nand \U$30861 ( \31238 , \9051 , \4376 );
nand \U$30862 ( \31239 , \31237 , \31238 );
nand \U$30863 ( \31240 , \31239 , \4381 );
nand \U$30864 ( \31241 , \31234 , \31240 );
xor \U$30865 ( \31242 , \31226 , \31241 );
not \U$30866 ( \31243 , \9534 );
not \U$30867 ( \31244 , RIc225f30_49);
not \U$30868 ( \31245 , \5216 );
or \U$30869 ( \31246 , \31244 , \31245 );
nand \U$30870 ( \31247 , \18459 , \9549 );
nand \U$30871 ( \31248 , \31246 , \31247 );
not \U$30872 ( \31249 , \31248 );
or \U$30873 ( \31250 , \31243 , \31249 );
not \U$30874 ( \31251 , RIc225f30_49);
not \U$30875 ( \31252 , \10220 );
or \U$30876 ( \31253 , \31251 , \31252 );
nand \U$30877 ( \31254 , \4407 , \9549 );
nand \U$30878 ( \31255 , \31253 , \31254 );
nand \U$30879 ( \31256 , \31255 , \9552 );
nand \U$30880 ( \31257 , \31250 , \31256 );
and \U$30881 ( \31258 , \31242 , \31257 );
and \U$30882 ( \31259 , \31226 , \31241 );
or \U$30883 ( \31260 , \31258 , \31259 );
or \U$30884 ( \31261 , RIc226bd8_22, RIc226b60_23);
nand \U$30885 ( \31262 , \31261 , \18367 );
and \U$30886 ( \31263 , RIc226bd8_22, RIc226b60_23);
nor \U$30887 ( \31264 , \31263 , \2383 );
and \U$30888 ( \31265 , \31262 , \31264 );
not \U$30889 ( \31266 , \2367 );
not \U$30890 ( \31267 , \30831 );
or \U$30891 ( \31268 , \31266 , \31267 );
or \U$30892 ( \31269 , \18367 , \2370 );
or \U$30893 ( \31270 , \18181 , RIc226c50_21);
nand \U$30894 ( \31271 , \31269 , \31270 );
nand \U$30895 ( \31272 , \31271 , \2391 );
nand \U$30896 ( \31273 , \31268 , \31272 );
xor \U$30897 ( \31274 , \31265 , \31273 );
not \U$30898 ( \31275 , \1930 );
not \U$30899 ( \31276 , \30840 );
or \U$30900 ( \31277 , \31275 , \31276 );
not \U$30901 ( \31278 , RIc226b60_23);
not \U$30902 ( \31279 , \17613 );
or \U$30903 ( \31280 , \31278 , \31279 );
not \U$30904 ( \31281 , \30679 );
nand \U$30905 ( \31282 , \31281 , \1927 );
nand \U$30906 ( \31283 , \31280 , \31282 );
nand \U$30907 ( \31284 , \31283 , \1914 );
nand \U$30908 ( \31285 , \31277 , \31284 );
xor \U$30909 ( \31286 , \31274 , \31285 );
not \U$30910 ( \31287 , \2138 );
not \U$30911 ( \31288 , RIc226980_27);
not \U$30912 ( \31289 , \16492 );
or \U$30913 ( \31290 , \31288 , \31289 );
nand \U$30914 ( \31291 , \20406 , \2150 );
nand \U$30915 ( \31292 , \31290 , \31291 );
not \U$30916 ( \31293 , \31292 );
or \U$30917 ( \31294 , \31287 , \31293 );
not \U$30918 ( \31295 , RIc226980_27);
not \U$30919 ( \31296 , \27990 );
or \U$30920 ( \31297 , \31295 , \31296 );
nand \U$30921 ( \31298 , \29423 , \2133 );
nand \U$30922 ( \31299 , \31297 , \31298 );
nand \U$30923 ( \31300 , \31299 , \2154 );
nand \U$30924 ( \31301 , \31294 , \31300 );
and \U$30925 ( \31302 , \31286 , \31301 );
and \U$30926 ( \31303 , \31274 , \31285 );
or \U$30927 ( \31304 , \31302 , \31303 );
not \U$30928 ( \31305 , \6307 );
not \U$30929 ( \31306 , RIc2263e0_39);
not \U$30930 ( \31307 , \8807 );
or \U$30931 ( \31308 , \31306 , \31307 );
nand \U$30932 ( \31309 , \10859 , \5498 );
nand \U$30933 ( \31310 , \31308 , \31309 );
not \U$30934 ( \31311 , \31310 );
or \U$30935 ( \31312 , \31305 , \31311 );
not \U$30936 ( \31313 , RIc2263e0_39);
not \U$30937 ( \31314 , \11565 );
or \U$30938 ( \31315 , \31313 , \31314 );
nand \U$30939 ( \31316 , \8952 , \8998 );
nand \U$30940 ( \31317 , \31315 , \31316 );
nand \U$30941 ( \31318 , \31317 , \6689 );
nand \U$30942 ( \31319 , \31312 , \31318 );
xor \U$30943 ( \31320 , \31304 , \31319 );
not \U$30944 ( \31321 , \9444 );
not \U$30945 ( \31322 , RIc225e40_51);
not \U$30946 ( \31323 , \4046 );
or \U$30947 ( \31324 , \31322 , \31323 );
nand \U$30948 ( \31325 , \3640 , \22140 );
nand \U$30949 ( \31326 , \31324 , \31325 );
not \U$30950 ( \31327 , \31326 );
or \U$30951 ( \31328 , \31321 , \31327 );
not \U$30952 ( \31329 , RIc225e40_51);
not \U$30953 ( \31330 , \13525 );
or \U$30954 ( \31331 , \31329 , \31330 );
nand \U$30955 ( \31332 , \13528 , \12423 );
nand \U$30956 ( \31333 , \31331 , \31332 );
nand \U$30957 ( \31334 , \31333 , \9459 );
nand \U$30958 ( \31335 , \31328 , \31334 );
and \U$30959 ( \31336 , \31320 , \31335 );
and \U$30960 ( \31337 , \31304 , \31319 );
or \U$30961 ( \31338 , \31336 , \31337 );
xor \U$30962 ( \31339 , \31260 , \31338 );
and \U$30963 ( \31340 , \31265 , \31273 );
not \U$30964 ( \31341 , \2195 );
not \U$30965 ( \31342 , RIc226a70_25);
not \U$30966 ( \31343 , \20693 );
or \U$30967 ( \31344 , \31342 , \31343 );
nand \U$30968 ( \31345 , \20694 , \2190 );
nand \U$30969 ( \31346 , \31344 , \31345 );
not \U$30970 ( \31347 , \31346 );
or \U$30971 ( \31348 , \31341 , \31347 );
nand \U$30972 ( \31349 , \2172 , \30692 );
nand \U$30973 ( \31350 , \31348 , \31349 );
xor \U$30974 ( \31351 , \31340 , \31350 );
not \U$30975 ( \31352 , \2154 );
not \U$30976 ( \31353 , \30869 );
or \U$30977 ( \31354 , \31352 , \31353 );
nand \U$30978 ( \31355 , \2138 , \31299 );
nand \U$30979 ( \31356 , \31354 , \31355 );
xor \U$30980 ( \31357 , \31351 , \31356 );
not \U$30981 ( \31358 , \11697 );
not \U$30982 ( \31359 , RIc225c60_55);
not \U$30983 ( \31360 , \9651 );
or \U$30984 ( \31361 , \31359 , \31360 );
nand \U$30985 ( \31362 , \4500 , \8767 );
nand \U$30986 ( \31363 , \31361 , \31362 );
not \U$30987 ( \31364 , \31363 );
or \U$30988 ( \31365 , \31358 , \31364 );
not \U$30989 ( \31366 , RIc225c60_55);
not \U$30990 ( \31367 , \9188 );
or \U$30991 ( \31368 , \31366 , \31367 );
nand \U$30992 ( \31369 , \9805 , \11108 );
nand \U$30993 ( \31370 , \31368 , \31369 );
nand \U$30994 ( \31371 , \31370 , \11038 );
nand \U$30995 ( \31372 , \31365 , \31371 );
xor \U$30996 ( \31373 , \31357 , \31372 );
not \U$30997 ( \31374 , \20862 );
not \U$30998 ( \31375 , RIc225990_61);
not \U$30999 ( \31376 , \9361 );
or \U$31000 ( \31377 , \31375 , \31376 );
nand \U$31001 ( \31378 , \9360 , \10338 );
nand \U$31002 ( \31379 , \31377 , \31378 );
not \U$31003 ( \31380 , \31379 );
or \U$31004 ( \31381 , \31374 , \31380 );
not \U$31005 ( \31382 , RIc225990_61);
not \U$31006 ( \31383 , \3035 );
or \U$31007 ( \31384 , \31382 , \31383 );
nand \U$31008 ( \31385 , \3036 , \12806 );
nand \U$31009 ( \31386 , \31384 , \31385 );
nand \U$31010 ( \31387 , \31386 , \15719 );
nand \U$31011 ( \31388 , \31381 , \31387 );
and \U$31012 ( \31389 , \31373 , \31388 );
and \U$31013 ( \31390 , \31357 , \31372 );
or \U$31014 ( \31391 , \31389 , \31390 );
and \U$31015 ( \31392 , \31339 , \31391 );
and \U$31016 ( \31393 , \31260 , \31338 );
or \U$31017 ( \31394 , \31392 , \31393 );
not \U$31018 ( \31395 , \31394 );
not \U$31019 ( \31396 , \9534 );
not \U$31020 ( \31397 , \31255 );
or \U$31021 ( \31398 , \31396 , \31397 );
nand \U$31022 ( \31399 , \30660 , \9552 );
nand \U$31023 ( \31400 , \31398 , \31399 );
not \U$31024 ( \31401 , \31400 );
not \U$31025 ( \31402 , \12698 );
not \U$31026 ( \31403 , \31402 );
not \U$31027 ( \31404 , \9100 );
and \U$31028 ( \31405 , \31403 , \31404 );
and \U$31029 ( \31406 , \15645 , \22795 );
nor \U$31030 ( \31407 , \31405 , \31406 );
not \U$31031 ( \31408 , \31407 );
not \U$31032 ( \31409 , \9383 );
and \U$31033 ( \31410 , \31408 , \31409 );
and \U$31034 ( \31411 , \30648 , \9398 );
nor \U$31035 ( \31412 , \31410 , \31411 );
not \U$31036 ( \31413 , \31412 );
not \U$31037 ( \31414 , \31413 );
or \U$31038 ( \31415 , \31401 , \31414 );
or \U$31039 ( \31416 , \31413 , \31400 );
not \U$31040 ( \31417 , \10001 );
not \U$31041 ( \31418 , RIc226020_47);
not \U$31042 ( \31419 , \10161 );
or \U$31043 ( \31420 , \31418 , \31419 );
nand \U$31044 ( \31421 , \5666 , \11607 );
nand \U$31045 ( \31422 , \31420 , \31421 );
not \U$31046 ( \31423 , \31422 );
or \U$31047 ( \31424 , \31417 , \31423 );
not \U$31048 ( \31425 , \30623 );
nand \U$31049 ( \31426 , \31425 , \12304 );
nand \U$31050 ( \31427 , \31424 , \31426 );
nand \U$31051 ( \31428 , \31416 , \31427 );
nand \U$31052 ( \31429 , \31415 , \31428 );
xor \U$31053 ( \31430 , \30674 , \30685 );
xor \U$31054 ( \31431 , \31430 , \30697 );
not \U$31055 ( \31432 , \9110 );
not \U$31056 ( \31433 , RIc226200_43);
not \U$31057 ( \31434 , \10142 );
or \U$31058 ( \31435 , \31433 , \31434 );
nand \U$31059 ( \31436 , \10310 , \9125 );
nand \U$31060 ( \31437 , \31435 , \31436 );
not \U$31061 ( \31438 , \31437 );
or \U$31062 ( \31439 , \31432 , \31438 );
nand \U$31063 ( \31440 , \30636 , \9129 );
nand \U$31064 ( \31441 , \31439 , \31440 );
xor \U$31065 ( \31442 , \31431 , \31441 );
not \U$31066 ( \31443 , \9690 );
not \U$31067 ( \31444 , RIc2262f0_41);
not \U$31068 ( \31445 , \12724 );
or \U$31069 ( \31446 , \31444 , \31445 );
not \U$31070 ( \31447 , \8857 );
nand \U$31071 ( \31448 , \31447 , \6303 );
nand \U$31072 ( \31449 , \31446 , \31448 );
not \U$31073 ( \31450 , \31449 );
or \U$31074 ( \31451 , \31443 , \31450 );
nand \U$31075 ( \31452 , \30716 , \9705 );
nand \U$31076 ( \31453 , \31451 , \31452 );
and \U$31077 ( \31454 , \31442 , \31453 );
and \U$31078 ( \31455 , \31431 , \31441 );
or \U$31079 ( \31456 , \31454 , \31455 );
and \U$31080 ( \31457 , \31429 , \31456 );
not \U$31081 ( \31458 , \31429 );
not \U$31082 ( \31459 , \31456 );
and \U$31083 ( \31460 , \31458 , \31459 );
nor \U$31084 ( \31461 , \31457 , \31460 );
not \U$31085 ( \31462 , \16891 );
not \U$31086 ( \31463 , RIc2258a0_63);
not \U$31087 ( \31464 , \24302 );
or \U$31088 ( \31465 , \31463 , \31464 );
not \U$31089 ( \31466 , RIc2258a0_63);
nand \U$31090 ( \31467 , \2014 , \31466 );
nand \U$31091 ( \31468 , \31465 , \31467 );
not \U$31092 ( \31469 , \31468 );
or \U$31093 ( \31470 , \31462 , \31469 );
nand \U$31094 ( \31471 , \31018 , RIc225828_64);
nand \U$31095 ( \31472 , \31470 , \31471 );
buf \U$31096 ( \31473 , \31472 );
not \U$31097 ( \31474 , \31473 );
not \U$31098 ( \31475 , \11974 );
not \U$31099 ( \31476 , \31003 );
or \U$31100 ( \31477 , \31475 , \31476 );
not \U$31101 ( \31478 , RIc225b70_57);
not \U$31102 ( \31479 , \3010 );
or \U$31103 ( \31480 , \31478 , \31479 );
nand \U$31104 ( \31481 , \4240 , \11033 );
nand \U$31105 ( \31482 , \31480 , \31481 );
nand \U$31106 ( \31483 , \31482 , \11965 );
nand \U$31107 ( \31484 , \31477 , \31483 );
not \U$31108 ( \31485 , \31484 );
or \U$31109 ( \31486 , \31474 , \31485 );
or \U$31110 ( \31487 , \31484 , \31473 );
not \U$31111 ( \31488 , \4383 );
not \U$31112 ( \31489 , \30982 );
or \U$31113 ( \31490 , \31488 , \31489 );
nand \U$31114 ( \31491 , \31232 , \4381 );
nand \U$31115 ( \31492 , \31490 , \31491 );
nand \U$31116 ( \31493 , \31487 , \31492 );
nand \U$31117 ( \31494 , \31486 , \31493 );
not \U$31118 ( \31495 , \31494 );
and \U$31119 ( \31496 , \31461 , \31495 );
not \U$31120 ( \31497 , \31461 );
and \U$31121 ( \31498 , \31497 , \31494 );
nor \U$31122 ( \31499 , \31496 , \31498 );
not \U$31123 ( \31500 , \31499 );
not \U$31124 ( \31501 , \31500 );
or \U$31125 ( \31502 , \31395 , \31501 );
not \U$31126 ( \31503 , \31394 );
nand \U$31127 ( \31504 , \31503 , \31499 );
xor \U$31128 ( \31505 , \31431 , \31441 );
xor \U$31129 ( \31506 , \31505 , \31453 );
not \U$31130 ( \31507 , \5509 );
not \U$31131 ( \31508 , RIc2264d0_37);
not \U$31132 ( \31509 , \8910 );
or \U$31133 ( \31510 , \31508 , \31509 );
nand \U$31134 ( \31511 , \9786 , \12522 );
nand \U$31135 ( \31512 , \31510 , \31511 );
not \U$31136 ( \31513 , \31512 );
or \U$31137 ( \31514 , \31507 , \31513 );
and \U$31138 ( \31515 , \11094 , RIc2264d0_37);
not \U$31139 ( \31516 , \11094 );
and \U$31140 ( \31517 , \31516 , \5504 );
or \U$31141 ( \31518 , \31515 , \31517 );
nand \U$31142 ( \31519 , \31518 , \5519 );
nand \U$31143 ( \31520 , \31514 , \31519 );
not \U$31144 ( \31521 , \9705 );
not \U$31145 ( \31522 , \31449 );
or \U$31146 ( \31523 , \31521 , \31522 );
not \U$31147 ( \31524 , RIc2262f0_41);
not \U$31148 ( \31525 , \9897 );
or \U$31149 ( \31526 , \31524 , \31525 );
nand \U$31150 ( \31527 , \20216 , \10679 );
nand \U$31151 ( \31528 , \31526 , \31527 );
nand \U$31152 ( \31529 , \31528 , \9690 );
nand \U$31153 ( \31530 , \31523 , \31529 );
xor \U$31154 ( \31531 , \31520 , \31530 );
not \U$31155 ( \31532 , \11965 );
not \U$31156 ( \31533 , RIc225b70_57);
not \U$31157 ( \31534 , \11068 );
or \U$31158 ( \31535 , \31533 , \31534 );
nand \U$31159 ( \31536 , \15490 , \12475 );
nand \U$31160 ( \31537 , \31535 , \31536 );
not \U$31161 ( \31538 , \31537 );
or \U$31162 ( \31539 , \31532 , \31538 );
nand \U$31163 ( \31540 , \31482 , \11974 );
nand \U$31164 ( \31541 , \31539 , \31540 );
and \U$31165 ( \31542 , \31531 , \31541 );
and \U$31166 ( \31543 , \31520 , \31530 );
or \U$31167 ( \31544 , \31542 , \31543 );
xor \U$31168 ( \31545 , \31506 , \31544 );
not \U$31169 ( \31546 , \16891 );
not \U$31170 ( \31547 , RIc2258a0_63);
not \U$31171 ( \31548 , \2587 );
or \U$31172 ( \31549 , \31547 , \31548 );
nand \U$31173 ( \31550 , \5809 , \31466 );
nand \U$31174 ( \31551 , \31549 , \31550 );
not \U$31175 ( \31552 , \31551 );
or \U$31176 ( \31553 , \31546 , \31552 );
nand \U$31177 ( \31554 , \31468 , RIc225828_64);
nand \U$31178 ( \31555 , \31553 , \31554 );
not \U$31179 ( \31556 , \9488 );
not \U$31180 ( \31557 , RIc225d50_53);
not \U$31181 ( \31558 , \17703 );
or \U$31182 ( \31559 , \31557 , \31558 );
not \U$31183 ( \31560 , \3726 );
nand \U$31184 ( \31561 , \31560 , \11391 );
nand \U$31185 ( \31562 , \31559 , \31561 );
not \U$31186 ( \31563 , \31562 );
or \U$31187 ( \31564 , \31556 , \31563 );
not \U$31188 ( \31565 , RIc225d50_53);
not \U$31189 ( \31566 , \5160 );
not \U$31190 ( \31567 , \31566 );
or \U$31191 ( \31568 , \31565 , \31567 );
nand \U$31192 ( \31569 , \22561 , \11585 );
nand \U$31193 ( \31570 , \31568 , \31569 );
nand \U$31194 ( \31571 , \31570 , \8788 );
nand \U$31195 ( \31572 , \31564 , \31571 );
xor \U$31196 ( \31573 , \31555 , \31572 );
not \U$31197 ( \31574 , \15164 );
and \U$31198 ( \31575 , RIc225a80_59, \3810 );
not \U$31199 ( \31576 , RIc225a80_59);
and \U$31200 ( \31577 , \31576 , \4564 );
or \U$31201 ( \31578 , \31575 , \31577 );
not \U$31202 ( \31579 , \31578 );
or \U$31203 ( \31580 , \31574 , \31579 );
and \U$31204 ( \31581 , RIc225a80_59, \2501 );
not \U$31205 ( \31582 , RIc225a80_59);
and \U$31206 ( \31583 , \31582 , \2500 );
or \U$31207 ( \31584 , \31581 , \31583 );
nand \U$31208 ( \31585 , \31584 , \18037 );
nand \U$31209 ( \31586 , \31580 , \31585 );
and \U$31210 ( \31587 , \31573 , \31586 );
and \U$31211 ( \31588 , \31555 , \31572 );
or \U$31212 ( \31589 , \31587 , \31588 );
and \U$31213 ( \31590 , \31545 , \31589 );
and \U$31214 ( \31591 , \31506 , \31544 );
or \U$31215 ( \31592 , \31590 , \31591 );
nand \U$31216 ( \31593 , \31504 , \31592 );
nand \U$31217 ( \31594 , \31502 , \31593 );
not \U$31218 ( \31595 , \31594 );
xor \U$31219 ( \31596 , \30811 , \30913 );
xor \U$31220 ( \31597 , \31596 , \30930 );
not \U$31221 ( \31598 , \31597 );
xor \U$31222 ( \31599 , \30861 , \30899 );
xor \U$31223 ( \31600 , \31599 , \30910 );
not \U$31224 ( \31601 , \31058 );
not \U$31225 ( \31602 , \31074 );
and \U$31226 ( \31603 , \31601 , \31602 );
and \U$31227 ( \31604 , \31058 , \31074 );
nor \U$31228 ( \31605 , \31603 , \31604 );
xnor \U$31229 ( \31606 , \31605 , \31069 );
or \U$31230 ( \31607 , \31600 , \31606 );
xor \U$31231 ( \31608 , \30822 , \30833 );
xor \U$31232 ( \31609 , \31608 , \30844 );
not \U$31233 ( \31610 , \2697 );
not \U$31234 ( \31611 , RIc2267a0_31);
not \U$31235 ( \31612 , \9276 );
or \U$31236 ( \31613 , \31611 , \31612 );
nand \U$31237 ( \31614 , \9275 , \9159 );
nand \U$31238 ( \31615 , \31613 , \31614 );
not \U$31239 ( \31616 , \31615 );
or \U$31240 ( \31617 , \31610 , \31616 );
nand \U$31241 ( \31618 , \30880 , \2710 );
nand \U$31242 ( \31619 , \31617 , \31618 );
xor \U$31243 ( \31620 , \31609 , \31619 );
not \U$31244 ( \31621 , \3631 );
not \U$31245 ( \31622 , \30895 );
or \U$31246 ( \31623 , \31621 , \31622 );
not \U$31247 ( \31624 , RIc2266b0_33);
not \U$31248 ( \31625 , \10814 );
or \U$31249 ( \31626 , \31624 , \31625 );
nand \U$31250 ( \31627 , \10110 , \6890 );
nand \U$31251 ( \31628 , \31626 , \31627 );
nand \U$31252 ( \31629 , \31628 , \3629 );
nand \U$31253 ( \31630 , \31623 , \31629 );
and \U$31254 ( \31631 , \31620 , \31630 );
and \U$31255 ( \31632 , \31609 , \31619 );
or \U$31256 ( \31633 , \31631 , \31632 );
xor \U$31257 ( \31634 , \30871 , \30884 );
xor \U$31258 ( \31635 , \30897 , \31634 );
xor \U$31259 ( \31636 , \31633 , \31635 );
not \U$31260 ( \31637 , \9110 );
not \U$31261 ( \31638 , RIc226200_43);
not \U$31262 ( \31639 , \8887 );
or \U$31263 ( \31640 , \31638 , \31639 );
nand \U$31264 ( \31641 , \17582 , \9106 );
nand \U$31265 ( \31642 , \31640 , \31641 );
not \U$31266 ( \31643 , \31642 );
or \U$31267 ( \31644 , \31637 , \31643 );
nand \U$31268 ( \31645 , \31437 , \9205 );
nand \U$31269 ( \31646 , \31644 , \31645 );
not \U$31270 ( \31647 , \9934 );
not \U$31271 ( \31648 , RIc226110_45);
not \U$31272 ( \31649 , \23758 );
or \U$31273 ( \31650 , \31648 , \31649 );
nand \U$31274 ( \31651 , \9740 , \9100 );
nand \U$31275 ( \31652 , \31650 , \31651 );
not \U$31276 ( \31653 , \31652 );
or \U$31277 ( \31654 , \31647 , \31653 );
not \U$31278 ( \31655 , \31407 );
nand \U$31279 ( \31656 , \31655 , \9398 );
nand \U$31280 ( \31657 , \31654 , \31656 );
or \U$31281 ( \31658 , \31646 , \31657 );
not \U$31282 ( \31659 , \9619 );
not \U$31283 ( \31660 , \31422 );
or \U$31284 ( \31661 , \31659 , \31660 );
not \U$31285 ( \31662 , RIc226020_47);
not \U$31286 ( \31663 , \10170 );
or \U$31287 ( \31664 , \31662 , \31663 );
nand \U$31288 ( \31665 , \6071 , \9373 );
nand \U$31289 ( \31666 , \31664 , \31665 );
nand \U$31290 ( \31667 , \10001 , \31666 );
nand \U$31291 ( \31668 , \31661 , \31667 );
nand \U$31292 ( \31669 , \31658 , \31668 );
nand \U$31293 ( \31670 , \31657 , \31646 );
nand \U$31294 ( \31671 , \31669 , \31670 );
and \U$31295 ( \31672 , \31636 , \31671 );
and \U$31296 ( \31673 , \31633 , \31635 );
or \U$31297 ( \31674 , \31672 , \31673 );
and \U$31298 ( \31675 , \31607 , \31674 );
and \U$31299 ( \31676 , \31600 , \31606 );
nor \U$31300 ( \31677 , \31675 , \31676 );
nand \U$31301 ( \31678 , \31598 , \31677 );
not \U$31302 ( \31679 , \31678 );
or \U$31303 ( \31680 , \31595 , \31679 );
not \U$31304 ( \31681 , \31677 );
nand \U$31305 ( \31682 , \31681 , \31597 );
nand \U$31306 ( \31683 , \31680 , \31682 );
xor \U$31307 ( \31684 , \31217 , \31683 );
xor \U$31308 ( \31685 , \30556 , \30583 );
xor \U$31309 ( \31686 , \31685 , \30590 );
xor \U$31310 ( \31687 , \30251 , \30227 );
xor \U$31311 ( \31688 , \31687 , \30238 );
xor \U$31312 ( \31689 , \31686 , \31688 );
xor \U$31313 ( \31690 , \30558 , \30567 );
xor \U$31314 ( \31691 , \31690 , \30580 );
xor \U$31315 ( \31692 , \30603 , \30614 );
xor \U$31316 ( \31693 , \31692 , \30625 );
xor \U$31317 ( \31694 , \31691 , \31693 );
not \U$31318 ( \31695 , \6688 );
not \U$31319 ( \31696 , \31310 );
or \U$31320 ( \31697 , \31695 , \31696 );
nand \U$31321 ( \31698 , \30706 , \6307 );
nand \U$31322 ( \31699 , \31697 , \31698 );
not \U$31323 ( \31700 , \31699 );
not \U$31324 ( \31701 , \5509 );
not \U$31325 ( \31702 , \31518 );
or \U$31326 ( \31703 , \31701 , \31702 );
nand \U$31327 ( \31704 , \30992 , \5519 );
nand \U$31328 ( \31705 , \31703 , \31704 );
not \U$31329 ( \31706 , \31705 );
or \U$31330 ( \31707 , \31700 , \31706 );
or \U$31331 ( \31708 , \31705 , \31699 );
xor \U$31332 ( \31709 , \31340 , \31350 );
and \U$31333 ( \31710 , \31709 , \31356 );
and \U$31334 ( \31711 , \31340 , \31350 );
or \U$31335 ( \31712 , \31710 , \31711 );
nand \U$31336 ( \31713 , \31708 , \31712 );
nand \U$31337 ( \31714 , \31707 , \31713 );
and \U$31338 ( \31715 , \31694 , \31714 );
and \U$31339 ( \31716 , \31691 , \31693 );
or \U$31340 ( \31717 , \31715 , \31716 );
and \U$31341 ( \31718 , \31689 , \31717 );
and \U$31342 ( \31719 , \31686 , \31688 );
or \U$31343 ( \31720 , \31718 , \31719 );
xor \U$31344 ( \31721 , \31130 , \31132 );
xor \U$31345 ( \31722 , \31721 , \31135 );
xor \U$31346 ( \31723 , \31720 , \31722 );
xor \U$31347 ( \31724 , \30628 , \30666 );
xor \U$31348 ( \31725 , \31724 , \30723 );
not \U$31349 ( \31726 , \31429 );
not \U$31350 ( \31727 , \31494 );
or \U$31351 ( \31728 , \31726 , \31727 );
or \U$31352 ( \31729 , \31494 , \31429 );
nand \U$31353 ( \31730 , \31729 , \31456 );
nand \U$31354 ( \31731 , \31728 , \31730 );
xor \U$31355 ( \31732 , \31725 , \31731 );
xor \U$31356 ( \31733 , \30700 , \30710 );
xor \U$31357 ( \31734 , \31733 , \30720 );
xor \U$31358 ( \31735 , \30640 , \30663 );
xnor \U$31359 ( \31736 , \31735 , \30650 );
xor \U$31360 ( \31737 , \31734 , \31736 );
not \U$31361 ( \31738 , \11118 );
not \U$31362 ( \31739 , \31370 );
or \U$31363 ( \31740 , \31738 , \31739 );
nand \U$31364 ( \31741 , \31042 , \11038 );
nand \U$31365 ( \31742 , \31740 , \31741 );
not \U$31366 ( \31743 , \9488 );
not \U$31367 ( \31744 , \31570 );
or \U$31368 ( \31745 , \31743 , \31744 );
nand \U$31369 ( \31746 , \31064 , \8788 );
nand \U$31370 ( \31747 , \31745 , \31746 );
xor \U$31371 ( \31748 , \31742 , \31747 );
not \U$31372 ( \31749 , \15719 );
not \U$31373 ( \31750 , \31379 );
or \U$31374 ( \31751 , \31749 , \31750 );
nand \U$31375 ( \31752 , \31029 , \20862 );
nand \U$31376 ( \31753 , \31751 , \31752 );
and \U$31377 ( \31754 , \31748 , \31753 );
and \U$31378 ( \31755 , \31742 , \31747 );
or \U$31379 ( \31756 , \31754 , \31755 );
and \U$31380 ( \31757 , \31737 , \31756 );
and \U$31381 ( \31758 , \31734 , \31736 );
or \U$31382 ( \31759 , \31757 , \31758 );
and \U$31383 ( \31760 , \31732 , \31759 );
and \U$31384 ( \31761 , \31725 , \31731 );
or \U$31385 ( \31762 , \31760 , \31761 );
xor \U$31386 ( \31763 , \31723 , \31762 );
xor \U$31387 ( \31764 , \31684 , \31763 );
xor \U$31388 ( \31765 , \31686 , \31688 );
xor \U$31389 ( \31766 , \31765 , \31717 );
xor \U$31390 ( \31767 , \31691 , \31693 );
xor \U$31391 ( \31768 , \31767 , \31714 );
xor \U$31392 ( \31769 , \31400 , \31412 );
xor \U$31393 ( \31770 , \31769 , \31427 );
not \U$31394 ( \31771 , \31770 );
xor \U$31395 ( \31772 , \31492 , \31472 );
xnor \U$31396 ( \31773 , \31772 , \31484 );
not \U$31397 ( \31774 , \31773 );
or \U$31398 ( \31775 , \31771 , \31774 );
xor \U$31399 ( \31776 , \31699 , \31712 );
xor \U$31400 ( \31777 , \31776 , \31705 );
nand \U$31401 ( \31778 , \31775 , \31777 );
not \U$31402 ( \31779 , \31770 );
not \U$31403 ( \31780 , \31773 );
nand \U$31404 ( \31781 , \31779 , \31780 );
nand \U$31405 ( \31782 , \31778 , \31781 );
xor \U$31406 ( \31783 , \31768 , \31782 );
xor \U$31407 ( \31784 , \31734 , \31736 );
xor \U$31408 ( \31785 , \31784 , \31756 );
and \U$31409 ( \31786 , \31783 , \31785 );
and \U$31410 ( \31787 , \31768 , \31782 );
or \U$31411 ( \31788 , \31786 , \31787 );
xor \U$31412 ( \31789 , \31766 , \31788 );
xor \U$31413 ( \31790 , \31725 , \31731 );
xor \U$31414 ( \31791 , \31790 , \31759 );
xor \U$31415 ( \31792 , \31789 , \31791 );
xor \U$31416 ( \31793 , \31609 , \31619 );
xor \U$31417 ( \31794 , \31793 , \31630 );
xor \U$31418 ( \31795 , \31226 , \31241 );
xor \U$31419 ( \31796 , \31795 , \31257 );
xor \U$31420 ( \31797 , \31794 , \31796 );
not \U$31421 ( \31798 , \9934 );
not \U$31422 ( \31799 , RIc226110_45);
not \U$31423 ( \31800 , \15699 );
or \U$31424 ( \31801 , \31799 , \31800 );
nand \U$31425 ( \31802 , \15700 , \9100 );
nand \U$31426 ( \31803 , \31801 , \31802 );
not \U$31427 ( \31804 , \31803 );
or \U$31428 ( \31805 , \31798 , \31804 );
nand \U$31429 ( \31806 , \31652 , \15183 );
nand \U$31430 ( \31807 , \31805 , \31806 );
not \U$31431 ( \31808 , \10953 );
not \U$31432 ( \31809 , \31666 );
or \U$31433 ( \31810 , \31808 , \31809 );
not \U$31434 ( \31811 , RIc226020_47);
not \U$31435 ( \31812 , \22928 );
or \U$31436 ( \31813 , \31811 , \31812 );
nand \U$31437 ( \31814 , \27798 , \11607 );
nand \U$31438 ( \31815 , \31813 , \31814 );
nand \U$31439 ( \31816 , \31815 , \9641 );
nand \U$31440 ( \31817 , \31810 , \31816 );
or \U$31441 ( \31818 , \31807 , \31817 );
not \U$31442 ( \31819 , \9552 );
not \U$31443 ( \31820 , \31248 );
or \U$31444 ( \31821 , \31819 , \31820 );
not \U$31445 ( \31822 , RIc225f30_49);
not \U$31446 ( \31823 , \20656 );
or \U$31447 ( \31824 , \31822 , \31823 );
nand \U$31448 ( \31825 , \19859 , \11289 );
nand \U$31449 ( \31826 , \31824 , \31825 );
nand \U$31450 ( \31827 , \31826 , \10445 );
nand \U$31451 ( \31828 , \31821 , \31827 );
nand \U$31452 ( \31829 , \31818 , \31828 );
nand \U$31453 ( \31830 , \31807 , \31817 );
nand \U$31454 ( \31831 , \31829 , \31830 );
and \U$31455 ( \31832 , \31797 , \31831 );
and \U$31456 ( \31833 , \31794 , \31796 );
or \U$31457 ( \31834 , \31832 , \31833 );
xor \U$31458 ( \31835 , \31260 , \31338 );
xor \U$31459 ( \31836 , \31835 , \31391 );
xor \U$31460 ( \31837 , \31834 , \31836 );
xor \U$31461 ( \31838 , \31304 , \31319 );
xor \U$31462 ( \31839 , \31838 , \31335 );
not \U$31463 ( \31840 , \9690 );
not \U$31464 ( \31841 , RIc2262f0_41);
buf \U$31465 ( \31842 , \8810 );
not \U$31466 ( \31843 , \31842 );
or \U$31467 ( \31844 , \31841 , \31843 );
nand \U$31468 ( \31845 , \8811 , \6303 );
nand \U$31469 ( \31846 , \31844 , \31845 );
not \U$31470 ( \31847 , \31846 );
or \U$31471 ( \31848 , \31840 , \31847 );
nand \U$31472 ( \31849 , \31528 , \9705 );
nand \U$31473 ( \31850 , \31848 , \31849 );
not \U$31474 ( \31851 , \6307 );
not \U$31475 ( \31852 , \31317 );
or \U$31476 ( \31853 , \31851 , \31852 );
not \U$31477 ( \31854 , RIc2263e0_39);
not \U$31478 ( \31855 , \11994 );
not \U$31479 ( \31856 , \31855 );
or \U$31480 ( \31857 , \31854 , \31856 );
nand \U$31481 ( \31858 , \21867 , \8990 );
nand \U$31482 ( \31859 , \31857 , \31858 );
nand \U$31483 ( \31860 , \31859 , \6688 );
nand \U$31484 ( \31861 , \31853 , \31860 );
xor \U$31485 ( \31862 , \31850 , \31861 );
or \U$31486 ( \31863 , RIc226ae8_24, RIc226a70_25);
nand \U$31487 ( \31864 , \31863 , \16248 );
and \U$31488 ( \31865 , RIc226ae8_24, RIc226a70_25);
nor \U$31489 ( \31866 , \31865 , \5637 );
and \U$31490 ( \31867 , \31864 , \31866 );
not \U$31491 ( \31868 , \1930 );
not \U$31492 ( \31869 , RIc226b60_23);
not \U$31493 ( \31870 , \16259 );
or \U$31494 ( \31871 , \31869 , \31870 );
nand \U$31495 ( \31872 , \16256 , \1927 );
nand \U$31496 ( \31873 , \31871 , \31872 );
not \U$31497 ( \31874 , \31873 );
or \U$31498 ( \31875 , \31868 , \31874 );
or \U$31499 ( \31876 , \16248 , \1911 );
or \U$31500 ( \31877 , \21954 , RIc226b60_23);
nand \U$31501 ( \31878 , \31876 , \31877 );
nand \U$31502 ( \31879 , \31878 , \1914 );
nand \U$31503 ( \31880 , \31875 , \31879 );
and \U$31504 ( \31881 , \31867 , \31880 );
not \U$31505 ( \31882 , \2154 );
not \U$31506 ( \31883 , \31292 );
or \U$31507 ( \31884 , \31882 , \31883 );
not \U$31508 ( \31885 , RIc226980_27);
not \U$31509 ( \31886 , \16042 );
or \U$31510 ( \31887 , \31885 , \31886 );
nand \U$31511 ( \31888 , \20694 , \2133 );
nand \U$31512 ( \31889 , \31887 , \31888 );
nand \U$31513 ( \31890 , \31889 , \2138 );
nand \U$31514 ( \31891 , \31884 , \31890 );
xor \U$31515 ( \31892 , \31881 , \31891 );
not \U$31516 ( \31893 , \2086 );
not \U$31517 ( \31894 , \10086 );
and \U$31518 ( \31895 , RIc226890_29, \31894 );
not \U$31519 ( \31896 , RIc226890_29);
and \U$31520 ( \31897 , \31896 , \21175 );
or \U$31521 ( \31898 , \31895 , \31897 );
not \U$31522 ( \31899 , \31898 );
or \U$31523 ( \31900 , \31893 , \31899 );
not \U$31524 ( \31901 , RIc226890_29);
not \U$31525 ( \31902 , \27990 );
or \U$31526 ( \31903 , \31901 , \31902 );
not \U$31527 ( \31904 , RIc226890_29);
nand \U$31528 ( \31905 , \31904 , \20701 );
nand \U$31529 ( \31906 , \31903 , \31905 );
nand \U$31530 ( \31907 , \31906 , \2078 );
nand \U$31531 ( \31908 , \31900 , \31907 );
and \U$31532 ( \31909 , \31892 , \31908 );
and \U$31533 ( \31910 , \31881 , \31891 );
or \U$31534 ( \31911 , \31909 , \31910 );
and \U$31535 ( \31912 , \31862 , \31911 );
and \U$31536 ( \31913 , \31850 , \31861 );
or \U$31537 ( \31914 , \31912 , \31913 );
xor \U$31538 ( \31915 , \31839 , \31914 );
not \U$31539 ( \31916 , \11577 );
not \U$31540 ( \31917 , \31562 );
or \U$31541 ( \31918 , \31916 , \31917 );
not \U$31542 ( \31919 , RIc225d50_53);
not \U$31543 ( \31920 , \4046 );
or \U$31544 ( \31921 , \31919 , \31920 );
nand \U$31545 ( \31922 , \15768 , \8782 );
nand \U$31546 ( \31923 , \31921 , \31922 );
nand \U$31547 ( \31924 , \31923 , \9488 );
nand \U$31548 ( \31925 , \31918 , \31924 );
not \U$31549 ( \31926 , \11117 );
not \U$31550 ( \31927 , RIc225c60_55);
not \U$31551 ( \31928 , \3116 );
or \U$31552 ( \31929 , \31927 , \31928 );
nand \U$31553 ( \31930 , \11320 , \8767 );
nand \U$31554 ( \31931 , \31929 , \31930 );
not \U$31555 ( \31932 , \31931 );
or \U$31556 ( \31933 , \31926 , \31932 );
nand \U$31557 ( \31934 , \31363 , \11038 );
nand \U$31558 ( \31935 , \31933 , \31934 );
xor \U$31559 ( \31936 , \31925 , \31935 );
not \U$31560 ( \31937 , RIc225828_64);
not \U$31561 ( \31938 , \31551 );
or \U$31562 ( \31939 , \31937 , \31938 );
not \U$31563 ( \31940 , RIc2258a0_63);
not \U$31564 ( \31941 , \4803 );
or \U$31565 ( \31942 , \31940 , \31941 );
nand \U$31566 ( \31943 , \22388 , \15620 );
nand \U$31567 ( \31944 , \31942 , \31943 );
nand \U$31568 ( \31945 , \31944 , \16891 );
nand \U$31569 ( \31946 , \31939 , \31945 );
and \U$31570 ( \31947 , \31936 , \31946 );
and \U$31571 ( \31948 , \31925 , \31935 );
or \U$31572 ( \31949 , \31947 , \31948 );
and \U$31573 ( \31950 , \31915 , \31949 );
and \U$31574 ( \31951 , \31839 , \31914 );
or \U$31575 ( \31952 , \31950 , \31951 );
and \U$31576 ( \31953 , \31837 , \31952 );
and \U$31577 ( \31954 , \31834 , \31836 );
or \U$31578 ( \31955 , \31953 , \31954 );
xor \U$31579 ( \31956 , \31633 , \31635 );
xor \U$31580 ( \31957 , \31956 , \31671 );
not \U$31581 ( \31958 , \11974 );
not \U$31582 ( \31959 , \31537 );
or \U$31583 ( \31960 , \31958 , \31959 );
not \U$31584 ( \31961 , RIc225b70_57);
not \U$31585 ( \31962 , \4227 );
or \U$31586 ( \31963 , \31961 , \31962 );
nand \U$31587 ( \31964 , \22197 , \12475 );
nand \U$31588 ( \31965 , \31963 , \31964 );
nand \U$31589 ( \31966 , \31965 , \11965 );
nand \U$31590 ( \31967 , \31960 , \31966 );
not \U$31591 ( \31968 , \31967 );
not \U$31592 ( \31969 , \15719 );
not \U$31593 ( \31970 , RIc225990_61);
not \U$31594 ( \31971 , \2501 );
or \U$31595 ( \31972 , \31970 , \31971 );
nand \U$31596 ( \31973 , \17122 , \12806 );
nand \U$31597 ( \31974 , \31972 , \31973 );
not \U$31598 ( \31975 , \31974 );
or \U$31599 ( \31976 , \31969 , \31975 );
nand \U$31600 ( \31977 , \31386 , \15729 );
nand \U$31601 ( \31978 , \31976 , \31977 );
not \U$31602 ( \31979 , \31978 );
or \U$31603 ( \31980 , \31968 , \31979 );
or \U$31604 ( \31981 , \31978 , \31967 );
not \U$31605 ( \31982 , \5519 );
not \U$31606 ( \31983 , \31512 );
or \U$31607 ( \31984 , \31982 , \31983 );
not \U$31608 ( \31985 , RIc2264d0_37);
not \U$31609 ( \31986 , \28026 );
or \U$31610 ( \31987 , \31985 , \31986 );
not \U$31611 ( \31988 , \11405 );
nand \U$31612 ( \31989 , \31988 , \4371 );
nand \U$31613 ( \31990 , \31987 , \31989 );
nand \U$31614 ( \31991 , \31990 , \5509 );
nand \U$31615 ( \31992 , \31984 , \31991 );
nand \U$31616 ( \31993 , \31981 , \31992 );
nand \U$31617 ( \31994 , \31980 , \31993 );
not \U$31618 ( \31995 , \31994 );
xor \U$31619 ( \31996 , \31520 , \31530 );
xor \U$31620 ( \31997 , \31996 , \31541 );
not \U$31621 ( \31998 , \31997 );
or \U$31622 ( \31999 , \31995 , \31998 );
or \U$31623 ( \32000 , \31994 , \31997 );
xor \U$31624 ( \32001 , \31657 , \31646 );
not \U$31625 ( \32002 , \31668 );
and \U$31626 ( \32003 , \32001 , \32002 );
not \U$31627 ( \32004 , \32001 );
and \U$31628 ( \32005 , \32004 , \31668 );
nor \U$31629 ( \32006 , \32003 , \32005 );
not \U$31630 ( \32007 , \32006 );
nand \U$31631 ( \32008 , \32000 , \32007 );
nand \U$31632 ( \32009 , \31999 , \32008 );
xor \U$31633 ( \32010 , \31957 , \32009 );
xor \U$31634 ( \32011 , \31357 , \31372 );
xor \U$31635 ( \32012 , \32011 , \31388 );
not \U$31636 ( \32013 , \2172 );
not \U$31637 ( \32014 , \31346 );
or \U$31638 ( \32015 , \32013 , \32014 );
not \U$31639 ( \32016 , RIc226a70_25);
not \U$31640 ( \32017 , \15444 );
or \U$31641 ( \32018 , \32016 , \32017 );
nand \U$31642 ( \32019 , \19721 , \1905 );
nand \U$31643 ( \32020 , \32018 , \32019 );
nand \U$31644 ( \32021 , \32020 , \2195 );
nand \U$31645 ( \32022 , \32015 , \32021 );
and \U$31646 ( \32023 , \16248 , \2367 );
not \U$31647 ( \32024 , \1930 );
not \U$31648 ( \32025 , \31283 );
or \U$31649 ( \32026 , \32024 , \32025 );
nand \U$31650 ( \32027 , \31873 , \1914 );
nand \U$31651 ( \32028 , \32026 , \32027 );
xor \U$31652 ( \32029 , \32023 , \32028 );
not \U$31653 ( \32030 , \2194 );
not \U$31654 ( \32031 , RIc226a70_25);
not \U$31655 ( \32032 , \15630 );
or \U$31656 ( \32033 , \32031 , \32032 );
nand \U$31657 ( \32034 , \12845 , \1905 );
nand \U$31658 ( \32035 , \32033 , \32034 );
not \U$31659 ( \32036 , \32035 );
or \U$31660 ( \32037 , \32030 , \32036 );
nand \U$31661 ( \32038 , \32020 , \2172 );
nand \U$31662 ( \32039 , \32037 , \32038 );
and \U$31663 ( \32040 , \32029 , \32039 );
and \U$31664 ( \32041 , \32023 , \32028 );
or \U$31665 ( \32042 , \32040 , \32041 );
xor \U$31666 ( \32043 , \32022 , \32042 );
not \U$31667 ( \32044 , \3629 );
not \U$31668 ( \32045 , RIc2266b0_33);
not \U$31669 ( \32046 , \9250 );
or \U$31670 ( \32047 , \32045 , \32046 );
nand \U$31671 ( \32048 , \9256 , \6890 );
nand \U$31672 ( \32049 , \32047 , \32048 );
not \U$31673 ( \32050 , \32049 );
or \U$31674 ( \32051 , \32044 , \32050 );
nand \U$31675 ( \32052 , \31628 , \3631 );
nand \U$31676 ( \32053 , \32051 , \32052 );
xor \U$31677 ( \32054 , \32043 , \32053 );
xor \U$31678 ( \32055 , \32023 , \32028 );
xor \U$31679 ( \32056 , \32055 , \32039 );
not \U$31680 ( \32057 , \3629 );
not \U$31681 ( \32058 , RIc2266b0_33);
not \U$31682 ( \32059 , \21156 );
or \U$31683 ( \32060 , \32058 , \32059 );
nand \U$31684 ( \32061 , \9275 , \16360 );
nand \U$31685 ( \32062 , \32060 , \32061 );
not \U$31686 ( \32063 , \32062 );
or \U$31687 ( \32064 , \32057 , \32063 );
nand \U$31688 ( \32065 , \32049 , \3631 );
nand \U$31689 ( \32066 , \32064 , \32065 );
xor \U$31690 ( \32067 , \32056 , \32066 );
not \U$31691 ( \32068 , \5519 );
not \U$31692 ( \32069 , \31990 );
or \U$31693 ( \32070 , \32068 , \32069 );
not \U$31694 ( \32071 , RIc2264d0_37);
not \U$31695 ( \32072 , \13465 );
or \U$31696 ( \32073 , \32071 , \32072 );
not \U$31697 ( \32074 , \9046 );
nand \U$31698 ( \32075 , \32074 , \5504 );
nand \U$31699 ( \32076 , \32073 , \32075 );
nand \U$31700 ( \32077 , \32076 , \5509 );
nand \U$31701 ( \32078 , \32070 , \32077 );
and \U$31702 ( \32079 , \32067 , \32078 );
and \U$31703 ( \32080 , \32056 , \32066 );
or \U$31704 ( \32081 , \32079 , \32080 );
xor \U$31705 ( \32082 , \32054 , \32081 );
not \U$31706 ( \32083 , \15164 );
and \U$31707 ( \32084 , RIc225a80_59, \2645 );
not \U$31708 ( \32085 , RIc225a80_59);
and \U$31709 ( \32086 , \32085 , \4240 );
or \U$31710 ( \32087 , \32084 , \32086 );
not \U$31711 ( \32088 , \32087 );
or \U$31712 ( \32089 , \32083 , \32088 );
nand \U$31713 ( \32090 , \31578 , \12670 );
nand \U$31714 ( \32091 , \32089 , \32090 );
and \U$31715 ( \32092 , \32082 , \32091 );
and \U$31716 ( \32093 , \32054 , \32081 );
or \U$31717 ( \32094 , \32092 , \32093 );
xor \U$31718 ( \32095 , \32012 , \32094 );
xor \U$31719 ( \32096 , \31555 , \31572 );
xor \U$31720 ( \32097 , \32096 , \31586 );
and \U$31721 ( \32098 , \32095 , \32097 );
and \U$31722 ( \32099 , \32012 , \32094 );
or \U$31723 ( \32100 , \32098 , \32099 );
and \U$31724 ( \32101 , \32010 , \32100 );
and \U$31725 ( \32102 , \31957 , \32009 );
or \U$31726 ( \32103 , \32101 , \32102 );
xor \U$31727 ( \32104 , \31955 , \32103 );
xor \U$31728 ( \32105 , \31394 , \31500 );
xor \U$31729 ( \32106 , \32105 , \31592 );
and \U$31730 ( \32107 , \32104 , \32106 );
and \U$31731 ( \32108 , \31955 , \32103 );
or \U$31732 ( \32109 , \32107 , \32108 );
xor \U$31733 ( \32110 , \31792 , \32109 );
xor \U$31734 ( \32111 , \30986 , \30996 );
xor \U$31735 ( \32112 , \32111 , \31007 );
and \U$31736 ( \32113 , \30906 , \9444 );
and \U$31737 ( \32114 , \31326 , \9459 );
nor \U$31738 ( \32115 , \32113 , \32114 );
not \U$31739 ( \32116 , \32115 );
not \U$31740 ( \32117 , \32116 );
and \U$31741 ( \32118 , \31056 , \12670 );
and \U$31742 ( \32119 , \31584 , \15164 );
nor \U$31743 ( \32120 , \32118 , \32119 );
not \U$31744 ( \32121 , \32120 );
not \U$31745 ( \32122 , \32121 );
or \U$31746 ( \32123 , \32117 , \32122 );
not \U$31747 ( \32124 , \32120 );
not \U$31748 ( \32125 , \32115 );
or \U$31749 ( \32126 , \32124 , \32125 );
xor \U$31750 ( \32127 , \30821 , \30847 );
xor \U$31751 ( \32128 , \32127 , \30858 );
nand \U$31752 ( \32129 , \32126 , \32128 );
nand \U$31753 ( \32130 , \32123 , \32129 );
xor \U$31754 ( \32131 , \32112 , \32130 );
xor \U$31755 ( \32132 , \31044 , \31031 );
xor \U$31756 ( \32133 , \32132 , \31020 );
xor \U$31757 ( \32134 , \32131 , \32133 );
xor \U$31758 ( \32135 , \32128 , \32116 );
xnor \U$31759 ( \32136 , \32135 , \32121 );
not \U$31760 ( \32137 , \32136 );
not \U$31761 ( \32138 , \32137 );
xor \U$31762 ( \32139 , \31742 , \31747 );
xor \U$31763 ( \32140 , \32139 , \31753 );
not \U$31764 ( \32141 , \32140 );
or \U$31765 ( \32142 , \32138 , \32141 );
or \U$31766 ( \32143 , \32140 , \32137 );
not \U$31767 ( \32144 , \9142 );
not \U$31768 ( \32145 , \31222 );
or \U$31769 ( \32146 , \32144 , \32145 );
nand \U$31770 ( \32147 , \31898 , \2078 );
nand \U$31771 ( \32148 , \32146 , \32147 );
not \U$31772 ( \32149 , \2697 );
not \U$31773 ( \32150 , RIc2267a0_31);
not \U$31774 ( \32151 , \10263 );
or \U$31775 ( \32152 , \32150 , \32151 );
nand \U$31776 ( \32153 , \10266 , \3648 );
nand \U$31777 ( \32154 , \32152 , \32153 );
not \U$31778 ( \32155 , \32154 );
or \U$31779 ( \32156 , \32149 , \32155 );
nand \U$31780 ( \32157 , \31615 , \2710 );
nand \U$31781 ( \32158 , \32156 , \32157 );
xor \U$31782 ( \32159 , \32148 , \32158 );
not \U$31783 ( \32160 , \5135 );
not \U$31784 ( \32161 , \31239 );
or \U$31785 ( \32162 , \32160 , \32161 );
not \U$31786 ( \32163 , RIc2265c0_35);
not \U$31787 ( \32164 , \9073 );
or \U$31788 ( \32165 , \32163 , \32164 );
nand \U$31789 ( \32166 , \10653 , \3620 );
nand \U$31790 ( \32167 , \32165 , \32166 );
nand \U$31791 ( \32168 , \32167 , \4381 );
nand \U$31792 ( \32169 , \32162 , \32168 );
and \U$31793 ( \32170 , \32159 , \32169 );
and \U$31794 ( \32171 , \32148 , \32158 );
or \U$31795 ( \32172 , \32170 , \32171 );
xor \U$31796 ( \32173 , \32022 , \32042 );
and \U$31797 ( \32174 , \32173 , \32053 );
and \U$31798 ( \32175 , \32022 , \32042 );
or \U$31799 ( \32176 , \32174 , \32175 );
xor \U$31800 ( \32177 , \32172 , \32176 );
xor \U$31801 ( \32178 , \31274 , \31285 );
xor \U$31802 ( \32179 , \32178 , \31301 );
not \U$31803 ( \32180 , \9129 );
not \U$31804 ( \32181 , \31642 );
or \U$31805 ( \32182 , \32180 , \32181 );
not \U$31806 ( \32183 , RIc226200_43);
not \U$31807 ( \32184 , \10322 );
or \U$31808 ( \32185 , \32183 , \32184 );
nand \U$31809 ( \32186 , \12727 , \9117 );
nand \U$31810 ( \32187 , \32185 , \32186 );
nand \U$31811 ( \32188 , \32187 , \9110 );
nand \U$31812 ( \32189 , \32182 , \32188 );
xor \U$31813 ( \32190 , \32179 , \32189 );
not \U$31814 ( \32191 , \9459 );
not \U$31815 ( \32192 , RIc225e40_51);
not \U$31816 ( \32193 , \9842 );
or \U$31817 ( \32194 , \32192 , \32193 );
nand \U$31818 ( \32195 , \4407 , \22140 );
nand \U$31819 ( \32196 , \32194 , \32195 );
not \U$31820 ( \32197 , \32196 );
or \U$31821 ( \32198 , \32191 , \32197 );
nand \U$31822 ( \32199 , \31333 , \9444 );
nand \U$31823 ( \32200 , \32198 , \32199 );
and \U$31824 ( \32201 , \32190 , \32200 );
and \U$31825 ( \32202 , \32179 , \32189 );
or \U$31826 ( \32203 , \32201 , \32202 );
and \U$31827 ( \32204 , \32177 , \32203 );
and \U$31828 ( \32205 , \32172 , \32176 );
or \U$31829 ( \32206 , \32204 , \32205 );
nand \U$31830 ( \32207 , \32143 , \32206 );
nand \U$31831 ( \32208 , \32142 , \32207 );
xor \U$31832 ( \32209 , \32134 , \32208 );
xor \U$31833 ( \32210 , \31606 , \31600 );
xor \U$31834 ( \32211 , \32210 , \31674 );
xor \U$31835 ( \32212 , \32209 , \32211 );
xor \U$31836 ( \32213 , \31768 , \31782 );
xor \U$31837 ( \32214 , \32213 , \31785 );
or \U$31838 ( \32215 , \32212 , \32214 );
xor \U$31839 ( \32216 , \31506 , \31544 );
xor \U$31840 ( \32217 , \32216 , \31589 );
not \U$31841 ( \32218 , \31780 );
and \U$31842 ( \32219 , \31777 , \31770 );
not \U$31843 ( \32220 , \31777 );
and \U$31844 ( \32221 , \32220 , \31779 );
nor \U$31845 ( \32222 , \32219 , \32221 );
not \U$31846 ( \32223 , \32222 );
or \U$31847 ( \32224 , \32218 , \32223 );
or \U$31848 ( \32225 , \32222 , \31780 );
nand \U$31849 ( \32226 , \32224 , \32225 );
xor \U$31850 ( \32227 , \32217 , \32226 );
xor \U$31851 ( \32228 , \32136 , \32140 );
xnor \U$31852 ( \32229 , \32228 , \32206 );
and \U$31853 ( \32230 , \32227 , \32229 );
and \U$31854 ( \32231 , \32217 , \32226 );
or \U$31855 ( \32232 , \32230 , \32231 );
nand \U$31856 ( \32233 , \32215 , \32232 );
nand \U$31857 ( \32234 , \32212 , \32214 );
nand \U$31858 ( \32235 , \32233 , \32234 );
and \U$31859 ( \32236 , \32110 , \32235 );
and \U$31860 ( \32237 , \31792 , \32109 );
or \U$31861 ( \32238 , \32236 , \32237 );
xor \U$31862 ( \32239 , \31764 , \32238 );
xor \U$31863 ( \32240 , \31766 , \31788 );
and \U$31864 ( \32241 , \32240 , \31791 );
and \U$31865 ( \32242 , \31766 , \31788 );
or \U$31866 ( \32243 , \32241 , \32242 );
xor \U$31867 ( \32244 , \30593 , \30725 );
xor \U$31868 ( \32245 , \32244 , \30743 );
xor \U$31869 ( \32246 , \32112 , \32130 );
and \U$31870 ( \32247 , \32246 , \32133 );
and \U$31871 ( \32248 , \32112 , \32130 );
or \U$31872 ( \32249 , \32247 , \32248 );
not \U$31873 ( \32250 , \32249 );
xor \U$31874 ( \32251 , \31010 , \31046 );
xor \U$31875 ( \32252 , \32251 , \31077 );
not \U$31876 ( \32253 , \32252 );
or \U$31877 ( \32254 , \32250 , \32253 );
or \U$31878 ( \32255 , \32252 , \32249 );
xor \U$31879 ( \32256 , \30728 , \30737 );
xor \U$31880 ( \32257 , \32256 , \30740 );
nand \U$31881 ( \32258 , \32255 , \32257 );
nand \U$31882 ( \32259 , \32254 , \32258 );
xor \U$31883 ( \32260 , \32245 , \32259 );
xor \U$31884 ( \32261 , \30973 , \30975 );
xor \U$31885 ( \32262 , \32261 , \31080 );
xor \U$31886 ( \32263 , \32260 , \32262 );
xor \U$31887 ( \32264 , \32243 , \32263 );
xor \U$31888 ( \32265 , \32257 , \32252 );
xnor \U$31889 ( \32266 , \32265 , \32249 );
not \U$31890 ( \32267 , \32266 );
not \U$31891 ( \32268 , \32267 );
xor \U$31892 ( \32269 , \31677 , \31597 );
xnor \U$31893 ( \32270 , \32269 , \31594 );
not \U$31894 ( \32271 , \32270 );
or \U$31895 ( \32272 , \32268 , \32271 );
or \U$31896 ( \32273 , \32270 , \32267 );
xor \U$31897 ( \32274 , \32134 , \32208 );
and \U$31898 ( \32275 , \32274 , \32211 );
and \U$31899 ( \32276 , \32134 , \32208 );
or \U$31900 ( \32277 , \32275 , \32276 );
nand \U$31901 ( \32278 , \32273 , \32277 );
nand \U$31902 ( \32279 , \32272 , \32278 );
xor \U$31903 ( \32280 , \32264 , \32279 );
and \U$31904 ( \32281 , \32239 , \32280 );
and \U$31905 ( \32282 , \31764 , \32238 );
or \U$31906 ( \32283 , \32281 , \32282 );
not \U$31907 ( \32284 , \32283 );
xor \U$31908 ( \32285 , \31113 , \31138 );
xnor \U$31909 ( \32286 , \32285 , \31109 );
xor \U$31910 ( \32287 , \31720 , \31722 );
and \U$31911 ( \32288 , \32287 , \31762 );
and \U$31912 ( \32289 , \31720 , \31722 );
or \U$31913 ( \32290 , \32288 , \32289 );
xor \U$31914 ( \32291 , \32286 , \32290 );
xor \U$31915 ( \32292 , \32245 , \32259 );
and \U$31916 ( \32293 , \32292 , \32262 );
and \U$31917 ( \32294 , \32245 , \32259 );
or \U$31918 ( \32295 , \32293 , \32294 );
xor \U$31919 ( \32296 , \32291 , \32295 );
xor \U$31920 ( \32297 , \32243 , \32263 );
and \U$31921 ( \32298 , \32297 , \32279 );
and \U$31922 ( \32299 , \32243 , \32263 );
or \U$31923 ( \32300 , \32298 , \32299 );
xor \U$31924 ( \32301 , \32296 , \32300 );
xor \U$31925 ( \32302 , \30554 , \30746 );
xor \U$31926 ( \32303 , \32302 , \30755 );
xor \U$31927 ( \32304 , \30936 , \31083 );
buf \U$31928 ( \32305 , \30968 );
xor \U$31929 ( \32306 , \32304 , \32305 );
xor \U$31930 ( \32307 , \32303 , \32306 );
xor \U$31931 ( \32308 , \31217 , \31683 );
and \U$31932 ( \32309 , \32308 , \31763 );
and \U$31933 ( \32310 , \31217 , \31683 );
or \U$31934 ( \32311 , \32309 , \32310 );
xor \U$31935 ( \32312 , \32307 , \32311 );
xor \U$31936 ( \32313 , \32301 , \32312 );
not \U$31937 ( \32314 , \32313 );
or \U$31938 ( \32315 , \32284 , \32314 );
xor \U$31939 ( \32316 , \31764 , \32238 );
xor \U$31940 ( \32317 , \32316 , \32280 );
xor \U$31941 ( \32318 , \31792 , \32109 );
xor \U$31942 ( \32319 , \32318 , \32235 );
not \U$31943 ( \32320 , \32319 );
and \U$31944 ( \32321 , \32277 , \32266 );
not \U$31945 ( \32322 , \32277 );
and \U$31946 ( \32323 , \32322 , \32267 );
nor \U$31947 ( \32324 , \32321 , \32323 );
not \U$31948 ( \32325 , \32324 );
not \U$31949 ( \32326 , \32270 );
or \U$31950 ( \32327 , \32325 , \32326 );
not \U$31951 ( \32328 , \32324 );
not \U$31952 ( \32329 , \32270 );
nand \U$31953 ( \32330 , \32328 , \32329 );
nand \U$31954 ( \32331 , \32327 , \32330 );
not \U$31955 ( \32332 , \32331 );
nand \U$31956 ( \32333 , \32320 , \32332 );
not \U$31957 ( \32334 , \32333 );
xor \U$31958 ( \32335 , \31955 , \32103 );
xor \U$31959 ( \32336 , \32335 , \32106 );
xor \U$31960 ( \32337 , \32148 , \32158 );
xor \U$31961 ( \32338 , \32337 , \32169 );
not \U$31962 ( \32339 , \32338 );
not \U$31963 ( \32340 , \9552 );
not \U$31964 ( \32341 , \31826 );
or \U$31965 ( \32342 , \32340 , \32341 );
not \U$31966 ( \32343 , RIc225f30_49);
not \U$31967 ( \32344 , \23773 );
or \U$31968 ( \32345 , \32343 , \32344 );
nand \U$31969 ( \32346 , \23776 , \11289 );
nand \U$31970 ( \32347 , \32345 , \32346 );
nand \U$31971 ( \32348 , \32347 , \10445 );
nand \U$31972 ( \32349 , \32342 , \32348 );
not \U$31973 ( \32350 , \4383 );
not \U$31974 ( \32351 , \32167 );
or \U$31975 ( \32352 , \32350 , \32351 );
not \U$31976 ( \32353 , RIc2265c0_35);
not \U$31977 ( \32354 , \10111 );
or \U$31978 ( \32355 , \32353 , \32354 );
nand \U$31979 ( \32356 , \10110 , \9587 );
nand \U$31980 ( \32357 , \32355 , \32356 );
nand \U$31981 ( \32358 , \32357 , \4381 );
nand \U$31982 ( \32359 , \32352 , \32358 );
not \U$31983 ( \32360 , \2710 );
not \U$31984 ( \32361 , \32154 );
or \U$31985 ( \32362 , \32360 , \32361 );
not \U$31986 ( \32363 , RIc2267a0_31);
not \U$31987 ( \32364 , \30574 );
or \U$31988 ( \32365 , \32363 , \32364 );
nand \U$31989 ( \32366 , \30573 , \2072 );
nand \U$31990 ( \32367 , \32365 , \32366 );
nand \U$31991 ( \32368 , \32367 , \2697 );
nand \U$31992 ( \32369 , \32362 , \32368 );
or \U$31993 ( \32370 , \32359 , \32369 );
and \U$31994 ( \32371 , \32349 , \32370 );
and \U$31995 ( \32372 , \32369 , \32359 );
nor \U$31996 ( \32373 , \32371 , \32372 );
nand \U$31997 ( \32374 , \32339 , \32373 );
not \U$31998 ( \32375 , \32374 );
xor \U$31999 ( \32376 , \31867 , \31880 );
not \U$32000 ( \32377 , \2172 );
not \U$32001 ( \32378 , \32035 );
or \U$32002 ( \32379 , \32377 , \32378 );
not \U$32003 ( \32380 , RIc226a70_25);
not \U$32004 ( \32381 , \15623 );
or \U$32005 ( \32382 , \32380 , \32381 );
nand \U$32006 ( \32383 , \20393 , \3982 );
nand \U$32007 ( \32384 , \32382 , \32383 );
nand \U$32008 ( \32385 , \32384 , \2194 );
nand \U$32009 ( \32386 , \32379 , \32385 );
xor \U$32010 ( \32387 , \32376 , \32386 );
not \U$32011 ( \32388 , \2154 );
not \U$32012 ( \32389 , \31889 );
or \U$32013 ( \32390 , \32388 , \32389 );
not \U$32014 ( \32391 , RIc226980_27);
not \U$32015 ( \32392 , \30815 );
or \U$32016 ( \32393 , \32391 , \32392 );
nand \U$32017 ( \32394 , \19721 , \2799 );
nand \U$32018 ( \32395 , \32393 , \32394 );
nand \U$32019 ( \32396 , \32395 , \2138 );
nand \U$32020 ( \32397 , \32390 , \32396 );
and \U$32021 ( \32398 , \32387 , \32397 );
and \U$32022 ( \32399 , \32376 , \32386 );
or \U$32023 ( \32400 , \32398 , \32399 );
not \U$32024 ( \32401 , \6688 );
not \U$32025 ( \32402 , RIc2263e0_39);
not \U$32026 ( \32403 , \8910 );
or \U$32027 ( \32404 , \32402 , \32403 );
nand \U$32028 ( \32405 , \17744 , \8990 );
nand \U$32029 ( \32406 , \32404 , \32405 );
not \U$32030 ( \32407 , \32406 );
or \U$32031 ( \32408 , \32401 , \32407 );
nand \U$32032 ( \32409 , \31859 , \6307 );
nand \U$32033 ( \32410 , \32408 , \32409 );
xor \U$32034 ( \32411 , \32400 , \32410 );
not \U$32035 ( \32412 , \9690 );
not \U$32036 ( \32413 , RIc2262f0_41);
not \U$32037 ( \32414 , \13370 );
or \U$32038 ( \32415 , \32413 , \32414 );
nand \U$32039 ( \32416 , \8952 , \9822 );
nand \U$32040 ( \32417 , \32415 , \32416 );
not \U$32041 ( \32418 , \32417 );
or \U$32042 ( \32419 , \32412 , \32418 );
not \U$32043 ( \32420 , \9817 );
nand \U$32044 ( \32421 , \32420 , \31846 );
nand \U$32045 ( \32422 , \32419 , \32421 );
and \U$32046 ( \32423 , \32411 , \32422 );
and \U$32047 ( \32424 , \32400 , \32410 );
or \U$32048 ( \32425 , \32423 , \32424 );
not \U$32049 ( \32426 , \32425 );
or \U$32050 ( \32427 , \32375 , \32426 );
not \U$32051 ( \32428 , \32373 );
nand \U$32052 ( \32429 , \32428 , \32338 );
nand \U$32053 ( \32430 , \32427 , \32429 );
xor \U$32054 ( \32431 , \32172 , \32176 );
xor \U$32055 ( \32432 , \32431 , \32203 );
xor \U$32056 ( \32433 , \32430 , \32432 );
xor \U$32057 ( \32434 , \31794 , \31796 );
xor \U$32058 ( \32435 , \32434 , \31831 );
and \U$32059 ( \32436 , \32433 , \32435 );
and \U$32060 ( \32437 , \32430 , \32432 );
or \U$32061 ( \32438 , \32436 , \32437 );
xor \U$32062 ( \32439 , \31834 , \31836 );
xor \U$32063 ( \32440 , \32439 , \31952 );
xor \U$32064 ( \32441 , \32438 , \32440 );
xor \U$32065 ( \32442 , \31957 , \32009 );
xor \U$32066 ( \32443 , \32442 , \32100 );
and \U$32067 ( \32444 , \32441 , \32443 );
and \U$32068 ( \32445 , \32438 , \32440 );
or \U$32069 ( \32446 , \32444 , \32445 );
or \U$32070 ( \32447 , \32336 , \32446 );
not \U$32071 ( \32448 , \9129 );
not \U$32072 ( \32449 , \32187 );
or \U$32073 ( \32450 , \32448 , \32449 );
not \U$32074 ( \32451 , RIc226200_43);
not \U$32075 ( \32452 , \8830 );
or \U$32076 ( \32453 , \32451 , \32452 );
nand \U$32077 ( \32454 , \20216 , \9106 );
nand \U$32078 ( \32455 , \32453 , \32454 );
nand \U$32079 ( \32456 , \32455 , \9110 );
nand \U$32080 ( \32457 , \32450 , \32456 );
not \U$32081 ( \32458 , \10953 );
not \U$32082 ( \32459 , \31815 );
or \U$32083 ( \32460 , \32458 , \32459 );
not \U$32084 ( \32461 , RIc226020_47);
not \U$32085 ( \32462 , \21438 );
or \U$32086 ( \32463 , \32461 , \32462 );
nand \U$32087 ( \32464 , \6720 , \11607 );
nand \U$32088 ( \32465 , \32463 , \32464 );
nand \U$32089 ( \32466 , \32465 , \9641 );
nand \U$32090 ( \32467 , \32460 , \32466 );
xor \U$32091 ( \32468 , \32457 , \32467 );
not \U$32092 ( \32469 , \9398 );
not \U$32093 ( \32470 , \31803 );
or \U$32094 ( \32471 , \32469 , \32470 );
not \U$32095 ( \32472 , RIc226110_45);
not \U$32096 ( \32473 , \16531 );
or \U$32097 ( \32474 , \32472 , \32473 );
nand \U$32098 ( \32475 , \8886 , \9379 );
nand \U$32099 ( \32476 , \32474 , \32475 );
nand \U$32100 ( \32477 , \32476 , \9934 );
nand \U$32101 ( \32478 , \32471 , \32477 );
and \U$32102 ( \32479 , \32468 , \32478 );
and \U$32103 ( \32480 , \32457 , \32467 );
or \U$32104 ( \32481 , \32479 , \32480 );
not \U$32105 ( \32482 , \32481 );
not \U$32106 ( \32483 , \32482 );
xor \U$32107 ( \32484 , \31817 , \31807 );
xnor \U$32108 ( \32485 , \32484 , \31828 );
not \U$32109 ( \32486 , \32485 );
or \U$32110 ( \32487 , \32483 , \32486 );
xor \U$32111 ( \32488 , \32179 , \32189 );
xor \U$32112 ( \32489 , \32488 , \32200 );
nand \U$32113 ( \32490 , \32487 , \32489 );
not \U$32114 ( \32491 , \32485 );
nand \U$32115 ( \32492 , \32491 , \32481 );
nand \U$32116 ( \32493 , \32490 , \32492 );
xor \U$32117 ( \32494 , \31850 , \31861 );
xor \U$32118 ( \32495 , \32494 , \31911 );
not \U$32119 ( \32496 , \9444 );
not \U$32120 ( \32497 , \32196 );
or \U$32121 ( \32498 , \32496 , \32497 );
not \U$32122 ( \32499 , RIc225e40_51);
not \U$32123 ( \32500 , \10230 );
or \U$32124 ( \32501 , \32499 , \32500 );
nand \U$32125 ( \32502 , \10231 , \22140 );
nand \U$32126 ( \32503 , \32501 , \32502 );
nand \U$32127 ( \32504 , \32503 , \9459 );
nand \U$32128 ( \32505 , \32498 , \32504 );
not \U$32129 ( \32506 , \12945 );
not \U$32130 ( \32507 , \31923 );
or \U$32131 ( \32508 , \32506 , \32507 );
not \U$32132 ( \32509 , RIc225d50_53);
not \U$32133 ( \32510 , \4414 );
or \U$32134 ( \32511 , \32509 , \32510 );
nand \U$32135 ( \32512 , \4418 , \11585 );
nand \U$32136 ( \32513 , \32511 , \32512 );
nand \U$32137 ( \32514 , \32513 , \9488 );
nand \U$32138 ( \32515 , \32508 , \32514 );
xor \U$32139 ( \32516 , \32505 , \32515 );
not \U$32140 ( \32517 , \11965 );
not \U$32141 ( \32518 , RIc225b70_57);
not \U$32142 ( \32519 , \15216 );
or \U$32143 ( \32520 , \32518 , \32519 );
nand \U$32144 ( \32521 , \10533 , \10074 );
nand \U$32145 ( \32522 , \32520 , \32521 );
not \U$32146 ( \32523 , \32522 );
or \U$32147 ( \32524 , \32517 , \32523 );
nand \U$32148 ( \32525 , \31965 , \11974 );
nand \U$32149 ( \32526 , \32524 , \32525 );
and \U$32150 ( \32527 , \32516 , \32526 );
and \U$32151 ( \32528 , \32505 , \32515 );
or \U$32152 ( \32529 , \32527 , \32528 );
xor \U$32153 ( \32530 , \32495 , \32529 );
xor \U$32154 ( \32531 , \31881 , \31891 );
xor \U$32155 ( \32532 , \32531 , \31908 );
not \U$32156 ( \32533 , \20862 );
not \U$32157 ( \32534 , \31974 );
or \U$32158 ( \32535 , \32533 , \32534 );
not \U$32159 ( \32536 , RIc225990_61);
not \U$32160 ( \32537 , \3810 );
or \U$32161 ( \32538 , \32536 , \32537 );
nand \U$32162 ( \32539 , \2720 , \10338 );
nand \U$32163 ( \32540 , \32538 , \32539 );
nand \U$32164 ( \32541 , \32540 , \15719 );
nand \U$32165 ( \32542 , \32535 , \32541 );
xor \U$32166 ( \32543 , \32532 , \32542 );
not \U$32167 ( \32544 , \13025 );
not \U$32168 ( \32545 , \31931 );
or \U$32169 ( \32546 , \32544 , \32545 );
not \U$32170 ( \32547 , RIc225c60_55);
not \U$32171 ( \32548 , \6439 );
or \U$32172 ( \32549 , \32547 , \32548 );
nand \U$32173 ( \32550 , \2981 , \11041 );
nand \U$32174 ( \32551 , \32549 , \32550 );
nand \U$32175 ( \32552 , \32551 , \11118 );
nand \U$32176 ( \32553 , \32546 , \32552 );
and \U$32177 ( \32554 , \32543 , \32553 );
and \U$32178 ( \32555 , \32532 , \32542 );
or \U$32179 ( \32556 , \32554 , \32555 );
and \U$32180 ( \32557 , \32530 , \32556 );
and \U$32181 ( \32558 , \32495 , \32529 );
or \U$32182 ( \32559 , \32557 , \32558 );
xor \U$32183 ( \32560 , \32493 , \32559 );
xor \U$32184 ( \32561 , \31925 , \31935 );
xor \U$32185 ( \32562 , \32561 , \31946 );
xnor \U$32186 ( \32563 , \31967 , \31992 );
not \U$32187 ( \32564 , \31978 );
and \U$32188 ( \32565 , \32563 , \32564 );
not \U$32189 ( \32566 , \32563 );
and \U$32190 ( \32567 , \32566 , \31978 );
nor \U$32191 ( \32568 , \32565 , \32567 );
or \U$32192 ( \32569 , \32562 , \32568 );
not \U$32193 ( \32570 , \2086 );
not \U$32194 ( \32571 , \31906 );
or \U$32195 ( \32572 , \32570 , \32571 );
and \U$32196 ( \32573 , RIc226890_29, \17625 );
not \U$32197 ( \32574 , RIc226890_29);
and \U$32198 ( \32575 , \32574 , \13497 );
or \U$32199 ( \32576 , \32573 , \32575 );
nand \U$32200 ( \32577 , \2078 , \32576 );
nand \U$32201 ( \32578 , \32572 , \32577 );
not \U$32202 ( \32579 , \1930 );
nor \U$32203 ( \32580 , \32579 , \18356 );
not \U$32204 ( \32581 , \2172 );
not \U$32205 ( \32582 , \32384 );
or \U$32206 ( \32583 , \32581 , \32582 );
not \U$32207 ( \32584 , RIc226a70_25);
not \U$32208 ( \32585 , \20528 );
or \U$32209 ( \32586 , \32584 , \32585 );
buf \U$32210 ( \32587 , \16259 );
not \U$32211 ( \32588 , \32587 );
nand \U$32212 ( \32589 , \32588 , \2190 );
nand \U$32213 ( \32590 , \32586 , \32589 );
nand \U$32214 ( \32591 , \32590 , \2194 );
nand \U$32215 ( \32592 , \32583 , \32591 );
xor \U$32216 ( \32593 , \32580 , \32592 );
not \U$32217 ( \32594 , \2138 );
not \U$32218 ( \32595 , RIc226980_27);
not \U$32219 ( \32596 , \15630 );
or \U$32220 ( \32597 , \32595 , \32596 );
nand \U$32221 ( \32598 , \15633 , \2799 );
nand \U$32222 ( \32599 , \32597 , \32598 );
not \U$32223 ( \32600 , \32599 );
or \U$32224 ( \32601 , \32594 , \32600 );
nand \U$32225 ( \32602 , \32395 , \2153 );
nand \U$32226 ( \32603 , \32601 , \32602 );
and \U$32227 ( \32604 , \32593 , \32603 );
and \U$32228 ( \32605 , \32580 , \32592 );
or \U$32229 ( \32606 , \32604 , \32605 );
xor \U$32230 ( \32607 , \32578 , \32606 );
not \U$32231 ( \32608 , \5509 );
not \U$32232 ( \32609 , RIc2264d0_37);
not \U$32233 ( \32610 , \10652 );
or \U$32234 ( \32611 , \32609 , \32610 );
not \U$32235 ( \32612 , \11478 );
nand \U$32236 ( \32613 , \32612 , \12522 );
nand \U$32237 ( \32614 , \32611 , \32613 );
not \U$32238 ( \32615 , \32614 );
or \U$32239 ( \32616 , \32608 , \32615 );
nand \U$32240 ( \32617 , \32076 , \5519 );
nand \U$32241 ( \32618 , \32616 , \32617 );
and \U$32242 ( \32619 , \32607 , \32618 );
and \U$32243 ( \32620 , \32578 , \32606 );
or \U$32244 ( \32621 , \32619 , \32620 );
not \U$32245 ( \32622 , \20159 );
not \U$32246 ( \32623 , RIc2258a0_63);
not \U$32247 ( \32624 , \5819 );
or \U$32248 ( \32625 , \32623 , \32624 );
nand \U$32249 ( \32626 , \2479 , \15620 );
nand \U$32250 ( \32627 , \32625 , \32626 );
not \U$32251 ( \32628 , \32627 );
or \U$32252 ( \32629 , \32622 , \32628 );
nand \U$32253 ( \32630 , \31944 , RIc225828_64);
nand \U$32254 ( \32631 , \32629 , \32630 );
xor \U$32255 ( \32632 , \32621 , \32631 );
not \U$32256 ( \32633 , \12670 );
not \U$32257 ( \32634 , \32087 );
or \U$32258 ( \32635 , \32633 , \32634 );
and \U$32259 ( \32636 , RIc225a80_59, \5527 );
not \U$32260 ( \32637 , RIc225a80_59);
and \U$32261 ( \32638 , \32637 , \2044 );
or \U$32262 ( \32639 , \32636 , \32638 );
nand \U$32263 ( \32640 , \32639 , \15164 );
nand \U$32264 ( \32641 , \32635 , \32640 );
and \U$32265 ( \32642 , \32632 , \32641 );
and \U$32266 ( \32643 , \32621 , \32631 );
or \U$32267 ( \32644 , \32642 , \32643 );
nand \U$32268 ( \32645 , \32569 , \32644 );
nand \U$32269 ( \32646 , \32562 , \32568 );
nand \U$32270 ( \32647 , \32645 , \32646 );
and \U$32271 ( \32648 , \32560 , \32647 );
and \U$32272 ( \32649 , \32493 , \32559 );
or \U$32273 ( \32650 , \32648 , \32649 );
xor \U$32274 ( \32651 , \31839 , \31914 );
xor \U$32275 ( \32652 , \32651 , \31949 );
and \U$32276 ( \32653 , \31994 , \32006 );
not \U$32277 ( \32654 , \31994 );
and \U$32278 ( \32655 , \32654 , \32007 );
or \U$32279 ( \32656 , \32653 , \32655 );
xor \U$32280 ( \32657 , \32656 , \31997 );
xor \U$32281 ( \32658 , \32652 , \32657 );
xor \U$32282 ( \32659 , \32054 , \32081 );
xor \U$32283 ( \32660 , \32659 , \32091 );
and \U$32284 ( \32661 , \32367 , \2710 );
not \U$32285 ( \32662 , RIc2267a0_31);
not \U$32286 ( \32663 , \12862 );
or \U$32287 ( \32664 , \32662 , \32663 );
nand \U$32288 ( \32665 , \10086 , \2072 );
nand \U$32289 ( \32666 , \32664 , \32665 );
and \U$32290 ( \32667 , \32666 , \2697 );
nor \U$32291 ( \32668 , \32661 , \32667 );
not \U$32292 ( \32669 , \32668 );
not \U$32293 ( \32670 , \3629 );
not \U$32294 ( \32671 , RIc2266b0_33);
not \U$32295 ( \32672 , \10263 );
or \U$32296 ( \32673 , \32671 , \32672 );
nand \U$32297 ( \32674 , \16998 , \2692 );
nand \U$32298 ( \32675 , \32673 , \32674 );
not \U$32299 ( \32676 , \32675 );
or \U$32300 ( \32677 , \32670 , \32676 );
nand \U$32301 ( \32678 , \32062 , \3631 );
nand \U$32302 ( \32679 , \32677 , \32678 );
not \U$32303 ( \32680 , \32679 );
not \U$32304 ( \32681 , \32680 );
or \U$32305 ( \32682 , \32669 , \32681 );
not \U$32306 ( \32683 , \4381 );
not \U$32307 ( \32684 , RIc2265c0_35);
not \U$32308 ( \32685 , \30875 );
or \U$32309 ( \32686 , \32684 , \32685 );
nand \U$32310 ( \32687 , \27239 , \3620 );
nand \U$32311 ( \32688 , \32686 , \32687 );
not \U$32312 ( \32689 , \32688 );
or \U$32313 ( \32690 , \32683 , \32689 );
nand \U$32314 ( \32691 , \32357 , \4383 );
nand \U$32315 ( \32692 , \32690 , \32691 );
nand \U$32316 ( \32693 , \32682 , \32692 );
not \U$32317 ( \32694 , \32668 );
nand \U$32318 ( \32695 , \32679 , \32694 );
nand \U$32319 ( \32696 , \32693 , \32695 );
xor \U$32320 ( \32697 , \32369 , \32359 );
xor \U$32321 ( \32698 , \32349 , \32697 );
xor \U$32322 ( \32699 , \32696 , \32698 );
xor \U$32323 ( \32700 , \32376 , \32386 );
xor \U$32324 ( \32701 , \32700 , \32397 );
not \U$32325 ( \32702 , \9641 );
and \U$32326 ( \32703 , \9731 , \9624 );
not \U$32327 ( \32704 , \9731 );
and \U$32328 ( \32705 , \32704 , RIc226020_47);
or \U$32329 ( \32706 , \32703 , \32705 );
not \U$32330 ( \32707 , \32706 );
or \U$32331 ( \32708 , \32702 , \32707 );
nand \U$32332 ( \32709 , \32465 , \10953 );
nand \U$32333 ( \32710 , \32708 , \32709 );
xor \U$32334 ( \32711 , \32701 , \32710 );
not \U$32335 ( \32712 , RIc225f30_49);
not \U$32336 ( \32713 , \6493 );
or \U$32337 ( \32714 , \32712 , \32713 );
nand \U$32338 ( \32715 , \27798 , \9549 );
nand \U$32339 ( \32716 , \32714 , \32715 );
not \U$32340 ( \32717 , \32716 );
or \U$32341 ( \32718 , \32717 , \9533 );
not \U$32342 ( \32719 , \32347 );
or \U$32343 ( \32720 , \32719 , \23415 );
nand \U$32344 ( \32721 , \32718 , \32720 );
and \U$32345 ( \32722 , \32711 , \32721 );
and \U$32346 ( \32723 , \32701 , \32710 );
or \U$32347 ( \32724 , \32722 , \32723 );
and \U$32348 ( \32725 , \32699 , \32724 );
and \U$32349 ( \32726 , \32696 , \32698 );
or \U$32350 ( \32727 , \32725 , \32726 );
xor \U$32351 ( \32728 , \32660 , \32727 );
xor \U$32352 ( \32729 , \32056 , \32066 );
xor \U$32353 ( \32730 , \32729 , \32078 );
not \U$32354 ( \32731 , \9110 );
not \U$32355 ( \32732 , RIc226200_43);
not \U$32356 ( \32733 , \8807 );
or \U$32357 ( \32734 , \32732 , \32733 );
nand \U$32358 ( \32735 , \10859 , \9106 );
nand \U$32359 ( \32736 , \32734 , \32735 );
not \U$32360 ( \32737 , \32736 );
or \U$32361 ( \32738 , \32731 , \32737 );
nand \U$32362 ( \32739 , \32455 , \9205 );
nand \U$32363 ( \32740 , \32738 , \32739 );
not \U$32364 ( \32741 , \32740 );
not \U$32365 ( \32742 , \9934 );
not \U$32366 ( \32743 , RIc226110_45);
not \U$32367 ( \32744 , \20674 );
or \U$32368 ( \32745 , \32743 , \32744 );
nand \U$32369 ( \32746 , \12727 , \9379 );
nand \U$32370 ( \32747 , \32745 , \32746 );
not \U$32371 ( \32748 , \32747 );
or \U$32372 ( \32749 , \32742 , \32748 );
nand \U$32373 ( \32750 , \32476 , \9398 );
nand \U$32374 ( \32751 , \32749 , \32750 );
not \U$32375 ( \32752 , \32751 );
or \U$32376 ( \32753 , \32741 , \32752 );
or \U$32377 ( \32754 , \32751 , \32740 );
not \U$32378 ( \32755 , \9816 );
not \U$32379 ( \32756 , \32417 );
or \U$32380 ( \32757 , \32755 , \32756 );
not \U$32381 ( \32758 , RIc2262f0_41);
not \U$32382 ( \32759 , \21866 );
or \U$32383 ( \32760 , \32758 , \32759 );
nand \U$32384 ( \32761 , \11095 , \6303 );
nand \U$32385 ( \32762 , \32760 , \32761 );
nand \U$32386 ( \32763 , \32762 , \9690 );
nand \U$32387 ( \32764 , \32757 , \32763 );
nand \U$32388 ( \32765 , \32754 , \32764 );
nand \U$32389 ( \32766 , \32753 , \32765 );
xor \U$32390 ( \32767 , \32730 , \32766 );
or \U$32391 ( \32768 , RIc2269f8_26, RIc226980_27);
nand \U$32392 ( \32769 , \32768 , \18367 );
and \U$32393 ( \32770 , RIc2269f8_26, RIc226980_27);
nor \U$32394 ( \32771 , \32770 , \1905 );
and \U$32395 ( \32772 , \32769 , \32771 );
not \U$32396 ( \32773 , \2172 );
not \U$32397 ( \32774 , \32590 );
or \U$32398 ( \32775 , \32773 , \32774 );
or \U$32399 ( \32776 , \16248 , \1905 );
or \U$32400 ( \32777 , \18356 , RIc226a70_25);
nand \U$32401 ( \32778 , \32776 , \32777 );
nand \U$32402 ( \32779 , \32778 , \2194 );
nand \U$32403 ( \32780 , \32775 , \32779 );
and \U$32404 ( \32781 , \32772 , \32780 );
not \U$32405 ( \32782 , \2078 );
and \U$32406 ( \32783 , RIc226890_29, \20693 );
not \U$32407 ( \32784 , RIc226890_29);
and \U$32408 ( \32785 , \32784 , \20694 );
or \U$32409 ( \32786 , \32783 , \32785 );
not \U$32410 ( \32787 , \32786 );
or \U$32411 ( \32788 , \32782 , \32787 );
nand \U$32412 ( \32789 , \32576 , \2086 );
nand \U$32413 ( \32790 , \32788 , \32789 );
xor \U$32414 ( \32791 , \32781 , \32790 );
not \U$32415 ( \32792 , \2710 );
not \U$32416 ( \32793 , \32666 );
or \U$32417 ( \32794 , \32792 , \32793 );
not \U$32418 ( \32795 , RIc2267a0_31);
not \U$32419 ( \32796 , \20702 );
or \U$32420 ( \32797 , \32795 , \32796 );
buf \U$32421 ( \32798 , \10370 );
nand \U$32422 ( \32799 , \32798 , \3648 );
nand \U$32423 ( \32800 , \32797 , \32799 );
nand \U$32424 ( \32801 , \32800 , \2697 );
nand \U$32425 ( \32802 , \32794 , \32801 );
and \U$32426 ( \32803 , \32791 , \32802 );
and \U$32427 ( \32804 , \32781 , \32790 );
or \U$32428 ( \32805 , \32803 , \32804 );
not \U$32429 ( \32806 , \6307 );
not \U$32430 ( \32807 , \32406 );
or \U$32431 ( \32808 , \32806 , \32807 );
not \U$32432 ( \32809 , RIc2263e0_39);
not \U$32433 ( \32810 , \9211 );
not \U$32434 ( \32811 , \32810 );
or \U$32435 ( \32812 , \32809 , \32811 );
not \U$32436 ( \32813 , \8925 );
nand \U$32437 ( \32814 , \32813 , \9573 );
nand \U$32438 ( \32815 , \32812 , \32814 );
nand \U$32439 ( \32816 , \32815 , \6688 );
nand \U$32440 ( \32817 , \32808 , \32816 );
xor \U$32441 ( \32818 , \32805 , \32817 );
not \U$32442 ( \32819 , \11577 );
not \U$32443 ( \32820 , \32513 );
or \U$32444 ( \32821 , \32819 , \32820 );
not \U$32445 ( \32822 , RIc225d50_53);
not \U$32446 ( \32823 , \6076 );
or \U$32447 ( \32824 , \32822 , \32823 );
nand \U$32448 ( \32825 , \4407 , \11585 );
nand \U$32449 ( \32826 , \32824 , \32825 );
nand \U$32450 ( \32827 , \32826 , \9488 );
nand \U$32451 ( \32828 , \32821 , \32827 );
and \U$32452 ( \32829 , \32818 , \32828 );
and \U$32453 ( \32830 , \32805 , \32817 );
or \U$32454 ( \32831 , \32829 , \32830 );
and \U$32455 ( \32832 , \32767 , \32831 );
and \U$32456 ( \32833 , \32730 , \32766 );
or \U$32457 ( \32834 , \32832 , \32833 );
and \U$32458 ( \32835 , \32728 , \32834 );
and \U$32459 ( \32836 , \32660 , \32727 );
or \U$32460 ( \32837 , \32835 , \32836 );
and \U$32461 ( \32838 , \32658 , \32837 );
and \U$32462 ( \32839 , \32652 , \32657 );
or \U$32463 ( \32840 , \32838 , \32839 );
or \U$32464 ( \32841 , \32650 , \32840 );
xor \U$32465 ( \32842 , \32217 , \32226 );
xor \U$32466 ( \32843 , \32842 , \32229 );
nand \U$32467 ( \32844 , \32841 , \32843 );
nand \U$32468 ( \32845 , \32650 , \32840 );
nand \U$32469 ( \32846 , \32844 , \32845 );
nand \U$32470 ( \32847 , \32447 , \32846 );
nand \U$32471 ( \32848 , \32336 , \32446 );
nand \U$32472 ( \32849 , \32847 , \32848 );
not \U$32473 ( \32850 , \32849 );
or \U$32474 ( \32851 , \32334 , \32850 );
nand \U$32475 ( \32852 , \32319 , \32331 );
nand \U$32476 ( \32853 , \32851 , \32852 );
nand \U$32477 ( \32854 , \32317 , \32853 );
nand \U$32478 ( \32855 , \32315 , \32854 );
not \U$32479 ( \32856 , \32313 );
not \U$32480 ( \32857 , \32283 );
nand \U$32481 ( \32858 , \32856 , \32857 );
nand \U$32482 ( \32859 , \32855 , \32858 );
xor \U$32483 ( \32860 , \32286 , \32290 );
and \U$32484 ( \32861 , \32860 , \32295 );
and \U$32485 ( \32862 , \32286 , \32290 );
or \U$32486 ( \32863 , \32861 , \32862 );
xor \U$32487 ( \32864 , \32303 , \32306 );
and \U$32488 ( \32865 , \32864 , \32311 );
and \U$32489 ( \32866 , \32303 , \32306 );
or \U$32490 ( \32867 , \32865 , \32866 );
xor \U$32491 ( \32868 , \32863 , \32867 );
not \U$32492 ( \32869 , \31178 );
not \U$32493 ( \32870 , \31171 );
not \U$32494 ( \32871 , \31174 );
and \U$32495 ( \32872 , \32870 , \32871 );
and \U$32496 ( \32873 , \31171 , \31174 );
nor \U$32497 ( \32874 , \32872 , \32873 );
not \U$32498 ( \32875 , \32874 );
or \U$32499 ( \32876 , \32869 , \32875 );
or \U$32500 ( \32877 , \32874 , \31178 );
nand \U$32501 ( \32878 , \32876 , \32877 );
xor \U$32502 ( \32879 , \32868 , \32878 );
not \U$32503 ( \32880 , \32879 );
xor \U$32504 ( \32881 , \32296 , \32300 );
and \U$32505 ( \32882 , \32881 , \32312 );
and \U$32506 ( \32883 , \32296 , \32300 );
or \U$32507 ( \32884 , \32882 , \32883 );
not \U$32508 ( \32885 , \32884 );
nand \U$32509 ( \32886 , \32880 , \32885 );
not \U$32510 ( \32887 , \32886 );
or \U$32511 ( \32888 , \32859 , \32887 );
xor \U$32512 ( \32889 , \31167 , \31182 );
xnor \U$32513 ( \32890 , \32889 , \31165 );
xor \U$32514 ( \32891 , \32863 , \32867 );
and \U$32515 ( \32892 , \32891 , \32878 );
and \U$32516 ( \32893 , \32863 , \32867 );
or \U$32517 ( \32894 , \32892 , \32893 );
nand \U$32518 ( \32895 , \32890 , \32894 );
nand \U$32519 ( \32896 , \32879 , \32884 );
and \U$32520 ( \32897 , \32895 , \32896 );
nand \U$32521 ( \32898 , \32888 , \32897 );
not \U$32522 ( \32899 , \32890 );
not \U$32523 ( \32900 , \32894 );
nand \U$32524 ( \32901 , \32899 , \32900 );
and \U$32525 ( \32902 , \32898 , \32901 );
nand \U$32526 ( \32903 , \31163 , \31185 );
and \U$32527 ( \32904 , \30139 , \30537 , \31193 , \32903 );
buf \U$32528 ( \32905 , \32904 );
nand \U$32529 ( \32906 , \32902 , \32905 );
and \U$32530 ( \32907 , \31207 , \32906 );
xor \U$32531 ( \32908 , \29225 , \29230 );
and \U$32532 ( \32909 , \32908 , \29236 );
and \U$32533 ( \32910 , \29225 , \29230 );
or \U$32534 ( \32911 , \32909 , \32910 );
not \U$32535 ( \32912 , \5135 );
not \U$32536 ( \32913 , \21892 );
or \U$32537 ( \32914 , \32912 , \32913 );
nand \U$32538 ( \32915 , \29245 , \5741 );
nand \U$32539 ( \32916 , \32914 , \32915 );
xor \U$32540 ( \32917 , \32911 , \32916 );
not \U$32541 ( \32918 , \15729 );
not \U$32542 ( \32919 , \22108 );
or \U$32543 ( \32920 , \32918 , \32919 );
nand \U$32544 ( \32921 , \28693 , \15719 );
nand \U$32545 ( \32922 , \32920 , \32921 );
and \U$32546 ( \32923 , \32917 , \32922 );
and \U$32547 ( \32924 , \32911 , \32916 );
or \U$32548 ( \32925 , \32923 , \32924 );
not \U$32549 ( \32926 , \2392 );
not \U$32550 ( \32927 , \28737 );
or \U$32551 ( \32928 , \32926 , \32927 );
nand \U$32552 ( \32929 , \21195 , \2367 );
nand \U$32553 ( \32930 , \32928 , \32929 );
not \U$32554 ( \32931 , \2534 );
not \U$32555 ( \32932 , \21133 );
or \U$32556 ( \32933 , \32931 , \32932 );
nand \U$32557 ( \32934 , \28838 , \2518 );
nand \U$32558 ( \32935 , \32933 , \32934 );
or \U$32559 ( \32936 , \32930 , \32935 );
xor \U$32560 ( \32937 , \21091 , \21108 );
xor \U$32561 ( \32938 , \32937 , \21124 );
nand \U$32562 ( \32939 , \32936 , \32938 );
nand \U$32563 ( \32940 , \32930 , \32935 );
nand \U$32564 ( \32941 , \32939 , \32940 );
not \U$32565 ( \32942 , RIc225828_64);
not \U$32566 ( \32943 , \21314 );
or \U$32567 ( \32944 , \32942 , \32943 );
not \U$32568 ( \32945 , RIc2258a0_63);
not \U$32569 ( \32946 , \1393 );
or \U$32570 ( \32947 , \32945 , \32946 );
not \U$32571 ( \32948 , \1392 );
nand \U$32572 ( \32949 , \32948 , \15620 );
nand \U$32573 ( \32950 , \32947 , \32949 );
nand \U$32574 ( \32951 , \32950 , \20159 );
nand \U$32575 ( \32952 , \32944 , \32951 );
xor \U$32576 ( \32953 , \32941 , \32952 );
not \U$32577 ( \32954 , \15164 );
and \U$32578 ( \32955 , RIc225a80_59, \4182 );
not \U$32579 ( \32956 , RIc225a80_59);
and \U$32580 ( \32957 , \32956 , \4183 );
or \U$32581 ( \32958 , \32955 , \32957 );
not \U$32582 ( \32959 , \32958 );
or \U$32583 ( \32960 , \32954 , \32959 );
nand \U$32584 ( \32961 , \21208 , \12670 );
nand \U$32585 ( \32962 , \32960 , \32961 );
xor \U$32586 ( \32963 , \32953 , \32962 );
xor \U$32587 ( \32964 , \32925 , \32963 );
and \U$32588 ( \32965 , \22057 , \22034 );
not \U$32589 ( \32966 , \22057 );
and \U$32590 ( \32967 , \32966 , \22033 );
nor \U$32591 ( \32968 , \32965 , \32967 );
buf \U$32592 ( \32969 , \22045 );
xor \U$32593 ( \32970 , \32968 , \32969 );
not \U$32594 ( \32971 , \32970 );
xor \U$32595 ( \32972 , \32964 , \32971 );
xor \U$32596 ( \32973 , \28840 , \28850 );
and \U$32597 ( \32974 , \32973 , \28861 );
and \U$32598 ( \32975 , \28840 , \28850 );
or \U$32599 ( \32976 , \32974 , \32975 );
xor \U$32600 ( \32977 , \28723 , \28728 );
and \U$32601 ( \32978 , \32977 , \28739 );
and \U$32602 ( \32979 , \28723 , \28728 );
or \U$32603 ( \32980 , \32978 , \32979 );
xor \U$32604 ( \32981 , \32976 , \32980 );
not \U$32605 ( \32982 , \29179 );
not \U$32606 ( \32983 , \29168 );
or \U$32607 ( \32984 , \32982 , \32983 );
or \U$32608 ( \32985 , \29168 , \29179 );
nand \U$32609 ( \32986 , \32985 , \29159 );
nand \U$32610 ( \32987 , \32984 , \32986 );
and \U$32611 ( \32988 , \32981 , \32987 );
and \U$32612 ( \32989 , \32976 , \32980 );
or \U$32613 ( \32990 , \32988 , \32989 );
not \U$32614 ( \32991 , \1945 );
not \U$32615 ( \32992 , \28857 );
or \U$32616 ( \32993 , \32991 , \32992 );
nand \U$32617 ( \32994 , \21152 , \1963 );
nand \U$32618 ( \32995 , \32993 , \32994 );
not \U$32619 ( \32996 , \1930 );
not \U$32620 ( \32997 , \21917 );
or \U$32621 ( \32998 , \32996 , \32997 );
nand \U$32622 ( \32999 , \28845 , \10214 );
nand \U$32623 ( \33000 , \32998 , \32999 );
xor \U$32624 ( \33001 , \32995 , \33000 );
not \U$32625 ( \33002 , \2710 );
not \U$32626 ( \33003 , \21989 );
or \U$32627 ( \33004 , \33002 , \33003 );
nand \U$32628 ( \33005 , \29175 , \2697 );
nand \U$32629 ( \33006 , \33004 , \33005 );
xor \U$32630 ( \33007 , \33001 , \33006 );
not \U$32631 ( \33008 , \29143 );
not \U$32632 ( \33009 , \29131 );
or \U$32633 ( \33010 , \33008 , \33009 );
nand \U$32634 ( \33011 , \33010 , \29122 );
not \U$32635 ( \33012 , \29131 );
nand \U$32636 ( \33013 , \33012 , \29142 );
nand \U$32637 ( \33014 , \33011 , \33013 );
xor \U$32638 ( \33015 , \33007 , \33014 );
xor \U$32639 ( \33016 , \29237 , \29247 );
and \U$32640 ( \33017 , \33016 , \29258 );
and \U$32641 ( \33018 , \29237 , \29247 );
or \U$32642 ( \33019 , \33017 , \33018 );
and \U$32643 ( \33020 , \33015 , \33019 );
and \U$32644 ( \33021 , \33007 , \33014 );
or \U$32645 ( \33022 , \33020 , \33021 );
xor \U$32646 ( \33023 , \32990 , \33022 );
xor \U$32647 ( \33024 , \32938 , \32935 );
xnor \U$32648 ( \33025 , \33024 , \32930 );
not \U$32649 ( \33026 , \33025 );
not \U$32650 ( \33027 , \33026 );
or \U$32651 ( \33028 , \29216 , \29195 );
nand \U$32652 ( \33029 , \33028 , \29205 );
nand \U$32653 ( \33030 , \29216 , \29195 );
nand \U$32654 ( \33031 , \33029 , \33030 );
not \U$32655 ( \33032 , \33031 );
or \U$32656 ( \33033 , \33027 , \33032 );
not \U$32657 ( \33034 , \33025 );
not \U$32658 ( \33035 , \33031 );
not \U$32659 ( \33036 , \33035 );
or \U$32660 ( \33037 , \33034 , \33036 );
xor \U$32661 ( \33038 , \28685 , \28695 );
and \U$32662 ( \33039 , \33038 , \28713 );
and \U$32663 ( \33040 , \28685 , \28695 );
or \U$32664 ( \33041 , \33039 , \33040 );
nand \U$32665 ( \33042 , \33037 , \33041 );
nand \U$32666 ( \33043 , \33033 , \33042 );
xor \U$32667 ( \33044 , \33023 , \33043 );
xor \U$32668 ( \33045 , \32972 , \33044 );
xor \U$32669 ( \33046 , \33007 , \33014 );
xor \U$32670 ( \33047 , \33046 , \33019 );
xor \U$32671 ( \33048 , \29259 , \29267 );
and \U$32672 ( \33049 , \33048 , \29274 );
and \U$32673 ( \33050 , \29259 , \29267 );
or \U$32674 ( \33051 , \33049 , \33050 );
xor \U$32675 ( \33052 , \33047 , \33051 );
xor \U$32676 ( \33053 , \29075 , \29079 );
and \U$32677 ( \33054 , \33053 , \29086 );
and \U$32678 ( \33055 , \29075 , \29079 );
or \U$32679 ( \33056 , \33054 , \33055 );
and \U$32680 ( \33057 , \33052 , \33056 );
and \U$32681 ( \33058 , \33047 , \33051 );
or \U$32682 ( \33059 , \33057 , \33058 );
xor \U$32683 ( \33060 , \33045 , \33059 );
xor \U$32684 ( \33061 , \33047 , \33051 );
xor \U$32685 ( \33062 , \33061 , \33056 );
not \U$32686 ( \33063 , \29222 );
not \U$32687 ( \33064 , \29218 );
or \U$32688 ( \33065 , \33063 , \33064 );
or \U$32689 ( \33066 , \29222 , \29218 );
nand \U$32690 ( \33067 , \33066 , \29275 );
nand \U$32691 ( \33068 , \33065 , \33067 );
xor \U$32692 ( \33069 , \33062 , \33068 );
not \U$32693 ( \33070 , \28635 );
nand \U$32694 ( \33071 , \33070 , \28658 );
and \U$32695 ( \33072 , \33071 , \28714 );
nor \U$32696 ( \33073 , \33070 , \28658 );
nor \U$32697 ( \33074 , \33072 , \33073 );
not \U$32698 ( \33075 , \33074 );
not \U$32699 ( \33076 , \33075 );
nand \U$32700 ( \33077 , \29180 , \29148 );
not \U$32701 ( \33078 , \33077 );
not \U$32702 ( \33079 , \29217 );
or \U$32703 ( \33080 , \33078 , \33079 );
not \U$32704 ( \33081 , \29148 );
nand \U$32705 ( \33082 , \33081 , \29181 );
nand \U$32706 ( \33083 , \33080 , \33082 );
not \U$32707 ( \33084 , \33083 );
not \U$32708 ( \33085 , \33084 );
or \U$32709 ( \33086 , \33076 , \33085 );
nand \U$32710 ( \33087 , \33083 , \33074 );
nand \U$32711 ( \33088 , \33086 , \33087 );
not \U$32712 ( \33089 , \9142 );
not \U$32713 ( \33090 , \21999 );
or \U$32714 ( \33091 , \33089 , \33090 );
nand \U$32715 ( \33092 , \29166 , \2784 );
nand \U$32716 ( \33093 , \33091 , \33092 );
not \U$32717 ( \33094 , \2138 );
not \U$32718 ( \33095 , \29155 );
or \U$32719 ( \33096 , \33094 , \33095 );
nand \U$32720 ( \33097 , \21907 , \2154 );
nand \U$32721 ( \33098 , \33096 , \33097 );
xor \U$32722 ( \33099 , \33093 , \33098 );
not \U$32723 ( \33100 , \2173 );
not \U$32724 ( \33101 , \21869 );
or \U$32725 ( \33102 , \33100 , \33101 );
nand \U$32726 ( \33103 , \29128 , \2195 );
nand \U$32727 ( \33104 , \33102 , \33103 );
xor \U$32728 ( \33105 , \33099 , \33104 );
not \U$32729 ( \33106 , \28784 );
not \U$32730 ( \33107 , \28808 );
or \U$32731 ( \33108 , \33106 , \33107 );
nand \U$32732 ( \33109 , \33108 , \28791 );
nand \U$32733 ( \33110 , \28807 , \28785 );
nand \U$32734 ( \33111 , \33109 , \33110 );
xor \U$32735 ( \33112 , \33105 , \33111 );
xor \U$32736 ( \33113 , \21959 , \21968 );
xor \U$32737 ( \33114 , \33113 , \21980 );
not \U$32738 ( \33115 , \16891 );
not \U$32739 ( \33116 , \28759 );
or \U$32740 ( \33117 , \33115 , \33116 );
nand \U$32741 ( \33118 , \32950 , RIc225828_64);
nand \U$32742 ( \33119 , \33117 , \33118 );
xor \U$32743 ( \33120 , \33114 , \33119 );
not \U$32744 ( \33121 , \9444 );
not \U$32745 ( \33122 , \22142 );
or \U$32746 ( \33123 , \33121 , \33122 );
nand \U$32747 ( \33124 , \28604 , \9459 );
nand \U$32748 ( \33125 , \33123 , \33124 );
xor \U$32749 ( \33126 , \33120 , \33125 );
xor \U$32750 ( \33127 , \33112 , \33126 );
and \U$32751 ( \33128 , \33088 , \33127 );
not \U$32752 ( \33129 , \33088 );
not \U$32753 ( \33130 , \33127 );
and \U$32754 ( \33131 , \33129 , \33130 );
nor \U$32755 ( \33132 , \33128 , \33131 );
and \U$32756 ( \33133 , \33069 , \33132 );
and \U$32757 ( \33134 , \33062 , \33068 );
or \U$32758 ( \33135 , \33133 , \33134 );
xor \U$32759 ( \33136 , \33060 , \33135 );
not \U$32760 ( \33137 , \33075 );
not \U$32761 ( \33138 , \33083 );
or \U$32762 ( \33139 , \33137 , \33138 );
not \U$32763 ( \33140 , \33074 );
not \U$32764 ( \33141 , \33084 );
or \U$32765 ( \33142 , \33140 , \33141 );
nand \U$32766 ( \33143 , \33142 , \33127 );
nand \U$32767 ( \33144 , \33139 , \33143 );
xor \U$32768 ( \33145 , \21090 , \21127 );
xor \U$32769 ( \33146 , \33145 , \21142 );
xor \U$32770 ( \33147 , \32995 , \33000 );
and \U$32771 ( \33148 , \33147 , \33006 );
and \U$32772 ( \33149 , \32995 , \33000 );
or \U$32773 ( \33150 , \33148 , \33149 );
xor \U$32774 ( \33151 , \33146 , \33150 );
xor \U$32775 ( \33152 , \33093 , \33098 );
and \U$32776 ( \33153 , \33152 , \33104 );
and \U$32777 ( \33154 , \33093 , \33098 );
or \U$32778 ( \33155 , \33153 , \33154 );
xor \U$32779 ( \33156 , \33151 , \33155 );
xor \U$32780 ( \33157 , \21162 , \21179 );
xor \U$32781 ( \33158 , \33157 , \21197 );
not \U$32782 ( \33159 , \5519 );
not \U$32783 ( \33160 , \21934 );
or \U$32784 ( \33161 , \33159 , \33160 );
nand \U$32785 ( \33162 , \29256 , \5509 );
nand \U$32786 ( \33163 , \33161 , \33162 );
not \U$32787 ( \33164 , \33163 );
not \U$32788 ( \33165 , \3629 );
not \U$32789 ( \33166 , \29140 );
or \U$32790 ( \33167 , \33165 , \33166 );
nand \U$32791 ( \33168 , \21882 , \3631 );
nand \U$32792 ( \33169 , \33167 , \33168 );
not \U$32793 ( \33170 , \33169 );
or \U$32794 ( \33171 , \33164 , \33170 );
not \U$32795 ( \33172 , \33169 );
not \U$32796 ( \33173 , \33172 );
not \U$32797 ( \33174 , \33163 );
not \U$32798 ( \33175 , \33174 );
or \U$32799 ( \33176 , \33173 , \33175 );
not \U$32800 ( \33177 , \6307 );
not \U$32801 ( \33178 , \22133 );
or \U$32802 ( \33179 , \33177 , \33178 );
nand \U$32803 ( \33180 , \29120 , \6688 );
nand \U$32804 ( \33181 , \33179 , \33180 );
nand \U$32805 ( \33182 , \33176 , \33181 );
nand \U$32806 ( \33183 , \33171 , \33182 );
xor \U$32807 ( \33184 , \33158 , \33183 );
not \U$32808 ( \33185 , \21920 );
not \U$32809 ( \33186 , \21924 );
or \U$32810 ( \33187 , \33185 , \33186 );
nand \U$32811 ( \33188 , \21911 , \21919 );
nand \U$32812 ( \33189 , \33187 , \33188 );
xor \U$32813 ( \33190 , \33189 , \21936 );
xor \U$32814 ( \33191 , \33184 , \33190 );
xor \U$32815 ( \33192 , \33156 , \33191 );
not \U$32816 ( \33193 , \33181 );
not \U$32817 ( \33194 , \33172 );
or \U$32818 ( \33195 , \33193 , \33194 );
or \U$32819 ( \33196 , \33181 , \33172 );
nand \U$32820 ( \33197 , \33195 , \33196 );
not \U$32821 ( \33198 , \33197 );
not \U$32822 ( \33199 , \33174 );
and \U$32823 ( \33200 , \33198 , \33199 );
and \U$32824 ( \33201 , \33197 , \33174 );
nor \U$32825 ( \33202 , \33200 , \33201 );
or \U$32826 ( \33203 , \28606 , \28619 );
nand \U$32827 ( \33204 , \33203 , \28634 );
nand \U$32828 ( \33205 , \28606 , \28619 );
nand \U$32829 ( \33206 , \33204 , \33205 );
not \U$32830 ( \33207 , \33206 );
and \U$32831 ( \33208 , \33202 , \33207 );
xor \U$32832 ( \33209 , \32911 , \32916 );
xor \U$32833 ( \33210 , \33209 , \32922 );
not \U$32834 ( \33211 , \33210 );
or \U$32835 ( \33212 , \33208 , \33211 );
not \U$32836 ( \33213 , \33202 );
nand \U$32837 ( \33214 , \33213 , \33206 );
nand \U$32838 ( \33215 , \33212 , \33214 );
xor \U$32839 ( \33216 , \33192 , \33215 );
xor \U$32840 ( \33217 , \33144 , \33216 );
not \U$32841 ( \33218 , \33105 );
not \U$32842 ( \33219 , \33111 );
or \U$32843 ( \33220 , \33218 , \33219 );
or \U$32844 ( \33221 , \33111 , \33105 );
nand \U$32845 ( \33222 , \33221 , \33126 );
nand \U$32846 ( \33223 , \33220 , \33222 );
xor \U$32847 ( \33224 , \28740 , \28744 );
and \U$32848 ( \33225 , \33224 , \28761 );
and \U$32849 ( \33226 , \28740 , \28744 );
or \U$32850 ( \33227 , \33225 , \33226 );
not \U$32851 ( \33228 , \9552 );
not \U$32852 ( \33229 , \22099 );
or \U$32853 ( \33230 , \33228 , \33229 );
nand \U$32854 ( \33231 , \28711 , \10445 );
nand \U$32855 ( \33232 , \33230 , \33231 );
not \U$32856 ( \33233 , \9641 );
not \U$32857 ( \33234 , \29201 );
or \U$32858 ( \33235 , \33233 , \33234 );
nand \U$32859 ( \33236 , \22055 , \12304 );
nand \U$32860 ( \33237 , \33235 , \33236 );
xor \U$32861 ( \33238 , \33232 , \33237 );
not \U$32862 ( \33239 , \11965 );
not \U$32863 ( \33240 , \29214 );
or \U$32864 ( \33241 , \33239 , \33240 );
nand \U$32865 ( \33242 , \22043 , \15267 );
nand \U$32866 ( \33243 , \33241 , \33242 );
and \U$32867 ( \33244 , \33238 , \33243 );
not \U$32868 ( \33245 , \33238 );
not \U$32869 ( \33246 , \33243 );
and \U$32870 ( \33247 , \33245 , \33246 );
nor \U$32871 ( \33248 , \33244 , \33247 );
xor \U$32872 ( \33249 , \33227 , \33248 );
not \U$32873 ( \33250 , \9398 );
not \U$32874 ( \33251 , \22029 );
or \U$32875 ( \33252 , \33250 , \33251 );
nand \U$32876 ( \33253 , \29193 , \9934 );
nand \U$32877 ( \33254 , \33252 , \33253 );
not \U$32878 ( \33255 , \9110 );
not \U$32879 ( \33256 , \28782 );
or \U$32880 ( \33257 , \33255 , \33256 );
nand \U$32881 ( \33258 , \22199 , \9205 );
nand \U$32882 ( \33259 , \33257 , \33258 );
xor \U$32883 ( \33260 , \33254 , \33259 );
not \U$32884 ( \33261 , \13025 );
not \U$32885 ( \33262 , \22176 );
or \U$32886 ( \33263 , \33261 , \33262 );
nand \U$32887 ( \33264 , \28805 , \11118 );
nand \U$32888 ( \33265 , \33263 , \33264 );
xor \U$32889 ( \33266 , \33260 , \33265 );
and \U$32890 ( \33267 , \33249 , \33266 );
and \U$32891 ( \33268 , \33227 , \33248 );
or \U$32892 ( \33269 , \33267 , \33268 );
xor \U$32893 ( \33270 , \33223 , \33269 );
xor \U$32894 ( \33271 , \33114 , \33119 );
and \U$32895 ( \33272 , \33271 , \33125 );
and \U$32896 ( \33273 , \33114 , \33119 );
or \U$32897 ( \33274 , \33272 , \33273 );
not \U$32898 ( \33275 , \33232 );
nand \U$32899 ( \33276 , \33275 , \33246 );
and \U$32900 ( \33277 , \33237 , \33276 );
and \U$32901 ( \33278 , \33232 , \33243 );
nor \U$32902 ( \33279 , \33277 , \33278 );
and \U$32903 ( \33280 , \33274 , \33279 );
not \U$32904 ( \33281 , \33274 );
not \U$32905 ( \33282 , \33279 );
and \U$32906 ( \33283 , \33281 , \33282 );
or \U$32907 ( \33284 , \33280 , \33283 );
not \U$32908 ( \33285 , \12670 );
not \U$32909 ( \33286 , \32958 );
or \U$32910 ( \33287 , \33285 , \33286 );
nand \U$32911 ( \33288 , \28617 , \15164 );
nand \U$32912 ( \33289 , \33287 , \33288 );
not \U$32913 ( \33290 , \33289 );
not \U$32914 ( \33291 , \12945 );
not \U$32915 ( \33292 , \22153 );
or \U$32916 ( \33293 , \33291 , \33292 );
nand \U$32917 ( \33294 , \28632 , \9488 );
nand \U$32918 ( \33295 , \33293 , \33294 );
not \U$32919 ( \33296 , \33295 );
nand \U$32920 ( \33297 , \33290 , \33296 );
not \U$32921 ( \33298 , \9690 );
not \U$32922 ( \33299 , \28787 );
or \U$32923 ( \33300 , \33298 , \33299 );
nand \U$32924 ( \33301 , \22187 , \9816 );
nand \U$32925 ( \33302 , \33300 , \33301 );
and \U$32926 ( \33303 , \33297 , \33302 );
nor \U$32927 ( \33304 , \33290 , \33296 );
nor \U$32928 ( \33305 , \33303 , \33304 );
not \U$32929 ( \33306 , \33305 );
xor \U$32930 ( \33307 , \33284 , \33306 );
xor \U$32931 ( \33308 , \33270 , \33307 );
xor \U$32932 ( \33309 , \33217 , \33308 );
xor \U$32933 ( \33310 , \33136 , \33309 );
xor \U$32934 ( \33311 , \33202 , \33207 );
and \U$32935 ( \33312 , \33311 , \33211 );
not \U$32936 ( \33313 , \33311 );
and \U$32937 ( \33314 , \33313 , \33210 );
nor \U$32938 ( \33315 , \33312 , \33314 );
not \U$32939 ( \33316 , \33315 );
not \U$32940 ( \33317 , \33316 );
xor \U$32941 ( \33318 , \33025 , \33041 );
xnor \U$32942 ( \33319 , \33318 , \33031 );
not \U$32943 ( \33320 , \33319 );
or \U$32944 ( \33321 , \33317 , \33320 );
or \U$32945 ( \33322 , \33316 , \33319 );
xor \U$32946 ( \33323 , \28762 , \28766 );
and \U$32947 ( \33324 , \33323 , \28813 );
and \U$32948 ( \33325 , \28762 , \28766 );
or \U$32949 ( \33326 , \33324 , \33325 );
nand \U$32950 ( \33327 , \33322 , \33326 );
nand \U$32951 ( \33328 , \33321 , \33327 );
xor \U$32952 ( \33329 , \28862 , \28866 );
and \U$32953 ( \33330 , \33329 , \28898 );
and \U$32954 ( \33331 , \28862 , \28866 );
or \U$32955 ( \33332 , \33330 , \33331 );
and \U$32956 ( \33333 , \33302 , \33295 );
not \U$32957 ( \33334 , \33302 );
and \U$32958 ( \33335 , \33334 , \33296 );
nor \U$32959 ( \33336 , \33333 , \33335 );
and \U$32960 ( \33337 , \33336 , \33289 );
not \U$32961 ( \33338 , \33336 );
and \U$32962 ( \33339 , \33338 , \33290 );
nor \U$32963 ( \33340 , \33337 , \33339 );
xor \U$32964 ( \33341 , \33332 , \33340 );
xor \U$32965 ( \33342 , \32976 , \32980 );
xor \U$32966 ( \33343 , \33342 , \32987 );
xnor \U$32967 ( \33344 , \33341 , \33343 );
not \U$32968 ( \33345 , \33344 );
not \U$32969 ( \33346 , \28899 );
nand \U$32970 ( \33347 , \33346 , \28830 );
and \U$32971 ( \33348 , \28912 , \33347 );
nor \U$32972 ( \33349 , \28830 , \28902 );
nor \U$32973 ( \33350 , \33348 , \33349 );
not \U$32974 ( \33351 , \33350 );
or \U$32975 ( \33352 , \33345 , \33351 );
xor \U$32976 ( \33353 , \33227 , \33248 );
xor \U$32977 ( \33354 , \33353 , \33266 );
nand \U$32978 ( \33355 , \33352 , \33354 );
not \U$32979 ( \33356 , \33350 );
not \U$32980 ( \33357 , \33344 );
nand \U$32981 ( \33358 , \33356 , \33357 );
nand \U$32982 ( \33359 , \33355 , \33358 );
xor \U$32983 ( \33360 , \33328 , \33359 );
xor \U$32984 ( \33361 , \21983 , \21993 );
xor \U$32985 ( \33362 , \33361 , \22003 );
xor \U$32986 ( \33363 , \21884 , \21896 );
xor \U$32987 ( \33364 , \33363 , \21873 );
xor \U$32988 ( \33365 , \33362 , \33364 );
xor \U$32989 ( \33366 , \33254 , \33259 );
and \U$32990 ( \33367 , \33366 , \33265 );
and \U$32991 ( \33368 , \33254 , \33259 );
or \U$32992 ( \33369 , \33367 , \33368 );
xnor \U$32993 ( \33370 , \33365 , \33369 );
not \U$32994 ( \33371 , \33343 );
buf \U$32995 ( \33372 , \33340 );
not \U$32996 ( \33373 , \33372 );
or \U$32997 ( \33374 , \33371 , \33373 );
or \U$32998 ( \33375 , \33372 , \33343 );
nand \U$32999 ( \33376 , \33375 , \33332 );
nand \U$33000 ( \33377 , \33374 , \33376 );
xor \U$33001 ( \33378 , \33370 , \33377 );
xor \U$33002 ( \33379 , \22135 , \22146 );
xor \U$33003 ( \33380 , \33379 , \22157 );
xor \U$33004 ( \33381 , \22091 , \22101 );
xor \U$33005 ( \33382 , \33381 , \22112 );
xor \U$33006 ( \33383 , \33380 , \33382 );
xor \U$33007 ( \33384 , \22180 , \22189 );
xor \U$33008 ( \33385 , \33384 , \22201 );
xor \U$33009 ( \33386 , \33383 , \33385 );
xor \U$33010 ( \33387 , \33378 , \33386 );
xnor \U$33011 ( \33388 , \33360 , \33387 );
not \U$33012 ( \33389 , \29087 );
not \U$33013 ( \33390 , \29095 );
or \U$33014 ( \33391 , \33389 , \33390 );
not \U$33015 ( \33392 , \29088 );
not \U$33016 ( \33393 , \29094 );
or \U$33017 ( \33394 , \33392 , \33393 );
nand \U$33018 ( \33395 , \33394 , \29106 );
nand \U$33019 ( \33396 , \33391 , \33395 );
not \U$33020 ( \33397 , \33396 );
not \U$33021 ( \33398 , \33397 );
and \U$33022 ( \33399 , \33319 , \33315 );
not \U$33023 ( \33400 , \33319 );
and \U$33024 ( \33401 , \33400 , \33316 );
nor \U$33025 ( \33402 , \33399 , \33401 );
xor \U$33026 ( \33403 , \33402 , \33326 );
not \U$33027 ( \33404 , \33403 );
or \U$33028 ( \33405 , \33398 , \33404 );
xor \U$33029 ( \33406 , \28719 , \28814 );
and \U$33030 ( \33407 , \33406 , \28819 );
and \U$33031 ( \33408 , \28719 , \28814 );
or \U$33032 ( \33409 , \33407 , \33408 );
nand \U$33033 ( \33410 , \33405 , \33409 );
not \U$33034 ( \33411 , \33397 );
not \U$33035 ( \33412 , \33403 );
nand \U$33036 ( \33413 , \33411 , \33412 );
nand \U$33037 ( \33414 , \33410 , \33413 );
not \U$33038 ( \33415 , \33414 );
and \U$33039 ( \33416 , \33388 , \33415 );
not \U$33040 ( \33417 , \33388 );
and \U$33041 ( \33418 , \33417 , \33414 );
nor \U$33042 ( \33419 , \33416 , \33418 );
not \U$33043 ( \33420 , \33357 );
not \U$33044 ( \33421 , \33420 );
not \U$33045 ( \33422 , \33354 );
and \U$33046 ( \33423 , \33350 , \33422 );
not \U$33047 ( \33424 , \33350 );
and \U$33048 ( \33425 , \33424 , \33354 );
nor \U$33049 ( \33426 , \33423 , \33425 );
not \U$33050 ( \33427 , \33426 );
or \U$33051 ( \33428 , \33421 , \33427 );
or \U$33052 ( \33429 , \33426 , \33420 );
nand \U$33053 ( \33430 , \33428 , \33429 );
not \U$33054 ( \33431 , \28913 );
not \U$33055 ( \33432 , \28917 );
or \U$33056 ( \33433 , \33431 , \33432 );
or \U$33057 ( \33434 , \28913 , \28917 );
nand \U$33058 ( \33435 , \33434 , \28922 );
nand \U$33059 ( \33436 , \33433 , \33435 );
xor \U$33060 ( \33437 , \33430 , \33436 );
xor \U$33061 ( \33438 , \33062 , \33068 );
xor \U$33062 ( \33439 , \33438 , \33132 );
and \U$33063 ( \33440 , \33437 , \33439 );
and \U$33064 ( \33441 , \33430 , \33436 );
or \U$33065 ( \33442 , \33440 , \33441 );
not \U$33066 ( \33443 , \33442 );
and \U$33067 ( \33444 , \33419 , \33443 );
not \U$33068 ( \33445 , \33419 );
and \U$33069 ( \33446 , \33445 , \33442 );
or \U$33070 ( \33447 , \33444 , \33446 );
xor \U$33071 ( \33448 , \33310 , \33447 );
xor \U$33072 ( \33449 , \29071 , \29111 );
and \U$33073 ( \33450 , \33449 , \29280 );
and \U$33074 ( \33451 , \29071 , \29111 );
or \U$33075 ( \33452 , \33450 , \33451 );
not \U$33076 ( \33453 , \33452 );
xor \U$33077 ( \33454 , \33396 , \33403 );
xnor \U$33078 ( \33455 , \33454 , \33409 );
not \U$33079 ( \33456 , \33455 );
nand \U$33080 ( \33457 , \33453 , \33456 );
not \U$33081 ( \33458 , \33457 );
xor \U$33082 ( \33459 , \33430 , \33436 );
xor \U$33083 ( \33460 , \33459 , \33439 );
not \U$33084 ( \33461 , \33460 );
or \U$33085 ( \33462 , \33458 , \33461 );
nand \U$33086 ( \33463 , \33455 , \33452 );
nand \U$33087 ( \33464 , \33462 , \33463 );
xnor \U$33088 ( \33465 , \33448 , \33464 );
not \U$33089 ( \33466 , \33465 );
not \U$33090 ( \33467 , \28820 );
not \U$33091 ( \33468 , \28935 );
or \U$33092 ( \33469 , \33467 , \33468 );
not \U$33093 ( \33470 , \28821 );
not \U$33094 ( \33471 , \28932 );
or \U$33095 ( \33472 , \33470 , \33471 );
nand \U$33096 ( \33473 , \33472 , \28924 );
nand \U$33097 ( \33474 , \33469 , \33473 );
not \U$33098 ( \33475 , \28949 );
not \U$33099 ( \33476 , \33475 );
not \U$33100 ( \33477 , \29281 );
or \U$33101 ( \33478 , \33476 , \33477 );
not \U$33102 ( \33479 , \28949 );
not \U$33103 ( \33480 , \29281 );
not \U$33104 ( \33481 , \33480 );
or \U$33105 ( \33482 , \33479 , \33481 );
nand \U$33106 ( \33483 , \33482 , \29587 );
nand \U$33107 ( \33484 , \33478 , \33483 );
xor \U$33108 ( \33485 , \33474 , \33484 );
not \U$33109 ( \33486 , \33460 );
and \U$33110 ( \33487 , \33452 , \33456 );
not \U$33111 ( \33488 , \33452 );
and \U$33112 ( \33489 , \33488 , \33455 );
nor \U$33113 ( \33490 , \33487 , \33489 );
not \U$33114 ( \33491 , \33490 );
or \U$33115 ( \33492 , \33486 , \33491 );
or \U$33116 ( \33493 , \33460 , \33490 );
nand \U$33117 ( \33494 , \33492 , \33493 );
and \U$33118 ( \33495 , \33485 , \33494 );
and \U$33119 ( \33496 , \33474 , \33484 );
or \U$33120 ( \33497 , \33495 , \33496 );
not \U$33121 ( \33498 , \33497 );
nand \U$33122 ( \33499 , \33466 , \33498 );
xor \U$33123 ( \33500 , \32990 , \33022 );
and \U$33124 ( \33501 , \33500 , \33043 );
and \U$33125 ( \33502 , \32990 , \33022 );
or \U$33126 ( \33503 , \33501 , \33502 );
xor \U$33127 ( \33504 , \33156 , \33191 );
and \U$33128 ( \33505 , \33504 , \33215 );
and \U$33129 ( \33506 , \33156 , \33191 );
or \U$33130 ( \33507 , \33505 , \33506 );
xor \U$33131 ( \33508 , \33503 , \33507 );
not \U$33132 ( \33509 , \22120 );
not \U$33133 ( \33510 , \22117 );
or \U$33134 ( \33511 , \33509 , \33510 );
or \U$33135 ( \33512 , \22117 , \22120 );
nand \U$33136 ( \33513 , \33511 , \33512 );
xor \U$33137 ( \33514 , \22115 , \33513 );
not \U$33138 ( \33515 , \22006 );
not \U$33139 ( \33516 , \21941 );
or \U$33140 ( \33517 , \33515 , \33516 );
not \U$33141 ( \33518 , \22006 );
nand \U$33142 ( \33519 , \33518 , \21938 );
nand \U$33143 ( \33520 , \33517 , \33519 );
and \U$33144 ( \33521 , \33520 , \21900 );
not \U$33145 ( \33522 , \33520 );
and \U$33146 ( \33523 , \33522 , \21899 );
nor \U$33147 ( \33524 , \33521 , \33523 );
xor \U$33148 ( \33525 , \33514 , \33524 );
not \U$33149 ( \33526 , \33364 );
not \U$33150 ( \33527 , \33369 );
or \U$33151 ( \33528 , \33526 , \33527 );
or \U$33152 ( \33529 , \33369 , \33364 );
nand \U$33153 ( \33530 , \33529 , \33362 );
nand \U$33154 ( \33531 , \33528 , \33530 );
xor \U$33155 ( \33532 , \33525 , \33531 );
xnor \U$33156 ( \33533 , \33508 , \33532 );
not \U$33157 ( \33534 , \33533 );
not \U$33158 ( \33535 , \33534 );
xor \U$33159 ( \33536 , \33144 , \33216 );
and \U$33160 ( \33537 , \33536 , \33308 );
and \U$33161 ( \33538 , \33144 , \33216 );
or \U$33162 ( \33539 , \33537 , \33538 );
not \U$33163 ( \33540 , \33539 );
not \U$33164 ( \33541 , \33540 );
or \U$33165 ( \33542 , \33535 , \33541 );
nand \U$33166 ( \33543 , \33539 , \33533 );
nand \U$33167 ( \33544 , \33542 , \33543 );
xor \U$33168 ( \33545 , \21145 , \21200 );
xor \U$33169 ( \33546 , \33545 , \21210 );
xor \U$33170 ( \33547 , \33158 , \33183 );
and \U$33171 ( \33548 , \33547 , \33190 );
and \U$33172 ( \33549 , \33158 , \33183 );
or \U$33173 ( \33550 , \33548 , \33549 );
xor \U$33174 ( \33551 , \33546 , \33550 );
not \U$33175 ( \33552 , \33282 );
not \U$33176 ( \33553 , \33306 );
or \U$33177 ( \33554 , \33552 , \33553 );
not \U$33178 ( \33555 , \33279 );
not \U$33179 ( \33556 , \33305 );
or \U$33180 ( \33557 , \33555 , \33556 );
nand \U$33181 ( \33558 , \33557 , \33274 );
nand \U$33182 ( \33559 , \33554 , \33558 );
xor \U$33183 ( \33560 , \33551 , \33559 );
xor \U$33184 ( \33561 , \33223 , \33269 );
and \U$33185 ( \33562 , \33561 , \33307 );
and \U$33186 ( \33563 , \33223 , \33269 );
or \U$33187 ( \33564 , \33562 , \33563 );
xor \U$33188 ( \33565 , \33560 , \33564 );
xor \U$33189 ( \33566 , \22020 , \22022 );
xor \U$33190 ( \33567 , \33566 , \22060 );
not \U$33191 ( \33568 , \32925 );
nand \U$33192 ( \33569 , \33568 , \32970 );
not \U$33193 ( \33570 , \33569 );
not \U$33194 ( \33571 , \32963 );
or \U$33195 ( \33572 , \33570 , \33571 );
nand \U$33196 ( \33573 , \32971 , \32925 );
nand \U$33197 ( \33574 , \33572 , \33573 );
xor \U$33198 ( \33575 , \33567 , \33574 );
xor \U$33199 ( \33576 , \33380 , \33382 );
and \U$33200 ( \33577 , \33576 , \33385 );
and \U$33201 ( \33578 , \33380 , \33382 );
or \U$33202 ( \33579 , \33577 , \33578 );
xor \U$33203 ( \33580 , \33575 , \33579 );
xnor \U$33204 ( \33581 , \33565 , \33580 );
xor \U$33205 ( \33582 , \33544 , \33581 );
not \U$33206 ( \33583 , \33443 );
buf \U$33207 ( \33584 , \33388 );
nor \U$33208 ( \33585 , \33584 , \33414 );
not \U$33209 ( \33586 , \33585 );
and \U$33210 ( \33587 , \33583 , \33586 );
and \U$33211 ( \33588 , \33584 , \33414 );
nor \U$33212 ( \33589 , \33587 , \33588 );
xor \U$33213 ( \33590 , \33582 , \33589 );
not \U$33214 ( \33591 , \33359 );
nand \U$33215 ( \33592 , \33591 , \33387 );
and \U$33216 ( \33593 , \33592 , \33328 );
not \U$33217 ( \33594 , \33359 );
nor \U$33218 ( \33595 , \33594 , \33387 );
nor \U$33219 ( \33596 , \33593 , \33595 );
not \U$33220 ( \33597 , \33377 );
not \U$33221 ( \33598 , \33386 );
or \U$33222 ( \33599 , \33597 , \33598 );
or \U$33223 ( \33600 , \33377 , \33386 );
not \U$33224 ( \33601 , \33370 );
nand \U$33225 ( \33602 , \33600 , \33601 );
nand \U$33226 ( \33603 , \33599 , \33602 );
xor \U$33227 ( \33604 , \22160 , \22169 );
xor \U$33228 ( \33605 , \33604 , \22204 );
not \U$33229 ( \33606 , \33605 );
not \U$33230 ( \33607 , \21273 );
not \U$33231 ( \33608 , \21301 );
not \U$33232 ( \33609 , \33608 );
or \U$33233 ( \33610 , \33607 , \33609 );
nand \U$33234 ( \33611 , \21301 , \21289 );
nand \U$33235 ( \33612 , \33610 , \33611 );
and \U$33236 ( \33613 , \33612 , \21285 );
not \U$33237 ( \33614 , \33612 );
and \U$33238 ( \33615 , \33614 , \21286 );
nor \U$33239 ( \33616 , \33613 , \33615 );
xor \U$33240 ( \33617 , \21388 , \21398 );
xor \U$33241 ( \33618 , \33617 , \21409 );
xor \U$33242 ( \33619 , \33616 , \33618 );
xor \U$33243 ( \33620 , \33146 , \33150 );
and \U$33244 ( \33621 , \33620 , \33155 );
and \U$33245 ( \33622 , \33146 , \33150 );
or \U$33246 ( \33623 , \33621 , \33622 );
xor \U$33247 ( \33624 , \33619 , \33623 );
not \U$33248 ( \33625 , \33624 );
or \U$33249 ( \33626 , \33606 , \33625 );
or \U$33250 ( \33627 , \33605 , \33624 );
nand \U$33251 ( \33628 , \33626 , \33627 );
and \U$33252 ( \33629 , \21327 , \21332 );
not \U$33253 ( \33630 , \21327 );
and \U$33254 ( \33631 , \33630 , \21333 );
nor \U$33255 ( \33632 , \33629 , \33631 );
not \U$33256 ( \33633 , \21316 );
and \U$33257 ( \33634 , \33632 , \33633 );
not \U$33258 ( \33635 , \33632 );
and \U$33259 ( \33636 , \33635 , \21316 );
nor \U$33260 ( \33637 , \33634 , \33636 );
xor \U$33261 ( \33638 , \32941 , \32952 );
and \U$33262 ( \33639 , \33638 , \32962 );
and \U$33263 ( \33640 , \32941 , \32952 );
or \U$33264 ( \33641 , \33639 , \33640 );
xor \U$33265 ( \33642 , \33637 , \33641 );
xor \U$33266 ( \33643 , \20901 , \20910 );
xor \U$33267 ( \33644 , \33643 , \20926 );
xor \U$33268 ( \33645 , \33642 , \33644 );
xor \U$33269 ( \33646 , \33628 , \33645 );
xor \U$33270 ( \33647 , \33603 , \33646 );
xor \U$33271 ( \33648 , \32972 , \33044 );
and \U$33272 ( \33649 , \33648 , \33059 );
and \U$33273 ( \33650 , \32972 , \33044 );
or \U$33274 ( \33651 , \33649 , \33650 );
xnor \U$33275 ( \33652 , \33647 , \33651 );
xor \U$33276 ( \33653 , \33596 , \33652 );
not \U$33277 ( \33654 , \33309 );
not \U$33278 ( \33655 , \33060 );
nand \U$33279 ( \33656 , \33654 , \33655 );
and \U$33280 ( \33657 , \33656 , \33135 );
nor \U$33281 ( \33658 , \33654 , \33655 );
nor \U$33282 ( \33659 , \33657 , \33658 );
xor \U$33283 ( \33660 , \33653 , \33659 );
xor \U$33284 ( \33661 , \33590 , \33660 );
not \U$33285 ( \33662 , \33310 );
buf \U$33286 ( \33663 , \33447 );
nand \U$33287 ( \33664 , \33662 , \33663 );
and \U$33288 ( \33665 , \33664 , \33464 );
not \U$33289 ( \33666 , \33310 );
nor \U$33290 ( \33667 , \33666 , \33663 );
nor \U$33291 ( \33668 , \33665 , \33667 );
nand \U$33292 ( \33669 , \33661 , \33668 );
xor \U$33293 ( \33670 , \33546 , \33550 );
and \U$33294 ( \33671 , \33670 , \33559 );
and \U$33295 ( \33672 , \33546 , \33550 );
or \U$33296 ( \33673 , \33671 , \33672 );
xor \U$33297 ( \33674 , \33514 , \33524 );
and \U$33298 ( \33675 , \33674 , \33531 );
and \U$33299 ( \33676 , \33514 , \33524 );
or \U$33300 ( \33677 , \33675 , \33676 );
xor \U$33301 ( \33678 , \33673 , \33677 );
xor \U$33302 ( \33679 , \33567 , \33574 );
and \U$33303 ( \33680 , \33679 , \33579 );
and \U$33304 ( \33681 , \33567 , \33574 );
or \U$33305 ( \33682 , \33680 , \33681 );
xor \U$33306 ( \33683 , \33678 , \33682 );
not \U$33307 ( \33684 , \33560 );
not \U$33308 ( \33685 , \33580 );
or \U$33309 ( \33686 , \33684 , \33685 );
or \U$33310 ( \33687 , \33580 , \33560 );
nand \U$33311 ( \33688 , \33687 , \33564 );
nand \U$33312 ( \33689 , \33686 , \33688 );
xor \U$33313 ( \33690 , \33683 , \33689 );
not \U$33314 ( \33691 , \22014 );
not \U$33315 ( \33692 , \22011 );
or \U$33316 ( \33693 , \33691 , \33692 );
or \U$33317 ( \33694 , \22011 , \22014 );
nand \U$33318 ( \33695 , \33693 , \33694 );
xor \U$33319 ( \33696 , \22063 , \33695 );
xor \U$33320 ( \33697 , \22125 , \22207 );
xor \U$33321 ( \33698 , \33697 , \22210 );
xor \U$33322 ( \33699 , \33696 , \33698 );
xor \U$33323 ( \33700 , \33637 , \33641 );
and \U$33324 ( \33701 , \33700 , \33644 );
and \U$33325 ( \33702 , \33637 , \33641 );
or \U$33326 ( \33703 , \33701 , \33702 );
xor \U$33327 ( \33704 , \21420 , \21412 );
xnor \U$33328 ( \33705 , \33704 , \21377 );
xor \U$33329 ( \33706 , \21303 , \21262 );
xnor \U$33330 ( \33707 , \33706 , \21335 );
and \U$33331 ( \33708 , \33705 , \33707 );
not \U$33332 ( \33709 , \33705 );
not \U$33333 ( \33710 , \33707 );
and \U$33334 ( \33711 , \33709 , \33710 );
nor \U$33335 ( \33712 , \33708 , \33711 );
xor \U$33336 ( \33713 , \33703 , \33712 );
xor \U$33337 ( \33714 , \33699 , \33713 );
xnor \U$33338 ( \33715 , \33690 , \33714 );
not \U$33339 ( \33716 , \33603 );
not \U$33340 ( \33717 , \33646 );
or \U$33341 ( \33718 , \33716 , \33717 );
or \U$33342 ( \33719 , \33646 , \33603 );
nand \U$33343 ( \33720 , \33719 , \33651 );
nand \U$33344 ( \33721 , \33718 , \33720 );
not \U$33345 ( \33722 , \33624 );
not \U$33346 ( \33723 , \33722 );
not \U$33347 ( \33724 , \33605 );
or \U$33348 ( \33725 , \33723 , \33724 );
not \U$33349 ( \33726 , \33605 );
not \U$33350 ( \33727 , \33726 );
not \U$33351 ( \33728 , \33624 );
or \U$33352 ( \33729 , \33727 , \33728 );
nand \U$33353 ( \33730 , \33729 , \33645 );
nand \U$33354 ( \33731 , \33725 , \33730 );
not \U$33355 ( \33732 , \33618 );
nand \U$33356 ( \33733 , \33732 , \33616 );
not \U$33357 ( \33734 , \33733 );
not \U$33358 ( \33735 , \33623 );
or \U$33359 ( \33736 , \33734 , \33735 );
not \U$33360 ( \33737 , \33616 );
nand \U$33361 ( \33738 , \33737 , \33618 );
nand \U$33362 ( \33739 , \33736 , \33738 );
xor \U$33363 ( \33740 , \21838 , \21840 );
xor \U$33364 ( \33741 , \33740 , \21850 );
xor \U$33365 ( \33742 , \33739 , \33741 );
xor \U$33366 ( \33743 , \21213 , \21215 );
xor \U$33367 ( \33744 , \33743 , \21218 );
xor \U$33368 ( \33745 , \33742 , \33744 );
xor \U$33369 ( \33746 , \33731 , \33745 );
or \U$33370 ( \33747 , \33503 , \33507 );
nand \U$33371 ( \33748 , \33747 , \33532 );
nand \U$33372 ( \33749 , \33503 , \33507 );
nand \U$33373 ( \33750 , \33748 , \33749 );
xor \U$33374 ( \33751 , \33746 , \33750 );
not \U$33375 ( \33752 , \33751 );
and \U$33376 ( \33753 , \33721 , \33752 );
not \U$33377 ( \33754 , \33721 );
and \U$33378 ( \33755 , \33754 , \33751 );
nor \U$33379 ( \33756 , \33753 , \33755 );
not \U$33380 ( \33757 , \33756 );
not \U$33381 ( \33758 , \33534 );
not \U$33382 ( \33759 , \33581 );
not \U$33383 ( \33760 , \33759 );
or \U$33384 ( \33761 , \33758 , \33760 );
not \U$33385 ( \33762 , \33533 );
not \U$33386 ( \33763 , \33581 );
or \U$33387 ( \33764 , \33762 , \33763 );
nand \U$33388 ( \33765 , \33764 , \33539 );
nand \U$33389 ( \33766 , \33761 , \33765 );
not \U$33390 ( \33767 , \33766 );
and \U$33391 ( \33768 , \33757 , \33767 );
and \U$33392 ( \33769 , \33766 , \33756 );
nor \U$33393 ( \33770 , \33768 , \33769 );
xor \U$33394 ( \33771 , \33715 , \33770 );
xor \U$33395 ( \33772 , \33596 , \33652 );
and \U$33396 ( \33773 , \33772 , \33659 );
and \U$33397 ( \33774 , \33596 , \33652 );
or \U$33398 ( \33775 , \33773 , \33774 );
xor \U$33399 ( \33776 , \33771 , \33775 );
xor \U$33400 ( \33777 , \33582 , \33589 );
and \U$33401 ( \33778 , \33777 , \33660 );
and \U$33402 ( \33779 , \33582 , \33589 );
or \U$33403 ( \33780 , \33778 , \33779 );
nand \U$33404 ( \33781 , \33776 , \33780 );
not \U$33405 ( \33782 , \29592 );
not \U$33406 ( \33783 , \28937 );
or \U$33407 ( \33784 , \33782 , \33783 );
nand \U$33408 ( \33785 , \33784 , \28590 );
not \U$33409 ( \33786 , \28937 );
nand \U$33410 ( \33787 , \33786 , \29593 );
nand \U$33411 ( \33788 , \33785 , \33787 );
not \U$33412 ( \33789 , \33788 );
xor \U$33413 ( \33790 , \33474 , \33484 );
xor \U$33414 ( \33791 , \33790 , \33494 );
not \U$33415 ( \33792 , \33791 );
nand \U$33416 ( \33793 , \33789 , \33792 );
and \U$33417 ( \33794 , \33499 , \33669 , \33781 , \33793 );
not \U$33418 ( \33795 , \33794 );
nor \U$33419 ( \33796 , \32907 , \33795 );
not \U$33420 ( \33797 , \33781 );
not \U$33421 ( \33798 , \33497 );
not \U$33422 ( \33799 , \33465 );
or \U$33423 ( \33800 , \33798 , \33799 );
nand \U$33424 ( \33801 , \33791 , \33788 );
nand \U$33425 ( \33802 , \33800 , \33801 );
nand \U$33426 ( \33803 , \33802 , \33499 );
not \U$33427 ( \33804 , \33669 );
or \U$33428 ( \33805 , \33803 , \33804 );
or \U$33429 ( \33806 , \33661 , \33668 );
nand \U$33430 ( \33807 , \33805 , \33806 );
not \U$33431 ( \33808 , \33807 );
or \U$33432 ( \33809 , \33797 , \33808 );
or \U$33433 ( \33810 , \33776 , \33780 );
nand \U$33434 ( \33811 , \33809 , \33810 );
or \U$33435 ( \33812 , \33796 , \33811 );
xor \U$33436 ( \33813 , \22084 , \22216 );
xnor \U$33437 ( \33814 , \33813 , \22213 );
xor \U$33438 ( \33815 , \33696 , \33698 );
and \U$33439 ( \33816 , \33815 , \33713 );
and \U$33440 ( \33817 , \33696 , \33698 );
or \U$33441 ( \33818 , \33816 , \33817 );
not \U$33442 ( \33819 , \33818 );
xor \U$33443 ( \33820 , \33814 , \33819 );
xor \U$33444 ( \33821 , \33739 , \33741 );
and \U$33445 ( \33822 , \33821 , \33744 );
and \U$33446 ( \33823 , \33739 , \33741 );
or \U$33447 ( \33824 , \33822 , \33823 );
not \U$33448 ( \33825 , \33710 );
not \U$33449 ( \33826 , \33705 );
not \U$33450 ( \33827 , \33826 );
or \U$33451 ( \33828 , \33825 , \33827 );
not \U$33452 ( \33829 , \33707 );
not \U$33453 ( \33830 , \33705 );
or \U$33454 ( \33831 , \33829 , \33830 );
nand \U$33455 ( \33832 , \33831 , \33703 );
nand \U$33456 ( \33833 , \33828 , \33832 );
xor \U$33457 ( \33834 , \33824 , \33833 );
xor \U$33458 ( \33835 , \20846 , \20879 );
xor \U$33459 ( \33836 , \33835 , \20955 );
xor \U$33460 ( \33837 , \33834 , \33836 );
xor \U$33461 ( \33838 , \33820 , \33837 );
not \U$33462 ( \33839 , \33721 );
nand \U$33463 ( \33840 , \33839 , \33752 );
not \U$33464 ( \33841 , \33840 );
not \U$33465 ( \33842 , \33766 );
or \U$33466 ( \33843 , \33841 , \33842 );
not \U$33467 ( \33844 , \33752 );
nand \U$33468 ( \33845 , \33844 , \33721 );
nand \U$33469 ( \33846 , \33843 , \33845 );
not \U$33470 ( \33847 , \33846 );
xor \U$33471 ( \33848 , \33838 , \33847 );
xor \U$33472 ( \33849 , \33731 , \33745 );
and \U$33473 ( \33850 , \33849 , \33750 );
and \U$33474 ( \33851 , \33731 , \33745 );
or \U$33475 ( \33852 , \33850 , \33851 );
not \U$33476 ( \33853 , \33852 );
xor \U$33477 ( \33854 , \21001 , \21078 );
xor \U$33478 ( \33855 , \33854 , \21221 );
xor \U$33479 ( \33856 , \21853 , \21860 );
xor \U$33480 ( \33857 , \33856 , \22065 );
xor \U$33481 ( \33858 , \33855 , \33857 );
xor \U$33482 ( \33859 , \33673 , \33677 );
and \U$33483 ( \33860 , \33859 , \33682 );
and \U$33484 ( \33861 , \33673 , \33677 );
or \U$33485 ( \33862 , \33860 , \33861 );
xor \U$33486 ( \33863 , \33858 , \33862 );
not \U$33487 ( \33864 , \33863 );
not \U$33488 ( \33865 , \33864 );
or \U$33489 ( \33866 , \33853 , \33865 );
not \U$33490 ( \33867 , \33852 );
nand \U$33491 ( \33868 , \33867 , \33863 );
nand \U$33492 ( \33869 , \33866 , \33868 );
not \U$33493 ( \33870 , \33683 );
not \U$33494 ( \33871 , \33714 );
or \U$33495 ( \33872 , \33870 , \33871 );
or \U$33496 ( \33873 , \33714 , \33683 );
nand \U$33497 ( \33874 , \33873 , \33689 );
nand \U$33498 ( \33875 , \33872 , \33874 );
not \U$33499 ( \33876 , \33875 );
and \U$33500 ( \33877 , \33869 , \33876 );
not \U$33501 ( \33878 , \33869 );
and \U$33502 ( \33879 , \33878 , \33875 );
nor \U$33503 ( \33880 , \33877 , \33879 );
xor \U$33504 ( \33881 , \33848 , \33880 );
xor \U$33505 ( \33882 , \33715 , \33770 );
and \U$33506 ( \33883 , \33882 , \33775 );
and \U$33507 ( \33884 , \33715 , \33770 );
or \U$33508 ( \33885 , \33883 , \33884 );
nand \U$33509 ( \33886 , \33881 , \33885 );
xor \U$33510 ( \33887 , \20844 , \20958 );
xor \U$33511 ( \33888 , \33887 , \21224 );
xor \U$33512 ( \33889 , \21663 , \21665 );
not \U$33513 ( \33890 , \33889 );
not \U$33514 ( \33891 , \33890 );
not \U$33515 ( \33892 , \21694 );
or \U$33516 ( \33893 , \33891 , \33892 );
not \U$33517 ( \33894 , \21694 );
nand \U$33518 ( \33895 , \33894 , \33889 );
nand \U$33519 ( \33896 , \33893 , \33895 );
xor \U$33520 ( \33897 , \33888 , \33896 );
not \U$33521 ( \33898 , \33833 );
not \U$33522 ( \33899 , \33836 );
or \U$33523 ( \33900 , \33898 , \33899 );
or \U$33524 ( \33901 , \33836 , \33833 );
nand \U$33525 ( \33902 , \33901 , \33824 );
nand \U$33526 ( \33903 , \33900 , \33902 );
and \U$33527 ( \33904 , \33897 , \33903 );
and \U$33528 ( \33905 , \33888 , \33896 );
nor \U$33529 ( \33906 , \33904 , \33905 );
xor \U$33530 ( \33907 , \33855 , \33857 );
and \U$33531 ( \33908 , \33907 , \33862 );
and \U$33532 ( \33909 , \33855 , \33857 );
or \U$33533 ( \33910 , \33908 , \33909 );
not \U$33534 ( \33911 , \33910 );
not \U$33535 ( \33912 , \22079 );
not \U$33536 ( \33913 , \22076 );
or \U$33537 ( \33914 , \33912 , \33913 );
nand \U$33538 ( \33915 , \22075 , \22068 );
nand \U$33539 ( \33916 , \33914 , \33915 );
not \U$33540 ( \33917 , \22218 );
and \U$33541 ( \33918 , \33916 , \33917 );
not \U$33542 ( \33919 , \33916 );
and \U$33543 ( \33920 , \33919 , \22218 );
nor \U$33544 ( \33921 , \33918 , \33920 );
nand \U$33545 ( \33922 , \33911 , \33921 );
not \U$33546 ( \33923 , \33922 );
xor \U$33547 ( \33924 , \33903 , \33888 );
xor \U$33548 ( \33925 , \33924 , \33896 );
not \U$33549 ( \33926 , \33925 );
or \U$33550 ( \33927 , \33923 , \33926 );
not \U$33551 ( \33928 , \33921 );
nand \U$33552 ( \33929 , \33928 , \33910 );
nand \U$33553 ( \33930 , \33927 , \33929 );
not \U$33554 ( \33931 , \33930 );
xor \U$33555 ( \33932 , \33906 , \33931 );
xor \U$33556 ( \33933 , \22220 , \22226 );
xor \U$33557 ( \33934 , \33933 , \22230 );
xor \U$33558 ( \33935 , \33932 , \33934 );
xor \U$33559 ( \33936 , \33910 , \33921 );
xnor \U$33560 ( \33937 , \33936 , \33925 );
not \U$33561 ( \33938 , \33814 );
nand \U$33562 ( \33939 , \33938 , \33819 );
not \U$33563 ( \33940 , \33939 );
not \U$33564 ( \33941 , \33837 );
or \U$33565 ( \33942 , \33940 , \33941 );
nand \U$33566 ( \33943 , \33818 , \33814 );
nand \U$33567 ( \33944 , \33942 , \33943 );
or \U$33568 ( \33945 , \33937 , \33944 );
not \U$33569 ( \33946 , \33875 );
not \U$33570 ( \33947 , \33852 );
nand \U$33571 ( \33948 , \33864 , \33947 );
not \U$33572 ( \33949 , \33948 );
or \U$33573 ( \33950 , \33946 , \33949 );
not \U$33574 ( \33951 , \33947 );
nand \U$33575 ( \33952 , \33951 , \33863 );
nand \U$33576 ( \33953 , \33950 , \33952 );
nand \U$33577 ( \33954 , \33945 , \33953 );
nand \U$33578 ( \33955 , \33937 , \33944 );
and \U$33579 ( \33956 , \33954 , \33955 );
nand \U$33580 ( \33957 , \33935 , \33956 );
xor \U$33581 ( \33958 , \33944 , \33953 );
xnor \U$33582 ( \33959 , \33958 , \33937 );
xor \U$33583 ( \33960 , \33838 , \33847 );
and \U$33584 ( \33961 , \33960 , \33880 );
and \U$33585 ( \33962 , \33838 , \33847 );
or \U$33586 ( \33963 , \33961 , \33962 );
nand \U$33587 ( \33964 , \33959 , \33963 );
xor \U$33588 ( \33965 , \33906 , \33931 );
and \U$33589 ( \33966 , \33965 , \33934 );
and \U$33590 ( \33967 , \33906 , \33931 );
or \U$33591 ( \33968 , \33966 , \33967 );
xor \U$33592 ( \33969 , \21824 , \22235 );
xnor \U$33593 ( \33970 , \33969 , \21835 );
nand \U$33594 ( \33971 , \33968 , \33970 );
and \U$33595 ( \33972 , \33886 , \33957 , \33964 , \33971 );
nand \U$33596 ( \33973 , \33812 , \33972 );
not \U$33597 ( \33974 , \13025 );
not \U$33598 ( \33975 , RIc225c60_55);
not \U$33599 ( \33976 , \6076 );
or \U$33600 ( \33977 , \33975 , \33976 );
nand \U$33601 ( \33978 , \4407 , \8767 );
nand \U$33602 ( \33979 , \33977 , \33978 );
not \U$33603 ( \33980 , \33979 );
or \U$33604 ( \33981 , \33974 , \33980 );
not \U$33605 ( \33982 , RIc225c60_55);
not \U$33606 ( \33983 , \9850 );
or \U$33607 ( \33984 , \33982 , \33983 );
nand \U$33608 ( \33985 , \10231 , \11108 );
nand \U$33609 ( \33986 , \33984 , \33985 );
nand \U$33610 ( \33987 , \33986 , \11118 );
nand \U$33611 ( \33988 , \33981 , \33987 );
not \U$33612 ( \33989 , \5135 );
not \U$33613 ( \33990 , RIc2265c0_35);
not \U$33614 ( \33991 , \10263 );
or \U$33615 ( \33992 , \33990 , \33991 );
nand \U$33616 ( \33993 , \16998 , \4376 );
nand \U$33617 ( \33994 , \33992 , \33993 );
not \U$33618 ( \33995 , \33994 );
or \U$33619 ( \33996 , \33989 , \33995 );
not \U$33620 ( \33997 , RIc2265c0_35);
not \U$33621 ( \33998 , \30574 );
or \U$33622 ( \33999 , \33997 , \33998 );
nand \U$33623 ( \34000 , \9320 , \3620 );
nand \U$33624 ( \34001 , \33999 , \34000 );
nand \U$33625 ( \34002 , \34001 , \4381 );
nand \U$33626 ( \34003 , \33996 , \34002 );
not \U$33627 ( \34004 , \5509 );
not \U$33628 ( \34005 , RIc2264d0_37);
not \U$33629 ( \34006 , \10800 );
or \U$33630 ( \34007 , \34005 , \34006 );
nand \U$33631 ( \34008 , \9275 , \5514 );
nand \U$33632 ( \34009 , \34007 , \34008 );
not \U$33633 ( \34010 , \34009 );
or \U$33634 ( \34011 , \34004 , \34010 );
not \U$33635 ( \34012 , RIc2264d0_37);
not \U$33636 ( \34013 , \17015 );
or \U$33637 ( \34014 , \34012 , \34013 );
nand \U$33638 ( \34015 , \30878 , \5504 );
nand \U$33639 ( \34016 , \34014 , \34015 );
nand \U$33640 ( \34017 , \34016 , \5519 );
nand \U$33641 ( \34018 , \34011 , \34017 );
not \U$33642 ( \34019 , \34018 );
and \U$33643 ( \34020 , \34003 , \34019 );
not \U$33644 ( \34021 , \34003 );
and \U$33645 ( \34022 , \34021 , \34018 );
or \U$33646 ( \34023 , \34020 , \34022 );
xor \U$33647 ( \34024 , \33988 , \34023 );
not \U$33648 ( \34025 , \12304 );
not \U$33649 ( \34026 , RIc226020_47);
not \U$33650 ( \34027 , \12724 );
or \U$33651 ( \34028 , \34026 , \34027 );
not \U$33652 ( \34029 , \10322 );
nand \U$33653 ( \34030 , \34029 , \9373 );
nand \U$33654 ( \34031 , \34028 , \34030 );
not \U$33655 ( \34032 , \34031 );
or \U$33656 ( \34033 , \34025 , \34032 );
not \U$33657 ( \34034 , RIc226020_47);
not \U$33658 ( \34035 , \20217 );
or \U$33659 ( \34036 , \34034 , \34035 );
nand \U$33660 ( \34037 , \22969 , \9624 );
nand \U$33661 ( \34038 , \34036 , \34037 );
nand \U$33662 ( \34039 , \34038 , \10001 );
nand \U$33663 ( \34040 , \34033 , \34039 );
not \U$33664 ( \34041 , \9384 );
not \U$33665 ( \34042 , RIc226110_45);
not \U$33666 ( \34043 , \8953 );
or \U$33667 ( \34044 , \34042 , \34043 );
nand \U$33668 ( \34045 , \20368 , \14390 );
nand \U$33669 ( \34046 , \34044 , \34045 );
not \U$33670 ( \34047 , \34046 );
or \U$33671 ( \34048 , \34041 , \34047 );
not \U$33672 ( \34049 , RIc226110_45);
not \U$33673 ( \34050 , \8807 );
or \U$33674 ( \34051 , \34049 , \34050 );
nand \U$33675 ( \34052 , \10859 , \9100 );
nand \U$33676 ( \34053 , \34051 , \34052 );
nand \U$33677 ( \34054 , \34053 , \9398 );
nand \U$33678 ( \34055 , \34048 , \34054 );
xor \U$33679 ( \34056 , \34040 , \34055 );
not \U$33680 ( \34057 , \9552 );
not \U$33681 ( \34058 , RIc225f30_49);
not \U$33682 ( \34059 , \10609 );
or \U$33683 ( \34060 , \34058 , \34059 );
nand \U$33684 ( \34061 , \20646 , \9549 );
nand \U$33685 ( \34062 , \34060 , \34061 );
not \U$33686 ( \34063 , \34062 );
or \U$33687 ( \34064 , \34057 , \34063 );
not \U$33688 ( \34065 , \9533 );
not \U$33689 ( \34066 , RIc225f30_49);
not \U$33690 ( \34067 , \8887 );
or \U$33691 ( \34068 , \34066 , \34067 );
nand \U$33692 ( \34069 , \16532 , \9541 );
nand \U$33693 ( \34070 , \34068 , \34069 );
nand \U$33694 ( \34071 , \34065 , \34070 );
nand \U$33695 ( \34072 , \34064 , \34071 );
xnor \U$33696 ( \34073 , \34056 , \34072 );
xor \U$33697 ( \34074 , \34024 , \34073 );
not \U$33698 ( \34075 , \15729 );
not \U$33699 ( \34076 , RIc225990_61);
not \U$33700 ( \34077 , \14476 );
or \U$33701 ( \34078 , \34076 , \34077 );
nand \U$33702 ( \34079 , \9189 , \12806 );
nand \U$33703 ( \34080 , \34078 , \34079 );
not \U$33704 ( \34081 , \34080 );
or \U$33705 ( \34082 , \34075 , \34081 );
not \U$33706 ( \34083 , RIc225990_61);
not \U$33707 ( \34084 , \3715 );
or \U$33708 ( \34085 , \34083 , \34084 );
nand \U$33709 ( \34086 , \4501 , \10338 );
nand \U$33710 ( \34087 , \34085 , \34086 );
nand \U$33711 ( \34088 , \34087 , \15719 );
nand \U$33712 ( \34089 , \34082 , \34088 );
not \U$33713 ( \34090 , \34089 );
not \U$33714 ( \34091 , \34090 );
not \U$33715 ( \34092 , \8788 );
not \U$33716 ( \34093 , RIc225d50_53);
not \U$33717 ( \34094 , \20656 );
or \U$33718 ( \34095 , \34093 , \34094 );
nand \U$33719 ( \34096 , \6726 , \11585 );
nand \U$33720 ( \34097 , \34095 , \34096 );
not \U$33721 ( \34098 , \34097 );
or \U$33722 ( \34099 , \34092 , \34098 );
not \U$33723 ( \34100 , RIc225d50_53);
not \U$33724 ( \34101 , \10170 );
or \U$33725 ( \34102 , \34100 , \34101 );
nand \U$33726 ( \34103 , \23776 , \8782 );
nand \U$33727 ( \34104 , \34102 , \34103 );
nand \U$33728 ( \34105 , \34104 , \8777 );
nand \U$33729 ( \34106 , \34099 , \34105 );
not \U$33730 ( \34107 , \34106 );
not \U$33731 ( \34108 , \9444 );
not \U$33732 ( \34109 , RIc225e40_51);
not \U$33733 ( \34110 , \22928 );
or \U$33734 ( \34111 , \34109 , \34110 );
nand \U$33735 ( \34112 , \6494 , \12423 );
nand \U$33736 ( \34113 , \34111 , \34112 );
not \U$33737 ( \34114 , \34113 );
or \U$33738 ( \34115 , \34108 , \34114 );
not \U$33739 ( \34116 , RIc225e40_51);
not \U$33740 ( \34117 , \21438 );
or \U$33741 ( \34118 , \34116 , \34117 );
nand \U$33742 ( \34119 , \9740 , \22140 );
nand \U$33743 ( \34120 , \34118 , \34119 );
nand \U$33744 ( \34121 , \34120 , \9459 );
nand \U$33745 ( \34122 , \34115 , \34121 );
not \U$33746 ( \34123 , \34122 );
not \U$33747 ( \34124 , \34123 );
or \U$33748 ( \34125 , \34107 , \34124 );
or \U$33749 ( \34126 , \34123 , \34106 );
nand \U$33750 ( \34127 , \34125 , \34126 );
not \U$33751 ( \34128 , \34127 );
and \U$33752 ( \34129 , \34091 , \34128 );
and \U$33753 ( \34130 , \34090 , \34127 );
nor \U$33754 ( \34131 , \34129 , \34130 );
xor \U$33755 ( \34132 , \34074 , \34131 );
not \U$33756 ( \34133 , \34132 );
not \U$33757 ( \34134 , \6688 );
not \U$33758 ( \34135 , RIc2263e0_39);
not \U$33759 ( \34136 , \30875 );
or \U$33760 ( \34137 , \34135 , \34136 );
nand \U$33761 ( \34138 , \30878 , \8990 );
nand \U$33762 ( \34139 , \34137 , \34138 );
not \U$33763 ( \34140 , \34139 );
or \U$33764 ( \34141 , \34134 , \34140 );
not \U$33765 ( \34142 , RIc2263e0_39);
not \U$33766 ( \34143 , \10814 );
or \U$33767 ( \34144 , \34142 , \34143 );
nand \U$33768 ( \34145 , \10110 , \5498 );
nand \U$33769 ( \34146 , \34144 , \34145 );
nand \U$33770 ( \34147 , \34146 , \6307 );
nand \U$33771 ( \34148 , \34141 , \34147 );
not \U$33772 ( \34149 , \5519 );
not \U$33773 ( \34150 , \34009 );
or \U$33774 ( \34151 , \34149 , \34150 );
not \U$33775 ( \34152 , RIc2264d0_37);
not \U$33776 ( \34153 , \9300 );
or \U$33777 ( \34154 , \34152 , \34153 );
nand \U$33778 ( \34155 , \10266 , \5504 );
nand \U$33779 ( \34156 , \34154 , \34155 );
nand \U$33780 ( \34157 , \34156 , \5509 );
nand \U$33781 ( \34158 , \34151 , \34157 );
xor \U$33782 ( \34159 , \34148 , \34158 );
not \U$33783 ( \34160 , \5135 );
not \U$33784 ( \34161 , \34001 );
or \U$33785 ( \34162 , \34160 , \34161 );
not \U$33786 ( \34163 , RIc2265c0_35);
not \U$33787 ( \34164 , \31894 );
or \U$33788 ( \34165 , \34163 , \34164 );
not \U$33789 ( \34166 , \20610 );
nand \U$33790 ( \34167 , \34166 , \4376 );
nand \U$33791 ( \34168 , \34165 , \34167 );
nand \U$33792 ( \34169 , \34168 , \5741 );
nand \U$33793 ( \34170 , \34162 , \34169 );
xnor \U$33794 ( \34171 , \34159 , \34170 );
not \U$33795 ( \34172 , \34171 );
not \U$33796 ( \34173 , \9458 );
not \U$33797 ( \34174 , RIc225e40_51);
not \U$33798 ( \34175 , \8886 );
not \U$33799 ( \34176 , \34175 );
or \U$33800 ( \34177 , \34174 , \34176 );
nand \U$33801 ( \34178 , \17582 , \11795 );
nand \U$33802 ( \34179 , \34177 , \34178 );
not \U$33803 ( \34180 , \34179 );
or \U$33804 ( \34181 , \34173 , \34180 );
not \U$33805 ( \34182 , RIc225e40_51);
not \U$33806 ( \34183 , \10142 );
or \U$33807 ( \34184 , \34182 , \34183 );
nand \U$33808 ( \34185 , \20646 , \22140 );
nand \U$33809 ( \34186 , \34184 , \34185 );
nand \U$33810 ( \34187 , \34186 , \9444 );
nand \U$33811 ( \34188 , \34181 , \34187 );
not \U$33812 ( \34189 , \8777 );
not \U$33813 ( \34190 , RIc225d50_53);
not \U$33814 ( \34191 , \21438 );
or \U$33815 ( \34192 , \34190 , \34191 );
nand \U$33816 ( \34193 , \30634 , \11391 );
nand \U$33817 ( \34194 , \34192 , \34193 );
not \U$33818 ( \34195 , \34194 );
or \U$33819 ( \34196 , \34189 , \34195 );
not \U$33820 ( \34197 , RIc225d50_53);
not \U$33821 ( \34198 , \10125 );
or \U$33822 ( \34199 , \34197 , \34198 );
or \U$33823 ( \34200 , \22928 , RIc225d50_53);
nand \U$33824 ( \34201 , \34199 , \34200 );
nand \U$33825 ( \34202 , \34201 , \9555 );
nand \U$33826 ( \34203 , \34196 , \34202 );
xor \U$33827 ( \34204 , \34188 , \34203 );
not \U$33828 ( \34205 , \15719 );
not \U$33829 ( \34206 , RIc225990_61);
not \U$33830 ( \34207 , \3726 );
or \U$33831 ( \34208 , \34206 , \34207 );
nand \U$33832 ( \34209 , \2980 , \10338 );
nand \U$33833 ( \34210 , \34208 , \34209 );
not \U$33834 ( \34211 , \34210 );
or \U$33835 ( \34212 , \34205 , \34211 );
and \U$33836 ( \34213 , \3119 , RIc225990_61);
not \U$33837 ( \34214 , \3119 );
and \U$33838 ( \34215 , \34214 , \10338 );
or \U$33839 ( \34216 , \34213 , \34215 );
nand \U$33840 ( \34217 , \34216 , \20862 );
nand \U$33841 ( \34218 , \34212 , \34217 );
and \U$33842 ( \34219 , \34204 , \34218 );
and \U$33843 ( \34220 , \34188 , \34203 );
or \U$33844 ( \34221 , \34219 , \34220 );
not \U$33845 ( \34222 , \34221 );
not \U$33846 ( \34223 , \34222 );
or \U$33847 ( \34224 , \34172 , \34223 );
or \U$33848 ( \34225 , RIc226908_28, RIc226890_29);
nand \U$33849 ( \34226 , \34225 , \16248 );
and \U$33850 ( \34227 , RIc226908_28, RIc226890_29);
nor \U$33851 ( \34228 , \34227 , \2150 );
and \U$33852 ( \34229 , \34226 , \34228 );
not \U$33853 ( \34230 , \2153 );
not \U$33854 ( \34231 , RIc226980_27);
not \U$33855 ( \34232 , \30827 );
or \U$33856 ( \34233 , \34231 , \34232 );
nand \U$33857 ( \34234 , \16482 , \2150 );
nand \U$33858 ( \34235 , \34233 , \34234 );
not \U$33859 ( \34236 , \34235 );
or \U$33860 ( \34237 , \34230 , \34236 );
or \U$33861 ( \34238 , \16248 , \2799 );
or \U$33862 ( \34239 , \21954 , RIc226980_27);
nand \U$33863 ( \34240 , \34238 , \34239 );
nand \U$33864 ( \34241 , \34240 , \2137 );
nand \U$33865 ( \34242 , \34237 , \34241 );
xor \U$33866 ( \34243 , \34229 , \34242 );
not \U$33867 ( \34244 , \2086 );
and \U$33868 ( \34245 , RIc226890_29, \12846 );
not \U$33869 ( \34246 , RIc226890_29);
and \U$33870 ( \34247 , \34246 , \18161 );
or \U$33871 ( \34248 , \34245 , \34247 );
not \U$33872 ( \34249 , \34248 );
or \U$33873 ( \34250 , \34244 , \34249 );
and \U$33874 ( \34251 , RIc226890_29, \13488 );
not \U$33875 ( \34252 , RIc226890_29);
and \U$33876 ( \34253 , \34252 , \30679 );
nor \U$33877 ( \34254 , \34251 , \34253 );
nand \U$33878 ( \34255 , \34254 , \2078 );
nand \U$33879 ( \34256 , \34250 , \34255 );
xor \U$33880 ( \34257 , \34243 , \34256 );
not \U$33881 ( \34258 , \3630 );
not \U$33882 ( \34259 , RIc2266b0_33);
not \U$33883 ( \34260 , \10198 );
or \U$33884 ( \34261 , \34259 , \34260 );
nand \U$33885 ( \34262 , \20701 , \5179 );
nand \U$33886 ( \34263 , \34261 , \34262 );
not \U$33887 ( \34264 , \34263 );
or \U$33888 ( \34265 , \34258 , \34264 );
not \U$33889 ( \34266 , RIc2266b0_33);
not \U$33890 ( \34267 , \13498 );
or \U$33891 ( \34268 , \34266 , \34267 );
nand \U$33892 ( \34269 , \13497 , \5179 );
nand \U$33893 ( \34270 , \34268 , \34269 );
nand \U$33894 ( \34271 , \34270 , \3629 );
nand \U$33895 ( \34272 , \34265 , \34271 );
xor \U$33896 ( \34273 , \34257 , \34272 );
not \U$33897 ( \34274 , \11697 );
not \U$33898 ( \34275 , RIc225c60_55);
not \U$33899 ( \34276 , \22893 );
not \U$33900 ( \34277 , \34276 );
or \U$33901 ( \34278 , \34275 , \34277 );
nand \U$33902 ( \34279 , \6726 , \8767 );
nand \U$33903 ( \34280 , \34278 , \34279 );
not \U$33904 ( \34281 , \34280 );
or \U$33905 ( \34282 , \34274 , \34281 );
nand \U$33906 ( \34283 , \33986 , \11038 );
nand \U$33907 ( \34284 , \34282 , \34283 );
xor \U$33908 ( \34285 , \34273 , \34284 );
not \U$33909 ( \34286 , \9534 );
not \U$33910 ( \34287 , RIc225f30_49);
not \U$33911 ( \34288 , \20674 );
or \U$33912 ( \34289 , \34287 , \34288 );
nand \U$33913 ( \34290 , \31447 , \9541 );
nand \U$33914 ( \34291 , \34289 , \34290 );
not \U$33915 ( \34292 , \34291 );
or \U$33916 ( \34293 , \34286 , \34292 );
nand \U$33917 ( \34294 , \34070 , \9552 );
nand \U$33918 ( \34295 , \34293 , \34294 );
not \U$33919 ( \34296 , \34295 );
xnor \U$33920 ( \34297 , \34285 , \34296 );
nand \U$33921 ( \34298 , \34224 , \34297 );
not \U$33922 ( \34299 , \34171 );
nand \U$33923 ( \34300 , \34299 , \34221 );
and \U$33924 ( \34301 , \34298 , \34300 );
not \U$33925 ( \34302 , \34301 );
not \U$33926 ( \34303 , \34302 );
or \U$33927 ( \34304 , \34133 , \34303 );
not \U$33928 ( \34305 , \34301 );
not \U$33929 ( \34306 , \34132 );
not \U$33930 ( \34307 , \34306 );
or \U$33931 ( \34308 , \34305 , \34307 );
and \U$33932 ( \34309 , \18367 , \2172 );
not \U$33933 ( \34310 , \2153 );
not \U$33934 ( \34311 , RIc226980_27);
not \U$33935 ( \34312 , \15623 );
or \U$33936 ( \34313 , \34311 , \34312 );
nand \U$33937 ( \34314 , \20393 , \2133 );
nand \U$33938 ( \34315 , \34313 , \34314 );
not \U$33939 ( \34316 , \34315 );
or \U$33940 ( \34317 , \34310 , \34316 );
nand \U$33941 ( \34318 , \34235 , \2137 );
nand \U$33942 ( \34319 , \34317 , \34318 );
xor \U$33943 ( \34320 , \34309 , \34319 );
not \U$33944 ( \34321 , \2086 );
and \U$33945 ( \34322 , RIc226890_29, \30815 );
not \U$33946 ( \34323 , RIc226890_29);
and \U$33947 ( \34324 , \34323 , \19721 );
or \U$33948 ( \34325 , \34322 , \34324 );
not \U$33949 ( \34326 , \34325 );
or \U$33950 ( \34327 , \34321 , \34326 );
nand \U$33951 ( \34328 , \34248 , \2078 );
nand \U$33952 ( \34329 , \34327 , \34328 );
xor \U$33953 ( \34330 , \34320 , \34329 );
not \U$33954 ( \34331 , \6307 );
not \U$33955 ( \34332 , RIc2263e0_39);
not \U$33956 ( \34333 , \19789 );
or \U$33957 ( \34334 , \34332 , \34333 );
nand \U$33958 ( \34335 , \32612 , \5498 );
nand \U$33959 ( \34336 , \34334 , \34335 );
not \U$33960 ( \34337 , \34336 );
or \U$33961 ( \34338 , \34331 , \34337 );
nand \U$33962 ( \34339 , \6688 , \34146 );
nand \U$33963 ( \34340 , \34338 , \34339 );
xor \U$33964 ( \34341 , \34330 , \34340 );
not \U$33965 ( \34342 , \9705 );
not \U$33966 ( \34343 , RIc2262f0_41);
buf \U$33967 ( \34344 , \9215 );
not \U$33968 ( \34345 , \34344 );
or \U$33969 ( \34346 , \34343 , \34345 );
nand \U$33970 ( \34347 , \9211 , \6303 );
nand \U$33971 ( \34348 , \34346 , \34347 );
not \U$33972 ( \34349 , \34348 );
or \U$33973 ( \34350 , \34342 , \34349 );
not \U$33974 ( \34351 , RIc2262f0_41);
not \U$33975 ( \34352 , \9046 );
or \U$33976 ( \34353 , \34351 , \34352 );
nand \U$33977 ( \34354 , \9051 , \6303 );
nand \U$33978 ( \34355 , \34353 , \34354 );
nand \U$33979 ( \34356 , \34355 , \9690 );
nand \U$33980 ( \34357 , \34350 , \34356 );
xor \U$33981 ( \34358 , \34341 , \34357 );
not \U$33982 ( \34359 , \9129 );
not \U$33983 ( \34360 , RIc226200_43);
not \U$33984 ( \34361 , \8910 );
or \U$33985 ( \34362 , \34360 , \34361 );
not \U$33986 ( \34363 , \8910 );
nand \U$33987 ( \34364 , \34363 , \9117 );
nand \U$33988 ( \34365 , \34362 , \34364 );
not \U$33989 ( \34366 , \34365 );
or \U$33990 ( \34367 , \34359 , \34366 );
not \U$33991 ( \34368 , RIc226200_43);
not \U$33992 ( \34369 , \32810 );
or \U$33993 ( \34370 , \34368 , \34369 );
not \U$33994 ( \34371 , \34344 );
nand \U$33995 ( \34372 , \34371 , \9125 );
nand \U$33996 ( \34373 , \34370 , \34372 );
nand \U$33997 ( \34374 , \34373 , \9110 );
nand \U$33998 ( \34375 , \34367 , \34374 );
not \U$33999 ( \34376 , \9398 );
not \U$34000 ( \34377 , \34046 );
or \U$34001 ( \34378 , \34376 , \34377 );
not \U$34002 ( \34379 , RIc226110_45);
not \U$34003 ( \34380 , \11094 );
or \U$34004 ( \34381 , \34379 , \34380 );
nand \U$34005 ( \34382 , \21867 , \10429 );
nand \U$34006 ( \34383 , \34381 , \34382 );
nand \U$34007 ( \34384 , \34383 , \9934 );
nand \U$34008 ( \34385 , \34378 , \34384 );
nor \U$34009 ( \34386 , \34375 , \34385 );
not \U$34010 ( \34387 , \10953 );
not \U$34011 ( \34388 , \34038 );
or \U$34012 ( \34389 , \34387 , \34388 );
not \U$34013 ( \34390 , RIc226020_47);
not \U$34014 ( \34391 , \10295 );
or \U$34015 ( \34392 , \34390 , \34391 );
not \U$34016 ( \34393 , \8807 );
nand \U$34017 ( \34394 , \34393 , \9624 );
nand \U$34018 ( \34395 , \34392 , \34394 );
nand \U$34019 ( \34396 , \34395 , \9641 );
nand \U$34020 ( \34397 , \34389 , \34396 );
not \U$34021 ( \34398 , \34397 );
or \U$34022 ( \34399 , \34386 , \34398 );
nand \U$34023 ( \34400 , \34375 , \34385 );
nand \U$34024 ( \34401 , \34399 , \34400 );
xor \U$34025 ( \34402 , \34358 , \34401 );
or \U$34026 ( \34403 , RIc226818_30, RIc2267a0_31);
nand \U$34027 ( \34404 , \34403 , \16248 );
and \U$34028 ( \34405 , RIc226818_30, RIc2267a0_31);
nor \U$34029 ( \34406 , \34405 , \19846 );
and \U$34030 ( \34407 , \34404 , \34406 );
not \U$34031 ( \34408 , \2086 );
and \U$34032 ( \34409 , RIc226890_29, \20528 );
not \U$34033 ( \34410 , RIc226890_29);
and \U$34034 ( \34411 , \34410 , \32588 );
or \U$34035 ( \34412 , \34409 , \34411 );
not \U$34036 ( \34413 , \34412 );
or \U$34037 ( \34414 , \34408 , \34413 );
not \U$34038 ( \34415 , \2077 );
and \U$34039 ( \34416 , RIc226890_29, \16248 );
not \U$34040 ( \34417 , RIc226890_29);
and \U$34041 ( \34418 , \34417 , \18356 );
nor \U$34042 ( \34419 , \34416 , \34418 );
nand \U$34043 ( \34420 , \34415 , \34419 );
nand \U$34044 ( \34421 , \34414 , \34420 );
and \U$34045 ( \34422 , \34407 , \34421 );
not \U$34046 ( \34423 , \3629 );
not \U$34047 ( \34424 , RIc2266b0_33);
not \U$34048 ( \34425 , \20690 );
or \U$34049 ( \34426 , \34424 , \34425 );
nand \U$34050 ( \34427 , \12756 , \6890 );
nand \U$34051 ( \34428 , \34426 , \34427 );
not \U$34052 ( \34429 , \34428 );
or \U$34053 ( \34430 , \34423 , \34429 );
nand \U$34054 ( \34431 , \34270 , \3631 );
nand \U$34055 ( \34432 , \34430 , \34431 );
xor \U$34056 ( \34433 , \34422 , \34432 );
not \U$34057 ( \34434 , \4383 );
not \U$34058 ( \34435 , \34168 );
or \U$34059 ( \34436 , \34434 , \34435 );
not \U$34060 ( \34437 , RIc2265c0_35);
not \U$34061 ( \34438 , \13211 );
or \U$34062 ( \34439 , \34437 , \34438 );
nand \U$34063 ( \34440 , \32798 , \4376 );
nand \U$34064 ( \34441 , \34439 , \34440 );
nand \U$34065 ( \34442 , \34441 , \4381 );
nand \U$34066 ( \34443 , \34436 , \34442 );
and \U$34067 ( \34444 , \34433 , \34443 );
and \U$34068 ( \34445 , \34422 , \34432 );
or \U$34069 ( \34446 , \34444 , \34445 );
not \U$34070 ( \34447 , \15267 );
not \U$34071 ( \34448 , RIc225b70_57);
not \U$34072 ( \34449 , \21512 );
or \U$34073 ( \34450 , \34448 , \34449 );
nand \U$34074 ( \34451 , \16519 , \12475 );
nand \U$34075 ( \34452 , \34450 , \34451 );
not \U$34076 ( \34453 , \34452 );
or \U$34077 ( \34454 , \34447 , \34453 );
not \U$34078 ( \34455 , RIc225b70_57);
not \U$34079 ( \34456 , \10220 );
or \U$34080 ( \34457 , \34455 , \34456 );
nand \U$34081 ( \34458 , \4406 , \10074 );
nand \U$34082 ( \34459 , \34457 , \34458 );
nand \U$34083 ( \34460 , \34459 , \11965 );
nand \U$34084 ( \34461 , \34454 , \34460 );
xor \U$34085 ( \34462 , \34446 , \34461 );
not \U$34086 ( \34463 , \8788 );
not \U$34087 ( \34464 , \34104 );
or \U$34088 ( \34465 , \34463 , \34464 );
nand \U$34089 ( \34466 , \34201 , \9488 );
nand \U$34090 ( \34467 , \34465 , \34466 );
and \U$34091 ( \34468 , \34462 , \34467 );
and \U$34092 ( \34469 , \34446 , \34461 );
or \U$34093 ( \34470 , \34468 , \34469 );
xor \U$34094 ( \34471 , \34402 , \34470 );
nand \U$34095 ( \34472 , \34308 , \34471 );
nand \U$34096 ( \34473 , \34304 , \34472 );
not \U$34097 ( \34474 , \34024 );
nand \U$34098 ( \34475 , \34474 , \34131 );
not \U$34099 ( \34476 , \34073 );
and \U$34100 ( \34477 , \34475 , \34476 );
not \U$34101 ( \34478 , \34024 );
nor \U$34102 ( \34479 , \34478 , \34131 );
nor \U$34103 ( \34480 , \34477 , \34479 );
not \U$34104 ( \34481 , \34480 );
not \U$34105 ( \34482 , \34481 );
not \U$34106 ( \34483 , \34482 );
not \U$34107 ( \34484 , \34148 );
not \U$34108 ( \34485 , \34158 );
or \U$34109 ( \34486 , \34484 , \34485 );
or \U$34110 ( \34487 , \34148 , \34158 );
nand \U$34111 ( \34488 , \34487 , \34170 );
nand \U$34112 ( \34489 , \34486 , \34488 );
not \U$34113 ( \34490 , \34489 );
not \U$34114 ( \34491 , \34284 );
nand \U$34115 ( \34492 , \34491 , \34296 );
and \U$34116 ( \34493 , \34492 , \34273 );
and \U$34117 ( \34494 , \34295 , \34284 );
nor \U$34118 ( \34495 , \34493 , \34494 );
nand \U$34119 ( \34496 , \34490 , \34495 );
not \U$34120 ( \34497 , \34496 );
not \U$34121 ( \34498 , \2710 );
not \U$34122 ( \34499 , RIc2267a0_31);
not \U$34123 ( \34500 , \20690 );
or \U$34124 ( \34501 , \34499 , \34500 );
not \U$34125 ( \34502 , \16042 );
nand \U$34126 ( \34503 , \34502 , \2072 );
nand \U$34127 ( \34504 , \34501 , \34503 );
not \U$34128 ( \34505 , \34504 );
or \U$34129 ( \34506 , \34498 , \34505 );
not \U$34130 ( \34507 , RIc2267a0_31);
not \U$34131 ( \34508 , \15444 );
or \U$34132 ( \34509 , \34507 , \34508 );
nand \U$34133 ( \34510 , \15443 , \3648 );
nand \U$34134 ( \34511 , \34509 , \34510 );
nand \U$34135 ( \34512 , \34511 , \2697 );
nand \U$34136 ( \34513 , \34506 , \34512 );
and \U$34137 ( \34514 , \18357 , \2153 );
not \U$34138 ( \34515 , \2086 );
not \U$34139 ( \34516 , \34254 );
or \U$34140 ( \34517 , \34515 , \34516 );
nand \U$34141 ( \34518 , \34412 , \2078 );
nand \U$34142 ( \34519 , \34517 , \34518 );
xor \U$34143 ( \34520 , \34514 , \34519 );
not \U$34144 ( \34521 , \2697 );
not \U$34145 ( \34522 , RIc2267a0_31);
not \U$34146 ( \34523 , \18161 );
not \U$34147 ( \34524 , \34523 );
or \U$34148 ( \34525 , \34522 , \34524 );
nand \U$34149 ( \34526 , \12845 , \2705 );
nand \U$34150 ( \34527 , \34525 , \34526 );
not \U$34151 ( \34528 , \34527 );
or \U$34152 ( \34529 , \34521 , \34528 );
nand \U$34153 ( \34530 , \34511 , \2710 );
nand \U$34154 ( \34531 , \34529 , \34530 );
and \U$34155 ( \34532 , \34520 , \34531 );
and \U$34156 ( \34533 , \34514 , \34519 );
or \U$34157 ( \34534 , \34532 , \34533 );
xor \U$34158 ( \34535 , \34513 , \34534 );
not \U$34159 ( \34536 , \9705 );
not \U$34160 ( \34537 , \34355 );
or \U$34161 ( \34538 , \34536 , \34537 );
not \U$34162 ( \34539 , RIc2262f0_41);
not \U$34163 ( \34540 , \11394 );
or \U$34164 ( \34541 , \34539 , \34540 );
nand \U$34165 ( \34542 , \10653 , \6303 );
nand \U$34166 ( \34543 , \34541 , \34542 );
nand \U$34167 ( \34544 , \34543 , \9690 );
nand \U$34168 ( \34545 , \34538 , \34544 );
and \U$34169 ( \34546 , \34535 , \34545 );
and \U$34170 ( \34547 , \34513 , \34534 );
or \U$34171 ( \34548 , \34546 , \34547 );
not \U$34172 ( \34549 , \34548 );
or \U$34173 ( \34550 , \34497 , \34549 );
not \U$34174 ( \34551 , \34495 );
nand \U$34175 ( \34552 , \34551 , \34489 );
nand \U$34176 ( \34553 , \34550 , \34552 );
xor \U$34177 ( \34554 , \34358 , \34401 );
and \U$34178 ( \34555 , \34554 , \34470 );
and \U$34179 ( \34556 , \34358 , \34401 );
or \U$34180 ( \34557 , \34555 , \34556 );
xor \U$34181 ( \34558 , \34553 , \34557 );
not \U$34182 ( \34559 , \34558 );
or \U$34183 ( \34560 , \34483 , \34559 );
or \U$34184 ( \34561 , \34558 , \34482 );
nand \U$34185 ( \34562 , \34560 , \34561 );
xor \U$34186 ( \34563 , \34473 , \34562 );
xor \U$34187 ( \34564 , \34330 , \34340 );
and \U$34188 ( \34565 , \34564 , \34357 );
and \U$34189 ( \34566 , \34330 , \34340 );
or \U$34190 ( \34567 , \34565 , \34566 );
not \U$34191 ( \34568 , \34003 );
nand \U$34192 ( \34569 , \34568 , \34019 );
not \U$34193 ( \34570 , \34569 );
not \U$34194 ( \34571 , \33988 );
or \U$34195 ( \34572 , \34570 , \34571 );
nand \U$34196 ( \34573 , \34018 , \34003 );
nand \U$34197 ( \34574 , \34572 , \34573 );
xor \U$34198 ( \34575 , \34567 , \34574 );
not \U$34199 ( \34576 , \3631 );
not \U$34200 ( \34577 , RIc2266b0_33);
not \U$34201 ( \34578 , \9321 );
or \U$34202 ( \34579 , \34577 , \34578 );
nand \U$34203 ( \34580 , \9320 , \9943 );
nand \U$34204 ( \34581 , \34579 , \34580 );
not \U$34205 ( \34582 , \34581 );
or \U$34206 ( \34583 , \34576 , \34582 );
and \U$34207 ( \34584 , RIc2266b0_33, \10086 );
not \U$34208 ( \34585 , RIc2266b0_33);
and \U$34209 ( \34586 , \34585 , \21172 );
nor \U$34210 ( \34587 , \34584 , \34586 );
nand \U$34211 ( \34588 , \34587 , \3629 );
nand \U$34212 ( \34589 , \34583 , \34588 );
not \U$34213 ( \34590 , \5509 );
not \U$34214 ( \34591 , \34016 );
or \U$34215 ( \34592 , \34590 , \34591 );
not \U$34216 ( \34593 , RIc2264d0_37);
not \U$34217 ( \34594 , \10814 );
or \U$34218 ( \34595 , \34593 , \34594 );
nand \U$34219 ( \34596 , \10110 , \5514 );
nand \U$34220 ( \34597 , \34595 , \34596 );
nand \U$34221 ( \34598 , \34597 , \5519 );
nand \U$34222 ( \34599 , \34592 , \34598 );
xor \U$34223 ( \34600 , \34589 , \34599 );
not \U$34224 ( \34601 , \4383 );
not \U$34225 ( \34602 , RIc2265c0_35);
not \U$34226 ( \34603 , \21156 );
or \U$34227 ( \34604 , \34602 , \34603 );
nand \U$34228 ( \34605 , \10976 , \4376 );
nand \U$34229 ( \34606 , \34604 , \34605 );
not \U$34230 ( \34607 , \34606 );
or \U$34231 ( \34608 , \34601 , \34607 );
nand \U$34232 ( \34609 , \33994 , \4381 );
nand \U$34233 ( \34610 , \34608 , \34609 );
xor \U$34234 ( \34611 , \34600 , \34610 );
xor \U$34235 ( \34612 , \34575 , \34611 );
not \U$34236 ( \34613 , \9816 );
not \U$34237 ( \34614 , RIc2262f0_41);
not \U$34238 ( \34615 , \8910 );
or \U$34239 ( \34616 , \34614 , \34615 );
not \U$34240 ( \34617 , \12403 );
nand \U$34241 ( \34618 , \34617 , \6303 );
nand \U$34242 ( \34619 , \34616 , \34618 );
not \U$34243 ( \34620 , \34619 );
or \U$34244 ( \34621 , \34613 , \34620 );
nand \U$34245 ( \34622 , \34348 , \9690 );
nand \U$34246 ( \34623 , \34621 , \34622 );
not \U$34247 ( \34624 , \11708 );
not \U$34248 ( \34625 , RIc225e40_51);
not \U$34249 ( \34626 , \10170 );
or \U$34250 ( \34627 , \34625 , \34626 );
not \U$34251 ( \34628 , \25704 );
nand \U$34252 ( \34629 , \34628 , \22140 );
nand \U$34253 ( \34630 , \34627 , \34629 );
not \U$34254 ( \34631 , \34630 );
or \U$34255 ( \34632 , \34624 , \34631 );
nand \U$34256 ( \34633 , \34113 , \9459 );
nand \U$34257 ( \34634 , \34632 , \34633 );
xor \U$34258 ( \34635 , \34623 , \34634 );
not \U$34259 ( \34636 , \8788 );
not \U$34260 ( \34637 , RIc225d50_53);
not \U$34261 ( \34638 , \10230 );
or \U$34262 ( \34639 , \34637 , \34638 );
not \U$34263 ( \34640 , \30619 );
nand \U$34264 ( \34641 , \34640 , \8782 );
nand \U$34265 ( \34642 , \34639 , \34641 );
not \U$34266 ( \34643 , \34642 );
or \U$34267 ( \34644 , \34636 , \34643 );
nand \U$34268 ( \34645 , \34097 , \9488 );
nand \U$34269 ( \34646 , \34644 , \34645 );
xor \U$34270 ( \34647 , \34635 , \34646 );
not \U$34271 ( \34648 , \34647 );
not \U$34272 ( \34649 , \34648 );
not \U$34273 ( \34650 , \34040 );
not \U$34274 ( \34651 , \34055 );
or \U$34275 ( \34652 , \34650 , \34651 );
or \U$34276 ( \34653 , \34055 , \34040 );
nand \U$34277 ( \34654 , \34653 , \34072 );
nand \U$34278 ( \34655 , \34652 , \34654 );
not \U$34279 ( \34656 , \11974 );
not \U$34280 ( \34657 , RIc225b70_57);
not \U$34281 ( \34658 , \4046 );
or \U$34282 ( \34659 , \34657 , \34658 );
nand \U$34283 ( \34660 , \15768 , \12475 );
nand \U$34284 ( \34661 , \34659 , \34660 );
not \U$34285 ( \34662 , \34661 );
or \U$34286 ( \34663 , \34656 , \34662 );
nand \U$34287 ( \34664 , \34452 , \11965 );
nand \U$34288 ( \34665 , \34663 , \34664 );
not \U$34289 ( \34666 , \9110 );
not \U$34290 ( \34667 , \34365 );
or \U$34291 ( \34668 , \34666 , \34667 );
not \U$34292 ( \34669 , RIc226200_43);
not \U$34293 ( \34670 , \21866 );
or \U$34294 ( \34671 , \34669 , \34670 );
nand \U$34295 ( \34672 , \21867 , \9106 );
nand \U$34296 ( \34673 , \34671 , \34672 );
nand \U$34297 ( \34674 , \34673 , \9205 );
nand \U$34298 ( \34675 , \34668 , \34674 );
or \U$34299 ( \34676 , \34665 , \34675 );
xor \U$34300 ( \34677 , \34243 , \34256 );
and \U$34301 ( \34678 , \34677 , \34272 );
and \U$34302 ( \34679 , \34243 , \34256 );
or \U$34303 ( \34680 , \34678 , \34679 );
nand \U$34304 ( \34681 , \34676 , \34680 );
nand \U$34305 ( \34682 , \34665 , \34675 );
nand \U$34306 ( \34683 , \34681 , \34682 );
xor \U$34307 ( \34684 , \34655 , \34683 );
not \U$34308 ( \34685 , \34684 );
or \U$34309 ( \34686 , \34649 , \34685 );
or \U$34310 ( \34687 , \34684 , \34648 );
nand \U$34311 ( \34688 , \34686 , \34687 );
xor \U$34312 ( \34689 , \34612 , \34688 );
xor \U$34313 ( \34690 , \32772 , \32780 );
not \U$34314 ( \34691 , \2154 );
not \U$34315 ( \34692 , \32599 );
or \U$34316 ( \34693 , \34691 , \34692 );
nand \U$34317 ( \34694 , \34315 , \2138 );
nand \U$34318 ( \34695 , \34693 , \34694 );
xor \U$34319 ( \34696 , \34690 , \34695 );
not \U$34320 ( \34697 , \2086 );
not \U$34321 ( \34698 , \32786 );
or \U$34322 ( \34699 , \34697 , \34698 );
nand \U$34323 ( \34700 , \34325 , \2078 );
nand \U$34324 ( \34701 , \34699 , \34700 );
xor \U$34325 ( \34702 , \34696 , \34701 );
not \U$34326 ( \34703 , \9532 );
not \U$34327 ( \34704 , \34062 );
or \U$34328 ( \34705 , \34703 , \34704 );
not \U$34329 ( \34706 , RIc225f30_49);
not \U$34330 ( \34707 , \6719 );
or \U$34331 ( \34708 , \34706 , \34707 );
not \U$34332 ( \34709 , \21438 );
nand \U$34333 ( \34710 , \34709 , \11289 );
nand \U$34334 ( \34711 , \34708 , \34710 );
nand \U$34335 ( \34712 , \34711 , \9552 );
nand \U$34336 ( \34713 , \34705 , \34712 );
xor \U$34337 ( \34714 , \34702 , \34713 );
not \U$34338 ( \34715 , \10001 );
not \U$34339 ( \34716 , \34031 );
or \U$34340 ( \34717 , \34715 , \34716 );
and \U$34341 ( \34718 , \11607 , \17582 );
not \U$34342 ( \34719 , \11607 );
and \U$34343 ( \34720 , \34719 , \8887 );
nor \U$34344 ( \34721 , \34718 , \34720 );
not \U$34345 ( \34722 , \34721 );
nand \U$34346 ( \34723 , \34722 , \9619 );
nand \U$34347 ( \34724 , \34717 , \34723 );
xor \U$34348 ( \34725 , \34714 , \34724 );
not \U$34349 ( \34726 , \34122 );
not \U$34350 ( \34727 , \34089 );
or \U$34351 ( \34728 , \34726 , \34727 );
or \U$34352 ( \34729 , \34089 , \34122 );
nand \U$34353 ( \34730 , \34729 , \34106 );
nand \U$34354 ( \34731 , \34728 , \34730 );
xor \U$34355 ( \34732 , \34725 , \34731 );
not \U$34356 ( \34733 , \15164 );
and \U$34357 ( \34734 , RIc225a80_59, \6439 );
not \U$34358 ( \34735 , RIc225a80_59);
and \U$34359 ( \34736 , \34735 , \2981 );
or \U$34360 ( \34737 , \34734 , \34736 );
not \U$34361 ( \34738 , \34737 );
or \U$34362 ( \34739 , \34733 , \34738 );
and \U$34363 ( \34740 , RIc225a80_59, \3121 );
not \U$34364 ( \34741 , RIc225a80_59);
and \U$34365 ( \34742 , \34741 , \5160 );
or \U$34366 ( \34743 , \34740 , \34742 );
nand \U$34367 ( \34744 , \34743 , \18037 );
nand \U$34368 ( \34745 , \34739 , \34744 );
not \U$34369 ( \34746 , \34745 );
not \U$34370 ( \34747 , RIc225828_64);
not \U$34371 ( \34748 , RIc2258a0_63);
not \U$34372 ( \34749 , \3010 );
or \U$34373 ( \34750 , \34748 , \34749 );
nand \U$34374 ( \34751 , \23331 , \16880 );
nand \U$34375 ( \34752 , \34750 , \34751 );
not \U$34376 ( \34753 , \34752 );
or \U$34377 ( \34754 , \34747 , \34753 );
not \U$34378 ( \34755 , RIc2258a0_63);
not \U$34379 ( \34756 , \3799 );
or \U$34380 ( \34757 , \34755 , \34756 );
nand \U$34381 ( \34758 , \2044 , \15620 );
nand \U$34382 ( \34759 , \34757 , \34758 );
nand \U$34383 ( \34760 , \34759 , \20159 );
nand \U$34384 ( \34761 , \34754 , \34760 );
not \U$34385 ( \34762 , \34761 );
or \U$34386 ( \34763 , \34746 , \34762 );
or \U$34387 ( \34764 , \34761 , \34745 );
and \U$34388 ( \34765 , \34229 , \34242 );
not \U$34389 ( \34766 , \2710 );
not \U$34390 ( \34767 , RIc2267a0_31);
not \U$34391 ( \34768 , \13498 );
or \U$34392 ( \34769 , \34767 , \34768 );
nand \U$34393 ( \34770 , \20406 , \3648 );
nand \U$34394 ( \34771 , \34769 , \34770 );
not \U$34395 ( \34772 , \34771 );
or \U$34396 ( \34773 , \34766 , \34772 );
nand \U$34397 ( \34774 , \34504 , \2697 );
nand \U$34398 ( \34775 , \34773 , \34774 );
xor \U$34399 ( \34776 , \34765 , \34775 );
not \U$34400 ( \34777 , \3631 );
not \U$34401 ( \34778 , \34587 );
or \U$34402 ( \34779 , \34777 , \34778 );
nand \U$34403 ( \34780 , \34263 , \3629 );
nand \U$34404 ( \34781 , \34779 , \34780 );
xor \U$34405 ( \34782 , \34776 , \34781 );
nand \U$34406 ( \34783 , \34764 , \34782 );
nand \U$34407 ( \34784 , \34763 , \34783 );
xor \U$34408 ( \34785 , \34732 , \34784 );
xor \U$34409 ( \34786 , \34689 , \34785 );
xor \U$34410 ( \34787 , \34563 , \34786 );
xor \U$34411 ( \34788 , \34171 , \34297 );
xnor \U$34412 ( \34789 , \34788 , \34221 );
xor \U$34413 ( \34790 , \34407 , \34421 );
not \U$34414 ( \34791 , \2710 );
not \U$34415 ( \34792 , \34527 );
or \U$34416 ( \34793 , \34791 , \34792 );
not \U$34417 ( \34794 , RIc2267a0_31);
not \U$34418 ( \34795 , \21094 );
or \U$34419 ( \34796 , \34794 , \34795 );
nand \U$34420 ( \34797 , \13488 , \2072 );
nand \U$34421 ( \34798 , \34796 , \34797 );
nand \U$34422 ( \34799 , \34798 , \2697 );
nand \U$34423 ( \34800 , \34793 , \34799 );
xor \U$34424 ( \34801 , \34790 , \34800 );
not \U$34425 ( \34802 , \5135 );
not \U$34426 ( \34803 , \34441 );
or \U$34427 ( \34804 , \34802 , \34803 );
not \U$34428 ( \34805 , RIc2265c0_35);
not \U$34429 ( \34806 , \16492 );
or \U$34430 ( \34807 , \34805 , \34806 );
nand \U$34431 ( \34808 , \10356 , \3620 );
nand \U$34432 ( \34809 , \34807 , \34808 );
nand \U$34433 ( \34810 , \34809 , \4380 );
nand \U$34434 ( \34811 , \34804 , \34810 );
and \U$34435 ( \34812 , \34801 , \34811 );
and \U$34436 ( \34813 , \34790 , \34800 );
or \U$34437 ( \34814 , \34812 , \34813 );
not \U$34438 ( \34815 , \12532 );
not \U$34439 ( \34816 , \34280 );
or \U$34440 ( \34817 , \34815 , \34816 );
not \U$34441 ( \34818 , RIc225c60_55);
not \U$34442 ( \34819 , \10170 );
or \U$34443 ( \34820 , \34818 , \34819 );
not \U$34444 ( \34821 , \17549 );
nand \U$34445 ( \34822 , \34821 , \11108 );
nand \U$34446 ( \34823 , \34820 , \34822 );
nand \U$34447 ( \34824 , \34823 , \11117 );
nand \U$34448 ( \34825 , \34817 , \34824 );
xor \U$34449 ( \34826 , \34814 , \34825 );
not \U$34450 ( \34827 , \15183 );
not \U$34451 ( \34828 , \34383 );
or \U$34452 ( \34829 , \34827 , \34828 );
not \U$34453 ( \34830 , RIc226110_45);
not \U$34454 ( \34831 , \8910 );
or \U$34455 ( \34832 , \34830 , \34831 );
nand \U$34456 ( \34833 , \9790 , \14660 );
nand \U$34457 ( \34834 , \34832 , \34833 );
nand \U$34458 ( \34835 , \34834 , \9934 );
nand \U$34459 ( \34836 , \34829 , \34835 );
xor \U$34460 ( \34837 , \34826 , \34836 );
xor \U$34461 ( \34838 , \34422 , \34432 );
xor \U$34462 ( \34839 , \34838 , \34443 );
not \U$34463 ( \34840 , \3631 );
not \U$34464 ( \34841 , \34428 );
or \U$34465 ( \34842 , \34840 , \34841 );
not \U$34466 ( \34843 , RIc2266b0_33);
not \U$34467 ( \34844 , \30815 );
or \U$34468 ( \34845 , \34843 , \34844 );
nand \U$34469 ( \34846 , \19721 , \16360 );
nand \U$34470 ( \34847 , \34845 , \34846 );
nand \U$34471 ( \34848 , \34847 , \3629 );
nand \U$34472 ( \34849 , \34842 , \34848 );
and \U$34473 ( \34850 , \16248 , \2086 );
not \U$34474 ( \34851 , \2710 );
not \U$34475 ( \34852 , \34798 );
or \U$34476 ( \34853 , \34851 , \34852 );
not \U$34477 ( \34854 , RIc2267a0_31);
not \U$34478 ( \34855 , \21102 );
or \U$34479 ( \34856 , \34854 , \34855 );
nand \U$34480 ( \34857 , \16482 , \2072 );
nand \U$34481 ( \34858 , \34856 , \34857 );
nand \U$34482 ( \34859 , \34858 , \2696 );
nand \U$34483 ( \34860 , \34853 , \34859 );
xor \U$34484 ( \34861 , \34850 , \34860 );
not \U$34485 ( \34862 , \3630 );
not \U$34486 ( \34863 , \34847 );
or \U$34487 ( \34864 , \34862 , \34863 );
not \U$34488 ( \34865 , RIc2266b0_33);
not \U$34489 ( \34866 , \18158 );
or \U$34490 ( \34867 , \34865 , \34866 );
nand \U$34491 ( \34868 , \18161 , \2692 );
nand \U$34492 ( \34869 , \34867 , \34868 );
nand \U$34493 ( \34870 , \34869 , \3629 );
nand \U$34494 ( \34871 , \34864 , \34870 );
and \U$34495 ( \34872 , \34861 , \34871 );
and \U$34496 ( \34873 , \34850 , \34860 );
or \U$34497 ( \34874 , \34872 , \34873 );
xor \U$34498 ( \34875 , \34849 , \34874 );
not \U$34499 ( \34876 , \9129 );
not \U$34500 ( \34877 , RIc226200_43);
not \U$34501 ( \34878 , \13465 );
or \U$34502 ( \34879 , \34877 , \34878 );
nand \U$34503 ( \34880 , \9051 , \9117 );
nand \U$34504 ( \34881 , \34879 , \34880 );
not \U$34505 ( \34882 , \34881 );
or \U$34506 ( \34883 , \34876 , \34882 );
not \U$34507 ( \34884 , RIc226200_43);
not \U$34508 ( \34885 , \19789 );
or \U$34509 ( \34886 , \34884 , \34885 );
nand \U$34510 ( \34887 , \32612 , \9117 );
nand \U$34511 ( \34888 , \34886 , \34887 );
nand \U$34512 ( \34889 , \34888 , \9110 );
nand \U$34513 ( \34890 , \34883 , \34889 );
and \U$34514 ( \34891 , \34875 , \34890 );
and \U$34515 ( \34892 , \34849 , \34874 );
or \U$34516 ( \34893 , \34891 , \34892 );
xor \U$34517 ( \34894 , \34839 , \34893 );
not \U$34518 ( \34895 , \20159 );
not \U$34519 ( \34896 , RIc2258a0_63);
not \U$34520 ( \34897 , \2104 );
or \U$34521 ( \34898 , \34896 , \34897 );
nand \U$34522 ( \34899 , \9654 , \16880 );
nand \U$34523 ( \34900 , \34898 , \34899 );
not \U$34524 ( \34901 , \34900 );
or \U$34525 ( \34902 , \34895 , \34901 );
not \U$34526 ( \34903 , RIc2258a0_63);
not \U$34527 ( \34904 , \4228 );
or \U$34528 ( \34905 , \34903 , \34904 );
nand \U$34529 ( \34906 , \13251 , \16880 );
nand \U$34530 ( \34907 , \34905 , \34906 );
nand \U$34531 ( \34908 , \34907 , RIc225828_64);
nand \U$34532 ( \34909 , \34902 , \34908 );
xor \U$34533 ( \34910 , \34894 , \34909 );
xor \U$34534 ( \34911 , \34837 , \34910 );
xor \U$34535 ( \34912 , \34849 , \34874 );
xor \U$34536 ( \34913 , \34912 , \34890 );
not \U$34537 ( \34914 , \6688 );
not \U$34538 ( \34915 , RIc2263e0_39);
not \U$34539 ( \34916 , \30574 );
or \U$34540 ( \34917 , \34915 , \34916 );
nand \U$34541 ( \34918 , \9324 , \8990 );
nand \U$34542 ( \34919 , \34917 , \34918 );
not \U$34543 ( \34920 , \34919 );
or \U$34544 ( \34921 , \34914 , \34920 );
not \U$34545 ( \34922 , RIc2263e0_39);
not \U$34546 ( \34923 , \9297 );
or \U$34547 ( \34924 , \34922 , \34923 );
nand \U$34548 ( \34925 , \10266 , \5498 );
nand \U$34549 ( \34926 , \34924 , \34925 );
nand \U$34550 ( \34927 , \34926 , \6307 );
nand \U$34551 ( \34928 , \34921 , \34927 );
not \U$34552 ( \34929 , \34928 );
not \U$34553 ( \34930 , \9110 );
not \U$34554 ( \34931 , RIc226200_43);
not \U$34555 ( \34932 , \10814 );
or \U$34556 ( \34933 , \34931 , \34932 );
nand \U$34557 ( \34934 , \10110 , \9117 );
nand \U$34558 ( \34935 , \34933 , \34934 );
not \U$34559 ( \34936 , \34935 );
or \U$34560 ( \34937 , \34930 , \34936 );
nand \U$34561 ( \34938 , \34888 , \9205 );
nand \U$34562 ( \34939 , \34937 , \34938 );
not \U$34563 ( \34940 , \34939 );
or \U$34564 ( \34941 , \34929 , \34940 );
or \U$34565 ( \34942 , \34939 , \34928 );
xor \U$34566 ( \34943 , \34850 , \34860 );
xor \U$34567 ( \34944 , \34943 , \34871 );
nand \U$34568 ( \34945 , \34942 , \34944 );
nand \U$34569 ( \34946 , \34941 , \34945 );
xor \U$34570 ( \34947 , \34913 , \34946 );
or \U$34571 ( \34948 , RIc226728_32, RIc2266b0_33);
nand \U$34572 ( \34949 , \34948 , \18357 );
and \U$34573 ( \34950 , RIc226728_32, RIc2266b0_33);
nor \U$34574 ( \34951 , \34950 , \2072 );
and \U$34575 ( \34952 , \34949 , \34951 );
not \U$34576 ( \34953 , \2710 );
not \U$34577 ( \34954 , \34858 );
or \U$34578 ( \34955 , \34953 , \34954 );
or \U$34579 ( \34956 , \18357 , \3648 );
or \U$34580 ( \34957 , \18356 , RIc2267a0_31);
nand \U$34581 ( \34958 , \34956 , \34957 );
nand \U$34582 ( \34959 , \34958 , \2696 );
nand \U$34583 ( \34960 , \34955 , \34959 );
xor \U$34584 ( \34961 , \34952 , \34960 );
not \U$34585 ( \34962 , \3630 );
not \U$34586 ( \34963 , \34869 );
or \U$34587 ( \34964 , \34962 , \34963 );
not \U$34588 ( \34965 , RIc2266b0_33);
not \U$34589 ( \34966 , \15623 );
or \U$34590 ( \34967 , \34965 , \34966 );
nand \U$34591 ( \34968 , \20393 , \5179 );
nand \U$34592 ( \34969 , \34967 , \34968 );
nand \U$34593 ( \34970 , \34969 , \3629 );
nand \U$34594 ( \34971 , \34964 , \34970 );
xor \U$34595 ( \34972 , \34961 , \34971 );
not \U$34596 ( \34973 , \5519 );
not \U$34597 ( \34974 , \5504 );
not \U$34598 ( \34975 , \20701 );
or \U$34599 ( \34976 , \34974 , \34975 );
not \U$34600 ( \34977 , \10370 );
nand \U$34601 ( \34978 , \34977 , RIc2264d0_37);
nand \U$34602 ( \34979 , \34976 , \34978 );
not \U$34603 ( \34980 , \34979 );
or \U$34604 ( \34981 , \34973 , \34980 );
not \U$34605 ( \34982 , RIc2264d0_37);
not \U$34606 ( \34983 , \17625 );
or \U$34607 ( \34984 , \34982 , \34983 );
nand \U$34608 ( \34985 , \13497 , \5504 );
nand \U$34609 ( \34986 , \34984 , \34985 );
nand \U$34610 ( \34987 , \34986 , \5509 );
nand \U$34611 ( \34988 , \34981 , \34987 );
and \U$34612 ( \34989 , \34972 , \34988 );
and \U$34613 ( \34990 , \34961 , \34971 );
or \U$34614 ( \34991 , \34989 , \34990 );
not \U$34615 ( \34992 , \11965 );
not \U$34616 ( \34993 , RIc225b70_57);
not \U$34617 ( \34994 , \9765 );
or \U$34618 ( \34995 , \34993 , \34994 );
nand \U$34619 ( \34996 , \9770 , \10074 );
nand \U$34620 ( \34997 , \34995 , \34996 );
not \U$34621 ( \34998 , \34997 );
or \U$34622 ( \34999 , \34992 , \34998 );
not \U$34623 ( \35000 , RIc225b70_57);
not \U$34624 ( \35001 , \5664 );
or \U$34625 ( \35002 , \35000 , \35001 );
nand \U$34626 ( \35003 , \5663 , \10074 );
nand \U$34627 ( \35004 , \35002 , \35003 );
nand \U$34628 ( \35005 , \35004 , \11974 );
nand \U$34629 ( \35006 , \34999 , \35005 );
xor \U$34630 ( \35007 , \34991 , \35006 );
not \U$34631 ( \35008 , \9488 );
not \U$34632 ( \35009 , RIc225d50_53);
not \U$34633 ( \35010 , \34175 );
or \U$34634 ( \35011 , \35009 , \35010 );
nand \U$34635 ( \35012 , \16532 , \8772 );
nand \U$34636 ( \35013 , \35011 , \35012 );
not \U$34637 ( \35014 , \35013 );
or \U$34638 ( \35015 , \35008 , \35014 );
not \U$34639 ( \35016 , RIc225d50_53);
not \U$34640 ( \35017 , \10307 );
or \U$34641 ( \35018 , \35016 , \35017 );
nand \U$34642 ( \35019 , \10141 , \8782 );
nand \U$34643 ( \35020 , \35018 , \35019 );
nand \U$34644 ( \35021 , \35020 , \8788 );
nand \U$34645 ( \35022 , \35015 , \35021 );
and \U$34646 ( \35023 , \35007 , \35022 );
and \U$34647 ( \35024 , \34991 , \35006 );
or \U$34648 ( \35025 , \35023 , \35024 );
and \U$34649 ( \35026 , \34947 , \35025 );
and \U$34650 ( \35027 , \34913 , \34946 );
or \U$34651 ( \35028 , \35026 , \35027 );
and \U$34652 ( \35029 , \34911 , \35028 );
and \U$34653 ( \35030 , \34837 , \34910 );
or \U$34654 ( \35031 , \35029 , \35030 );
xor \U$34655 ( \35032 , \34789 , \35031 );
xor \U$34656 ( \35033 , \34446 , \34461 );
xor \U$34657 ( \35034 , \35033 , \34467 );
xor \U$34658 ( \35035 , \34375 , \34398 );
xor \U$34659 ( \35036 , \35035 , \34385 );
and \U$34660 ( \35037 , \35034 , \35036 );
not \U$34661 ( \35038 , \35034 );
not \U$34662 ( \35039 , \35036 );
and \U$34663 ( \35040 , \35038 , \35039 );
or \U$34664 ( \35041 , \35037 , \35040 );
not \U$34665 ( \35042 , \9444 );
not \U$34666 ( \35043 , \34120 );
or \U$34667 ( \35044 , \35042 , \35043 );
nand \U$34668 ( \35045 , \34186 , \9459 );
nand \U$34669 ( \35046 , \35044 , \35045 );
not \U$34670 ( \35047 , \20862 );
not \U$34671 ( \35048 , \34087 );
or \U$34672 ( \35049 , \35047 , \35048 );
nand \U$34673 ( \35050 , \34216 , \15719 );
nand \U$34674 ( \35051 , \35049 , \35050 );
xor \U$34675 ( \35052 , \35046 , \35051 );
not \U$34676 ( \35053 , \20159 );
not \U$34677 ( \35054 , \34907 );
or \U$34678 ( \35055 , \35053 , \35054 );
nand \U$34679 ( \35056 , \34759 , RIc225828_64);
nand \U$34680 ( \35057 , \35055 , \35056 );
xnor \U$34681 ( \35058 , \35052 , \35057 );
xnor \U$34682 ( \35059 , \35041 , \35058 );
and \U$34683 ( \35060 , \35032 , \35059 );
and \U$34684 ( \35061 , \34789 , \35031 );
or \U$34685 ( \35062 , \35060 , \35061 );
not \U$34686 ( \35063 , \35062 );
not \U$34687 ( \35064 , \35036 );
not \U$34688 ( \35065 , \35058 );
or \U$34689 ( \35066 , \35064 , \35065 );
nand \U$34690 ( \35067 , \35066 , \35034 );
not \U$34691 ( \35068 , \35058 );
nand \U$34692 ( \35069 , \35068 , \35039 );
nand \U$34693 ( \35070 , \35067 , \35069 );
not \U$34694 ( \35071 , \35070 );
xor \U$34695 ( \35072 , \34680 , \34675 );
xnor \U$34696 ( \35073 , \35072 , \34665 );
not \U$34697 ( \35074 , \35057 );
not \U$34698 ( \35075 , \35051 );
or \U$34699 ( \35076 , \35074 , \35075 );
or \U$34700 ( \35077 , \35051 , \35057 );
nand \U$34701 ( \35078 , \35077 , \35046 );
nand \U$34702 ( \35079 , \35076 , \35078 );
xor \U$34703 ( \35080 , \35073 , \35079 );
xor \U$34704 ( \35081 , \34513 , \34534 );
xor \U$34705 ( \35082 , \35081 , \34545 );
not \U$34706 ( \35083 , \35082 );
not \U$34707 ( \35084 , \18037 );
not \U$34708 ( \35085 , \34737 );
or \U$34709 ( \35086 , \35084 , \35085 );
not \U$34710 ( \35087 , RIc225a80_59);
not \U$34711 ( \35088 , \14299 );
or \U$34712 ( \35089 , \35087 , \35088 );
or \U$34713 ( \35090 , \4049 , RIc225a80_59);
nand \U$34714 ( \35091 , \35089 , \35090 );
nand \U$34715 ( \35092 , \35091 , \15164 );
nand \U$34716 ( \35093 , \35086 , \35092 );
not \U$34717 ( \35094 , \35093 );
or \U$34718 ( \35095 , \35083 , \35094 );
or \U$34719 ( \35096 , \35093 , \35082 );
xor \U$34720 ( \35097 , \34514 , \34519 );
xor \U$34721 ( \35098 , \35097 , \34531 );
not \U$34722 ( \35099 , \6307 );
not \U$34723 ( \35100 , \34139 );
or \U$34724 ( \35101 , \35099 , \35100 );
not \U$34725 ( \35102 , RIc2263e0_39);
not \U$34726 ( \35103 , \10800 );
or \U$34727 ( \35104 , \35102 , \35103 );
nand \U$34728 ( \35105 , \9274 , \5498 );
nand \U$34729 ( \35106 , \35104 , \35105 );
nand \U$34730 ( \35107 , \35106 , \6688 );
nand \U$34731 ( \35108 , \35101 , \35107 );
xor \U$34732 ( \35109 , \35098 , \35108 );
not \U$34733 ( \35110 , \9205 );
not \U$34734 ( \35111 , \34373 );
or \U$34735 ( \35112 , \35110 , \35111 );
nand \U$34736 ( \35113 , \34881 , \9110 );
nand \U$34737 ( \35114 , \35112 , \35113 );
and \U$34738 ( \35115 , \35109 , \35114 );
and \U$34739 ( \35116 , \35098 , \35108 );
or \U$34740 ( \35117 , \35115 , \35116 );
nand \U$34741 ( \35118 , \35096 , \35117 );
nand \U$34742 ( \35119 , \35095 , \35118 );
xnor \U$34743 ( \35120 , \35080 , \35119 );
not \U$34744 ( \35121 , \35120 );
not \U$34745 ( \35122 , \35121 );
or \U$34746 ( \35123 , \35071 , \35122 );
not \U$34747 ( \35124 , \35070 );
nand \U$34748 ( \35125 , \35124 , \35120 );
nand \U$34749 ( \35126 , \35123 , \35125 );
xor \U$34750 ( \35127 , \34839 , \34893 );
and \U$34751 ( \35128 , \35127 , \34909 );
and \U$34752 ( \35129 , \34839 , \34893 );
or \U$34753 ( \35130 , \35128 , \35129 );
not \U$34754 ( \35131 , \6688 );
not \U$34755 ( \35132 , \34926 );
or \U$34756 ( \35133 , \35131 , \35132 );
nand \U$34757 ( \35134 , \35106 , \6307 );
nand \U$34758 ( \35135 , \35133 , \35134 );
not \U$34759 ( \35136 , \9705 );
not \U$34760 ( \35137 , RIc2262f0_41);
not \U$34761 ( \35138 , \10814 );
or \U$34762 ( \35139 , \35137 , \35138 );
nand \U$34763 ( \35140 , \10110 , \6303 );
nand \U$34764 ( \35141 , \35139 , \35140 );
not \U$34765 ( \35142 , \35141 );
or \U$34766 ( \35143 , \35136 , \35142 );
not \U$34767 ( \35144 , RIc2262f0_41);
not \U$34768 ( \35145 , \9250 );
or \U$34769 ( \35146 , \35144 , \35145 );
nand \U$34770 ( \35147 , \17014 , \6303 );
nand \U$34771 ( \35148 , \35146 , \35147 );
nand \U$34772 ( \35149 , \35148 , \9690 );
nand \U$34773 ( \35150 , \35143 , \35149 );
xor \U$34774 ( \35151 , \35135 , \35150 );
not \U$34775 ( \35152 , \5519 );
not \U$34776 ( \35153 , RIc2264d0_37);
not \U$34777 ( \35154 , \12100 );
or \U$34778 ( \35155 , \35153 , \35154 );
nand \U$34779 ( \35156 , \9324 , \4371 );
nand \U$34780 ( \35157 , \35155 , \35156 );
not \U$34781 ( \35158 , \35157 );
or \U$34782 ( \35159 , \35152 , \35158 );
and \U$34783 ( \35160 , RIc2264d0_37, \21172 );
not \U$34784 ( \35161 , RIc2264d0_37);
and \U$34785 ( \35162 , \35161 , \10086 );
nor \U$34786 ( \35163 , \35160 , \35162 );
not \U$34787 ( \35164 , \35163 );
nand \U$34788 ( \35165 , \35164 , \5509 );
nand \U$34789 ( \35166 , \35159 , \35165 );
and \U$34790 ( \35167 , \35151 , \35166 );
and \U$34791 ( \35168 , \35135 , \35150 );
or \U$34792 ( \35169 , \35167 , \35168 );
not \U$34793 ( \35170 , RIc225b70_57);
not \U$34794 ( \35171 , \10230 );
or \U$34795 ( \35172 , \35170 , \35171 );
nand \U$34796 ( \35173 , \13515 , \11033 );
nand \U$34797 ( \35174 , \35172 , \35173 );
and \U$34798 ( \35175 , \35174 , \11974 );
and \U$34799 ( \35176 , \35004 , \11965 );
nor \U$34800 ( \35177 , \35175 , \35176 );
not \U$34801 ( \35178 , \35177 );
not \U$34802 ( \35179 , \35178 );
not \U$34803 ( \35180 , \9398 );
not \U$34804 ( \35181 , \34834 );
or \U$34805 ( \35182 , \35180 , \35181 );
not \U$34806 ( \35183 , RIc226110_45);
not \U$34807 ( \35184 , \11405 );
or \U$34808 ( \35185 , \35183 , \35184 );
not \U$34809 ( \35186 , \13129 );
nand \U$34810 ( \35187 , \35186 , \9379 );
nand \U$34811 ( \35188 , \35185 , \35187 );
nand \U$34812 ( \35189 , \35188 , \9934 );
nand \U$34813 ( \35190 , \35182 , \35189 );
not \U$34814 ( \35191 , \35190 );
or \U$34815 ( \35192 , \35179 , \35191 );
not \U$34816 ( \35193 , \35177 );
not \U$34817 ( \35194 , \35190 );
not \U$34818 ( \35195 , \35194 );
or \U$34819 ( \35196 , \35193 , \35195 );
not \U$34820 ( \35197 , \10001 );
not \U$34821 ( \35198 , RIc226020_47);
not \U$34822 ( \35199 , \21866 );
or \U$34823 ( \35200 , \35198 , \35199 );
nand \U$34824 ( \35201 , \8979 , \9624 );
nand \U$34825 ( \35202 , \35200 , \35201 );
not \U$34826 ( \35203 , \35202 );
or \U$34827 ( \35204 , \35197 , \35203 );
not \U$34828 ( \35205 , RIc226020_47);
not \U$34829 ( \35206 , \8953 );
or \U$34830 ( \35207 , \35205 , \35206 );
nand \U$34831 ( \35208 , \8952 , \9624 );
nand \U$34832 ( \35209 , \35207 , \35208 );
nand \U$34833 ( \35210 , \35209 , \10953 );
nand \U$34834 ( \35211 , \35204 , \35210 );
nand \U$34835 ( \35212 , \35196 , \35211 );
nand \U$34836 ( \35213 , \35192 , \35212 );
xor \U$34837 ( \35214 , \35169 , \35213 );
xor \U$34838 ( \35215 , \34790 , \34800 );
xor \U$34839 ( \35216 , \35215 , \34811 );
not \U$34840 ( \35217 , \9552 );
not \U$34841 ( \35218 , RIc225f30_49);
not \U$34842 ( \35219 , \20217 );
or \U$34843 ( \35220 , \35218 , \35219 );
nand \U$34844 ( \35221 , \20216 , \28163 );
nand \U$34845 ( \35222 , \35220 , \35221 );
not \U$34846 ( \35223 , \35222 );
or \U$34847 ( \35224 , \35217 , \35223 );
not \U$34848 ( \35225 , RIc225f30_49);
not \U$34849 ( \35226 , \10858 );
or \U$34850 ( \35227 , \35225 , \35226 );
nand \U$34851 ( \35228 , \23042 , \9541 );
nand \U$34852 ( \35229 , \35227 , \35228 );
nand \U$34853 ( \35230 , \35229 , \9534 );
nand \U$34854 ( \35231 , \35224 , \35230 );
xor \U$34855 ( \35232 , \35216 , \35231 );
not \U$34856 ( \35233 , \15164 );
and \U$34857 ( \35234 , RIc225a80_59, \9842 );
not \U$34858 ( \35235 , RIc225a80_59);
and \U$34859 ( \35236 , \35235 , \22991 );
or \U$34860 ( \35237 , \35234 , \35236 );
not \U$34861 ( \35238 , \35237 );
or \U$34862 ( \35239 , \35233 , \35238 );
and \U$34863 ( \35240 , RIc225a80_59, \4417 );
not \U$34864 ( \35241 , RIc225a80_59);
and \U$34865 ( \35242 , \35241 , \16519 );
or \U$34866 ( \35243 , \35240 , \35242 );
nand \U$34867 ( \35244 , \35243 , \12670 );
nand \U$34868 ( \35245 , \35239 , \35244 );
and \U$34869 ( \35246 , \35232 , \35245 );
and \U$34870 ( \35247 , \35216 , \35231 );
or \U$34871 ( \35248 , \35246 , \35247 );
and \U$34872 ( \35249 , \35214 , \35248 );
and \U$34873 ( \35250 , \35169 , \35213 );
or \U$34874 ( \35251 , \35249 , \35250 );
xor \U$34875 ( \35252 , \35130 , \35251 );
xor \U$34876 ( \35253 , \35098 , \35108 );
xor \U$34877 ( \35254 , \35253 , \35114 );
not \U$34878 ( \35255 , \5509 );
not \U$34879 ( \35256 , \35157 );
or \U$34880 ( \35257 , \35255 , \35256 );
nand \U$34881 ( \35258 , \34156 , \5519 );
nand \U$34882 ( \35259 , \35257 , \35258 );
not \U$34883 ( \35260 , \9816 );
not \U$34884 ( \35261 , \34543 );
or \U$34885 ( \35262 , \35260 , \35261 );
nand \U$34886 ( \35263 , \35141 , \9690 );
nand \U$34887 ( \35264 , \35262 , \35263 );
xor \U$34888 ( \35265 , \35259 , \35264 );
not \U$34889 ( \35266 , \9552 );
not \U$34890 ( \35267 , \34291 );
or \U$34891 ( \35268 , \35266 , \35267 );
nand \U$34892 ( \35269 , \35222 , \9534 );
nand \U$34893 ( \35270 , \35268 , \35269 );
xor \U$34894 ( \35271 , \35265 , \35270 );
xor \U$34895 ( \35272 , \35254 , \35271 );
not \U$34896 ( \35273 , \8777 );
not \U$34897 ( \35274 , \35020 );
or \U$34898 ( \35275 , \35273 , \35274 );
nand \U$34899 ( \35276 , \8788 , \34194 );
nand \U$34900 ( \35277 , \35275 , \35276 );
not \U$34901 ( \35278 , \11697 );
not \U$34902 ( \35279 , RIc225c60_55);
not \U$34903 ( \35280 , \14192 );
or \U$34904 ( \35281 , \35279 , \35280 );
nand \U$34905 ( \35282 , \6492 , \11108 );
nand \U$34906 ( \35283 , \35281 , \35282 );
not \U$34907 ( \35284 , \35283 );
or \U$34908 ( \35285 , \35278 , \35284 );
nand \U$34909 ( \35286 , \34823 , \11038 );
nand \U$34910 ( \35287 , \35285 , \35286 );
or \U$34911 ( \35288 , \35277 , \35287 );
and \U$34912 ( \35289 , \34952 , \34960 );
not \U$34913 ( \35290 , \4381 );
not \U$34914 ( \35291 , RIc2265c0_35);
not \U$34915 ( \35292 , \13198 );
or \U$34916 ( \35293 , \35291 , \35292 );
nand \U$34917 ( \35294 , \12755 , \3620 );
nand \U$34918 ( \35295 , \35293 , \35294 );
not \U$34919 ( \35296 , \35295 );
or \U$34920 ( \35297 , \35290 , \35296 );
nand \U$34921 ( \35298 , \34809 , \4383 );
nand \U$34922 ( \35299 , \35297 , \35298 );
xor \U$34923 ( \35300 , \35289 , \35299 );
not \U$34924 ( \35301 , \34979 );
not \U$34925 ( \35302 , \5509 );
or \U$34926 ( \35303 , \35301 , \35302 );
or \U$34927 ( \35304 , \35163 , \5556 );
nand \U$34928 ( \35305 , \35303 , \35304 );
and \U$34929 ( \35306 , \35300 , \35305 );
and \U$34930 ( \35307 , \35289 , \35299 );
or \U$34931 ( \35308 , \35306 , \35307 );
nand \U$34932 ( \35309 , \35288 , \35308 );
nand \U$34933 ( \35310 , \35287 , \35277 );
nand \U$34934 ( \35311 , \35309 , \35310 );
and \U$34935 ( \35312 , \35272 , \35311 );
and \U$34936 ( \35313 , \35254 , \35271 );
or \U$34937 ( \35314 , \35312 , \35313 );
and \U$34938 ( \35315 , \35252 , \35314 );
and \U$34939 ( \35316 , \35130 , \35251 );
or \U$34940 ( \35317 , \35315 , \35316 );
not \U$34941 ( \35318 , \35317 );
and \U$34942 ( \35319 , \35126 , \35318 );
not \U$34943 ( \35320 , \35126 );
and \U$34944 ( \35321 , \35320 , \35317 );
nor \U$34945 ( \35322 , \35319 , \35321 );
nand \U$34946 ( \35323 , \35063 , \35322 );
not \U$34947 ( \35324 , \35323 );
xor \U$34948 ( \35325 , \35130 , \35251 );
xor \U$34949 ( \35326 , \35325 , \35314 );
not \U$34950 ( \35327 , \35326 );
xor \U$34951 ( \35328 , \35169 , \35213 );
xor \U$34952 ( \35329 , \35328 , \35248 );
not \U$34953 ( \35330 , \11974 );
not \U$34954 ( \35331 , \34459 );
or \U$34955 ( \35332 , \35330 , \35331 );
nand \U$34956 ( \35333 , \35174 , \11965 );
nand \U$34957 ( \35334 , \35332 , \35333 );
not \U$34958 ( \35335 , \9619 );
not \U$34959 ( \35336 , \34395 );
or \U$34960 ( \35337 , \35335 , \35336 );
nand \U$34961 ( \35338 , \35209 , \10001 );
nand \U$34962 ( \35339 , \35337 , \35338 );
xor \U$34963 ( \35340 , \35334 , \35339 );
not \U$34964 ( \35341 , \12670 );
not \U$34965 ( \35342 , \35091 );
or \U$34966 ( \35343 , \35341 , \35342 );
nand \U$34967 ( \35344 , \35243 , \15164 );
nand \U$34968 ( \35345 , \35343 , \35344 );
xor \U$34969 ( \35346 , \35340 , \35345 );
xor \U$34970 ( \35347 , \34188 , \34203 );
xor \U$34971 ( \35348 , \35347 , \34218 );
xor \U$34972 ( \35349 , \35346 , \35348 );
not \U$34973 ( \35350 , \9459 );
not \U$34974 ( \35351 , RIc225e40_51);
not \U$34975 ( \35352 , \20674 );
or \U$34976 ( \35353 , \35351 , \35352 );
nand \U$34977 ( \35354 , \12727 , \12423 );
nand \U$34978 ( \35355 , \35353 , \35354 );
not \U$34979 ( \35356 , \35355 );
or \U$34980 ( \35357 , \35350 , \35356 );
nand \U$34981 ( \35358 , \34179 , \9444 );
nand \U$34982 ( \35359 , \35357 , \35358 );
not \U$34983 ( \35360 , \20862 );
not \U$34984 ( \35361 , \34210 );
or \U$34985 ( \35362 , \35360 , \35361 );
not \U$34986 ( \35363 , RIc225990_61);
not \U$34987 ( \35364 , \19926 );
or \U$34988 ( \35365 , \35363 , \35364 );
nand \U$34989 ( \35366 , \3641 , \12806 );
nand \U$34990 ( \35367 , \35365 , \35366 );
nand \U$34991 ( \35368 , \35367 , \15719 );
nand \U$34992 ( \35369 , \35362 , \35368 );
xor \U$34993 ( \35370 , \35359 , \35369 );
not \U$34994 ( \35371 , RIc225828_64);
not \U$34995 ( \35372 , \34900 );
or \U$34996 ( \35373 , \35371 , \35372 );
not \U$34997 ( \35374 , RIc2258a0_63);
not \U$34998 ( \35375 , \31566 );
or \U$34999 ( \35376 , \35374 , \35375 );
not \U$35000 ( \35377 , \9513 );
nand \U$35001 ( \35378 , \35377 , \28750 );
nand \U$35002 ( \35379 , \35376 , \35378 );
nand \U$35003 ( \35380 , \35379 , \20159 );
nand \U$35004 ( \35381 , \35373 , \35380 );
and \U$35005 ( \35382 , \35370 , \35381 );
and \U$35006 ( \35383 , \35359 , \35369 );
or \U$35007 ( \35384 , \35382 , \35383 );
xor \U$35008 ( \35385 , \35349 , \35384 );
xor \U$35009 ( \35386 , \35329 , \35385 );
xor \U$35010 ( \35387 , \35289 , \35299 );
xor \U$35011 ( \35388 , \35387 , \35305 );
not \U$35012 ( \35389 , \35388 );
not \U$35013 ( \35390 , \6307 );
not \U$35014 ( \35391 , \34919 );
or \U$35015 ( \35392 , \35390 , \35391 );
not \U$35016 ( \35393 , RIc2263e0_39);
not \U$35017 ( \35394 , \21172 );
or \U$35018 ( \35395 , \35393 , \35394 );
nand \U$35019 ( \35396 , \10086 , \8990 );
nand \U$35020 ( \35397 , \35395 , \35396 );
nand \U$35021 ( \35398 , \35397 , \6688 );
nand \U$35022 ( \35399 , \35392 , \35398 );
not \U$35023 ( \35400 , \35399 );
not \U$35024 ( \35401 , \9398 );
not \U$35025 ( \35402 , RIc226110_45);
not \U$35026 ( \35403 , \9046 );
or \U$35027 ( \35404 , \35402 , \35403 );
nand \U$35028 ( \35405 , \9051 , \9379 );
nand \U$35029 ( \35406 , \35404 , \35405 );
not \U$35030 ( \35407 , \35406 );
or \U$35031 ( \35408 , \35401 , \35407 );
not \U$35032 ( \35409 , RIc226110_45);
not \U$35033 ( \35410 , \19789 );
or \U$35034 ( \35411 , \35409 , \35410 );
nand \U$35035 ( \35412 , \32612 , \9100 );
nand \U$35036 ( \35413 , \35411 , \35412 );
nand \U$35037 ( \35414 , \35413 , \9382 );
nand \U$35038 ( \35415 , \35408 , \35414 );
not \U$35039 ( \35416 , \35415 );
or \U$35040 ( \35417 , \35400 , \35416 );
or \U$35041 ( \35418 , \35415 , \35399 );
not \U$35042 ( \35419 , \9705 );
not \U$35043 ( \35420 , RIc2262f0_41);
not \U$35044 ( \35421 , \10800 );
or \U$35045 ( \35422 , \35420 , \35421 );
nand \U$35046 ( \35423 , \9275 , \6303 );
nand \U$35047 ( \35424 , \35422 , \35423 );
not \U$35048 ( \35425 , \35424 );
or \U$35049 ( \35426 , \35419 , \35425 );
not \U$35050 ( \35427 , RIc2262f0_41);
not \U$35051 ( \35428 , \30069 );
or \U$35052 ( \35429 , \35427 , \35428 );
nand \U$35053 ( \35430 , \21150 , \6303 );
nand \U$35054 ( \35431 , \35429 , \35430 );
nand \U$35055 ( \35432 , \35431 , \9690 );
nand \U$35056 ( \35433 , \35426 , \35432 );
nand \U$35057 ( \35434 , \35418 , \35433 );
nand \U$35058 ( \35435 , \35417 , \35434 );
not \U$35059 ( \35436 , \35435 );
or \U$35060 ( \35437 , \35389 , \35436 );
or \U$35061 ( \35438 , \35435 , \35388 );
not \U$35062 ( \35439 , \4383 );
not \U$35063 ( \35440 , \35295 );
or \U$35064 ( \35441 , \35439 , \35440 );
not \U$35065 ( \35442 , RIc2265c0_35);
not \U$35066 ( \35443 , \15444 );
or \U$35067 ( \35444 , \35442 , \35443 );
nand \U$35068 ( \35445 , \15443 , \4376 );
nand \U$35069 ( \35446 , \35444 , \35445 );
nand \U$35070 ( \35447 , \35446 , \5741 );
nand \U$35071 ( \35448 , \35441 , \35447 );
and \U$35072 ( \35449 , \16248 , \2710 );
not \U$35073 ( \35450 , \3630 );
not \U$35074 ( \35451 , \34969 );
or \U$35075 ( \35452 , \35450 , \35451 );
and \U$35076 ( \35453 , \2692 , \20528 );
not \U$35077 ( \35454 , \2692 );
not \U$35078 ( \35455 , \21102 );
and \U$35079 ( \35456 , \35454 , \35455 );
nor \U$35080 ( \35457 , \35453 , \35456 );
nand \U$35081 ( \35458 , \35457 , \3628 );
nand \U$35082 ( \35459 , \35452 , \35458 );
xor \U$35083 ( \35460 , \35449 , \35459 );
not \U$35084 ( \35461 , \4382 );
not \U$35085 ( \35462 , \35446 );
or \U$35086 ( \35463 , \35461 , \35462 );
not \U$35087 ( \35464 , RIc2265c0_35);
not \U$35088 ( \35465 , \12846 );
or \U$35089 ( \35466 , \35464 , \35465 );
nand \U$35090 ( \35467 , \18161 , \3620 );
nand \U$35091 ( \35468 , \35466 , \35467 );
nand \U$35092 ( \35469 , \35468 , \4381 );
nand \U$35093 ( \35470 , \35463 , \35469 );
and \U$35094 ( \35471 , \35460 , \35470 );
and \U$35095 ( \35472 , \35449 , \35459 );
or \U$35096 ( \35473 , \35471 , \35472 );
xor \U$35097 ( \35474 , \35448 , \35473 );
not \U$35098 ( \35475 , \9110 );
not \U$35099 ( \35476 , RIc226200_43);
not \U$35100 ( \35477 , \11488 );
or \U$35101 ( \35478 , \35476 , \35477 );
not \U$35102 ( \35479 , \30875 );
nand \U$35103 ( \35480 , \35479 , \9117 );
nand \U$35104 ( \35481 , \35478 , \35480 );
not \U$35105 ( \35482 , \35481 );
or \U$35106 ( \35483 , \35475 , \35482 );
nand \U$35107 ( \35484 , \34935 , \9129 );
nand \U$35108 ( \35485 , \35483 , \35484 );
and \U$35109 ( \35486 , \35474 , \35485 );
and \U$35110 ( \35487 , \35448 , \35473 );
or \U$35111 ( \35488 , \35486 , \35487 );
nand \U$35112 ( \35489 , \35438 , \35488 );
nand \U$35113 ( \35490 , \35437 , \35489 );
not \U$35114 ( \35491 , \15164 );
and \U$35115 ( \35492 , RIc225a80_59, \10230 );
not \U$35116 ( \35493 , RIc225a80_59);
and \U$35117 ( \35494 , \35493 , \34640 );
or \U$35118 ( \35495 , \35492 , \35494 );
not \U$35119 ( \35496 , \35495 );
or \U$35120 ( \35497 , \35491 , \35496 );
nand \U$35121 ( \35498 , \35237 , \12670 );
nand \U$35122 ( \35499 , \35497 , \35498 );
not \U$35123 ( \35500 , \11708 );
not \U$35124 ( \35501 , \35355 );
or \U$35125 ( \35502 , \35500 , \35501 );
not \U$35126 ( \35503 , RIc225e40_51);
not \U$35127 ( \35504 , \9897 );
or \U$35128 ( \35505 , \35503 , \35504 );
not \U$35129 ( \35506 , \28149 );
nand \U$35130 ( \35507 , \35506 , \22140 );
nand \U$35131 ( \35508 , \35505 , \35507 );
nand \U$35132 ( \35509 , \35508 , \9459 );
nand \U$35133 ( \35510 , \35502 , \35509 );
xor \U$35134 ( \35511 , \35499 , \35510 );
not \U$35135 ( \35512 , \20159 );
not \U$35136 ( \35513 , RIc2258a0_63);
not \U$35137 ( \35514 , \6439 );
or \U$35138 ( \35515 , \35513 , \35514 );
not \U$35139 ( \35516 , \3727 );
nand \U$35140 ( \35517 , \35516 , \15620 );
nand \U$35141 ( \35518 , \35515 , \35517 );
not \U$35142 ( \35519 , \35518 );
or \U$35143 ( \35520 , \35512 , \35519 );
nand \U$35144 ( \35521 , \35379 , RIc225828_64);
nand \U$35145 ( \35522 , \35520 , \35521 );
and \U$35146 ( \35523 , \35511 , \35522 );
and \U$35147 ( \35524 , \35499 , \35510 );
or \U$35148 ( \35525 , \35523 , \35524 );
xor \U$35149 ( \35526 , \35490 , \35525 );
xor \U$35150 ( \35527 , \35359 , \35369 );
xor \U$35151 ( \35528 , \35527 , \35381 );
and \U$35152 ( \35529 , \35526 , \35528 );
and \U$35153 ( \35530 , \35490 , \35525 );
or \U$35154 ( \35531 , \35529 , \35530 );
and \U$35155 ( \35532 , \35386 , \35531 );
and \U$35156 ( \35533 , \35329 , \35385 );
or \U$35157 ( \35534 , \35532 , \35533 );
not \U$35158 ( \35535 , \35534 );
or \U$35159 ( \35536 , \35327 , \35535 );
or \U$35160 ( \35537 , \35534 , \35326 );
xor \U$35161 ( \35538 , \35135 , \35150 );
xor \U$35162 ( \35539 , \35538 , \35166 );
not \U$35163 ( \35540 , \9690 );
not \U$35164 ( \35541 , \35424 );
or \U$35165 ( \35542 , \35540 , \35541 );
nand \U$35166 ( \35543 , \35148 , \9816 );
nand \U$35167 ( \35544 , \35542 , \35543 );
not \U$35168 ( \35545 , \9398 );
not \U$35169 ( \35546 , \35188 );
or \U$35170 ( \35547 , \35545 , \35546 );
nand \U$35171 ( \35548 , \35406 , \9934 );
nand \U$35172 ( \35549 , \35547 , \35548 );
or \U$35173 ( \35550 , \35544 , \35549 );
not \U$35174 ( \35551 , \9534 );
and \U$35175 ( \35552 , RIc225f30_49, \13370 );
not \U$35176 ( \35553 , RIc225f30_49);
and \U$35177 ( \35554 , \35553 , \20368 );
or \U$35178 ( \35555 , \35552 , \35554 );
not \U$35179 ( \35556 , \35555 );
or \U$35180 ( \35557 , \35551 , \35556 );
nand \U$35181 ( \35558 , \35229 , \9552 );
nand \U$35182 ( \35559 , \35557 , \35558 );
nand \U$35183 ( \35560 , \35550 , \35559 );
nand \U$35184 ( \35561 , \35549 , \35544 );
nand \U$35185 ( \35562 , \35560 , \35561 );
xor \U$35186 ( \35563 , \35539 , \35562 );
not \U$35187 ( \35564 , \11117 );
not \U$35188 ( \35565 , RIc225c60_55);
not \U$35189 ( \35566 , \21438 );
or \U$35190 ( \35567 , \35565 , \35566 );
nand \U$35191 ( \35568 , \34709 , \11041 );
nand \U$35192 ( \35569 , \35567 , \35568 );
not \U$35193 ( \35570 , \35569 );
or \U$35194 ( \35571 , \35564 , \35570 );
nand \U$35195 ( \35572 , \35283 , \11038 );
nand \U$35196 ( \35573 , \35571 , \35572 );
not \U$35197 ( \35574 , \15729 );
not \U$35198 ( \35575 , \35367 );
or \U$35199 ( \35576 , \35574 , \35575 );
not \U$35200 ( \35577 , RIc225990_61);
not \U$35201 ( \35578 , \4414 );
or \U$35202 ( \35579 , \35577 , \35578 );
nand \U$35203 ( \35580 , \4418 , \10338 );
nand \U$35204 ( \35581 , \35579 , \35580 );
nand \U$35205 ( \35582 , \35581 , \15719 );
nand \U$35206 ( \35583 , \35576 , \35582 );
nor \U$35207 ( \35584 , \35573 , \35583 );
and \U$35208 ( \35585 , \35202 , \10953 );
not \U$35209 ( \35586 , RIc226020_47);
not \U$35210 ( \35587 , \9787 );
or \U$35211 ( \35588 , \35586 , \35587 );
nand \U$35212 ( \35589 , \17744 , \9373 );
nand \U$35213 ( \35590 , \35588 , \35589 );
not \U$35214 ( \35591 , \35590 );
nor \U$35215 ( \35592 , \35591 , \9640 );
nor \U$35216 ( \35593 , \35585 , \35592 );
or \U$35217 ( \35594 , \35584 , \35593 );
nand \U$35218 ( \35595 , \35583 , \35573 );
nand \U$35219 ( \35596 , \35594 , \35595 );
and \U$35220 ( \35597 , \35563 , \35596 );
and \U$35221 ( \35598 , \35539 , \35562 );
or \U$35222 ( \35599 , \35597 , \35598 );
xor \U$35223 ( \35600 , \35308 , \35277 );
xnor \U$35224 ( \35601 , \35600 , \35287 );
not \U$35225 ( \35602 , \35601 );
not \U$35226 ( \35603 , \35602 );
and \U$35227 ( \35604 , \35211 , \35190 );
not \U$35228 ( \35605 , \35211 );
and \U$35229 ( \35606 , \35605 , \35194 );
nor \U$35230 ( \35607 , \35604 , \35606 );
and \U$35231 ( \35608 , \35607 , \35177 );
not \U$35232 ( \35609 , \35607 );
and \U$35233 ( \35610 , \35609 , \35178 );
nor \U$35234 ( \35611 , \35608 , \35610 );
not \U$35235 ( \35612 , \35611 );
not \U$35236 ( \35613 , \35612 );
or \U$35237 ( \35614 , \35603 , \35613 );
not \U$35238 ( \35615 , \35601 );
not \U$35239 ( \35616 , \35611 );
or \U$35240 ( \35617 , \35615 , \35616 );
xor \U$35241 ( \35618 , \35216 , \35231 );
xor \U$35242 ( \35619 , \35618 , \35245 );
nand \U$35243 ( \35620 , \35617 , \35619 );
nand \U$35244 ( \35621 , \35614 , \35620 );
xor \U$35245 ( \35622 , \35599 , \35621 );
xor \U$35246 ( \35623 , \35254 , \35271 );
xor \U$35247 ( \35624 , \35623 , \35311 );
and \U$35248 ( \35625 , \35622 , \35624 );
and \U$35249 ( \35626 , \35599 , \35621 );
or \U$35250 ( \35627 , \35625 , \35626 );
nand \U$35251 ( \35628 , \35537 , \35627 );
nand \U$35252 ( \35629 , \35536 , \35628 );
not \U$35253 ( \35630 , \35629 );
or \U$35254 ( \35631 , \35324 , \35630 );
not \U$35255 ( \35632 , \35322 );
nand \U$35256 ( \35633 , \35632 , \35062 );
nand \U$35257 ( \35634 , \35631 , \35633 );
xor \U$35258 ( \35635 , \34787 , \35634 );
not \U$35259 ( \35636 , \35070 );
not \U$35260 ( \35637 , \35120 );
or \U$35261 ( \35638 , \35636 , \35637 );
not \U$35262 ( \35639 , \35124 );
not \U$35263 ( \35640 , \35121 );
or \U$35264 ( \35641 , \35639 , \35640 );
nand \U$35265 ( \35642 , \35641 , \35317 );
nand \U$35266 ( \35643 , \35638 , \35642 );
xor \U$35267 ( \35644 , \34782 , \34761 );
xnor \U$35268 ( \35645 , \35644 , \34745 );
not \U$35269 ( \35646 , \35645 );
not \U$35270 ( \35647 , \35646 );
xor \U$35271 ( \35648 , \34548 , \34489 );
xor \U$35272 ( \35649 , \34495 , \35648 );
not \U$35273 ( \35650 , \35649 );
not \U$35274 ( \35651 , \35650 );
or \U$35275 ( \35652 , \35647 , \35651 );
not \U$35276 ( \35653 , \35645 );
not \U$35277 ( \35654 , \35649 );
or \U$35278 ( \35655 , \35653 , \35654 );
xor \U$35279 ( \35656 , \35259 , \35264 );
and \U$35280 ( \35657 , \35656 , \35270 );
and \U$35281 ( \35658 , \35259 , \35264 );
or \U$35282 ( \35659 , \35657 , \35658 );
not \U$35283 ( \35660 , \35659 );
xor \U$35284 ( \35661 , \35334 , \35339 );
and \U$35285 ( \35662 , \35661 , \35345 );
and \U$35286 ( \35663 , \35334 , \35339 );
or \U$35287 ( \35664 , \35662 , \35663 );
not \U$35288 ( \35665 , \35664 );
or \U$35289 ( \35666 , \35660 , \35665 );
or \U$35290 ( \35667 , \35664 , \35659 );
xor \U$35291 ( \35668 , \34814 , \34825 );
and \U$35292 ( \35669 , \35668 , \34836 );
and \U$35293 ( \35670 , \34814 , \34825 );
or \U$35294 ( \35671 , \35669 , \35670 );
nand \U$35295 ( \35672 , \35667 , \35671 );
nand \U$35296 ( \35673 , \35666 , \35672 );
nand \U$35297 ( \35674 , \35655 , \35673 );
nand \U$35298 ( \35675 , \35652 , \35674 );
not \U$35299 ( \35676 , \35079 );
nand \U$35300 ( \35677 , \35676 , \35073 );
and \U$35301 ( \35678 , \35677 , \35119 );
not \U$35302 ( \35679 , \35079 );
nor \U$35303 ( \35680 , \35679 , \35073 );
nor \U$35304 ( \35681 , \35678 , \35680 );
not \U$35305 ( \35682 , \35681 );
and \U$35306 ( \35683 , \35675 , \35682 );
not \U$35307 ( \35684 , \35675 );
and \U$35308 ( \35685 , \35684 , \35681 );
nor \U$35309 ( \35686 , \35683 , \35685 );
xor \U$35310 ( \35687 , \34765 , \34775 );
and \U$35311 ( \35688 , \35687 , \34781 );
and \U$35312 ( \35689 , \34765 , \34775 );
or \U$35313 ( \35690 , \35688 , \35689 );
not \U$35314 ( \35691 , \9129 );
not \U$35315 ( \35692 , \9125 );
not \U$35316 ( \35693 , \8952 );
or \U$35317 ( \35694 , \35692 , \35693 );
not \U$35318 ( \35695 , \9916 );
nand \U$35319 ( \35696 , \35695 , RIc226200_43);
nand \U$35320 ( \35697 , \35694 , \35696 );
not \U$35321 ( \35698 , \35697 );
or \U$35322 ( \35699 , \35691 , \35698 );
nand \U$35323 ( \35700 , \34673 , \9110 );
nand \U$35324 ( \35701 , \35699 , \35700 );
xor \U$35325 ( \35702 , \35690 , \35701 );
not \U$35326 ( \35703 , \9398 );
not \U$35327 ( \35704 , RIc226110_45);
not \U$35328 ( \35705 , \28149 );
or \U$35329 ( \35706 , \35704 , \35705 );
nand \U$35330 ( \35707 , \10289 , \14660 );
nand \U$35331 ( \35708 , \35706 , \35707 );
not \U$35332 ( \35709 , \35708 );
or \U$35333 ( \35710 , \35703 , \35709 );
nand \U$35334 ( \35711 , \34053 , \9384 );
nand \U$35335 ( \35712 , \35710 , \35711 );
xor \U$35336 ( \35713 , \35702 , \35712 );
not \U$35337 ( \35714 , \2697 );
not \U$35338 ( \35715 , \34771 );
or \U$35339 ( \35716 , \35714 , \35715 );
nand \U$35340 ( \35717 , \32800 , \2710 );
nand \U$35341 ( \35718 , \35716 , \35717 );
xor \U$35342 ( \35719 , \34309 , \34319 );
and \U$35343 ( \35720 , \35719 , \34329 );
and \U$35344 ( \35721 , \34309 , \34319 );
or \U$35345 ( \35722 , \35720 , \35721 );
xor \U$35346 ( \35723 , \35718 , \35722 );
not \U$35347 ( \35724 , \6307 );
not \U$35348 ( \35725 , RIc2263e0_39);
not \U$35349 ( \35726 , \10643 );
or \U$35350 ( \35727 , \35725 , \35726 );
nand \U$35351 ( \35728 , \9225 , \9573 );
nand \U$35352 ( \35729 , \35727 , \35728 );
not \U$35353 ( \35730 , \35729 );
or \U$35354 ( \35731 , \35724 , \35730 );
nand \U$35355 ( \35732 , \34336 , \6688 );
nand \U$35356 ( \35733 , \35731 , \35732 );
xor \U$35357 ( \35734 , \35723 , \35733 );
not \U$35358 ( \35735 , \15729 );
not \U$35359 ( \35736 , RIc225990_61);
not \U$35360 ( \35737 , \3799 );
or \U$35361 ( \35738 , \35736 , \35737 );
nand \U$35362 ( \35739 , \20183 , \12806 );
nand \U$35363 ( \35740 , \35738 , \35739 );
not \U$35364 ( \35741 , \35740 );
or \U$35365 ( \35742 , \35735 , \35741 );
nand \U$35366 ( \35743 , \34080 , \15719 );
nand \U$35367 ( \35744 , \35742 , \35743 );
xor \U$35368 ( \35745 , \35734 , \35744 );
not \U$35369 ( \35746 , \18037 );
and \U$35370 ( \35747 , RIc225a80_59, \2104 );
not \U$35371 ( \35748 , RIc225a80_59);
and \U$35372 ( \35749 , \35748 , \4501 );
or \U$35373 ( \35750 , \35747 , \35749 );
not \U$35374 ( \35751 , \35750 );
or \U$35375 ( \35752 , \35746 , \35751 );
nand \U$35376 ( \35753 , \34743 , \15164 );
nand \U$35377 ( \35754 , \35752 , \35753 );
xor \U$35378 ( \35755 , \35745 , \35754 );
xor \U$35379 ( \35756 , \35713 , \35755 );
not \U$35380 ( \35757 , \13025 );
xor \U$35381 ( \35758 , \4418 , \16788 );
nor \U$35382 ( \35759 , \35757 , \35758 );
and \U$35383 ( \35760 , \33979 , \11118 );
nor \U$35384 ( \35761 , \35759 , \35760 );
not \U$35385 ( \35762 , \3732 );
not \U$35386 ( \35763 , \10074 );
or \U$35387 ( \35764 , \35762 , \35763 );
not \U$35388 ( \35765 , \2981 );
nand \U$35389 ( \35766 , \35765 , RIc225b70_57);
nand \U$35390 ( \35767 , \35764 , \35766 );
and \U$35391 ( \35768 , \35767 , \15267 );
and \U$35392 ( \35769 , \34661 , \11965 );
nor \U$35393 ( \35770 , \35768 , \35769 );
xor \U$35394 ( \35771 , \35761 , \35770 );
and \U$35395 ( \35772 , \34752 , \20159 );
not \U$35396 ( \35773 , RIc2258a0_63);
not \U$35397 ( \35774 , \2671 );
or \U$35398 ( \35775 , \35773 , \35774 );
nand \U$35399 ( \35776 , \2720 , \15620 );
nand \U$35400 ( \35777 , \35775 , \35776 );
not \U$35401 ( \35778 , \35777 );
nor \U$35402 ( \35779 , \35778 , \16882 );
nor \U$35403 ( \35780 , \35772 , \35779 );
xor \U$35404 ( \35781 , \35771 , \35780 );
not \U$35405 ( \35782 , \35781 );
xnor \U$35406 ( \35783 , \35756 , \35782 );
not \U$35407 ( \35784 , \35783 );
xor \U$35408 ( \35785 , \35686 , \35784 );
xor \U$35409 ( \35786 , \35643 , \35785 );
xor \U$35410 ( \35787 , \34471 , \34132 );
xnor \U$35411 ( \35788 , \35787 , \34302 );
not \U$35412 ( \35789 , \35788 );
not \U$35413 ( \35790 , \35789 );
xor \U$35414 ( \35791 , \35645 , \35673 );
and \U$35415 ( \35792 , \35791 , \35649 );
not \U$35416 ( \35793 , \35791 );
and \U$35417 ( \35794 , \35793 , \35650 );
nor \U$35418 ( \35795 , \35792 , \35794 );
not \U$35419 ( \35796 , \35795 );
or \U$35420 ( \35797 , \35790 , \35796 );
not \U$35421 ( \35798 , \35795 );
not \U$35422 ( \35799 , \35798 );
not \U$35423 ( \35800 , \35788 );
or \U$35424 ( \35801 , \35799 , \35800 );
xor \U$35425 ( \35802 , \35082 , \35117 );
xor \U$35426 ( \35803 , \35802 , \35093 );
xor \U$35427 ( \35804 , \35346 , \35348 );
and \U$35428 ( \35805 , \35804 , \35384 );
and \U$35429 ( \35806 , \35346 , \35348 );
or \U$35430 ( \35807 , \35805 , \35806 );
xor \U$35431 ( \35808 , \35803 , \35807 );
xor \U$35432 ( \35809 , \35664 , \35671 );
xor \U$35433 ( \35810 , \35809 , \35659 );
and \U$35434 ( \35811 , \35808 , \35810 );
and \U$35435 ( \35812 , \35803 , \35807 );
or \U$35436 ( \35813 , \35811 , \35812 );
nand \U$35437 ( \35814 , \35801 , \35813 );
nand \U$35438 ( \35815 , \35797 , \35814 );
xor \U$35439 ( \35816 , \35786 , \35815 );
xnor \U$35440 ( \35817 , \35635 , \35816 );
xor \U$35441 ( \35818 , \35795 , \35813 );
not \U$35442 ( \35819 , \35789 );
xor \U$35443 ( \35820 , \35818 , \35819 );
xor \U$35444 ( \35821 , \35803 , \35807 );
xor \U$35445 ( \35822 , \35821 , \35810 );
xor \U$35446 ( \35823 , \34789 , \35031 );
xor \U$35447 ( \35824 , \35823 , \35059 );
xor \U$35448 ( \35825 , \35822 , \35824 );
xor \U$35449 ( \35826 , \34837 , \34910 );
xor \U$35450 ( \35827 , \35826 , \35028 );
xor \U$35451 ( \35828 , \34913 , \34946 );
xor \U$35452 ( \35829 , \35828 , \35025 );
xor \U$35453 ( \35830 , \35544 , \35549 );
xnor \U$35454 ( \35831 , \35830 , \35559 );
not \U$35455 ( \35832 , \35831 );
not \U$35456 ( \35833 , \35832 );
not \U$35457 ( \35834 , \10953 );
not \U$35458 ( \35835 , \35590 );
or \U$35459 ( \35836 , \35834 , \35835 );
and \U$35460 ( \35837 , RIc226020_47, \9211 );
not \U$35461 ( \35838 , RIc226020_47);
and \U$35462 ( \35839 , \35838 , \32810 );
nor \U$35463 ( \35840 , \35837 , \35839 );
nand \U$35464 ( \35841 , \35840 , \9641 );
nand \U$35465 ( \35842 , \35836 , \35841 );
not \U$35466 ( \35843 , \35842 );
not \U$35467 ( \35844 , RIc225f30_49);
not \U$35468 ( \35845 , \8975 );
or \U$35469 ( \35846 , \35844 , \35845 );
nand \U$35470 ( \35847 , \11095 , \9549 );
nand \U$35471 ( \35848 , \35846 , \35847 );
not \U$35472 ( \35849 , \35848 );
not \U$35473 ( \35850 , \35849 );
not \U$35474 ( \35851 , \9533 );
and \U$35475 ( \35852 , \35850 , \35851 );
and \U$35476 ( \35853 , \35555 , \9552 );
nor \U$35477 ( \35854 , \35852 , \35853 );
nand \U$35478 ( \35855 , \35843 , \35854 );
xor \U$35479 ( \35856 , \34961 , \34971 );
xor \U$35480 ( \35857 , \35856 , \34988 );
and \U$35481 ( \35858 , \35855 , \35857 );
not \U$35482 ( \35859 , \35842 );
nor \U$35483 ( \35860 , \35859 , \35854 );
nor \U$35484 ( \35861 , \35858 , \35860 );
not \U$35485 ( \35862 , \35861 );
not \U$35486 ( \35863 , \35862 );
or \U$35487 ( \35864 , \35833 , \35863 );
not \U$35488 ( \35865 , \35831 );
not \U$35489 ( \35866 , \35861 );
or \U$35490 ( \35867 , \35865 , \35866 );
or \U$35491 ( \35868 , RIc226638_34, RIc2265c0_35);
nand \U$35492 ( \35869 , \35868 , \18367 );
and \U$35493 ( \35870 , RIc226638_34, RIc2265c0_35);
nor \U$35494 ( \35871 , \35870 , \2692 );
and \U$35495 ( \35872 , \35869 , \35871 );
not \U$35496 ( \35873 , \3630 );
not \U$35497 ( \35874 , \35457 );
or \U$35498 ( \35875 , \35873 , \35874 );
or \U$35499 ( \35876 , \16248 , \2692 );
or \U$35500 ( \35877 , \21954 , RIc2266b0_33);
nand \U$35501 ( \35878 , \35876 , \35877 );
nand \U$35502 ( \35879 , \35878 , \3628 );
nand \U$35503 ( \35880 , \35875 , \35879 );
and \U$35504 ( \35881 , \35872 , \35880 );
not \U$35505 ( \35882 , \5509 );
not \U$35506 ( \35883 , RIc2264d0_37);
not \U$35507 ( \35884 , \16042 );
or \U$35508 ( \35885 , \35883 , \35884 );
nand \U$35509 ( \35886 , \20694 , \5504 );
nand \U$35510 ( \35887 , \35885 , \35886 );
not \U$35511 ( \35888 , \35887 );
or \U$35512 ( \35889 , \35882 , \35888 );
nand \U$35513 ( \35890 , \34986 , \5519 );
nand \U$35514 ( \35891 , \35889 , \35890 );
xor \U$35515 ( \35892 , \35881 , \35891 );
not \U$35516 ( \35893 , \6307 );
not \U$35517 ( \35894 , \35397 );
or \U$35518 ( \35895 , \35893 , \35894 );
not \U$35519 ( \35896 , \27990 );
and \U$35520 ( \35897 , \35896 , \8990 );
not \U$35521 ( \35898 , \35896 );
and \U$35522 ( \35899 , \35898 , RIc2263e0_39);
or \U$35523 ( \35900 , \35897 , \35899 );
nand \U$35524 ( \35901 , \35900 , \6688 );
nand \U$35525 ( \35902 , \35895 , \35901 );
and \U$35526 ( \35903 , \35892 , \35902 );
and \U$35527 ( \35904 , \35881 , \35891 );
or \U$35528 ( \35905 , \35903 , \35904 );
not \U$35529 ( \35906 , \11038 );
not \U$35530 ( \35907 , \35569 );
or \U$35531 ( \35908 , \35906 , \35907 );
not \U$35532 ( \35909 , RIc225c60_55);
not \U$35533 ( \35910 , \10142 );
or \U$35534 ( \35911 , \35909 , \35910 );
nand \U$35535 ( \35912 , \10310 , \11041 );
nand \U$35536 ( \35913 , \35911 , \35912 );
nand \U$35537 ( \35914 , \35913 , \11697 );
nand \U$35538 ( \35915 , \35908 , \35914 );
xor \U$35539 ( \35916 , \35905 , \35915 );
not \U$35540 ( \35917 , \20862 );
not \U$35541 ( \35918 , \35581 );
or \U$35542 ( \35919 , \35917 , \35918 );
not \U$35543 ( \35920 , RIc225990_61);
not \U$35544 ( \35921 , \18450 );
or \U$35545 ( \35922 , \35920 , \35921 );
nand \U$35546 ( \35923 , \4407 , \10338 );
nand \U$35547 ( \35924 , \35922 , \35923 );
nand \U$35548 ( \35925 , \35924 , \15719 );
nand \U$35549 ( \35926 , \35919 , \35925 );
and \U$35550 ( \35927 , \35916 , \35926 );
and \U$35551 ( \35928 , \35905 , \35915 );
or \U$35552 ( \35929 , \35927 , \35928 );
nand \U$35553 ( \35930 , \35867 , \35929 );
nand \U$35554 ( \35931 , \35864 , \35930 );
xor \U$35555 ( \35932 , \35829 , \35931 );
xor \U$35556 ( \35933 , \35539 , \35562 );
xor \U$35557 ( \35934 , \35933 , \35596 );
and \U$35558 ( \35935 , \35932 , \35934 );
and \U$35559 ( \35936 , \35829 , \35931 );
or \U$35560 ( \35937 , \35935 , \35936 );
xor \U$35561 ( \35938 , \35827 , \35937 );
and \U$35562 ( \35939 , \35619 , \35602 );
not \U$35563 ( \35940 , \35619 );
and \U$35564 ( \35941 , \35940 , \35601 );
nor \U$35565 ( \35942 , \35939 , \35941 );
buf \U$35566 ( \35943 , \35612 );
xnor \U$35567 ( \35944 , \35942 , \35943 );
not \U$35568 ( \35945 , \35944 );
not \U$35569 ( \35946 , \35945 );
not \U$35570 ( \35947 , \12670 );
not \U$35571 ( \35948 , \35495 );
or \U$35572 ( \35949 , \35947 , \35948 );
and \U$35573 ( \35950 , RIc225a80_59, \10161 );
not \U$35574 ( \35951 , RIc225a80_59);
and \U$35575 ( \35952 , \35951 , \19859 );
or \U$35576 ( \35953 , \35950 , \35952 );
nand \U$35577 ( \35954 , \35953 , \15164 );
nand \U$35578 ( \35955 , \35949 , \35954 );
not \U$35579 ( \35956 , \35955 );
not \U$35580 ( \35957 , \11974 );
not \U$35581 ( \35958 , \34997 );
or \U$35582 ( \35959 , \35957 , \35958 );
and \U$35583 ( \35960 , RIc225b70_57, \10125 );
not \U$35584 ( \35961 , RIc225b70_57);
and \U$35585 ( \35962 , \35961 , \6494 );
or \U$35586 ( \35963 , \35960 , \35962 );
nand \U$35587 ( \35964 , \35963 , \11965 );
nand \U$35588 ( \35965 , \35959 , \35964 );
not \U$35589 ( \35966 , \35965 );
or \U$35590 ( \35967 , \35956 , \35966 );
or \U$35591 ( \35968 , \35965 , \35955 );
not \U$35592 ( \35969 , \8788 );
not \U$35593 ( \35970 , \35013 );
or \U$35594 ( \35971 , \35969 , \35970 );
not \U$35595 ( \35972 , RIc225d50_53);
not \U$35596 ( \35973 , \20674 );
or \U$35597 ( \35974 , \35972 , \35973 );
nand \U$35598 ( \35975 , \12727 , \8782 );
nand \U$35599 ( \35976 , \35974 , \35975 );
nand \U$35600 ( \35977 , \35976 , \9488 );
nand \U$35601 ( \35978 , \35971 , \35977 );
nand \U$35602 ( \35979 , \35968 , \35978 );
nand \U$35603 ( \35980 , \35967 , \35979 );
not \U$35604 ( \35981 , \35980 );
xor \U$35605 ( \35982 , \35583 , \35573 );
xor \U$35606 ( \35983 , \35982 , \35593 );
nand \U$35607 ( \35984 , \35981 , \35983 );
xor \U$35608 ( \35985 , \34944 , \34928 );
xnor \U$35609 ( \35986 , \35985 , \34939 );
not \U$35610 ( \35987 , \35986 );
and \U$35611 ( \35988 , \35984 , \35987 );
not \U$35612 ( \35989 , \35980 );
nor \U$35613 ( \35990 , \35983 , \35989 );
nor \U$35614 ( \35991 , \35988 , \35990 );
not \U$35615 ( \35992 , \35991 );
not \U$35616 ( \35993 , \35992 );
or \U$35617 ( \35994 , \35946 , \35993 );
not \U$35618 ( \35995 , \35991 );
not \U$35619 ( \35996 , \35944 );
or \U$35620 ( \35997 , \35995 , \35996 );
xor \U$35621 ( \35998 , \34991 , \35006 );
xor \U$35622 ( \35999 , \35998 , \35022 );
not \U$35623 ( \36000 , \9444 );
not \U$35624 ( \36001 , \35508 );
or \U$35625 ( \36002 , \36000 , \36001 );
not \U$35626 ( \36003 , RIc225e40_51);
not \U$35627 ( \36004 , \31842 );
or \U$35628 ( \36005 , \36003 , \36004 );
nand \U$35629 ( \36006 , \8811 , \9450 );
nand \U$35630 ( \36007 , \36005 , \36006 );
nand \U$35631 ( \36008 , \36007 , \9459 );
nand \U$35632 ( \36009 , \36002 , \36008 );
xor \U$35633 ( \36010 , \35449 , \35459 );
xor \U$35634 ( \36011 , \36010 , \35470 );
not \U$35635 ( \36012 , \9934 );
not \U$35636 ( \36013 , RIc226110_45);
not \U$35637 ( \36014 , \10814 );
or \U$35638 ( \36015 , \36013 , \36014 );
nand \U$35639 ( \36016 , \10110 , \14390 );
nand \U$35640 ( \36017 , \36015 , \36016 );
not \U$35641 ( \36018 , \36017 );
or \U$35642 ( \36019 , \36012 , \36018 );
nand \U$35643 ( \36020 , \35413 , \11825 );
nand \U$35644 ( \36021 , \36019 , \36020 );
xor \U$35645 ( \36022 , \36011 , \36021 );
not \U$35646 ( \36023 , \9129 );
not \U$35647 ( \36024 , \35481 );
or \U$35648 ( \36025 , \36023 , \36024 );
not \U$35649 ( \36026 , RIc226200_43);
not \U$35650 ( \36027 , \10975 );
or \U$35651 ( \36028 , \36026 , \36027 );
not \U$35652 ( \36029 , \29689 );
nand \U$35653 ( \36030 , \36029 , \9106 );
nand \U$35654 ( \36031 , \36028 , \36030 );
nand \U$35655 ( \36032 , \36031 , \9110 );
nand \U$35656 ( \36033 , \36025 , \36032 );
and \U$35657 ( \36034 , \36022 , \36033 );
and \U$35658 ( \36035 , \36011 , \36021 );
or \U$35659 ( \36036 , \36034 , \36035 );
xor \U$35660 ( \36037 , \36009 , \36036 );
not \U$35661 ( \36038 , RIc225828_64);
not \U$35662 ( \36039 , \35518 );
or \U$35663 ( \36040 , \36038 , \36039 );
not \U$35664 ( \36041 , RIc2258a0_63);
not \U$35665 ( \36042 , \4046 );
or \U$35666 ( \36043 , \36041 , \36042 );
nand \U$35667 ( \36044 , \3641 , \15620 );
nand \U$35668 ( \36045 , \36043 , \36044 );
nand \U$35669 ( \36046 , \36045 , \20159 );
nand \U$35670 ( \36047 , \36040 , \36046 );
and \U$35671 ( \36048 , \36037 , \36047 );
and \U$35672 ( \36049 , \36009 , \36036 );
or \U$35673 ( \36050 , \36048 , \36049 );
xor \U$35674 ( \36051 , \35999 , \36050 );
xor \U$35675 ( \36052 , \35499 , \35510 );
xor \U$35676 ( \36053 , \36052 , \35522 );
and \U$35677 ( \36054 , \36051 , \36053 );
and \U$35678 ( \36055 , \35999 , \36050 );
or \U$35679 ( \36056 , \36054 , \36055 );
nand \U$35680 ( \36057 , \35997 , \36056 );
nand \U$35681 ( \36058 , \35994 , \36057 );
and \U$35682 ( \36059 , \35938 , \36058 );
and \U$35683 ( \36060 , \35827 , \35937 );
or \U$35684 ( \36061 , \36059 , \36060 );
and \U$35685 ( \36062 , \35825 , \36061 );
and \U$35686 ( \36063 , \35822 , \35824 );
or \U$35687 ( \36064 , \36062 , \36063 );
not \U$35688 ( \36065 , \36064 );
xor \U$35689 ( \36066 , \35820 , \36065 );
xnor \U$35690 ( \36067 , \35062 , \35322 );
not \U$35691 ( \36068 , \35629 );
and \U$35692 ( \36069 , \36067 , \36068 );
not \U$35693 ( \36070 , \36067 );
and \U$35694 ( \36071 , \36070 , \35629 );
nor \U$35695 ( \36072 , \36069 , \36071 );
and \U$35696 ( \36073 , \36066 , \36072 );
and \U$35697 ( \36074 , \35820 , \36065 );
or \U$35698 ( \36075 , \36073 , \36074 );
nand \U$35699 ( \36076 , \35817 , \36075 );
not \U$35700 ( \36077 , \36076 );
xor \U$35701 ( \36078 , \35820 , \36065 );
xor \U$35702 ( \36079 , \36078 , \36072 );
xor \U$35703 ( \36080 , \35822 , \35824 );
xor \U$35704 ( \36081 , \36080 , \36061 );
not \U$35705 ( \36082 , \36081 );
xor \U$35706 ( \36083 , \35627 , \35326 );
xnor \U$35707 ( \36084 , \36083 , \35534 );
nand \U$35708 ( \36085 , \36082 , \36084 );
xor \U$35709 ( \36086 , \35599 , \35621 );
xor \U$35710 ( \36087 , \36086 , \35624 );
xor \U$35711 ( \36088 , \35329 , \35385 );
xor \U$35712 ( \36089 , \36088 , \35531 );
or \U$35713 ( \36090 , \36087 , \36089 );
xor \U$35714 ( \36091 , \35490 , \35525 );
xor \U$35715 ( \36092 , \36091 , \35528 );
not \U$35716 ( \36093 , \36092 );
xor \U$35717 ( \36094 , \35829 , \35931 );
xor \U$35718 ( \36095 , \36094 , \35934 );
not \U$35719 ( \36096 , \36095 );
or \U$35720 ( \36097 , \36093 , \36096 );
or \U$35721 ( \36098 , \36095 , \36092 );
xor \U$35722 ( \36099 , \35399 , \35415 );
xor \U$35723 ( \36100 , \36099 , \35433 );
not \U$35724 ( \36101 , \11697 );
not \U$35725 ( \36102 , RIc225c60_55);
not \U$35726 ( \36103 , \16531 );
or \U$35727 ( \36104 , \36102 , \36103 );
nand \U$35728 ( \36105 , \16532 , \11041 );
nand \U$35729 ( \36106 , \36104 , \36105 );
not \U$35730 ( \36107 , \36106 );
or \U$35731 ( \36108 , \36101 , \36107 );
nand \U$35732 ( \36109 , \35913 , \11038 );
nand \U$35733 ( \36110 , \36108 , \36109 );
not \U$35734 ( \36111 , \36110 );
not \U$35735 ( \36112 , RIc225828_64);
not \U$35736 ( \36113 , \36045 );
or \U$35737 ( \36114 , \36112 , \36113 );
not \U$35738 ( \36115 , RIc2258a0_63);
not \U$35739 ( \36116 , \4414 );
or \U$35740 ( \36117 , \36115 , \36116 );
not \U$35741 ( \36118 , \4417 );
nand \U$35742 ( \36119 , \36118 , \16880 );
nand \U$35743 ( \36120 , \36117 , \36119 );
nand \U$35744 ( \36121 , \36120 , \20159 );
nand \U$35745 ( \36122 , \36114 , \36121 );
not \U$35746 ( \36123 , \36122 );
or \U$35747 ( \36124 , \36111 , \36123 );
or \U$35748 ( \36125 , \36122 , \36110 );
not \U$35749 ( \36126 , \9488 );
not \U$35750 ( \36127 , RIc225d50_53);
not \U$35751 ( \36128 , \20217 );
or \U$35752 ( \36129 , \36127 , \36128 );
nand \U$35753 ( \36130 , \20216 , \11585 );
nand \U$35754 ( \36131 , \36129 , \36130 );
not \U$35755 ( \36132 , \36131 );
or \U$35756 ( \36133 , \36126 , \36132 );
nand \U$35757 ( \36134 , \35976 , \11577 );
nand \U$35758 ( \36135 , \36133 , \36134 );
nand \U$35759 ( \36136 , \36125 , \36135 );
nand \U$35760 ( \36137 , \36124 , \36136 );
xor \U$35761 ( \36138 , \36100 , \36137 );
xor \U$35762 ( \36139 , \35857 , \35842 );
xnor \U$35763 ( \36140 , \36139 , \35854 );
and \U$35764 ( \36141 , \36138 , \36140 );
and \U$35765 ( \36142 , \36100 , \36137 );
or \U$35766 ( \36143 , \36141 , \36142 );
not \U$35767 ( \36144 , \36143 );
xor \U$35768 ( \36145 , \35905 , \35915 );
xor \U$35769 ( \36146 , \36145 , \35926 );
not \U$35770 ( \36147 , \36146 );
xor \U$35771 ( \36148 , \35978 , \35965 );
xnor \U$35772 ( \36149 , \36148 , \35955 );
nand \U$35773 ( \36150 , \36147 , \36149 );
xor \U$35774 ( \36151 , \35881 , \35891 );
xor \U$35775 ( \36152 , \36151 , \35902 );
not \U$35776 ( \36153 , \18037 );
not \U$35777 ( \36154 , \35953 );
or \U$35778 ( \36155 , \36153 , \36154 );
and \U$35779 ( \36156 , RIc225a80_59, \16555 );
not \U$35780 ( \36157 , RIc225a80_59);
and \U$35781 ( \36158 , \36157 , \23776 );
or \U$35782 ( \36159 , \36156 , \36158 );
nand \U$35783 ( \36160 , \36159 , \15164 );
nand \U$35784 ( \36161 , \36155 , \36160 );
xor \U$35785 ( \36162 , \36152 , \36161 );
not \U$35786 ( \36163 , \9459 );
not \U$35787 ( \36164 , RIc225e40_51);
not \U$35788 ( \36165 , \20367 );
or \U$35789 ( \36166 , \36164 , \36165 );
nand \U$35790 ( \36167 , \8952 , \11795 );
nand \U$35791 ( \36168 , \36166 , \36167 );
not \U$35792 ( \36169 , \36168 );
or \U$35793 ( \36170 , \36163 , \36169 );
nand \U$35794 ( \36171 , \36007 , \9445 );
nand \U$35795 ( \36172 , \36170 , \36171 );
and \U$35796 ( \36173 , \36162 , \36172 );
and \U$35797 ( \36174 , \36152 , \36161 );
or \U$35798 ( \36175 , \36173 , \36174 );
and \U$35799 ( \36176 , \36150 , \36175 );
not \U$35800 ( \36177 , \36146 );
nor \U$35801 ( \36178 , \36177 , \36149 );
nor \U$35802 ( \36179 , \36176 , \36178 );
not \U$35803 ( \36180 , \36179 );
not \U$35804 ( \36181 , \36180 );
or \U$35805 ( \36182 , \36144 , \36181 );
not \U$35806 ( \36183 , \36143 );
not \U$35807 ( \36184 , \36183 );
not \U$35808 ( \36185 , \36179 );
or \U$35809 ( \36186 , \36184 , \36185 );
not \U$35810 ( \36187 , \35987 );
not \U$35811 ( \36188 , \35989 );
or \U$35812 ( \36189 , \36187 , \36188 );
nand \U$35813 ( \36190 , \35980 , \35986 );
nand \U$35814 ( \36191 , \36189 , \36190 );
xnor \U$35815 ( \36192 , \36191 , \35983 );
nand \U$35816 ( \36193 , \36186 , \36192 );
nand \U$35817 ( \36194 , \36182 , \36193 );
nand \U$35818 ( \36195 , \36098 , \36194 );
nand \U$35819 ( \36196 , \36097 , \36195 );
nand \U$35820 ( \36197 , \36090 , \36196 );
nand \U$35821 ( \36198 , \36089 , \36087 );
nand \U$35822 ( \36199 , \36197 , \36198 );
buf \U$35823 ( \36200 , \36199 );
and \U$35824 ( \36201 , \36085 , \36200 );
not \U$35825 ( \36202 , \36081 );
nor \U$35826 ( \36203 , \36202 , \36084 );
nor \U$35827 ( \36204 , \36201 , \36203 );
nand \U$35828 ( \36205 , \36079 , \36204 );
not \U$35829 ( \36206 , \36205 );
not \U$35830 ( \36207 , \36199 );
not \U$35831 ( \36208 , \36084 );
and \U$35832 ( \36209 , \36207 , \36208 );
and \U$35833 ( \36210 , \36199 , \36084 );
nor \U$35834 ( \36211 , \36209 , \36210 );
xnor \U$35835 ( \36212 , \36211 , \36081 );
xor \U$35836 ( \36213 , \35827 , \35937 );
xor \U$35837 ( \36214 , \36213 , \36058 );
not \U$35838 ( \36215 , \36214 );
not \U$35839 ( \36216 , \36215 );
xor \U$35840 ( \36217 , \36087 , \36089 );
xnor \U$35841 ( \36218 , \36217 , \36196 );
not \U$35842 ( \36219 , \36218 );
or \U$35843 ( \36220 , \36216 , \36219 );
xor \U$35844 ( \36221 , \35388 , \35488 );
xor \U$35845 ( \36222 , \36221 , \35435 );
xor \U$35846 ( \36223 , \35448 , \35473 );
xor \U$35847 ( \36224 , \36223 , \35485 );
not \U$35848 ( \36225 , \9690 );
not \U$35849 ( \36226 , RIc2262f0_41);
not \U$35850 ( \36227 , \9321 );
or \U$35851 ( \36228 , \36226 , \36227 );
nand \U$35852 ( \36229 , \9320 , \6303 );
nand \U$35853 ( \36230 , \36228 , \36229 );
not \U$35854 ( \36231 , \36230 );
or \U$35855 ( \36232 , \36225 , \36231 );
nand \U$35856 ( \36233 , \35431 , \9816 );
nand \U$35857 ( \36234 , \36232 , \36233 );
not \U$35858 ( \36235 , \9619 );
not \U$35859 ( \36236 , \35840 );
or \U$35860 ( \36237 , \36235 , \36236 );
and \U$35861 ( \36238 , RIc226020_47, \21183 );
not \U$35862 ( \36239 , RIc226020_47);
and \U$35863 ( \36240 , \36239 , \9051 );
or \U$35864 ( \36241 , \36238 , \36240 );
nand \U$35865 ( \36242 , \36241 , \9641 );
nand \U$35866 ( \36243 , \36237 , \36242 );
xor \U$35867 ( \36244 , \36234 , \36243 );
not \U$35868 ( \36245 , \10445 );
not \U$35869 ( \36246 , RIc225f30_49);
not \U$35870 ( \36247 , \9787 );
or \U$35871 ( \36248 , \36246 , \36247 );
nand \U$35872 ( \36249 , \17744 , \9549 );
nand \U$35873 ( \36250 , \36248 , \36249 );
not \U$35874 ( \36251 , \36250 );
or \U$35875 ( \36252 , \36245 , \36251 );
nand \U$35876 ( \36253 , \35848 , \9552 );
nand \U$35877 ( \36254 , \36252 , \36253 );
and \U$35878 ( \36255 , \36244 , \36254 );
and \U$35879 ( \36256 , \36234 , \36243 );
or \U$35880 ( \36257 , \36255 , \36256 );
xor \U$35881 ( \36258 , \36224 , \36257 );
xor \U$35882 ( \36259 , \35872 , \35880 );
not \U$35883 ( \36260 , \36259 );
and \U$35884 ( \36261 , \35468 , \5135 );
and \U$35885 ( \36262 , \3620 , \21094 );
not \U$35886 ( \36263 , \3620 );
and \U$35887 ( \36264 , \36263 , \31281 );
nor \U$35888 ( \36265 , \36262 , \36264 );
not \U$35889 ( \36266 , \36265 );
nor \U$35890 ( \36267 , \36266 , \5740 );
nor \U$35891 ( \36268 , \36261 , \36267 );
nand \U$35892 ( \36269 , \36260 , \36268 );
not \U$35893 ( \36270 , \36269 );
not \U$35894 ( \36271 , \6688 );
not \U$35895 ( \36272 , RIc2263e0_39);
not \U$35896 ( \36273 , \20406 );
not \U$35897 ( \36274 , \36273 );
or \U$35898 ( \36275 , \36272 , \36274 );
nand \U$35899 ( \36276 , \13497 , \5498 );
nand \U$35900 ( \36277 , \36275 , \36276 );
not \U$35901 ( \36278 , \36277 );
or \U$35902 ( \36279 , \36271 , \36278 );
nand \U$35903 ( \36280 , \35900 , \6307 );
nand \U$35904 ( \36281 , \36279 , \36280 );
not \U$35905 ( \36282 , \36281 );
or \U$35906 ( \36283 , \36270 , \36282 );
not \U$35907 ( \36284 , \36268 );
nand \U$35908 ( \36285 , \36284 , \36259 );
nand \U$35909 ( \36286 , \36283 , \36285 );
not \U$35910 ( \36287 , \15729 );
not \U$35911 ( \36288 , \35924 );
or \U$35912 ( \36289 , \36287 , \36288 );
not \U$35913 ( \36290 , RIc225990_61);
not \U$35914 ( \36291 , \9850 );
or \U$35915 ( \36292 , \36290 , \36291 );
nand \U$35916 ( \36293 , \10231 , \10338 );
nand \U$35917 ( \36294 , \36292 , \36293 );
nand \U$35918 ( \36295 , \36294 , \15719 );
nand \U$35919 ( \36296 , \36289 , \36295 );
xor \U$35920 ( \36297 , \36286 , \36296 );
not \U$35921 ( \36298 , \15267 );
not \U$35922 ( \36299 , \35963 );
or \U$35923 ( \36300 , \36298 , \36299 );
not \U$35924 ( \36301 , RIc225b70_57);
not \U$35925 ( \36302 , \6719 );
or \U$35926 ( \36303 , \36301 , \36302 );
nand \U$35927 ( \36304 , \6720 , \11033 );
nand \U$35928 ( \36305 , \36303 , \36304 );
nand \U$35929 ( \36306 , \36305 , \11965 );
nand \U$35930 ( \36307 , \36300 , \36306 );
and \U$35931 ( \36308 , \36297 , \36307 );
and \U$35932 ( \36309 , \36286 , \36296 );
or \U$35933 ( \36310 , \36308 , \36309 );
and \U$35934 ( \36311 , \36258 , \36310 );
and \U$35935 ( \36312 , \36224 , \36257 );
or \U$35936 ( \36313 , \36311 , \36312 );
xor \U$35937 ( \36314 , \36222 , \36313 );
and \U$35938 ( \36315 , \35929 , \35831 );
not \U$35939 ( \36316 , \35929 );
and \U$35940 ( \36317 , \36316 , \35832 );
nor \U$35941 ( \36318 , \36315 , \36317 );
xnor \U$35942 ( \36319 , \35862 , \36318 );
and \U$35943 ( \36320 , \36314 , \36319 );
and \U$35944 ( \36321 , \36222 , \36313 );
or \U$35945 ( \36322 , \36320 , \36321 );
not \U$35946 ( \36323 , \35992 );
not \U$35947 ( \36324 , \36056 );
not \U$35948 ( \36325 , \36324 );
or \U$35949 ( \36326 , \36323 , \36325 );
nand \U$35950 ( \36327 , \36056 , \35991 );
nand \U$35951 ( \36328 , \36326 , \36327 );
and \U$35952 ( \36329 , \36328 , \35945 );
not \U$35953 ( \36330 , \36328 );
and \U$35954 ( \36331 , \36330 , \35944 );
nor \U$35955 ( \36332 , \36329 , \36331 );
xor \U$35956 ( \36333 , \36322 , \36332 );
xor \U$35957 ( \36334 , \35999 , \36050 );
xor \U$35958 ( \36335 , \36334 , \36053 );
xor \U$35959 ( \36336 , \36009 , \36036 );
xor \U$35960 ( \36337 , \36336 , \36047 );
not \U$35961 ( \36338 , \5519 );
not \U$35962 ( \36339 , \35887 );
or \U$35963 ( \36340 , \36338 , \36339 );
not \U$35964 ( \36341 , RIc2264d0_37);
not \U$35965 ( \36342 , \20519 );
or \U$35966 ( \36343 , \36341 , \36342 );
nand \U$35967 ( \36344 , \19721 , \5504 );
nand \U$35968 ( \36345 , \36343 , \36344 );
nand \U$35969 ( \36346 , \36345 , \5509 );
nand \U$35970 ( \36347 , \36340 , \36346 );
and \U$35971 ( \36348 , \18357 , \3630 );
not \U$35972 ( \36349 , \4381 );
and \U$35973 ( \36350 , \4376 , \20528 );
not \U$35974 ( \36351 , \4376 );
and \U$35975 ( \36352 , \36351 , \16256 );
nor \U$35976 ( \36353 , \36350 , \36352 );
not \U$35977 ( \36354 , \36353 );
or \U$35978 ( \36355 , \36349 , \36354 );
nand \U$35979 ( \36356 , \36265 , \4382 );
nand \U$35980 ( \36357 , \36355 , \36356 );
xor \U$35981 ( \36358 , \36348 , \36357 );
not \U$35982 ( \36359 , \5509 );
not \U$35983 ( \36360 , RIc2264d0_37);
not \U$35984 ( \36361 , \34523 );
or \U$35985 ( \36362 , \36360 , \36361 );
nand \U$35986 ( \36363 , \15633 , \5514 );
nand \U$35987 ( \36364 , \36362 , \36363 );
not \U$35988 ( \36365 , \36364 );
or \U$35989 ( \36366 , \36359 , \36365 );
nand \U$35990 ( \36367 , \36345 , \5519 );
nand \U$35991 ( \36368 , \36366 , \36367 );
and \U$35992 ( \36369 , \36358 , \36368 );
and \U$35993 ( \36370 , \36348 , \36357 );
or \U$35994 ( \36371 , \36369 , \36370 );
xor \U$35995 ( \36372 , \36347 , \36371 );
not \U$35996 ( \36373 , \9398 );
not \U$35997 ( \36374 , \36017 );
or \U$35998 ( \36375 , \36373 , \36374 );
not \U$35999 ( \36376 , \9256 );
not \U$36000 ( \36377 , \22795 );
and \U$36001 ( \36378 , \36376 , \36377 );
and \U$36002 ( \36379 , \27239 , \9100 );
nor \U$36003 ( \36380 , \36378 , \36379 );
not \U$36004 ( \36381 , \36380 );
nand \U$36005 ( \36382 , \36381 , \9384 );
nand \U$36006 ( \36383 , \36375 , \36382 );
and \U$36007 ( \36384 , \36372 , \36383 );
and \U$36008 ( \36385 , \36347 , \36371 );
or \U$36009 ( \36386 , \36384 , \36385 );
not \U$36010 ( \36387 , \9205 );
not \U$36011 ( \36388 , \36031 );
or \U$36012 ( \36389 , \36387 , \36388 );
not \U$36013 ( \36390 , RIc226200_43);
not \U$36014 ( \36391 , \9300 );
or \U$36015 ( \36392 , \36390 , \36391 );
nand \U$36016 ( \36393 , \21150 , \9117 );
nand \U$36017 ( \36394 , \36392 , \36393 );
nand \U$36018 ( \36395 , \36394 , \9110 );
nand \U$36019 ( \36396 , \36389 , \36395 );
not \U$36020 ( \36397 , \9705 );
not \U$36021 ( \36398 , \36230 );
or \U$36022 ( \36399 , \36397 , \36398 );
not \U$36023 ( \36400 , RIc2262f0_41);
not \U$36024 ( \36401 , \31894 );
or \U$36025 ( \36402 , \36400 , \36401 );
nand \U$36026 ( \36403 , \10086 , \17820 );
nand \U$36027 ( \36404 , \36402 , \36403 );
nand \U$36028 ( \36405 , \36404 , \9690 );
nand \U$36029 ( \36406 , \36399 , \36405 );
xor \U$36030 ( \36407 , \36396 , \36406 );
not \U$36031 ( \36408 , \10001 );
not \U$36032 ( \36409 , RIc226020_47);
not \U$36033 ( \36410 , \11394 );
or \U$36034 ( \36411 , \36409 , \36410 );
not \U$36035 ( \36412 , \9073 );
nand \U$36036 ( \36413 , \36412 , \9624 );
nand \U$36037 ( \36414 , \36411 , \36413 );
not \U$36038 ( \36415 , \36414 );
or \U$36039 ( \36416 , \36408 , \36415 );
nand \U$36040 ( \36417 , \36241 , \10953 );
nand \U$36041 ( \36418 , \36416 , \36417 );
and \U$36042 ( \36419 , \36407 , \36418 );
and \U$36043 ( \36420 , \36396 , \36406 );
or \U$36044 ( \36421 , \36419 , \36420 );
xor \U$36045 ( \36422 , \36386 , \36421 );
xor \U$36046 ( \36423 , \36234 , \36243 );
xor \U$36047 ( \36424 , \36423 , \36254 );
and \U$36048 ( \36425 , \36422 , \36424 );
and \U$36049 ( \36426 , \36386 , \36421 );
or \U$36050 ( \36427 , \36425 , \36426 );
xor \U$36051 ( \36428 , \36337 , \36427 );
xor \U$36052 ( \36429 , \36011 , \36021 );
xor \U$36053 ( \36430 , \36429 , \36033 );
not \U$36054 ( \36431 , \16891 );
not \U$36055 ( \36432 , RIc2258a0_63);
not \U$36056 ( \36433 , \24549 );
or \U$36057 ( \36434 , \36432 , \36433 );
not \U$36058 ( \36435 , \9842 );
nand \U$36059 ( \36436 , \36435 , \16880 );
nand \U$36060 ( \36437 , \36434 , \36436 );
not \U$36061 ( \36438 , \36437 );
or \U$36062 ( \36439 , \36431 , \36438 );
nand \U$36063 ( \36440 , \36120 , RIc225828_64);
nand \U$36064 ( \36441 , \36439 , \36440 );
not \U$36065 ( \36442 , \36441 );
not \U$36066 ( \36443 , \15164 );
and \U$36067 ( \36444 , RIc225a80_59, \6493 );
not \U$36068 ( \36445 , RIc225a80_59);
and \U$36069 ( \36446 , \36445 , \27798 );
or \U$36070 ( \36447 , \36444 , \36446 );
not \U$36071 ( \36448 , \36447 );
or \U$36072 ( \36449 , \36443 , \36448 );
nand \U$36073 ( \36450 , \36159 , \12670 );
nand \U$36074 ( \36451 , \36449 , \36450 );
not \U$36075 ( \36452 , \36451 );
or \U$36076 ( \36453 , \36442 , \36452 );
or \U$36077 ( \36454 , \36441 , \36451 );
not \U$36078 ( \36455 , \9488 );
not \U$36079 ( \36456 , RIc225d50_53);
not \U$36080 ( \36457 , \31842 );
or \U$36081 ( \36458 , \36456 , \36457 );
nand \U$36082 ( \36459 , \8811 , \8782 );
nand \U$36083 ( \36460 , \36458 , \36459 );
not \U$36084 ( \36461 , \36460 );
or \U$36085 ( \36462 , \36455 , \36461 );
nand \U$36086 ( \36463 , \36131 , \11577 );
nand \U$36087 ( \36464 , \36462 , \36463 );
nand \U$36088 ( \36465 , \36454 , \36464 );
nand \U$36089 ( \36466 , \36453 , \36465 );
xor \U$36090 ( \36467 , \36430 , \36466 );
not \U$36091 ( \36468 , \11965 );
not \U$36092 ( \36469 , RIc225b70_57);
not \U$36093 ( \36470 , \10609 );
or \U$36094 ( \36471 , \36469 , \36470 );
nand \U$36095 ( \36472 , \15700 , \10074 );
nand \U$36096 ( \36473 , \36471 , \36472 );
not \U$36097 ( \36474 , \36473 );
or \U$36098 ( \36475 , \36468 , \36474 );
nand \U$36099 ( \36476 , \36305 , \11974 );
nand \U$36100 ( \36477 , \36475 , \36476 );
not \U$36101 ( \36478 , \36477 );
not \U$36102 ( \36479 , \11117 );
not \U$36103 ( \36480 , RIc225c60_55);
not \U$36104 ( \36481 , \12724 );
or \U$36105 ( \36482 , \36480 , \36481 );
nand \U$36106 ( \36483 , \31447 , \11108 );
nand \U$36107 ( \36484 , \36482 , \36483 );
not \U$36108 ( \36485 , \36484 );
or \U$36109 ( \36486 , \36479 , \36485 );
nand \U$36110 ( \36487 , \36106 , \12532 );
nand \U$36111 ( \36488 , \36486 , \36487 );
not \U$36112 ( \36489 , \36488 );
or \U$36113 ( \36490 , \36478 , \36489 );
or \U$36114 ( \36491 , \36488 , \36477 );
or \U$36115 ( \36492 , RIc226548_36, RIc2264d0_37);
nand \U$36116 ( \36493 , \36492 , \18367 );
and \U$36117 ( \36494 , RIc226548_36, RIc2264d0_37);
nor \U$36118 ( \36495 , \36494 , \3620 );
and \U$36119 ( \36496 , \36493 , \36495 );
not \U$36120 ( \36497 , \4382 );
not \U$36121 ( \36498 , \36353 );
or \U$36122 ( \36499 , \36497 , \36498 );
or \U$36123 ( \36500 , \18367 , \3620 );
or \U$36124 ( \36501 , \21954 , RIc2265c0_35);
nand \U$36125 ( \36502 , \36500 , \36501 );
nand \U$36126 ( \36503 , \36502 , \4380 );
nand \U$36127 ( \36504 , \36499 , \36503 );
and \U$36128 ( \36505 , \36496 , \36504 );
not \U$36129 ( \36506 , \6307 );
not \U$36130 ( \36507 , \36277 );
or \U$36131 ( \36508 , \36506 , \36507 );
not \U$36132 ( \36509 , RIc2263e0_39);
not \U$36133 ( \36510 , \20690 );
or \U$36134 ( \36511 , \36509 , \36510 );
nand \U$36135 ( \36512 , \12756 , \8990 );
nand \U$36136 ( \36513 , \36511 , \36512 );
nand \U$36137 ( \36514 , \36513 , \6688 );
nand \U$36138 ( \36515 , \36508 , \36514 );
xor \U$36139 ( \36516 , \36505 , \36515 );
not \U$36140 ( \36517 , \9705 );
not \U$36141 ( \36518 , \36404 );
or \U$36142 ( \36519 , \36517 , \36518 );
not \U$36143 ( \36520 , RIc2262f0_41);
not \U$36144 ( \36521 , \10199 );
or \U$36145 ( \36522 , \36520 , \36521 );
nand \U$36146 ( \36523 , \35896 , \6303 );
nand \U$36147 ( \36524 , \36522 , \36523 );
nand \U$36148 ( \36525 , \36524 , \9690 );
nand \U$36149 ( \36526 , \36519 , \36525 );
and \U$36150 ( \36527 , \36516 , \36526 );
and \U$36151 ( \36528 , \36505 , \36515 );
or \U$36152 ( \36529 , \36527 , \36528 );
nand \U$36153 ( \36530 , \36491 , \36529 );
nand \U$36154 ( \36531 , \36490 , \36530 );
and \U$36155 ( \36532 , \36467 , \36531 );
and \U$36156 ( \36533 , \36430 , \36466 );
or \U$36157 ( \36534 , \36532 , \36533 );
and \U$36158 ( \36535 , \36428 , \36534 );
and \U$36159 ( \36536 , \36337 , \36427 );
or \U$36160 ( \36537 , \36535 , \36536 );
xor \U$36161 ( \36538 , \36335 , \36537 );
xor \U$36162 ( \36539 , \36224 , \36257 );
xor \U$36163 ( \36540 , \36539 , \36310 );
not \U$36164 ( \36541 , \9552 );
not \U$36165 ( \36542 , \36250 );
or \U$36166 ( \36543 , \36541 , \36542 );
not \U$36167 ( \36544 , RIc225f30_49);
not \U$36168 ( \36545 , \34344 );
or \U$36169 ( \36546 , \36544 , \36545 );
nand \U$36170 ( \36547 , \9216 , \9549 );
nand \U$36171 ( \36548 , \36546 , \36547 );
nand \U$36172 ( \36549 , \36548 , \9534 );
nand \U$36173 ( \36550 , \36543 , \36549 );
not \U$36174 ( \36551 , \36550 );
not \U$36175 ( \36552 , \15719 );
not \U$36176 ( \36553 , RIc225990_61);
not \U$36177 ( \36554 , \10161 );
or \U$36178 ( \36555 , \36553 , \36554 );
nand \U$36179 ( \36556 , \6726 , \12806 );
nand \U$36180 ( \36557 , \36555 , \36556 );
not \U$36181 ( \36558 , \36557 );
or \U$36182 ( \36559 , \36552 , \36558 );
nand \U$36183 ( \36560 , \36294 , \20862 );
nand \U$36184 ( \36561 , \36559 , \36560 );
not \U$36185 ( \36562 , \36561 );
or \U$36186 ( \36563 , \36551 , \36562 );
or \U$36187 ( \36564 , \36561 , \36550 );
xor \U$36188 ( \36565 , \36259 , \36284 );
xnor \U$36189 ( \36566 , \36565 , \36281 );
not \U$36190 ( \36567 , \36566 );
nand \U$36191 ( \36568 , \36564 , \36567 );
nand \U$36192 ( \36569 , \36563 , \36568 );
xor \U$36193 ( \36570 , \36286 , \36296 );
xor \U$36194 ( \36571 , \36570 , \36307 );
xor \U$36195 ( \36572 , \36569 , \36571 );
xor \U$36196 ( \36573 , \36152 , \36161 );
xor \U$36197 ( \36574 , \36573 , \36172 );
and \U$36198 ( \36575 , \36572 , \36574 );
and \U$36199 ( \36576 , \36569 , \36571 );
or \U$36200 ( \36577 , \36575 , \36576 );
xor \U$36201 ( \36578 , \36540 , \36577 );
xor \U$36202 ( \36579 , \36100 , \36137 );
xor \U$36203 ( \36580 , \36579 , \36140 );
and \U$36204 ( \36581 , \36578 , \36580 );
and \U$36205 ( \36582 , \36540 , \36577 );
or \U$36206 ( \36583 , \36581 , \36582 );
and \U$36207 ( \36584 , \36538 , \36583 );
and \U$36208 ( \36585 , \36335 , \36537 );
or \U$36209 ( \36586 , \36584 , \36585 );
and \U$36210 ( \36587 , \36333 , \36586 );
and \U$36211 ( \36588 , \36322 , \36332 );
or \U$36212 ( \36589 , \36587 , \36588 );
nand \U$36213 ( \36590 , \36220 , \36589 );
or \U$36214 ( \36591 , \36218 , \36215 );
nand \U$36215 ( \36592 , \36590 , \36591 );
nor \U$36216 ( \36593 , \36212 , \36592 );
xor \U$36217 ( \36594 , \36214 , \36218 );
xnor \U$36218 ( \36595 , \36594 , \36589 );
and \U$36219 ( \36596 , \36095 , \36092 );
not \U$36220 ( \36597 , \36095 );
not \U$36221 ( \36598 , \36092 );
and \U$36222 ( \36599 , \36597 , \36598 );
nor \U$36223 ( \36600 , \36596 , \36599 );
buf \U$36224 ( \36601 , \36194 );
xor \U$36225 ( \36602 , \36600 , \36601 );
xor \U$36226 ( \36603 , \36143 , \36180 );
xor \U$36227 ( \36604 , \36603 , \36192 );
not \U$36228 ( \36605 , \36604 );
xor \U$36229 ( \36606 , \36222 , \36313 );
xor \U$36230 ( \36607 , \36606 , \36319 );
not \U$36231 ( \36608 , \36607 );
nand \U$36232 ( \36609 , \36605 , \36608 );
not \U$36233 ( \36610 , \36609 );
xor \U$36234 ( \36611 , \36335 , \36537 );
xor \U$36235 ( \36612 , \36611 , \36583 );
not \U$36236 ( \36613 , \36612 );
or \U$36237 ( \36614 , \36610 , \36613 );
nand \U$36238 ( \36615 , \36604 , \36607 );
nand \U$36239 ( \36616 , \36614 , \36615 );
xor \U$36240 ( \36617 , \36602 , \36616 );
xor \U$36241 ( \36618 , \36322 , \36332 );
xor \U$36242 ( \36619 , \36618 , \36586 );
and \U$36243 ( \36620 , \36617 , \36619 );
and \U$36244 ( \36621 , \36602 , \36616 );
or \U$36245 ( \36622 , \36620 , \36621 );
nand \U$36246 ( \36623 , \36595 , \36622 );
or \U$36247 ( \36624 , \36593 , \36623 );
nand \U$36248 ( \36625 , \36212 , \36592 );
nand \U$36249 ( \36626 , \36624 , \36625 );
not \U$36250 ( \36627 , \36626 );
or \U$36251 ( \36628 , \36206 , \36627 );
or \U$36252 ( \36629 , \36079 , \36204 );
nand \U$36253 ( \36630 , \36628 , \36629 );
not \U$36254 ( \36631 , \36630 );
or \U$36255 ( \36632 , \36077 , \36631 );
or \U$36256 ( \36633 , \35817 , \36075 );
nand \U$36257 ( \36634 , \36632 , \36633 );
not \U$36258 ( \36635 , \36595 );
not \U$36259 ( \36636 , \36622 );
nand \U$36260 ( \36637 , \36635 , \36636 );
not \U$36261 ( \36638 , \36637 );
nor \U$36262 ( \36639 , \36638 , \36593 );
nand \U$36263 ( \36640 , \36639 , \36076 , \36205 );
xor \U$36264 ( \36641 , \36175 , \36146 );
xnor \U$36265 ( \36642 , \36641 , \36149 );
xor \U$36266 ( \36643 , \36135 , \36110 );
xor \U$36267 ( \36644 , \36643 , \36122 );
not \U$36268 ( \36645 , \9459 );
not \U$36269 ( \36646 , RIc225e40_51);
not \U$36270 ( \36647 , \11094 );
or \U$36271 ( \36648 , \36646 , \36647 );
nand \U$36272 ( \36649 , \11095 , \22140 );
nand \U$36273 ( \36650 , \36648 , \36649 );
not \U$36274 ( \36651 , \36650 );
or \U$36275 ( \36652 , \36645 , \36651 );
nand \U$36276 ( \36653 , \36168 , \11708 );
nand \U$36277 ( \36654 , \36652 , \36653 );
xor \U$36278 ( \36655 , \36347 , \36371 );
xor \U$36279 ( \36656 , \36655 , \36383 );
or \U$36280 ( \36657 , \36654 , \36656 );
xor \U$36281 ( \36658 , \36348 , \36357 );
xor \U$36282 ( \36659 , \36658 , \36368 );
not \U$36283 ( \36660 , RIc226110_45);
not \U$36284 ( \36661 , \9276 );
or \U$36285 ( \36662 , \36660 , \36661 );
nand \U$36286 ( \36663 , \10976 , \10429 );
nand \U$36287 ( \36664 , \36662 , \36663 );
not \U$36288 ( \36665 , \36664 );
or \U$36289 ( \36666 , \36665 , \9383 );
not \U$36290 ( \36667 , \11825 );
or \U$36291 ( \36668 , \36380 , \36667 );
nand \U$36292 ( \36669 , \36666 , \36668 );
xor \U$36293 ( \36670 , \36659 , \36669 );
not \U$36294 ( \36671 , \10953 );
not \U$36295 ( \36672 , \36414 );
or \U$36296 ( \36673 , \36671 , \36672 );
not \U$36297 ( \36674 , RIc226020_47);
not \U$36298 ( \36675 , \10111 );
or \U$36299 ( \36676 , \36674 , \36675 );
nand \U$36300 ( \36677 , \10110 , \11607 );
nand \U$36301 ( \36678 , \36676 , \36677 );
nand \U$36302 ( \36679 , \36678 , \9641 );
nand \U$36303 ( \36680 , \36673 , \36679 );
and \U$36304 ( \36681 , \36670 , \36680 );
and \U$36305 ( \36682 , \36659 , \36669 );
or \U$36306 ( \36683 , \36681 , \36682 );
nand \U$36307 ( \36684 , \36657 , \36683 );
nand \U$36308 ( \36685 , \36654 , \36656 );
nand \U$36309 ( \36686 , \36684 , \36685 );
xor \U$36310 ( \36687 , \36644 , \36686 );
xor \U$36311 ( \36688 , \36386 , \36421 );
xor \U$36312 ( \36689 , \36688 , \36424 );
and \U$36313 ( \36690 , \36687 , \36689 );
and \U$36314 ( \36691 , \36644 , \36686 );
or \U$36315 ( \36692 , \36690 , \36691 );
xor \U$36316 ( \36693 , \36642 , \36692 );
xor \U$36317 ( \36694 , \36430 , \36466 );
xor \U$36318 ( \36695 , \36694 , \36531 );
not \U$36319 ( \36696 , \9129 );
not \U$36320 ( \36697 , \36394 );
or \U$36321 ( \36698 , \36696 , \36697 );
not \U$36322 ( \36699 , RIc226200_43);
not \U$36323 ( \36700 , \9321 );
or \U$36324 ( \36701 , \36699 , \36700 );
nand \U$36325 ( \36702 , \9320 , \13805 );
nand \U$36326 ( \36703 , \36701 , \36702 );
nand \U$36327 ( \36704 , \36703 , \9110 );
nand \U$36328 ( \36705 , \36698 , \36704 );
not \U$36329 ( \36706 , \36705 );
not \U$36330 ( \36707 , \11965 );
not \U$36331 ( \36708 , RIc225b70_57);
not \U$36332 ( \36709 , \8887 );
or \U$36333 ( \36710 , \36708 , \36709 );
nand \U$36334 ( \36711 , \17582 , \11033 );
nand \U$36335 ( \36712 , \36710 , \36711 );
not \U$36336 ( \36713 , \36712 );
or \U$36337 ( \36714 , \36707 , \36713 );
nand \U$36338 ( \36715 , \36473 , \11974 );
nand \U$36339 ( \36716 , \36714 , \36715 );
not \U$36340 ( \36717 , \36716 );
or \U$36341 ( \36718 , \36706 , \36717 );
or \U$36342 ( \36719 , \36716 , \36705 );
and \U$36343 ( \36720 , \9541 , \9051 );
not \U$36344 ( \36721 , \9541 );
and \U$36345 ( \36722 , \36721 , \21183 );
nor \U$36346 ( \36723 , \36720 , \36722 );
not \U$36347 ( \36724 , \36723 );
not \U$36348 ( \36725 , \9533 );
and \U$36349 ( \36726 , \36724 , \36725 );
and \U$36350 ( \36727 , \36548 , \9552 );
nor \U$36351 ( \36728 , \36726 , \36727 );
not \U$36352 ( \36729 , \36728 );
nand \U$36353 ( \36730 , \36719 , \36729 );
nand \U$36354 ( \36731 , \36718 , \36730 );
not \U$36355 ( \36732 , \36731 );
not \U$36356 ( \36733 , \36732 );
not \U$36357 ( \36734 , \13025 );
not \U$36358 ( \36735 , \36484 );
or \U$36359 ( \36736 , \36734 , \36735 );
not \U$36360 ( \36737 , RIc225c60_55);
not \U$36361 ( \36738 , \9897 );
or \U$36362 ( \36739 , \36737 , \36738 );
nand \U$36363 ( \36740 , \22969 , \11108 );
nand \U$36364 ( \36741 , \36739 , \36740 );
nand \U$36365 ( \36742 , \36741 , \11117 );
nand \U$36366 ( \36743 , \36736 , \36742 );
not \U$36367 ( \36744 , \36743 );
not \U$36368 ( \36745 , \15164 );
xnor \U$36369 ( \36746 , RIc225a80_59, \6719 );
not \U$36370 ( \36747 , \36746 );
or \U$36371 ( \36748 , \36745 , \36747 );
nand \U$36372 ( \36749 , \36447 , \12670 );
nand \U$36373 ( \36750 , \36748 , \36749 );
not \U$36374 ( \36751 , \36750 );
nand \U$36375 ( \36752 , \36744 , \36751 );
not \U$36376 ( \36753 , \9488 );
not \U$36377 ( \36754 , RIc225d50_53);
not \U$36378 ( \36755 , \13370 );
or \U$36379 ( \36756 , \36754 , \36755 );
not \U$36380 ( \36757 , \9912 );
nand \U$36381 ( \36758 , \36757 , \8782 );
nand \U$36382 ( \36759 , \36756 , \36758 );
not \U$36383 ( \36760 , \36759 );
or \U$36384 ( \36761 , \36753 , \36760 );
nand \U$36385 ( \36762 , \36460 , \8788 );
nand \U$36386 ( \36763 , \36761 , \36762 );
and \U$36387 ( \36764 , \36752 , \36763 );
not \U$36388 ( \36765 , \36743 );
nor \U$36389 ( \36766 , \36765 , \36751 );
nor \U$36390 ( \36767 , \36764 , \36766 );
not \U$36391 ( \36768 , \36767 );
or \U$36392 ( \36769 , \36733 , \36768 );
xor \U$36393 ( \36770 , \36496 , \36504 );
not \U$36394 ( \36771 , \5519 );
not \U$36395 ( \36772 , \36364 );
or \U$36396 ( \36773 , \36771 , \36772 );
not \U$36397 ( \36774 , RIc2264d0_37);
not \U$36398 ( \36775 , \15623 );
or \U$36399 ( \36776 , \36774 , \36775 );
nand \U$36400 ( \36777 , \13488 , \12522 );
nand \U$36401 ( \36778 , \36776 , \36777 );
nand \U$36402 ( \36779 , \36778 , \5509 );
nand \U$36403 ( \36780 , \36773 , \36779 );
xor \U$36404 ( \36781 , \36770 , \36780 );
not \U$36405 ( \36782 , \9690 );
not \U$36406 ( \36783 , RIc2262f0_41);
not \U$36407 ( \36784 , \17625 );
or \U$36408 ( \36785 , \36783 , \36784 );
nand \U$36409 ( \36786 , \20406 , \6303 );
nand \U$36410 ( \36787 , \36785 , \36786 );
not \U$36411 ( \36788 , \36787 );
or \U$36412 ( \36789 , \36782 , \36788 );
nand \U$36413 ( \36790 , \36524 , \9705 );
nand \U$36414 ( \36791 , \36789 , \36790 );
and \U$36415 ( \36792 , \36781 , \36791 );
and \U$36416 ( \36793 , \36770 , \36780 );
or \U$36417 ( \36794 , \36792 , \36793 );
not \U$36418 ( \36795 , \15729 );
not \U$36419 ( \36796 , \36557 );
or \U$36420 ( \36797 , \36795 , \36796 );
not \U$36421 ( \36798 , RIc225990_61);
not \U$36422 ( \36799 , \16555 );
or \U$36423 ( \36800 , \36798 , \36799 );
not \U$36424 ( \36801 , \10170 );
nand \U$36425 ( \36802 , \36801 , \10338 );
nand \U$36426 ( \36803 , \36800 , \36802 );
nand \U$36427 ( \36804 , \36803 , \15719 );
nand \U$36428 ( \36805 , \36797 , \36804 );
xor \U$36429 ( \36806 , \36794 , \36805 );
not \U$36430 ( \36807 , RIc225828_64);
not \U$36431 ( \36808 , \36437 );
or \U$36432 ( \36809 , \36807 , \36808 );
and \U$36433 ( \36810 , \5216 , RIc2258a0_63);
not \U$36434 ( \36811 , \5216 );
and \U$36435 ( \36812 , \36811 , \15620 );
or \U$36436 ( \36813 , \36810 , \36812 );
nand \U$36437 ( \36814 , \36813 , \16891 );
nand \U$36438 ( \36815 , \36809 , \36814 );
and \U$36439 ( \36816 , \36806 , \36815 );
and \U$36440 ( \36817 , \36794 , \36805 );
or \U$36441 ( \36818 , \36816 , \36817 );
nand \U$36442 ( \36819 , \36769 , \36818 );
not \U$36443 ( \36820 , \36767 );
nand \U$36444 ( \36821 , \36820 , \36731 );
nand \U$36445 ( \36822 , \36819 , \36821 );
xor \U$36446 ( \36823 , \36695 , \36822 );
xor \U$36447 ( \36824 , \36464 , \36451 );
xor \U$36448 ( \36825 , \36824 , \36441 );
xor \U$36449 ( \36826 , \36396 , \36406 );
xor \U$36450 ( \36827 , \36826 , \36418 );
or \U$36451 ( \36828 , \36825 , \36827 );
xor \U$36452 ( \36829 , \36488 , \36477 );
xor \U$36453 ( \36830 , \36829 , \36529 );
nand \U$36454 ( \36831 , \36828 , \36830 );
nand \U$36455 ( \36832 , \36825 , \36827 );
nand \U$36456 ( \36833 , \36831 , \36832 );
and \U$36457 ( \36834 , \36823 , \36833 );
and \U$36458 ( \36835 , \36695 , \36822 );
or \U$36459 ( \36836 , \36834 , \36835 );
xor \U$36460 ( \36837 , \36693 , \36836 );
not \U$36461 ( \36838 , \9382 );
not \U$36462 ( \36839 , RIc226110_45);
not \U$36463 ( \36840 , \9297 );
or \U$36464 ( \36841 , \36839 , \36840 );
nand \U$36465 ( \36842 , \16998 , \9100 );
nand \U$36466 ( \36843 , \36841 , \36842 );
not \U$36467 ( \36844 , \36843 );
or \U$36468 ( \36845 , \36838 , \36844 );
nand \U$36469 ( \36846 , \36664 , \9398 );
nand \U$36470 ( \36847 , \36845 , \36846 );
not \U$36471 ( \36848 , \9129 );
not \U$36472 ( \36849 , \36703 );
or \U$36473 ( \36850 , \36848 , \36849 );
not \U$36474 ( \36851 , RIc226200_43);
not \U$36475 ( \36852 , \16945 );
or \U$36476 ( \36853 , \36851 , \36852 );
nand \U$36477 ( \36854 , \10086 , \9125 );
nand \U$36478 ( \36855 , \36853 , \36854 );
nand \U$36479 ( \36856 , \36855 , \9110 );
nand \U$36480 ( \36857 , \36850 , \36856 );
or \U$36481 ( \36858 , \36847 , \36857 );
not \U$36482 ( \36859 , RIc225f30_49);
not \U$36483 ( \36860 , \10652 );
or \U$36484 ( \36861 , \36859 , \36860 );
nand \U$36485 ( \36862 , \10653 , \11289 );
nand \U$36486 ( \36863 , \36861 , \36862 );
not \U$36487 ( \36864 , \36863 );
not \U$36488 ( \36865 , \10445 );
or \U$36489 ( \36866 , \36864 , \36865 );
not \U$36490 ( \36867 , \36723 );
nand \U$36491 ( \36868 , \36867 , \9552 );
nand \U$36492 ( \36869 , \36866 , \36868 );
and \U$36493 ( \36870 , \36858 , \36869 );
and \U$36494 ( \36871 , \36847 , \36857 );
nor \U$36495 ( \36872 , \36870 , \36871 );
not \U$36496 ( \36873 , \36728 );
not \U$36497 ( \36874 , \36705 );
and \U$36498 ( \36875 , \36873 , \36874 );
and \U$36499 ( \36876 , \36728 , \36705 );
nor \U$36500 ( \36877 , \36875 , \36876 );
xor \U$36501 ( \36878 , \36877 , \36716 );
xor \U$36502 ( \36879 , \36872 , \36878 );
not \U$36503 ( \36880 , RIc225828_64);
not \U$36504 ( \36881 , \36813 );
or \U$36505 ( \36882 , \36880 , \36881 );
not \U$36506 ( \36883 , RIc2258a0_63);
not \U$36507 ( \36884 , \34276 );
or \U$36508 ( \36885 , \36883 , \36884 );
nand \U$36509 ( \36886 , \22893 , \15620 );
nand \U$36510 ( \36887 , \36885 , \36886 );
nand \U$36511 ( \36888 , \36887 , \16891 );
nand \U$36512 ( \36889 , \36882 , \36888 );
not \U$36513 ( \36890 , \36889 );
not \U$36514 ( \36891 , \11974 );
not \U$36515 ( \36892 , \36712 );
or \U$36516 ( \36893 , \36891 , \36892 );
not \U$36517 ( \36894 , RIc225b70_57);
not \U$36518 ( \36895 , \12724 );
or \U$36519 ( \36896 , \36894 , \36895 );
nand \U$36520 ( \36897 , \8856 , \15262 );
nand \U$36521 ( \36898 , \36896 , \36897 );
nand \U$36522 ( \36899 , \36898 , \11965 );
nand \U$36523 ( \36900 , \36893 , \36899 );
not \U$36524 ( \36901 , \36900 );
nand \U$36525 ( \36902 , \36890 , \36901 );
xor \U$36526 ( \36903 , \36770 , \36780 );
xor \U$36527 ( \36904 , \36903 , \36791 );
and \U$36528 ( \36905 , \36902 , \36904 );
and \U$36529 ( \36906 , \36900 , \36889 );
nor \U$36530 ( \36907 , \36905 , \36906 );
and \U$36531 ( \36908 , \36879 , \36907 );
and \U$36532 ( \36909 , \36872 , \36878 );
or \U$36533 ( \36910 , \36908 , \36909 );
not \U$36534 ( \36911 , \36910 );
xor \U$36535 ( \36912 , \36731 , \36818 );
xor \U$36536 ( \36913 , \36912 , \36767 );
not \U$36537 ( \36914 , \36913 );
or \U$36538 ( \36915 , \36911 , \36914 );
not \U$36539 ( \36916 , \36683 );
not \U$36540 ( \36917 , \36654 );
not \U$36541 ( \36918 , \36917 );
and \U$36542 ( \36919 , \36916 , \36918 );
and \U$36543 ( \36920 , \36683 , \36917 );
nor \U$36544 ( \36921 , \36919 , \36920 );
xor \U$36545 ( \36922 , \36921 , \36656 );
not \U$36546 ( \36923 , \36922 );
nand \U$36547 ( \36924 , \36915 , \36923 );
not \U$36548 ( \36925 , \36913 );
not \U$36549 ( \36926 , \36910 );
nand \U$36550 ( \36927 , \36925 , \36926 );
and \U$36551 ( \36928 , \36924 , \36927 );
not \U$36552 ( \36929 , \36928 );
not \U$36553 ( \36930 , \36929 );
xor \U$36554 ( \36931 , \36695 , \36822 );
xor \U$36555 ( \36932 , \36931 , \36833 );
not \U$36556 ( \36933 , \36932 );
or \U$36557 ( \36934 , \36930 , \36933 );
or \U$36558 ( \36935 , \36932 , \36929 );
xor \U$36559 ( \36936 , \36827 , \36830 );
xnor \U$36560 ( \36937 , \36936 , \36825 );
not \U$36561 ( \36938 , \36937 );
not \U$36562 ( \36939 , \36938 );
xor \U$36563 ( \36940 , \36794 , \36805 );
xor \U$36564 ( \36941 , \36940 , \36815 );
xor \U$36565 ( \36942 , \36505 , \36515 );
xor \U$36566 ( \36943 , \36942 , \36526 );
not \U$36567 ( \36944 , \9444 );
not \U$36568 ( \36945 , \36650 );
or \U$36569 ( \36946 , \36944 , \36945 );
not \U$36570 ( \36947 , RIc225e40_51);
not \U$36571 ( \36948 , \12403 );
or \U$36572 ( \36949 , \36947 , \36948 );
nand \U$36573 ( \36950 , \17744 , \9450 );
nand \U$36574 ( \36951 , \36949 , \36950 );
nand \U$36575 ( \36952 , \36951 , \9458 );
nand \U$36576 ( \36953 , \36946 , \36952 );
xor \U$36577 ( \36954 , \36943 , \36953 );
not \U$36578 ( \36955 , \6307 );
not \U$36579 ( \36956 , \36513 );
or \U$36580 ( \36957 , \36955 , \36956 );
not \U$36581 ( \36958 , RIc2263e0_39);
not \U$36582 ( \36959 , \15444 );
or \U$36583 ( \36960 , \36958 , \36959 );
nand \U$36584 ( \36961 , \12825 , \25483 );
nand \U$36585 ( \36962 , \36960 , \36961 );
nand \U$36586 ( \36963 , \36962 , \6688 );
nand \U$36587 ( \36964 , \36957 , \36963 );
and \U$36588 ( \36965 , \16248 , \4382 );
not \U$36589 ( \36966 , \5519 );
not \U$36590 ( \36967 , \36778 );
or \U$36591 ( \36968 , \36966 , \36967 );
and \U$36592 ( \36969 , RIc2264d0_37, \16256 );
not \U$36593 ( \36970 , RIc2264d0_37);
and \U$36594 ( \36971 , \36970 , \21102 );
nor \U$36595 ( \36972 , \36969 , \36971 );
nand \U$36596 ( \36973 , \36972 , \5508 );
nand \U$36597 ( \36974 , \36968 , \36973 );
xor \U$36598 ( \36975 , \36965 , \36974 );
not \U$36599 ( \36976 , \6306 );
not \U$36600 ( \36977 , \36962 );
or \U$36601 ( \36978 , \36976 , \36977 );
not \U$36602 ( \36979 , RIc2263e0_39);
not \U$36603 ( \36980 , \18158 );
or \U$36604 ( \36981 , \36979 , \36980 );
nand \U$36605 ( \36982 , \15633 , \9573 );
nand \U$36606 ( \36983 , \36981 , \36982 );
nand \U$36607 ( \36984 , \36983 , \6312 );
nand \U$36608 ( \36985 , \36978 , \36984 );
and \U$36609 ( \36986 , \36975 , \36985 );
and \U$36610 ( \36987 , \36965 , \36974 );
or \U$36611 ( \36988 , \36986 , \36987 );
xor \U$36612 ( \36989 , \36964 , \36988 );
not \U$36613 ( \36990 , \10001 );
not \U$36614 ( \36991 , RIc226020_47);
not \U$36615 ( \36992 , \30875 );
or \U$36616 ( \36993 , \36991 , \36992 );
nand \U$36617 ( \36994 , \35479 , \11607 );
nand \U$36618 ( \36995 , \36993 , \36994 );
not \U$36619 ( \36996 , \36995 );
or \U$36620 ( \36997 , \36990 , \36996 );
nand \U$36621 ( \36998 , \36678 , \9619 );
nand \U$36622 ( \36999 , \36997 , \36998 );
and \U$36623 ( \37000 , \36989 , \36999 );
and \U$36624 ( \37001 , \36964 , \36988 );
or \U$36625 ( \37002 , \37000 , \37001 );
xor \U$36626 ( \37003 , \36954 , \37002 );
xor \U$36627 ( \37004 , \36941 , \37003 );
xor \U$36628 ( \37005 , \36743 , \36751 );
xnor \U$36629 ( \37006 , \37005 , \36763 );
and \U$36630 ( \37007 , \37004 , \37006 );
and \U$36631 ( \37008 , \36941 , \37003 );
or \U$36632 ( \37009 , \37007 , \37008 );
not \U$36633 ( \37010 , \37009 );
or \U$36634 ( \37011 , \36939 , \37010 );
or \U$36635 ( \37012 , \37009 , \36938 );
xor \U$36636 ( \37013 , \36943 , \36953 );
and \U$36637 ( \37014 , \37013 , \37002 );
and \U$36638 ( \37015 , \36943 , \36953 );
or \U$36639 ( \37016 , \37014 , \37015 );
not \U$36640 ( \37017 , \37016 );
xor \U$36641 ( \37018 , \36550 , \36566 );
xnor \U$36642 ( \37019 , \37018 , \36561 );
not \U$36643 ( \37020 , \37019 );
and \U$36644 ( \37021 , \37017 , \37020 );
not \U$36645 ( \37022 , \37017 );
and \U$36646 ( \37023 , \37022 , \37019 );
nor \U$36647 ( \37024 , \37021 , \37023 );
xor \U$36648 ( \37025 , \36659 , \36669 );
xor \U$36649 ( \37026 , \37025 , \36680 );
not \U$36650 ( \37027 , \37026 );
not \U$36651 ( \37028 , \9445 );
not \U$36652 ( \37029 , \36951 );
or \U$36653 ( \37030 , \37028 , \37029 );
not \U$36654 ( \37031 , RIc225e40_51);
not \U$36655 ( \37032 , \32810 );
or \U$36656 ( \37033 , \37031 , \37032 );
not \U$36657 ( \37034 , \28026 );
nand \U$36658 ( \37035 , \37034 , \22140 );
nand \U$36659 ( \37036 , \37033 , \37035 );
nand \U$36660 ( \37037 , \37036 , \9459 );
nand \U$36661 ( \37038 , \37030 , \37037 );
not \U$36662 ( \37039 , \12670 );
not \U$36663 ( \37040 , \36746 );
or \U$36664 ( \37041 , \37039 , \37040 );
xnor \U$36665 ( \37042 , RIc225a80_59, \10609 );
nand \U$36666 ( \37043 , \37042 , \15164 );
nand \U$36667 ( \37044 , \37041 , \37043 );
xor \U$36668 ( \37045 , \37038 , \37044 );
not \U$36669 ( \37046 , \11577 );
not \U$36670 ( \37047 , \36759 );
or \U$36671 ( \37048 , \37046 , \37047 );
not \U$36672 ( \37049 , RIc225d50_53);
not \U$36673 ( \37050 , \31855 );
or \U$36674 ( \37051 , \37049 , \37050 );
nand \U$36675 ( \37052 , \11095 , \8782 );
nand \U$36676 ( \37053 , \37051 , \37052 );
nand \U$36677 ( \37054 , \37053 , \9488 );
nand \U$36678 ( \37055 , \37048 , \37054 );
and \U$36679 ( \37056 , \37045 , \37055 );
and \U$36680 ( \37057 , \37038 , \37044 );
or \U$36681 ( \37058 , \37056 , \37057 );
not \U$36682 ( \37059 , \37058 );
or \U$36683 ( \37060 , \37027 , \37059 );
or \U$36684 ( \37061 , \37058 , \37026 );
or \U$36685 ( \37062 , RIc226458_38, RIc2263e0_39);
nand \U$36686 ( \37063 , \37062 , \18357 );
and \U$36687 ( \37064 , RIc226458_38, RIc2263e0_39);
nor \U$36688 ( \37065 , \37064 , \4371 );
and \U$36689 ( \37066 , \37063 , \37065 );
not \U$36690 ( \37067 , \5519 );
not \U$36691 ( \37068 , \36972 );
or \U$36692 ( \37069 , \37067 , \37068 );
and \U$36693 ( \37070 , \21954 , RIc2264d0_37);
and \U$36694 ( \37071 , \16248 , \5504 );
nor \U$36695 ( \37072 , \37070 , \37071 );
or \U$36696 ( \37073 , \37072 , \5507 );
nand \U$36697 ( \37074 , \37069 , \37073 );
and \U$36698 ( \37075 , \37066 , \37074 );
not \U$36699 ( \37076 , \9705 );
not \U$36700 ( \37077 , \36787 );
or \U$36701 ( \37078 , \37076 , \37077 );
not \U$36702 ( \37079 , RIc2262f0_41);
not \U$36703 ( \37080 , \20693 );
or \U$36704 ( \37081 , \37079 , \37080 );
nand \U$36705 ( \37082 , \12755 , \17820 );
nand \U$36706 ( \37083 , \37081 , \37082 );
nand \U$36707 ( \37084 , \37083 , \9690 );
nand \U$36708 ( \37085 , \37078 , \37084 );
xor \U$36709 ( \37086 , \37075 , \37085 );
not \U$36710 ( \37087 , \9129 );
not \U$36711 ( \37088 , \36855 );
or \U$36712 ( \37089 , \37087 , \37088 );
not \U$36713 ( \37090 , RIc226200_43);
not \U$36714 ( \37091 , \20702 );
or \U$36715 ( \37092 , \37090 , \37091 );
nand \U$36716 ( \37093 , \21976 , \9106 );
nand \U$36717 ( \37094 , \37092 , \37093 );
nand \U$36718 ( \37095 , \37094 , \9110 );
nand \U$36719 ( \37096 , \37089 , \37095 );
and \U$36720 ( \37097 , \37086 , \37096 );
and \U$36721 ( \37098 , \37075 , \37085 );
or \U$36722 ( \37099 , \37097 , \37098 );
not \U$36723 ( \37100 , \15729 );
not \U$36724 ( \37101 , \36803 );
or \U$36725 ( \37102 , \37100 , \37101 );
not \U$36726 ( \37103 , RIc225990_61);
not \U$36727 ( \37104 , \10125 );
or \U$36728 ( \37105 , \37103 , \37104 );
nand \U$36729 ( \37106 , \27798 , \12806 );
nand \U$36730 ( \37107 , \37105 , \37106 );
nand \U$36731 ( \37108 , \37107 , \15719 );
nand \U$36732 ( \37109 , \37102 , \37108 );
xor \U$36733 ( \37110 , \37099 , \37109 );
not \U$36734 ( \37111 , \12532 );
not \U$36735 ( \37112 , \36741 );
or \U$36736 ( \37113 , \37111 , \37112 );
not \U$36737 ( \37114 , RIc225c60_55);
not \U$36738 ( \37115 , \8810 );
or \U$36739 ( \37116 , \37114 , \37115 );
nand \U$36740 ( \37117 , \8811 , \11041 );
nand \U$36741 ( \37118 , \37116 , \37117 );
nand \U$36742 ( \37119 , \37118 , \11118 );
nand \U$36743 ( \37120 , \37113 , \37119 );
and \U$36744 ( \37121 , \37110 , \37120 );
and \U$36745 ( \37122 , \37099 , \37109 );
or \U$36746 ( \37123 , \37121 , \37122 );
nand \U$36747 ( \37124 , \37061 , \37123 );
nand \U$36748 ( \37125 , \37060 , \37124 );
xor \U$36749 ( \37126 , \37024 , \37125 );
nand \U$36750 ( \37127 , \37012 , \37126 );
nand \U$36751 ( \37128 , \37011 , \37127 );
nand \U$36752 ( \37129 , \36935 , \37128 );
nand \U$36753 ( \37130 , \36934 , \37129 );
xor \U$36754 ( \37131 , \36837 , \37130 );
xor \U$36755 ( \37132 , \36337 , \36427 );
xor \U$36756 ( \37133 , \37132 , \36534 );
xor \U$36757 ( \37134 , \36540 , \36577 );
xor \U$36758 ( \37135 , \37134 , \36580 );
xor \U$36759 ( \37136 , \37133 , \37135 );
xor \U$36760 ( \37137 , \36569 , \36571 );
xor \U$36761 ( \37138 , \37137 , \36574 );
xor \U$36762 ( \37139 , \36644 , \36686 );
xor \U$36763 ( \37140 , \37139 , \36689 );
xor \U$36764 ( \37141 , \37138 , \37140 );
nand \U$36765 ( \37142 , \37017 , \37020 );
not \U$36766 ( \37143 , \37142 );
not \U$36767 ( \37144 , \37125 );
or \U$36768 ( \37145 , \37143 , \37144 );
nand \U$36769 ( \37146 , \37016 , \37019 );
nand \U$36770 ( \37147 , \37145 , \37146 );
and \U$36771 ( \37148 , \37141 , \37147 );
and \U$36772 ( \37149 , \37138 , \37140 );
or \U$36773 ( \37150 , \37148 , \37149 );
xor \U$36774 ( \37151 , \37136 , \37150 );
xor \U$36775 ( \37152 , \37131 , \37151 );
not \U$36776 ( \37153 , \36932 );
not \U$36777 ( \37154 , \36928 );
or \U$36778 ( \37155 , \37153 , \37154 );
or \U$36779 ( \37156 , \36928 , \36932 );
nand \U$36780 ( \37157 , \37155 , \37156 );
and \U$36781 ( \37158 , \37157 , \37128 );
not \U$36782 ( \37159 , \37157 );
not \U$36783 ( \37160 , \37128 );
and \U$36784 ( \37161 , \37159 , \37160 );
nor \U$36785 ( \37162 , \37158 , \37161 );
not \U$36786 ( \37163 , \37162 );
xor \U$36787 ( \37164 , \37138 , \37140 );
xor \U$36788 ( \37165 , \37164 , \37147 );
not \U$36789 ( \37166 , \37165 );
xor \U$36790 ( \37167 , \36847 , \36857 );
and \U$36791 ( \37168 , \37167 , \36869 );
not \U$36792 ( \37169 , \37167 );
not \U$36793 ( \37170 , \36869 );
and \U$36794 ( \37171 , \37169 , \37170 );
nor \U$36795 ( \37172 , \37168 , \37171 );
not \U$36796 ( \37173 , \37172 );
not \U$36797 ( \37174 , RIc225828_64);
not \U$36798 ( \37175 , \36887 );
or \U$36799 ( \37176 , \37174 , \37175 );
and \U$36800 ( \37177 , RIc2258a0_63, \9765 );
not \U$36801 ( \37178 , RIc2258a0_63);
and \U$36802 ( \37179 , \37178 , \34821 );
or \U$36803 ( \37180 , \37177 , \37179 );
nand \U$36804 ( \37181 , \37180 , \16891 );
nand \U$36805 ( \37182 , \37176 , \37181 );
not \U$36806 ( \37183 , \37182 );
not \U$36807 ( \37184 , \12670 );
not \U$36808 ( \37185 , \37042 );
or \U$36809 ( \37186 , \37184 , \37185 );
and \U$36810 ( \37187 , RIc225a80_59, \8887 );
not \U$36811 ( \37188 , RIc225a80_59);
and \U$36812 ( \37189 , \37188 , \17582 );
or \U$36813 ( \37190 , \37187 , \37189 );
nand \U$36814 ( \37191 , \37190 , \15164 );
nand \U$36815 ( \37192 , \37186 , \37191 );
not \U$36816 ( \37193 , \37192 );
or \U$36817 ( \37194 , \37183 , \37193 );
or \U$36818 ( \37195 , \37192 , \37182 );
not \U$36819 ( \37196 , \8788 );
not \U$36820 ( \37197 , \37053 );
or \U$36821 ( \37198 , \37196 , \37197 );
not \U$36822 ( \37199 , RIc225d50_53);
not \U$36823 ( \37200 , \8910 );
or \U$36824 ( \37201 , \37199 , \37200 );
nand \U$36825 ( \37202 , \34363 , \8782 );
nand \U$36826 ( \37203 , \37201 , \37202 );
nand \U$36827 ( \37204 , \37203 , \9488 );
nand \U$36828 ( \37205 , \37198 , \37204 );
nand \U$36829 ( \37206 , \37195 , \37205 );
nand \U$36830 ( \37207 , \37194 , \37206 );
not \U$36831 ( \37208 , \37207 );
or \U$36832 ( \37209 , \37173 , \37208 );
or \U$36833 ( \37210 , \37207 , \37172 );
not \U$36834 ( \37211 , \9934 );
not \U$36835 ( \37212 , RIc226110_45);
not \U$36836 ( \37213 , \12100 );
or \U$36837 ( \37214 , \37212 , \37213 );
nand \U$36838 ( \37215 , \9324 , \14390 );
nand \U$36839 ( \37216 , \37214 , \37215 );
not \U$36840 ( \37217 , \37216 );
or \U$36841 ( \37218 , \37211 , \37217 );
nand \U$36842 ( \37219 , \36843 , \9398 );
nand \U$36843 ( \37220 , \37218 , \37219 );
not \U$36844 ( \37221 , \9552 );
not \U$36845 ( \37222 , \36863 );
or \U$36846 ( \37223 , \37221 , \37222 );
not \U$36847 ( \37224 , RIc225f30_49);
not \U$36848 ( \37225 , \10111 );
or \U$36849 ( \37226 , \37224 , \37225 );
nand \U$36850 ( \37227 , \10110 , \9549 );
nand \U$36851 ( \37228 , \37226 , \37227 );
nand \U$36852 ( \37229 , \9532 , \37228 );
nand \U$36853 ( \37230 , \37223 , \37229 );
xor \U$36854 ( \37231 , \37220 , \37230 );
not \U$36855 ( \37232 , \11974 );
not \U$36856 ( \37233 , \36898 );
or \U$36857 ( \37234 , \37232 , \37233 );
not \U$36858 ( \37235 , RIc225b70_57);
not \U$36859 ( \37236 , \20217 );
or \U$36860 ( \37237 , \37235 , \37236 );
nand \U$36861 ( \37238 , \22969 , \11033 );
nand \U$36862 ( \37239 , \37237 , \37238 );
nand \U$36863 ( \37240 , \37239 , \11965 );
nand \U$36864 ( \37241 , \37234 , \37240 );
and \U$36865 ( \37242 , \37231 , \37241 );
and \U$36866 ( \37243 , \37220 , \37230 );
or \U$36867 ( \37244 , \37242 , \37243 );
nand \U$36868 ( \37245 , \37210 , \37244 );
nand \U$36869 ( \37246 , \37209 , \37245 );
not \U$36870 ( \37247 , \37246 );
xor \U$36871 ( \37248 , \37066 , \37074 );
not \U$36872 ( \37249 , \6307 );
not \U$36873 ( \37250 , \36983 );
or \U$36874 ( \37251 , \37249 , \37250 );
and \U$36875 ( \37252 , \8990 , \21094 );
not \U$36876 ( \37253 , \8990 );
and \U$36877 ( \37254 , \37253 , \20393 );
nor \U$36878 ( \37255 , \37252 , \37254 );
nand \U$36879 ( \37256 , \37255 , \6312 );
nand \U$36880 ( \37257 , \37251 , \37256 );
xor \U$36881 ( \37258 , \37248 , \37257 );
not \U$36882 ( \37259 , \9705 );
not \U$36883 ( \37260 , \37083 );
or \U$36884 ( \37261 , \37259 , \37260 );
not \U$36885 ( \37262 , RIc2262f0_41);
not \U$36886 ( \37263 , \18167 );
or \U$36887 ( \37264 , \37262 , \37263 );
nand \U$36888 ( \37265 , \19721 , \6303 );
nand \U$36889 ( \37266 , \37264 , \37265 );
nand \U$36890 ( \37267 , \37266 , \9690 );
nand \U$36891 ( \37268 , \37261 , \37267 );
and \U$36892 ( \37269 , \37258 , \37268 );
and \U$36893 ( \37270 , \37248 , \37257 );
or \U$36894 ( \37271 , \37269 , \37270 );
not \U$36895 ( \37272 , \15719 );
not \U$36896 ( \37273 , RIc225990_61);
not \U$36897 ( \37274 , \6719 );
or \U$36898 ( \37275 , \37273 , \37274 );
nand \U$36899 ( \37276 , \6720 , \10338 );
nand \U$36900 ( \37277 , \37275 , \37276 );
not \U$36901 ( \37278 , \37277 );
or \U$36902 ( \37279 , \37272 , \37278 );
nand \U$36903 ( \37280 , \37107 , \15729 );
nand \U$36904 ( \37281 , \37279 , \37280 );
xor \U$36905 ( \37282 , \37271 , \37281 );
not \U$36906 ( \37283 , \12532 );
not \U$36907 ( \37284 , \37118 );
or \U$36908 ( \37285 , \37283 , \37284 );
not \U$36909 ( \37286 , RIc225c60_55);
not \U$36910 ( \37287 , \20367 );
or \U$36911 ( \37288 , \37286 , \37287 );
nand \U$36912 ( \37289 , \8952 , \11108 );
nand \U$36913 ( \37290 , \37288 , \37289 );
nand \U$36914 ( \37291 , \37290 , \11117 );
nand \U$36915 ( \37292 , \37285 , \37291 );
and \U$36916 ( \37293 , \37282 , \37292 );
and \U$36917 ( \37294 , \37271 , \37281 );
or \U$36918 ( \37295 , \37293 , \37294 );
not \U$36919 ( \37296 , \37295 );
xor \U$36920 ( \37297 , \36965 , \36974 );
xor \U$36921 ( \37298 , \37297 , \36985 );
not \U$36922 ( \37299 , \9641 );
not \U$36923 ( \37300 , RIc226020_47);
not \U$36924 ( \37301 , \21156 );
or \U$36925 ( \37302 , \37300 , \37301 );
nand \U$36926 ( \37303 , \10976 , \11607 );
nand \U$36927 ( \37304 , \37302 , \37303 );
not \U$36928 ( \37305 , \37304 );
or \U$36929 ( \37306 , \37299 , \37305 );
nand \U$36930 ( \37307 , \36995 , \9619 );
nand \U$36931 ( \37308 , \37306 , \37307 );
xor \U$36932 ( \37309 , \37298 , \37308 );
not \U$36933 ( \37310 , \9445 );
not \U$36934 ( \37311 , \37036 );
or \U$36935 ( \37312 , \37310 , \37311 );
not \U$36936 ( \37313 , RIc225e40_51);
not \U$36937 ( \37314 , \13465 );
or \U$36938 ( \37315 , \37313 , \37314 );
nand \U$36939 ( \37316 , \9051 , \11795 );
nand \U$36940 ( \37317 , \37315 , \37316 );
nand \U$36941 ( \37318 , \37317 , \9459 );
nand \U$36942 ( \37319 , \37312 , \37318 );
and \U$36943 ( \37320 , \37309 , \37319 );
and \U$36944 ( \37321 , \37298 , \37308 );
or \U$36945 ( \37322 , \37320 , \37321 );
not \U$36946 ( \37323 , \37322 );
xor \U$36947 ( \37324 , \36964 , \36988 );
xor \U$36948 ( \37325 , \37324 , \36999 );
not \U$36949 ( \37326 , \37325 );
nand \U$36950 ( \37327 , \37323 , \37326 );
not \U$36951 ( \37328 , \37327 );
or \U$36952 ( \37329 , \37296 , \37328 );
not \U$36953 ( \37330 , \37326 );
nand \U$36954 ( \37331 , \37330 , \37322 );
nand \U$36955 ( \37332 , \37329 , \37331 );
not \U$36956 ( \37333 , \37332 );
nand \U$36957 ( \37334 , \37247 , \37333 );
xor \U$36958 ( \37335 , \37026 , \37123 );
xnor \U$36959 ( \37336 , \37335 , \37058 );
not \U$36960 ( \37337 , \37336 );
and \U$36961 ( \37338 , \37334 , \37337 );
nor \U$36962 ( \37339 , \37247 , \37333 );
nor \U$36963 ( \37340 , \37338 , \37339 );
not \U$36964 ( \37341 , \37340 );
not \U$36965 ( \37342 , \37341 );
xor \U$36966 ( \37343 , \36872 , \36878 );
xor \U$36967 ( \37344 , \37343 , \36907 );
not \U$36968 ( \37345 , \37344 );
not \U$36969 ( \37346 , \37345 );
xor \U$36970 ( \37347 , \37038 , \37044 );
xor \U$36971 ( \37348 , \37347 , \37055 );
xor \U$36972 ( \37349 , \37099 , \37109 );
xor \U$36973 ( \37350 , \37349 , \37120 );
or \U$36974 ( \37351 , \37348 , \37350 );
xor \U$36975 ( \37352 , \36904 , \36889 );
xnor \U$36976 ( \37353 , \37352 , \36901 );
and \U$36977 ( \37354 , \37351 , \37353 );
and \U$36978 ( \37355 , \37350 , \37348 );
nor \U$36979 ( \37356 , \37354 , \37355 );
not \U$36980 ( \37357 , \37356 );
not \U$36981 ( \37358 , \37357 );
or \U$36982 ( \37359 , \37346 , \37358 );
xor \U$36983 ( \37360 , \36941 , \37003 );
xor \U$36984 ( \37361 , \37360 , \37006 );
nand \U$36985 ( \37362 , \37356 , \37344 );
nand \U$36986 ( \37363 , \37361 , \37362 );
nand \U$36987 ( \37364 , \37359 , \37363 );
not \U$36988 ( \37365 , \37364 );
or \U$36989 ( \37366 , \37342 , \37365 );
not \U$36990 ( \37367 , \37364 );
not \U$36991 ( \37368 , \37367 );
not \U$36992 ( \37369 , \37340 );
or \U$36993 ( \37370 , \37368 , \37369 );
xor \U$36994 ( \37371 , \36922 , \36926 );
xnor \U$36995 ( \37372 , \37371 , \36925 );
nand \U$36996 ( \37373 , \37370 , \37372 );
nand \U$36997 ( \37374 , \37366 , \37373 );
not \U$36998 ( \37375 , \37374 );
nand \U$36999 ( \37376 , \37166 , \37375 );
not \U$37000 ( \37377 , \37376 );
or \U$37001 ( \37378 , \37163 , \37377 );
nand \U$37002 ( \37379 , \37374 , \37165 );
nand \U$37003 ( \37380 , \37378 , \37379 );
nand \U$37004 ( \37381 , \37152 , \37380 );
not \U$37005 ( \37382 , \37381 );
not \U$37006 ( \37383 , \37375 );
not \U$37007 ( \37384 , \37165 );
or \U$37008 ( \37385 , \37383 , \37384 );
or \U$37009 ( \37386 , \37375 , \37165 );
nand \U$37010 ( \37387 , \37385 , \37386 );
xor \U$37011 ( \37388 , \37387 , \37162 );
xor \U$37012 ( \37389 , \37075 , \37085 );
xor \U$37013 ( \37390 , \37389 , \37096 );
not \U$37014 ( \37391 , \9129 );
not \U$37015 ( \37392 , \37094 );
or \U$37016 ( \37393 , \37391 , \37392 );
not \U$37017 ( \37394 , RIc226200_43);
not \U$37018 ( \37395 , \13498 );
or \U$37019 ( \37396 , \37394 , \37395 );
not \U$37020 ( \37397 , \21084 );
nand \U$37021 ( \37398 , \37397 , \9125 );
nand \U$37022 ( \37399 , \37396 , \37398 );
nand \U$37023 ( \37400 , \37399 , \9110 );
nand \U$37024 ( \37401 , \37393 , \37400 );
and \U$37025 ( \37402 , \16248 , \5519 );
not \U$37026 ( \37403 , \6306 );
not \U$37027 ( \37404 , \37255 );
or \U$37028 ( \37405 , \37403 , \37404 );
and \U$37029 ( \37406 , RIc2263e0_39, \16482 );
not \U$37030 ( \37407 , RIc2263e0_39);
and \U$37031 ( \37408 , \37407 , \21102 );
nor \U$37032 ( \37409 , \37406 , \37408 );
nand \U$37033 ( \37410 , \37409 , \6312 );
nand \U$37034 ( \37411 , \37405 , \37410 );
xor \U$37035 ( \37412 , \37402 , \37411 );
not \U$37036 ( \37413 , \9689 );
not \U$37037 ( \37414 , RIc2262f0_41);
not \U$37038 ( \37415 , \12846 );
or \U$37039 ( \37416 , \37414 , \37415 );
nand \U$37040 ( \37417 , \12845 , \6303 );
nand \U$37041 ( \37418 , \37416 , \37417 );
not \U$37042 ( \37419 , \37418 );
or \U$37043 ( \37420 , \37413 , \37419 );
nand \U$37044 ( \37421 , \37266 , \9705 );
nand \U$37045 ( \37422 , \37420 , \37421 );
and \U$37046 ( \37423 , \37412 , \37422 );
and \U$37047 ( \37424 , \37402 , \37411 );
or \U$37048 ( \37425 , \37423 , \37424 );
xor \U$37049 ( \37426 , \37401 , \37425 );
not \U$37050 ( \37427 , \9444 );
not \U$37051 ( \37428 , \37317 );
or \U$37052 ( \37429 , \37427 , \37428 );
not \U$37053 ( \37430 , RIc225e40_51);
not \U$37054 ( \37431 , \9073 );
or \U$37055 ( \37432 , \37430 , \37431 );
nand \U$37056 ( \37433 , \9072 , \12423 );
nand \U$37057 ( \37434 , \37432 , \37433 );
nand \U$37058 ( \37435 , \37434 , \9458 );
nand \U$37059 ( \37436 , \37429 , \37435 );
and \U$37060 ( \37437 , \37426 , \37436 );
and \U$37061 ( \37438 , \37401 , \37425 );
or \U$37062 ( \37439 , \37437 , \37438 );
xor \U$37063 ( \37440 , \37390 , \37439 );
not \U$37064 ( \37441 , \9398 );
not \U$37065 ( \37442 , \37216 );
or \U$37066 ( \37443 , \37441 , \37442 );
not \U$37067 ( \37444 , RIc226110_45);
not \U$37068 ( \37445 , \16945 );
or \U$37069 ( \37446 , \37444 , \37445 );
nand \U$37070 ( \37447 , \10086 , \9379 );
nand \U$37071 ( \37448 , \37446 , \37447 );
nand \U$37072 ( \37449 , \37448 , \9382 );
nand \U$37073 ( \37450 , \37443 , \37449 );
not \U$37074 ( \37451 , \9534 );
not \U$37075 ( \37452 , RIc225f30_49);
not \U$37076 ( \37453 , \9250 );
or \U$37077 ( \37454 , \37452 , \37453 );
nand \U$37078 ( \37455 , \9256 , \11289 );
nand \U$37079 ( \37456 , \37454 , \37455 );
not \U$37080 ( \37457 , \37456 );
or \U$37081 ( \37458 , \37451 , \37457 );
nand \U$37082 ( \37459 , \9552 , \37228 );
nand \U$37083 ( \37460 , \37458 , \37459 );
xor \U$37084 ( \37461 , \37450 , \37460 );
not \U$37085 ( \37462 , \10001 );
not \U$37086 ( \37463 , RIc226020_47);
not \U$37087 ( \37464 , \9300 );
or \U$37088 ( \37465 , \37463 , \37464 );
nand \U$37089 ( \37466 , \9299 , \9624 );
nand \U$37090 ( \37467 , \37465 , \37466 );
not \U$37091 ( \37468 , \37467 );
or \U$37092 ( \37469 , \37462 , \37468 );
nand \U$37093 ( \37470 , \37304 , \9619 );
nand \U$37094 ( \37471 , \37469 , \37470 );
and \U$37095 ( \37472 , \37461 , \37471 );
and \U$37096 ( \37473 , \37450 , \37460 );
or \U$37097 ( \37474 , \37472 , \37473 );
and \U$37098 ( \37475 , \37440 , \37474 );
and \U$37099 ( \37476 , \37390 , \37439 );
or \U$37100 ( \37477 , \37475 , \37476 );
xor \U$37101 ( \37478 , \37220 , \37230 );
xor \U$37102 ( \37479 , \37478 , \37241 );
not \U$37103 ( \37480 , \9555 );
not \U$37104 ( \37481 , \37203 );
or \U$37105 ( \37482 , \37480 , \37481 );
and \U$37106 ( \37483 , RIc225d50_53, \9211 );
not \U$37107 ( \37484 , RIc225d50_53);
and \U$37108 ( \37485 , \37484 , \8925 );
nor \U$37109 ( \37486 , \37483 , \37485 );
nand \U$37110 ( \37487 , \37486 , \8777 );
nand \U$37111 ( \37488 , \37482 , \37487 );
not \U$37112 ( \37489 , \37488 );
not \U$37113 ( \37490 , \16891 );
not \U$37114 ( \37491 , RIc2258a0_63);
not \U$37115 ( \37492 , \6493 );
or \U$37116 ( \37493 , \37491 , \37492 );
not \U$37117 ( \37494 , RIc2258a0_63);
nand \U$37118 ( \37495 , \6494 , \37494 );
nand \U$37119 ( \37496 , \37493 , \37495 );
not \U$37120 ( \37497 , \37496 );
or \U$37121 ( \37498 , \37490 , \37497 );
nand \U$37122 ( \37499 , \37180 , RIc225828_64);
nand \U$37123 ( \37500 , \37498 , \37499 );
not \U$37124 ( \37501 , \37500 );
or \U$37125 ( \37502 , \37489 , \37501 );
or \U$37126 ( \37503 , \37500 , \37488 );
not \U$37127 ( \37504 , \13025 );
not \U$37128 ( \37505 , \37290 );
or \U$37129 ( \37506 , \37504 , \37505 );
and \U$37130 ( \37507 , \8975 , RIc225c60_55);
not \U$37131 ( \37508 , \8975 );
and \U$37132 ( \37509 , \37508 , \11108 );
or \U$37133 ( \37510 , \37507 , \37509 );
nand \U$37134 ( \37511 , \37510 , \11117 );
nand \U$37135 ( \37512 , \37506 , \37511 );
nand \U$37136 ( \37513 , \37503 , \37512 );
nand \U$37137 ( \37514 , \37502 , \37513 );
xor \U$37138 ( \37515 , \37479 , \37514 );
not \U$37139 ( \37516 , \11965 );
not \U$37140 ( \37517 , RIc225b70_57);
not \U$37141 ( \37518 , \10858 );
or \U$37142 ( \37519 , \37517 , \37518 );
nand \U$37143 ( \37520 , \23042 , \11033 );
nand \U$37144 ( \37521 , \37519 , \37520 );
not \U$37145 ( \37522 , \37521 );
or \U$37146 ( \37523 , \37516 , \37522 );
nand \U$37147 ( \37524 , \37239 , \11974 );
nand \U$37148 ( \37525 , \37523 , \37524 );
or \U$37149 ( \37526 , RIc226368_40, RIc2262f0_41);
nand \U$37150 ( \37527 , \37526 , \18357 );
and \U$37151 ( \37528 , RIc226368_40, RIc2262f0_41);
nor \U$37152 ( \37529 , \37528 , \8998 );
and \U$37153 ( \37530 , \37527 , \37529 );
not \U$37154 ( \37531 , \6306 );
not \U$37155 ( \37532 , \37409 );
or \U$37156 ( \37533 , \37531 , \37532 );
and \U$37157 ( \37534 , RIc2263e0_39, \16248 );
not \U$37158 ( \37535 , RIc2263e0_39);
and \U$37159 ( \37536 , \37535 , \18181 );
nor \U$37160 ( \37537 , \37534 , \37536 );
nand \U$37161 ( \37538 , \37537 , \6312 );
nand \U$37162 ( \37539 , \37533 , \37538 );
and \U$37163 ( \37540 , \37530 , \37539 );
not \U$37164 ( \37541 , \9110 );
not \U$37165 ( \37542 , RIc226200_43);
not \U$37166 ( \37543 , \13198 );
or \U$37167 ( \37544 , \37542 , \37543 );
nand \U$37168 ( \37545 , \12755 , \9117 );
nand \U$37169 ( \37546 , \37544 , \37545 );
not \U$37170 ( \37547 , \37546 );
or \U$37171 ( \37548 , \37541 , \37547 );
nand \U$37172 ( \37549 , \37399 , \9128 );
nand \U$37173 ( \37550 , \37548 , \37549 );
xor \U$37174 ( \37551 , \37540 , \37550 );
not \U$37175 ( \37552 , \9398 );
not \U$37176 ( \37553 , \37448 );
or \U$37177 ( \37554 , \37552 , \37553 );
not \U$37178 ( \37555 , RIc226110_45);
not \U$37179 ( \37556 , \10198 );
or \U$37180 ( \37557 , \37555 , \37556 );
not \U$37181 ( \37558 , \13211 );
nand \U$37182 ( \37559 , \37558 , \9100 );
nand \U$37183 ( \37560 , \37557 , \37559 );
nand \U$37184 ( \37561 , \37560 , \9934 );
nand \U$37185 ( \37562 , \37554 , \37561 );
and \U$37186 ( \37563 , \37551 , \37562 );
and \U$37187 ( \37564 , \37540 , \37550 );
or \U$37188 ( \37565 , \37563 , \37564 );
xor \U$37189 ( \37566 , \37525 , \37565 );
not \U$37190 ( \37567 , \15729 );
not \U$37191 ( \37568 , \37277 );
or \U$37192 ( \37569 , \37567 , \37568 );
not \U$37193 ( \37570 , RIc225990_61);
not \U$37194 ( \37571 , \15699 );
or \U$37195 ( \37572 , \37570 , \37571 );
nand \U$37196 ( \37573 , \10310 , \10338 );
nand \U$37197 ( \37574 , \37572 , \37573 );
nand \U$37198 ( \37575 , \37574 , \15719 );
nand \U$37199 ( \37576 , \37569 , \37575 );
and \U$37200 ( \37577 , \37566 , \37576 );
and \U$37201 ( \37578 , \37525 , \37565 );
or \U$37202 ( \37579 , \37577 , \37578 );
and \U$37203 ( \37580 , \37515 , \37579 );
and \U$37204 ( \37581 , \37479 , \37514 );
or \U$37205 ( \37582 , \37580 , \37581 );
xor \U$37206 ( \37583 , \37477 , \37582 );
and \U$37207 ( \37584 , \37322 , \37325 );
not \U$37208 ( \37585 , \37322 );
and \U$37209 ( \37586 , \37585 , \37326 );
nor \U$37210 ( \37587 , \37584 , \37586 );
xor \U$37211 ( \37588 , \37587 , \37295 );
and \U$37212 ( \37589 , \37583 , \37588 );
and \U$37213 ( \37590 , \37477 , \37582 );
or \U$37214 ( \37591 , \37589 , \37590 );
not \U$37215 ( \37592 , \37591 );
xor \U$37216 ( \37593 , \37332 , \37246 );
xnor \U$37217 ( \37594 , \37593 , \37336 );
not \U$37218 ( \37595 , \37594 );
or \U$37219 ( \37596 , \37592 , \37595 );
or \U$37220 ( \37597 , \37591 , \37594 );
xor \U$37221 ( \37598 , \37172 , \37244 );
xnor \U$37222 ( \37599 , \37598 , \37207 );
not \U$37223 ( \37600 , \37599 );
not \U$37224 ( \37601 , \37600 );
xor \U$37225 ( \37602 , \37350 , \37348 );
xor \U$37226 ( \37603 , \37602 , \37353 );
not \U$37227 ( \37604 , \37603 );
or \U$37228 ( \37605 , \37601 , \37604 );
or \U$37229 ( \37606 , \37603 , \37600 );
xor \U$37230 ( \37607 , \37298 , \37308 );
xor \U$37231 ( \37608 , \37607 , \37319 );
not \U$37232 ( \37609 , \37608 );
xor \U$37233 ( \37610 , \37182 , \37192 );
not \U$37234 ( \37611 , \37205 );
and \U$37235 ( \37612 , \37610 , \37611 );
not \U$37236 ( \37613 , \37610 );
and \U$37237 ( \37614 , \37613 , \37205 );
nor \U$37238 ( \37615 , \37612 , \37614 );
nand \U$37239 ( \37616 , \37609 , \37615 );
xor \U$37240 ( \37617 , \37271 , \37281 );
xor \U$37241 ( \37618 , \37617 , \37292 );
and \U$37242 ( \37619 , \37616 , \37618 );
not \U$37243 ( \37620 , \37608 );
nor \U$37244 ( \37621 , \37620 , \37615 );
nor \U$37245 ( \37622 , \37619 , \37621 );
not \U$37246 ( \37623 , \37622 );
nand \U$37247 ( \37624 , \37606 , \37623 );
nand \U$37248 ( \37625 , \37605 , \37624 );
nand \U$37249 ( \37626 , \37597 , \37625 );
nand \U$37250 ( \37627 , \37596 , \37626 );
and \U$37251 ( \37628 , \37009 , \36938 );
not \U$37252 ( \37629 , \37009 );
and \U$37253 ( \37630 , \37629 , \36937 );
nor \U$37254 ( \37631 , \37628 , \37630 );
xor \U$37255 ( \37632 , \37631 , \37126 );
or \U$37256 ( \37633 , \37627 , \37632 );
xor \U$37257 ( \37634 , \37364 , \37341 );
xor \U$37258 ( \37635 , \37634 , \37372 );
nand \U$37259 ( \37636 , \37633 , \37635 );
nand \U$37260 ( \37637 , \37627 , \37632 );
nand \U$37261 ( \37638 , \37636 , \37637 );
nand \U$37262 ( \37639 , \37388 , \37638 );
not \U$37263 ( \37640 , \37639 );
or \U$37264 ( \37641 , \37382 , \37640 );
or \U$37265 ( \37642 , \37152 , \37380 );
nand \U$37266 ( \37643 , \37641 , \37642 );
xor \U$37267 ( \37644 , \36642 , \36692 );
and \U$37268 ( \37645 , \37644 , \36836 );
and \U$37269 ( \37646 , \36642 , \36692 );
or \U$37270 ( \37647 , \37645 , \37646 );
xor \U$37271 ( \37648 , \37133 , \37135 );
and \U$37272 ( \37649 , \37648 , \37150 );
and \U$37273 ( \37650 , \37133 , \37135 );
or \U$37274 ( \37651 , \37649 , \37650 );
xor \U$37275 ( \37652 , \37647 , \37651 );
and \U$37276 ( \37653 , \36604 , \36607 );
not \U$37277 ( \37654 , \36604 );
and \U$37278 ( \37655 , \37654 , \36608 );
nor \U$37279 ( \37656 , \37653 , \37655 );
and \U$37280 ( \37657 , \37656 , \36612 );
not \U$37281 ( \37658 , \37656 );
not \U$37282 ( \37659 , \36612 );
and \U$37283 ( \37660 , \37658 , \37659 );
nor \U$37284 ( \37661 , \37657 , \37660 );
xor \U$37285 ( \37662 , \37652 , \37661 );
xor \U$37286 ( \37663 , \36837 , \37130 );
and \U$37287 ( \37664 , \37663 , \37151 );
and \U$37288 ( \37665 , \36837 , \37130 );
or \U$37289 ( \37666 , \37664 , \37665 );
nor \U$37290 ( \37667 , \37662 , \37666 );
or \U$37291 ( \37668 , \37643 , \37667 );
nand \U$37292 ( \37669 , \37662 , \37666 );
nand \U$37293 ( \37670 , \37668 , \37669 );
xor \U$37294 ( \37671 , \36602 , \36616 );
xor \U$37295 ( \37672 , \37671 , \36619 );
not \U$37296 ( \37673 , \37672 );
xor \U$37297 ( \37674 , \37647 , \37651 );
and \U$37298 ( \37675 , \37674 , \37661 );
and \U$37299 ( \37676 , \37647 , \37651 );
or \U$37300 ( \37677 , \37675 , \37676 );
not \U$37301 ( \37678 , \37677 );
nand \U$37302 ( \37679 , \37673 , \37678 );
and \U$37303 ( \37680 , \37670 , \37679 );
not \U$37304 ( \37681 , \37672 );
nor \U$37305 ( \37682 , \37681 , \37678 );
nor \U$37306 ( \37683 , \37680 , \37682 );
nor \U$37307 ( \37684 , \36640 , \37683 );
nor \U$37308 ( \37685 , \36634 , \37684 );
xor \U$37309 ( \37686 , \32578 , \32606 );
xor \U$37310 ( \37687 , \37686 , \32618 );
xor \U$37311 ( \37688 , \32580 , \32592 );
xor \U$37312 ( \37689 , \37688 , \32603 );
not \U$37313 ( \37690 , \3631 );
not \U$37314 ( \37691 , \32675 );
or \U$37315 ( \37692 , \37690 , \37691 );
nand \U$37316 ( \37693 , \34581 , \3629 );
nand \U$37317 ( \37694 , \37692 , \37693 );
xor \U$37318 ( \37695 , \37689 , \37694 );
not \U$37319 ( \37696 , \6307 );
not \U$37320 ( \37697 , \32815 );
or \U$37321 ( \37698 , \37696 , \37697 );
nand \U$37322 ( \37699 , \35729 , \6689 );
nand \U$37323 ( \37700 , \37698 , \37699 );
and \U$37324 ( \37701 , \37695 , \37700 );
and \U$37325 ( \37702 , \37689 , \37694 );
or \U$37326 ( \37703 , \37701 , \37702 );
xor \U$37327 ( \37704 , \37687 , \37703 );
not \U$37328 ( \37705 , \32694 );
not \U$37329 ( \37706 , \32680 );
or \U$37330 ( \37707 , \37705 , \37706 );
nand \U$37331 ( \37708 , \32679 , \32668 );
nand \U$37332 ( \37709 , \37707 , \37708 );
xnor \U$37333 ( \37710 , \37709 , \32692 );
xor \U$37334 ( \37711 , \37704 , \37710 );
not \U$37335 ( \37712 , \5135 );
not \U$37336 ( \37713 , \32688 );
or \U$37337 ( \37714 , \37712 , \37713 );
nand \U$37338 ( \37715 , \34606 , \5741 );
nand \U$37339 ( \37716 , \37714 , \37715 );
not \U$37340 ( \37717 , \5519 );
not \U$37341 ( \37718 , \32614 );
or \U$37342 ( \37719 , \37717 , \37718 );
nand \U$37343 ( \37720 , \34597 , \5509 );
nand \U$37344 ( \37721 , \37719 , \37720 );
xor \U$37345 ( \37722 , \37716 , \37721 );
not \U$37346 ( \37723 , \9534 );
not \U$37347 ( \37724 , \34711 );
or \U$37348 ( \37725 , \37723 , \37724 );
nand \U$37349 ( \37726 , \32716 , \9552 );
nand \U$37350 ( \37727 , \37725 , \37726 );
and \U$37351 ( \37728 , \37722 , \37727 );
and \U$37352 ( \37729 , \37716 , \37721 );
or \U$37353 ( \37730 , \37728 , \37729 );
xor \U$37354 ( \37731 , \34690 , \34695 );
and \U$37355 ( \37732 , \37731 , \34701 );
and \U$37356 ( \37733 , \34690 , \34695 );
or \U$37357 ( \37734 , \37732 , \37733 );
not \U$37358 ( \37735 , \9488 );
not \U$37359 ( \37736 , \34642 );
or \U$37360 ( \37737 , \37735 , \37736 );
nand \U$37361 ( \37738 , \32826 , \8788 );
nand \U$37362 ( \37739 , \37737 , \37738 );
xor \U$37363 ( \37740 , \37734 , \37739 );
not \U$37364 ( \37741 , \9690 );
not \U$37365 ( \37742 , \34619 );
or \U$37366 ( \37743 , \37741 , \37742 );
nand \U$37367 ( \37744 , \32762 , \9705 );
nand \U$37368 ( \37745 , \37743 , \37744 );
and \U$37369 ( \37746 , \37740 , \37745 );
and \U$37370 ( \37747 , \37734 , \37739 );
or \U$37371 ( \37748 , \37746 , \37747 );
xor \U$37372 ( \37749 , \37730 , \37748 );
and \U$37373 ( \37750 , \35697 , \9110 );
and \U$37374 ( \37751 , \32736 , \9129 );
nor \U$37375 ( \37752 , \37750 , \37751 );
and \U$37376 ( \37753 , \35708 , \9934 );
and \U$37377 ( \37754 , \32747 , \9398 );
nor \U$37378 ( \37755 , \37753 , \37754 );
xor \U$37379 ( \37756 , \37752 , \37755 );
not \U$37380 ( \37757 , \34721 );
not \U$37381 ( \37758 , \9640 );
and \U$37382 ( \37759 , \37757 , \37758 );
and \U$37383 ( \37760 , \32706 , \12304 );
nor \U$37384 ( \37761 , \37759 , \37760 );
and \U$37385 ( \37762 , \37756 , \37761 );
and \U$37386 ( \37763 , \37752 , \37755 );
or \U$37387 ( \37764 , \37762 , \37763 );
not \U$37388 ( \37765 , \37764 );
xnor \U$37389 ( \37766 , \37749 , \37765 );
xor \U$37390 ( \37767 , \37711 , \37766 );
xor \U$37391 ( \37768 , \35761 , \35770 );
and \U$37392 ( \37769 , \37768 , \35780 );
and \U$37393 ( \37770 , \35761 , \35770 );
or \U$37394 ( \37771 , \37769 , \37770 );
xor \U$37395 ( \37772 , \37752 , \37755 );
xor \U$37396 ( \37773 , \37772 , \37761 );
nand \U$37397 ( \37774 , \37771 , \37773 );
xor \U$37398 ( \37775 , \37734 , \37739 );
xor \U$37399 ( \37776 , \37775 , \37745 );
and \U$37400 ( \37777 , \37774 , \37776 );
nor \U$37401 ( \37778 , \37771 , \37773 );
nor \U$37402 ( \37779 , \37777 , \37778 );
xor \U$37403 ( \37780 , \37767 , \37779 );
not \U$37404 ( \37781 , \37780 );
not \U$37405 ( \37782 , \37781 );
not \U$37406 ( \37783 , \35782 );
not \U$37407 ( \37784 , \35713 );
or \U$37408 ( \37785 , \37783 , \37784 );
not \U$37409 ( \37786 , \35713 );
not \U$37410 ( \37787 , \37786 );
not \U$37411 ( \37788 , \35781 );
or \U$37412 ( \37789 , \37787 , \37788 );
nand \U$37413 ( \37790 , \37789 , \35755 );
nand \U$37414 ( \37791 , \37785 , \37790 );
not \U$37415 ( \37792 , \37791 );
xor \U$37416 ( \37793 , \37689 , \37694 );
xor \U$37417 ( \37794 , \37793 , \37700 );
xor \U$37418 ( \37795 , \37716 , \37721 );
xor \U$37419 ( \37796 , \37795 , \37727 );
xor \U$37420 ( \37797 , \37794 , \37796 );
xor \U$37421 ( \37798 , \35690 , \35701 );
and \U$37422 ( \37799 , \37798 , \35712 );
and \U$37423 ( \37800 , \35690 , \35701 );
or \U$37424 ( \37801 , \37799 , \37800 );
xnor \U$37425 ( \37802 , \37797 , \37801 );
nand \U$37426 ( \37803 , \37792 , \37802 );
xor \U$37427 ( \37804 , \34623 , \34634 );
and \U$37428 ( \37805 , \37804 , \34646 );
and \U$37429 ( \37806 , \34623 , \34634 );
or \U$37430 ( \37807 , \37805 , \37806 );
xor \U$37431 ( \37808 , \34702 , \34713 );
and \U$37432 ( \37809 , \37808 , \34724 );
and \U$37433 ( \37810 , \34702 , \34713 );
or \U$37434 ( \37811 , \37809 , \37810 );
xor \U$37435 ( \37812 , \37807 , \37811 );
not \U$37436 ( \37813 , \13025 );
not \U$37437 ( \37814 , RIc225c60_55);
not \U$37438 ( \37815 , \19926 );
or \U$37439 ( \37816 , \37814 , \37815 );
nand \U$37440 ( \37817 , \4050 , \11041 );
nand \U$37441 ( \37818 , \37816 , \37817 );
not \U$37442 ( \37819 , \37818 );
or \U$37443 ( \37820 , \37813 , \37819 );
not \U$37444 ( \37821 , \35758 );
nand \U$37445 ( \37822 , \37821 , \11118 );
nand \U$37446 ( \37823 , \37820 , \37822 );
not \U$37447 ( \37824 , \9444 );
not \U$37448 ( \37825 , RIc225e40_51);
not \U$37449 ( \37826 , \20656 );
or \U$37450 ( \37827 , \37825 , \37826 );
not \U$37451 ( \37828 , \5664 );
nand \U$37452 ( \37829 , \37828 , \11795 );
nand \U$37453 ( \37830 , \37827 , \37829 );
not \U$37454 ( \37831 , \37830 );
or \U$37455 ( \37832 , \37824 , \37831 );
nand \U$37456 ( \37833 , \34630 , \9459 );
nand \U$37457 ( \37834 , \37832 , \37833 );
xor \U$37458 ( \37835 , \37823 , \37834 );
not \U$37459 ( \37836 , \11965 );
not \U$37460 ( \37837 , \35767 );
or \U$37461 ( \37838 , \37836 , \37837 );
not \U$37462 ( \37839 , RIc225b70_57);
not \U$37463 ( \37840 , \15755 );
or \U$37464 ( \37841 , \37839 , \37840 );
nand \U$37465 ( \37842 , \11320 , \11033 );
nand \U$37466 ( \37843 , \37841 , \37842 );
nand \U$37467 ( \37844 , \37843 , \15267 );
nand \U$37468 ( \37845 , \37838 , \37844 );
xor \U$37469 ( \37846 , \37835 , \37845 );
xor \U$37470 ( \37847 , \37812 , \37846 );
and \U$37471 ( \37848 , \37803 , \37847 );
not \U$37472 ( \37849 , \37791 );
nor \U$37473 ( \37850 , \37849 , \37802 );
nor \U$37474 ( \37851 , \37848 , \37850 );
not \U$37475 ( \37852 , \37851 );
or \U$37476 ( \37853 , \37782 , \37852 );
not \U$37477 ( \37854 , \37851 );
nand \U$37478 ( \37855 , \37854 , \37780 );
nand \U$37479 ( \37856 , \37853 , \37855 );
xor \U$37480 ( \37857 , \37807 , \37811 );
and \U$37481 ( \37858 , \37857 , \37846 );
and \U$37482 ( \37859 , \37807 , \37811 );
or \U$37483 ( \37860 , \37858 , \37859 );
xor \U$37484 ( \37861 , \32764 , \32740 );
xor \U$37485 ( \37862 , \37861 , \32751 );
xor \U$37486 ( \37863 , \32781 , \32790 );
xor \U$37487 ( \37864 , \37863 , \32802 );
not \U$37488 ( \37865 , \15719 );
not \U$37489 ( \37866 , \35740 );
or \U$37490 ( \37867 , \37865 , \37866 );
not \U$37491 ( \37868 , RIc225990_61);
not \U$37492 ( \37869 , \3010 );
or \U$37493 ( \37870 , \37868 , \37869 );
nand \U$37494 ( \37871 , \17966 , \12806 );
nand \U$37495 ( \37872 , \37870 , \37871 );
nand \U$37496 ( \37873 , \37872 , \15729 );
nand \U$37497 ( \37874 , \37867 , \37873 );
xor \U$37498 ( \37875 , \37864 , \37874 );
not \U$37499 ( \37876 , \20159 );
not \U$37500 ( \37877 , \35777 );
or \U$37501 ( \37878 , \37876 , \37877 );
not \U$37502 ( \37879 , RIc2258a0_63);
not \U$37503 ( \37880 , \2501 );
or \U$37504 ( \37881 , \37879 , \37880 );
nand \U$37505 ( \37882 , \17122 , \16880 );
nand \U$37506 ( \37883 , \37881 , \37882 );
nand \U$37507 ( \37884 , \37883 , RIc225828_64);
nand \U$37508 ( \37885 , \37878 , \37884 );
and \U$37509 ( \37886 , \37875 , \37885 );
and \U$37510 ( \37887 , \37864 , \37874 );
or \U$37511 ( \37888 , \37886 , \37887 );
xor \U$37512 ( \37889 , \37862 , \37888 );
xor \U$37513 ( \37890 , \34589 , \34599 );
and \U$37514 ( \37891 , \37890 , \34610 );
and \U$37515 ( \37892 , \34589 , \34599 );
or \U$37516 ( \37893 , \37891 , \37892 );
xor \U$37517 ( \37894 , \35718 , \35722 );
and \U$37518 ( \37895 , \37894 , \35733 );
and \U$37519 ( \37896 , \35718 , \35722 );
or \U$37520 ( \37897 , \37895 , \37896 );
xor \U$37521 ( \37898 , \37893 , \37897 );
not \U$37522 ( \37899 , \15164 );
not \U$37523 ( \37900 , \35750 );
or \U$37524 ( \37901 , \37899 , \37900 );
and \U$37525 ( \37902 , RIc225a80_59, \2635 );
not \U$37526 ( \37903 , RIc225a80_59);
and \U$37527 ( \37904 , \37903 , \5386 );
or \U$37528 ( \37905 , \37902 , \37904 );
nand \U$37529 ( \37906 , \37905 , \12670 );
nand \U$37530 ( \37907 , \37901 , \37906 );
and \U$37531 ( \37908 , \37898 , \37907 );
and \U$37532 ( \37909 , \37893 , \37897 );
or \U$37533 ( \37910 , \37908 , \37909 );
xor \U$37534 ( \37911 , \37889 , \37910 );
xor \U$37535 ( \37912 , \37860 , \37911 );
xor \U$37536 ( \37913 , \32805 , \32817 );
xor \U$37537 ( \37914 , \37913 , \32828 );
xor \U$37538 ( \37915 , \32701 , \32710 );
xor \U$37539 ( \37916 , \37915 , \32721 );
xor \U$37540 ( \37917 , \37914 , \37916 );
xor \U$37541 ( \37918 , \37823 , \37834 );
and \U$37542 ( \37919 , \37918 , \37845 );
and \U$37543 ( \37920 , \37823 , \37834 );
or \U$37544 ( \37921 , \37919 , \37920 );
xor \U$37545 ( \37922 , \37917 , \37921 );
xor \U$37546 ( \37923 , \37912 , \37922 );
xnor \U$37547 ( \37924 , \37856 , \37923 );
xor \U$37548 ( \37925 , \37776 , \37773 );
xor \U$37549 ( \37926 , \37925 , \37771 );
not \U$37550 ( \37927 , \37926 );
not \U$37551 ( \37928 , \34611 );
not \U$37552 ( \37929 , \34574 );
or \U$37553 ( \37930 , \37928 , \37929 );
or \U$37554 ( \37931 , \34574 , \34611 );
nand \U$37555 ( \37932 , \37931 , \34567 );
nand \U$37556 ( \37933 , \37930 , \37932 );
xor \U$37557 ( \37934 , \35734 , \35744 );
and \U$37558 ( \37935 , \37934 , \35754 );
and \U$37559 ( \37936 , \35734 , \35744 );
or \U$37560 ( \37937 , \37935 , \37936 );
xor \U$37561 ( \37938 , \37933 , \37937 );
xor \U$37562 ( \37939 , \37864 , \37874 );
xor \U$37563 ( \37940 , \37939 , \37885 );
xor \U$37564 ( \37941 , \37938 , \37940 );
not \U$37565 ( \37942 , \37941 );
or \U$37566 ( \37943 , \37927 , \37942 );
not \U$37567 ( \37944 , \34557 );
nand \U$37568 ( \37945 , \34480 , \37944 );
and \U$37569 ( \37946 , \37945 , \34553 );
nor \U$37570 ( \37947 , \37944 , \34480 );
nor \U$37571 ( \37948 , \37946 , \37947 );
not \U$37572 ( \37949 , \37948 );
or \U$37573 ( \37950 , \37941 , \37926 );
nand \U$37574 ( \37951 , \37949 , \37950 );
nand \U$37575 ( \37952 , \37943 , \37951 );
xor \U$37576 ( \37953 , \37933 , \37937 );
and \U$37577 ( \37954 , \37953 , \37940 );
and \U$37578 ( \37955 , \37933 , \37937 );
or \U$37579 ( \37956 , \37954 , \37955 );
not \U$37580 ( \37957 , \9459 );
not \U$37581 ( \37958 , \37830 );
or \U$37582 ( \37959 , \37957 , \37958 );
nand \U$37583 ( \37960 , \32503 , \9444 );
nand \U$37584 ( \37961 , \37959 , \37960 );
not \U$37585 ( \37962 , \11965 );
not \U$37586 ( \37963 , \37843 );
or \U$37587 ( \37964 , \37962 , \37963 );
nand \U$37588 ( \37965 , \32522 , \11974 );
nand \U$37589 ( \37966 , \37964 , \37965 );
xor \U$37590 ( \37967 , \37961 , \37966 );
not \U$37591 ( \37968 , \15729 );
not \U$37592 ( \37969 , \32540 );
or \U$37593 ( \37970 , \37968 , \37969 );
nand \U$37594 ( \37971 , \37872 , \15719 );
nand \U$37595 ( \37972 , \37970 , \37971 );
xor \U$37596 ( \37973 , \37967 , \37972 );
not \U$37597 ( \37974 , RIc225828_64);
not \U$37598 ( \37975 , \32627 );
or \U$37599 ( \37976 , \37974 , \37975 );
nand \U$37600 ( \37977 , \37883 , \16891 );
nand \U$37601 ( \37978 , \37976 , \37977 );
not \U$37602 ( \37979 , \13025 );
not \U$37603 ( \37980 , \32551 );
or \U$37604 ( \37981 , \37979 , \37980 );
nand \U$37605 ( \37982 , \37818 , \11118 );
nand \U$37606 ( \37983 , \37981 , \37982 );
xor \U$37607 ( \37984 , \37978 , \37983 );
not \U$37608 ( \37985 , \15164 );
not \U$37609 ( \37986 , \37905 );
or \U$37610 ( \37987 , \37985 , \37986 );
nand \U$37611 ( \37988 , \32639 , \12670 );
nand \U$37612 ( \37989 , \37987 , \37988 );
xor \U$37613 ( \37990 , \37984 , \37989 );
xor \U$37614 ( \37991 , \37973 , \37990 );
or \U$37615 ( \37992 , \37794 , \37796 );
nand \U$37616 ( \37993 , \37992 , \37801 );
nand \U$37617 ( \37994 , \37796 , \37794 );
nand \U$37618 ( \37995 , \37993 , \37994 );
xor \U$37619 ( \37996 , \37991 , \37995 );
xor \U$37620 ( \37997 , \37956 , \37996 );
not \U$37621 ( \37998 , \34655 );
not \U$37622 ( \37999 , \34647 );
or \U$37623 ( \38000 , \37998 , \37999 );
or \U$37624 ( \38001 , \34655 , \34647 );
nand \U$37625 ( \38002 , \38001 , \34683 );
nand \U$37626 ( \38003 , \38000 , \38002 );
xor \U$37627 ( \38004 , \37893 , \37897 );
xor \U$37628 ( \38005 , \38004 , \37907 );
or \U$37629 ( \38006 , \38003 , \38005 );
not \U$37630 ( \38007 , \38006 );
xor \U$37631 ( \38008 , \34725 , \34731 );
and \U$37632 ( \38009 , \38008 , \34784 );
and \U$37633 ( \38010 , \34725 , \34731 );
or \U$37634 ( \38011 , \38009 , \38010 );
not \U$37635 ( \38012 , \38011 );
or \U$37636 ( \38013 , \38007 , \38012 );
nand \U$37637 ( \38014 , \38003 , \38005 );
nand \U$37638 ( \38015 , \38013 , \38014 );
xor \U$37639 ( \38016 , \37997 , \38015 );
xor \U$37640 ( \38017 , \37952 , \38016 );
xor \U$37641 ( \38018 , \38005 , \38003 );
xnor \U$37642 ( \38019 , \38018 , \38011 );
not \U$37643 ( \38020 , \38019 );
not \U$37644 ( \38021 , \38020 );
xor \U$37645 ( \38022 , \34612 , \34688 );
and \U$37646 ( \38023 , \38022 , \34785 );
and \U$37647 ( \38024 , \34612 , \34688 );
or \U$37648 ( \38025 , \38023 , \38024 );
not \U$37649 ( \38026 , \38025 );
or \U$37650 ( \38027 , \38021 , \38026 );
xor \U$37651 ( \38028 , \37802 , \37847 );
xnor \U$37652 ( \38029 , \38028 , \37791 );
not \U$37653 ( \38030 , \38025 );
nand \U$37654 ( \38031 , \38030 , \38019 );
nand \U$37655 ( \38032 , \38029 , \38031 );
nand \U$37656 ( \38033 , \38027 , \38032 );
xnor \U$37657 ( \38034 , \38017 , \38033 );
xor \U$37658 ( \38035 , \37924 , \38034 );
not \U$37659 ( \38036 , \34562 );
not \U$37660 ( \38037 , \34473 );
or \U$37661 ( \38038 , \38036 , \38037 );
or \U$37662 ( \38039 , \34473 , \34562 );
nand \U$37663 ( \38040 , \38039 , \34786 );
nand \U$37664 ( \38041 , \38038 , \38040 );
not \U$37665 ( \38042 , \35682 );
not \U$37666 ( \38043 , \35784 );
or \U$37667 ( \38044 , \38042 , \38043 );
not \U$37668 ( \38045 , \35681 );
not \U$37669 ( \38046 , \35783 );
or \U$37670 ( \38047 , \38045 , \38046 );
nand \U$37671 ( \38048 , \38047 , \35675 );
nand \U$37672 ( \38049 , \38044 , \38048 );
or \U$37673 ( \38050 , \38041 , \38049 );
xor \U$37674 ( \38051 , \37941 , \37926 );
xor \U$37675 ( \38052 , \38051 , \37948 );
not \U$37676 ( \38053 , \38052 );
nand \U$37677 ( \38054 , \38050 , \38053 );
nand \U$37678 ( \38055 , \38041 , \38049 );
and \U$37679 ( \38056 , \38054 , \38055 );
xor \U$37680 ( \38057 , \38035 , \38056 );
xor \U$37681 ( \38058 , \35643 , \35785 );
and \U$37682 ( \38059 , \38058 , \35815 );
and \U$37683 ( \38060 , \35643 , \35785 );
or \U$37684 ( \38061 , \38059 , \38060 );
xor \U$37685 ( \38062 , \38025 , \38020 );
xor \U$37686 ( \38063 , \38062 , \38029 );
or \U$37687 ( \38064 , \38061 , \38063 );
xor \U$37688 ( \38065 , \38049 , \38052 );
xnor \U$37689 ( \38066 , \38065 , \38041 );
buf \U$37690 ( \38067 , \38066 );
and \U$37691 ( \38068 , \38064 , \38067 );
and \U$37692 ( \38069 , \38061 , \38063 );
nor \U$37693 ( \38070 , \38068 , \38069 );
nand \U$37694 ( \38071 , \38057 , \38070 );
xor \U$37695 ( \38072 , \32730 , \32766 );
xor \U$37696 ( \38073 , \38072 , \32831 );
xor \U$37697 ( \38074 , \32696 , \32698 );
xor \U$37698 ( \38075 , \38074 , \32724 );
xor \U$37699 ( \38076 , \38073 , \38075 );
xor \U$37700 ( \38077 , \37914 , \37916 );
and \U$37701 ( \38078 , \38077 , \37921 );
and \U$37702 ( \38079 , \37914 , \37916 );
or \U$37703 ( \38080 , \38078 , \38079 );
xor \U$37704 ( \38081 , \38076 , \38080 );
xor \U$37705 ( \38082 , \37860 , \37911 );
and \U$37706 ( \38083 , \38082 , \37922 );
and \U$37707 ( \38084 , \37860 , \37911 );
or \U$37708 ( \38085 , \38083 , \38084 );
xor \U$37709 ( \38086 , \38081 , \38085 );
or \U$37710 ( \38087 , \37862 , \37888 );
nand \U$37711 ( \38088 , \38087 , \37910 );
nand \U$37712 ( \38089 , \37888 , \37862 );
nand \U$37713 ( \38090 , \38088 , \38089 );
xor \U$37714 ( \38091 , \37961 , \37966 );
and \U$37715 ( \38092 , \38091 , \37972 );
and \U$37716 ( \38093 , \37961 , \37966 );
or \U$37717 ( \38094 , \38092 , \38093 );
xor \U$37718 ( \38095 , \32457 , \32467 );
xor \U$37719 ( \38096 , \38095 , \32478 );
xor \U$37720 ( \38097 , \38094 , \38096 );
xor \U$37721 ( \38098 , \32505 , \32515 );
xor \U$37722 ( \38099 , \38098 , \32526 );
xnor \U$37723 ( \38100 , \38097 , \38099 );
and \U$37724 ( \38101 , \38090 , \38100 );
not \U$37725 ( \38102 , \38090 );
not \U$37726 ( \38103 , \38100 );
and \U$37727 ( \38104 , \38102 , \38103 );
or \U$37728 ( \38105 , \38101 , \38104 );
xor \U$37729 ( \38106 , \32400 , \32410 );
xor \U$37730 ( \38107 , \38106 , \32422 );
xor \U$37731 ( \38108 , \37978 , \37983 );
and \U$37732 ( \38109 , \38108 , \37989 );
and \U$37733 ( \38110 , \37978 , \37983 );
or \U$37734 ( \38111 , \38109 , \38110 );
xor \U$37735 ( \38112 , \38107 , \38111 );
xor \U$37736 ( \38113 , \32621 , \32631 );
xor \U$37737 ( \38114 , \38113 , \32641 );
xor \U$37738 ( \38115 , \38112 , \38114 );
not \U$37739 ( \38116 , \38115 );
and \U$37740 ( \38117 , \38105 , \38116 );
not \U$37741 ( \38118 , \38105 );
and \U$37742 ( \38119 , \38118 , \38115 );
nor \U$37743 ( \38120 , \38117 , \38119 );
xnor \U$37744 ( \38121 , \38086 , \38120 );
not \U$37745 ( \38122 , \37952 );
not \U$37746 ( \38123 , \38016 );
or \U$37747 ( \38124 , \38122 , \38123 );
or \U$37748 ( \38125 , \37952 , \38016 );
nand \U$37749 ( \38126 , \38125 , \38033 );
nand \U$37750 ( \38127 , \38124 , \38126 );
xor \U$37751 ( \38128 , \38121 , \38127 );
xor \U$37752 ( \38129 , \37956 , \37996 );
and \U$37753 ( \38130 , \38129 , \38015 );
and \U$37754 ( \38131 , \37956 , \37996 );
or \U$37755 ( \38132 , \38130 , \38131 );
or \U$37756 ( \38133 , \37990 , \37973 );
and \U$37757 ( \38134 , \38133 , \37995 );
and \U$37758 ( \38135 , \37973 , \37990 );
nor \U$37759 ( \38136 , \38134 , \38135 );
not \U$37760 ( \38137 , \37687 );
nand \U$37761 ( \38138 , \38137 , \37710 );
and \U$37762 ( \38139 , \38138 , \37703 );
not \U$37763 ( \38140 , \37687 );
nor \U$37764 ( \38141 , \38140 , \37710 );
nor \U$37765 ( \38142 , \38139 , \38141 );
xor \U$37766 ( \38143 , \32532 , \32542 );
xor \U$37767 ( \38144 , \38143 , \32553 );
xor \U$37768 ( \38145 , \38142 , \38144 );
not \U$37769 ( \38146 , \37730 );
not \U$37770 ( \38147 , \38146 );
not \U$37771 ( \38148 , \37764 );
or \U$37772 ( \38149 , \38147 , \38148 );
nand \U$37773 ( \38150 , \38149 , \37748 );
nand \U$37774 ( \38151 , \37765 , \37730 );
nand \U$37775 ( \38152 , \38150 , \38151 );
xor \U$37776 ( \38153 , \38145 , \38152 );
xor \U$37777 ( \38154 , \38136 , \38153 );
xor \U$37778 ( \38155 , \37711 , \37766 );
and \U$37779 ( \38156 , \38155 , \37779 );
and \U$37780 ( \38157 , \37711 , \37766 );
or \U$37781 ( \38158 , \38156 , \38157 );
xor \U$37782 ( \38159 , \38154 , \38158 );
xor \U$37783 ( \38160 , \38132 , \38159 );
not \U$37784 ( \38161 , \37854 );
not \U$37785 ( \38162 , \37781 );
or \U$37786 ( \38163 , \38161 , \38162 );
not \U$37787 ( \38164 , \37780 );
not \U$37788 ( \38165 , \37851 );
or \U$37789 ( \38166 , \38164 , \38165 );
nand \U$37790 ( \38167 , \38166 , \37923 );
nand \U$37791 ( \38168 , \38163 , \38167 );
xnor \U$37792 ( \38169 , \38160 , \38168 );
xnor \U$37793 ( \38170 , \38128 , \38169 );
xor \U$37794 ( \38171 , \37924 , \38034 );
and \U$37795 ( \38172 , \38171 , \38056 );
and \U$37796 ( \38173 , \37924 , \38034 );
or \U$37797 ( \38174 , \38172 , \38173 );
nand \U$37798 ( \38175 , \38170 , \38174 );
xor \U$37799 ( \38176 , \38063 , \38066 );
xor \U$37800 ( \38177 , \38176 , \38061 );
not \U$37801 ( \38178 , \38177 );
buf \U$37802 ( \38179 , \34787 );
or \U$37803 ( \38180 , \38179 , \35816 );
nand \U$37804 ( \38181 , \38180 , \35634 );
nand \U$37805 ( \38182 , \38179 , \35816 );
nand \U$37806 ( \38183 , \38181 , \38182 );
not \U$37807 ( \38184 , \38183 );
nand \U$37808 ( \38185 , \38178 , \38184 );
and \U$37809 ( \38186 , \32562 , \32644 );
not \U$37810 ( \38187 , \32562 );
not \U$37811 ( \38188 , \32644 );
and \U$37812 ( \38189 , \38187 , \38188 );
nor \U$37813 ( \38190 , \38186 , \38189 );
not \U$37814 ( \38191 , \32568 );
and \U$37815 ( \38192 , \38190 , \38191 );
not \U$37816 ( \38193 , \38190 );
and \U$37817 ( \38194 , \38193 , \32568 );
nor \U$37818 ( \38195 , \38192 , \38194 );
xor \U$37819 ( \38196 , \32481 , \32489 );
xor \U$37820 ( \38197 , \38196 , \32485 );
xor \U$37821 ( \38198 , \38107 , \38111 );
and \U$37822 ( \38199 , \38198 , \38114 );
and \U$37823 ( \38200 , \38107 , \38111 );
or \U$37824 ( \38201 , \38199 , \38200 );
or \U$37825 ( \38202 , \38197 , \38201 );
nand \U$37826 ( \38203 , \38201 , \38197 );
nand \U$37827 ( \38204 , \38202 , \38203 );
not \U$37828 ( \38205 , \38204 );
xor \U$37829 ( \38206 , \38195 , \38205 );
buf \U$37830 ( \38207 , \38206 );
not \U$37831 ( \38208 , \38090 );
not \U$37832 ( \38209 , \38103 );
or \U$37833 ( \38210 , \38208 , \38209 );
or \U$37834 ( \38211 , \38090 , \38103 );
nand \U$37835 ( \38212 , \38211 , \38115 );
nand \U$37836 ( \38213 , \38210 , \38212 );
not \U$37837 ( \38214 , \38096 );
not \U$37838 ( \38215 , \38094 );
or \U$37839 ( \38216 , \38214 , \38215 );
or \U$37840 ( \38217 , \38096 , \38094 );
nand \U$37841 ( \38218 , \38217 , \38099 );
nand \U$37842 ( \38219 , \38216 , \38218 );
xor \U$37843 ( \38220 , \32338 , \32373 );
xor \U$37844 ( \38221 , \38220 , \32425 );
not \U$37845 ( \38222 , \38221 );
and \U$37846 ( \38223 , \38219 , \38222 );
not \U$37847 ( \38224 , \38219 );
and \U$37848 ( \38225 , \38224 , \38221 );
or \U$37849 ( \38226 , \38223 , \38225 );
xor \U$37850 ( \38227 , \32495 , \32529 );
xor \U$37851 ( \38228 , \38227 , \32556 );
xor \U$37852 ( \38229 , \38226 , \38228 );
not \U$37853 ( \38230 , \38229 );
and \U$37854 ( \38231 , \38213 , \38230 );
not \U$37855 ( \38232 , \38213 );
and \U$37856 ( \38233 , \38232 , \38229 );
nor \U$37857 ( \38234 , \38231 , \38233 );
xnor \U$37858 ( \38235 , \38207 , \38234 );
not \U$37859 ( \38236 , \38132 );
not \U$37860 ( \38237 , \38236 );
not \U$37861 ( \38238 , \38159 );
or \U$37862 ( \38239 , \38237 , \38238 );
nand \U$37863 ( \38240 , \38239 , \38168 );
not \U$37864 ( \38241 , \38240 );
nor \U$37865 ( \38242 , \38159 , \38236 );
nor \U$37866 ( \38243 , \38241 , \38242 );
xor \U$37867 ( \38244 , \38235 , \38243 );
xor \U$37868 ( \38245 , \38136 , \38153 );
and \U$37869 ( \38246 , \38245 , \38158 );
and \U$37870 ( \38247 , \38136 , \38153 );
or \U$37871 ( \38248 , \38246 , \38247 );
not \U$37872 ( \38249 , \38152 );
not \U$37873 ( \38250 , \38144 );
nand \U$37874 ( \38251 , \38250 , \38142 );
not \U$37875 ( \38252 , \38251 );
or \U$37876 ( \38253 , \38249 , \38252 );
not \U$37877 ( \38254 , \38142 );
nand \U$37878 ( \38255 , \38254 , \38144 );
nand \U$37879 ( \38256 , \38253 , \38255 );
xor \U$37880 ( \38257 , \32660 , \32727 );
xor \U$37881 ( \38258 , \38257 , \32834 );
xor \U$37882 ( \38259 , \38256 , \38258 );
xor \U$37883 ( \38260 , \38073 , \38075 );
and \U$37884 ( \38261 , \38260 , \38080 );
and \U$37885 ( \38262 , \38073 , \38075 );
or \U$37886 ( \38263 , \38261 , \38262 );
xnor \U$37887 ( \38264 , \38259 , \38263 );
xor \U$37888 ( \38265 , \38248 , \38264 );
not \U$37889 ( \38266 , \38081 );
nand \U$37890 ( \38267 , \38120 , \38266 );
and \U$37891 ( \38268 , \38267 , \38085 );
nor \U$37892 ( \38269 , \38120 , \38266 );
nor \U$37893 ( \38270 , \38268 , \38269 );
xor \U$37894 ( \38271 , \38265 , \38270 );
xor \U$37895 ( \38272 , \38244 , \38271 );
or \U$37896 ( \38273 , \38127 , \38121 );
and \U$37897 ( \38274 , \38169 , \38273 );
and \U$37898 ( \38275 , \38127 , \38121 );
nor \U$37899 ( \38276 , \38274 , \38275 );
nand \U$37900 ( \38277 , \38272 , \38276 );
and \U$37901 ( \38278 , \38071 , \38175 , \38185 , \38277 );
not \U$37902 ( \38279 , \38278 );
nor \U$37903 ( \38280 , \37685 , \38279 );
nand \U$37904 ( \38281 , \38177 , \38183 );
not \U$37905 ( \38282 , \38281 );
nand \U$37906 ( \38283 , \38282 , \38071 );
or \U$37907 ( \38284 , \38057 , \38070 );
nand \U$37908 ( \38285 , \38283 , \38284 );
nand \U$37909 ( \38286 , \38285 , \38175 );
not \U$37910 ( \38287 , \38170 );
not \U$37911 ( \38288 , \38174 );
nand \U$37912 ( \38289 , \38287 , \38288 );
not \U$37913 ( \38290 , \38272 );
not \U$37914 ( \38291 , \38276 );
nand \U$37915 ( \38292 , \38290 , \38291 );
and \U$37916 ( \38293 , \38289 , \38292 );
and \U$37917 ( \38294 , \38286 , \38293 );
not \U$37918 ( \38295 , \38277 );
nor \U$37919 ( \38296 , \38294 , \38295 );
or \U$37920 ( \38297 , \38280 , \38296 );
xor \U$37921 ( \38298 , \32214 , \32232 );
xnor \U$37922 ( \38299 , \38298 , \32212 );
xor \U$37923 ( \38300 , \32012 , \32094 );
xor \U$37924 ( \38301 , \38300 , \32097 );
xor \U$37925 ( \38302 , \32430 , \32432 );
xor \U$37926 ( \38303 , \38302 , \32435 );
xor \U$37927 ( \38304 , \38301 , \38303 );
not \U$37928 ( \38305 , \38222 );
not \U$37929 ( \38306 , \38219 );
or \U$37930 ( \38307 , \38305 , \38306 );
not \U$37931 ( \38308 , \38219 );
nand \U$37932 ( \38309 , \38308 , \38221 );
nand \U$37933 ( \38310 , \38309 , \38228 );
nand \U$37934 ( \38311 , \38307 , \38310 );
and \U$37935 ( \38312 , \38304 , \38311 );
and \U$37936 ( \38313 , \38301 , \38303 );
or \U$37937 ( \38314 , \38312 , \38313 );
not \U$37938 ( \38315 , \38314 );
xor \U$37939 ( \38316 , \32438 , \32440 );
xor \U$37940 ( \38317 , \38316 , \32443 );
not \U$37941 ( \38318 , \38317 );
or \U$37942 ( \38319 , \38315 , \38318 );
or \U$37943 ( \38320 , \38314 , \38317 );
xor \U$37944 ( \38321 , \32652 , \32657 );
xor \U$37945 ( \38322 , \38321 , \32837 );
xor \U$37946 ( \38323 , \32493 , \32559 );
xor \U$37947 ( \38324 , \38323 , \32647 );
or \U$37948 ( \38325 , \38322 , \38324 );
nand \U$37949 ( \38326 , \38195 , \38197 );
and \U$37950 ( \38327 , \38326 , \38201 );
nor \U$37951 ( \38328 , \38195 , \38197 );
nor \U$37952 ( \38329 , \38327 , \38328 );
not \U$37953 ( \38330 , \38329 );
nand \U$37954 ( \38331 , \38325 , \38330 );
nand \U$37955 ( \38332 , \38322 , \38324 );
nand \U$37956 ( \38333 , \38331 , \38332 );
nand \U$37957 ( \38334 , \38320 , \38333 );
nand \U$37958 ( \38335 , \38319 , \38334 );
not \U$37959 ( \38336 , \38335 );
xor \U$37960 ( \38337 , \38299 , \38336 );
xor \U$37961 ( \38338 , \32446 , \32336 );
xnor \U$37962 ( \38339 , \38338 , \32846 );
xor \U$37963 ( \38340 , \38337 , \38339 );
xor \U$37964 ( \38341 , \32840 , \32650 );
not \U$37965 ( \38342 , \32843 );
and \U$37966 ( \38343 , \38341 , \38342 );
not \U$37967 ( \38344 , \38341 );
and \U$37968 ( \38345 , \38344 , \32843 );
nor \U$37969 ( \38346 , \38343 , \38345 );
not \U$37970 ( \38347 , \38256 );
not \U$37971 ( \38348 , \38258 );
or \U$37972 ( \38349 , \38347 , \38348 );
or \U$37973 ( \38350 , \38258 , \38256 );
nand \U$37974 ( \38351 , \38350 , \38263 );
nand \U$37975 ( \38352 , \38349 , \38351 );
xor \U$37976 ( \38353 , \38301 , \38303 );
xor \U$37977 ( \38354 , \38353 , \38311 );
or \U$37978 ( \38355 , \38352 , \38354 );
not \U$37979 ( \38356 , \38213 );
nand \U$37980 ( \38357 , \38356 , \38229 );
not \U$37981 ( \38358 , \38357 );
not \U$37982 ( \38359 , \38206 );
or \U$37983 ( \38360 , \38358 , \38359 );
nand \U$37984 ( \38361 , \38213 , \38230 );
nand \U$37985 ( \38362 , \38360 , \38361 );
nand \U$37986 ( \38363 , \38355 , \38362 );
nand \U$37987 ( \38364 , \38354 , \38352 );
and \U$37988 ( \38365 , \38363 , \38364 );
xor \U$37989 ( \38366 , \38346 , \38365 );
xor \U$37990 ( \38367 , \38314 , \38317 );
xnor \U$37991 ( \38368 , \38367 , \38333 );
and \U$37992 ( \38369 , \38366 , \38368 );
and \U$37993 ( \38370 , \38346 , \38365 );
or \U$37994 ( \38371 , \38369 , \38370 );
nand \U$37995 ( \38372 , \38340 , \38371 );
xor \U$37996 ( \38373 , \38346 , \38365 );
xor \U$37997 ( \38374 , \38373 , \38368 );
not \U$37998 ( \38375 , \38329 );
not \U$37999 ( \38376 , \38322 );
or \U$38000 ( \38377 , \38375 , \38376 );
or \U$38001 ( \38378 , \38322 , \38329 );
nand \U$38002 ( \38379 , \38377 , \38378 );
not \U$38003 ( \38380 , \38324 );
and \U$38004 ( \38381 , \38379 , \38380 );
not \U$38005 ( \38382 , \38379 );
and \U$38006 ( \38383 , \38382 , \38324 );
nor \U$38007 ( \38384 , \38381 , \38383 );
xor \U$38008 ( \38385 , \38248 , \38264 );
and \U$38009 ( \38386 , \38385 , \38270 );
and \U$38010 ( \38387 , \38248 , \38264 );
or \U$38011 ( \38388 , \38386 , \38387 );
xor \U$38012 ( \38389 , \38384 , \38388 );
xor \U$38013 ( \38390 , \38352 , \38354 );
xnor \U$38014 ( \38391 , \38390 , \38362 );
and \U$38015 ( \38392 , \38389 , \38391 );
and \U$38016 ( \38393 , \38384 , \38388 );
or \U$38017 ( \38394 , \38392 , \38393 );
nand \U$38018 ( \38395 , \38374 , \38394 );
xor \U$38019 ( \38396 , \32331 , \32849 );
xnor \U$38020 ( \38397 , \38396 , \32319 );
xor \U$38021 ( \38398 , \38299 , \38336 );
and \U$38022 ( \38399 , \38398 , \38339 );
and \U$38023 ( \38400 , \38299 , \38336 );
or \U$38024 ( \38401 , \38399 , \38400 );
nand \U$38025 ( \38402 , \38397 , \38401 );
xor \U$38026 ( \38403 , \38384 , \38388 );
xor \U$38027 ( \38404 , \38403 , \38391 );
xor \U$38028 ( \38405 , \38235 , \38243 );
and \U$38029 ( \38406 , \38405 , \38271 );
and \U$38030 ( \38407 , \38235 , \38243 );
or \U$38031 ( \38408 , \38406 , \38407 );
nand \U$38032 ( \38409 , \38404 , \38408 );
and \U$38033 ( \38410 , \38372 , \38395 , \38402 , \38409 );
buf \U$38034 ( \38411 , \38410 );
nand \U$38035 ( \38412 , \38297 , \38411 );
not \U$38036 ( \38413 , \38412 );
nand \U$38037 ( \38414 , \32886 , \32901 );
not \U$38038 ( \38415 , \32317 );
not \U$38039 ( \38416 , \32853 );
nand \U$38040 ( \38417 , \38415 , \38416 );
nand \U$38041 ( \38418 , \32858 , \38417 );
nor \U$38042 ( \38419 , \38414 , \38418 );
and \U$38043 ( \38420 , \32904 , \38419 );
and \U$38044 ( \38421 , \33794 , \38420 );
nand \U$38045 ( \38422 , \38413 , \38421 , \33972 );
not \U$38046 ( \38423 , \37388 );
not \U$38047 ( \38424 , \37638 );
nand \U$38048 ( \38425 , \38423 , \38424 );
and \U$38049 ( \38426 , \37642 , \38425 );
not \U$38050 ( \38427 , \37667 );
and \U$38051 ( \38428 , \38426 , \37679 , \38427 );
buf \U$38052 ( \38429 , \36205 );
and \U$38053 ( \38430 , \38428 , \36639 , \36076 , \38429 );
and \U$38054 ( \38431 , \38430 , \38278 , \38410 );
xor \U$38055 ( \38432 , \37450 , \37460 );
xor \U$38056 ( \38433 , \38432 , \37471 );
xor \U$38057 ( \38434 , \37401 , \37425 );
xor \U$38058 ( \38435 , \38434 , \37436 );
xor \U$38059 ( \38436 , \38433 , \38435 );
not \U$38060 ( \38437 , \15729 );
not \U$38061 ( \38438 , \37574 );
or \U$38062 ( \38439 , \38437 , \38438 );
not \U$38063 ( \38440 , RIc225990_61);
not \U$38064 ( \38441 , \34175 );
or \U$38065 ( \38442 , \38440 , \38441 );
nand \U$38066 ( \38443 , \16532 , \12806 );
nand \U$38067 ( \38444 , \38442 , \38443 );
nand \U$38068 ( \38445 , \38444 , \15719 );
nand \U$38069 ( \38446 , \38439 , \38445 );
not \U$38070 ( \38447 , \38446 );
not \U$38071 ( \38448 , \11974 );
not \U$38072 ( \38449 , \37521 );
or \U$38073 ( \38450 , \38448 , \38449 );
not \U$38074 ( \38451 , RIc225b70_57);
not \U$38075 ( \38452 , \9912 );
or \U$38076 ( \38453 , \38451 , \38452 );
nand \U$38077 ( \38454 , \8952 , \11033 );
nand \U$38078 ( \38455 , \38453 , \38454 );
nand \U$38079 ( \38456 , \38455 , \11965 );
nand \U$38080 ( \38457 , \38450 , \38456 );
not \U$38081 ( \38458 , \38457 );
or \U$38082 ( \38459 , \38447 , \38458 );
or \U$38083 ( \38460 , \38457 , \38446 );
xor \U$38084 ( \38461 , \37530 , \37539 );
not \U$38085 ( \38462 , \9705 );
not \U$38086 ( \38463 , \37418 );
or \U$38087 ( \38464 , \38462 , \38463 );
not \U$38088 ( \38465 , RIc2262f0_41);
not \U$38089 ( \38466 , \15623 );
or \U$38090 ( \38467 , \38465 , \38466 );
nand \U$38091 ( \38468 , \21097 , \12937 );
nand \U$38092 ( \38469 , \38467 , \38468 );
nand \U$38093 ( \38470 , \38469 , \9689 );
nand \U$38094 ( \38471 , \38464 , \38470 );
xor \U$38095 ( \38472 , \38461 , \38471 );
not \U$38096 ( \38473 , \9129 );
not \U$38097 ( \38474 , \37546 );
or \U$38098 ( \38475 , \38473 , \38474 );
not \U$38099 ( \38476 , \19721 );
not \U$38100 ( \38477 , \12456 );
and \U$38101 ( \38478 , \38476 , \38477 );
and \U$38102 ( \38479 , \19721 , \12456 );
nor \U$38103 ( \38480 , \38478 , \38479 );
not \U$38104 ( \38481 , \38480 );
nand \U$38105 ( \38482 , \38481 , \9110 );
nand \U$38106 ( \38483 , \38475 , \38482 );
and \U$38107 ( \38484 , \38472 , \38483 );
and \U$38108 ( \38485 , \38461 , \38471 );
or \U$38109 ( \38486 , \38484 , \38485 );
nand \U$38110 ( \38487 , \38460 , \38486 );
nand \U$38111 ( \38488 , \38459 , \38487 );
xor \U$38112 ( \38489 , \38436 , \38488 );
xor \U$38113 ( \38490 , \37540 , \37550 );
xor \U$38114 ( \38491 , \38490 , \37562 );
not \U$38115 ( \38492 , \16891 );
not \U$38116 ( \38493 , RIc2258a0_63);
not \U$38117 ( \38494 , \23758 );
or \U$38118 ( \38495 , \38493 , \38494 );
nand \U$38119 ( \38496 , \6720 , \16880 );
nand \U$38120 ( \38497 , \38495 , \38496 );
not \U$38121 ( \38498 , \38497 );
or \U$38122 ( \38499 , \38492 , \38498 );
nand \U$38123 ( \38500 , \37496 , RIc225828_64);
nand \U$38124 ( \38501 , \38499 , \38500 );
xor \U$38125 ( \38502 , \38491 , \38501 );
not \U$38126 ( \38503 , \11697 );
not \U$38127 ( \38504 , RIc225c60_55);
not \U$38128 ( \38505 , \8910 );
or \U$38129 ( \38506 , \38504 , \38505 );
nand \U$38130 ( \38507 , \17744 , \11041 );
nand \U$38131 ( \38508 , \38506 , \38507 );
not \U$38132 ( \38509 , \38508 );
or \U$38133 ( \38510 , \38503 , \38509 );
nand \U$38134 ( \38511 , \37510 , \11038 );
nand \U$38135 ( \38512 , \38510 , \38511 );
xor \U$38136 ( \38513 , \38502 , \38512 );
not \U$38137 ( \38514 , \38513 );
not \U$38138 ( \38515 , \38514 );
xor \U$38139 ( \38516 , \38486 , \38446 );
xnor \U$38140 ( \38517 , \38516 , \38457 );
not \U$38141 ( \38518 , \38517 );
or \U$38142 ( \38519 , \38515 , \38518 );
not \U$38143 ( \38520 , \9934 );
not \U$38144 ( \38521 , RIc226110_45);
not \U$38145 ( \38522 , \20406 );
not \U$38146 ( \38523 , \38522 );
or \U$38147 ( \38524 , \38521 , \38523 );
not \U$38148 ( \38525 , \13498 );
nand \U$38149 ( \38526 , \38525 , \9379 );
nand \U$38150 ( \38527 , \38524 , \38526 );
not \U$38151 ( \38528 , \38527 );
or \U$38152 ( \38529 , \38520 , \38528 );
nand \U$38153 ( \38530 , \37560 , \9398 );
nand \U$38154 ( \38531 , \38529 , \38530 );
and \U$38155 ( \38532 , \16248 , \6306 );
not \U$38156 ( \38533 , \9705 );
not \U$38157 ( \38534 , \38469 );
or \U$38158 ( \38535 , \38533 , \38534 );
not \U$38159 ( \38536 , RIc2262f0_41);
not \U$38160 ( \38537 , \30827 );
or \U$38161 ( \38538 , \38536 , \38537 );
nand \U$38162 ( \38539 , \16482 , \12937 );
nand \U$38163 ( \38540 , \38538 , \38539 );
nand \U$38164 ( \38541 , \38540 , \9689 );
nand \U$38165 ( \38542 , \38535 , \38541 );
xor \U$38166 ( \38543 , \38532 , \38542 );
not \U$38167 ( \38544 , \9110 );
not \U$38168 ( \38545 , RIc226200_43);
not \U$38169 ( \38546 , \15630 );
or \U$38170 ( \38547 , \38545 , \38546 );
nand \U$38171 ( \38548 , \12844 , \9117 );
nand \U$38172 ( \38549 , \38547 , \38548 );
not \U$38173 ( \38550 , \38549 );
or \U$38174 ( \38551 , \38544 , \38550 );
not \U$38175 ( \38552 , \9128 );
or \U$38176 ( \38553 , \38480 , \38552 );
nand \U$38177 ( \38554 , \38551 , \38553 );
and \U$38178 ( \38555 , \38543 , \38554 );
and \U$38179 ( \38556 , \38532 , \38542 );
or \U$38180 ( \38557 , \38555 , \38556 );
xor \U$38181 ( \38558 , \38531 , \38557 );
not \U$38182 ( \38559 , \9619 );
not \U$38183 ( \38560 , RIc226020_47);
not \U$38184 ( \38561 , \13442 );
or \U$38185 ( \38562 , \38560 , \38561 );
nand \U$38186 ( \38563 , \9320 , \9624 );
nand \U$38187 ( \38564 , \38562 , \38563 );
not \U$38188 ( \38565 , \38564 );
or \U$38189 ( \38566 , \38559 , \38565 );
not \U$38190 ( \38567 , RIc226020_47);
not \U$38191 ( \38568 , \10360 );
or \U$38192 ( \38569 , \38567 , \38568 );
nand \U$38193 ( \38570 , \10086 , \9624 );
nand \U$38194 ( \38571 , \38569 , \38570 );
nand \U$38195 ( \38572 , \38571 , \9639 );
nand \U$38196 ( \38573 , \38566 , \38572 );
xor \U$38197 ( \38574 , \38558 , \38573 );
not \U$38198 ( \38575 , \16891 );
not \U$38199 ( \38576 , RIc2258a0_63);
not \U$38200 ( \38577 , \10142 );
or \U$38201 ( \38578 , \38576 , \38577 );
nand \U$38202 ( \38579 , \10141 , \16880 );
nand \U$38203 ( \38580 , \38578 , \38579 );
not \U$38204 ( \38581 , \38580 );
or \U$38205 ( \38582 , \38575 , \38581 );
nand \U$38206 ( \38583 , \38497 , RIc225828_64);
nand \U$38207 ( \38584 , \38582 , \38583 );
xor \U$38208 ( \38585 , \38574 , \38584 );
xor \U$38209 ( \38586 , \38532 , \38542 );
xor \U$38210 ( \38587 , \38586 , \38554 );
not \U$38211 ( \38588 , \9552 );
not \U$38212 ( \38589 , RIc225f30_49);
not \U$38213 ( \38590 , \9300 );
or \U$38214 ( \38591 , \38589 , \38590 );
nand \U$38215 ( \38592 , \21150 , \9541 );
nand \U$38216 ( \38593 , \38591 , \38592 );
not \U$38217 ( \38594 , \38593 );
or \U$38218 ( \38595 , \38588 , \38594 );
not \U$38219 ( \38596 , RIc225f30_49);
not \U$38220 ( \38597 , \9321 );
or \U$38221 ( \38598 , \38596 , \38597 );
nand \U$38222 ( \38599 , \9324 , \9549 );
nand \U$38223 ( \38600 , \38598 , \38599 );
nand \U$38224 ( \38601 , \38600 , \9532 );
nand \U$38225 ( \38602 , \38595 , \38601 );
xor \U$38226 ( \38603 , \38587 , \38602 );
not \U$38227 ( \38604 , \11038 );
not \U$38228 ( \38605 , RIc225c60_55);
not \U$38229 ( \38606 , \32810 );
or \U$38230 ( \38607 , \38605 , \38606 );
nand \U$38231 ( \38608 , \34371 , \11108 );
nand \U$38232 ( \38609 , \38607 , \38608 );
not \U$38233 ( \38610 , \38609 );
or \U$38234 ( \38611 , \38604 , \38610 );
not \U$38235 ( \38612 , RIc225c60_55);
not \U$38236 ( \38613 , \10645 );
or \U$38237 ( \38614 , \38612 , \38613 );
nand \U$38238 ( \38615 , \9050 , \8767 );
nand \U$38239 ( \38616 , \38614 , \38615 );
nand \U$38240 ( \38617 , \38616 , \11697 );
nand \U$38241 ( \38618 , \38611 , \38617 );
and \U$38242 ( \38619 , \38603 , \38618 );
and \U$38243 ( \38620 , \38587 , \38602 );
or \U$38244 ( \38621 , \38619 , \38620 );
and \U$38245 ( \38622 , \38585 , \38621 );
and \U$38246 ( \38623 , \38574 , \38584 );
or \U$38247 ( \38624 , \38622 , \38623 );
nand \U$38248 ( \38625 , \38519 , \38624 );
not \U$38249 ( \38626 , \38514 );
not \U$38250 ( \38627 , \38517 );
nand \U$38251 ( \38628 , \38626 , \38627 );
nand \U$38252 ( \38629 , \38625 , \38628 );
xor \U$38253 ( \38630 , \38489 , \38629 );
xor \U$38254 ( \38631 , \37402 , \37411 );
xor \U$38255 ( \38632 , \38631 , \37422 );
not \U$38256 ( \38633 , \12304 );
not \U$38257 ( \38634 , \37467 );
or \U$38258 ( \38635 , \38633 , \38634 );
nand \U$38259 ( \38636 , \38564 , \9641 );
nand \U$38260 ( \38637 , \38635 , \38636 );
xor \U$38261 ( \38638 , \38632 , \38637 );
not \U$38262 ( \38639 , \8788 );
not \U$38263 ( \38640 , \37486 );
or \U$38264 ( \38641 , \38639 , \38640 );
not \U$38265 ( \38642 , RIc225d50_53);
buf \U$38266 ( \38643 , \10643 );
not \U$38267 ( \38644 , \38643 );
or \U$38268 ( \38645 , \38642 , \38644 );
nand \U$38269 ( \38646 , \14608 , \8782 );
nand \U$38270 ( \38647 , \38645 , \38646 );
nand \U$38271 ( \38648 , \38647 , \9488 );
nand \U$38272 ( \38649 , \38641 , \38648 );
xor \U$38273 ( \38650 , \38638 , \38649 );
or \U$38274 ( \38651 , RIc226278_42, RIc226200_43);
nand \U$38275 ( \38652 , \38651 , \18357 );
and \U$38276 ( \38653 , RIc226278_42, RIc226200_43);
nor \U$38277 ( \38654 , \38653 , \6303 );
and \U$38278 ( \38655 , \38652 , \38654 );
not \U$38279 ( \38656 , \9705 );
not \U$38280 ( \38657 , \38540 );
or \U$38281 ( \38658 , \38656 , \38657 );
or \U$38282 ( \38659 , \18182 , \9822 );
or \U$38283 ( \38660 , \18181 , RIc2262f0_41);
nand \U$38284 ( \38661 , \38659 , \38660 );
nand \U$38285 ( \38662 , \38661 , \9689 );
nand \U$38286 ( \38663 , \38658 , \38662 );
and \U$38287 ( \38664 , \38655 , \38663 );
not \U$38288 ( \38665 , \9398 );
not \U$38289 ( \38666 , \38527 );
or \U$38290 ( \38667 , \38665 , \38666 );
not \U$38291 ( \38668 , RIc226110_45);
not \U$38292 ( \38669 , \16042 );
or \U$38293 ( \38670 , \38668 , \38669 );
nand \U$38294 ( \38671 , \20694 , \14660 );
nand \U$38295 ( \38672 , \38670 , \38671 );
nand \U$38296 ( \38673 , \38672 , \9934 );
nand \U$38297 ( \38674 , \38667 , \38673 );
xor \U$38298 ( \38675 , \38664 , \38674 );
not \U$38299 ( \38676 , \9619 );
not \U$38300 ( \38677 , \38571 );
or \U$38301 ( \38678 , \38676 , \38677 );
not \U$38302 ( \38679 , RIc226020_47);
not \U$38303 ( \38680 , \13211 );
or \U$38304 ( \38681 , \38679 , \38680 );
nand \U$38305 ( \38682 , \29423 , \9624 );
nand \U$38306 ( \38683 , \38681 , \38682 );
nand \U$38307 ( \38684 , \38683 , \9639 );
nand \U$38308 ( \38685 , \38678 , \38684 );
and \U$38309 ( \38686 , \38675 , \38685 );
and \U$38310 ( \38687 , \38664 , \38674 );
or \U$38311 ( \38688 , \38686 , \38687 );
not \U$38312 ( \38689 , \15729 );
not \U$38313 ( \38690 , \38444 );
or \U$38314 ( \38691 , \38689 , \38690 );
not \U$38315 ( \38692 , RIc225990_61);
not \U$38316 ( \38693 , \8857 );
or \U$38317 ( \38694 , \38692 , \38693 );
nand \U$38318 ( \38695 , \12727 , \12806 );
nand \U$38319 ( \38696 , \38694 , \38695 );
nand \U$38320 ( \38697 , \38696 , \15719 );
nand \U$38321 ( \38698 , \38691 , \38697 );
xor \U$38322 ( \38699 , \38688 , \38698 );
not \U$38323 ( \38700 , \11965 );
not \U$38324 ( \38701 , RIc225b70_57);
not \U$38325 ( \38702 , \8975 );
or \U$38326 ( \38703 , \38701 , \38702 );
nand \U$38327 ( \38704 , \8979 , \12475 );
nand \U$38328 ( \38705 , \38703 , \38704 );
not \U$38329 ( \38706 , \38705 );
or \U$38330 ( \38707 , \38700 , \38706 );
nand \U$38331 ( \38708 , \38455 , \11974 );
nand \U$38332 ( \38709 , \38707 , \38708 );
and \U$38333 ( \38710 , \38699 , \38709 );
and \U$38334 ( \38711 , \38688 , \38698 );
or \U$38335 ( \38712 , \38710 , \38711 );
xor \U$38336 ( \38713 , \38650 , \38712 );
xor \U$38337 ( \38714 , \38461 , \38471 );
xor \U$38338 ( \38715 , \38714 , \38483 );
not \U$38339 ( \38716 , \12532 );
not \U$38340 ( \38717 , \38508 );
or \U$38341 ( \38718 , \38716 , \38717 );
nand \U$38342 ( \38719 , \38609 , \11118 );
nand \U$38343 ( \38720 , \38718 , \38719 );
xor \U$38344 ( \38721 , \38715 , \38720 );
not \U$38345 ( \38722 , \12670 );
and \U$38346 ( \38723 , RIc225a80_59, \9897 );
not \U$38347 ( \38724 , RIc225a80_59);
and \U$38348 ( \38725 , \38724 , \20216 );
or \U$38349 ( \38726 , \38723 , \38725 );
not \U$38350 ( \38727 , \38726 );
or \U$38351 ( \38728 , \38722 , \38727 );
and \U$38352 ( \38729 , RIc225a80_59, \8810 );
not \U$38353 ( \38730 , RIc225a80_59);
and \U$38354 ( \38731 , \38730 , \10859 );
or \U$38355 ( \38732 , \38729 , \38731 );
nand \U$38356 ( \38733 , \38732 , \15164 );
nand \U$38357 ( \38734 , \38728 , \38733 );
and \U$38358 ( \38735 , \38721 , \38734 );
and \U$38359 ( \38736 , \38715 , \38720 );
or \U$38360 ( \38737 , \38735 , \38736 );
and \U$38361 ( \38738 , \38713 , \38737 );
and \U$38362 ( \38739 , \38650 , \38712 );
or \U$38363 ( \38740 , \38738 , \38739 );
xor \U$38364 ( \38741 , \38630 , \38740 );
xor \U$38365 ( \38742 , \38664 , \38674 );
xor \U$38366 ( \38743 , \38742 , \38685 );
not \U$38367 ( \38744 , \38743 );
not \U$38368 ( \38745 , \8777 );
not \U$38369 ( \38746 , RIc225d50_53);
not \U$38370 ( \38747 , \9250 );
or \U$38371 ( \38748 , \38746 , \38747 );
nand \U$38372 ( \38749 , \17018 , \8782 );
nand \U$38373 ( \38750 , \38748 , \38749 );
not \U$38374 ( \38751 , \38750 );
or \U$38375 ( \38752 , \38745 , \38751 );
not \U$38376 ( \38753 , RIc225d50_53);
not \U$38377 ( \38754 , \10814 );
or \U$38378 ( \38755 , \38753 , \38754 );
nand \U$38379 ( \38756 , \10110 , \8782 );
nand \U$38380 ( \38757 , \38755 , \38756 );
nand \U$38381 ( \38758 , \38757 , \8788 );
nand \U$38382 ( \38759 , \38752 , \38758 );
not \U$38383 ( \38760 , \11038 );
not \U$38384 ( \38761 , \38616 );
or \U$38385 ( \38762 , \38760 , \38761 );
not \U$38386 ( \38763 , RIc225c60_55);
not \U$38387 ( \38764 , \10654 );
or \U$38388 ( \38765 , \38763 , \38764 );
nand \U$38389 ( \38766 , \9072 , \16788 );
nand \U$38390 ( \38767 , \38765 , \38766 );
nand \U$38391 ( \38768 , \38767 , \11045 );
nand \U$38392 ( \38769 , \38762 , \38768 );
nor \U$38393 ( \38770 , \38759 , \38769 );
not \U$38394 ( \38771 , \9459 );
not \U$38395 ( \38772 , RIc225e40_51);
not \U$38396 ( \38773 , \10263 );
or \U$38397 ( \38774 , \38772 , \38773 );
nand \U$38398 ( \38775 , \30852 , \22140 );
nand \U$38399 ( \38776 , \38774 , \38775 );
not \U$38400 ( \38777 , \38776 );
or \U$38401 ( \38778 , \38771 , \38777 );
not \U$38402 ( \38779 , RIc225e40_51);
not \U$38403 ( \38780 , \13453 );
or \U$38404 ( \38781 , \38779 , \38780 );
nand \U$38405 ( \38782 , \10976 , \22140 );
nand \U$38406 ( \38783 , \38781 , \38782 );
nand \U$38407 ( \38784 , \38783 , \9444 );
nand \U$38408 ( \38785 , \38778 , \38784 );
not \U$38409 ( \38786 , \38785 );
or \U$38410 ( \38787 , \38770 , \38786 );
nand \U$38411 ( \38788 , \38769 , \38759 );
nand \U$38412 ( \38789 , \38787 , \38788 );
not \U$38413 ( \38790 , \38789 );
or \U$38414 ( \38791 , \38744 , \38790 );
or \U$38415 ( \38792 , \38789 , \38743 );
xor \U$38416 ( \38793 , \38655 , \38663 );
not \U$38417 ( \38794 , \9128 );
not \U$38418 ( \38795 , \38549 );
or \U$38419 ( \38796 , \38794 , \38795 );
not \U$38420 ( \38797 , RIc226200_43);
not \U$38421 ( \38798 , \20392 );
or \U$38422 ( \38799 , \38797 , \38798 );
nand \U$38423 ( \38800 , \21097 , \9117 );
nand \U$38424 ( \38801 , \38799 , \38800 );
nand \U$38425 ( \38802 , \38801 , \9110 );
nand \U$38426 ( \38803 , \38796 , \38802 );
xor \U$38427 ( \38804 , \38793 , \38803 );
not \U$38428 ( \38805 , \9619 );
not \U$38429 ( \38806 , \38683 );
or \U$38430 ( \38807 , \38805 , \38806 );
not \U$38431 ( \38808 , RIc226020_47);
not \U$38432 ( \38809 , \36273 );
or \U$38433 ( \38810 , \38808 , \38809 );
nand \U$38434 ( \38811 , \20406 , \9624 );
nand \U$38435 ( \38812 , \38810 , \38811 );
nand \U$38436 ( \38813 , \38812 , \9639 );
nand \U$38437 ( \38814 , \38807 , \38813 );
and \U$38438 ( \38815 , \38804 , \38814 );
and \U$38439 ( \38816 , \38793 , \38803 );
or \U$38440 ( \38817 , \38815 , \38816 );
nand \U$38441 ( \38818 , \38792 , \38817 );
nand \U$38442 ( \38819 , \38791 , \38818 );
xor \U$38443 ( \38820 , \38688 , \38698 );
xor \U$38444 ( \38821 , \38820 , \38709 );
xor \U$38445 ( \38822 , \38819 , \38821 );
xor \U$38446 ( \38823 , \38715 , \38720 );
xor \U$38447 ( \38824 , \38823 , \38734 );
and \U$38448 ( \38825 , \38822 , \38824 );
and \U$38449 ( \38826 , \38819 , \38821 );
or \U$38450 ( \38827 , \38825 , \38826 );
not \U$38451 ( \38828 , \38827 );
not \U$38452 ( \38829 , \38514 );
not \U$38453 ( \38830 , \38627 );
or \U$38454 ( \38831 , \38829 , \38830 );
nand \U$38455 ( \38832 , \38513 , \38517 );
nand \U$38456 ( \38833 , \38831 , \38832 );
and \U$38457 ( \38834 , \38833 , \38624 );
not \U$38458 ( \38835 , \38833 );
not \U$38459 ( \38836 , \38624 );
and \U$38460 ( \38837 , \38835 , \38836 );
nor \U$38461 ( \38838 , \38834 , \38837 );
not \U$38462 ( \38839 , \38838 );
nand \U$38463 ( \38840 , \38828 , \38839 );
not \U$38464 ( \38841 , \38840 );
xor \U$38465 ( \38842 , \38574 , \38584 );
xor \U$38466 ( \38843 , \38842 , \38621 );
not \U$38467 ( \38844 , \9398 );
not \U$38468 ( \38845 , \38672 );
or \U$38469 ( \38846 , \38844 , \38845 );
not \U$38470 ( \38847 , RIc226110_45);
not \U$38471 ( \38848 , \30815 );
or \U$38472 ( \38849 , \38847 , \38848 );
nand \U$38473 ( \38850 , \15443 , \14660 );
nand \U$38474 ( \38851 , \38849 , \38850 );
nand \U$38475 ( \38852 , \38851 , \9382 );
nand \U$38476 ( \38853 , \38846 , \38852 );
not \U$38477 ( \38854 , \38853 );
and \U$38478 ( \38855 , \38600 , \9552 );
not \U$38479 ( \38856 , RIc225f30_49);
not \U$38480 ( \38857 , \21172 );
or \U$38481 ( \38858 , \38856 , \38857 );
nand \U$38482 ( \38859 , \10086 , \9549 );
nand \U$38483 ( \38860 , \38858 , \38859 );
and \U$38484 ( \38861 , \38860 , \9532 );
nor \U$38485 ( \38862 , \38855 , \38861 );
nand \U$38486 ( \38863 , \38854 , \38862 );
not \U$38487 ( \38864 , \38863 );
and \U$38488 ( \38865 , \16248 , \9705 );
not \U$38489 ( \38866 , \9128 );
not \U$38490 ( \38867 , \38801 );
or \U$38491 ( \38868 , \38866 , \38867 );
not \U$38492 ( \38869 , RIc226200_43);
not \U$38493 ( \38870 , \16259 );
or \U$38494 ( \38871 , \38869 , \38870 );
nand \U$38495 ( \38872 , \16256 , \9117 );
nand \U$38496 ( \38873 , \38871 , \38872 );
not \U$38497 ( \38874 , \9109 );
nand \U$38498 ( \38875 , \38873 , \38874 );
nand \U$38499 ( \38876 , \38868 , \38875 );
xor \U$38500 ( \38877 , \38865 , \38876 );
not \U$38501 ( \38878 , \9382 );
not \U$38502 ( \38879 , RIc226110_45);
not \U$38503 ( \38880 , \12846 );
or \U$38504 ( \38881 , \38879 , \38880 );
nand \U$38505 ( \38882 , \18161 , \14390 );
nand \U$38506 ( \38883 , \38881 , \38882 );
not \U$38507 ( \38884 , \38883 );
or \U$38508 ( \38885 , \38878 , \38884 );
nand \U$38509 ( \38886 , \38851 , \9398 );
nand \U$38510 ( \38887 , \38885 , \38886 );
and \U$38511 ( \38888 , \38877 , \38887 );
and \U$38512 ( \38889 , \38865 , \38876 );
or \U$38513 ( \38890 , \38888 , \38889 );
not \U$38514 ( \38891 , \38890 );
or \U$38515 ( \38892 , \38864 , \38891 );
not \U$38516 ( \38893 , \38862 );
nand \U$38517 ( \38894 , \38893 , \38853 );
nand \U$38518 ( \38895 , \38892 , \38894 );
not \U$38519 ( \38896 , \38895 );
not \U$38520 ( \38897 , \9459 );
not \U$38521 ( \38898 , \38783 );
or \U$38522 ( \38899 , \38897 , \38898 );
not \U$38523 ( \38900 , RIc225e40_51);
not \U$38524 ( \38901 , \9250 );
or \U$38525 ( \38902 , \38900 , \38901 );
nand \U$38526 ( \38903 , \17014 , \12423 );
nand \U$38527 ( \38904 , \38902 , \38903 );
nand \U$38528 ( \38905 , \38904 , \9445 );
nand \U$38529 ( \38906 , \38899 , \38905 );
not \U$38530 ( \38907 , \8777 );
not \U$38531 ( \38908 , \38757 );
or \U$38532 ( \38909 , \38907 , \38908 );
not \U$38533 ( \38910 , RIc225d50_53);
not \U$38534 ( \38911 , \9073 );
or \U$38535 ( \38912 , \38910 , \38911 );
nand \U$38536 ( \38913 , \9072 , \8782 );
nand \U$38537 ( \38914 , \38912 , \38913 );
nand \U$38538 ( \38915 , \38914 , \9555 );
nand \U$38539 ( \38916 , \38909 , \38915 );
xor \U$38540 ( \38917 , \38906 , \38916 );
not \U$38541 ( \38918 , \11974 );
not \U$38542 ( \38919 , \38705 );
or \U$38543 ( \38920 , \38918 , \38919 );
not \U$38544 ( \38921 , RIc225b70_57);
not \U$38545 ( \38922 , \8910 );
or \U$38546 ( \38923 , \38921 , \38922 );
nand \U$38547 ( \38924 , \12406 , \11033 );
nand \U$38548 ( \38925 , \38923 , \38924 );
nand \U$38549 ( \38926 , \38925 , \11965 );
nand \U$38550 ( \38927 , \38920 , \38926 );
xor \U$38551 ( \38928 , \38917 , \38927 );
not \U$38552 ( \38929 , \38928 );
or \U$38553 ( \38930 , \38896 , \38929 );
or \U$38554 ( \38931 , \38928 , \38895 );
xor \U$38555 ( \38932 , \38793 , \38803 );
xor \U$38556 ( \38933 , \38932 , \38814 );
not \U$38557 ( \38934 , \9552 );
not \U$38558 ( \38935 , \38860 );
or \U$38559 ( \38936 , \38934 , \38935 );
not \U$38560 ( \38937 , RIc225f30_49);
not \U$38561 ( \38938 , \20702 );
or \U$38562 ( \38939 , \38937 , \38938 );
nand \U$38563 ( \38940 , \35896 , \11289 );
nand \U$38564 ( \38941 , \38939 , \38940 );
nand \U$38565 ( \38942 , \38941 , \9532 );
nand \U$38566 ( \38943 , \38936 , \38942 );
not \U$38567 ( \38944 , \38943 );
not \U$38568 ( \38945 , \38812 );
not \U$38569 ( \38946 , \38945 );
not \U$38570 ( \38947 , \22984 );
and \U$38571 ( \38948 , \38946 , \38947 );
not \U$38572 ( \38949 , \11607 );
not \U$38573 ( \38950 , \12756 );
or \U$38574 ( \38951 , \38949 , \38950 );
not \U$38575 ( \38952 , \20694 );
nand \U$38576 ( \38953 , \38952 , RIc226020_47);
nand \U$38577 ( \38954 , \38951 , \38953 );
and \U$38578 ( \38955 , \38954 , \9639 );
nor \U$38579 ( \38956 , \38948 , \38955 );
nand \U$38580 ( \38957 , \38944 , \38956 );
not \U$38581 ( \38958 , \38957 );
or \U$38582 ( \38959 , RIc226188_44, RIc226110_45);
nand \U$38583 ( \38960 , \38959 , \18357 );
and \U$38584 ( \38961 , RIc226188_44, RIc226110_45);
nor \U$38585 ( \38962 , \38961 , \12456 );
and \U$38586 ( \38963 , \38960 , \38962 );
not \U$38587 ( \38964 , \9128 );
not \U$38588 ( \38965 , \38873 );
or \U$38589 ( \38966 , \38964 , \38965 );
or \U$38590 ( \38967 , \16248 , \9125 );
or \U$38591 ( \38968 , \18356 , RIc226200_43);
nand \U$38592 ( \38969 , \38967 , \38968 );
nand \U$38593 ( \38970 , \38969 , \38874 );
nand \U$38594 ( \38971 , \38966 , \38970 );
and \U$38595 ( \38972 , \38963 , \38971 );
not \U$38596 ( \38973 , \38972 );
or \U$38597 ( \38974 , \38958 , \38973 );
not \U$38598 ( \38975 , \38956 );
nand \U$38599 ( \38976 , \38943 , \38975 );
nand \U$38600 ( \38977 , \38974 , \38976 );
xor \U$38601 ( \38978 , \38933 , \38977 );
not \U$38602 ( \38979 , \15164 );
and \U$38603 ( \38980 , RIc225a80_59, \31855 );
not \U$38604 ( \38981 , RIc225a80_59);
and \U$38605 ( \38982 , \38981 , \21867 );
or \U$38606 ( \38983 , \38980 , \38982 );
not \U$38607 ( \38984 , \38983 );
or \U$38608 ( \38985 , \38979 , \38984 );
and \U$38609 ( \38986 , RIc225a80_59, \13370 );
not \U$38610 ( \38987 , RIc225a80_59);
and \U$38611 ( \38988 , \38987 , \8952 );
or \U$38612 ( \38989 , \38986 , \38988 );
nand \U$38613 ( \38990 , \38989 , \12670 );
nand \U$38614 ( \38991 , \38985 , \38990 );
and \U$38615 ( \38992 , \38978 , \38991 );
and \U$38616 ( \38993 , \38933 , \38977 );
or \U$38617 ( \38994 , \38992 , \38993 );
nand \U$38618 ( \38995 , \38931 , \38994 );
nand \U$38619 ( \38996 , \38930 , \38995 );
xor \U$38620 ( \38997 , \38843 , \38996 );
xor \U$38621 ( \38998 , \38587 , \38602 );
xor \U$38622 ( \38999 , \38998 , \38618 );
not \U$38623 ( \39000 , RIc225b70_57);
not \U$38624 ( \39001 , \9212 );
or \U$38625 ( \39002 , \39000 , \39001 );
nand \U$38626 ( \39003 , \9216 , \12475 );
nand \U$38627 ( \39004 , \39002 , \39003 );
not \U$38628 ( \39005 , \39004 );
not \U$38629 ( \39006 , \39005 );
not \U$38630 ( \39007 , \29044 );
and \U$38631 ( \39008 , \39006 , \39007 );
and \U$38632 ( \39009 , \38925 , \11974 );
nor \U$38633 ( \39010 , \39008 , \39009 );
not \U$38634 ( \39011 , \39010 );
not \U$38635 ( \39012 , RIc2258a0_63);
not \U$38636 ( \39013 , \20674 );
or \U$38637 ( \39014 , \39012 , \39013 );
not \U$38638 ( \39015 , \10322 );
nand \U$38639 ( \39016 , \39015 , \15620 );
nand \U$38640 ( \39017 , \39014 , \39016 );
and \U$38641 ( \39018 , \39017 , \16891 );
not \U$38642 ( \39019 , RIc2258a0_63);
not \U$38643 ( \39020 , \34175 );
or \U$38644 ( \39021 , \39019 , \39020 );
nand \U$38645 ( \39022 , \17582 , \16880 );
nand \U$38646 ( \39023 , \39021 , \39022 );
and \U$38647 ( \39024 , \39023 , RIc225828_64);
nor \U$38648 ( \39025 , \39018 , \39024 );
not \U$38649 ( \39026 , \39025 );
or \U$38650 ( \39027 , \39011 , \39026 );
not \U$38651 ( \39028 , \15719 );
not \U$38652 ( \39029 , RIc225990_61);
not \U$38653 ( \39030 , \10858 );
or \U$38654 ( \39031 , \39029 , \39030 );
nand \U$38655 ( \39032 , \8811 , \10338 );
nand \U$38656 ( \39033 , \39031 , \39032 );
not \U$38657 ( \39034 , \39033 );
or \U$38658 ( \39035 , \39028 , \39034 );
not \U$38659 ( \39036 , RIc225990_61);
not \U$38660 ( \39037 , \20217 );
or \U$38661 ( \39038 , \39036 , \39037 );
nand \U$38662 ( \39039 , \22969 , \10338 );
nand \U$38663 ( \39040 , \39038 , \39039 );
nand \U$38664 ( \39041 , \39040 , \15729 );
nand \U$38665 ( \39042 , \39035 , \39041 );
nand \U$38666 ( \39043 , \39027 , \39042 );
or \U$38667 ( \39044 , \39010 , \39025 );
nand \U$38668 ( \39045 , \39043 , \39044 );
xor \U$38669 ( \39046 , \38999 , \39045 );
not \U$38670 ( \39047 , \15719 );
not \U$38671 ( \39048 , \39040 );
or \U$38672 ( \39049 , \39047 , \39048 );
nand \U$38673 ( \39050 , \38696 , \15729 );
nand \U$38674 ( \39051 , \39049 , \39050 );
not \U$38675 ( \39052 , \15164 );
not \U$38676 ( \39053 , \38989 );
or \U$38677 ( \39054 , \39052 , \39053 );
nand \U$38678 ( \39055 , \38732 , \12670 );
nand \U$38679 ( \39056 , \39054 , \39055 );
xor \U$38680 ( \39057 , \39051 , \39056 );
not \U$38681 ( \39058 , RIc225828_64);
not \U$38682 ( \39059 , \38580 );
or \U$38683 ( \39060 , \39058 , \39059 );
nand \U$38684 ( \39061 , \39023 , \16891 );
nand \U$38685 ( \39062 , \39060 , \39061 );
xor \U$38686 ( \39063 , \39057 , \39062 );
and \U$38687 ( \39064 , \39046 , \39063 );
and \U$38688 ( \39065 , \38999 , \39045 );
or \U$38689 ( \39066 , \39064 , \39065 );
and \U$38690 ( \39067 , \38997 , \39066 );
and \U$38691 ( \39068 , \38843 , \38996 );
or \U$38692 ( \39069 , \39067 , \39068 );
not \U$38693 ( \39070 , \39069 );
or \U$38694 ( \39071 , \38841 , \39070 );
nand \U$38695 ( \39072 , \38827 , \38838 );
nand \U$38696 ( \39073 , \39071 , \39072 );
xor \U$38697 ( \39074 , \38741 , \39073 );
not \U$38698 ( \39075 , \10445 );
not \U$38699 ( \39076 , RIc225f30_49);
not \U$38700 ( \39077 , \10975 );
or \U$38701 ( \39078 , \39076 , \39077 );
nand \U$38702 ( \39079 , \9275 , \9549 );
nand \U$38703 ( \39080 , \39078 , \39079 );
not \U$38704 ( \39081 , \39080 );
or \U$38705 ( \39082 , \39075 , \39081 );
nand \U$38706 ( \39083 , \37456 , \9552 );
nand \U$38707 ( \39084 , \39082 , \39083 );
not \U$38708 ( \39085 , \9459 );
not \U$38709 ( \39086 , RIc225e40_51);
not \U$38710 ( \39087 , \10111 );
or \U$38711 ( \39088 , \39086 , \39087 );
nand \U$38712 ( \39089 , \10110 , \12423 );
nand \U$38713 ( \39090 , \39088 , \39089 );
not \U$38714 ( \39091 , \39090 );
or \U$38715 ( \39092 , \39085 , \39091 );
nand \U$38716 ( \39093 , \37434 , \9445 );
nand \U$38717 ( \39094 , \39092 , \39093 );
xor \U$38718 ( \39095 , \39084 , \39094 );
not \U$38719 ( \39096 , \12670 );
and \U$38720 ( \39097 , RIc225a80_59, \12724 );
not \U$38721 ( \39098 , RIc225a80_59);
and \U$38722 ( \39099 , \39098 , \31447 );
or \U$38723 ( \39100 , \39097 , \39099 );
not \U$38724 ( \39101 , \39100 );
or \U$38725 ( \39102 , \39096 , \39101 );
nand \U$38726 ( \39103 , \38726 , \15164 );
nand \U$38727 ( \39104 , \39102 , \39103 );
and \U$38728 ( \39105 , \39095 , \39104 );
and \U$38729 ( \39106 , \39084 , \39094 );
or \U$38730 ( \39107 , \39105 , \39106 );
xor \U$38731 ( \39108 , \38512 , \38501 );
and \U$38732 ( \39109 , \39108 , \38491 );
and \U$38733 ( \39110 , \38512 , \38501 );
nor \U$38734 ( \39111 , \39109 , \39110 );
not \U$38735 ( \39112 , \39111 );
xor \U$38736 ( \39113 , \39107 , \39112 );
xor \U$38737 ( \39114 , \37525 , \37565 );
xor \U$38738 ( \39115 , \39114 , \37576 );
xor \U$38739 ( \39116 , \39113 , \39115 );
xor \U$38740 ( \39117 , \37512 , \37500 );
xor \U$38741 ( \39118 , \39117 , \37488 );
xor \U$38742 ( \39119 , \37248 , \37257 );
xor \U$38743 ( \39120 , \39119 , \37268 );
not \U$38744 ( \39121 , \15164 );
not \U$38745 ( \39122 , \39100 );
or \U$38746 ( \39123 , \39121 , \39122 );
nand \U$38747 ( \39124 , \37190 , \12670 );
nand \U$38748 ( \39125 , \39123 , \39124 );
xor \U$38749 ( \39126 , \39120 , \39125 );
xor \U$38750 ( \39127 , \38632 , \38637 );
and \U$38751 ( \39128 , \39127 , \38649 );
and \U$38752 ( \39129 , \38632 , \38637 );
or \U$38753 ( \39130 , \39128 , \39129 );
xor \U$38754 ( \39131 , \39126 , \39130 );
xor \U$38755 ( \39132 , \39118 , \39131 );
xor \U$38756 ( \39133 , \38531 , \38557 );
and \U$38757 ( \39134 , \39133 , \38573 );
and \U$38758 ( \39135 , \38531 , \38557 );
or \U$38759 ( \39136 , \39134 , \39135 );
not \U$38760 ( \39137 , \9444 );
not \U$38761 ( \39138 , \39090 );
or \U$38762 ( \39139 , \39137 , \39138 );
nand \U$38763 ( \39140 , \38904 , \9458 );
nand \U$38764 ( \39141 , \39139 , \39140 );
not \U$38765 ( \39142 , \9532 );
not \U$38766 ( \39143 , \38593 );
or \U$38767 ( \39144 , \39142 , \39143 );
nand \U$38768 ( \39145 , \39080 , \9552 );
nand \U$38769 ( \39146 , \39144 , \39145 );
xor \U$38770 ( \39147 , \39141 , \39146 );
not \U$38771 ( \39148 , \11577 );
not \U$38772 ( \39149 , \38647 );
or \U$38773 ( \39150 , \39148 , \39149 );
nand \U$38774 ( \39151 , \38914 , \8777 );
nand \U$38775 ( \39152 , \39150 , \39151 );
and \U$38776 ( \39153 , \39147 , \39152 );
and \U$38777 ( \39154 , \39141 , \39146 );
or \U$38778 ( \39155 , \39153 , \39154 );
xor \U$38779 ( \39156 , \39136 , \39155 );
xor \U$38780 ( \39157 , \39084 , \39094 );
xor \U$38781 ( \39158 , \39157 , \39104 );
and \U$38782 ( \39159 , \39156 , \39158 );
and \U$38783 ( \39160 , \39136 , \39155 );
or \U$38784 ( \39161 , \39159 , \39160 );
xor \U$38785 ( \39162 , \39132 , \39161 );
xor \U$38786 ( \39163 , \39116 , \39162 );
xor \U$38787 ( \39164 , \39141 , \39146 );
xor \U$38788 ( \39165 , \39164 , \39152 );
xor \U$38789 ( \39166 , \38906 , \38916 );
and \U$38790 ( \39167 , \39166 , \38927 );
and \U$38791 ( \39168 , \38906 , \38916 );
or \U$38792 ( \39169 , \39167 , \39168 );
xor \U$38793 ( \39170 , \39165 , \39169 );
xor \U$38794 ( \39171 , \39051 , \39056 );
and \U$38795 ( \39172 , \39171 , \39062 );
and \U$38796 ( \39173 , \39051 , \39056 );
or \U$38797 ( \39174 , \39172 , \39173 );
and \U$38798 ( \39175 , \39170 , \39174 );
and \U$38799 ( \39176 , \39165 , \39169 );
or \U$38800 ( \39177 , \39175 , \39176 );
xor \U$38801 ( \39178 , \39136 , \39155 );
xor \U$38802 ( \39179 , \39178 , \39158 );
or \U$38803 ( \39180 , \39177 , \39179 );
xor \U$38804 ( \39181 , \38650 , \38712 );
xor \U$38805 ( \39182 , \39181 , \38737 );
nand \U$38806 ( \39183 , \39180 , \39182 );
nand \U$38807 ( \39184 , \39177 , \39179 );
nand \U$38808 ( \39185 , \39183 , \39184 );
xor \U$38809 ( \39186 , \39163 , \39185 );
xnor \U$38810 ( \39187 , \39074 , \39186 );
xor \U$38811 ( \39188 , \39179 , \39177 );
xnor \U$38812 ( \39189 , \39188 , \39182 );
not \U$38813 ( \39190 , \39069 );
and \U$38814 ( \39191 , \38827 , \38839 );
not \U$38815 ( \39192 , \38827 );
and \U$38816 ( \39193 , \39192 , \38838 );
nor \U$38817 ( \39194 , \39191 , \39193 );
not \U$38818 ( \39195 , \39194 );
and \U$38819 ( \39196 , \39190 , \39195 );
and \U$38820 ( \39197 , \39069 , \39194 );
nor \U$38821 ( \39198 , \39196 , \39197 );
xor \U$38822 ( \39199 , \39189 , \39198 );
xor \U$38823 ( \39200 , \38819 , \38821 );
xor \U$38824 ( \39201 , \39200 , \38824 );
xor \U$38825 ( \39202 , \39165 , \39169 );
xor \U$38826 ( \39203 , \39202 , \39174 );
or \U$38827 ( \39204 , \39201 , \39203 );
xor \U$38828 ( \39205 , \38843 , \38996 );
xor \U$38829 ( \39206 , \39205 , \39066 );
nand \U$38830 ( \39207 , \39204 , \39206 );
nand \U$38831 ( \39208 , \39201 , \39203 );
and \U$38832 ( \39209 , \39207 , \39208 );
and \U$38833 ( \39210 , \39199 , \39209 );
and \U$38834 ( \39211 , \39189 , \39198 );
or \U$38835 ( \39212 , \39210 , \39211 );
nand \U$38836 ( \39213 , \39187 , \39212 );
not \U$38837 ( \39214 , \39213 );
xor \U$38838 ( \39215 , \39189 , \39198 );
xor \U$38839 ( \39216 , \39215 , \39209 );
xnor \U$38840 ( \39217 , \39201 , \39203 );
not \U$38841 ( \39218 , \39217 );
not \U$38842 ( \39219 , \39206 );
or \U$38843 ( \39220 , \39218 , \39219 );
or \U$38844 ( \39221 , \39206 , \39217 );
nand \U$38845 ( \39222 , \39220 , \39221 );
not \U$38846 ( \39223 , RIc225828_64);
not \U$38847 ( \39224 , \39017 );
or \U$38848 ( \39225 , \39223 , \39224 );
not \U$38849 ( \39226 , RIc2258a0_63);
not \U$38850 ( \39227 , \20217 );
or \U$38851 ( \39228 , \39226 , \39227 );
nand \U$38852 ( \39229 , \20216 , \15620 );
nand \U$38853 ( \39230 , \39228 , \39229 );
nand \U$38854 ( \39231 , \39230 , \16891 );
nand \U$38855 ( \39232 , \39225 , \39231 );
not \U$38856 ( \39233 , \12670 );
not \U$38857 ( \39234 , \38983 );
or \U$38858 ( \39235 , \39233 , \39234 );
and \U$38859 ( \39236 , RIc225a80_59, \12403 );
not \U$38860 ( \39237 , RIc225a80_59);
and \U$38861 ( \39238 , \39237 , \17744 );
or \U$38862 ( \39239 , \39236 , \39238 );
nand \U$38863 ( \39240 , \39239 , \15164 );
nand \U$38864 ( \39241 , \39235 , \39240 );
xor \U$38865 ( \39242 , \39232 , \39241 );
xor \U$38866 ( \39243 , \38963 , \38971 );
not \U$38867 ( \39244 , \9398 );
not \U$38868 ( \39245 , \38883 );
or \U$38869 ( \39246 , \39244 , \39245 );
not \U$38870 ( \39247 , RIc226110_45);
not \U$38871 ( \39248 , \30679 );
or \U$38872 ( \39249 , \39247 , \39248 );
nand \U$38873 ( \39250 , \13488 , \9379 );
nand \U$38874 ( \39251 , \39249 , \39250 );
nand \U$38875 ( \39252 , \39251 , \9382 );
nand \U$38876 ( \39253 , \39246 , \39252 );
xor \U$38877 ( \39254 , \39243 , \39253 );
not \U$38878 ( \39255 , \9552 );
not \U$38879 ( \39256 , \38941 );
or \U$38880 ( \39257 , \39255 , \39256 );
not \U$38881 ( \39258 , RIc225f30_49);
not \U$38882 ( \39259 , \13498 );
or \U$38883 ( \39260 , \39258 , \39259 );
not \U$38884 ( \39261 , \38522 );
nand \U$38885 ( \39262 , \39261 , \11289 );
nand \U$38886 ( \39263 , \39260 , \39262 );
nand \U$38887 ( \39264 , \39263 , \9534 );
nand \U$38888 ( \39265 , \39257 , \39264 );
and \U$38889 ( \39266 , \39254 , \39265 );
and \U$38890 ( \39267 , \39243 , \39253 );
or \U$38891 ( \39268 , \39266 , \39267 );
and \U$38892 ( \39269 , \39242 , \39268 );
and \U$38893 ( \39270 , \39232 , \39241 );
or \U$38894 ( \39271 , \39269 , \39270 );
not \U$38895 ( \39272 , \39271 );
not \U$38896 ( \39273 , \9444 );
not \U$38897 ( \39274 , \38776 );
or \U$38898 ( \39275 , \39273 , \39274 );
not \U$38899 ( \39276 , RIc225e40_51);
not \U$38900 ( \39277 , \9321 );
or \U$38901 ( \39278 , \39276 , \39277 );
nand \U$38902 ( \39279 , \9320 , \22140 );
nand \U$38903 ( \39280 , \39278 , \39279 );
nand \U$38904 ( \39281 , \39280 , \9459 );
nand \U$38905 ( \39282 , \39275 , \39281 );
not \U$38906 ( \39283 , \39282 );
not \U$38907 ( \39284 , \15719 );
not \U$38908 ( \39285 , RIc225990_61);
not \U$38909 ( \39286 , \13370 );
or \U$38910 ( \39287 , \39285 , \39286 );
nand \U$38911 ( \39288 , \8952 , \12806 );
nand \U$38912 ( \39289 , \39287 , \39288 );
not \U$38913 ( \39290 , \39289 );
or \U$38914 ( \39291 , \39284 , \39290 );
nand \U$38915 ( \39292 , \39033 , \15729 );
nand \U$38916 ( \39293 , \39291 , \39292 );
not \U$38917 ( \39294 , \39293 );
or \U$38918 ( \39295 , \39283 , \39294 );
or \U$38919 ( \39296 , \39293 , \39282 );
not \U$38920 ( \39297 , \8788 );
not \U$38921 ( \39298 , \38750 );
or \U$38922 ( \39299 , \39297 , \39298 );
not \U$38923 ( \39300 , \8776 );
not \U$38924 ( \39301 , RIc225d50_53);
not \U$38925 ( \39302 , \10975 );
or \U$38926 ( \39303 , \39301 , \39302 );
nand \U$38927 ( \39304 , \9275 , \8782 );
nand \U$38928 ( \39305 , \39303 , \39304 );
nand \U$38929 ( \39306 , \39300 , \39305 );
nand \U$38930 ( \39307 , \39299 , \39306 );
nand \U$38931 ( \39308 , \39296 , \39307 );
nand \U$38932 ( \39309 , \39295 , \39308 );
not \U$38933 ( \39310 , \39309 );
or \U$38934 ( \39311 , \39272 , \39310 );
or \U$38935 ( \39312 , \39309 , \39271 );
xor \U$38936 ( \39313 , \38933 , \38977 );
xor \U$38937 ( \39314 , \39313 , \38991 );
nand \U$38938 ( \39315 , \39312 , \39314 );
nand \U$38939 ( \39316 , \39311 , \39315 );
not \U$38940 ( \39317 , \39316 );
xor \U$38941 ( \39318 , \38895 , \38928 );
xnor \U$38942 ( \39319 , \39318 , \38994 );
not \U$38943 ( \39320 , \39319 );
not \U$38944 ( \39321 , \39320 );
or \U$38945 ( \39322 , \39317 , \39321 );
xor \U$38946 ( \39323 , \39042 , \39010 );
xnor \U$38947 ( \39324 , \39323 , \39025 );
not \U$38948 ( \39325 , \11038 );
not \U$38949 ( \39326 , RIc225c60_55);
not \U$38950 ( \39327 , \10814 );
or \U$38951 ( \39328 , \39326 , \39327 );
nand \U$38952 ( \39329 , \10110 , \11108 );
nand \U$38953 ( \39330 , \39328 , \39329 );
not \U$38954 ( \39331 , \39330 );
or \U$38955 ( \39332 , \39325 , \39331 );
not \U$38956 ( \39333 , RIc225c60_55);
not \U$38957 ( \39334 , \17015 );
or \U$38958 ( \39335 , \39333 , \39334 );
nand \U$38959 ( \39336 , \30878 , \11108 );
nand \U$38960 ( \39337 , \39335 , \39336 );
nand \U$38961 ( \39338 , \39337 , \11117 );
nand \U$38962 ( \39339 , \39332 , \39338 );
not \U$38963 ( \39340 , \9488 );
not \U$38964 ( \39341 , RIc225d50_53);
not \U$38965 ( \39342 , \9297 );
or \U$38966 ( \39343 , \39341 , \39342 );
nand \U$38967 ( \39344 , \30852 , \11391 );
nand \U$38968 ( \39345 , \39343 , \39344 );
not \U$38969 ( \39346 , \39345 );
or \U$38970 ( \39347 , \39340 , \39346 );
nand \U$38971 ( \39348 , \39305 , \8788 );
nand \U$38972 ( \39349 , \39347 , \39348 );
or \U$38973 ( \39350 , \39339 , \39349 );
not \U$38974 ( \39351 , \9445 );
not \U$38975 ( \39352 , \39280 );
or \U$38976 ( \39353 , \39351 , \39352 );
not \U$38977 ( \39354 , RIc225e40_51);
not \U$38978 ( \39355 , \10360 );
or \U$38979 ( \39356 , \39354 , \39355 );
nand \U$38980 ( \39357 , \10086 , \12423 );
nand \U$38981 ( \39358 , \39356 , \39357 );
nand \U$38982 ( \39359 , \39358 , \9459 );
nand \U$38983 ( \39360 , \39353 , \39359 );
nand \U$38984 ( \39361 , \39350 , \39360 );
nand \U$38985 ( \39362 , \39349 , \39339 );
and \U$38986 ( \39363 , \39361 , \39362 );
xor \U$38987 ( \39364 , \38972 , \38975 );
xnor \U$38988 ( \39365 , \39364 , \38943 );
nand \U$38989 ( \39366 , \39363 , \39365 );
not \U$38990 ( \39367 , \9619 );
not \U$38991 ( \39368 , \38954 );
or \U$38992 ( \39369 , \39367 , \39368 );
not \U$38993 ( \39370 , RIc226020_47);
not \U$38994 ( \39371 , \20519 );
or \U$38995 ( \39372 , \39370 , \39371 );
nand \U$38996 ( \39373 , \12825 , \9373 );
nand \U$38997 ( \39374 , \39372 , \39373 );
nand \U$38998 ( \39375 , \39374 , \9639 );
nand \U$38999 ( \39376 , \39369 , \39375 );
not \U$39000 ( \39377 , \11974 );
not \U$39001 ( \39378 , RIc225b70_57);
not \U$39002 ( \39379 , \38643 );
or \U$39003 ( \39380 , \39378 , \39379 );
nand \U$39004 ( \39381 , \14608 , \10074 );
nand \U$39005 ( \39382 , \39380 , \39381 );
not \U$39006 ( \39383 , \39382 );
or \U$39007 ( \39384 , \39377 , \39383 );
not \U$39008 ( \39385 , RIc225b70_57);
not \U$39009 ( \39386 , \9073 );
or \U$39010 ( \39387 , \39385 , \39386 );
nand \U$39011 ( \39388 , \9072 , \15262 );
nand \U$39012 ( \39389 , \39387 , \39388 );
nand \U$39013 ( \39390 , \39389 , \11965 );
nand \U$39014 ( \39391 , \39384 , \39390 );
or \U$39015 ( \39392 , \39376 , \39391 );
and \U$39016 ( \39393 , \18357 , \9128 );
not \U$39017 ( \39394 , \9398 );
not \U$39018 ( \39395 , \39251 );
or \U$39019 ( \39396 , \39394 , \39395 );
and \U$39020 ( \39397 , RIc226110_45, \32588 );
not \U$39021 ( \39398 , RIc226110_45);
and \U$39022 ( \39399 , \39398 , \20528 );
nor \U$39023 ( \39400 , \39397 , \39399 );
nand \U$39024 ( \39401 , \39400 , \9382 );
nand \U$39025 ( \39402 , \39396 , \39401 );
xor \U$39026 ( \39403 , \39393 , \39402 );
not \U$39027 ( \39404 , \9619 );
not \U$39028 ( \39405 , \39374 );
or \U$39029 ( \39406 , \39404 , \39405 );
not \U$39030 ( \39407 , RIc226020_47);
not \U$39031 ( \39408 , \15630 );
or \U$39032 ( \39409 , \39407 , \39408 );
nand \U$39033 ( \39410 , \15633 , \9624 );
nand \U$39034 ( \39411 , \39409 , \39410 );
nand \U$39035 ( \39412 , \39411 , \9639 );
nand \U$39036 ( \39413 , \39406 , \39412 );
and \U$39037 ( \39414 , \39403 , \39413 );
and \U$39038 ( \39415 , \39393 , \39402 );
or \U$39039 ( \39416 , \39414 , \39415 );
nand \U$39040 ( \39417 , \39392 , \39416 );
nand \U$39041 ( \39418 , \39391 , \39376 );
nand \U$39042 ( \39419 , \39417 , \39418 );
and \U$39043 ( \39420 , \39366 , \39419 );
nor \U$39044 ( \39421 , \39363 , \39365 );
nor \U$39045 ( \39422 , \39420 , \39421 );
nand \U$39046 ( \39423 , \39324 , \39422 );
not \U$39047 ( \39424 , \39423 );
xnor \U$39048 ( \39425 , \39307 , \39282 );
xor \U$39049 ( \39426 , \39293 , \39425 );
not \U$39050 ( \39427 , \39426 );
not \U$39051 ( \39428 , \39427 );
xor \U$39052 ( \39429 , \38865 , \38876 );
xor \U$39053 ( \39430 , \39429 , \38887 );
not \U$39054 ( \39431 , \11965 );
not \U$39055 ( \39432 , \39382 );
or \U$39056 ( \39433 , \39431 , \39432 );
nand \U$39057 ( \39434 , \39004 , \11974 );
nand \U$39058 ( \39435 , \39433 , \39434 );
xor \U$39059 ( \39436 , \39430 , \39435 );
not \U$39060 ( \39437 , \11038 );
not \U$39061 ( \39438 , \38767 );
or \U$39062 ( \39439 , \39437 , \39438 );
nand \U$39063 ( \39440 , \11117 , \39330 );
nand \U$39064 ( \39441 , \39439 , \39440 );
xor \U$39065 ( \39442 , \39436 , \39441 );
not \U$39066 ( \39443 , \39442 );
or \U$39067 ( \39444 , \39428 , \39443 );
not \U$39068 ( \39445 , \39442 );
not \U$39069 ( \39446 , \39445 );
not \U$39070 ( \39447 , \39426 );
or \U$39071 ( \39448 , \39446 , \39447 );
not \U$39072 ( \39449 , \20159 );
not \U$39073 ( \39450 , RIc2258a0_63);
not \U$39074 ( \39451 , \8810 );
or \U$39075 ( \39452 , \39450 , \39451 );
or \U$39076 ( \39453 , \31842 , RIc2258a0_63);
nand \U$39077 ( \39454 , \39452 , \39453 );
not \U$39078 ( \39455 , \39454 );
or \U$39079 ( \39456 , \39449 , \39455 );
nand \U$39080 ( \39457 , \39230 , RIc225828_64);
nand \U$39081 ( \39458 , \39456 , \39457 );
not \U$39082 ( \39459 , \20862 );
not \U$39083 ( \39460 , \39289 );
or \U$39084 ( \39461 , \39459 , \39460 );
not \U$39085 ( \39462 , RIc225990_61);
not \U$39086 ( \39463 , \11094 );
or \U$39087 ( \39464 , \39462 , \39463 );
nand \U$39088 ( \39465 , \11994 , \10338 );
nand \U$39089 ( \39466 , \39464 , \39465 );
nand \U$39090 ( \39467 , \39466 , \15719 );
nand \U$39091 ( \39468 , \39461 , \39467 );
or \U$39092 ( \39469 , \39458 , \39468 );
xor \U$39093 ( \39470 , \39243 , \39253 );
xor \U$39094 ( \39471 , \39470 , \39265 );
nand \U$39095 ( \39472 , \39469 , \39471 );
nand \U$39096 ( \39473 , \39458 , \39468 );
nand \U$39097 ( \39474 , \39472 , \39473 );
nand \U$39098 ( \39475 , \39448 , \39474 );
nand \U$39099 ( \39476 , \39444 , \39475 );
not \U$39100 ( \39477 , \39476 );
or \U$39101 ( \39478 , \39424 , \39477 );
not \U$39102 ( \39479 , \39422 );
not \U$39103 ( \39480 , \39324 );
nand \U$39104 ( \39481 , \39479 , \39480 );
nand \U$39105 ( \39482 , \39478 , \39481 );
not \U$39106 ( \39483 , \39316 );
nand \U$39107 ( \39484 , \39319 , \39483 );
nand \U$39108 ( \39485 , \39482 , \39484 );
nand \U$39109 ( \39486 , \39322 , \39485 );
not \U$39110 ( \39487 , \39486 );
xor \U$39111 ( \39488 , \38999 , \39045 );
xor \U$39112 ( \39489 , \39488 , \39063 );
xor \U$39113 ( \39490 , \38890 , \38853 );
xnor \U$39114 ( \39491 , \39490 , \38893 );
not \U$39115 ( \39492 , \39491 );
xor \U$39116 ( \39493 , \38769 , \38759 );
and \U$39117 ( \39494 , \39493 , \38786 );
not \U$39118 ( \39495 , \39493 );
and \U$39119 ( \39496 , \39495 , \38785 );
nor \U$39120 ( \39497 , \39494 , \39496 );
not \U$39121 ( \39498 , \39497 );
or \U$39122 ( \39499 , \39492 , \39498 );
xor \U$39123 ( \39500 , \39430 , \39435 );
and \U$39124 ( \39501 , \39500 , \39441 );
and \U$39125 ( \39502 , \39430 , \39435 );
or \U$39126 ( \39503 , \39501 , \39502 );
nand \U$39127 ( \39504 , \39499 , \39503 );
not \U$39128 ( \39505 , \39497 );
not \U$39129 ( \39506 , \39491 );
nand \U$39130 ( \39507 , \39505 , \39506 );
nand \U$39131 ( \39508 , \39504 , \39507 );
not \U$39132 ( \39509 , \39508 );
xor \U$39133 ( \39510 , \38817 , \38743 );
xnor \U$39134 ( \39511 , \39510 , \38789 );
nand \U$39135 ( \39512 , \39509 , \39511 );
and \U$39136 ( \39513 , \39489 , \39512 );
not \U$39137 ( \39514 , \39508 );
nor \U$39138 ( \39515 , \39514 , \39511 );
nor \U$39139 ( \39516 , \39513 , \39515 );
nand \U$39140 ( \39517 , \39487 , \39516 );
and \U$39141 ( \39518 , \39222 , \39517 );
not \U$39142 ( \39519 , \39486 );
nor \U$39143 ( \39520 , \39519 , \39516 );
nor \U$39144 ( \39521 , \39518 , \39520 );
nand \U$39145 ( \39522 , \39216 , \39521 );
not \U$39146 ( \39523 , \39522 );
not \U$39147 ( \39524 , \39222 );
not \U$39148 ( \39525 , \39486 );
not \U$39149 ( \39526 , \39516 );
and \U$39150 ( \39527 , \39525 , \39526 );
and \U$39151 ( \39528 , \39486 , \39516 );
nor \U$39152 ( \39529 , \39527 , \39528 );
not \U$39153 ( \39530 , \39529 );
and \U$39154 ( \39531 , \39524 , \39530 );
and \U$39155 ( \39532 , \39222 , \39529 );
nor \U$39156 ( \39533 , \39531 , \39532 );
not \U$39157 ( \39534 , \39508 );
not \U$39158 ( \39535 , \39511 );
and \U$39159 ( \39536 , \39534 , \39535 );
and \U$39160 ( \39537 , \39508 , \39511 );
nor \U$39161 ( \39538 , \39536 , \39537 );
xor \U$39162 ( \39539 , \39489 , \39538 );
not \U$39163 ( \39540 , \39320 );
not \U$39164 ( \39541 , \39483 );
or \U$39165 ( \39542 , \39540 , \39541 );
nand \U$39166 ( \39543 , \39319 , \39316 );
nand \U$39167 ( \39544 , \39542 , \39543 );
not \U$39168 ( \39545 , \39482 );
and \U$39169 ( \39546 , \39544 , \39545 );
not \U$39170 ( \39547 , \39544 );
and \U$39171 ( \39548 , \39547 , \39482 );
nor \U$39172 ( \39549 , \39546 , \39548 );
xor \U$39173 ( \39550 , \39539 , \39549 );
xor \U$39174 ( \39551 , \39506 , \39503 );
xor \U$39175 ( \39552 , \39551 , \39505 );
xor \U$39176 ( \39553 , \39309 , \39271 );
xor \U$39177 ( \39554 , \39553 , \39314 );
or \U$39178 ( \39555 , \39552 , \39554 );
not \U$39179 ( \39556 , \9552 );
not \U$39180 ( \39557 , \39263 );
or \U$39181 ( \39558 , \39556 , \39557 );
not \U$39182 ( \39559 , RIc225f30_49);
not \U$39183 ( \39560 , \20693 );
or \U$39184 ( \39561 , \39559 , \39560 );
nand \U$39185 ( \39562 , \12756 , \28163 );
nand \U$39186 ( \39563 , \39561 , \39562 );
nand \U$39187 ( \39564 , \39563 , \10445 );
nand \U$39188 ( \39565 , \39558 , \39564 );
not \U$39189 ( \39566 , \39565 );
not \U$39190 ( \39567 , \9444 );
not \U$39191 ( \39568 , \39358 );
or \U$39192 ( \39569 , \39567 , \39568 );
not \U$39193 ( \39570 , RIc225e40_51);
not \U$39194 ( \39571 , \27990 );
or \U$39195 ( \39572 , \39570 , \39571 );
nand \U$39196 ( \39573 , \35896 , \12423 );
nand \U$39197 ( \39574 , \39572 , \39573 );
nand \U$39198 ( \39575 , \39574 , \9458 );
nand \U$39199 ( \39576 , \39569 , \39575 );
not \U$39200 ( \39577 , \39576 );
nand \U$39201 ( \39578 , \39566 , \39577 );
or \U$39202 ( \39579 , RIc226098_46, RIc226020_47);
nand \U$39203 ( \39580 , \39579 , \18367 );
and \U$39204 ( \39581 , RIc226098_46, RIc226020_47);
nor \U$39205 ( \39582 , \39581 , \9100 );
and \U$39206 ( \39583 , \39580 , \39582 );
not \U$39207 ( \39584 , \9398 );
not \U$39208 ( \39585 , \39400 );
or \U$39209 ( \39586 , \39584 , \39585 );
and \U$39210 ( \39587 , \16248 , RIc226110_45);
not \U$39211 ( \39588 , \16248 );
and \U$39212 ( \39589 , \39588 , \14390 );
nor \U$39213 ( \39590 , \39587 , \39589 );
nand \U$39214 ( \39591 , \39590 , \9382 );
nand \U$39215 ( \39592 , \39586 , \39591 );
and \U$39216 ( \39593 , \39583 , \39592 );
and \U$39217 ( \39594 , \39578 , \39593 );
not \U$39218 ( \39595 , \39565 );
nor \U$39219 ( \39596 , \39595 , \39577 );
nor \U$39220 ( \39597 , \39594 , \39596 );
xor \U$39221 ( \39598 , \39416 , \39376 );
xnor \U$39222 ( \39599 , \39598 , \39391 );
xor \U$39223 ( \39600 , \39597 , \39599 );
and \U$39224 ( \39601 , \39239 , \18037 );
and \U$39225 ( \39602 , RIc225a80_59, \32810 );
not \U$39226 ( \39603 , RIc225a80_59);
and \U$39227 ( \39604 , \39603 , \32813 );
or \U$39228 ( \39605 , \39602 , \39604 );
not \U$39229 ( \39606 , \39605 );
nor \U$39230 ( \39607 , \39606 , \16439 );
nor \U$39231 ( \39608 , \39601 , \39607 );
and \U$39232 ( \39609 , \39600 , \39608 );
and \U$39233 ( \39610 , \39597 , \39599 );
or \U$39234 ( \39611 , \39609 , \39610 );
not \U$39235 ( \39612 , \39611 );
not \U$39236 ( \39613 , \39612 );
xor \U$39237 ( \39614 , \39232 , \39241 );
xor \U$39238 ( \39615 , \39614 , \39268 );
not \U$39239 ( \39616 , \39615 );
or \U$39240 ( \39617 , \39613 , \39616 );
or \U$39241 ( \39618 , \39615 , \39612 );
xor \U$39242 ( \39619 , \39393 , \39402 );
xor \U$39243 ( \39620 , \39619 , \39413 );
not \U$39244 ( \39621 , \11118 );
not \U$39245 ( \39622 , RIc225c60_55);
not \U$39246 ( \39623 , \9276 );
or \U$39247 ( \39624 , \39622 , \39623 );
nand \U$39248 ( \39625 , \36029 , \11108 );
nand \U$39249 ( \39626 , \39624 , \39625 );
not \U$39250 ( \39627 , \39626 );
or \U$39251 ( \39628 , \39621 , \39627 );
nand \U$39252 ( \39629 , \39337 , \13024 );
nand \U$39253 ( \39630 , \39628 , \39629 );
xor \U$39254 ( \39631 , \39620 , \39630 );
not \U$39255 ( \39632 , \11965 );
not \U$39256 ( \39633 , RIc225b70_57);
not \U$39257 ( \39634 , \13223 );
or \U$39258 ( \39635 , \39633 , \39634 );
nand \U$39259 ( \39636 , \10110 , \10074 );
nand \U$39260 ( \39637 , \39635 , \39636 );
not \U$39261 ( \39638 , \39637 );
or \U$39262 ( \39639 , \39632 , \39638 );
nand \U$39263 ( \39640 , \39389 , \11974 );
nand \U$39264 ( \39641 , \39639 , \39640 );
and \U$39265 ( \39642 , \39631 , \39641 );
and \U$39266 ( \39643 , \39620 , \39630 );
or \U$39267 ( \39644 , \39642 , \39643 );
not \U$39268 ( \39645 , \9488 );
not \U$39269 ( \39646 , RIc225d50_53);
not \U$39270 ( \39647 , \9321 );
or \U$39271 ( \39648 , \39646 , \39647 );
nand \U$39272 ( \39649 , \9320 , \11391 );
nand \U$39273 ( \39650 , \39648 , \39649 );
not \U$39274 ( \39651 , \39650 );
or \U$39275 ( \39652 , \39645 , \39651 );
nand \U$39276 ( \39653 , \39345 , \9555 );
nand \U$39277 ( \39654 , \39652 , \39653 );
not \U$39278 ( \39655 , \12670 );
not \U$39279 ( \39656 , \39605 );
or \U$39280 ( \39657 , \39655 , \39656 );
and \U$39281 ( \39658 , RIc225a80_59, \13465 );
not \U$39282 ( \39659 , RIc225a80_59);
and \U$39283 ( \39660 , \39659 , \10644 );
or \U$39284 ( \39661 , \39658 , \39660 );
nand \U$39285 ( \39662 , \39661 , \15164 );
nand \U$39286 ( \39663 , \39657 , \39662 );
xor \U$39287 ( \39664 , \39654 , \39663 );
not \U$39288 ( \39665 , \15719 );
not \U$39289 ( \39666 , RIc225990_61);
not \U$39290 ( \39667 , \8910 );
or \U$39291 ( \39668 , \39666 , \39667 );
nand \U$39292 ( \39669 , \34363 , \10338 );
nand \U$39293 ( \39670 , \39668 , \39669 );
not \U$39294 ( \39671 , \39670 );
or \U$39295 ( \39672 , \39665 , \39671 );
nand \U$39296 ( \39673 , \39466 , \20862 );
nand \U$39297 ( \39674 , \39672 , \39673 );
and \U$39298 ( \39675 , \39664 , \39674 );
and \U$39299 ( \39676 , \39654 , \39663 );
or \U$39300 ( \39677 , \39675 , \39676 );
xor \U$39301 ( \39678 , \39644 , \39677 );
xor \U$39302 ( \39679 , \39349 , \39339 );
xor \U$39303 ( \39680 , \39679 , \39360 );
and \U$39304 ( \39681 , \39678 , \39680 );
and \U$39305 ( \39682 , \39644 , \39677 );
or \U$39306 ( \39683 , \39681 , \39682 );
nand \U$39307 ( \39684 , \39618 , \39683 );
nand \U$39308 ( \39685 , \39617 , \39684 );
and \U$39309 ( \39686 , \39555 , \39685 );
and \U$39310 ( \39687 , \39552 , \39554 );
nor \U$39311 ( \39688 , \39686 , \39687 );
and \U$39312 ( \39689 , \39550 , \39688 );
and \U$39313 ( \39690 , \39539 , \39549 );
or \U$39314 ( \39691 , \39689 , \39690 );
nand \U$39315 ( \39692 , \39533 , \39691 );
xor \U$39316 ( \39693 , \39419 , \39363 );
xor \U$39317 ( \39694 , \39693 , \39365 );
not \U$39318 ( \39695 , \39694 );
not \U$39319 ( \39696 , \39695 );
xor \U$39320 ( \39697 , \39442 , \39427 );
xnor \U$39321 ( \39698 , \39697 , \39474 );
not \U$39322 ( \39699 , \39698 );
or \U$39323 ( \39700 , \39696 , \39699 );
xor \U$39324 ( \39701 , \39597 , \39599 );
xor \U$39325 ( \39702 , \39701 , \39608 );
not \U$39326 ( \39703 , \39702 );
not \U$39327 ( \39704 , \39703 );
xor \U$39328 ( \39705 , \39471 , \39468 );
xnor \U$39329 ( \39706 , \39705 , \39458 );
not \U$39330 ( \39707 , \39706 );
not \U$39331 ( \39708 , \39707 );
or \U$39332 ( \39709 , \39704 , \39708 );
not \U$39333 ( \39710 , \39702 );
not \U$39334 ( \39711 , \39706 );
or \U$39335 ( \39712 , \39710 , \39711 );
xor \U$39336 ( \39713 , \39583 , \39592 );
not \U$39337 ( \39714 , \9619 );
not \U$39338 ( \39715 , \39411 );
or \U$39339 ( \39716 , \39714 , \39715 );
and \U$39340 ( \39717 , \11607 , \17613 );
not \U$39341 ( \39718 , \11607 );
and \U$39342 ( \39719 , \39718 , \13488 );
nor \U$39343 ( \39720 , \39717 , \39719 );
nand \U$39344 ( \39721 , \39720 , \9639 );
nand \U$39345 ( \39722 , \39716 , \39721 );
xor \U$39346 ( \39723 , \39713 , \39722 );
not \U$39347 ( \39724 , \9552 );
not \U$39348 ( \39725 , \39563 );
or \U$39349 ( \39726 , \39724 , \39725 );
not \U$39350 ( \39727 , RIc225f30_49);
not \U$39351 ( \39728 , \30815 );
or \U$39352 ( \39729 , \39727 , \39728 );
nand \U$39353 ( \39730 , \19721 , \11289 );
nand \U$39354 ( \39731 , \39729 , \39730 );
nand \U$39355 ( \39732 , \39731 , \9532 );
nand \U$39356 ( \39733 , \39726 , \39732 );
and \U$39357 ( \39734 , \39723 , \39733 );
and \U$39358 ( \39735 , \39713 , \39722 );
or \U$39359 ( \39736 , \39734 , \39735 );
xor \U$39360 ( \39737 , \39593 , \39565 );
xnor \U$39361 ( \39738 , \39737 , \39577 );
xor \U$39362 ( \39739 , \39736 , \39738 );
not \U$39363 ( \39740 , \20159 );
not \U$39364 ( \39741 , RIc2258a0_63);
not \U$39365 ( \39742 , \13370 );
or \U$39366 ( \39743 , \39741 , \39742 );
not \U$39367 ( \39744 , RIc2258a0_63);
nand \U$39368 ( \39745 , \8952 , \39744 );
nand \U$39369 ( \39746 , \39743 , \39745 );
not \U$39370 ( \39747 , \39746 );
or \U$39371 ( \39748 , \39740 , \39747 );
nand \U$39372 ( \39749 , \39454 , RIc225828_64);
nand \U$39373 ( \39750 , \39748 , \39749 );
and \U$39374 ( \39751 , \39739 , \39750 );
and \U$39375 ( \39752 , \39736 , \39738 );
or \U$39376 ( \39753 , \39751 , \39752 );
nand \U$39377 ( \39754 , \39712 , \39753 );
nand \U$39378 ( \39755 , \39709 , \39754 );
nand \U$39379 ( \39756 , \39700 , \39755 );
not \U$39380 ( \39757 , \39698 );
nand \U$39381 ( \39758 , \39757 , \39694 );
nand \U$39382 ( \39759 , \39756 , \39758 );
not \U$39383 ( \39760 , \39759 );
buf \U$39384 ( \39761 , \39476 );
not \U$39385 ( \39762 , \39761 );
xor \U$39386 ( \39763 , \39480 , \39422 );
not \U$39387 ( \39764 , \39763 );
or \U$39388 ( \39765 , \39762 , \39764 );
or \U$39389 ( \39766 , \39763 , \39761 );
nand \U$39390 ( \39767 , \39765 , \39766 );
not \U$39391 ( \39768 , \39767 );
nand \U$39392 ( \39769 , \39760 , \39768 );
not \U$39393 ( \39770 , \39685 );
not \U$39394 ( \39771 , \39770 );
xor \U$39395 ( \39772 , \39552 , \39554 );
not \U$39396 ( \39773 , \39772 );
or \U$39397 ( \39774 , \39771 , \39773 );
or \U$39398 ( \39775 , \39772 , \39770 );
nand \U$39399 ( \39776 , \39774 , \39775 );
and \U$39400 ( \39777 , \39769 , \39776 );
and \U$39401 ( \39778 , \39767 , \39759 );
nor \U$39402 ( \39779 , \39777 , \39778 );
xor \U$39403 ( \39780 , \39539 , \39549 );
xor \U$39404 ( \39781 , \39780 , \39688 );
nor \U$39405 ( \39782 , \39779 , \39781 );
nand \U$39406 ( \39783 , \39692 , \39782 );
not \U$39407 ( \39784 , \39533 );
not \U$39408 ( \39785 , \39691 );
nand \U$39409 ( \39786 , \39784 , \39785 );
nand \U$39410 ( \39787 , \39783 , \39786 );
not \U$39411 ( \39788 , \39787 );
or \U$39412 ( \39789 , \39523 , \39788 );
not \U$39413 ( \39790 , \39216 );
not \U$39414 ( \39791 , \39521 );
nand \U$39415 ( \39792 , \39790 , \39791 );
nand \U$39416 ( \39793 , \39789 , \39792 );
not \U$39417 ( \39794 , \39793 );
or \U$39418 ( \39795 , \39214 , \39794 );
or \U$39419 ( \39796 , \39187 , \39212 );
nand \U$39420 ( \39797 , \39795 , \39796 );
nand \U$39421 ( \39798 , \39781 , \39779 );
and \U$39422 ( \39799 , \39692 , \39798 );
nand \U$39423 ( \39800 , \39799 , \39213 , \39522 );
xor \U$39424 ( \39801 , \39753 , \39706 );
xnor \U$39425 ( \39802 , \39801 , \39703 );
and \U$39426 ( \39803 , \18357 , \9398 );
not \U$39427 ( \39804 , \9619 );
not \U$39428 ( \39805 , \39720 );
or \U$39429 ( \39806 , \39804 , \39805 );
and \U$39430 ( \39807 , \9624 , \32587 );
not \U$39431 ( \39808 , \9624 );
and \U$39432 ( \39809 , \39808 , \16482 );
nor \U$39433 ( \39810 , \39807 , \39809 );
nand \U$39434 ( \39811 , \39810 , \9639 );
nand \U$39435 ( \39812 , \39806 , \39811 );
xor \U$39436 ( \39813 , \39803 , \39812 );
not \U$39437 ( \39814 , \9532 );
not \U$39438 ( \39815 , RIc225f30_49);
not \U$39439 ( \39816 , \12846 );
or \U$39440 ( \39817 , \39815 , \39816 );
nand \U$39441 ( \39818 , \18161 , \9549 );
nand \U$39442 ( \39819 , \39817 , \39818 );
not \U$39443 ( \39820 , \39819 );
or \U$39444 ( \39821 , \39814 , \39820 );
nand \U$39445 ( \39822 , \39731 , \9552 );
nand \U$39446 ( \39823 , \39821 , \39822 );
and \U$39447 ( \39824 , \39813 , \39823 );
and \U$39448 ( \39825 , \39803 , \39812 );
or \U$39449 ( \39826 , \39824 , \39825 );
not \U$39450 ( \39827 , \9444 );
not \U$39451 ( \39828 , \39574 );
or \U$39452 ( \39829 , \39827 , \39828 );
not \U$39453 ( \39830 , RIc225e40_51);
not \U$39454 ( \39831 , \13498 );
or \U$39455 ( \39832 , \39830 , \39831 );
nand \U$39456 ( \39833 , \37397 , \12423 );
nand \U$39457 ( \39834 , \39832 , \39833 );
nand \U$39458 ( \39835 , \39834 , \9459 );
nand \U$39459 ( \39836 , \39829 , \39835 );
xor \U$39460 ( \39837 , \39826 , \39836 );
not \U$39461 ( \39838 , \11965 );
not \U$39462 ( \39839 , RIc225b70_57);
not \U$39463 ( \39840 , \11488 );
or \U$39464 ( \39841 , \39839 , \39840 );
nand \U$39465 ( \39842 , \35479 , \12475 );
nand \U$39466 ( \39843 , \39841 , \39842 );
not \U$39467 ( \39844 , \39843 );
or \U$39468 ( \39845 , \39838 , \39844 );
nand \U$39469 ( \39846 , \39637 , \15267 );
nand \U$39470 ( \39847 , \39845 , \39846 );
xor \U$39471 ( \39848 , \39837 , \39847 );
not \U$39472 ( \39849 , \39848 );
not \U$39473 ( \39850 , RIc225828_64);
not \U$39474 ( \39851 , \39746 );
or \U$39475 ( \39852 , \39850 , \39851 );
not \U$39476 ( \39853 , RIc2258a0_63);
not \U$39477 ( \39854 , \11094 );
or \U$39478 ( \39855 , \39853 , \39854 );
nand \U$39479 ( \39856 , \11994 , \15620 );
nand \U$39480 ( \39857 , \39855 , \39856 );
nand \U$39481 ( \39858 , \39857 , \20159 );
nand \U$39482 ( \39859 , \39852 , \39858 );
not \U$39483 ( \39860 , \39859 );
or \U$39484 ( \39861 , \39849 , \39860 );
or \U$39485 ( \39862 , \39859 , \39848 );
xor \U$39486 ( \39863 , \39803 , \39812 );
xor \U$39487 ( \39864 , \39863 , \39823 );
not \U$39488 ( \39865 , \11965 );
not \U$39489 ( \39866 , RIc225b70_57);
not \U$39490 ( \39867 , \10975 );
or \U$39491 ( \39868 , \39866 , \39867 );
nand \U$39492 ( \39869 , \9275 , \15262 );
nand \U$39493 ( \39870 , \39868 , \39869 );
not \U$39494 ( \39871 , \39870 );
or \U$39495 ( \39872 , \39865 , \39871 );
nand \U$39496 ( \39873 , \39843 , \11974 );
nand \U$39497 ( \39874 , \39872 , \39873 );
xor \U$39498 ( \39875 , \39864 , \39874 );
not \U$39499 ( \39876 , \11038 );
not \U$39500 ( \39877 , RIc225c60_55);
not \U$39501 ( \39878 , \10263 );
or \U$39502 ( \39879 , \39877 , \39878 );
nand \U$39503 ( \39880 , \16998 , \11108 );
nand \U$39504 ( \39881 , \39879 , \39880 );
not \U$39505 ( \39882 , \39881 );
or \U$39506 ( \39883 , \39876 , \39882 );
not \U$39507 ( \39884 , RIc225c60_55);
not \U$39508 ( \39885 , \9321 );
or \U$39509 ( \39886 , \39884 , \39885 );
nand \U$39510 ( \39887 , \9320 , \11041 );
nand \U$39511 ( \39888 , \39886 , \39887 );
nand \U$39512 ( \39889 , \39888 , \11117 );
nand \U$39513 ( \39890 , \39883 , \39889 );
and \U$39514 ( \39891 , \39875 , \39890 );
and \U$39515 ( \39892 , \39864 , \39874 );
or \U$39516 ( \39893 , \39891 , \39892 );
nand \U$39517 ( \39894 , \39862 , \39893 );
nand \U$39518 ( \39895 , \39861 , \39894 );
not \U$39519 ( \39896 , \15164 );
and \U$39520 ( \39897 , RIc225a80_59, \10652 );
not \U$39521 ( \39898 , RIc225a80_59);
and \U$39522 ( \39899 , \39898 , \32612 );
or \U$39523 ( \39900 , \39897 , \39899 );
not \U$39524 ( \39901 , \39900 );
or \U$39525 ( \39902 , \39896 , \39901 );
nand \U$39526 ( \39903 , \39661 , \12670 );
nand \U$39527 ( \39904 , \39902 , \39903 );
not \U$39528 ( \39905 , \11045 );
not \U$39529 ( \39906 , \39881 );
or \U$39530 ( \39907 , \39905 , \39906 );
nand \U$39531 ( \39908 , \39626 , \11038 );
nand \U$39532 ( \39909 , \39907 , \39908 );
nor \U$39533 ( \39910 , \39904 , \39909 );
and \U$39534 ( \39911 , \39650 , \9555 );
not \U$39535 ( \39912 , RIc225d50_53);
not \U$39536 ( \39913 , \10360 );
or \U$39537 ( \39914 , \39912 , \39913 );
nand \U$39538 ( \39915 , \10086 , \8782 );
nand \U$39539 ( \39916 , \39914 , \39915 );
and \U$39540 ( \39917 , \39916 , \8777 );
nor \U$39541 ( \39918 , \39911 , \39917 );
or \U$39542 ( \39919 , \39910 , \39918 );
nand \U$39543 ( \39920 , \39904 , \39909 );
nand \U$39544 ( \39921 , \39919 , \39920 );
xor \U$39545 ( \39922 , \39826 , \39836 );
and \U$39546 ( \39923 , \39922 , \39847 );
and \U$39547 ( \39924 , \39826 , \39836 );
or \U$39548 ( \39925 , \39923 , \39924 );
xor \U$39549 ( \39926 , \39921 , \39925 );
xor \U$39550 ( \39927 , \39620 , \39630 );
xor \U$39551 ( \39928 , \39927 , \39641 );
xor \U$39552 ( \39929 , \39926 , \39928 );
xor \U$39553 ( \39930 , \39895 , \39929 );
xor \U$39554 ( \39931 , \39904 , \39909 );
xnor \U$39555 ( \39932 , \39931 , \39918 );
xor \U$39556 ( \39933 , \39713 , \39722 );
xor \U$39557 ( \39934 , \39933 , \39733 );
or \U$39558 ( \39935 , RIc225fa8_48, RIc225f30_49);
nand \U$39559 ( \39936 , \39935 , \18367 );
and \U$39560 ( \39937 , RIc225fa8_48, RIc225f30_49);
nor \U$39561 ( \39938 , \39937 , \9373 );
and \U$39562 ( \39939 , \39936 , \39938 );
not \U$39563 ( \39940 , \9619 );
not \U$39564 ( \39941 , \39810 );
or \U$39565 ( \39942 , \39940 , \39941 );
and \U$39566 ( \39943 , \18366 , RIc226020_47);
and \U$39567 ( \39944 , \18357 , \11607 );
nor \U$39568 ( \39945 , \39943 , \39944 );
or \U$39569 ( \39946 , \39945 , \9640 );
nand \U$39570 ( \39947 , \39942 , \39946 );
and \U$39571 ( \39948 , \39939 , \39947 );
not \U$39572 ( \39949 , \9459 );
and \U$39573 ( \39950 , \16042 , RIc225e40_51);
not \U$39574 ( \39951 , \16042 );
and \U$39575 ( \39952 , \39951 , \12423 );
or \U$39576 ( \39953 , \39950 , \39952 );
not \U$39577 ( \39954 , \39953 );
or \U$39578 ( \39955 , \39949 , \39954 );
nand \U$39579 ( \39956 , \39834 , \9444 );
nand \U$39580 ( \39957 , \39955 , \39956 );
xor \U$39581 ( \39958 , \39948 , \39957 );
not \U$39582 ( \39959 , \8788 );
not \U$39583 ( \39960 , \39916 );
or \U$39584 ( \39961 , \39959 , \39960 );
and \U$39585 ( \39962 , \13211 , RIc225d50_53);
not \U$39586 ( \39963 , \13211 );
and \U$39587 ( \39964 , \39963 , \8772 );
or \U$39588 ( \39965 , \39962 , \39964 );
nand \U$39589 ( \39966 , \39965 , \8777 );
nand \U$39590 ( \39967 , \39961 , \39966 );
and \U$39591 ( \39968 , \39958 , \39967 );
and \U$39592 ( \39969 , \39948 , \39957 );
or \U$39593 ( \39970 , \39968 , \39969 );
xor \U$39594 ( \39971 , \39934 , \39970 );
not \U$39595 ( \39972 , \20862 );
not \U$39596 ( \39973 , \39670 );
or \U$39597 ( \39974 , \39972 , \39973 );
not \U$39598 ( \39975 , RIc225990_61);
not \U$39599 ( \39976 , \8925 );
or \U$39600 ( \39977 , \39975 , \39976 );
not \U$39601 ( \39978 , \32810 );
nand \U$39602 ( \39979 , \39978 , \12806 );
nand \U$39603 ( \39980 , \39977 , \39979 );
nand \U$39604 ( \39981 , \39980 , \15719 );
nand \U$39605 ( \39982 , \39974 , \39981 );
xor \U$39606 ( \39983 , \39971 , \39982 );
xor \U$39607 ( \39984 , \39932 , \39983 );
not \U$39608 ( \39985 , \12670 );
not \U$39609 ( \39986 , \39900 );
or \U$39610 ( \39987 , \39985 , \39986 );
and \U$39611 ( \39988 , RIc225a80_59, \13223 );
not \U$39612 ( \39989 , RIc225a80_59);
and \U$39613 ( \39990 , \39989 , \10110 );
or \U$39614 ( \39991 , \39988 , \39990 );
nand \U$39615 ( \39992 , \39991 , \15164 );
nand \U$39616 ( \39993 , \39987 , \39992 );
not \U$39617 ( \39994 , \15729 );
not \U$39618 ( \39995 , \39980 );
or \U$39619 ( \39996 , \39994 , \39995 );
not \U$39620 ( \39997 , RIc225990_61);
not \U$39621 ( \39998 , \38643 );
or \U$39622 ( \39999 , \39997 , \39998 );
nand \U$39623 ( \40000 , \14608 , \10338 );
nand \U$39624 ( \40001 , \39999 , \40000 );
nand \U$39625 ( \40002 , \40001 , \15719 );
nand \U$39626 ( \40003 , \39996 , \40002 );
xor \U$39627 ( \40004 , \39993 , \40003 );
not \U$39628 ( \40005 , \16891 );
not \U$39629 ( \40006 , RIc2258a0_63);
not \U$39630 ( \40007 , \8910 );
or \U$39631 ( \40008 , \40006 , \40007 );
nand \U$39632 ( \40009 , \34363 , \16880 );
nand \U$39633 ( \40010 , \40008 , \40009 );
not \U$39634 ( \40011 , \40010 );
or \U$39635 ( \40012 , \40005 , \40011 );
nand \U$39636 ( \40013 , \39857 , RIc225828_64);
nand \U$39637 ( \40014 , \40012 , \40013 );
and \U$39638 ( \40015 , \40004 , \40014 );
and \U$39639 ( \40016 , \39993 , \40003 );
or \U$39640 ( \40017 , \40015 , \40016 );
and \U$39641 ( \40018 , \39984 , \40017 );
and \U$39642 ( \40019 , \39932 , \39983 );
or \U$39643 ( \40020 , \40018 , \40019 );
and \U$39644 ( \40021 , \39930 , \40020 );
and \U$39645 ( \40022 , \39895 , \39929 );
or \U$39646 ( \40023 , \40021 , \40022 );
xor \U$39647 ( \40024 , \39802 , \40023 );
xor \U$39648 ( \40025 , \39921 , \39925 );
and \U$39649 ( \40026 , \40025 , \39928 );
and \U$39650 ( \40027 , \39921 , \39925 );
or \U$39651 ( \40028 , \40026 , \40027 );
xor \U$39652 ( \40029 , \39644 , \39677 );
xor \U$39653 ( \40030 , \40029 , \39680 );
xor \U$39654 ( \40031 , \40028 , \40030 );
xor \U$39655 ( \40032 , \39654 , \39663 );
xor \U$39656 ( \40033 , \40032 , \39674 );
not \U$39657 ( \40034 , \40033 );
not \U$39658 ( \40035 , \40034 );
xor \U$39659 ( \40036 , \39934 , \39970 );
and \U$39660 ( \40037 , \40036 , \39982 );
and \U$39661 ( \40038 , \39934 , \39970 );
or \U$39662 ( \40039 , \40037 , \40038 );
not \U$39663 ( \40040 , \40039 );
not \U$39664 ( \40041 , \40040 );
or \U$39665 ( \40042 , \40035 , \40041 );
xor \U$39666 ( \40043 , \39736 , \39738 );
xor \U$39667 ( \40044 , \40043 , \39750 );
nand \U$39668 ( \40045 , \40042 , \40044 );
nand \U$39669 ( \40046 , \40039 , \40033 );
nand \U$39670 ( \40047 , \40045 , \40046 );
xor \U$39671 ( \40048 , \40031 , \40047 );
xor \U$39672 ( \40049 , \40024 , \40048 );
and \U$39673 ( \40050 , \40039 , \40033 );
not \U$39674 ( \40051 , \40039 );
and \U$39675 ( \40052 , \40051 , \40034 );
nor \U$39676 ( \40053 , \40050 , \40052 );
xor \U$39677 ( \40054 , \40053 , \40044 );
xor \U$39678 ( \40055 , \39895 , \39929 );
xor \U$39679 ( \40056 , \40055 , \40020 );
xor \U$39680 ( \40057 , \40054 , \40056 );
xor \U$39681 ( \40058 , \39939 , \39947 );
not \U$39682 ( \40059 , \9552 );
not \U$39683 ( \40060 , \39819 );
or \U$39684 ( \40061 , \40059 , \40060 );
and \U$39685 ( \40062 , \9549 , \21097 );
not \U$39686 ( \40063 , \9549 );
and \U$39687 ( \40064 , \40063 , \15623 );
nor \U$39688 ( \40065 , \40062 , \40064 );
or \U$39689 ( \40066 , \40065 , \9533 );
nand \U$39690 ( \40067 , \40061 , \40066 );
xor \U$39691 ( \40068 , \40058 , \40067 );
not \U$39692 ( \40069 , \8777 );
not \U$39693 ( \40070 , RIc225d50_53);
not \U$39694 ( \40071 , \37397 );
not \U$39695 ( \40072 , \40071 );
or \U$39696 ( \40073 , \40070 , \40072 );
not \U$39697 ( \40074 , \21084 );
nand \U$39698 ( \40075 , \40074 , \11391 );
nand \U$39699 ( \40076 , \40073 , \40075 );
not \U$39700 ( \40077 , \40076 );
or \U$39701 ( \40078 , \40069 , \40077 );
nand \U$39702 ( \40079 , \39965 , \8788 );
nand \U$39703 ( \40080 , \40078 , \40079 );
and \U$39704 ( \40081 , \40068 , \40080 );
and \U$39705 ( \40082 , \40058 , \40067 );
or \U$39706 ( \40083 , \40081 , \40082 );
xor \U$39707 ( \40084 , \39948 , \39957 );
xor \U$39708 ( \40085 , \40084 , \39967 );
xor \U$39709 ( \40086 , \40083 , \40085 );
not \U$39710 ( \40087 , \9445 );
not \U$39711 ( \40088 , \39953 );
or \U$39712 ( \40089 , \40087 , \40088 );
not \U$39713 ( \40090 , RIc225e40_51);
not \U$39714 ( \40091 , \18167 );
or \U$39715 ( \40092 , \40090 , \40091 );
not \U$39716 ( \40093 , \30815 );
nand \U$39717 ( \40094 , \40093 , \9450 );
nand \U$39718 ( \40095 , \40092 , \40094 );
nand \U$39719 ( \40096 , \40095 , \9459 );
nand \U$39720 ( \40097 , \40089 , \40096 );
and \U$39721 ( \40098 , \18367 , \9619 );
not \U$39722 ( \40099 , \9532 );
not \U$39723 ( \40100 , RIc225f30_49);
not \U$39724 ( \40101 , \30827 );
or \U$39725 ( \40102 , \40100 , \40101 );
nand \U$39726 ( \40103 , \16256 , \11289 );
nand \U$39727 ( \40104 , \40102 , \40103 );
not \U$39728 ( \40105 , \40104 );
or \U$39729 ( \40106 , \40099 , \40105 );
or \U$39730 ( \40107 , \40065 , \23415 );
nand \U$39731 ( \40108 , \40106 , \40107 );
xor \U$39732 ( \40109 , \40098 , \40108 );
not \U$39733 ( \40110 , \9458 );
not \U$39734 ( \40111 , RIc225e40_51);
not \U$39735 ( \40112 , \15630 );
or \U$39736 ( \40113 , \40111 , \40112 );
nand \U$39737 ( \40114 , \18161 , \22140 );
nand \U$39738 ( \40115 , \40113 , \40114 );
not \U$39739 ( \40116 , \40115 );
or \U$39740 ( \40117 , \40110 , \40116 );
nand \U$39741 ( \40118 , \40095 , \9444 );
nand \U$39742 ( \40119 , \40117 , \40118 );
and \U$39743 ( \40120 , \40109 , \40119 );
and \U$39744 ( \40121 , \40098 , \40108 );
or \U$39745 ( \40122 , \40120 , \40121 );
xor \U$39746 ( \40123 , \40097 , \40122 );
not \U$39747 ( \40124 , \11974 );
not \U$39748 ( \40125 , \39870 );
or \U$39749 ( \40126 , \40124 , \40125 );
not \U$39750 ( \40127 , RIc225b70_57);
not \U$39751 ( \40128 , \30069 );
or \U$39752 ( \40129 , \40127 , \40128 );
nand \U$39753 ( \40130 , \9299 , \15262 );
nand \U$39754 ( \40131 , \40129 , \40130 );
nand \U$39755 ( \40132 , \40131 , \11965 );
nand \U$39756 ( \40133 , \40126 , \40132 );
and \U$39757 ( \40134 , \40123 , \40133 );
and \U$39758 ( \40135 , \40097 , \40122 );
or \U$39759 ( \40136 , \40134 , \40135 );
and \U$39760 ( \40137 , \40086 , \40136 );
and \U$39761 ( \40138 , \40083 , \40085 );
or \U$39762 ( \40139 , \40137 , \40138 );
not \U$39763 ( \40140 , \39848 );
not \U$39764 ( \40141 , \40140 );
not \U$39765 ( \40142 , \39859 );
not \U$39766 ( \40143 , \39893 );
not \U$39767 ( \40144 , \40143 );
or \U$39768 ( \40145 , \40142 , \40144 );
or \U$39769 ( \40146 , \39859 , \40143 );
nand \U$39770 ( \40147 , \40145 , \40146 );
not \U$39771 ( \40148 , \40147 );
or \U$39772 ( \40149 , \40141 , \40148 );
or \U$39773 ( \40150 , \40147 , \40140 );
nand \U$39774 ( \40151 , \40149 , \40150 );
xor \U$39775 ( \40152 , \40139 , \40151 );
xor \U$39776 ( \40153 , \39993 , \40003 );
xor \U$39777 ( \40154 , \40153 , \40014 );
not \U$39778 ( \40155 , \15719 );
not \U$39779 ( \40156 , RIc225990_61);
not \U$39780 ( \40157 , \11394 );
or \U$39781 ( \40158 , \40156 , \40157 );
nand \U$39782 ( \40159 , \9072 , \10338 );
nand \U$39783 ( \40160 , \40158 , \40159 );
not \U$39784 ( \40161 , \40160 );
or \U$39785 ( \40162 , \40155 , \40161 );
nand \U$39786 ( \40163 , \40001 , \15729 );
nand \U$39787 ( \40164 , \40162 , \40163 );
not \U$39788 ( \40165 , \40164 );
not \U$39789 ( \40166 , \12665 );
and \U$39790 ( \40167 , RIc225a80_59, \9251 );
not \U$39791 ( \40168 , RIc225a80_59);
and \U$39792 ( \40169 , \40168 , \30878 );
or \U$39793 ( \40170 , \40167 , \40169 );
not \U$39794 ( \40171 , \40170 );
or \U$39795 ( \40172 , \40166 , \40171 );
nand \U$39796 ( \40173 , \39991 , \12670 );
nand \U$39797 ( \40174 , \40172 , \40173 );
not \U$39798 ( \40175 , \40174 );
or \U$39799 ( \40176 , \40165 , \40175 );
or \U$39800 ( \40177 , \40164 , \40174 );
and \U$39801 ( \40178 , \39888 , \13024 );
not \U$39802 ( \40179 , RIc225c60_55);
not \U$39803 ( \40180 , \31894 );
or \U$39804 ( \40181 , \40179 , \40180 );
not \U$39805 ( \40182 , \10360 );
nand \U$39806 ( \40183 , \40182 , \11041 );
nand \U$39807 ( \40184 , \40181 , \40183 );
and \U$39808 ( \40185 , \40184 , \11117 );
nor \U$39809 ( \40186 , \40178 , \40185 );
not \U$39810 ( \40187 , \40186 );
nand \U$39811 ( \40188 , \40177 , \40187 );
nand \U$39812 ( \40189 , \40176 , \40188 );
or \U$39813 ( \40190 , \40154 , \40189 );
not \U$39814 ( \40191 , \40190 );
xor \U$39815 ( \40192 , \40058 , \40067 );
xor \U$39816 ( \40193 , \40192 , \40080 );
or \U$39817 ( \40194 , RIc225eb8_50, RIc225e40_51);
nand \U$39818 ( \40195 , \40194 , \18367 );
and \U$39819 ( \40196 , RIc225eb8_50, RIc225e40_51);
nor \U$39820 ( \40197 , \40196 , \9541 );
and \U$39821 ( \40198 , \40195 , \40197 );
not \U$39822 ( \40199 , \9552 );
not \U$39823 ( \40200 , \40104 );
or \U$39824 ( \40201 , \40199 , \40200 );
or \U$39825 ( \40202 , \18357 , \9541 );
or \U$39826 ( \40203 , \18356 , RIc225f30_49);
nand \U$39827 ( \40204 , \40202 , \40203 );
nand \U$39828 ( \40205 , \40204 , \9532 );
nand \U$39829 ( \40206 , \40201 , \40205 );
and \U$39830 ( \40207 , \40198 , \40206 );
not \U$39831 ( \40208 , \8777 );
not \U$39832 ( \40209 , RIc225d50_53);
not \U$39833 ( \40210 , \20690 );
or \U$39834 ( \40211 , \40209 , \40210 );
nand \U$39835 ( \40212 , \20694 , \11585 );
nand \U$39836 ( \40213 , \40211 , \40212 );
not \U$39837 ( \40214 , \40213 );
or \U$39838 ( \40215 , \40208 , \40214 );
nand \U$39839 ( \40216 , \40076 , \8788 );
nand \U$39840 ( \40217 , \40215 , \40216 );
xor \U$39841 ( \40218 , \40207 , \40217 );
not \U$39842 ( \40219 , \12532 );
not \U$39843 ( \40220 , \40184 );
or \U$39844 ( \40221 , \40219 , \40220 );
and \U$39845 ( \40222 , RIc225c60_55, \10199 );
not \U$39846 ( \40223 , RIc225c60_55);
and \U$39847 ( \40224 , \40223 , \35896 );
or \U$39848 ( \40225 , \40222 , \40224 );
nand \U$39849 ( \40226 , \40225 , \11117 );
nand \U$39850 ( \40227 , \40221 , \40226 );
and \U$39851 ( \40228 , \40218 , \40227 );
and \U$39852 ( \40229 , \40207 , \40217 );
or \U$39853 ( \40230 , \40228 , \40229 );
xor \U$39854 ( \40231 , \40193 , \40230 );
not \U$39855 ( \40232 , RIc225828_64);
not \U$39856 ( \40233 , \40010 );
or \U$39857 ( \40234 , \40232 , \40233 );
and \U$39858 ( \40235 , \8925 , RIc2258a0_63);
not \U$39859 ( \40236 , \8925 );
and \U$39860 ( \40237 , \40236 , \15620 );
or \U$39861 ( \40238 , \40235 , \40237 );
nand \U$39862 ( \40239 , \40238 , \20159 );
nand \U$39863 ( \40240 , \40234 , \40239 );
and \U$39864 ( \40241 , \40231 , \40240 );
and \U$39865 ( \40242 , \40193 , \40230 );
or \U$39866 ( \40243 , \40241 , \40242 );
not \U$39867 ( \40244 , \40243 );
or \U$39868 ( \40245 , \40191 , \40244 );
nand \U$39869 ( \40246 , \40154 , \40189 );
nand \U$39870 ( \40247 , \40245 , \40246 );
and \U$39871 ( \40248 , \40152 , \40247 );
and \U$39872 ( \40249 , \40139 , \40151 );
or \U$39873 ( \40250 , \40248 , \40249 );
and \U$39874 ( \40251 , \40057 , \40250 );
and \U$39875 ( \40252 , \40054 , \40056 );
or \U$39876 ( \40253 , \40251 , \40252 );
nand \U$39877 ( \40254 , \40049 , \40253 );
xor \U$39878 ( \40255 , \40054 , \40056 );
xor \U$39879 ( \40256 , \40255 , \40250 );
xor \U$39880 ( \40257 , \39932 , \39983 );
xor \U$39881 ( \40258 , \40257 , \40017 );
not \U$39882 ( \40259 , \40258 );
xor \U$39883 ( \40260 , \39864 , \39874 );
xor \U$39884 ( \40261 , \40260 , \39890 );
not \U$39885 ( \40262 , \40261 );
xor \U$39886 ( \40263 , \40083 , \40085 );
xor \U$39887 ( \40264 , \40263 , \40136 );
not \U$39888 ( \40265 , \40264 );
or \U$39889 ( \40266 , \40262 , \40265 );
or \U$39890 ( \40267 , \40264 , \40261 );
xor \U$39891 ( \40268 , \40097 , \40122 );
xor \U$39892 ( \40269 , \40268 , \40133 );
xor \U$39893 ( \40270 , \40198 , \40206 );
not \U$39894 ( \40271 , \9444 );
not \U$39895 ( \40272 , \40115 );
or \U$39896 ( \40273 , \40271 , \40272 );
and \U$39897 ( \40274 , \22140 , \17613 );
not \U$39898 ( \40275 , \22140 );
and \U$39899 ( \40276 , \40275 , \21097 );
nor \U$39900 ( \40277 , \40274 , \40276 );
nand \U$39901 ( \40278 , \40277 , \9458 );
nand \U$39902 ( \40279 , \40273 , \40278 );
xor \U$39903 ( \40280 , \40270 , \40279 );
not \U$39904 ( \40281 , \8788 );
not \U$39905 ( \40282 , \40213 );
or \U$39906 ( \40283 , \40281 , \40282 );
not \U$39907 ( \40284 , RIc225d50_53);
not \U$39908 ( \40285 , \20519 );
or \U$39909 ( \40286 , \40284 , \40285 );
not \U$39910 ( \40287 , \20519 );
nand \U$39911 ( \40288 , \40287 , \11391 );
nand \U$39912 ( \40289 , \40286 , \40288 );
nand \U$39913 ( \40290 , \40289 , \8777 );
nand \U$39914 ( \40291 , \40283 , \40290 );
and \U$39915 ( \40292 , \40280 , \40291 );
and \U$39916 ( \40293 , \40270 , \40279 );
or \U$39917 ( \40294 , \40292 , \40293 );
not \U$39918 ( \40295 , \12670 );
not \U$39919 ( \40296 , \40170 );
or \U$39920 ( \40297 , \40295 , \40296 );
and \U$39921 ( \40298 , RIc225a80_59, \10975 );
not \U$39922 ( \40299 , RIc225a80_59);
and \U$39923 ( \40300 , \40299 , \9274 );
or \U$39924 ( \40301 , \40298 , \40300 );
nand \U$39925 ( \40302 , \40301 , \12665 );
nand \U$39926 ( \40303 , \40297 , \40302 );
xor \U$39927 ( \40304 , \40294 , \40303 );
not \U$39928 ( \40305 , \15729 );
not \U$39929 ( \40306 , \40160 );
or \U$39930 ( \40307 , \40305 , \40306 );
and \U$39931 ( \40308 , \10111 , RIc225990_61);
not \U$39932 ( \40309 , \10111 );
and \U$39933 ( \40310 , \40309 , \12806 );
or \U$39934 ( \40311 , \40308 , \40310 );
nand \U$39935 ( \40312 , \40311 , \15719 );
nand \U$39936 ( \40313 , \40307 , \40312 );
and \U$39937 ( \40314 , \40304 , \40313 );
and \U$39938 ( \40315 , \40294 , \40303 );
or \U$39939 ( \40316 , \40314 , \40315 );
xor \U$39940 ( \40317 , \40269 , \40316 );
xor \U$39941 ( \40318 , \40098 , \40108 );
xor \U$39942 ( \40319 , \40318 , \40119 );
not \U$39943 ( \40320 , \15267 );
not \U$39944 ( \40321 , \40131 );
or \U$39945 ( \40322 , \40320 , \40321 );
not \U$39946 ( \40323 , RIc225b70_57);
not \U$39947 ( \40324 , \9321 );
or \U$39948 ( \40325 , \40323 , \40324 );
nand \U$39949 ( \40326 , \9320 , \15262 );
nand \U$39950 ( \40327 , \40325 , \40326 );
nand \U$39951 ( \40328 , \40327 , \11965 );
nand \U$39952 ( \40329 , \40322 , \40328 );
xor \U$39953 ( \40330 , \40319 , \40329 );
not \U$39954 ( \40331 , RIc225828_64);
not \U$39955 ( \40332 , \40238 );
or \U$39956 ( \40333 , \40331 , \40332 );
not \U$39957 ( \40334 , RIc2258a0_63);
not \U$39958 ( \40335 , \38643 );
or \U$39959 ( \40336 , \40334 , \40335 );
nand \U$39960 ( \40337 , \14608 , \37494 );
nand \U$39961 ( \40338 , \40336 , \40337 );
nand \U$39962 ( \40339 , \40338 , \16891 );
nand \U$39963 ( \40340 , \40333 , \40339 );
and \U$39964 ( \40341 , \40330 , \40340 );
and \U$39965 ( \40342 , \40319 , \40329 );
or \U$39966 ( \40343 , \40341 , \40342 );
and \U$39967 ( \40344 , \40317 , \40343 );
and \U$39968 ( \40345 , \40269 , \40316 );
or \U$39969 ( \40346 , \40344 , \40345 );
nand \U$39970 ( \40347 , \40267 , \40346 );
nand \U$39971 ( \40348 , \40266 , \40347 );
not \U$39972 ( \40349 , \40348 );
nand \U$39973 ( \40350 , \40259 , \40349 );
not \U$39974 ( \40351 , \40350 );
xor \U$39975 ( \40352 , \40139 , \40151 );
xor \U$39976 ( \40353 , \40352 , \40247 );
not \U$39977 ( \40354 , \40353 );
or \U$39978 ( \40355 , \40351 , \40354 );
nand \U$39979 ( \40356 , \40258 , \40348 );
nand \U$39980 ( \40357 , \40355 , \40356 );
nand \U$39981 ( \40358 , \40256 , \40357 );
nand \U$39982 ( \40359 , \40254 , \40358 );
or \U$39983 ( \40360 , \40049 , \40253 );
nand \U$39984 ( \40361 , \40359 , \40360 );
xor \U$39985 ( \40362 , \39694 , \39757 );
xnor \U$39986 ( \40363 , \40362 , \39755 );
not \U$39987 ( \40364 , \40363 );
not \U$39988 ( \40365 , \39611 );
not \U$39989 ( \40366 , \39615 );
or \U$39990 ( \40367 , \40365 , \40366 );
or \U$39991 ( \40368 , \39615 , \39611 );
nand \U$39992 ( \40369 , \40367 , \40368 );
xnor \U$39993 ( \40370 , \40369 , \39683 );
not \U$39994 ( \40371 , \40370 );
xor \U$39995 ( \40372 , \40028 , \40030 );
and \U$39996 ( \40373 , \40372 , \40047 );
and \U$39997 ( \40374 , \40028 , \40030 );
or \U$39998 ( \40375 , \40373 , \40374 );
not \U$39999 ( \40376 , \40375 );
or \U$40000 ( \40377 , \40371 , \40376 );
or \U$40001 ( \40378 , \40375 , \40370 );
nand \U$40002 ( \40379 , \40377 , \40378 );
not \U$40003 ( \40380 , \40379 );
or \U$40004 ( \40381 , \40364 , \40380 );
or \U$40005 ( \40382 , \40363 , \40379 );
nand \U$40006 ( \40383 , \40381 , \40382 );
xor \U$40007 ( \40384 , \39802 , \40023 );
and \U$40008 ( \40385 , \40384 , \40048 );
and \U$40009 ( \40386 , \39802 , \40023 );
or \U$40010 ( \40387 , \40385 , \40386 );
nor \U$40011 ( \40388 , \40383 , \40387 );
or \U$40012 ( \40389 , \40361 , \40388 );
nand \U$40013 ( \40390 , \40383 , \40387 );
nand \U$40014 ( \40391 , \40389 , \40390 );
not \U$40015 ( \40392 , \39768 );
not \U$40016 ( \40393 , \39759 );
or \U$40017 ( \40394 , \40392 , \40393 );
or \U$40018 ( \40395 , \39759 , \39768 );
nand \U$40019 ( \40396 , \40394 , \40395 );
xnor \U$40020 ( \40397 , \40396 , \39776 );
nand \U$40021 ( \40398 , \40363 , \40370 );
and \U$40022 ( \40399 , \40398 , \40375 );
nor \U$40023 ( \40400 , \40363 , \40370 );
nor \U$40024 ( \40401 , \40399 , \40400 );
nand \U$40025 ( \40402 , \40397 , \40401 );
and \U$40026 ( \40403 , \40391 , \40402 );
nor \U$40027 ( \40404 , \40397 , \40401 );
nor \U$40028 ( \40405 , \40403 , \40404 );
nor \U$40029 ( \40406 , \39800 , \40405 );
nor \U$40030 ( \40407 , \39797 , \40406 );
not \U$40031 ( \40408 , \40407 );
not \U$40032 ( \40409 , \39800 );
xor \U$40033 ( \40410 , \40269 , \40316 );
xor \U$40034 ( \40411 , \40410 , \40343 );
xor \U$40035 ( \40412 , \40294 , \40303 );
xor \U$40036 ( \40413 , \40412 , \40313 );
xor \U$40037 ( \40414 , \40319 , \40329 );
xor \U$40038 ( \40415 , \40414 , \40340 );
xor \U$40039 ( \40416 , \40413 , \40415 );
xor \U$40040 ( \40417 , \40270 , \40279 );
xor \U$40041 ( \40418 , \40417 , \40291 );
or \U$40042 ( \40419 , RIc225dc8_52, RIc225d50_53);
nand \U$40043 ( \40420 , \40419 , \18182 );
and \U$40044 ( \40421 , RIc225dc8_52, RIc225d50_53);
nor \U$40045 ( \40422 , \40421 , \11795 );
and \U$40046 ( \40423 , \40420 , \40422 );
not \U$40047 ( \40424 , \9444 );
and \U$40048 ( \40425 , RIc225e40_51, \32588 );
not \U$40049 ( \40426 , RIc225e40_51);
and \U$40050 ( \40427 , \40426 , \16259 );
nor \U$40051 ( \40428 , \40425 , \40427 );
not \U$40052 ( \40429 , \40428 );
or \U$40053 ( \40430 , \40424 , \40429 );
or \U$40054 ( \40431 , \18367 , \11795 );
or \U$40055 ( \40432 , \18356 , RIc225e40_51);
nand \U$40056 ( \40433 , \40431 , \40432 );
nand \U$40057 ( \40434 , \40433 , \9457 );
nand \U$40058 ( \40435 , \40430 , \40434 );
and \U$40059 ( \40436 , \40423 , \40435 );
not \U$40060 ( \40437 , \11038 );
not \U$40061 ( \40438 , RIc225c60_55);
not \U$40062 ( \40439 , \21084 );
or \U$40063 ( \40440 , \40438 , \40439 );
buf \U$40064 ( \40441 , \37397 );
nand \U$40065 ( \40442 , \40441 , \11108 );
nand \U$40066 ( \40443 , \40440 , \40442 );
not \U$40067 ( \40444 , \40443 );
or \U$40068 ( \40445 , \40437 , \40444 );
not \U$40069 ( \40446 , RIc225c60_55);
not \U$40070 ( \40447 , \20690 );
or \U$40071 ( \40448 , \40446 , \40447 );
nand \U$40072 ( \40449 , \12756 , \8767 );
nand \U$40073 ( \40450 , \40448 , \40449 );
nand \U$40074 ( \40451 , \40450 , \11117 );
nand \U$40075 ( \40452 , \40445 , \40451 );
xor \U$40076 ( \40453 , \40436 , \40452 );
not \U$40077 ( \40454 , \15267 );
buf \U$40078 ( \40455 , \10086 );
and \U$40079 ( \40456 , RIc225b70_57, \40455 );
not \U$40080 ( \40457 , RIc225b70_57);
not \U$40081 ( \40458 , \40455 );
and \U$40082 ( \40459 , \40457 , \40458 );
nor \U$40083 ( \40460 , \40456 , \40459 );
not \U$40084 ( \40461 , \40460 );
or \U$40085 ( \40462 , \40454 , \40461 );
and \U$40086 ( \40463 , \11033 , \10199 );
not \U$40087 ( \40464 , \11033 );
and \U$40088 ( \40465 , \40464 , \35896 );
nor \U$40089 ( \40466 , \40463 , \40465 );
nand \U$40090 ( \40467 , \40466 , \11965 );
nand \U$40091 ( \40468 , \40462 , \40467 );
and \U$40092 ( \40469 , \40453 , \40468 );
and \U$40093 ( \40470 , \40436 , \40452 );
or \U$40094 ( \40471 , \40469 , \40470 );
xor \U$40095 ( \40472 , \40418 , \40471 );
and \U$40096 ( \40473 , \18367 , \9552 );
not \U$40097 ( \40474 , \9458 );
not \U$40098 ( \40475 , \40428 );
or \U$40099 ( \40476 , \40474 , \40475 );
nand \U$40100 ( \40477 , \40277 , \9444 );
nand \U$40101 ( \40478 , \40476 , \40477 );
xor \U$40102 ( \40479 , \40473 , \40478 );
not \U$40103 ( \40480 , \8777 );
not \U$40104 ( \40481 , RIc225d50_53);
not \U$40105 ( \40482 , \12846 );
or \U$40106 ( \40483 , \40481 , \40482 );
nand \U$40107 ( \40484 , \18161 , \8772 );
nand \U$40108 ( \40485 , \40483 , \40484 );
not \U$40109 ( \40486 , \40485 );
or \U$40110 ( \40487 , \40480 , \40486 );
nand \U$40111 ( \40488 , \40289 , \8788 );
nand \U$40112 ( \40489 , \40487 , \40488 );
xor \U$40113 ( \40490 , \40479 , \40489 );
not \U$40114 ( \40491 , \12670 );
xnor \U$40115 ( \40492 , RIc225a80_59, \30069 );
not \U$40116 ( \40493 , \40492 );
or \U$40117 ( \40494 , \40491 , \40493 );
and \U$40118 ( \40495 , RIc225a80_59, \12100 );
not \U$40119 ( \40496 , RIc225a80_59);
and \U$40120 ( \40497 , \40496 , \9320 );
or \U$40121 ( \40498 , \40495 , \40497 );
nand \U$40122 ( \40499 , \40498 , \15164 );
nand \U$40123 ( \40500 , \40494 , \40499 );
xor \U$40124 ( \40501 , \40490 , \40500 );
not \U$40125 ( \40502 , \20862 );
not \U$40126 ( \40503 , RIc225990_61);
not \U$40127 ( \40504 , \9251 );
or \U$40128 ( \40505 , \40503 , \40504 );
nand \U$40129 ( \40506 , \35479 , \12806 );
nand \U$40130 ( \40507 , \40505 , \40506 );
not \U$40131 ( \40508 , \40507 );
or \U$40132 ( \40509 , \40502 , \40508 );
not \U$40133 ( \40510 , RIc225990_61);
not \U$40134 ( \40511 , \10975 );
or \U$40135 ( \40512 , \40510 , \40511 );
nand \U$40136 ( \40513 , \9274 , \10338 );
nand \U$40137 ( \40514 , \40512 , \40513 );
nand \U$40138 ( \40515 , \40514 , \15719 );
nand \U$40139 ( \40516 , \40509 , \40515 );
and \U$40140 ( \40517 , \40501 , \40516 );
and \U$40141 ( \40518 , \40490 , \40500 );
or \U$40142 ( \40519 , \40517 , \40518 );
and \U$40143 ( \40520 , \40472 , \40519 );
and \U$40144 ( \40521 , \40418 , \40471 );
or \U$40145 ( \40522 , \40520 , \40521 );
and \U$40146 ( \40523 , \40416 , \40522 );
and \U$40147 ( \40524 , \40413 , \40415 );
or \U$40148 ( \40525 , \40523 , \40524 );
not \U$40149 ( \40526 , \40525 );
xor \U$40150 ( \40527 , \40411 , \40526 );
xnor \U$40151 ( \40528 , \40186 , \40174 );
xor \U$40152 ( \40529 , \40528 , \40164 );
xor \U$40153 ( \40530 , \40193 , \40230 );
xor \U$40154 ( \40531 , \40530 , \40240 );
xor \U$40155 ( \40532 , \40529 , \40531 );
xor \U$40156 ( \40533 , \40207 , \40217 );
xor \U$40157 ( \40534 , \40533 , \40227 );
not \U$40158 ( \40535 , \11117 );
not \U$40159 ( \40536 , \40443 );
or \U$40160 ( \40537 , \40535 , \40536 );
nand \U$40161 ( \40538 , \40225 , \13024 );
nand \U$40162 ( \40539 , \40537 , \40538 );
xor \U$40163 ( \40540 , \40473 , \40478 );
and \U$40164 ( \40541 , \40540 , \40489 );
and \U$40165 ( \40542 , \40473 , \40478 );
or \U$40166 ( \40543 , \40541 , \40542 );
xor \U$40167 ( \40544 , \40539 , \40543 );
not \U$40168 ( \40545 , \40327 );
not \U$40169 ( \40546 , \11974 );
or \U$40170 ( \40547 , \40545 , \40546 );
nand \U$40171 ( \40548 , \40460 , \11965 );
nand \U$40172 ( \40549 , \40547 , \40548 );
and \U$40173 ( \40550 , \40544 , \40549 );
and \U$40174 ( \40551 , \40539 , \40543 );
or \U$40175 ( \40552 , \40550 , \40551 );
xor \U$40176 ( \40553 , \40534 , \40552 );
not \U$40177 ( \40554 , \15729 );
not \U$40178 ( \40555 , \40311 );
or \U$40179 ( \40556 , \40554 , \40555 );
nand \U$40180 ( \40557 , \40507 , \15719 );
nand \U$40181 ( \40558 , \40556 , \40557 );
not \U$40182 ( \40559 , \40558 );
not \U$40183 ( \40560 , RIc225828_64);
not \U$40184 ( \40561 , \40338 );
or \U$40185 ( \40562 , \40560 , \40561 );
not \U$40186 ( \40563 , RIc2258a0_63);
not \U$40187 ( \40564 , \9073 );
or \U$40188 ( \40565 , \40563 , \40564 );
nand \U$40189 ( \40566 , \9072 , \16880 );
nand \U$40190 ( \40567 , \40565 , \40566 );
nand \U$40191 ( \40568 , \40567 , \16891 );
nand \U$40192 ( \40569 , \40562 , \40568 );
not \U$40193 ( \40570 , \40569 );
or \U$40194 ( \40571 , \40559 , \40570 );
or \U$40195 ( \40572 , \40569 , \40558 );
not \U$40196 ( \40573 , \12670 );
not \U$40197 ( \40574 , \40301 );
or \U$40198 ( \40575 , \40573 , \40574 );
nand \U$40199 ( \40576 , \40492 , \15164 );
nand \U$40200 ( \40577 , \40575 , \40576 );
nand \U$40201 ( \40578 , \40572 , \40577 );
nand \U$40202 ( \40579 , \40571 , \40578 );
and \U$40203 ( \40580 , \40553 , \40579 );
and \U$40204 ( \40581 , \40534 , \40552 );
or \U$40205 ( \40582 , \40580 , \40581 );
xor \U$40206 ( \40583 , \40532 , \40582 );
xnor \U$40207 ( \40584 , \40527 , \40583 );
xor \U$40208 ( \40585 , \40534 , \40552 );
xor \U$40209 ( \40586 , \40585 , \40579 );
xor \U$40210 ( \40587 , \40539 , \40543 );
xor \U$40211 ( \40588 , \40587 , \40549 );
not \U$40212 ( \40589 , \40588 );
xor \U$40213 ( \40590 , \40569 , \40558 );
xnor \U$40214 ( \40591 , \40590 , \40577 );
not \U$40215 ( \40592 , \40591 );
not \U$40216 ( \40593 , \40592 );
or \U$40217 ( \40594 , \40589 , \40593 );
or \U$40218 ( \40595 , \40592 , \40588 );
xor \U$40219 ( \40596 , \40423 , \40435 );
not \U$40220 ( \40597 , \8788 );
not \U$40221 ( \40598 , \40485 );
or \U$40222 ( \40599 , \40597 , \40598 );
and \U$40223 ( \40600 , RIc225d50_53, \20393 );
not \U$40224 ( \40601 , RIc225d50_53);
and \U$40225 ( \40602 , \40601 , \30679 );
nor \U$40226 ( \40603 , \40600 , \40602 );
nand \U$40227 ( \40604 , \40603 , \8777 );
nand \U$40228 ( \40605 , \40599 , \40604 );
xor \U$40229 ( \40606 , \40596 , \40605 );
not \U$40230 ( \40607 , \11038 );
not \U$40231 ( \40608 , \40450 );
or \U$40232 ( \40609 , \40607 , \40608 );
and \U$40233 ( \40610 , RIc225c60_55, \40287 );
not \U$40234 ( \40611 , RIc225c60_55);
and \U$40235 ( \40612 , \40611 , \15444 );
nor \U$40236 ( \40613 , \40610 , \40612 );
nand \U$40237 ( \40614 , \40613 , \11045 );
nand \U$40238 ( \40615 , \40609 , \40614 );
and \U$40239 ( \40616 , \40606 , \40615 );
and \U$40240 ( \40617 , \40596 , \40605 );
or \U$40241 ( \40618 , \40616 , \40617 );
not \U$40242 ( \40619 , RIc225828_64);
not \U$40243 ( \40620 , \40567 );
or \U$40244 ( \40621 , \40619 , \40620 );
not \U$40245 ( \40622 , RIc2258a0_63);
not \U$40246 ( \40623 , \10111 );
or \U$40247 ( \40624 , \40622 , \40623 );
nand \U$40248 ( \40625 , \10110 , \16880 );
nand \U$40249 ( \40626 , \40624 , \40625 );
nand \U$40250 ( \40627 , \40626 , \16891 );
nand \U$40251 ( \40628 , \40621 , \40627 );
xor \U$40252 ( \40629 , \40618 , \40628 );
xor \U$40253 ( \40630 , \40436 , \40452 );
xor \U$40254 ( \40631 , \40630 , \40468 );
and \U$40255 ( \40632 , \40629 , \40631 );
and \U$40256 ( \40633 , \40618 , \40628 );
or \U$40257 ( \40634 , \40632 , \40633 );
nand \U$40258 ( \40635 , \40595 , \40634 );
nand \U$40259 ( \40636 , \40594 , \40635 );
xor \U$40260 ( \40637 , \40586 , \40636 );
xor \U$40261 ( \40638 , \40413 , \40415 );
xor \U$40262 ( \40639 , \40638 , \40522 );
and \U$40263 ( \40640 , \40637 , \40639 );
and \U$40264 ( \40641 , \40586 , \40636 );
or \U$40265 ( \40642 , \40640 , \40641 );
or \U$40266 ( \40643 , \40584 , \40642 );
nand \U$40267 ( \40644 , \40584 , \40642 );
xor \U$40268 ( \40645 , \40586 , \40636 );
xor \U$40269 ( \40646 , \40645 , \40639 );
xor \U$40270 ( \40647 , \40418 , \40471 );
xor \U$40271 ( \40648 , \40647 , \40519 );
not \U$40272 ( \40649 , \40648 );
not \U$40273 ( \40650 , \40649 );
xor \U$40274 ( \40651 , \40588 , \40591 );
xor \U$40275 ( \40652 , \40651 , \40634 );
not \U$40276 ( \40653 , \40652 );
or \U$40277 ( \40654 , \40650 , \40653 );
not \U$40278 ( \40655 , \11965 );
not \U$40279 ( \40656 , RIc225b70_57);
not \U$40280 ( \40657 , \40441 );
not \U$40281 ( \40658 , \40657 );
or \U$40282 ( \40659 , \40656 , \40658 );
nand \U$40283 ( \40660 , \40074 , \12475 );
nand \U$40284 ( \40661 , \40659 , \40660 );
not \U$40285 ( \40662 , \40661 );
or \U$40286 ( \40663 , \40655 , \40662 );
nand \U$40287 ( \40664 , \40466 , \11974 );
nand \U$40288 ( \40665 , \40663 , \40664 );
and \U$40289 ( \40666 , \18357 , \9444 );
not \U$40290 ( \40667 , \8788 );
not \U$40291 ( \40668 , \40603 );
or \U$40292 ( \40669 , \40667 , \40668 );
and \U$40293 ( \40670 , RIc225d50_53, \16256 );
not \U$40294 ( \40671 , RIc225d50_53);
and \U$40295 ( \40672 , \40671 , \32587 );
nor \U$40296 ( \40673 , \40670 , \40672 );
nand \U$40297 ( \40674 , \40673 , \8777 );
nand \U$40298 ( \40675 , \40669 , \40674 );
xor \U$40299 ( \40676 , \40666 , \40675 );
not \U$40300 ( \40677 , \11045 );
not \U$40301 ( \40678 , RIc225c60_55);
not \U$40302 ( \40679 , \12846 );
or \U$40303 ( \40680 , \40678 , \40679 );
nand \U$40304 ( \40681 , \18161 , \11041 );
nand \U$40305 ( \40682 , \40680 , \40681 );
not \U$40306 ( \40683 , \40682 );
or \U$40307 ( \40684 , \40677 , \40683 );
nand \U$40308 ( \40685 , \40613 , \11038 );
nand \U$40309 ( \40686 , \40684 , \40685 );
and \U$40310 ( \40687 , \40676 , \40686 );
and \U$40311 ( \40688 , \40666 , \40675 );
or \U$40312 ( \40689 , \40687 , \40688 );
xor \U$40313 ( \40690 , \40665 , \40689 );
not \U$40314 ( \40691 , \15719 );
not \U$40315 ( \40692 , RIc225990_61);
not \U$40316 ( \40693 , \30069 );
or \U$40317 ( \40694 , \40692 , \40693 );
nand \U$40318 ( \40695 , \9299 , \10338 );
nand \U$40319 ( \40696 , \40694 , \40695 );
not \U$40320 ( \40697 , \40696 );
or \U$40321 ( \40698 , \40691 , \40697 );
nand \U$40322 ( \40699 , \15729 , \40514 );
nand \U$40323 ( \40700 , \40698 , \40699 );
and \U$40324 ( \40701 , \40690 , \40700 );
and \U$40325 ( \40702 , \40665 , \40689 );
or \U$40326 ( \40703 , \40701 , \40702 );
xor \U$40327 ( \40704 , \40490 , \40500 );
xor \U$40328 ( \40705 , \40704 , \40516 );
xor \U$40329 ( \40706 , \40703 , \40705 );
xor \U$40330 ( \40707 , \40596 , \40605 );
xor \U$40331 ( \40708 , \40707 , \40615 );
not \U$40332 ( \40709 , \12670 );
not \U$40333 ( \40710 , \40498 );
or \U$40334 ( \40711 , \40709 , \40710 );
and \U$40335 ( \40712 , RIc225a80_59, \40455 );
not \U$40336 ( \40713 , RIc225a80_59);
and \U$40337 ( \40714 , \40713 , \31894 );
nor \U$40338 ( \40715 , \40712 , \40714 );
nand \U$40339 ( \40716 , \40715 , \15164 );
nand \U$40340 ( \40717 , \40711 , \40716 );
xor \U$40341 ( \40718 , \40708 , \40717 );
not \U$40342 ( \40719 , \16891 );
not \U$40343 ( \40720 , RIc2258a0_63);
not \U$40344 ( \40721 , \11488 );
or \U$40345 ( \40722 , \40720 , \40721 );
nand \U$40346 ( \40723 , \30878 , \16880 );
nand \U$40347 ( \40724 , \40722 , \40723 );
not \U$40348 ( \40725 , \40724 );
or \U$40349 ( \40726 , \40719 , \40725 );
nand \U$40350 ( \40727 , \40626 , RIc225828_64);
nand \U$40351 ( \40728 , \40726 , \40727 );
and \U$40352 ( \40729 , \40718 , \40728 );
and \U$40353 ( \40730 , \40708 , \40717 );
or \U$40354 ( \40731 , \40729 , \40730 );
and \U$40355 ( \40732 , \40706 , \40731 );
and \U$40356 ( \40733 , \40703 , \40705 );
or \U$40357 ( \40734 , \40732 , \40733 );
nand \U$40358 ( \40735 , \40654 , \40734 );
not \U$40359 ( \40736 , \40652 );
nand \U$40360 ( \40737 , \40736 , \40648 );
nand \U$40361 ( \40738 , \40735 , \40737 );
nand \U$40362 ( \40739 , \40646 , \40738 );
nand \U$40363 ( \40740 , \40644 , \40739 );
nand \U$40364 ( \40741 , \40643 , \40740 );
xor \U$40365 ( \40742 , \40189 , \40243 );
xnor \U$40366 ( \40743 , \40742 , \40154 );
xor \U$40367 ( \40744 , \40529 , \40531 );
and \U$40368 ( \40745 , \40744 , \40582 );
and \U$40369 ( \40746 , \40529 , \40531 );
or \U$40370 ( \40747 , \40745 , \40746 );
not \U$40371 ( \40748 , \40747 );
xor \U$40372 ( \40749 , \40743 , \40748 );
xor \U$40373 ( \40750 , \40261 , \40264 );
xnor \U$40374 ( \40751 , \40750 , \40346 );
xor \U$40375 ( \40752 , \40749 , \40751 );
not \U$40376 ( \40753 , \40411 );
nand \U$40377 ( \40754 , \40753 , \40526 );
and \U$40378 ( \40755 , \40583 , \40754 );
nor \U$40379 ( \40756 , \40526 , \40753 );
nor \U$40380 ( \40757 , \40755 , \40756 );
nand \U$40381 ( \40758 , \40752 , \40757 );
not \U$40382 ( \40759 , \40758 );
nor \U$40383 ( \40760 , \40741 , \40759 );
nor \U$40384 ( \40761 , \40752 , \40757 );
or \U$40385 ( \40762 , \40760 , \40761 );
not \U$40386 ( \40763 , \40349 );
not \U$40387 ( \40764 , \40258 );
or \U$40388 ( \40765 , \40763 , \40764 );
nand \U$40389 ( \40766 , \40259 , \40348 );
nand \U$40390 ( \40767 , \40765 , \40766 );
xnor \U$40391 ( \40768 , \40767 , \40353 );
xor \U$40392 ( \40769 , \40743 , \40748 );
and \U$40393 ( \40770 , \40769 , \40751 );
and \U$40394 ( \40771 , \40743 , \40748 );
or \U$40395 ( \40772 , \40770 , \40771 );
nand \U$40396 ( \40773 , \40768 , \40772 );
nand \U$40397 ( \40774 , \40762 , \40773 );
or \U$40398 ( \40775 , \40646 , \40738 );
and \U$40399 ( \40776 , \40775 , \40643 );
xor \U$40400 ( \40777 , \40618 , \40628 );
xor \U$40401 ( \40778 , \40777 , \40631 );
not \U$40402 ( \40779 , \40778 );
or \U$40403 ( \40780 , RIc225cd8_54, RIc225c60_55);
nand \U$40404 ( \40781 , \40780 , \18367 );
and \U$40405 ( \40782 , RIc225cd8_54, RIc225c60_55);
nor \U$40406 ( \40783 , \40782 , \8782 );
and \U$40407 ( \40784 , \40781 , \40783 );
not \U$40408 ( \40785 , \40673 );
not \U$40409 ( \40786 , \8788 );
or \U$40410 ( \40787 , \40785 , \40786 );
and \U$40411 ( \40788 , \18356 , RIc225d50_53);
and \U$40412 ( \40789 , \18357 , \8782 );
nor \U$40413 ( \40790 , \40788 , \40789 );
or \U$40414 ( \40791 , \40790 , \8776 );
nand \U$40415 ( \40792 , \40787 , \40791 );
and \U$40416 ( \40793 , \40784 , \40792 );
not \U$40417 ( \40794 , \11974 );
not \U$40418 ( \40795 , \40661 );
or \U$40419 ( \40796 , \40794 , \40795 );
not \U$40420 ( \40797 , RIc225b70_57);
not \U$40421 ( \40798 , \20690 );
or \U$40422 ( \40799 , \40797 , \40798 );
nand \U$40423 ( \40800 , \12756 , \12475 );
nand \U$40424 ( \40801 , \40799 , \40800 );
nand \U$40425 ( \40802 , \40801 , \11965 );
nand \U$40426 ( \40803 , \40796 , \40802 );
xor \U$40427 ( \40804 , \40793 , \40803 );
not \U$40428 ( \40805 , \12670 );
not \U$40429 ( \40806 , \40715 );
or \U$40430 ( \40807 , \40805 , \40806 );
and \U$40431 ( \40808 , \17064 , \27990 );
not \U$40432 ( \40809 , \17064 );
not \U$40433 ( \40810 , \10199 );
and \U$40434 ( \40811 , \40809 , \40810 );
nor \U$40435 ( \40812 , \40808 , \40811 );
nand \U$40436 ( \40813 , \40812 , \15164 );
nand \U$40437 ( \40814 , \40807 , \40813 );
and \U$40438 ( \40815 , \40804 , \40814 );
and \U$40439 ( \40816 , \40793 , \40803 );
or \U$40440 ( \40817 , \40815 , \40816 );
xor \U$40441 ( \40818 , \40665 , \40689 );
xor \U$40442 ( \40819 , \40818 , \40700 );
xor \U$40443 ( \40820 , \40817 , \40819 );
not \U$40444 ( \40821 , \15719 );
and \U$40445 ( \40822 , \9321 , RIc225990_61);
not \U$40446 ( \40823 , \9321 );
and \U$40447 ( \40824 , \40823 , \12806 );
or \U$40448 ( \40825 , \40822 , \40824 );
not \U$40449 ( \40826 , \40825 );
or \U$40450 ( \40827 , \40821 , \40826 );
nand \U$40451 ( \40828 , \40696 , \15729 );
nand \U$40452 ( \40829 , \40827 , \40828 );
xor \U$40453 ( \40830 , \40666 , \40675 );
xor \U$40454 ( \40831 , \40830 , \40686 );
and \U$40455 ( \40832 , \40829 , \40831 );
not \U$40456 ( \40833 , RIc225828_64);
not \U$40457 ( \40834 , \40724 );
or \U$40458 ( \40835 , \40833 , \40834 );
not \U$40459 ( \40836 , RIc2258a0_63);
not \U$40460 ( \40837 , \10975 );
or \U$40461 ( \40838 , \40836 , \40837 );
nand \U$40462 ( \40839 , \9274 , \15620 );
nand \U$40463 ( \40840 , \40838 , \40839 );
nand \U$40464 ( \40841 , \40840 , \16891 );
nand \U$40465 ( \40842 , \40835 , \40841 );
xor \U$40466 ( \40843 , \40666 , \40675 );
xor \U$40467 ( \40844 , \40843 , \40686 );
and \U$40468 ( \40845 , \40842 , \40844 );
and \U$40469 ( \40846 , \40829 , \40842 );
or \U$40470 ( \40847 , \40832 , \40845 , \40846 );
and \U$40471 ( \40848 , \40820 , \40847 );
and \U$40472 ( \40849 , \40817 , \40819 );
or \U$40473 ( \40850 , \40848 , \40849 );
not \U$40474 ( \40851 , \40850 );
or \U$40475 ( \40852 , \40779 , \40851 );
not \U$40476 ( \40853 , \40778 );
not \U$40477 ( \40854 , \40853 );
not \U$40478 ( \40855 , \40850 );
not \U$40479 ( \40856 , \40855 );
or \U$40480 ( \40857 , \40854 , \40856 );
xor \U$40481 ( \40858 , \40703 , \40705 );
xor \U$40482 ( \40859 , \40858 , \40731 );
nand \U$40483 ( \40860 , \40857 , \40859 );
nand \U$40484 ( \40861 , \40852 , \40860 );
not \U$40485 ( \40862 , \40861 );
and \U$40486 ( \40863 , \40734 , \40648 );
not \U$40487 ( \40864 , \40734 );
and \U$40488 ( \40865 , \40864 , \40649 );
nor \U$40489 ( \40866 , \40863 , \40865 );
and \U$40490 ( \40867 , \40866 , \40652 );
not \U$40491 ( \40868 , \40866 );
and \U$40492 ( \40869 , \40868 , \40736 );
nor \U$40493 ( \40870 , \40867 , \40869 );
nand \U$40494 ( \40871 , \40862 , \40870 );
and \U$40495 ( \40872 , \40850 , \40853 );
not \U$40496 ( \40873 , \40850 );
and \U$40497 ( \40874 , \40873 , \40778 );
or \U$40498 ( \40875 , \40872 , \40874 );
not \U$40499 ( \40876 , \40859 );
and \U$40500 ( \40877 , \40875 , \40876 );
not \U$40501 ( \40878 , \40875 );
and \U$40502 ( \40879 , \40878 , \40859 );
nor \U$40503 ( \40880 , \40877 , \40879 );
xor \U$40504 ( \40881 , \40817 , \40819 );
xor \U$40505 ( \40882 , \40881 , \40847 );
xor \U$40506 ( \40883 , \40784 , \40792 );
not \U$40507 ( \40884 , \11038 );
not \U$40508 ( \40885 , \40682 );
or \U$40509 ( \40886 , \40884 , \40885 );
and \U$40510 ( \40887 , \15623 , RIc225c60_55);
and \U$40511 ( \40888 , \21097 , \8767 );
nor \U$40512 ( \40889 , \40887 , \40888 );
or \U$40513 ( \40890 , \40889 , \11046 );
nand \U$40514 ( \40891 , \40886 , \40890 );
xor \U$40515 ( \40892 , \40883 , \40891 );
not \U$40516 ( \40893 , \11974 );
not \U$40517 ( \40894 , \40801 );
or \U$40518 ( \40895 , \40893 , \40894 );
and \U$40519 ( \40896 , \18167 , RIc225b70_57);
and \U$40520 ( \40897 , \40093 , \12475 );
nor \U$40521 ( \40898 , \40896 , \40897 );
not \U$40522 ( \40899 , \40898 );
nand \U$40523 ( \40900 , \40899 , \11965 );
nand \U$40524 ( \40901 , \40895 , \40900 );
and \U$40525 ( \40902 , \40892 , \40901 );
and \U$40526 ( \40903 , \40883 , \40891 );
or \U$40527 ( \40904 , \40902 , \40903 );
xor \U$40528 ( \40905 , \40793 , \40803 );
xor \U$40529 ( \40906 , \40905 , \40814 );
xor \U$40530 ( \40907 , \40904 , \40906 );
not \U$40531 ( \40908 , \12665 );
and \U$40532 ( \40909 , \17064 , \40657 );
not \U$40533 ( \40910 , \17064 );
and \U$40534 ( \40911 , \40910 , \40074 );
nor \U$40535 ( \40912 , \40909 , \40911 );
not \U$40536 ( \40913 , \40912 );
or \U$40537 ( \40914 , \40908 , \40913 );
nand \U$40538 ( \40915 , \40812 , \12670 );
nand \U$40539 ( \40916 , \40914 , \40915 );
not \U$40540 ( \40917 , \18367 );
nor \U$40541 ( \40918 , \40917 , \8787 );
and \U$40542 ( \40919 , RIc225c60_55, \32588 );
not \U$40543 ( \40920 , RIc225c60_55);
and \U$40544 ( \40921 , \40920 , \20528 );
nor \U$40545 ( \40922 , \40919 , \40921 );
not \U$40546 ( \40923 , \40922 );
or \U$40547 ( \40924 , \40923 , \11046 );
or \U$40548 ( \40925 , \40889 , \11039 );
nand \U$40549 ( \40926 , \40924 , \40925 );
xor \U$40550 ( \40927 , \40918 , \40926 );
not \U$40551 ( \40928 , \11965 );
and \U$40552 ( \40929 , RIc225b70_57, \12845 );
not \U$40553 ( \40930 , RIc225b70_57);
and \U$40554 ( \40931 , \40930 , \12846 );
nor \U$40555 ( \40932 , \40929 , \40931 );
not \U$40556 ( \40933 , \40932 );
or \U$40557 ( \40934 , \40928 , \40933 );
not \U$40558 ( \40935 , \10072 );
or \U$40559 ( \40936 , \40898 , \40935 );
nand \U$40560 ( \40937 , \40934 , \40936 );
and \U$40561 ( \40938 , \40927 , \40937 );
and \U$40562 ( \40939 , \40918 , \40926 );
or \U$40563 ( \40940 , \40938 , \40939 );
xor \U$40564 ( \40941 , \40916 , \40940 );
not \U$40565 ( \40942 , \20862 );
not \U$40566 ( \40943 , \40825 );
or \U$40567 ( \40944 , \40942 , \40943 );
and \U$40568 ( \40945 , RIc225990_61, \40455 );
not \U$40569 ( \40946 , RIc225990_61);
and \U$40570 ( \40947 , \40946 , \40458 );
nor \U$40571 ( \40948 , \40945 , \40947 );
nand \U$40572 ( \40949 , \40948 , \15719 );
nand \U$40573 ( \40950 , \40944 , \40949 );
and \U$40574 ( \40951 , \40941 , \40950 );
and \U$40575 ( \40952 , \40916 , \40940 );
or \U$40576 ( \40953 , \40951 , \40952 );
and \U$40577 ( \40954 , \40907 , \40953 );
and \U$40578 ( \40955 , \40904 , \40906 );
or \U$40579 ( \40956 , \40954 , \40955 );
xor \U$40580 ( \40957 , \40708 , \40717 );
xor \U$40581 ( \40958 , \40957 , \40728 );
or \U$40582 ( \40959 , \40956 , \40958 );
and \U$40583 ( \40960 , \40882 , \40959 );
and \U$40584 ( \40961 , \40958 , \40956 );
nor \U$40585 ( \40962 , \40960 , \40961 );
nand \U$40586 ( \40963 , \40880 , \40962 );
and \U$40587 ( \40964 , \40871 , \40963 );
or \U$40588 ( \40965 , RIc225be8_56, RIc225b70_57);
nand \U$40589 ( \40966 , \40965 , \18367 );
and \U$40590 ( \40967 , RIc225be8_56, RIc225b70_57);
nor \U$40591 ( \40968 , \40967 , \8767 );
and \U$40592 ( \40969 , \40966 , \40968 );
not \U$40593 ( \40970 , \11045 );
or \U$40594 ( \40971 , \18182 , \11108 );
or \U$40595 ( \40972 , \18366 , RIc225c60_55);
nand \U$40596 ( \40973 , \40971 , \40972 );
not \U$40597 ( \40974 , \40973 );
or \U$40598 ( \40975 , \40970 , \40974 );
nand \U$40599 ( \40976 , \40922 , \11038 );
nand \U$40600 ( \40977 , \40975 , \40976 );
and \U$40601 ( \40978 , \40969 , \40977 );
not \U$40602 ( \40979 , \15164 );
and \U$40603 ( \40980 , RIc225a80_59, \20690 );
not \U$40604 ( \40981 , RIc225a80_59);
and \U$40605 ( \40982 , \40981 , \12756 );
or \U$40606 ( \40983 , \40980 , \40982 );
not \U$40607 ( \40984 , \40983 );
or \U$40608 ( \40985 , \40979 , \40984 );
nand \U$40609 ( \40986 , \40912 , \12670 );
nand \U$40610 ( \40987 , \40985 , \40986 );
xor \U$40611 ( \40988 , \40978 , \40987 );
not \U$40612 ( \40989 , \15729 );
not \U$40613 ( \40990 , \40948 );
or \U$40614 ( \40991 , \40989 , \40990 );
not \U$40615 ( \40992 , RIc225990_61);
not \U$40616 ( \40993 , \10199 );
or \U$40617 ( \40994 , \40992 , \40993 );
nand \U$40618 ( \40995 , \21976 , \12806 );
nand \U$40619 ( \40996 , \40994 , \40995 );
nand \U$40620 ( \40997 , \40996 , \15719 );
nand \U$40621 ( \40998 , \40991 , \40997 );
xor \U$40622 ( \40999 , \40988 , \40998 );
not \U$40623 ( \41000 , \40999 );
not \U$40624 ( \41001 , \12670 );
not \U$40625 ( \41002 , \40983 );
or \U$40626 ( \41003 , \41001 , \41002 );
and \U$40627 ( \41004 , RIc225a80_59, \40287 );
not \U$40628 ( \41005 , RIc225a80_59);
and \U$40629 ( \41006 , \41005 , \20519 );
nor \U$40630 ( \41007 , \41004 , \41006 );
nand \U$40631 ( \41008 , \41007 , \12665 );
nand \U$40632 ( \41009 , \41003 , \41008 );
nand \U$40633 ( \41010 , \18367 , \11038 );
not \U$40634 ( \41011 , \41010 );
not \U$40635 ( \41012 , \41011 );
not \U$40636 ( \41013 , \10072 );
and \U$40637 ( \41014 , RIc225b70_57, \20393 );
not \U$40638 ( \41015 , RIc225b70_57);
and \U$40639 ( \41016 , \41015 , \20392 );
nor \U$40640 ( \41017 , \41014 , \41016 );
not \U$40641 ( \41018 , \41017 );
or \U$40642 ( \41019 , \41013 , \41018 );
and \U$40643 ( \41020 , RIc225b70_57, \16482 );
not \U$40644 ( \41021 , RIc225b70_57);
and \U$40645 ( \41022 , \41021 , \16259 );
nor \U$40646 ( \41023 , \41020 , \41022 );
nand \U$40647 ( \41024 , \41023 , \10077 );
nand \U$40648 ( \41025 , \41019 , \41024 );
not \U$40649 ( \41026 , \41025 );
or \U$40650 ( \41027 , \41012 , \41026 );
not \U$40651 ( \41028 , \12665 );
not \U$40652 ( \41029 , RIc225a80_59);
not \U$40653 ( \41030 , \15630 );
or \U$40654 ( \41031 , \41029 , \41030 );
not \U$40655 ( \41032 , RIc225a80_59);
nand \U$40656 ( \41033 , \41032 , \12845 );
nand \U$40657 ( \41034 , \41031 , \41033 );
not \U$40658 ( \41035 , \41034 );
or \U$40659 ( \41036 , \41028 , \41035 );
nand \U$40660 ( \41037 , \10342 , \41007 );
nand \U$40661 ( \41038 , \41036 , \41037 );
not \U$40662 ( \41039 , \41025 );
nand \U$40663 ( \41040 , \41039 , \41010 );
nand \U$40664 ( \41041 , \41038 , \41040 );
nand \U$40665 ( \41042 , \41027 , \41041 );
xor \U$40666 ( \41043 , \41009 , \41042 );
not \U$40667 ( \41044 , RIc225828_64);
not \U$40668 ( \41045 , RIc2258a0_63);
not \U$40669 ( \41046 , \12100 );
or \U$40670 ( \41047 , \41045 , \41046 );
nand \U$40671 ( \41048 , \30573 , \15620 );
nand \U$40672 ( \41049 , \41047 , \41048 );
not \U$40673 ( \41050 , \41049 );
or \U$40674 ( \41051 , \41044 , \41050 );
not \U$40675 ( \41052 , RIc2258a0_63);
not \U$40676 ( \41053 , \21172 );
or \U$40677 ( \41054 , \41052 , \41053 );
nand \U$40678 ( \41055 , \10086 , \16880 );
nand \U$40679 ( \41056 , \41054 , \41055 );
nand \U$40680 ( \41057 , \41056 , \16891 );
nand \U$40681 ( \41058 , \41051 , \41057 );
and \U$40682 ( \41059 , \41043 , \41058 );
and \U$40683 ( \41060 , \41009 , \41042 );
or \U$40684 ( \41061 , \41059 , \41060 );
not \U$40685 ( \41062 , \41061 );
or \U$40686 ( \41063 , \41000 , \41062 );
or \U$40687 ( \41064 , \41061 , \40999 );
xor \U$40688 ( \41065 , \40918 , \40926 );
xor \U$40689 ( \41066 , \41065 , \40937 );
xor \U$40690 ( \41067 , \40969 , \40977 );
not \U$40691 ( \41068 , \10072 );
not \U$40692 ( \41069 , \40932 );
or \U$40693 ( \41070 , \41068 , \41069 );
nand \U$40694 ( \41071 , \41017 , \11965 );
nand \U$40695 ( \41072 , \41070 , \41071 );
xor \U$40696 ( \41073 , \41067 , \41072 );
not \U$40697 ( \41074 , \15729 );
not \U$40698 ( \41075 , \40996 );
or \U$40699 ( \41076 , \41074 , \41075 );
not \U$40700 ( \41077 , RIc225990_61);
not \U$40701 ( \41078 , \40071 );
or \U$40702 ( \41079 , \41077 , \41078 );
nand \U$40703 ( \41080 , \40441 , \10338 );
nand \U$40704 ( \41081 , \41079 , \41080 );
nand \U$40705 ( \41082 , \41081 , \15719 );
nand \U$40706 ( \41083 , \41076 , \41082 );
and \U$40707 ( \41084 , \41073 , \41083 );
and \U$40708 ( \41085 , \41067 , \41072 );
or \U$40709 ( \41086 , \41084 , \41085 );
xor \U$40710 ( \41087 , \41066 , \41086 );
not \U$40711 ( \41088 , \20159 );
not \U$40712 ( \41089 , \41049 );
or \U$40713 ( \41090 , \41088 , \41089 );
xor \U$40714 ( \41091 , \16880 , \30069 );
nand \U$40715 ( \41092 , \41091 , RIc225828_64);
nand \U$40716 ( \41093 , \41090 , \41092 );
xor \U$40717 ( \41094 , \41087 , \41093 );
nand \U$40718 ( \41095 , \41064 , \41094 );
nand \U$40719 ( \41096 , \41063 , \41095 );
xor \U$40720 ( \41097 , \40916 , \40940 );
xor \U$40721 ( \41098 , \41097 , \40950 );
xor \U$40722 ( \41099 , \41066 , \41086 );
and \U$40723 ( \41100 , \41099 , \41093 );
and \U$40724 ( \41101 , \41066 , \41086 );
or \U$40725 ( \41102 , \41100 , \41101 );
xor \U$40726 ( \41103 , \41098 , \41102 );
xor \U$40727 ( \41104 , \40978 , \40987 );
and \U$40728 ( \41105 , \41104 , \40998 );
and \U$40729 ( \41106 , \40978 , \40987 );
or \U$40730 ( \41107 , \41105 , \41106 );
not \U$40731 ( \41108 , \20159 );
not \U$40732 ( \41109 , \41091 );
or \U$40733 ( \41110 , \41108 , \41109 );
nand \U$40734 ( \41111 , RIc225828_64, \40840 );
nand \U$40735 ( \41112 , \41110 , \41111 );
xor \U$40736 ( \41113 , \41107 , \41112 );
xor \U$40737 ( \41114 , \40883 , \40891 );
xor \U$40738 ( \41115 , \41114 , \40901 );
xor \U$40739 ( \41116 , \41113 , \41115 );
xor \U$40740 ( \41117 , \41103 , \41116 );
xor \U$40741 ( \41118 , \41096 , \41117 );
xor \U$40742 ( \41119 , \41067 , \41072 );
xor \U$40743 ( \41120 , \41119 , \41083 );
not \U$40744 ( \41121 , \41120 );
xor \U$40745 ( \41122 , \41009 , \41042 );
xor \U$40746 ( \41123 , \41122 , \41058 );
not \U$40747 ( \41124 , \41123 );
or \U$40748 ( \41125 , \41121 , \41124 );
or \U$40749 ( \41126 , \41123 , \41120 );
not \U$40750 ( \41127 , RIc225828_64);
not \U$40751 ( \41128 , \41056 );
or \U$40752 ( \41129 , \41127 , \41128 );
not \U$40753 ( \41130 , RIc2258a0_63);
not \U$40754 ( \41131 , \27990 );
or \U$40755 ( \41132 , \41130 , \41131 );
nand \U$40756 ( \41133 , \21976 , \16880 );
nand \U$40757 ( \41134 , \41132 , \41133 );
nand \U$40758 ( \41135 , \41134 , \16891 );
nand \U$40759 ( \41136 , \41129 , \41135 );
not \U$40760 ( \41137 , \15719 );
not \U$40761 ( \41138 , RIc225990_61);
not \U$40762 ( \41139 , \16042 );
or \U$40763 ( \41140 , \41138 , \41139 );
nand \U$40764 ( \41141 , \12756 , \10338 );
nand \U$40765 ( \41142 , \41140 , \41141 );
not \U$40766 ( \41143 , \41142 );
or \U$40767 ( \41144 , \41137 , \41143 );
nand \U$40768 ( \41145 , \41081 , \15729 );
nand \U$40769 ( \41146 , \41144 , \41145 );
or \U$40770 ( \41147 , \41136 , \41146 );
not \U$40771 ( \41148 , \10072 );
not \U$40772 ( \41149 , \41023 );
or \U$40773 ( \41150 , \41148 , \41149 );
or \U$40774 ( \41151 , \18357 , \10074 );
or \U$40775 ( \41152 , \18356 , RIc225b70_57);
nand \U$40776 ( \41153 , \41151 , \41152 );
nand \U$40777 ( \41154 , \41153 , \10077 );
nand \U$40778 ( \41155 , \41150 , \41154 );
or \U$40779 ( \41156 , RIc225af8_58, RIc225a80_59);
nand \U$40780 ( \41157 , \41156 , \18367 );
and \U$40781 ( \41158 , RIc225af8_58, RIc225a80_59);
nor \U$40782 ( \41159 , \41158 , \15262 );
and \U$40783 ( \41160 , \41157 , \41159 );
nand \U$40784 ( \41161 , \41155 , \41160 );
not \U$40785 ( \41162 , \41161 );
nand \U$40786 ( \41163 , \41147 , \41162 );
nand \U$40787 ( \41164 , \41136 , \41146 );
nand \U$40788 ( \41165 , \41163 , \41164 );
nand \U$40789 ( \41166 , \41126 , \41165 );
nand \U$40790 ( \41167 , \41125 , \41166 );
not \U$40791 ( \41168 , \41167 );
xor \U$40792 ( \41169 , \40999 , \41061 );
xnor \U$40793 ( \41170 , \41169 , \41094 );
nand \U$40794 ( \41171 , \41168 , \41170 );
not \U$40795 ( \41172 , \41171 );
and \U$40796 ( \41173 , \41025 , \41010 );
not \U$40797 ( \41174 , \41025 );
and \U$40798 ( \41175 , \41174 , \41011 );
nor \U$40799 ( \41176 , \41173 , \41175 );
not \U$40800 ( \41177 , \41176 );
not \U$40801 ( \41178 , \41038 );
and \U$40802 ( \41179 , \41177 , \41178 );
and \U$40803 ( \41180 , \41038 , \41176 );
nor \U$40804 ( \41181 , \41179 , \41180 );
not \U$40805 ( \41182 , \10342 );
not \U$40806 ( \41183 , \41034 );
or \U$40807 ( \41184 , \41182 , \41183 );
and \U$40808 ( \41185 , RIc225a80_59, \21097 );
not \U$40809 ( \41186 , RIc225a80_59);
and \U$40810 ( \41187 , \41186 , \21094 );
nor \U$40811 ( \41188 , \41185 , \41187 );
nand \U$40812 ( \41189 , \41188 , \12665 );
nand \U$40813 ( \41190 , \41184 , \41189 );
not \U$40814 ( \41191 , \15729 );
not \U$40815 ( \41192 , \41142 );
or \U$40816 ( \41193 , \41191 , \41192 );
not \U$40817 ( \41194 , RIc225990_61);
not \U$40818 ( \41195 , \30815 );
or \U$40819 ( \41196 , \41194 , \41195 );
nand \U$40820 ( \41197 , \19721 , \12806 );
nand \U$40821 ( \41198 , \41196 , \41197 );
nand \U$40822 ( \41199 , \41198 , \15719 );
nand \U$40823 ( \41200 , \41193 , \41199 );
or \U$40824 ( \41201 , \41190 , \41200 );
xor \U$40825 ( \41202 , \41155 , \41160 );
nand \U$40826 ( \41203 , \41201 , \41202 );
nand \U$40827 ( \41204 , \41200 , \41190 );
and \U$40828 ( \41205 , \41203 , \41204 );
xor \U$40829 ( \41206 , \41181 , \41205 );
xor \U$40830 ( \41207 , \41161 , \41146 );
xor \U$40831 ( \41208 , \41207 , \41136 );
xor \U$40832 ( \41209 , \41206 , \41208 );
and \U$40833 ( \41210 , \18367 , \10072 );
not \U$40834 ( \41211 , \10342 );
not \U$40835 ( \41212 , \41188 );
or \U$40836 ( \41213 , \41211 , \41212 );
and \U$40837 ( \41214 , RIc225a80_59, \16482 );
not \U$40838 ( \41215 , RIc225a80_59);
and \U$40839 ( \41216 , \41215 , \30827 );
nor \U$40840 ( \41217 , \41214 , \41216 );
nand \U$40841 ( \41218 , \41217 , \12665 );
nand \U$40842 ( \41219 , \41213 , \41218 );
xor \U$40843 ( \41220 , \41210 , \41219 );
not \U$40844 ( \41221 , \12803 );
not \U$40845 ( \41222 , \41198 );
or \U$40846 ( \41223 , \41221 , \41222 );
and \U$40847 ( \41224 , RIc225990_61, \12844 );
not \U$40848 ( \41225 , RIc225990_61);
and \U$40849 ( \41226 , \41225 , \12846 );
nor \U$40850 ( \41227 , \41224 , \41226 );
nand \U$40851 ( \41228 , \41227 , \15719 );
nand \U$40852 ( \41229 , \41223 , \41228 );
and \U$40853 ( \41230 , \41220 , \41229 );
and \U$40854 ( \41231 , \41210 , \41219 );
or \U$40855 ( \41232 , \41230 , \41231 );
not \U$40856 ( \41233 , \16891 );
not \U$40857 ( \41234 , RIc2258a0_63);
not \U$40858 ( \41235 , \21084 );
or \U$40859 ( \41236 , \41234 , \41235 );
not \U$40860 ( \41237 , \40071 );
nand \U$40861 ( \41238 , \41237 , \16880 );
nand \U$40862 ( \41239 , \41236 , \41238 );
not \U$40863 ( \41240 , \41239 );
or \U$40864 ( \41241 , \41233 , \41240 );
nand \U$40865 ( \41242 , \41134 , RIc225828_64);
nand \U$40866 ( \41243 , \41241 , \41242 );
or \U$40867 ( \41244 , \41232 , \41243 );
xor \U$40868 ( \41245 , \41190 , \41202 );
xor \U$40869 ( \41246 , \41245 , \41200 );
nand \U$40870 ( \41247 , \41244 , \41246 );
nand \U$40871 ( \41248 , \41232 , \41243 );
and \U$40872 ( \41249 , \41247 , \41248 );
nand \U$40873 ( \41250 , \41209 , \41249 );
not \U$40874 ( \41251 , \41165 );
not \U$40875 ( \41252 , \41251 );
not \U$40876 ( \41253 , \41120 );
and \U$40877 ( \41254 , \41252 , \41253 );
and \U$40878 ( \41255 , \41251 , \41120 );
nor \U$40879 ( \41256 , \41254 , \41255 );
not \U$40880 ( \41257 , \41256 );
not \U$40881 ( \41258 , \41123 );
and \U$40882 ( \41259 , \41257 , \41258 );
and \U$40883 ( \41260 , \41123 , \41256 );
nor \U$40884 ( \41261 , \41259 , \41260 );
xor \U$40885 ( \41262 , \41181 , \41205 );
and \U$40886 ( \41263 , \41262 , \41208 );
and \U$40887 ( \41264 , \41181 , \41205 );
or \U$40888 ( \41265 , \41263 , \41264 );
nand \U$40889 ( \41266 , \41261 , \41265 );
and \U$40890 ( \41267 , \41250 , \41266 );
not \U$40891 ( \41268 , \41267 );
or \U$40892 ( \41269 , RIc225a08_60, RIc225990_61);
nand \U$40893 ( \41270 , \41269 , \18367 );
and \U$40894 ( \41271 , RIc225a08_60, RIc225990_61);
nor \U$40895 ( \41272 , \41271 , \17064 );
and \U$40896 ( \41273 , \41270 , \41272 );
not \U$40897 ( \41274 , \10342 );
not \U$40898 ( \41275 , \41217 );
or \U$40899 ( \41276 , \41274 , \41275 );
and \U$40900 ( \41277 , RIc225a80_59, \18366 );
not \U$40901 ( \41278 , RIc225a80_59);
and \U$40902 ( \41279 , \41278 , \16248 );
nor \U$40903 ( \41280 , \41277 , \41279 );
not \U$40904 ( \41281 , \10341 );
or \U$40905 ( \41282 , \41280 , \41281 );
nand \U$40906 ( \41283 , \41276 , \41282 );
and \U$40907 ( \41284 , \41273 , \41283 );
not \U$40908 ( \41285 , RIc225828_64);
not \U$40909 ( \41286 , \41239 );
or \U$40910 ( \41287 , \41285 , \41286 );
and \U$40911 ( \41288 , RIc2258a0_63, \34502 );
not \U$40912 ( \41289 , RIc2258a0_63);
and \U$40913 ( \41290 , \41289 , \20693 );
nor \U$40914 ( \41291 , \41288 , \41290 );
nand \U$40915 ( \41292 , \41291 , \16891 );
nand \U$40916 ( \41293 , \41287 , \41292 );
xor \U$40917 ( \41294 , \41284 , \41293 );
xor \U$40918 ( \41295 , \41210 , \41219 );
xor \U$40919 ( \41296 , \41295 , \41229 );
and \U$40920 ( \41297 , \41294 , \41296 );
and \U$40921 ( \41298 , \41284 , \41293 );
or \U$40922 ( \41299 , \41297 , \41298 );
xor \U$40923 ( \41300 , \41243 , \41232 );
xor \U$40924 ( \41301 , \41300 , \41246 );
xor \U$40925 ( \41302 , \41299 , \41301 );
not \U$40926 ( \41303 , \12803 );
not \U$40927 ( \41304 , \41227 );
or \U$40928 ( \41305 , \41303 , \41304 );
and \U$40929 ( \41306 , RIc225990_61, \13487 );
not \U$40930 ( \41307 , RIc225990_61);
and \U$40931 ( \41308 , \41307 , \30679 );
nor \U$40932 ( \41309 , \41306 , \41308 );
nand \U$40933 ( \41310 , \41309 , \15719 );
nand \U$40934 ( \41311 , \41305 , \41310 );
xor \U$40935 ( \41312 , \41273 , \41283 );
xor \U$40936 ( \41313 , \41311 , \41312 );
not \U$40937 ( \41314 , RIc225828_64);
not \U$40938 ( \41315 , \41291 );
or \U$40939 ( \41316 , \41314 , \41315 );
not \U$40940 ( \41317 , RIc2258a0_63);
not \U$40941 ( \41318 , \15444 );
or \U$40942 ( \41319 , \41317 , \41318 );
nand \U$40943 ( \41320 , \19721 , \39744 );
nand \U$40944 ( \41321 , \41319 , \41320 );
nand \U$40945 ( \41322 , \41321 , \16891 );
nand \U$40946 ( \41323 , \41316 , \41322 );
and \U$40947 ( \41324 , \41313 , \41323 );
and \U$40948 ( \41325 , \41311 , \41312 );
or \U$40949 ( \41326 , \41324 , \41325 );
xor \U$40950 ( \41327 , \41284 , \41293 );
xor \U$40951 ( \41328 , \41327 , \41296 );
xor \U$40952 ( \41329 , \41326 , \41328 );
and \U$40953 ( \41330 , \16248 , \10342 );
not \U$40954 ( \41331 , \12803 );
not \U$40955 ( \41332 , \41309 );
or \U$40956 ( \41333 , \41331 , \41332 );
and \U$40957 ( \41334 , \16256 , RIc225990_61);
not \U$40958 ( \41335 , \16256 );
and \U$40959 ( \41336 , \41335 , \12806 );
nor \U$40960 ( \41337 , \41334 , \41336 );
nand \U$40961 ( \41338 , \41337 , \12811 );
nand \U$40962 ( \41339 , \41333 , \41338 );
xor \U$40963 ( \41340 , \41330 , \41339 );
not \U$40964 ( \41341 , RIc225828_64);
not \U$40965 ( \41342 , \41321 );
or \U$40966 ( \41343 , \41341 , \41342 );
not \U$40967 ( \41344 , RIc2258a0_63);
not \U$40968 ( \41345 , \15629 );
or \U$40969 ( \41346 , \41344 , \41345 );
nand \U$40970 ( \41347 , \12845 , \37494 );
nand \U$40971 ( \41348 , \41346 , \41347 );
nand \U$40972 ( \41349 , \41348 , \16890 );
nand \U$40973 ( \41350 , \41343 , \41349 );
and \U$40974 ( \41351 , \41340 , \41350 );
and \U$40975 ( \41352 , \41330 , \41339 );
or \U$40976 ( \41353 , \41351 , \41352 );
xor \U$40977 ( \41354 , \41311 , \41312 );
xor \U$40978 ( \41355 , \41354 , \41323 );
xor \U$40979 ( \41356 , \41353 , \41355 );
or \U$40980 ( \41357 , RIc225918_62, RIc2258a0_63);
nand \U$40981 ( \41358 , \41357 , \18357 );
and \U$40982 ( \41359 , RIc225918_62, RIc2258a0_63);
nor \U$40983 ( \41360 , \41359 , \12806 );
and \U$40984 ( \41361 , \41358 , \41360 );
not \U$40985 ( \41362 , \12811 );
or \U$40986 ( \41363 , \18367 , \10338 );
or \U$40987 ( \41364 , \18181 , RIc225990_61);
nand \U$40988 ( \41365 , \41363 , \41364 );
not \U$40989 ( \41366 , \41365 );
or \U$40990 ( \41367 , \41362 , \41366 );
nand \U$40991 ( \41368 , \41337 , \12803 );
nand \U$40992 ( \41369 , \41367 , \41368 );
and \U$40993 ( \41370 , \41361 , \41369 );
not \U$40994 ( \41371 , \41348 );
or \U$40995 ( \41372 , \41371 , \16882 );
not \U$40996 ( \41373 , \13487 );
not \U$40997 ( \41374 , \16880 );
and \U$40998 ( \41375 , \41373 , \41374 );
and \U$40999 ( \41376 , \13487 , \28750 );
nor \U$41000 ( \41377 , \41375 , \41376 );
not \U$41001 ( \41378 , \41377 );
nand \U$41002 ( \41379 , \41378 , \16890 );
nand \U$41003 ( \41380 , \41372 , \41379 );
xor \U$41004 ( \41381 , \41361 , \41369 );
nor \U$41005 ( \41382 , \41380 , \41381 );
nor \U$41006 ( \41383 , \18181 , \12804 );
not \U$41007 ( \41384 , \16248 );
not \U$41008 ( \41385 , \16889 );
and \U$41009 ( \41386 , \41384 , \41385 );
and \U$41010 ( \41387 , RIc2258a0_63, \16259 );
not \U$41011 ( \41388 , RIc2258a0_63);
and \U$41012 ( \41389 , \41388 , \16256 );
or \U$41013 ( \41390 , \41387 , \41389 );
and \U$41014 ( \41391 , \41390 , RIc225828_64);
nor \U$41015 ( \41392 , \41386 , \41391 );
and \U$41016 ( \41393 , \16248 , RIc225828_64);
not \U$41017 ( \41394 , \41393 );
nand \U$41018 ( \41395 , \41394 , RIc2258a0_63);
nor \U$41019 ( \41396 , \41392 , \41395 );
xor \U$41020 ( \41397 , \41383 , \41396 );
or \U$41021 ( \41398 , \41377 , \16882 );
nand \U$41022 ( \41399 , \41390 , \16890 );
nand \U$41023 ( \41400 , \41398 , \41399 );
and \U$41024 ( \41401 , \41397 , \41400 );
and \U$41025 ( \41402 , \41383 , \41396 );
or \U$41026 ( \41403 , \41401 , \41402 );
not \U$41027 ( \41404 , \41403 );
or \U$41028 ( \41405 , \41382 , \41404 );
nand \U$41029 ( \41406 , \41380 , \41381 );
nand \U$41030 ( \41407 , \41405 , \41406 );
xor \U$41031 ( \41408 , \41370 , \41407 );
xor \U$41032 ( \41409 , \41330 , \41339 );
xor \U$41033 ( \41410 , \41409 , \41350 );
and \U$41034 ( \41411 , \41408 , \41410 );
and \U$41035 ( \41412 , \41370 , \41407 );
or \U$41036 ( \41413 , \41411 , \41412 );
and \U$41037 ( \41414 , \41356 , \41413 );
and \U$41038 ( \41415 , \41353 , \41355 );
or \U$41039 ( \41416 , \41414 , \41415 );
and \U$41040 ( \41417 , \41329 , \41416 );
and \U$41041 ( \41418 , \41326 , \41328 );
or \U$41042 ( \41419 , \41417 , \41418 );
and \U$41043 ( \41420 , \41302 , \41419 );
and \U$41044 ( \41421 , \41299 , \41301 );
or \U$41045 ( \41422 , \41420 , \41421 );
not \U$41046 ( \41423 , \41422 );
or \U$41047 ( \41424 , \41268 , \41423 );
nor \U$41048 ( \41425 , \41209 , \41249 );
nand \U$41049 ( \41426 , \41266 , \41425 );
not \U$41050 ( \41427 , \41261 );
not \U$41051 ( \41428 , \41265 );
nand \U$41052 ( \41429 , \41427 , \41428 );
and \U$41053 ( \41430 , \41426 , \41429 );
nand \U$41054 ( \41431 , \41424 , \41430 );
not \U$41055 ( \41432 , \41431 );
or \U$41056 ( \41433 , \41172 , \41432 );
not \U$41057 ( \41434 , \41170 );
nand \U$41058 ( \41435 , \41434 , \41167 );
nand \U$41059 ( \41436 , \41433 , \41435 );
and \U$41060 ( \41437 , \41118 , \41436 );
and \U$41061 ( \41438 , \41096 , \41117 );
or \U$41062 ( \41439 , \41437 , \41438 );
xor \U$41063 ( \41440 , \40958 , \40956 );
xor \U$41064 ( \41441 , \40882 , \41440 );
xor \U$41065 ( \41442 , \40666 , \40675 );
xor \U$41066 ( \41443 , \41442 , \40686 );
xor \U$41067 ( \41444 , \40829 , \40842 );
xor \U$41068 ( \41445 , \41443 , \41444 );
xor \U$41069 ( \41446 , \41107 , \41112 );
and \U$41070 ( \41447 , \41446 , \41115 );
and \U$41071 ( \41448 , \41107 , \41112 );
or \U$41072 ( \41449 , \41447 , \41448 );
xor \U$41073 ( \41450 , \41445 , \41449 );
xor \U$41074 ( \41451 , \40904 , \40906 );
xor \U$41075 ( \41452 , \41451 , \40953 );
and \U$41076 ( \41453 , \41450 , \41452 );
and \U$41077 ( \41454 , \41445 , \41449 );
or \U$41078 ( \41455 , \41453 , \41454 );
nor \U$41079 ( \41456 , \41441 , \41455 );
xor \U$41080 ( \41457 , \41445 , \41449 );
xor \U$41081 ( \41458 , \41457 , \41452 );
xor \U$41082 ( \41459 , \41098 , \41102 );
and \U$41083 ( \41460 , \41459 , \41116 );
and \U$41084 ( \41461 , \41098 , \41102 );
or \U$41085 ( \41462 , \41460 , \41461 );
nor \U$41086 ( \41463 , \41458 , \41462 );
nor \U$41087 ( \41464 , \41456 , \41463 );
nand \U$41088 ( \41465 , \40964 , \41439 , \41464 );
not \U$41089 ( \41466 , \40963 );
nand \U$41090 ( \41467 , \41458 , \41462 );
or \U$41091 ( \41468 , \41456 , \41467 );
nand \U$41092 ( \41469 , \41441 , \41455 );
nand \U$41093 ( \41470 , \41468 , \41469 );
not \U$41094 ( \41471 , \41470 );
or \U$41095 ( \41472 , \41466 , \41471 );
not \U$41096 ( \41473 , \40880 );
not \U$41097 ( \41474 , \40962 );
nand \U$41098 ( \41475 , \41473 , \41474 );
nand \U$41099 ( \41476 , \41472 , \41475 );
buf \U$41100 ( \41477 , \40871 );
nand \U$41101 ( \41478 , \41476 , \41477 );
not \U$41102 ( \41479 , \40870 );
nand \U$41103 ( \41480 , \41479 , \40861 );
nand \U$41104 ( \41481 , \41465 , \41478 , \41480 );
and \U$41105 ( \41482 , \40773 , \40758 );
nand \U$41106 ( \41483 , \40776 , \41481 , \41482 );
or \U$41107 ( \41484 , \40768 , \40772 );
nand \U$41108 ( \41485 , \40774 , \41483 , \41484 );
or \U$41109 ( \41486 , \40256 , \40357 );
and \U$41110 ( \41487 , \40360 , \41486 );
not \U$41111 ( \41488 , \40388 );
and \U$41112 ( \41489 , \40402 , \41487 , \41488 );
nand \U$41113 ( \41490 , \40409 , \41485 , \41489 );
not \U$41114 ( \41491 , \41490 );
or \U$41115 ( \41492 , \40408 , \41491 );
xor \U$41116 ( \41493 , \37479 , \37514 );
xor \U$41117 ( \41494 , \41493 , \37579 );
not \U$41118 ( \41495 , \41494 );
xor \U$41119 ( \41496 , \37608 , \37618 );
xor \U$41120 ( \41497 , \41496 , \37615 );
not \U$41121 ( \41498 , \41497 );
not \U$41122 ( \41499 , \41498 );
or \U$41123 ( \41500 , \41495 , \41499 );
not \U$41124 ( \41501 , \41494 );
not \U$41125 ( \41502 , \41501 );
not \U$41126 ( \41503 , \41497 );
or \U$41127 ( \41504 , \41502 , \41503 );
not \U$41128 ( \41505 , \39107 );
nand \U$41129 ( \41506 , \41505 , \39111 );
not \U$41130 ( \41507 , \41506 );
not \U$41131 ( \41508 , \39115 );
or \U$41132 ( \41509 , \41507 , \41508 );
nand \U$41133 ( \41510 , \39112 , \39107 );
nand \U$41134 ( \41511 , \41509 , \41510 );
nand \U$41135 ( \41512 , \41504 , \41511 );
nand \U$41136 ( \41513 , \41500 , \41512 );
xor \U$41137 ( \41514 , \39118 , \39131 );
and \U$41138 ( \41515 , \41514 , \39161 );
and \U$41139 ( \41516 , \39118 , \39131 );
or \U$41140 ( \41517 , \41515 , \41516 );
xor \U$41141 ( \41518 , \37390 , \37439 );
xor \U$41142 ( \41519 , \41518 , \37474 );
xor \U$41143 ( \41520 , \39120 , \39125 );
and \U$41144 ( \41521 , \41520 , \39130 );
and \U$41145 ( \41522 , \39120 , \39125 );
or \U$41146 ( \41523 , \41521 , \41522 );
xor \U$41147 ( \41524 , \41519 , \41523 );
xor \U$41148 ( \41525 , \38433 , \38435 );
and \U$41149 ( \41526 , \41525 , \38488 );
and \U$41150 ( \41527 , \38433 , \38435 );
or \U$41151 ( \41528 , \41526 , \41527 );
xor \U$41152 ( \41529 , \41524 , \41528 );
xor \U$41153 ( \41530 , \41517 , \41529 );
xor \U$41154 ( \41531 , \38489 , \38629 );
and \U$41155 ( \41532 , \41531 , \38740 );
and \U$41156 ( \41533 , \38489 , \38629 );
or \U$41157 ( \41534 , \41532 , \41533 );
and \U$41158 ( \41535 , \41530 , \41534 );
and \U$41159 ( \41536 , \41517 , \41529 );
or \U$41160 ( \41537 , \41535 , \41536 );
xor \U$41161 ( \41538 , \41513 , \41537 );
not \U$41162 ( \41539 , \37622 );
not \U$41163 ( \41540 , \37600 );
or \U$41164 ( \41541 , \41539 , \41540 );
nand \U$41165 ( \41542 , \37623 , \37599 );
nand \U$41166 ( \41543 , \41541 , \41542 );
not \U$41167 ( \41544 , \37603 );
and \U$41168 ( \41545 , \41543 , \41544 );
not \U$41169 ( \41546 , \41543 );
and \U$41170 ( \41547 , \41546 , \37603 );
nor \U$41171 ( \41548 , \41545 , \41547 );
not \U$41172 ( \41549 , \41548 );
not \U$41173 ( \41550 , \41549 );
not \U$41174 ( \41551 , \41528 );
not \U$41175 ( \41552 , \41519 );
nand \U$41176 ( \41553 , \41551 , \41552 );
and \U$41177 ( \41554 , \41553 , \41523 );
not \U$41178 ( \41555 , \41528 );
nor \U$41179 ( \41556 , \41555 , \41552 );
nor \U$41180 ( \41557 , \41554 , \41556 );
not \U$41181 ( \41558 , \41557 );
xor \U$41182 ( \41559 , \37477 , \37582 );
xor \U$41183 ( \41560 , \41559 , \37588 );
not \U$41184 ( \41561 , \41560 );
or \U$41185 ( \41562 , \41558 , \41561 );
or \U$41186 ( \41563 , \41560 , \41557 );
nand \U$41187 ( \41564 , \41562 , \41563 );
not \U$41188 ( \41565 , \41564 );
not \U$41189 ( \41566 , \41565 );
or \U$41190 ( \41567 , \41550 , \41566 );
nand \U$41191 ( \41568 , \41548 , \41564 );
nand \U$41192 ( \41569 , \41567 , \41568 );
xor \U$41193 ( \41570 , \41538 , \41569 );
not \U$41194 ( \41571 , \41570 );
xor \U$41195 ( \41572 , \41517 , \41529 );
xor \U$41196 ( \41573 , \41572 , \41534 );
not \U$41197 ( \41574 , \41573 );
not \U$41198 ( \41575 , \41494 );
not \U$41199 ( \41576 , \41511 );
not \U$41200 ( \41577 , \41576 );
or \U$41201 ( \41578 , \41575 , \41577 );
or \U$41202 ( \41579 , \41576 , \41494 );
nand \U$41203 ( \41580 , \41578 , \41579 );
and \U$41204 ( \41581 , \41580 , \41497 );
not \U$41205 ( \41582 , \41580 );
and \U$41206 ( \41583 , \41582 , \41498 );
nor \U$41207 ( \41584 , \41581 , \41583 );
nand \U$41208 ( \41585 , \41574 , \41584 );
xor \U$41209 ( \41586 , \39116 , \39162 );
and \U$41210 ( \41587 , \41586 , \39185 );
and \U$41211 ( \41588 , \39116 , \39162 );
or \U$41212 ( \41589 , \41587 , \41588 );
and \U$41213 ( \41590 , \41585 , \41589 );
not \U$41214 ( \41591 , \41573 );
nor \U$41215 ( \41592 , \41591 , \41584 );
nor \U$41216 ( \41593 , \41590 , \41592 );
nand \U$41217 ( \41594 , \41571 , \41593 );
xor \U$41218 ( \41595 , \41584 , \41589 );
xnor \U$41219 ( \41596 , \41595 , \41573 );
or \U$41220 ( \41597 , \39186 , \38741 );
not \U$41221 ( \41598 , \41597 );
not \U$41222 ( \41599 , \39073 );
or \U$41223 ( \41600 , \41598 , \41599 );
nand \U$41224 ( \41601 , \39186 , \38741 );
nand \U$41225 ( \41602 , \41600 , \41601 );
or \U$41226 ( \41603 , \41596 , \41602 );
and \U$41227 ( \41604 , \41594 , \41603 );
and \U$41228 ( \41605 , \37357 , \37345 );
not \U$41229 ( \41606 , \37357 );
and \U$41230 ( \41607 , \41606 , \37344 );
nor \U$41231 ( \41608 , \41605 , \41607 );
xnor \U$41232 ( \41609 , \41608 , \37361 );
not \U$41233 ( \41610 , \41560 );
nand \U$41234 ( \41611 , \41610 , \41557 );
not \U$41235 ( \41612 , \41611 );
not \U$41236 ( \41613 , \41549 );
or \U$41237 ( \41614 , \41612 , \41613 );
not \U$41238 ( \41615 , \41557 );
nand \U$41239 ( \41616 , \41615 , \41560 );
nand \U$41240 ( \41617 , \41614 , \41616 );
not \U$41241 ( \41618 , \41617 );
xor \U$41242 ( \41619 , \41609 , \41618 );
xor \U$41243 ( \41620 , \37591 , \37594 );
xnor \U$41244 ( \41621 , \41620 , \37625 );
xor \U$41245 ( \41622 , \41619 , \41621 );
not \U$41246 ( \41623 , \41513 );
not \U$41247 ( \41624 , \41569 );
nand \U$41248 ( \41625 , \41623 , \41624 );
and \U$41249 ( \41626 , \41625 , \41537 );
not \U$41250 ( \41627 , \41513 );
nor \U$41251 ( \41628 , \41627 , \41624 );
nor \U$41252 ( \41629 , \41626 , \41628 );
nand \U$41253 ( \41630 , \41622 , \41629 );
xor \U$41254 ( \41631 , \41609 , \41618 );
and \U$41255 ( \41632 , \41631 , \41621 );
and \U$41256 ( \41633 , \41609 , \41618 );
or \U$41257 ( \41634 , \41632 , \41633 );
xor \U$41258 ( \41635 , \37632 , \37627 );
xnor \U$41259 ( \41636 , \41635 , \37635 );
nand \U$41260 ( \41637 , \41634 , \41636 );
and \U$41261 ( \41638 , \41604 , \41630 , \41637 );
nand \U$41262 ( \41639 , \41492 , \41638 );
not \U$41263 ( \41640 , \41630 );
not \U$41264 ( \41641 , \41594 );
and \U$41265 ( \41642 , \41596 , \41602 );
not \U$41266 ( \41643 , \41642 );
or \U$41267 ( \41644 , \41641 , \41643 );
not \U$41268 ( \41645 , \41593 );
buf \U$41269 ( \41646 , \41570 );
nand \U$41270 ( \41647 , \41645 , \41646 );
nand \U$41271 ( \41648 , \41644 , \41647 );
not \U$41272 ( \41649 , \41648 );
or \U$41273 ( \41650 , \41640 , \41649 );
or \U$41274 ( \41651 , \41622 , \41629 );
nand \U$41275 ( \41652 , \41650 , \41651 );
and \U$41276 ( \41653 , \41652 , \41637 );
nor \U$41277 ( \41654 , \41634 , \41636 );
nor \U$41278 ( \41655 , \41653 , \41654 );
nand \U$41279 ( \41656 , \41639 , \41655 );
and \U$41280 ( \41657 , \38431 , \41656 );
buf \U$41281 ( \41658 , \38402 );
not \U$41282 ( \41659 , \41658 );
not \U$41283 ( \41660 , \38372 );
nor \U$41284 ( \41661 , \38404 , \38408 );
nand \U$41285 ( \41662 , \38395 , \41661 );
not \U$41286 ( \41663 , \38374 );
not \U$41287 ( \41664 , \38394 );
nand \U$41288 ( \41665 , \41663 , \41664 );
nand \U$41289 ( \41666 , \41662 , \41665 );
not \U$41290 ( \41667 , \41666 );
or \U$41291 ( \41668 , \41660 , \41667 );
or \U$41292 ( \41669 , \38340 , \38371 );
nand \U$41293 ( \41670 , \41668 , \41669 );
not \U$41294 ( \41671 , \41670 );
or \U$41295 ( \41672 , \41659 , \41671 );
or \U$41296 ( \41673 , \38397 , \38401 );
nand \U$41297 ( \41674 , \41672 , \41673 );
nor \U$41298 ( \41675 , \41657 , \41674 );
not \U$41299 ( \41676 , \41675 );
nand \U$41300 ( \41677 , \38421 , \41676 , \33972 );
nor \U$41301 ( \41678 , \33881 , \33885 );
nand \U$41302 ( \41679 , \33964 , \41678 );
not \U$41303 ( \41680 , \33959 );
not \U$41304 ( \41681 , \33963 );
nand \U$41305 ( \41682 , \41680 , \41681 );
nand \U$41306 ( \41683 , \41679 , \41682 );
nor \U$41307 ( \41684 , \33935 , \33956 );
or \U$41308 ( \41685 , \41683 , \41684 );
and \U$41309 ( \41686 , \33971 , \33957 );
nand \U$41310 ( \41687 , \41685 , \41686 );
or \U$41311 ( \41688 , \33970 , \33968 );
and \U$41312 ( \41689 , \41687 , \41688 );
nand \U$41313 ( \41690 , \33973 , \38422 , \41677 , \41689 );
not \U$41314 ( \41691 , \41690 );
not \U$41315 ( \41692 , \17457 );
buf \U$41316 ( \41693 , \22243 );
not \U$41317 ( \41694 , \22252 );
or \U$41318 ( \41695 , \21815 , \22238 );
and \U$41319 ( \41696 , \20831 , \41693 , \41694 , \41695 );
nand \U$41320 ( \41697 , \41692 , \22264 , \15100 , \41696 );
nor \U$41321 ( \41698 , \26611 , \41697 );
not \U$41322 ( \41699 , \41698 );
or \U$41323 ( \41700 , \41691 , \41699 );
not \U$41324 ( \41701 , \26602 );
or \U$41325 ( \41702 , \26546 , \26550 );
not \U$41326 ( \41703 , \26587 );
or \U$41327 ( \41704 , \41702 , \41703 );
or \U$41328 ( \41705 , \26582 , \26586 );
nand \U$41329 ( \41706 , \41704 , \41705 );
not \U$41330 ( \41707 , \41706 );
or \U$41331 ( \41708 , \41701 , \41707 );
or \U$41332 ( \41709 , \26597 , \26601 );
nand \U$41333 ( \41710 , \41708 , \41709 );
and \U$41334 ( \41711 , \41710 , \26609 );
nor \U$41335 ( \41712 , \26604 , \26608 );
nor \U$41336 ( \41713 , \41711 , \41712 );
nand \U$41337 ( \41714 , \41700 , \41713 );
nor \U$41338 ( \41715 , \26671 , \41714 );
not \U$41339 ( \41716 , \41715 );
not \U$41340 ( \41717 , \41716 );
or \U$41341 ( \41718 , \8766 , \41717 );
not \U$41342 ( \41719 , \8257 );
not \U$41343 ( \41720 , \41719 );
not \U$41344 ( \41721 , \7991 );
not \U$41345 ( \41722 , \8128 );
not \U$41346 ( \41723 , \5109 );
not \U$41347 ( \41724 , \6947 );
not \U$41348 ( \41725 , \5913 );
and \U$41349 ( \41726 , \6251 , \6937 );
nand \U$41350 ( \41727 , \41726 , \6244 );
not \U$41351 ( \41728 , \5916 );
not \U$41352 ( \41729 , \6243 );
nand \U$41353 ( \41730 , \41728 , \41729 );
nand \U$41354 ( \41731 , \41727 , \41730 );
not \U$41355 ( \41732 , \41731 );
or \U$41356 ( \41733 , \41725 , \41732 );
or \U$41357 ( \41734 , \5450 , \5912 );
nand \U$41358 ( \41735 , \41733 , \41734 );
not \U$41359 ( \41736 , \41735 );
or \U$41360 ( \41737 , \41724 , \41736 );
or \U$41361 ( \41738 , \6942 , \6946 );
nand \U$41362 ( \41739 , \41737 , \41738 );
not \U$41363 ( \41740 , \41739 );
or \U$41364 ( \41741 , \41723 , \41740 );
not \U$41365 ( \41742 , \5100 );
not \U$41366 ( \41743 , \5107 );
nand \U$41367 ( \41744 , \4276 , \4649 );
or \U$41368 ( \41745 , \41744 , \4273 );
nand \U$41369 ( \41746 , \3892 , \4272 );
nand \U$41370 ( \41747 , \41745 , \41746 );
not \U$41371 ( \41748 , \41747 );
or \U$41372 ( \41749 , \41743 , \41748 );
or \U$41373 ( \41750 , \5102 , \5106 );
nand \U$41374 ( \41751 , \41749 , \41750 );
not \U$41375 ( \41752 , \41751 );
or \U$41376 ( \41753 , \41742 , \41752 );
or \U$41377 ( \41754 , \5079 , \5099 );
nand \U$41378 ( \41755 , \41753 , \41754 );
not \U$41379 ( \41756 , \41755 );
nand \U$41380 ( \41757 , \41741 , \41756 );
not \U$41381 ( \41758 , \41757 );
or \U$41382 ( \41759 , \41722 , \41758 );
not \U$41383 ( \41760 , \8119 );
nor \U$41384 ( \41761 , \8092 , \8096 );
not \U$41385 ( \41762 , \41761 );
not \U$41386 ( \41763 , \8090 );
or \U$41387 ( \41764 , \41762 , \41763 );
not \U$41388 ( \41765 , \8067 );
not \U$41389 ( \41766 , \8089 );
nand \U$41390 ( \41767 , \41765 , \41766 );
nand \U$41391 ( \41768 , \41764 , \41767 );
not \U$41392 ( \41769 , \41768 );
or \U$41393 ( \41770 , \41760 , \41769 );
not \U$41394 ( \41771 , \8118 );
nand \U$41395 ( \41772 , \41771 , \8106 );
nand \U$41396 ( \41773 , \41770 , \41772 );
and \U$41397 ( \41774 , \41773 , \8126 );
nor \U$41398 ( \41775 , \8121 , \8125 );
nor \U$41399 ( \41776 , \41774 , \41775 );
nand \U$41400 ( \41777 , \41759 , \41776 );
not \U$41401 ( \41778 , \41777 );
or \U$41402 ( \41779 , \41721 , \41778 );
not \U$41403 ( \41780 , \7990 );
not \U$41404 ( \41781 , \41780 );
not \U$41405 ( \41782 , \7712 );
nand \U$41406 ( \41783 , \41782 , \7667 );
not \U$41407 ( \41784 , \7857 );
or \U$41408 ( \41785 , \41783 , \41784 );
nand \U$41409 ( \41786 , \7852 , \7856 );
nand \U$41410 ( \41787 , \41785 , \41786 );
not \U$41411 ( \41788 , \41787 );
or \U$41412 ( \41789 , \41781 , \41788 );
nand \U$41413 ( \41790 , \7985 , \7989 );
nand \U$41414 ( \41791 , \41789 , \41790 );
not \U$41415 ( \41792 , \41791 );
nand \U$41416 ( \41793 , \41779 , \41792 );
not \U$41417 ( \41794 , \41793 );
or \U$41418 ( \41795 , \41720 , \41794 );
nand \U$41419 ( \41796 , \8256 , \8133 );
nand \U$41420 ( \41797 , \41795 , \41796 );
not \U$41421 ( \41798 , \8764 );
and \U$41422 ( \41799 , \41797 , \41798 );
not \U$41423 ( \41800 , \8763 );
and \U$41424 ( \41801 , \8735 , \8750 );
not \U$41425 ( \41802 , \41801 );
not \U$41426 ( \41803 , \8661 );
not \U$41427 ( \41804 , \8583 );
nand \U$41428 ( \41805 , \8372 , \8376 );
or \U$41429 ( \41806 , \41805 , \8485 );
nand \U$41430 ( \41807 , \8480 , \8484 );
nand \U$41431 ( \41808 , \41806 , \41807 );
not \U$41432 ( \41809 , \41808 );
or \U$41433 ( \41810 , \41804 , \41809 );
nand \U$41434 ( \41811 , \8578 , \8582 );
nand \U$41435 ( \41812 , \41810 , \41811 );
not \U$41436 ( \41813 , \41812 );
or \U$41437 ( \41814 , \41803 , \41813 );
nand \U$41438 ( \41815 , \8587 , \8660 );
nand \U$41439 ( \41816 , \41814 , \41815 );
not \U$41440 ( \41817 , \41816 );
or \U$41441 ( \41818 , \41802 , \41817 );
nand \U$41442 ( \41819 , \8700 , \8704 );
or \U$41443 ( \41820 , \41819 , \8734 );
nand \U$41444 ( \41821 , \8729 , \8733 );
nand \U$41445 ( \41822 , \41820 , \41821 );
and \U$41446 ( \41823 , \41822 , \8750 );
and \U$41447 ( \41824 , \8745 , \8749 );
nor \U$41448 ( \41825 , \41823 , \41824 );
nand \U$41449 ( \41826 , \41818 , \41825 );
not \U$41450 ( \41827 , \41826 );
or \U$41451 ( \41828 , \41800 , \41827 );
nand \U$41452 ( \41829 , \8758 , \8762 );
nand \U$41453 ( \41830 , \41828 , \41829 );
nor \U$41454 ( \41831 , \41799 , \41830 );
nand \U$41455 ( \41832 , \41718 , \41831 );
not \U$41456 ( \41833 , \41832 );
or \U$41457 ( \41834 , \1902 , \41833 );
not \U$41458 ( \41835 , \1866 );
nand \U$41459 ( \41836 , \1664 , \1792 );
nor \U$41460 ( \41837 , \41836 , \1829 );
and \U$41461 ( \41838 , \1828 , \1824 );
nor \U$41462 ( \41839 , \41837 , \41838 );
or \U$41463 ( \41840 , \41839 , \1852 );
nand \U$41464 ( \41841 , \1843 , \1851 );
nand \U$41465 ( \41842 , \41840 , \41841 );
not \U$41466 ( \41843 , \41842 );
or \U$41467 ( \41844 , \41835 , \41843 );
nand \U$41468 ( \41845 , \1861 , \1865 );
nand \U$41469 ( \41846 , \41844 , \41845 );
and \U$41470 ( \41847 , \41846 , \1288 );
nand \U$41471 ( \41848 , \1188 , \1249 );
or \U$41472 ( \41849 , \41848 , \1287 );
nand \U$41473 ( \41850 , \1259 , \1286 );
nand \U$41474 ( \41851 , \41849 , \41850 );
nor \U$41475 ( \41852 , \41847 , \41851 );
not \U$41476 ( \41853 , \41852 );
not \U$41477 ( \41854 , \1900 );
and \U$41478 ( \41855 , \41853 , \41854 );
and \U$41479 ( \41856 , \1875 , \1899 );
nor \U$41480 ( \41857 , \41855 , \41856 );
nand \U$41481 ( \41858 , \41834 , \41857 );
xor \U$41482 ( \41859 , \1892 , \1893 );
and \U$41483 ( \41860 , \41859 , \1898 );
and \U$41484 ( \41861 , \1892 , \1893 );
or \U$41485 ( \41862 , \41860 , \41861 );
nand \U$41486 ( \41863 , \1271 , RIc2275b0_1);
not \U$41487 ( \41864 , \41863 );
not \U$41488 ( \41865 , \1877 );
not \U$41489 ( \41866 , \855 );
and \U$41490 ( \41867 , \41865 , \41866 );
and \U$41491 ( \41868 , \1579 , RIc2275b0_1);
nor \U$41492 ( \41869 , \41867 , \41868 );
not \U$41493 ( \41870 , \41869 );
or \U$41494 ( \41871 , \41864 , \41870 );
or \U$41495 ( \41872 , \41869 , \41863 );
nand \U$41496 ( \41873 , \41871 , \41872 );
not \U$41497 ( \41874 , \41873 );
and \U$41498 ( \41875 , \1879 , \1885 );
nor \U$41499 ( \41876 , \41875 , \1887 );
not \U$41500 ( \41877 , \41876 );
or \U$41501 ( \41878 , \41874 , \41877 );
or \U$41502 ( \41879 , \41876 , \41873 );
nand \U$41503 ( \41880 , \41878 , \41879 );
xor \U$41504 ( \41881 , \41862 , \41880 );
xnor \U$41505 ( \41882 , \41858 , \41881 );
xor \U$41506 ( \41883 , RIc22c560_231, RIc22cb78_244);
xnor \U$41507 ( \41884 , RIc22c218_224, RIc22b660_199);
xnor \U$41508 ( \41885 , \41883 , \41884 );
xor \U$41509 ( \41886 , RIc22b840_203, RIc22cd58_248);
xor \U$41510 ( \41887 , RIc22b9a8_206, RIc22c038_220);
xor \U$41511 ( \41888 , \41886 , \41887 );
xor \U$41512 ( \41889 , \41885 , \41888 );
xnor \U$41513 ( \41890 , RIc22c0b0_221, RIc22b930_205);
xor \U$41514 ( \41891 , RIc22c740_235, RIc22cc68_246);
xor \U$41515 ( \41892 , \41890 , \41891 );
xor \U$41516 ( \41893 , RIc22bc00_211, RIc22cce0_247);
xnor \U$41517 ( \41894 , RIc22bed0_217, RIc22bcf0_213);
xnor \U$41518 ( \41895 , \41893 , \41894 );
xor \U$41519 ( \41896 , \41892 , \41895 );
xor \U$41520 ( \41897 , \41889 , \41896 );
not \U$41521 ( \41898 , \41897 );
xor \U$41522 ( \41899 , RIc22c8a8_238, RIc22ba20_207);
xor \U$41523 ( \41900 , RIc22c4e8_230, RIc22ce48_250);
xnor \U$41524 ( \41901 , \41899 , \41900 );
xor \U$41525 ( \41902 , RIc22b480_195, RIc22cfb0_253);
not \U$41526 ( \41903 , \41902 );
not \U$41527 ( \41904 , RIc22b6d8_200);
xor \U$41528 ( \41905 , RIc22c998_240, \41904 );
not \U$41529 ( \41906 , \41905 );
or \U$41530 ( \41907 , \41903 , \41906 );
or \U$41531 ( \41908 , \41905 , \41902 );
nand \U$41532 ( \41909 , \41907 , \41908 );
or \U$41533 ( \41910 , \41901 , \41909 );
nand \U$41534 ( \41911 , \41901 , \41909 );
nand \U$41535 ( \41912 , \41910 , \41911 );
xor \U$41536 ( \41913 , RIc22b8b8_204, RIc22c920_239);
xor \U$41537 ( \41914 , RIc22b7c8_202, RIc22c128_222);
xor \U$41538 ( \41915 , \41913 , \41914 );
xor \U$41539 ( \41916 , RIc22c6c8_234, RIc22d028_254);
xnor \U$41540 ( \41917 , RIc22c650_233, RIc22c5d8_232);
xnor \U$41541 ( \41918 , \41916 , \41917 );
xor \U$41542 ( \41919 , \41915 , \41918 );
xor \U$41543 ( \41920 , \41912 , \41919 );
not \U$41544 ( \41921 , \41920 );
and \U$41545 ( \41922 , \41898 , \41921 );
and \U$41546 ( \41923 , \41897 , \41920 );
nor \U$41547 ( \41924 , \41922 , \41923 );
xnor \U$41548 ( \41925 , RIc22bde0_215, RIc22bd68_214);
xor \U$41549 ( \41926 , RIc22be58_216, RIc22c7b8_236);
xor \U$41550 ( \41927 , \41925 , \41926 );
xor \U$41551 ( \41928 , RIc22b408_194, RIc22d0a0_255);
xor \U$41552 ( \41929 , RIc22b750_201, RIc22c1a0_223);
xor \U$41553 ( \41930 , \41928 , \41929 );
or \U$41554 ( \41931 , \41927 , \41930 );
nand \U$41555 ( \41932 , \41927 , \41930 );
nand \U$41556 ( \41933 , \41931 , \41932 );
xor \U$41557 ( \41934 , RIc22bb88_210, RIc22cf38_252);
xor \U$41558 ( \41935 , RIc22bc78_212, RIc22c830_237);
xor \U$41559 ( \41936 , \41934 , \41935 );
not \U$41560 ( \41937 , \41936 );
xnor \U$41561 ( \41938 , RIc22c290_225, RIc22b5e8_198);
not \U$41562 ( \41939 , \41938 );
xor \U$41563 ( \41940 , RIc22cbf0_245, RIc22cec0_251);
not \U$41564 ( \41941 , \41940 );
and \U$41565 ( \41942 , \41939 , \41941 );
and \U$41566 ( \41943 , \41938 , \41940 );
nor \U$41567 ( \41944 , \41942 , \41943 );
not \U$41568 ( \41945 , \41944 );
or \U$41569 ( \41946 , \41937 , \41945 );
or \U$41570 ( \41947 , \41944 , \41936 );
nand \U$41571 ( \41948 , \41946 , \41947 );
xnor \U$41572 ( \41949 , \41933 , \41948 );
not \U$41573 ( \41950 , \41949 );
xnor \U$41574 ( \41951 , RIc22bf48_218, RIc22bb10_209);
xor \U$41575 ( \41952 , RIc22c3f8_228, RIc22ca88_242);
xor \U$41576 ( \41953 , \41951 , \41952 );
xor \U$41577 ( \41954 , RIc22b4f8_196, RIc22cdd0_249);
xor \U$41578 ( \41955 , RIc22ba98_208, RIc22bfc0_219);
xor \U$41579 ( \41956 , \41954 , \41955 );
or \U$41580 ( \41957 , \41953 , \41956 );
nand \U$41581 ( \41958 , \41953 , \41956 );
nand \U$41582 ( \41959 , \41957 , \41958 );
xor \U$41583 ( \41960 , RIc22ca10_241, RIc22b570_197);
xor \U$41584 ( \41961 , RIc22c470_229, RIc22cb00_243);
xnor \U$41585 ( \41962 , \41960 , \41961 );
xor \U$41586 ( \41963 , RIc22b390_193, RIc22d118_256);
not \U$41587 ( \41964 , \41963 );
xnor \U$41588 ( \41965 , RIc22c380_227, RIc22c308_226);
not \U$41589 ( \41966 , \41965 );
or \U$41590 ( \41967 , \41964 , \41966 );
or \U$41591 ( \41968 , \41965 , \41963 );
nand \U$41592 ( \41969 , \41967 , \41968 );
xor \U$41593 ( \41970 , \41962 , \41969 );
xnor \U$41594 ( \41971 , \41959 , \41970 );
not \U$41595 ( \41972 , \41971 );
or \U$41596 ( \41973 , \41950 , \41972 );
or \U$41597 ( \41974 , \41971 , \41949 );
nand \U$41598 ( \41975 , \41973 , \41974 );
xor \U$41599 ( \41976 , \41924 , \41975 );
not \U$41600 ( \41977 , \41976 );
not \U$41601 ( \41978 , \41977 );
not \U$41602 ( \41979 , \41978 );
buf \U$41603 ( \41980 , \41979 );
buf \U$41604 ( \41981 , \41980 );
not \U$41605 ( \41982 , \41981 );
nor \U$41606 ( \41983 , \41882 , \41982 );
buf \U$41607 ( \41984 , \41983 );
not \U$41608 ( \41985 , \1867 );
and \U$41609 ( \41986 , \41798 , \41985 , \1288 );
not \U$41610 ( \41987 , \41986 );
not \U$41611 ( \41988 , \8259 );
not \U$41612 ( \41989 , \41988 );
not \U$41613 ( \41990 , \41716 );
or \U$41614 ( \41991 , \41989 , \41990 );
not \U$41615 ( \41992 , \41797 );
nand \U$41616 ( \41993 , \41991 , \41992 );
not \U$41617 ( \41994 , \41993 );
or \U$41618 ( \41995 , \41987 , \41994 );
not \U$41619 ( \41996 , \41985 );
not \U$41620 ( \41997 , \41830 );
or \U$41621 ( \41998 , \41996 , \41997 );
not \U$41622 ( \41999 , \41846 );
nand \U$41623 ( \42000 , \41998 , \41999 );
and \U$41624 ( \42001 , \42000 , \1288 );
nor \U$41625 ( \42002 , \42001 , \41851 );
nand \U$41626 ( \42003 , \41995 , \42002 );
nor \U$41627 ( \42004 , \41856 , \1900 );
xnor \U$41628 ( \42005 , \42003 , \42004 );
nor \U$41629 ( \42006 , \42005 , \41982 );
buf \U$41630 ( \42007 , \42006 );
and \U$41631 ( \42008 , \41798 , \41985 , \1250 );
not \U$41632 ( \42009 , \42008 );
not \U$41633 ( \42010 , \41993 );
or \U$41634 ( \42011 , \42009 , \42010 );
and \U$41635 ( \42012 , \42000 , \1250 );
not \U$41636 ( \42013 , \41848 );
nor \U$41637 ( \42014 , \42012 , \42013 );
nand \U$41638 ( \42015 , \42011 , \42014 );
not \U$41639 ( \42016 , \1287 );
nand \U$41640 ( \42017 , \42016 , \41850 );
xor \U$41641 ( \42018 , \42015 , \42017 );
nor \U$41642 ( \42019 , \42018 , \41982 );
buf \U$41643 ( \42020 , \42019 );
not \U$41644 ( \42021 , \41985 );
not \U$41645 ( \42022 , \41832 );
or \U$41646 ( \42023 , \42021 , \42022 );
nand \U$41647 ( \42024 , \42023 , \41999 );
nand \U$41648 ( \42025 , \1250 , \41848 );
xor \U$41649 ( \42026 , \42024 , \42025 );
nor \U$41650 ( \42027 , \42026 , \41982 );
buf \U$41651 ( \42028 , \42027 );
not \U$41652 ( \42029 , \1853 );
nor \U$41653 ( \42030 , \42029 , \8764 );
not \U$41654 ( \42031 , \42030 );
not \U$41655 ( \42032 , \41993 );
or \U$41656 ( \42033 , \42031 , \42032 );
and \U$41657 ( \42034 , \41830 , \1853 );
nor \U$41658 ( \42035 , \42034 , \41842 );
nand \U$41659 ( \42036 , \42033 , \42035 );
nand \U$41660 ( \42037 , \1866 , \41845 );
xor \U$41661 ( \42038 , \42036 , \42037 );
nor \U$41662 ( \42039 , \42038 , \41982 );
buf \U$41663 ( \42040 , \42039 );
not \U$41664 ( \42041 , \1830 );
not \U$41665 ( \42042 , \41832 );
or \U$41666 ( \42043 , \42041 , \42042 );
nand \U$41667 ( \42044 , \42043 , \41839 );
not \U$41668 ( \42045 , \1852 );
nand \U$41669 ( \42046 , \42045 , \41841 );
xor \U$41670 ( \42047 , \42044 , \42046 );
nor \U$41671 ( \42048 , \42047 , \41982 );
buf \U$41672 ( \42049 , \42048 );
not \U$41673 ( \42050 , \1793 );
not \U$41674 ( \42051 , \42050 );
not \U$41675 ( \42052 , \41832 );
or \U$41676 ( \42053 , \42051 , \42052 );
nand \U$41677 ( \42054 , \42053 , \41836 );
nor \U$41678 ( \42055 , \41838 , \1829 );
xnor \U$41679 ( \42056 , \42054 , \42055 );
nor \U$41680 ( \42057 , \42056 , \41982 );
buf \U$41681 ( \42058 , \42057 );
nand \U$41682 ( \42059 , \41836 , \42050 );
xnor \U$41683 ( \42060 , \41832 , \42059 );
not \U$41684 ( \42061 , \42060 );
nor \U$41685 ( \42062 , \42061 , \41982 );
buf \U$41686 ( \42063 , \42062 );
and \U$41687 ( \42064 , \8662 , \41801 );
not \U$41688 ( \42065 , \42064 );
not \U$41689 ( \42066 , \41993 );
or \U$41690 ( \42067 , \42065 , \42066 );
not \U$41691 ( \42068 , \41826 );
nand \U$41692 ( \42069 , \42067 , \42068 );
nand \U$41693 ( \42070 , \8763 , \41829 );
xor \U$41694 ( \42071 , \42069 , \42070 );
nor \U$41695 ( \42072 , \42071 , \41982 );
buf \U$41696 ( \42073 , \42072 );
not \U$41697 ( \42074 , \8735 );
not \U$41698 ( \42075 , \8662 );
or \U$41699 ( \42076 , \26671 , \41714 );
and \U$41700 ( \42077 , \42076 , \41988 );
not \U$41701 ( \42078 , \42077 );
or \U$41702 ( \42079 , \42075 , \42078 );
and \U$41703 ( \42080 , \8662 , \41797 );
nor \U$41704 ( \42081 , \42080 , \41816 );
nand \U$41705 ( \42082 , \42079 , \42081 );
not \U$41706 ( \42083 , \42082 );
or \U$41707 ( \42084 , \42074 , \42083 );
not \U$41708 ( \42085 , \41822 );
nand \U$41709 ( \42086 , \42084 , \42085 );
not \U$41710 ( \42087 , \41824 );
nand \U$41711 ( \42088 , \42087 , \8750 );
xor \U$41712 ( \42089 , \42086 , \42088 );
nor \U$41713 ( \42090 , \42089 , \41982 );
buf \U$41714 ( \42091 , \42090 );
not \U$41715 ( \42092 , \8705 );
not \U$41716 ( \42093 , \42092 );
not \U$41717 ( \42094 , \42082 );
or \U$41718 ( \42095 , \42093 , \42094 );
nand \U$41719 ( \42096 , \42095 , \41819 );
not \U$41720 ( \42097 , \8734 );
nand \U$41721 ( \42098 , \42097 , \41821 );
xor \U$41722 ( \42099 , \42096 , \42098 );
nor \U$41723 ( \42100 , \42099 , \41982 );
buf \U$41724 ( \42101 , \42100 );
not \U$41725 ( \42102 , \8662 );
not \U$41726 ( \42103 , \42077 );
or \U$41727 ( \42104 , \42102 , \42103 );
nand \U$41728 ( \42105 , \42104 , \42081 );
nand \U$41729 ( \42106 , \41819 , \42092 );
xor \U$41730 ( \42107 , \42105 , \42106 );
nor \U$41731 ( \42108 , \42107 , \41982 );
buf \U$41732 ( \42109 , \42108 );
not \U$41733 ( \42110 , \8583 );
not \U$41734 ( \42111 , \8486 );
not \U$41735 ( \42112 , \42077 );
or \U$41736 ( \42113 , \42111 , \42112 );
and \U$41737 ( \42114 , \8486 , \41797 );
nor \U$41738 ( \42115 , \42114 , \41808 );
nand \U$41739 ( \42116 , \42113 , \42115 );
not \U$41740 ( \42117 , \42116 );
or \U$41741 ( \42118 , \42110 , \42117 );
nand \U$41742 ( \42119 , \42118 , \41811 );
nand \U$41743 ( \42120 , \8661 , \41815 );
xor \U$41744 ( \42121 , \42119 , \42120 );
nor \U$41745 ( \42122 , \42121 , \41982 );
buf \U$41746 ( \42123 , \42122 );
nand \U$41747 ( \42124 , \41811 , \8583 );
xor \U$41748 ( \42125 , \42116 , \42124 );
nor \U$41749 ( \42126 , \42125 , \41982 );
buf \U$41750 ( \42127 , \42126 );
not \U$41751 ( \42128 , \8377 );
not \U$41752 ( \42129 , \42128 );
not \U$41753 ( \42130 , \41993 );
or \U$41754 ( \42131 , \42129 , \42130 );
nand \U$41755 ( \42132 , \42131 , \41805 );
not \U$41756 ( \42133 , \8485 );
nand \U$41757 ( \42134 , \42133 , \41807 );
xor \U$41758 ( \42135 , \42132 , \42134 );
nor \U$41759 ( \42136 , \42135 , \41982 );
buf \U$41760 ( \42137 , \42136 );
nand \U$41761 ( \42138 , \41805 , \42128 );
xor \U$41762 ( \42139 , \41993 , \42138 );
nor \U$41763 ( \42140 , \42139 , \41982 );
buf \U$41764 ( \42141 , \42140 );
not \U$41765 ( \42142 , \8129 );
not \U$41766 ( \42143 , \42142 );
not \U$41767 ( \42144 , \6949 );
not \U$41768 ( \42145 , \41716 );
or \U$41769 ( \42146 , \42144 , \42145 );
buf \U$41770 ( \42147 , \41757 );
not \U$41771 ( \42148 , \42147 );
nand \U$41772 ( \42149 , \42146 , \42148 );
not \U$41773 ( \42150 , \42149 );
or \U$41774 ( \42151 , \42143 , \42150 );
not \U$41775 ( \42152 , \41776 );
and \U$41776 ( \42153 , \42152 , \7991 );
nor \U$41777 ( \42154 , \42153 , \41791 );
nand \U$41778 ( \42155 , \42151 , \42154 );
nand \U$41779 ( \42156 , \41719 , \41796 );
xor \U$41780 ( \42157 , \42155 , \42156 );
nor \U$41781 ( \42158 , \42157 , \41982 );
buf \U$41782 ( \42159 , \42158 );
not \U$41783 ( \42160 , \7858 );
not \U$41784 ( \42161 , \42160 );
not \U$41785 ( \42162 , \8128 );
and \U$41786 ( \42163 , \42076 , \6949 );
not \U$41787 ( \42164 , \42163 );
or \U$41788 ( \42165 , \42162 , \42164 );
not \U$41789 ( \42166 , \41777 );
nand \U$41790 ( \42167 , \42165 , \42166 );
not \U$41791 ( \42168 , \42167 );
or \U$41792 ( \42169 , \42161 , \42168 );
not \U$41793 ( \42170 , \41787 );
nand \U$41794 ( \42171 , \42169 , \42170 );
nand \U$41795 ( \42172 , \41780 , \41790 );
xor \U$41796 ( \42173 , \42171 , \42172 );
nor \U$41797 ( \42174 , \42173 , \41982 );
buf \U$41798 ( \42175 , \42174 );
not \U$41799 ( \42176 , \7713 );
not \U$41800 ( \42177 , \42167 );
or \U$41801 ( \42178 , \42176 , \42177 );
nand \U$41802 ( \42179 , \42178 , \41783 );
nand \U$41803 ( \42180 , \41786 , \7857 );
xor \U$41804 ( \42181 , \42179 , \42180 );
nor \U$41805 ( \42182 , \42181 , \41982 );
buf \U$41806 ( \42183 , \42182 );
nand \U$41807 ( \42184 , \41783 , \7713 );
xnor \U$41808 ( \42185 , \42167 , \42184 );
not \U$41809 ( \42186 , \42185 );
nor \U$41810 ( \42187 , \42186 , \41982 );
buf \U$41811 ( \42188 , \42187 );
not \U$41812 ( \42189 , \8119 );
not \U$41813 ( \42190 , \8098 );
not \U$41814 ( \42191 , \42190 );
not \U$41815 ( \42192 , \42163 );
or \U$41816 ( \42193 , \42191 , \42192 );
and \U$41817 ( \42194 , \42147 , \42190 );
nor \U$41818 ( \42195 , \42194 , \41768 );
nand \U$41819 ( \42196 , \42193 , \42195 );
not \U$41820 ( \42197 , \42196 );
or \U$41821 ( \42198 , \42189 , \42197 );
nand \U$41822 ( \42199 , \42198 , \41772 );
not \U$41823 ( \42200 , \41775 );
nand \U$41824 ( \42201 , \42200 , \8126 );
xor \U$41825 ( \42202 , \42199 , \42201 );
nor \U$41826 ( \42203 , \42202 , \41982 );
buf \U$41827 ( \42204 , \42203 );
nand \U$41828 ( \42205 , \41772 , \8119 );
xor \U$41829 ( \42206 , \42196 , \42205 );
nor \U$41830 ( \42207 , \42206 , \41982 );
buf \U$41831 ( \42208 , \42207 );
not \U$41832 ( \42209 , \8097 );
not \U$41833 ( \42210 , \42149 );
or \U$41834 ( \42211 , \42209 , \42210 );
not \U$41835 ( \42212 , \41761 );
nand \U$41836 ( \42213 , \42211 , \42212 );
nand \U$41837 ( \42214 , \41767 , \8090 );
xor \U$41838 ( \42215 , \42213 , \42214 );
nor \U$41839 ( \42216 , \42215 , \41982 );
buf \U$41840 ( \42217 , \42216 );
nand \U$41841 ( \42218 , \42212 , \8097 );
xor \U$41842 ( \42219 , \42149 , \42218 );
nor \U$41843 ( \42220 , \42219 , \41982 );
buf \U$41844 ( \42221 , \42220 );
not \U$41845 ( \42222 , \4651 );
buf \U$41846 ( \42223 , \41739 );
nand \U$41847 ( \42224 , \42222 , \42223 );
not \U$41848 ( \42225 , \42224 );
nor \U$41849 ( \42226 , \6948 , \4651 );
nand \U$41850 ( \42227 , \41716 , \42226 );
not \U$41851 ( \42228 , \42227 );
or \U$41852 ( \42229 , \42225 , \42228 );
nand \U$41853 ( \42230 , \42229 , \5107 );
not \U$41854 ( \42231 , \41751 );
nand \U$41855 ( \42232 , \42230 , \42231 );
nand \U$41856 ( \42233 , \41754 , \5100 );
xor \U$41857 ( \42234 , \42232 , \42233 );
nor \U$41858 ( \42235 , \42234 , \41982 );
buf \U$41859 ( \42236 , \42235 );
not \U$41860 ( \42237 , \42226 );
not \U$41861 ( \42238 , \41716 );
or \U$41862 ( \42239 , \42237 , \42238 );
not \U$41863 ( \42240 , \42224 );
nor \U$41864 ( \42241 , \42240 , \41747 );
nand \U$41865 ( \42242 , \42239 , \42241 );
nand \U$41866 ( \42243 , \5107 , \41750 );
xor \U$41867 ( \42244 , \42242 , \42243 );
nor \U$41868 ( \42245 , \42244 , \41982 );
buf \U$41869 ( \42246 , \42245 );
not \U$41870 ( \42247 , \4650 );
not \U$41871 ( \42248 , \6948 );
not \U$41872 ( \42249 , \42248 );
not \U$41873 ( \42250 , \41716 );
or \U$41874 ( \42251 , \42249 , \42250 );
not \U$41875 ( \42252 , \42223 );
nand \U$41876 ( \42253 , \42251 , \42252 );
not \U$41877 ( \42254 , \42253 );
or \U$41878 ( \42255 , \42247 , \42254 );
nand \U$41879 ( \42256 , \42255 , \41744 );
not \U$41880 ( \42257 , \4273 );
nand \U$41881 ( \42258 , \42257 , \41746 );
xor \U$41882 ( \42259 , \42256 , \42258 );
nor \U$41883 ( \42260 , \42259 , \41982 );
buf \U$41884 ( \42261 , \42260 );
nand \U$41885 ( \42262 , \41744 , \4650 );
xor \U$41886 ( \42263 , \42253 , \42262 );
nor \U$41887 ( \42264 , \42263 , \41982 );
buf \U$41888 ( \42265 , \42264 );
not \U$41889 ( \42266 , \6940 );
not \U$41890 ( \42267 , \41716 );
or \U$41891 ( \42268 , \42266 , \42267 );
not \U$41892 ( \42269 , \41735 );
nand \U$41893 ( \42270 , \42268 , \42269 );
nand \U$41894 ( \42271 , \41738 , \6947 );
xor \U$41895 ( \42272 , \42270 , \42271 );
nor \U$41896 ( \42273 , \42272 , \41982 );
buf \U$41897 ( \42274 , \42273 );
not \U$41898 ( \42275 , \6939 );
not \U$41899 ( \42276 , \42275 );
not \U$41900 ( \42277 , \41716 );
or \U$41901 ( \42278 , \42276 , \42277 );
not \U$41902 ( \42279 , \41731 );
nand \U$41903 ( \42280 , \42278 , \42279 );
nand \U$41904 ( \42281 , \41734 , \5913 );
xor \U$41905 ( \42282 , \42280 , \42281 );
nor \U$41906 ( \42283 , \42282 , \41982 );
buf \U$41907 ( \42284 , \42283 );
not \U$41908 ( \42285 , \6938 );
not \U$41909 ( \42286 , \41716 );
or \U$41910 ( \42287 , \42285 , \42286 );
not \U$41911 ( \42288 , \41726 );
nand \U$41912 ( \42289 , \42287 , \42288 );
nand \U$41913 ( \42290 , \41730 , \6245 );
xor \U$41914 ( \42291 , \42289 , \42290 );
nor \U$41915 ( \42292 , \42291 , \41982 );
buf \U$41916 ( \42293 , \42292 );
not \U$41917 ( \42294 , \41981 );
nand \U$41918 ( \42295 , \42288 , \6938 );
xor \U$41919 ( \42296 , \42295 , \41716 );
nor \U$41920 ( \42297 , \42294 , \42296 );
buf \U$41921 ( \42298 , \42297 );
buf \U$41922 ( \42299 , \26496 );
and \U$41923 ( \42300 , \26551 , \26587 , \26602 );
and \U$41924 ( \42301 , \42299 , \42300 );
not \U$41925 ( \42302 , \42301 );
buf \U$41926 ( \42303 , \25824 );
not \U$41927 ( \42304 , \42303 );
not \U$41928 ( \42305 , \41697 );
not \U$41929 ( \42306 , \42305 );
buf \U$41930 ( \42307 , \41690 );
not \U$41931 ( \42308 , \42307 );
or \U$41932 ( \42309 , \42306 , \42308 );
buf \U$41933 ( \42310 , \22307 );
not \U$41934 ( \42311 , \42310 );
nand \U$41935 ( \42312 , \42309 , \42311 );
not \U$41936 ( \42313 , \42312 );
or \U$41937 ( \42314 , \42304 , \42313 );
buf \U$41938 ( \42315 , \26651 );
not \U$41939 ( \42316 , \42315 );
nand \U$41940 ( \42317 , \42314 , \42316 );
not \U$41941 ( \42318 , \42317 );
or \U$41942 ( \42319 , \42302 , \42318 );
not \U$41943 ( \42320 , \26668 );
and \U$41944 ( \42321 , \42320 , \42300 );
nor \U$41945 ( \42322 , \42321 , \41710 );
nand \U$41946 ( \42323 , \42319 , \42322 );
not \U$41947 ( \42324 , \41712 );
nand \U$41948 ( \42325 , \42324 , \26609 );
xor \U$41949 ( \42326 , \42323 , \42325 );
nor \U$41950 ( \42327 , \42326 , \41982 );
buf \U$41951 ( \42328 , \42327 );
not \U$41952 ( \42329 , \26551 );
nor \U$41953 ( \42330 , \42329 , \41703 );
not \U$41954 ( \42331 , \42330 );
and \U$41955 ( \42332 , \42303 , \42299 );
not \U$41956 ( \42333 , \42332 );
not \U$41957 ( \42334 , \42312 );
or \U$41958 ( \42335 , \42333 , \42334 );
not \U$41959 ( \42336 , \26669 );
nand \U$41960 ( \42337 , \42335 , \42336 );
not \U$41961 ( \42338 , \42337 );
or \U$41962 ( \42339 , \42331 , \42338 );
not \U$41963 ( \42340 , \41706 );
nand \U$41964 ( \42341 , \42339 , \42340 );
nand \U$41965 ( \42342 , \41709 , \26602 );
xor \U$41966 ( \42343 , \42341 , \42342 );
nor \U$41967 ( \42344 , \42343 , \41982 );
buf \U$41968 ( \42345 , \42344 );
not \U$41969 ( \42346 , \42337 );
not \U$41970 ( \42347 , \26551 );
or \U$41971 ( \42348 , \42346 , \42347 );
nand \U$41972 ( \42349 , \42348 , \41702 );
nand \U$41973 ( \42350 , \41705 , \26587 );
xor \U$41974 ( \42351 , \42349 , \42350 );
nor \U$41975 ( \42352 , \42351 , \41982 );
buf \U$41976 ( \42353 , \42352 );
nand \U$41977 ( \42354 , \41702 , \26551 );
xor \U$41978 ( \42355 , \42337 , \42354 );
nor \U$41979 ( \42356 , \42355 , \41982 );
buf \U$41980 ( \42357 , \42356 );
buf \U$41981 ( \42358 , \26304 );
buf \U$41982 ( \42359 , \26419 );
and \U$41983 ( \42360 , \42303 , \42358 , \42359 );
not \U$41984 ( \42361 , \42360 );
not \U$41985 ( \42362 , \42305 );
not \U$41986 ( \42363 , \42307 );
or \U$41987 ( \42364 , \42362 , \42363 );
not \U$41988 ( \42365 , \42310 );
nand \U$41989 ( \42366 , \42364 , \42365 );
not \U$41990 ( \42367 , \42366 );
or \U$41991 ( \42368 , \42361 , \42367 );
not \U$41992 ( \42369 , \42358 );
not \U$41993 ( \42370 , \42315 );
or \U$41994 ( \42371 , \42369 , \42370 );
not \U$41995 ( \42372 , \26660 );
nand \U$41996 ( \42373 , \42371 , \42372 );
and \U$41997 ( \42374 , \42373 , \42359 );
not \U$41998 ( \42375 , \26663 );
nor \U$41999 ( \42376 , \42374 , \42375 );
nand \U$42000 ( \42377 , \42368 , \42376 );
not \U$42001 ( \42378 , \26667 );
nand \U$42002 ( \42379 , \42378 , \26665 );
xor \U$42003 ( \42380 , \42377 , \42379 );
nor \U$42004 ( \42381 , \42380 , \41982 );
buf \U$42005 ( \42382 , \42381 );
not \U$42006 ( \42383 , \42358 );
not \U$42007 ( \42384 , \42317 );
or \U$42008 ( \42385 , \42383 , \42384 );
nand \U$42009 ( \42386 , \42385 , \42372 );
nand \U$42010 ( \42387 , \26663 , \42359 );
xor \U$42011 ( \42388 , \42386 , \42387 );
nor \U$42012 ( \42389 , \42388 , \41982 );
buf \U$42013 ( \42390 , \42389 );
buf \U$42014 ( \42391 , \26303 );
not \U$42015 ( \42392 , \42391 );
not \U$42016 ( \42393 , \42317 );
or \U$42017 ( \42394 , \42392 , \42393 );
not \U$42018 ( \42395 , \26656 );
nand \U$42019 ( \42396 , \42394 , \42395 );
nand \U$42020 ( \42397 , \26296 , \26659 );
xor \U$42021 ( \42398 , \42396 , \42397 );
nor \U$42022 ( \42399 , \42398 , \41982 );
buf \U$42023 ( \42400 , \42399 );
not \U$42024 ( \42401 , \42317 );
nand \U$42025 ( \42402 , \42395 , \42391 );
not \U$42026 ( \42403 , \42402 );
or \U$42027 ( \42404 , \42401 , \42403 );
or \U$42028 ( \42405 , \42402 , \42317 );
nand \U$42029 ( \42406 , \42404 , \42405 );
and \U$42030 ( \42407 , \42406 , \41981 );
buf \U$42031 ( \42408 , \42407 );
not \U$42032 ( \42409 , \25014 );
buf \U$42033 ( \42410 , \25430 );
and \U$42034 ( \42411 , \42409 , \42410 );
not \U$42035 ( \42412 , \42411 );
buf \U$42036 ( \42413 , \24153 );
and \U$42037 ( \42414 , \42366 , \42413 );
not \U$42038 ( \42415 , \42414 );
or \U$42039 ( \42416 , \42412 , \42415 );
not \U$42040 ( \42417 , \42409 );
buf \U$42041 ( \42418 , \26632 );
not \U$42042 ( \42419 , \42418 );
or \U$42043 ( \42420 , \42417 , \42419 );
not \U$42044 ( \42421 , \26642 );
nand \U$42045 ( \42422 , \42420 , \42421 );
and \U$42046 ( \42423 , \42422 , \42410 );
not \U$42047 ( \42424 , \26645 );
nor \U$42048 ( \42425 , \42423 , \42424 );
nand \U$42049 ( \42426 , \42416 , \42425 );
not \U$42050 ( \42427 , \26649 );
nand \U$42051 ( \42428 , \42427 , \26647 );
xor \U$42052 ( \42429 , \42426 , \42428 );
nor \U$42053 ( \42430 , \42429 , \41982 );
buf \U$42054 ( \42431 , \42430 );
not \U$42055 ( \42432 , \42409 );
not \U$42056 ( \42433 , \42413 );
not \U$42057 ( \42434 , \42312 );
or \U$42058 ( \42435 , \42433 , \42434 );
not \U$42059 ( \42436 , \42418 );
nand \U$42060 ( \42437 , \42435 , \42436 );
not \U$42061 ( \42438 , \42437 );
or \U$42062 ( \42439 , \42432 , \42438 );
nand \U$42063 ( \42440 , \42439 , \42421 );
nand \U$42064 ( \42441 , \42410 , \26645 );
xor \U$42065 ( \42442 , \42440 , \42441 );
nor \U$42066 ( \42443 , \42442 , \41982 );
buf \U$42067 ( \42444 , \42443 );
not \U$42068 ( \42445 , \25013 );
not \U$42069 ( \42446 , \42437 );
or \U$42070 ( \42447 , \42445 , \42446 );
buf \U$42071 ( \42448 , \26638 );
nand \U$42072 ( \42449 , \42447 , \42448 );
not \U$42073 ( \42450 , \26637 );
nand \U$42074 ( \42451 , \42450 , \26641 );
xor \U$42075 ( \42452 , \42449 , \42451 );
nor \U$42076 ( \42453 , \42452 , \41982 );
buf \U$42077 ( \42454 , \42453 );
not \U$42078 ( \42455 , \42437 );
nand \U$42079 ( \42456 , \42448 , \25013 );
not \U$42080 ( \42457 , \42456 );
or \U$42081 ( \42458 , \42455 , \42457 );
or \U$42082 ( \42459 , \42456 , \42437 );
nand \U$42083 ( \42460 , \42458 , \42459 );
and \U$42084 ( \42461 , \42460 , \41981 );
buf \U$42085 ( \42462 , \42461 );
and \U$42086 ( \42463 , \24128 , \24152 );
nand \U$42087 ( \42464 , \42366 , \42463 );
not \U$42088 ( \42465 , \24135 );
or \U$42089 ( \42466 , \42464 , \42465 );
not \U$42090 ( \42467 , \26628 );
nand \U$42091 ( \42468 , \42466 , \42467 );
nand \U$42092 ( \42469 , \24070 , \26631 );
xor \U$42093 ( \42470 , \42468 , \42469 );
nor \U$42094 ( \42471 , \42470 , \41982 );
buf \U$42095 ( \42472 , \42471 );
not \U$42096 ( \42473 , \26624 );
nand \U$42097 ( \42474 , \42464 , \42473 );
nand \U$42098 ( \42475 , \26627 , \24135 );
xor \U$42099 ( \42476 , \42474 , \42475 );
nor \U$42100 ( \42477 , \42476 , \41982 );
buf \U$42101 ( \42478 , \42477 );
nand \U$42102 ( \42479 , \26623 , \24128 );
not \U$42103 ( \42480 , \24152 );
not \U$42104 ( \42481 , \42366 );
or \U$42105 ( \42482 , \42480 , \42481 );
buf \U$42106 ( \42483 , \26618 );
nand \U$42107 ( \42484 , \42482 , \42483 );
xor \U$42108 ( \42485 , \42479 , \42484 );
nor \U$42109 ( \42486 , \42485 , \41982 );
buf \U$42110 ( \42487 , \42486 );
not \U$42111 ( \42488 , \42366 );
nand \U$42112 ( \42489 , \42483 , \24152 );
not \U$42113 ( \42490 , \42489 );
or \U$42114 ( \42491 , \42488 , \42490 );
or \U$42115 ( \42492 , \42489 , \42366 );
nand \U$42116 ( \42493 , \42491 , \42492 );
and \U$42117 ( \42494 , \42493 , \41981 );
buf \U$42118 ( \42495 , \42494 );
not \U$42119 ( \42496 , \15098 );
nor \U$42120 ( \42497 , \17457 , \14093 );
not \U$42121 ( \42498 , \42497 );
buf \U$42122 ( \42499 , \22262 );
and \U$42123 ( \42500 , \22263 , \42499 );
buf \U$42124 ( \42501 , \18889 );
and \U$42125 ( \42502 , \41696 , \42500 , \20024 , \42501 );
not \U$42126 ( \42503 , \42502 );
not \U$42127 ( \42504 , \42307 );
or \U$42128 ( \42505 , \42503 , \42504 );
not \U$42129 ( \42506 , \22266 );
nand \U$42130 ( \42507 , \42505 , \42506 );
not \U$42131 ( \42508 , \42507 );
or \U$42132 ( \42509 , \42498 , \42508 );
buf \U$42133 ( \42510 , \22285 );
not \U$42134 ( \42511 , \14093 );
and \U$42135 ( \42512 , \42510 , \42511 );
nor \U$42136 ( \42513 , \42512 , \22295 );
nand \U$42137 ( \42514 , \42509 , \42513 );
not \U$42138 ( \42515 , \42514 );
or \U$42139 ( \42516 , \42496 , \42515 );
nand \U$42140 ( \42517 , \42516 , \22299 );
not \U$42141 ( \42518 , \22303 );
nand \U$42142 ( \42519 , \42518 , \22301 );
xor \U$42143 ( \42520 , \42517 , \42519 );
nor \U$42144 ( \42521 , \42520 , \41982 );
buf \U$42145 ( \42522 , \42521 );
nand \U$42146 ( \42523 , \15098 , \22299 );
xor \U$42147 ( \42524 , \42514 , \42523 );
nor \U$42148 ( \42525 , \42524 , \41982 );
buf \U$42149 ( \42526 , \42525 );
not \U$42150 ( \42527 , \13561 );
not \U$42151 ( \42528 , \41692 );
not \U$42152 ( \42529 , \42507 );
or \U$42153 ( \42530 , \42528 , \42529 );
not \U$42154 ( \42531 , \42510 );
nand \U$42155 ( \42532 , \42530 , \42531 );
not \U$42156 ( \42533 , \42532 );
or \U$42157 ( \42534 , \42527 , \42533 );
buf \U$42158 ( \42535 , \22290 );
nand \U$42159 ( \42536 , \42534 , \42535 );
nand \U$42160 ( \42537 , \22294 , \14092 );
xor \U$42161 ( \42538 , \42536 , \42537 );
nor \U$42162 ( \42539 , \42538 , \41982 );
buf \U$42163 ( \42540 , \42539 );
nand \U$42164 ( \42541 , \42535 , \13561 );
xor \U$42165 ( \42542 , \42532 , \42541 );
nor \U$42166 ( \42543 , \42542 , \41982 );
buf \U$42167 ( \42544 , \42543 );
nand \U$42168 ( \42545 , \17445 , \16740 );
nor \U$42169 ( \42546 , \42545 , \16194 );
not \U$42170 ( \42547 , \42546 );
buf \U$42171 ( \42548 , \42507 );
not \U$42172 ( \42549 , \42548 );
or \U$42173 ( \42550 , \42547 , \42549 );
not \U$42174 ( \42551 , \22279 );
nand \U$42175 ( \42552 , \42550 , \42551 );
nand \U$42176 ( \42553 , \17456 , \22284 );
xor \U$42177 ( \42554 , \42552 , \42553 );
nor \U$42178 ( \42555 , \42554 , \41982 );
buf \U$42179 ( \42556 , \42555 );
not \U$42180 ( \42557 , \42545 );
not \U$42181 ( \42558 , \42557 );
not \U$42182 ( \42559 , \42548 );
or \U$42183 ( \42560 , \42558 , \42559 );
buf \U$42184 ( \42561 , \22276 );
nand \U$42185 ( \42562 , \42560 , \42561 );
not \U$42186 ( \42563 , \16194 );
nand \U$42187 ( \42564 , \42563 , \22278 );
xor \U$42188 ( \42565 , \42562 , \42564 );
nor \U$42189 ( \42566 , \42565 , \41982 );
buf \U$42190 ( \42567 , \42566 );
not \U$42191 ( \42568 , \17445 );
not \U$42192 ( \42569 , \42548 );
or \U$42193 ( \42570 , \42568 , \42569 );
buf \U$42194 ( \42571 , \22274 );
nand \U$42195 ( \42572 , \42570 , \42571 );
not \U$42196 ( \42573 , \16737 );
not \U$42197 ( \42574 , \16197 );
or \U$42198 ( \42575 , \42573 , \42574 );
nand \U$42199 ( \42576 , \42575 , \16740 );
xor \U$42200 ( \42577 , \42572 , \42576 );
nor \U$42201 ( \42578 , \42577 , \41982 );
buf \U$42202 ( \42579 , \42578 );
nand \U$42203 ( \42580 , \42571 , \17445 );
not \U$42204 ( \42581 , \42580 );
not \U$42205 ( \42582 , \42548 );
or \U$42206 ( \42583 , \42581 , \42582 );
or \U$42207 ( \42584 , \42548 , \42580 );
nand \U$42208 ( \42585 , \42583 , \42584 );
and \U$42209 ( \42586 , \42585 , \41981 );
buf \U$42210 ( \42587 , \42586 );
and \U$42211 ( \42588 , \42500 , \42501 );
not \U$42212 ( \42589 , \42588 );
not \U$42213 ( \42590 , \41696 );
not \U$42214 ( \42591 , \42307 );
or \U$42215 ( \42592 , \42590 , \42591 );
not \U$42216 ( \42593 , \22261 );
nand \U$42217 ( \42594 , \42592 , \42593 );
not \U$42218 ( \42595 , \42594 );
or \U$42219 ( \42596 , \42589 , \42595 );
not \U$42220 ( \42597 , \20014 );
nand \U$42221 ( \42598 , \42596 , \42597 );
not \U$42222 ( \42599 , \20026 );
nand \U$42223 ( \42600 , \42599 , \20024 );
xor \U$42224 ( \42601 , \42598 , \42600 );
nor \U$42225 ( \42602 , \42601 , \41982 );
buf \U$42226 ( \42603 , \42602 );
not \U$42227 ( \42604 , \42500 );
not \U$42228 ( \42605 , \42594 );
or \U$42229 ( \42606 , \42604 , \42605 );
not \U$42230 ( \42607 , \20010 );
nand \U$42231 ( \42608 , \42606 , \42607 );
nand \U$42232 ( \42609 , \20013 , \42501 );
xor \U$42233 ( \42610 , \42608 , \42609 );
nor \U$42234 ( \42611 , \42610 , \41982 );
buf \U$42235 ( \42612 , \42611 );
not \U$42236 ( \42613 , \22263 );
not \U$42237 ( \42614 , \42594 );
or \U$42238 ( \42615 , \42613 , \42614 );
not \U$42239 ( \42616 , \19996 );
nand \U$42240 ( \42617 , \42615 , \42616 );
nand \U$42241 ( \42618 , \20009 , \42499 );
xor \U$42242 ( \42619 , \42617 , \42618 );
nor \U$42243 ( \42620 , \42619 , \41982 );
buf \U$42244 ( \42621 , \42620 );
not \U$42245 ( \42622 , \42594 );
nand \U$42246 ( \42623 , \22263 , \42616 );
not \U$42247 ( \42624 , \42623 );
or \U$42248 ( \42625 , \42622 , \42624 );
or \U$42249 ( \42626 , \42623 , \42594 );
nand \U$42250 ( \42627 , \42625 , \42626 );
and \U$42251 ( \42628 , \42627 , \41981 );
buf \U$42252 ( \42629 , \42628 );
not \U$42253 ( \42630 , \41694 );
buf \U$42254 ( \42631 , \41695 );
and \U$42255 ( \42632 , \41693 , \42631 );
not \U$42256 ( \42633 , \42632 );
buf \U$42257 ( \42634 , \42307 );
not \U$42258 ( \42635 , \42634 );
or \U$42259 ( \42636 , \42633 , \42635 );
buf \U$42260 ( \42637 , \22244 );
nand \U$42261 ( \42638 , \42636 , \42637 );
not \U$42262 ( \42639 , \42638 );
or \U$42263 ( \42640 , \42630 , \42639 );
buf \U$42264 ( \42641 , \22254 );
nand \U$42265 ( \42642 , \42640 , \42641 );
nand \U$42266 ( \42643 , \22260 , \20831 );
xor \U$42267 ( \42644 , \42642 , \42643 );
nor \U$42268 ( \42645 , \42644 , \41982 );
buf \U$42269 ( \42646 , \42645 );
nand \U$42270 ( \42647 , \42641 , \41694 );
xor \U$42271 ( \42648 , \42638 , \42647 );
not \U$42272 ( \42649 , \41980 );
nor \U$42273 ( \42650 , \42648 , \42649 );
buf \U$42274 ( \42651 , \42650 );
not \U$42275 ( \42652 , \42631 );
not \U$42276 ( \42653 , \42307 );
or \U$42277 ( \42654 , \42652 , \42653 );
buf \U$42278 ( \42655 , \22239 );
nand \U$42279 ( \42656 , \42654 , \42655 );
not \U$42280 ( \42657 , \22242 );
not \U$42281 ( \42658 , \42657 );
not \U$42282 ( \42659 , \21811 );
or \U$42283 ( \42660 , \42658 , \42659 );
nand \U$42284 ( \42661 , \42660 , \41693 );
xor \U$42285 ( \42662 , \42656 , \42661 );
nor \U$42286 ( \42663 , \42662 , \41982 );
buf \U$42287 ( \42664 , \42663 );
not \U$42288 ( \42665 , \42307 );
nand \U$42289 ( \42666 , \42655 , \42631 );
not \U$42290 ( \42667 , \42666 );
or \U$42291 ( \42668 , \42665 , \42667 );
or \U$42292 ( \42669 , \42634 , \42666 );
nand \U$42293 ( \42670 , \42668 , \42669 );
and \U$42294 ( \42671 , \42670 , \41979 );
buf \U$42295 ( \42672 , \42671 );
not \U$42296 ( \42673 , RIc2275b0_1);
nor \U$42297 ( \42674 , \42673 , \41980 );
not \U$42298 ( \42675 , \42674 );
nand \U$42299 ( \42676 , \33971 , \41688 );
not \U$42300 ( \42677 , \42676 );
not \U$42301 ( \42678 , \33957 );
and \U$42302 ( \42679 , \33964 , \33886 );
not \U$42303 ( \42680 , \42679 );
not \U$42304 ( \42681 , \33795 );
nand \U$42305 ( \42682 , \38412 , \41675 );
not \U$42306 ( \42683 , \42682 );
not \U$42307 ( \42684 , \38420 );
or \U$42308 ( \42685 , \42683 , \42684 );
and \U$42309 ( \42686 , \31207 , \32906 );
nand \U$42310 ( \42687 , \42685 , \42686 );
nand \U$42311 ( \42688 , \42681 , \42687 );
not \U$42312 ( \42689 , \33811 );
nand \U$42313 ( \42690 , \42688 , \42689 );
not \U$42314 ( \42691 , \42690 );
or \U$42315 ( \42692 , \42680 , \42691 );
not \U$42316 ( \42693 , \41683 );
nand \U$42317 ( \42694 , \42692 , \42693 );
not \U$42318 ( \42695 , \42694 );
or \U$42319 ( \42696 , \42678 , \42695 );
not \U$42320 ( \42697 , \41684 );
nand \U$42321 ( \42698 , \42696 , \42697 );
not \U$42322 ( \42699 , \42698 );
or \U$42323 ( \42700 , \42677 , \42699 );
or \U$42324 ( \42701 , \42698 , \42676 );
nand \U$42325 ( \42702 , \42700 , \42701 );
nand \U$42326 ( \42703 , \42702 , \41981 );
nand \U$42327 ( \42704 , \42675 , \42703 );
buf \U$42328 ( \42705 , \42704 );
not \U$42329 ( \42706 , RIc227538_2);
nor \U$42330 ( \42707 , \42706 , \41979 );
not \U$42331 ( \42708 , \42707 );
nand \U$42332 ( \42709 , \42697 , \33957 );
not \U$42333 ( \42710 , \42709 );
not \U$42334 ( \42711 , \42694 );
or \U$42335 ( \42712 , \42710 , \42711 );
or \U$42336 ( \42713 , \42694 , \42709 );
nand \U$42337 ( \42714 , \42712 , \42713 );
nand \U$42338 ( \42715 , \42714 , \41981 );
nand \U$42339 ( \42716 , \42708 , \42715 );
buf \U$42340 ( \42717 , \42716 );
not \U$42341 ( \42718 , RIc2274c0_3);
nor \U$42342 ( \42719 , \42718 , \41979 );
not \U$42343 ( \42720 , \42719 );
nand \U$42344 ( \42721 , \41682 , \33964 );
not \U$42345 ( \42722 , \42721 );
not \U$42346 ( \42723 , \33886 );
not \U$42347 ( \42724 , \42690 );
or \U$42348 ( \42725 , \42723 , \42724 );
not \U$42349 ( \42726 , \41678 );
nand \U$42350 ( \42727 , \42725 , \42726 );
not \U$42351 ( \42728 , \42727 );
or \U$42352 ( \42729 , \42722 , \42728 );
or \U$42353 ( \42730 , \42727 , \42721 );
nand \U$42354 ( \42731 , \42729 , \42730 );
nand \U$42355 ( \42732 , \42731 , \41981 );
nand \U$42356 ( \42733 , \42720 , \42732 );
buf \U$42357 ( \42734 , \42733 );
not \U$42358 ( \42735 , RIc227448_4);
nor \U$42359 ( \42736 , \42735 , \41979 );
not \U$42360 ( \42737 , \42736 );
nand \U$42361 ( \42738 , \33886 , \42726 );
not \U$42362 ( \42739 , \42738 );
not \U$42363 ( \42740 , \42690 );
or \U$42364 ( \42741 , \42739 , \42740 );
or \U$42365 ( \42742 , \42738 , \42690 );
nand \U$42366 ( \42743 , \42741 , \42742 );
nand \U$42367 ( \42744 , \42743 , \41980 );
nand \U$42368 ( \42745 , \42737 , \42744 );
buf \U$42369 ( \42746 , \42745 );
not \U$42370 ( \42747 , RIc2273d0_5);
nor \U$42371 ( \42748 , \42747 , \41980 );
not \U$42372 ( \42749 , \42748 );
not \U$42373 ( \42750 , \33669 );
buf \U$42374 ( \42751 , \33499 );
buf \U$42375 ( \42752 , \33793 );
and \U$42376 ( \42753 , \42751 , \42752 );
not \U$42377 ( \42754 , \42753 );
not \U$42378 ( \42755 , \42687 );
or \U$42379 ( \42756 , \42754 , \42755 );
nand \U$42380 ( \42757 , \42756 , \33803 );
not \U$42381 ( \42758 , \42757 );
or \U$42382 ( \42759 , \42750 , \42758 );
nand \U$42383 ( \42760 , \42759 , \33806 );
nand \U$42384 ( \42761 , \33810 , \33781 );
not \U$42385 ( \42762 , \42761 );
and \U$42386 ( \42763 , \42760 , \42762 );
not \U$42387 ( \42764 , \42760 );
and \U$42388 ( \42765 , \42764 , \42761 );
nor \U$42389 ( \42766 , \42763 , \42765 );
nand \U$42390 ( \42767 , \42766 , \41981 );
nand \U$42391 ( \42768 , \42749 , \42767 );
buf \U$42392 ( \42769 , \42768 );
not \U$42393 ( \42770 , RIc227358_6);
nor \U$42394 ( \42771 , \42770 , \41979 );
not \U$42395 ( \42772 , \42771 );
not \U$42396 ( \42773 , \33804 );
nand \U$42397 ( \42774 , \42773 , \33806 );
not \U$42398 ( \42775 , \42774 );
and \U$42399 ( \42776 , \42757 , \42775 );
not \U$42400 ( \42777 , \42757 );
and \U$42401 ( \42778 , \42777 , \42774 );
nor \U$42402 ( \42779 , \42776 , \42778 );
nand \U$42403 ( \42780 , \42779 , \41980 );
nand \U$42404 ( \42781 , \42772 , \42780 );
buf \U$42405 ( \42782 , \42781 );
not \U$42406 ( \42783 , RIc2272e0_7);
nor \U$42407 ( \42784 , \42783 , \41979 );
not \U$42408 ( \42785 , \42784 );
not \U$42409 ( \42786 , \42752 );
not \U$42410 ( \42787 , \42687 );
or \U$42411 ( \42788 , \42786 , \42787 );
nand \U$42412 ( \42789 , \42788 , \33801 );
not \U$42413 ( \42790 , \33497 );
not \U$42414 ( \42791 , \33465 );
or \U$42415 ( \42792 , \42790 , \42791 );
nand \U$42416 ( \42793 , \42792 , \42751 );
not \U$42417 ( \42794 , \42793 );
and \U$42418 ( \42795 , \42789 , \42794 );
not \U$42419 ( \42796 , \42789 );
and \U$42420 ( \42797 , \42796 , \42793 );
nor \U$42421 ( \42798 , \42795 , \42797 );
nand \U$42422 ( \42799 , \42798 , \41979 );
nand \U$42423 ( \42800 , \42785 , \42799 );
buf \U$42424 ( \42801 , \42800 );
not \U$42425 ( \42802 , \41979 );
nand \U$42426 ( \42803 , \33801 , \42752 );
xnor \U$42427 ( \42804 , \42803 , \42687 );
not \U$42428 ( \42805 , \42804 );
or \U$42429 ( \42806 , \42802 , \42805 );
nand \U$42430 ( \42807 , \41978 , RIc227268_8);
nand \U$42431 ( \42808 , \42806 , \42807 );
buf \U$42432 ( \42809 , \42808 );
not \U$42433 ( \42810 , RIc2271f0_9);
nor \U$42434 ( \42811 , \42810 , \41979 );
not \U$42435 ( \42812 , \42811 );
nand \U$42436 ( \42813 , \31205 , \30140 );
not \U$42437 ( \42814 , \42813 );
buf \U$42438 ( \42815 , \30537 );
not \U$42439 ( \42816 , \42815 );
buf \U$42440 ( \42817 , \31193 );
and \U$42441 ( \42818 , \32903 , \42817 );
not \U$42442 ( \42819 , \42818 );
nor \U$42443 ( \42820 , \38414 , \38418 );
not \U$42444 ( \42821 , \42820 );
not \U$42445 ( \42822 , \42682 );
or \U$42446 ( \42823 , \42821 , \42822 );
not \U$42447 ( \42824 , \32902 );
nand \U$42448 ( \42825 , \42823 , \42824 );
not \U$42449 ( \42826 , \42825 );
or \U$42450 ( \42827 , \42819 , \42826 );
not \U$42451 ( \42828 , \31196 );
nand \U$42452 ( \42829 , \42827 , \42828 );
not \U$42453 ( \42830 , \42829 );
or \U$42454 ( \42831 , \42816 , \42830 );
nand \U$42455 ( \42832 , \42831 , \31201 );
not \U$42456 ( \42833 , \42832 );
or \U$42457 ( \42834 , \42814 , \42833 );
or \U$42458 ( \42835 , \42832 , \42813 );
nand \U$42459 ( \42836 , \42834 , \42835 );
nand \U$42460 ( \42837 , \42836 , \41981 );
nand \U$42461 ( \42838 , \42812 , \42837 );
buf \U$42462 ( \42839 , \42838 );
not \U$42463 ( \42840 , RIc227178_10);
nor \U$42464 ( \42841 , \42840 , \41979 );
not \U$42465 ( \42842 , \42841 );
nand \U$42466 ( \42843 , \31201 , \42815 );
not \U$42467 ( \42844 , \42843 );
not \U$42468 ( \42845 , \42829 );
or \U$42469 ( \42846 , \42844 , \42845 );
or \U$42470 ( \42847 , \42829 , \42843 );
nand \U$42471 ( \42848 , \42846 , \42847 );
nand \U$42472 ( \42849 , \41980 , \42848 );
nand \U$42473 ( \42850 , \42842 , \42849 );
buf \U$42474 ( \42851 , \42850 );
not \U$42475 ( \42852 , RIc227100_11);
nor \U$42476 ( \42853 , \42852 , \41979 );
not \U$42477 ( \42854 , \42853 );
not \U$42478 ( \42855 , \32903 );
not \U$42479 ( \42856 , \42825 );
or \U$42480 ( \42857 , \42855 , \42856 );
not \U$42481 ( \42858 , \31186 );
nand \U$42482 ( \42859 , \42857 , \42858 );
nand \U$42483 ( \42860 , \31195 , \42817 );
not \U$42484 ( \42861 , \42860 );
and \U$42485 ( \42862 , \42859 , \42861 );
not \U$42486 ( \42863 , \42859 );
and \U$42487 ( \42864 , \42863 , \42860 );
nor \U$42488 ( \42865 , \42862 , \42864 );
nand \U$42489 ( \42866 , \42865 , \41980 );
nand \U$42490 ( \42867 , \42854 , \42866 );
buf \U$42491 ( \42868 , \42867 );
not \U$42492 ( \42869 , \41979 );
nand \U$42493 ( \42870 , \32903 , \42858 );
not \U$42494 ( \42871 , \42870 );
not \U$42495 ( \42872 , \42825 );
or \U$42496 ( \42873 , \42871 , \42872 );
or \U$42497 ( \42874 , \42870 , \42825 );
nand \U$42498 ( \42875 , \42873 , \42874 );
not \U$42499 ( \42876 , \42875 );
or \U$42500 ( \42877 , \42869 , \42876 );
nand \U$42501 ( \42878 , \41978 , RIc227088_12);
nand \U$42502 ( \42879 , \42877 , \42878 );
buf \U$42503 ( \42880 , \42879 );
not \U$42504 ( \42881 , RIc227010_13);
nor \U$42505 ( \42882 , \42881 , \41979 );
not \U$42506 ( \42883 , \42882 );
not \U$42507 ( \42884 , \32887 );
not \U$42508 ( \42885 , \42884 );
not \U$42509 ( \42886 , \38418 );
not \U$42510 ( \42887 , \42886 );
not \U$42511 ( \42888 , \42682 );
or \U$42512 ( \42889 , \42887 , \42888 );
nand \U$42513 ( \42890 , \42889 , \32859 );
not \U$42514 ( \42891 , \42890 );
or \U$42515 ( \42892 , \42885 , \42891 );
nand \U$42516 ( \42893 , \42892 , \32896 );
nand \U$42517 ( \42894 , \32895 , \32901 );
not \U$42518 ( \42895 , \42894 );
and \U$42519 ( \42896 , \42893 , \42895 );
not \U$42520 ( \42897 , \42893 );
and \U$42521 ( \42898 , \42897 , \42894 );
nor \U$42522 ( \42899 , \42896 , \42898 );
nand \U$42523 ( \42900 , \42899 , \41979 );
nand \U$42524 ( \42901 , \42883 , \42900 );
buf \U$42525 ( \42902 , \42901 );
not \U$42526 ( \42903 , \41979 );
nand \U$42527 ( \42904 , \32896 , \42884 );
not \U$42528 ( \42905 , \42904 );
not \U$42529 ( \42906 , \42890 );
or \U$42530 ( \42907 , \42905 , \42906 );
or \U$42531 ( \42908 , \42904 , \42890 );
nand \U$42532 ( \42909 , \42907 , \42908 );
not \U$42533 ( \42910 , \42909 );
or \U$42534 ( \42911 , \42903 , \42910 );
nand \U$42535 ( \42912 , \41978 , RIc226f98_14);
nand \U$42536 ( \42913 , \42911 , \42912 );
buf \U$42537 ( \42914 , \42913 );
not \U$42538 ( \42915 , \41979 );
not \U$42539 ( \42916 , \32283 );
not \U$42540 ( \42917 , \32313 );
or \U$42541 ( \42918 , \42916 , \42917 );
nand \U$42542 ( \42919 , \42918 , \32858 );
not \U$42543 ( \42920 , \42919 );
buf \U$42544 ( \42921 , \38417 );
not \U$42545 ( \42922 , \42921 );
not \U$42546 ( \42923 , \42682 );
or \U$42547 ( \42924 , \42922 , \42923 );
nand \U$42548 ( \42925 , \42924 , \32854 );
not \U$42549 ( \42926 , \42925 );
or \U$42550 ( \42927 , \42920 , \42926 );
or \U$42551 ( \42928 , \42925 , \42919 );
nand \U$42552 ( \42929 , \42927 , \42928 );
not \U$42553 ( \42930 , \42929 );
or \U$42554 ( \42931 , \42915 , \42930 );
nand \U$42555 ( \42932 , \41978 , RIc226f20_15);
nand \U$42556 ( \42933 , \42931 , \42932 );
buf \U$42557 ( \42934 , \42933 );
and \U$42558 ( \42935 , \41978 , RIc226ea8_16);
not \U$42559 ( \42936 , \41978 );
nand \U$42560 ( \42937 , \32854 , \42921 );
xnor \U$42561 ( \42938 , \42682 , \42937 );
and \U$42562 ( \42939 , \42936 , \42938 );
or \U$42563 ( \42940 , \42935 , \42939 );
buf \U$42564 ( \42941 , \42940 );
not \U$42565 ( \42942 , RIc226e30_17);
nor \U$42566 ( \42943 , \42942 , \41979 );
not \U$42567 ( \42944 , \42943 );
nand \U$42568 ( \42945 , \41673 , \41658 );
not \U$42569 ( \42946 , \42945 );
not \U$42570 ( \42947 , \38372 );
buf \U$42571 ( \42948 , \38395 );
buf \U$42572 ( \42949 , \38409 );
and \U$42573 ( \42950 , \42948 , \42949 );
not \U$42574 ( \42951 , \42950 );
not \U$42575 ( \42952 , \38278 );
not \U$42576 ( \42953 , \38430 );
not \U$42577 ( \42954 , \41656 );
or \U$42578 ( \42955 , \42953 , \42954 );
nand \U$42579 ( \42956 , \42955 , \37685 );
not \U$42580 ( \42957 , \42956 );
or \U$42581 ( \42958 , \42952 , \42957 );
not \U$42582 ( \42959 , \38296 );
nand \U$42583 ( \42960 , \42958 , \42959 );
not \U$42584 ( \42961 , \42960 );
or \U$42585 ( \42962 , \42951 , \42961 );
not \U$42586 ( \42963 , \41666 );
nand \U$42587 ( \42964 , \42962 , \42963 );
not \U$42588 ( \42965 , \42964 );
or \U$42589 ( \42966 , \42947 , \42965 );
nand \U$42590 ( \42967 , \42966 , \41669 );
not \U$42591 ( \42968 , \42967 );
or \U$42592 ( \42969 , \42946 , \42968 );
or \U$42593 ( \42970 , \42967 , \42945 );
nand \U$42594 ( \42971 , \42969 , \42970 );
nand \U$42595 ( \42972 , \42971 , \41979 );
nand \U$42596 ( \42973 , \42944 , \42972 );
buf \U$42597 ( \42974 , \42973 );
nand \U$42598 ( \42975 , \41669 , \38372 );
not \U$42599 ( \42976 , \42975 );
not \U$42600 ( \42977 , \42964 );
or \U$42601 ( \42978 , \42976 , \42977 );
or \U$42602 ( \42979 , \42964 , \42975 );
nand \U$42603 ( \42980 , \42978 , \42979 );
and \U$42604 ( \42981 , \41979 , \42980 );
not \U$42605 ( \42982 , \41979 );
and \U$42606 ( \42983 , \42982 , RIc226db8_18);
or \U$42607 ( \42984 , \42981 , \42983 );
buf \U$42608 ( \42985 , \42984 );
buf \U$42609 ( \42986 , \41665 );
nand \U$42610 ( \42987 , \42986 , \42948 );
not \U$42611 ( \42988 , \42987 );
not \U$42612 ( \42989 , \42949 );
not \U$42613 ( \42990 , \42960 );
or \U$42614 ( \42991 , \42989 , \42990 );
not \U$42615 ( \42992 , \41661 );
nand \U$42616 ( \42993 , \42991 , \42992 );
not \U$42617 ( \42994 , \42993 );
or \U$42618 ( \42995 , \42988 , \42994 );
or \U$42619 ( \42996 , \42993 , \42987 );
nand \U$42620 ( \42997 , \42995 , \42996 );
and \U$42621 ( \42998 , \41979 , \42997 );
not \U$42622 ( \42999 , \41979 );
and \U$42623 ( \43000 , \42999 , RIc226d40_19);
or \U$42624 ( \43001 , \42998 , \43000 );
buf \U$42625 ( \43002 , \43001 );
nand \U$42626 ( \43003 , \42992 , \42949 );
xnor \U$42627 ( \43004 , \42960 , \43003 );
and \U$42628 ( \43005 , \41979 , \43004 );
not \U$42629 ( \43006 , \41979 );
and \U$42630 ( \43007 , \43006 , RIc226cc8_20);
or \U$42631 ( \43008 , \43005 , \43007 );
buf \U$42632 ( \43009 , \43008 );
nand \U$42633 ( \43010 , \38292 , \38277 );
not \U$42634 ( \43011 , \43010 );
not \U$42635 ( \43012 , \38175 );
buf \U$42636 ( \43013 , \38185 );
and \U$42637 ( \43014 , \38071 , \43013 );
not \U$42638 ( \43015 , \43014 );
not \U$42639 ( \43016 , \42956 );
or \U$42640 ( \43017 , \43015 , \43016 );
not \U$42641 ( \43018 , \38285 );
nand \U$42642 ( \43019 , \43017 , \43018 );
not \U$42643 ( \43020 , \43019 );
or \U$42644 ( \43021 , \43012 , \43020 );
nand \U$42645 ( \43022 , \43021 , \38289 );
not \U$42646 ( \43023 , \43022 );
or \U$42647 ( \43024 , \43011 , \43023 );
or \U$42648 ( \43025 , \43022 , \43010 );
nand \U$42649 ( \43026 , \43024 , \43025 );
and \U$42650 ( \43027 , \41979 , \43026 );
not \U$42651 ( \43028 , \41979 );
and \U$42652 ( \43029 , \43028 , RIc226c50_21);
or \U$42653 ( \43030 , \43027 , \43029 );
buf \U$42654 ( \43031 , \43030 );
nand \U$42655 ( \43032 , \38289 , \38175 );
not \U$42656 ( \43033 , \43032 );
not \U$42657 ( \43034 , \43019 );
or \U$42658 ( \43035 , \43033 , \43034 );
or \U$42659 ( \43036 , \43019 , \43032 );
nand \U$42660 ( \43037 , \43035 , \43036 );
and \U$42661 ( \43038 , \41979 , \43037 );
not \U$42662 ( \43039 , \41979 );
and \U$42663 ( \43040 , \43039 , RIc226bd8_22);
or \U$42664 ( \43041 , \43038 , \43040 );
buf \U$42665 ( \43042 , \43041 );
not \U$42666 ( \43043 , RIc226b60_23);
nor \U$42667 ( \43044 , \43043 , \41979 );
not \U$42668 ( \43045 , \43044 );
nand \U$42669 ( \43046 , \38284 , \38071 );
not \U$42670 ( \43047 , \43046 );
not \U$42671 ( \43048 , \43013 );
not \U$42672 ( \43049 , \42956 );
or \U$42673 ( \43050 , \43048 , \43049 );
nand \U$42674 ( \43051 , \43050 , \38281 );
not \U$42675 ( \43052 , \43051 );
or \U$42676 ( \43053 , \43047 , \43052 );
or \U$42677 ( \43054 , \43051 , \43046 );
nand \U$42678 ( \43055 , \43053 , \43054 );
nand \U$42679 ( \43056 , \43055 , \41979 );
nand \U$42680 ( \43057 , \43045 , \43056 );
buf \U$42681 ( \43058 , \43057 );
nand \U$42682 ( \43059 , \38281 , \43013 );
xnor \U$42683 ( \43060 , \42956 , \43059 );
and \U$42684 ( \43061 , \41979 , \43060 );
not \U$42685 ( \43062 , \41979 );
and \U$42686 ( \43063 , \43062 , RIc226ae8_24);
or \U$42687 ( \43064 , \43061 , \43063 );
buf \U$42688 ( \43065 , \43064 );
nand \U$42689 ( \43066 , \36633 , \36076 );
not \U$42690 ( \43067 , \43066 );
not \U$42691 ( \43068 , \38429 );
not \U$42692 ( \43069 , \36639 );
not \U$42693 ( \43070 , \38428 );
not \U$42694 ( \43071 , \41656 );
or \U$42695 ( \43072 , \43070 , \43071 );
nand \U$42696 ( \43073 , \43072 , \37683 );
not \U$42697 ( \43074 , \43073 );
or \U$42698 ( \43075 , \43069 , \43074 );
not \U$42699 ( \43076 , \36626 );
nand \U$42700 ( \43077 , \43075 , \43076 );
not \U$42701 ( \43078 , \43077 );
or \U$42702 ( \43079 , \43068 , \43078 );
buf \U$42703 ( \43080 , \36629 );
nand \U$42704 ( \43081 , \43079 , \43080 );
not \U$42705 ( \43082 , \43081 );
or \U$42706 ( \43083 , \43067 , \43082 );
or \U$42707 ( \43084 , \43081 , \43066 );
nand \U$42708 ( \43085 , \43083 , \43084 );
and \U$42709 ( \43086 , \41979 , \43085 );
not \U$42710 ( \43087 , \41979 );
and \U$42711 ( \43088 , \43087 , RIc226a70_25);
or \U$42712 ( \43089 , \43086 , \43088 );
buf \U$42713 ( \43090 , \43089 );
nand \U$42714 ( \43091 , \43080 , \38429 );
not \U$42715 ( \43092 , \43091 );
not \U$42716 ( \43093 , \43077 );
or \U$42717 ( \43094 , \43092 , \43093 );
or \U$42718 ( \43095 , \43077 , \43091 );
nand \U$42719 ( \43096 , \43094 , \43095 );
and \U$42720 ( \43097 , \41979 , \43096 );
not \U$42721 ( \43098 , \41979 );
and \U$42722 ( \43099 , \43098 , RIc2269f8_26);
or \U$42723 ( \43100 , \43097 , \43099 );
buf \U$42724 ( \43101 , \43100 );
not \U$42725 ( \43102 , \36593 );
nand \U$42726 ( \43103 , \43102 , \36625 );
not \U$42727 ( \43104 , \43103 );
not \U$42728 ( \43105 , \36637 );
not \U$42729 ( \43106 , \43073 );
or \U$42730 ( \43107 , \43105 , \43106 );
nand \U$42731 ( \43108 , \43107 , \36623 );
not \U$42732 ( \43109 , \43108 );
or \U$42733 ( \43110 , \43104 , \43109 );
or \U$42734 ( \43111 , \43108 , \43103 );
nand \U$42735 ( \43112 , \43110 , \43111 );
and \U$42736 ( \43113 , \41979 , \43112 );
not \U$42737 ( \43114 , \41979 );
and \U$42738 ( \43115 , \43114 , RIc226980_27);
or \U$42739 ( \43116 , \43113 , \43115 );
buf \U$42740 ( \43117 , \43116 );
not \U$42741 ( \43118 , RIc226908_28);
nor \U$42742 ( \43119 , \43118 , \41979 );
not \U$42743 ( \43120 , \43119 );
nand \U$42744 ( \43121 , \36623 , \36637 );
not \U$42745 ( \43122 , \43121 );
not \U$42746 ( \43123 , \43073 );
or \U$42747 ( \43124 , \43122 , \43123 );
or \U$42748 ( \43125 , \43073 , \43121 );
nand \U$42749 ( \43126 , \43124 , \43125 );
nand \U$42750 ( \43127 , \43126 , \41979 );
nand \U$42751 ( \43128 , \43120 , \43127 );
buf \U$42752 ( \43129 , \43128 );
not \U$42753 ( \43130 , RIc226890_29);
nor \U$42754 ( \43131 , \43130 , \41979 );
not \U$42755 ( \43132 , \43131 );
not \U$42756 ( \43133 , \37682 );
nand \U$42757 ( \43134 , \43133 , \37679 );
not \U$42758 ( \43135 , \43134 );
not \U$42759 ( \43136 , \38427 );
not \U$42760 ( \43137 , \38426 );
not \U$42761 ( \43138 , \41656 );
or \U$42762 ( \43139 , \43137 , \43138 );
nand \U$42763 ( \43140 , \43139 , \37643 );
not \U$42764 ( \43141 , \43140 );
or \U$42765 ( \43142 , \43136 , \43141 );
nand \U$42766 ( \43143 , \43142 , \37669 );
not \U$42767 ( \43144 , \43143 );
or \U$42768 ( \43145 , \43135 , \43144 );
or \U$42769 ( \43146 , \43143 , \43134 );
nand \U$42770 ( \43147 , \43145 , \43146 );
nand \U$42771 ( \43148 , \43147 , \41979 );
nand \U$42772 ( \43149 , \43132 , \43148 );
buf \U$42773 ( \43150 , \43149 );
not \U$42774 ( \43151 , RIc226818_30);
nor \U$42775 ( \43152 , \43151 , \41979 );
not \U$42776 ( \43153 , \43152 );
nand \U$42777 ( \43154 , \37669 , \38427 );
not \U$42778 ( \43155 , \43154 );
not \U$42779 ( \43156 , \43140 );
or \U$42780 ( \43157 , \43155 , \43156 );
or \U$42781 ( \43158 , \43140 , \43154 );
nand \U$42782 ( \43159 , \43157 , \43158 );
nand \U$42783 ( \43160 , \43159 , \41979 );
nand \U$42784 ( \43161 , \43153 , \43160 );
buf \U$42785 ( \43162 , \43161 );
not \U$42786 ( \43163 , RIc2267a0_31);
nor \U$42787 ( \43164 , \43163 , \41979 );
not \U$42788 ( \43165 , \43164 );
nand \U$42789 ( \43166 , \37381 , \37642 );
not \U$42790 ( \43167 , \43166 );
not \U$42791 ( \43168 , \38425 );
not \U$42792 ( \43169 , \41656 );
or \U$42793 ( \43170 , \43168 , \43169 );
buf \U$42794 ( \43171 , \37639 );
nand \U$42795 ( \43172 , \43170 , \43171 );
not \U$42796 ( \43173 , \43172 );
or \U$42797 ( \43174 , \43167 , \43173 );
or \U$42798 ( \43175 , \43172 , \43166 );
nand \U$42799 ( \43176 , \43174 , \43175 );
nand \U$42800 ( \43177 , \43176 , \41979 );
nand \U$42801 ( \43178 , \43165 , \43177 );
buf \U$42802 ( \43179 , \43178 );
nand \U$42803 ( \43180 , \38425 , \43171 );
xnor \U$42804 ( \43181 , \41656 , \43180 );
and \U$42805 ( \43182 , \41979 , \43181 );
not \U$42806 ( \43183 , \41979 );
and \U$42807 ( \43184 , \43183 , RIc226728_32);
or \U$42808 ( \43185 , \43182 , \43184 );
buf \U$42809 ( \43186 , \43185 );
not \U$42810 ( \43187 , RIc2266b0_33);
nor \U$42811 ( \43188 , \43187 , \41979 );
not \U$42812 ( \43189 , \43188 );
not \U$42813 ( \43190 , \41654 );
nand \U$42814 ( \43191 , \43190 , \41637 );
not \U$42815 ( \43192 , \43191 );
not \U$42816 ( \43193 , \41630 );
not \U$42817 ( \43194 , \41604 );
not \U$42818 ( \43195 , \40409 );
not \U$42819 ( \43196 , \41485 );
not \U$42820 ( \43197 , \41489 );
or \U$42821 ( \43198 , \43196 , \43197 );
nand \U$42822 ( \43199 , \43198 , \40405 );
not \U$42823 ( \43200 , \43199 );
or \U$42824 ( \43201 , \43195 , \43200 );
not \U$42825 ( \43202 , \39797 );
nand \U$42826 ( \43203 , \43201 , \43202 );
not \U$42827 ( \43204 , \43203 );
or \U$42828 ( \43205 , \43194 , \43204 );
not \U$42829 ( \43206 , \41648 );
nand \U$42830 ( \43207 , \43205 , \43206 );
not \U$42831 ( \43208 , \43207 );
or \U$42832 ( \43209 , \43193 , \43208 );
nand \U$42833 ( \43210 , \43209 , \41651 );
not \U$42834 ( \43211 , \43210 );
or \U$42835 ( \43212 , \43192 , \43211 );
or \U$42836 ( \43213 , \43210 , \43191 );
nand \U$42837 ( \43214 , \43212 , \43213 );
nand \U$42838 ( \43215 , \43214 , \41979 );
nand \U$42839 ( \43216 , \43189 , \43215 );
buf \U$42840 ( \43217 , \43216 );
not \U$42841 ( \43218 , \41979 );
and \U$42842 ( \43219 , \43218 , RIc226638_34);
not \U$42843 ( \43220 , \43218 );
nand \U$42844 ( \43221 , \41651 , \41630 );
not \U$42845 ( \43222 , \43221 );
not \U$42846 ( \43223 , \43207 );
or \U$42847 ( \43224 , \43222 , \43223 );
or \U$42848 ( \43225 , \43221 , \43207 );
nand \U$42849 ( \43226 , \43224 , \43225 );
and \U$42850 ( \43227 , \43220 , \43226 );
or \U$42851 ( \43228 , \43219 , \43227 );
buf \U$42852 ( \43229 , \43228 );
and \U$42853 ( \43230 , \43218 , \4376 );
not \U$42854 ( \43231 , \43218 );
not \U$42855 ( \43232 , \41603 );
not \U$42856 ( \43233 , \43203 );
or \U$42857 ( \43234 , \43232 , \43233 );
not \U$42858 ( \43235 , \41642 );
nand \U$42859 ( \43236 , \43234 , \43235 );
nand \U$42860 ( \43237 , \41647 , \41594 );
xor \U$42861 ( \43238 , \43236 , \43237 );
and \U$42862 ( \43239 , \43231 , \43238 );
nor \U$42863 ( \43240 , \43230 , \43239 );
buf \U$42864 ( \43241 , \43240 );
and \U$42865 ( \43242 , \43218 , RIc226548_36);
not \U$42866 ( \43243 , \43218 );
nand \U$42867 ( \43244 , \43235 , \41603 );
not \U$42868 ( \43245 , \43244 );
not \U$42869 ( \43246 , \43203 );
or \U$42870 ( \43247 , \43245 , \43246 );
or \U$42871 ( \43248 , \43244 , \43203 );
nand \U$42872 ( \43249 , \43247 , \43248 );
and \U$42873 ( \43250 , \43243 , \43249 );
or \U$42874 ( \43251 , \43242 , \43250 );
buf \U$42875 ( \43252 , \43251 );
not \U$42876 ( \43253 , RIc2264d0_37);
nor \U$42877 ( \43254 , \43253 , \41979 );
not \U$42878 ( \43255 , \43254 );
not \U$42879 ( \43256 , \39522 );
not \U$42880 ( \43257 , \39799 );
not \U$42881 ( \43258 , \43199 );
or \U$42882 ( \43259 , \43257 , \43258 );
not \U$42883 ( \43260 , \39787 );
nand \U$42884 ( \43261 , \43259 , \43260 );
not \U$42885 ( \43262 , \43261 );
or \U$42886 ( \43263 , \43256 , \43262 );
nand \U$42887 ( \43264 , \43263 , \39792 );
nand \U$42888 ( \43265 , \39796 , \39213 );
not \U$42889 ( \43266 , \43265 );
and \U$42890 ( \43267 , \43264 , \43266 );
not \U$42891 ( \43268 , \43264 );
and \U$42892 ( \43269 , \43268 , \43265 );
nor \U$42893 ( \43270 , \43267 , \43269 );
nand \U$42894 ( \43271 , \43270 , \41979 );
nand \U$42895 ( \43272 , \43255 , \43271 );
buf \U$42896 ( \43273 , \43272 );
and \U$42897 ( \43274 , \43218 , RIc226458_38);
not \U$42898 ( \43275 , \43218 );
nand \U$42899 ( \43276 , \39792 , \39522 );
xnor \U$42900 ( \43277 , \43261 , \43276 );
and \U$42901 ( \43278 , \43275 , \43277 );
or \U$42902 ( \43279 , \43274 , \43278 );
buf \U$42903 ( \43280 , \43279 );
and \U$42904 ( \43281 , \43218 , RIc2263e0_39);
not \U$42905 ( \43282 , \43218 );
nand \U$42906 ( \43283 , \39786 , \39692 );
not \U$42907 ( \43284 , \43283 );
not \U$42908 ( \43285 , \39798 );
not \U$42909 ( \43286 , \43199 );
or \U$42910 ( \43287 , \43285 , \43286 );
not \U$42911 ( \43288 , \39782 );
nand \U$42912 ( \43289 , \43287 , \43288 );
not \U$42913 ( \43290 , \43289 );
or \U$42914 ( \43291 , \43284 , \43290 );
or \U$42915 ( \43292 , \43289 , \43283 );
nand \U$42916 ( \43293 , \43291 , \43292 );
and \U$42917 ( \43294 , \43282 , \43293 );
or \U$42918 ( \43295 , \43281 , \43294 );
buf \U$42919 ( \43296 , \43295 );
and \U$42920 ( \43297 , \43218 , RIc226368_40);
not \U$42921 ( \43298 , \43218 );
and \U$42922 ( \43299 , \43288 , \39798 );
xor \U$42923 ( \43300 , \43199 , \43299 );
and \U$42924 ( \43301 , \43298 , \43300 );
or \U$42925 ( \43302 , \43297 , \43301 );
buf \U$42926 ( \43303 , \43302 );
not \U$42927 ( \43304 , RIc2262f0_41);
nor \U$42928 ( \43305 , \43304 , \41979 );
not \U$42929 ( \43306 , \43305 );
not \U$42930 ( \43307 , \41488 );
not \U$42931 ( \43308 , \41487 );
not \U$42932 ( \43309 , \41485 );
or \U$42933 ( \43310 , \43308 , \43309 );
nand \U$42934 ( \43311 , \43310 , \40361 );
not \U$42935 ( \43312 , \43311 );
or \U$42936 ( \43313 , \43307 , \43312 );
nand \U$42937 ( \43314 , \43313 , \40390 );
not \U$42938 ( \43315 , \40404 );
nand \U$42939 ( \43316 , \43315 , \40402 );
not \U$42940 ( \43317 , \43316 );
and \U$42941 ( \43318 , \43314 , \43317 );
not \U$42942 ( \43319 , \43314 );
and \U$42943 ( \43320 , \43319 , \43316 );
nor \U$42944 ( \43321 , \43318 , \43320 );
nand \U$42945 ( \43322 , \43321 , \41979 );
nand \U$42946 ( \43323 , \43306 , \43322 );
buf \U$42947 ( \43324 , \43323 );
and \U$42948 ( \43325 , \43218 , RIc226278_42);
not \U$42949 ( \43326 , \43218 );
not \U$42950 ( \43327 , \40388 );
nand \U$42951 ( \43328 , \43327 , \40390 );
xnor \U$42952 ( \43329 , \43311 , \43328 );
and \U$42953 ( \43330 , \43326 , \43329 );
or \U$42954 ( \43331 , \43325 , \43330 );
buf \U$42955 ( \43332 , \43331 );
and \U$42956 ( \43333 , \43218 , RIc226200_43);
not \U$42957 ( \43334 , \43218 );
not \U$42958 ( \43335 , \41486 );
not \U$42959 ( \43336 , \41485 );
or \U$42960 ( \43337 , \43335 , \43336 );
nand \U$42961 ( \43338 , \43337 , \40358 );
nand \U$42962 ( \43339 , \40254 , \40360 );
not \U$42963 ( \43340 , \43339 );
and \U$42964 ( \43341 , \43338 , \43340 );
not \U$42965 ( \43342 , \43338 );
and \U$42966 ( \43343 , \43342 , \43339 );
nor \U$42967 ( \43344 , \43341 , \43343 );
and \U$42968 ( \43345 , \43334 , \43344 );
or \U$42969 ( \43346 , \43333 , \43345 );
buf \U$42970 ( \43347 , \43346 );
and \U$42971 ( \43348 , \43218 , RIc226188_44);
not \U$42972 ( \43349 , \43218 );
and \U$42973 ( \43350 , \40358 , \41486 );
xor \U$42974 ( \43351 , \41485 , \43350 );
and \U$42975 ( \43352 , \43349 , \43351 );
or \U$42976 ( \43353 , \43348 , \43352 );
buf \U$42977 ( \43354 , \43353 );
not \U$42978 ( \43355 , RIc226110_45);
nor \U$42979 ( \43356 , \43355 , \41979 );
not \U$42980 ( \43357 , \43356 );
not \U$42981 ( \43358 , \40758 );
not \U$42982 ( \43359 , \41481 );
not \U$42983 ( \43360 , \40776 );
or \U$42984 ( \43361 , \43359 , \43360 );
nand \U$42985 ( \43362 , \43361 , \40741 );
not \U$42986 ( \43363 , \43362 );
or \U$42987 ( \43364 , \43358 , \43363 );
not \U$42988 ( \43365 , \40761 );
nand \U$42989 ( \43366 , \43364 , \43365 );
nand \U$42990 ( \43367 , \41484 , \40773 );
not \U$42991 ( \43368 , \43367 );
and \U$42992 ( \43369 , \43366 , \43368 );
not \U$42993 ( \43370 , \43366 );
and \U$42994 ( \43371 , \43370 , \43367 );
nor \U$42995 ( \43372 , \43369 , \43371 );
nand \U$42996 ( \43373 , \43372 , \41979 );
nand \U$42997 ( \43374 , \43357 , \43373 );
buf \U$42998 ( \43375 , \43374 );
not \U$42999 ( \43376 , \41979 );
not \U$43000 ( \43377 , \40761 );
nand \U$43001 ( \43378 , \43377 , \40758 );
not \U$43002 ( \43379 , \43378 );
not \U$43003 ( \43380 , \43362 );
or \U$43004 ( \43381 , \43379 , \43380 );
or \U$43005 ( \43382 , \43362 , \43378 );
nand \U$43006 ( \43383 , \43381 , \43382 );
not \U$43007 ( \43384 , \43383 );
or \U$43008 ( \43385 , \43376 , \43384 );
nand \U$43009 ( \43386 , \43218 , RIc226098_46);
nand \U$43010 ( \43387 , \43385 , \43386 );
buf \U$43011 ( \43388 , \43387 );
not \U$43012 ( \43389 , \41979 );
not \U$43013 ( \43390 , \41481 );
not \U$43014 ( \43391 , \40775 );
or \U$43015 ( \43392 , \43390 , \43391 );
nand \U$43016 ( \43393 , \43392 , \40739 );
not \U$43017 ( \43394 , \43393 );
nand \U$43018 ( \43395 , \40644 , \40643 );
not \U$43019 ( \43396 , \43395 );
or \U$43020 ( \43397 , \43394 , \43396 );
or \U$43021 ( \43398 , \43395 , \43393 );
nand \U$43022 ( \43399 , \43397 , \43398 );
not \U$43023 ( \43400 , \43399 );
or \U$43024 ( \43401 , \43389 , \43400 );
nand \U$43025 ( \43402 , \43218 , RIc226020_47);
nand \U$43026 ( \43403 , \43401 , \43402 );
buf \U$43027 ( \43404 , \43403 );
and \U$43028 ( \43405 , \43218 , RIc225fa8_48);
not \U$43029 ( \43406 , \43218 );
nand \U$43030 ( \43407 , \40739 , \40775 );
xor \U$43031 ( \43408 , \43390 , \43407 );
and \U$43032 ( \43409 , \43406 , \43408 );
or \U$43033 ( \43410 , \43405 , \43409 );
buf \U$43034 ( \43411 , \43410 );
and \U$43035 ( \43412 , \43218 , RIc225f30_49);
not \U$43036 ( \43413 , \43218 );
not \U$43037 ( \43414 , \40963 );
not \U$43038 ( \43415 , \41464 );
not \U$43039 ( \43416 , \41439 );
or \U$43040 ( \43417 , \43415 , \43416 );
not \U$43041 ( \43418 , \41470 );
nand \U$43042 ( \43419 , \43417 , \43418 );
not \U$43043 ( \43420 , \43419 );
or \U$43044 ( \43421 , \43414 , \43420 );
nand \U$43045 ( \43422 , \43421 , \41475 );
nand \U$43046 ( \43423 , \41480 , \41477 );
not \U$43047 ( \43424 , \43423 );
and \U$43048 ( \43425 , \43422 , \43424 );
not \U$43049 ( \43426 , \43422 );
and \U$43050 ( \43427 , \43426 , \43423 );
nor \U$43051 ( \43428 , \43425 , \43427 );
and \U$43052 ( \43429 , \43413 , \43428 );
or \U$43053 ( \43430 , \43412 , \43429 );
buf \U$43054 ( \43431 , \43430 );
and \U$43055 ( \43432 , \43218 , RIc225eb8_50);
not \U$43056 ( \43433 , \43218 );
nand \U$43057 ( \43434 , \40963 , \41475 );
xnor \U$43058 ( \43435 , \43419 , \43434 );
and \U$43059 ( \43436 , \43433 , \43435 );
or \U$43060 ( \43437 , \43432 , \43436 );
buf \U$43061 ( \43438 , \43437 );
and \U$43062 ( \43439 , \43218 , RIc225e40_51);
not \U$43063 ( \43440 , \43218 );
not \U$43064 ( \43441 , \41463 );
not \U$43065 ( \43442 , \43441 );
not \U$43066 ( \43443 , \41439 );
or \U$43067 ( \43444 , \43442 , \43443 );
nand \U$43068 ( \43445 , \43444 , \41467 );
not \U$43069 ( \43446 , \41456 );
nand \U$43070 ( \43447 , \43446 , \41469 );
xnor \U$43071 ( \43448 , \43445 , \43447 );
and \U$43072 ( \43449 , \43440 , \43448 );
or \U$43073 ( \43450 , \43439 , \43449 );
buf \U$43074 ( \43451 , \43450 );
not \U$43075 ( \43452 , \41979 );
nand \U$43076 ( \43453 , \43441 , \41467 );
not \U$43077 ( \43454 , \43453 );
not \U$43078 ( \43455 , \41439 );
or \U$43079 ( \43456 , \43454 , \43455 );
or \U$43080 ( \43457 , \41439 , \43453 );
nand \U$43081 ( \43458 , \43456 , \43457 );
not \U$43082 ( \43459 , \43458 );
or \U$43083 ( \43460 , \43452 , \43459 );
nand \U$43084 ( \43461 , \43218 , RIc225dc8_52);
nand \U$43085 ( \43462 , \43460 , \43461 );
buf \U$43086 ( \43463 , \43462 );
not \U$43087 ( \43464 , \41979 );
xor \U$43088 ( \43465 , \41096 , \41117 );
xor \U$43089 ( \43466 , \43465 , \41436 );
not \U$43090 ( \43467 , \43466 );
or \U$43091 ( \43468 , \43464 , \43467 );
nand \U$43092 ( \43469 , \43218 , RIc225d50_53);
nand \U$43093 ( \43470 , \43468 , \43469 );
buf \U$43094 ( \43471 , \43470 );
not \U$43095 ( \43472 , \41978 );
not \U$43096 ( \43473 , RIc225cd8_54);
or \U$43097 ( \43474 , \43472 , \43473 );
nand \U$43098 ( \43475 , \41435 , \41171 );
xnor \U$43099 ( \43476 , \41431 , \43475 );
nand \U$43100 ( \43477 , \43476 , \41979 );
nand \U$43101 ( \43478 , \43474 , \43477 );
buf \U$43102 ( \43479 , \43478 );
and \U$43103 ( \43480 , \41978 , RIc225c60_55);
not \U$43104 ( \43481 , \41978 );
nand \U$43105 ( \43482 , \41422 , \41250 );
not \U$43106 ( \43483 , \41425 );
nand \U$43107 ( \43484 , \43482 , \43483 );
nand \U$43108 ( \43485 , \41266 , \41429 );
xnor \U$43109 ( \43486 , \43484 , \43485 );
and \U$43110 ( \43487 , \43481 , \43486 );
or \U$43111 ( \43488 , \43480 , \43487 );
buf \U$43112 ( \43489 , \43488 );
endmodule

