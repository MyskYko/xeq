//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RIbb2d630_69,RIbb317d0_133,RIbb2d5b8_70,RIbb31848_134,RIbb2d540_71,RIbb318c0_135,RIbb2d4c8_72,RIbb31938_136,RIbb2d720_67,
        RIbb316e0_131,RIbb2d6a8_68,RIbb31758_132,RIbb2d798_66,RIbb31668_130,RIbb2d810_65,RIbb315f0_129,RIbb2cfa0_83,RIbb31e60_147,RIbb2cf28_84,
        RIbb31ed8_148,RIbb2d090_81,RIbb31d70_145,RIbb2d018_82,RIbb31de8_146,RIbb2caf0_93,RIbb32310_157,RIbb2ca78_94,RIbb32388_158,RIbb2ca00_95,
        RIbb32400_159,RIbb2c988_96,RIbb32478_160,RIbb2cc58_90,RIbb321a8_154,RIbb2ccd0_89,RIbb32130_153,RIbb2cbe0_91,RIbb32220_155,RIbb2cb68_92,
        RIbb32298_156,RIbb2cdc0_87,RIbb32040_151,RIbb2cd48_88,RIbb320b8_152,RIbb2ceb0_85,RIbb31f50_149,RIbb2ce38_86,RIbb31fc8_150,RIbb2d360_75,
        RIbb31aa0_139,RIbb2d2e8_76,RIbb31b18_140,RIbb2d3d8_74,RIbb31a28_138,RIbb2d450_73,RIbb319b0_137,RIbb2d180_79,RIbb31c80_143,RIbb2d108_80,
        RIbb31cf8_144,RIbb2d270_77,RIbb31b90_141,RIbb2d1f8_78,RIbb31c08_142,RIbb2be48_120,RIbb32fb8_184,RIbb2bec0_119,RIbb32f40_183,RIbb2bfb0_117,
        RIbb32e50_181,RIbb2bf38_118,RIbb32ec8_182,RIbb2c0a0_115,RIbb32d60_179,RIbb2c028_116,RIbb32dd8_180,RIbb2c118_114,RIbb32ce8_178,RIbb2c190_113,
        RIbb32c70_177,RIbb2bbf0_125,RIbb33210_189,RIbb2bb78_126,RIbb33288_190,RIbb31578_128,RIbb33378_192,RIbb31500_127,RIbb33300_191,RIbb2bce0_123,
        RIbb33120_187,RIbb2bc68_124,RIbb33198_188,RIbb2bdd0_121,RIbb33030_185,RIbb2bd58_122,RIbb330a8_186,RIbb2c370_109,RIbb32a90_173,RIbb2c280_111,
        RIbb32b80_175,RIbb2c460_107,RIbb329a0_171,RIbb2c550_105,RIbb328b0_169,RIbb2c2f8_110,RIbb32b08_174,RIbb2c3e8_108,RIbb32a18_172,RIbb2c208_112,
        RIbb32bf8_176,RIbb2c4d8_106,RIbb32928_170,RIbb2c640_103,RIbb327c0_167,RIbb2c5c8_104,RIbb32838_168,RIbb2c6b8_102,RIbb32748_166,RIbb2c730_101,
        RIbb326d0_165,RIbb2c898_98,RIbb32568_162,RIbb2c910_97,RIbb324f0_161,RIbb2c7a8_100,RIbb32658_164,RIbb2c820_99,RIbb325e0_163,RIbb2ee90_17,
        RIbb2ee18_18,RIbb2eda0_19,RIbb2ed28_20,RIbb2ecb0_21,RIbb2f070_13,RIbb2eff8_14,RIbb2ef80_15,RIbb2f160_11,RIbb2f0e8_12,RIbb2f340_7,
        RIbb2f3b8_6,RIbb2f430_5,RIbb2f520_3,RIbb2f4a8_4,RIbb2f610_1,RIbb2f598_2,RIbb2ef08_16,RIbb2f250_9,RIbb2f1d8_10,RIbb2f2c8_8,
        RIbb2ec38_22,RIbb2ebc0_23,RIbb2e8f0_29,RIbb2e878_30,RIbb2e800_31,RIbb2e788_32,RIbb2e710_33,RIbb2e9e0_27,RIbb2ea58_26,RIbb2ead0_25,
        RIbb2eb48_24,RIbb2e968_28,RIbb2e698_34,RIbb2e620_35,RIbb2e5a8_36,RIbb2e530_37,RIbb2e440_39,RIbb2e4b8_38,RIbb2e3c8_40,RIbb2e350_41,
        RIbb2e260_43,RIbb2e2d8_42,RIbb2e1e8_44,RIbb2e170_45,RIbb2e0f8_46,RIbb2e080_47,RIbb2e008_48,RIbb2df90_49,RIbb2df18_50,RIbb2dea0_51,
        RIbb2ddb0_53,RIbb2de28_52,RIbb2dd38_54,RIbb2dcc0_55,RIbb2dbd0_57,RIbb2dc48_56,RIbb2db58_58,RIbb2dae0_59,RIbb2da68_60,RIbb2d9f0_61,
        RIbb2d900_63,RIbb2d978_62,RIbb2d888_64,RIbb345c0_231,RIbb34bd8_244,RIbb336c0_199,RIbb34278_224,RIbb338a0_203,RIbb34db8_248,RIbb34098_220,
        RIbb33a08_206,RIbb34110_221,RIbb33990_205,RIbb347a0_235,RIbb34cc8_246,RIbb33c60_211,RIbb34d40_247,RIbb33f30_217,RIbb33d50_213,RIbb34548_230,
        RIbb34ea8_250,RIbb34908_238,RIbb33a80_207,RIbb334e0_195,RIbb35010_253,RIbb33738_200,RIbb349f8_240,RIbb33918_204,RIbb34980_239,RIbb33828_202,
        RIbb34188_222,RIbb34728_234,RIbb35088_254,RIbb346b0_233,RIbb34638_232,RIbb34458_228,RIbb34ae8_242,RIbb33b70_209,RIbb33fa8_218,RIbb33558_196,
        RIbb34e30_249,RIbb33af8_208,RIbb34020_219,RIbb333f0_193,RIbb35178_256,RIbb343e0_227,RIbb34368_226,RIbb34a70_241,RIbb335d0_197,RIbb344d0_229,
        RIbb34b60_243,RIbb33be8_210,RIbb34f98_252,RIbb33cd8_212,RIbb34890_237,RIbb342f0_225,RIbb33648_198,RIbb34c50_245,RIbb34f20_251,RIbb33468_194,
        RIbb35100_255,RIbb337b0_201,RIbb34200_223,RIbb33eb8_216,RIbb34818_236,RIbb33dc8_214,RIbb33e40_215,R_109_95e4d78,R_10a_95e4e20,R_10c_95e4f70,
        R_10f_95e5168,R_111_95e52b8,R_119_95e57f8,R_11c_95e59f0,R_11d_95e5a98,R_11f_95e5be8,R_122_95e5de0,R_123_95e5e88,R_124_95e5f30,R_125_95e5fd8,
        R_127_95e6128,R_128_95e61d0,R_129_95e6278,R_12b_95e63c8,R_12c_95e6470,R_12e_95e65c0,R_12f_95e6668,R_130_95e6710,R_131_95e67b8,R_135_95e6a58,
        R_136_95e6b00,R_137_95e6ba8,R_138_95e6c50,R_139_95e6cf8,R_13b_95e6e48,R_13d_95e6f98,R_13e_95e7040,R_13f_95e70e8,R_140_95e7190,R_141_95e7238,
        R_143_95e7388,R_144_95e7430,R_145_95e74d8,R_146_95e7580,R_147_95e7628,R_148_95e76d0,R_149_95e7778,R_14a_95e7820,R_14b_95e78c8,R_14c_95e7970,
        R_14d_95e7a18,R_14e_95e7ac0,R_14f_95e7b68,R_150_95e7c10,R_151_95e7cb8,R_152_95e7d60,R_153_95e7e08,R_154_95e7eb0,R_155_95e7f58,R_156_95e8000,
        R_157_95e80a8,R_158_95e8150,R_159_95e81f8,R_15a_95e82a0,R_15b_95e8348,R_15c_95e83f0,R_15d_95e8498,R_15e_95e8540,R_15f_95e85e8,R_160_95e8690,
        R_161_95e8738,R_162_95e87e0,R_163_95e8888,R_164_95e8930,R_165_95e89d8,R_166_95e8a80,R_167_95e8b28,R_168_95e8bd0,R_169_95e8c78,R_16a_95e8d20,
        R_16b_95e8dc8,R_16c_95e8e70,R_16d_95e8f18,R_16e_95e8fc0,R_16f_95e9068,R_170_95e9110,R_171_95e91b8,R_172_95e9260,R_173_95e9308,R_174_95e93b0,
        R_175_95e9458,R_176_95e9500);
input RIbb2d630_69,RIbb317d0_133,RIbb2d5b8_70,RIbb31848_134,RIbb2d540_71,RIbb318c0_135,RIbb2d4c8_72,RIbb31938_136,RIbb2d720_67,
        RIbb316e0_131,RIbb2d6a8_68,RIbb31758_132,RIbb2d798_66,RIbb31668_130,RIbb2d810_65,RIbb315f0_129,RIbb2cfa0_83,RIbb31e60_147,RIbb2cf28_84,
        RIbb31ed8_148,RIbb2d090_81,RIbb31d70_145,RIbb2d018_82,RIbb31de8_146,RIbb2caf0_93,RIbb32310_157,RIbb2ca78_94,RIbb32388_158,RIbb2ca00_95,
        RIbb32400_159,RIbb2c988_96,RIbb32478_160,RIbb2cc58_90,RIbb321a8_154,RIbb2ccd0_89,RIbb32130_153,RIbb2cbe0_91,RIbb32220_155,RIbb2cb68_92,
        RIbb32298_156,RIbb2cdc0_87,RIbb32040_151,RIbb2cd48_88,RIbb320b8_152,RIbb2ceb0_85,RIbb31f50_149,RIbb2ce38_86,RIbb31fc8_150,RIbb2d360_75,
        RIbb31aa0_139,RIbb2d2e8_76,RIbb31b18_140,RIbb2d3d8_74,RIbb31a28_138,RIbb2d450_73,RIbb319b0_137,RIbb2d180_79,RIbb31c80_143,RIbb2d108_80,
        RIbb31cf8_144,RIbb2d270_77,RIbb31b90_141,RIbb2d1f8_78,RIbb31c08_142,RIbb2be48_120,RIbb32fb8_184,RIbb2bec0_119,RIbb32f40_183,RIbb2bfb0_117,
        RIbb32e50_181,RIbb2bf38_118,RIbb32ec8_182,RIbb2c0a0_115,RIbb32d60_179,RIbb2c028_116,RIbb32dd8_180,RIbb2c118_114,RIbb32ce8_178,RIbb2c190_113,
        RIbb32c70_177,RIbb2bbf0_125,RIbb33210_189,RIbb2bb78_126,RIbb33288_190,RIbb31578_128,RIbb33378_192,RIbb31500_127,RIbb33300_191,RIbb2bce0_123,
        RIbb33120_187,RIbb2bc68_124,RIbb33198_188,RIbb2bdd0_121,RIbb33030_185,RIbb2bd58_122,RIbb330a8_186,RIbb2c370_109,RIbb32a90_173,RIbb2c280_111,
        RIbb32b80_175,RIbb2c460_107,RIbb329a0_171,RIbb2c550_105,RIbb328b0_169,RIbb2c2f8_110,RIbb32b08_174,RIbb2c3e8_108,RIbb32a18_172,RIbb2c208_112,
        RIbb32bf8_176,RIbb2c4d8_106,RIbb32928_170,RIbb2c640_103,RIbb327c0_167,RIbb2c5c8_104,RIbb32838_168,RIbb2c6b8_102,RIbb32748_166,RIbb2c730_101,
        RIbb326d0_165,RIbb2c898_98,RIbb32568_162,RIbb2c910_97,RIbb324f0_161,RIbb2c7a8_100,RIbb32658_164,RIbb2c820_99,RIbb325e0_163,RIbb2ee90_17,
        RIbb2ee18_18,RIbb2eda0_19,RIbb2ed28_20,RIbb2ecb0_21,RIbb2f070_13,RIbb2eff8_14,RIbb2ef80_15,RIbb2f160_11,RIbb2f0e8_12,RIbb2f340_7,
        RIbb2f3b8_6,RIbb2f430_5,RIbb2f520_3,RIbb2f4a8_4,RIbb2f610_1,RIbb2f598_2,RIbb2ef08_16,RIbb2f250_9,RIbb2f1d8_10,RIbb2f2c8_8,
        RIbb2ec38_22,RIbb2ebc0_23,RIbb2e8f0_29,RIbb2e878_30,RIbb2e800_31,RIbb2e788_32,RIbb2e710_33,RIbb2e9e0_27,RIbb2ea58_26,RIbb2ead0_25,
        RIbb2eb48_24,RIbb2e968_28,RIbb2e698_34,RIbb2e620_35,RIbb2e5a8_36,RIbb2e530_37,RIbb2e440_39,RIbb2e4b8_38,RIbb2e3c8_40,RIbb2e350_41,
        RIbb2e260_43,RIbb2e2d8_42,RIbb2e1e8_44,RIbb2e170_45,RIbb2e0f8_46,RIbb2e080_47,RIbb2e008_48,RIbb2df90_49,RIbb2df18_50,RIbb2dea0_51,
        RIbb2ddb0_53,RIbb2de28_52,RIbb2dd38_54,RIbb2dcc0_55,RIbb2dbd0_57,RIbb2dc48_56,RIbb2db58_58,RIbb2dae0_59,RIbb2da68_60,RIbb2d9f0_61,
        RIbb2d900_63,RIbb2d978_62,RIbb2d888_64,RIbb345c0_231,RIbb34bd8_244,RIbb336c0_199,RIbb34278_224,RIbb338a0_203,RIbb34db8_248,RIbb34098_220,
        RIbb33a08_206,RIbb34110_221,RIbb33990_205,RIbb347a0_235,RIbb34cc8_246,RIbb33c60_211,RIbb34d40_247,RIbb33f30_217,RIbb33d50_213,RIbb34548_230,
        RIbb34ea8_250,RIbb34908_238,RIbb33a80_207,RIbb334e0_195,RIbb35010_253,RIbb33738_200,RIbb349f8_240,RIbb33918_204,RIbb34980_239,RIbb33828_202,
        RIbb34188_222,RIbb34728_234,RIbb35088_254,RIbb346b0_233,RIbb34638_232,RIbb34458_228,RIbb34ae8_242,RIbb33b70_209,RIbb33fa8_218,RIbb33558_196,
        RIbb34e30_249,RIbb33af8_208,RIbb34020_219,RIbb333f0_193,RIbb35178_256,RIbb343e0_227,RIbb34368_226,RIbb34a70_241,RIbb335d0_197,RIbb344d0_229,
        RIbb34b60_243,RIbb33be8_210,RIbb34f98_252,RIbb33cd8_212,RIbb34890_237,RIbb342f0_225,RIbb33648_198,RIbb34c50_245,RIbb34f20_251,RIbb33468_194,
        RIbb35100_255,RIbb337b0_201,RIbb34200_223,RIbb33eb8_216,RIbb34818_236,RIbb33dc8_214,RIbb33e40_215;
output R_109_95e4d78,R_10a_95e4e20,R_10c_95e4f70,R_10f_95e5168,R_111_95e52b8,R_119_95e57f8,R_11c_95e59f0,R_11d_95e5a98,R_11f_95e5be8,
        R_122_95e5de0,R_123_95e5e88,R_124_95e5f30,R_125_95e5fd8,R_127_95e6128,R_128_95e61d0,R_129_95e6278,R_12b_95e63c8,R_12c_95e6470,R_12e_95e65c0,
        R_12f_95e6668,R_130_95e6710,R_131_95e67b8,R_135_95e6a58,R_136_95e6b00,R_137_95e6ba8,R_138_95e6c50,R_139_95e6cf8,R_13b_95e6e48,R_13d_95e6f98,
        R_13e_95e7040,R_13f_95e70e8,R_140_95e7190,R_141_95e7238,R_143_95e7388,R_144_95e7430,R_145_95e74d8,R_146_95e7580,R_147_95e7628,R_148_95e76d0,
        R_149_95e7778,R_14a_95e7820,R_14b_95e78c8,R_14c_95e7970,R_14d_95e7a18,R_14e_95e7ac0,R_14f_95e7b68,R_150_95e7c10,R_151_95e7cb8,R_152_95e7d60,
        R_153_95e7e08,R_154_95e7eb0,R_155_95e7f58,R_156_95e8000,R_157_95e80a8,R_158_95e8150,R_159_95e81f8,R_15a_95e82a0,R_15b_95e8348,R_15c_95e83f0,
        R_15d_95e8498,R_15e_95e8540,R_15f_95e85e8,R_160_95e8690,R_161_95e8738,R_162_95e87e0,R_163_95e8888,R_164_95e8930,R_165_95e89d8,R_166_95e8a80,
        R_167_95e8b28,R_168_95e8bd0,R_169_95e8c78,R_16a_95e8d20,R_16b_95e8dc8,R_16c_95e8e70,R_16d_95e8f18,R_16e_95e8fc0,R_16f_95e9068,R_170_95e9110,
        R_171_95e91b8,R_172_95e9260,R_173_95e9308,R_174_95e93b0,R_175_95e9458,R_176_95e9500;

wire \342_ZERO , \343_ONE , \344 , \345 , \346 , \347 , \348 , \349 , \350 ,
         \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 ,
         \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 ,
         \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 ,
         \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 ,
         \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 ,
         \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 ,
         \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 ,
         \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 ,
         \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 ,
         \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 ,
         \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 ,
         \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 ,
         \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 ,
         \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 ,
         \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 ,
         \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 ,
         \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 ,
         \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 ,
         \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 ,
         \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 ,
         \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 ,
         \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 ,
         \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 ,
         \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 ,
         \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 ,
         \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 ,
         \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 ,
         \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 ,
         \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 ,
         \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 ,
         \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 ,
         \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 ,
         \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 ,
         \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 ,
         \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 ,
         \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 ,
         \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 ,
         \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 ,
         \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 ,
         \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 ,
         \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 ,
         \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 ,
         \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 ,
         \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 ,
         \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 ,
         \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 ,
         \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 ,
         \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 ,
         \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 ,
         \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 ,
         \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 ,
         \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 ,
         \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 ,
         \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 ,
         \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 ,
         \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 ,
         \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 ,
         \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 ,
         \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 ,
         \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 ,
         \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 ,
         \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 ,
         \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 ,
         \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 ,
         \991 , \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 ,
         \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 ,
         \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 ,
         \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 ,
         \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 ,
         \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 ,
         \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 ,
         \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 ,
         \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 ,
         \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 ,
         \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 ,
         \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 ,
         \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 ,
         \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 ,
         \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 ,
         \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 ,
         \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 ,
         \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 ,
         \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 ,
         \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 ,
         \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 ,
         \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 ,
         \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 ,
         \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 ,
         \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 ,
         \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 ,
         \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 ,
         \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 ,
         \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 ,
         \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 ,
         \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 ,
         \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 ,
         \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 ,
         \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 ,
         \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 ,
         \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 ,
         \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 ,
         \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 ,
         \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 ,
         \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 ,
         \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 ,
         \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 ,
         \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 ,
         \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 ,
         \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 ,
         \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 ,
         \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 ,
         \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 ,
         \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 ,
         \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 ,
         \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 ,
         \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 ,
         \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 ,
         \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 ,
         \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 ,
         \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 ,
         \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 ,
         \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 ,
         \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 ,
         \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 ,
         \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 ,
         \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 ,
         \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 ,
         \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 ,
         \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 ,
         \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 ,
         \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 ,
         \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 ,
         \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 ,
         \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 ,
         \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 ,
         \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 ,
         \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 ,
         \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 ,
         \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 ,
         \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 ,
         \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 ,
         \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 ,
         \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 ,
         \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 ,
         \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 ,
         \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 ,
         \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 ,
         \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 ,
         \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 ,
         \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 ,
         \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 ,
         \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 ,
         \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 ,
         \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 ,
         \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 ,
         \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 ,
         \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 ,
         \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 ,
         \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 ,
         \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 ,
         \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 ,
         \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 ,
         \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 ,
         \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 ,
         \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 ,
         \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 ,
         \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 ,
         \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 ,
         \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 ,
         \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 ,
         \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 ,
         \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 ,
         \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 ,
         \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 ,
         \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 ,
         \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 ,
         \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 ,
         \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 ,
         \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 ,
         \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 ,
         \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 ,
         \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 ,
         \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 ,
         \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 ,
         \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 ,
         \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 ,
         \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 ,
         \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 ,
         \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 ,
         \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 ,
         \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 ,
         \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 ,
         \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 ,
         \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 ,
         \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 ,
         \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 ,
         \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 ,
         \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 ,
         \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 ,
         \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 ,
         \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 ,
         \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 ,
         \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 ,
         \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 ,
         \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 ,
         \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 ,
         \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 ,
         \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 ,
         \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 ,
         \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 ,
         \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 ,
         \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 ,
         \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 ,
         \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 ,
         \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 ,
         \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 ,
         \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 ,
         \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 ,
         \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 ,
         \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 ,
         \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 ,
         \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 ,
         \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 ,
         \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 ,
         \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 ,
         \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 ,
         \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 ,
         \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 ,
         \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 ,
         \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 ,
         \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 ,
         \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 ,
         \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 ,
         \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 ,
         \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 ,
         \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 ,
         \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 ,
         \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 ,
         \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 ,
         \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 ,
         \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 ,
         \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 ,
         \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 ,
         \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 ,
         \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 ,
         \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 ,
         \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 ,
         \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 ,
         \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 ,
         \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 ,
         \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 ,
         \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 ,
         \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 ,
         \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 ,
         \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 ,
         \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 ,
         \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 ,
         \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 ,
         \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 ,
         \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 ,
         \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 ,
         \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 ,
         \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 ,
         \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 ,
         \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 ,
         \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 ,
         \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 ,
         \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 ,
         \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 ,
         \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 ,
         \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 ,
         \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 ,
         \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 ,
         \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 ,
         \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 ,
         \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 ,
         \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 ,
         \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 ,
         \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 ,
         \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 ,
         \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 ,
         \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 ,
         \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 ,
         \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 ,
         \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 ,
         \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 ,
         \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 ,
         \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 ,
         \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 ,
         \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 ,
         \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 ,
         \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 ,
         \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 ,
         \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 ,
         \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 ,
         \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 ,
         \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 ,
         \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 ,
         \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 ,
         \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 ,
         \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 ,
         \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 ,
         \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 ,
         \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 ,
         \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 ,
         \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 ,
         \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 ,
         \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 ,
         \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 ,
         \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 ,
         \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 ,
         \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 ,
         \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 ,
         \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 ,
         \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 ,
         \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 ,
         \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 ,
         \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 ,
         \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 ,
         \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 ,
         \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 ,
         \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 ,
         \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 ,
         \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 ,
         \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 ,
         \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 ,
         \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 ,
         \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 ,
         \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 ,
         \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 ,
         \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 ,
         \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 ,
         \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 ,
         \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 ,
         \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 ,
         \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 ,
         \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 ,
         \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 ,
         \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 ,
         \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 ,
         \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 ,
         \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 ,
         \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 ,
         \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 ,
         \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 ,
         \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 ,
         \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 ,
         \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 ,
         \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 ,
         \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 ,
         \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 ,
         \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 ,
         \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 ,
         \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 ,
         \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 ,
         \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 ,
         \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 ,
         \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 ,
         \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 ,
         \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 ,
         \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 ,
         \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 ,
         \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 ,
         \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 ,
         \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 ,
         \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 ,
         \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 ,
         \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 ,
         \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 ,
         \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 ,
         \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 ,
         \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 ,
         \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 ,
         \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 ,
         \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 ,
         \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 ,
         \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 ,
         \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 ,
         \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 ,
         \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 ,
         \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 ,
         \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 ,
         \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 ,
         \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 ,
         \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 ,
         \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 ,
         \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 ,
         \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 ,
         \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 ,
         \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 ,
         \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 ,
         \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 ,
         \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 ,
         \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 ,
         \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 ,
         \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 ,
         \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 ,
         \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 ,
         \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 ,
         \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 ,
         \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 ,
         \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 ,
         \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 ,
         \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 ,
         \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 ,
         \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 ,
         \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 ,
         \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 ,
         \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 ,
         \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 ,
         \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 ,
         \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 ,
         \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 ,
         \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 ,
         \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 ,
         \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 ,
         \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 ,
         \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 ,
         \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 ,
         \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 ,
         \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 ,
         \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 ,
         \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 ,
         \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 ,
         \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 ,
         \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 ,
         \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 ,
         \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 ,
         \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 ,
         \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 ,
         \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 ,
         \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 ,
         \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 ,
         \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 ,
         \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 ,
         \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 ,
         \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 ,
         \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 ,
         \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 ,
         \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 ,
         \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 ,
         \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 ,
         \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 ,
         \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 ,
         \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 ,
         \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 ,
         \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 ,
         \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 ,
         \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 ,
         \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 ,
         \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 ,
         \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 ,
         \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 ,
         \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 ,
         \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 ,
         \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 ,
         \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 ,
         \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 ,
         \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 ,
         \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 ,
         \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 ,
         \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 ,
         \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 ,
         \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 ,
         \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 ,
         \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 ,
         \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 ,
         \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 ,
         \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 ,
         \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 ,
         \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 ,
         \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 ,
         \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 ,
         \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 ,
         \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 ,
         \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 ,
         \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 ,
         \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 ,
         \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 ,
         \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 ,
         \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 ,
         \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 ,
         \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 ,
         \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 ,
         \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 ,
         \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 ,
         \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 ,
         \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 ,
         \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 ,
         \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 ,
         \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 ,
         \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 ,
         \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 ,
         \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 ,
         \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 ,
         \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 ,
         \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 ,
         \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 ,
         \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 ,
         \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 ,
         \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 ,
         \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 ,
         \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 ,
         \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 ,
         \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 ,
         \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 ,
         \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 ,
         \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 ,
         \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 ,
         \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 ,
         \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 ,
         \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 ,
         \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 ,
         \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 ,
         \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 ,
         \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 ,
         \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 ,
         \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 ,
         \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 ,
         \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 ,
         \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 ,
         \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 ,
         \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 ,
         \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 ,
         \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 ,
         \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 ,
         \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 ,
         \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 ,
         \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 ,
         \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 ,
         \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 ,
         \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 ,
         \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 ,
         \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 ,
         \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 ,
         \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 ,
         \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 ,
         \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 ,
         \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 ,
         \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 ,
         \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 ,
         \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 ,
         \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 ,
         \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 ,
         \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 ,
         \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 ,
         \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 ,
         \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 ,
         \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 ,
         \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 ,
         \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 ,
         \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 ,
         \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 ,
         \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 ,
         \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 ,
         \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 ,
         \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 ,
         \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 ,
         \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 ,
         \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 ,
         \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 ,
         \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 ,
         \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 ,
         \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 ,
         \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 ,
         \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 ,
         \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 ,
         \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 ,
         \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 ,
         \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 ,
         \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 ,
         \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 ,
         \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 ,
         \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 ,
         \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 ,
         \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 ,
         \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 ,
         \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 ,
         \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 ,
         \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 ,
         \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 ,
         \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 ,
         \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 ,
         \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 ,
         \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 ,
         \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 ,
         \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 ,
         \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 ,
         \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 ,
         \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 ,
         \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 ,
         \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 ,
         \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 ,
         \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 ,
         \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 ,
         \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 ,
         \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 ,
         \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 ,
         \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 ,
         \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 ,
         \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 ,
         \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 ,
         \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 ,
         \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 ,
         \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 ,
         \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 ,
         \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 ,
         \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 ,
         \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 ,
         \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 ,
         \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 ,
         \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 ,
         \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 ,
         \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 ,
         \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 ,
         \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 ,
         \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 ,
         \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 ,
         \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 ,
         \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 ,
         \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 ,
         \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 ,
         \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 ,
         \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 ,
         \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 ,
         \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 ,
         \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 ,
         \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 ,
         \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 ,
         \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 ,
         \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 ,
         \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 ,
         \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 ,
         \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 ,
         \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 ,
         \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 ,
         \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 ,
         \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 ,
         \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 ,
         \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 ,
         \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 ,
         \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 ,
         \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 ,
         \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 ,
         \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 ,
         \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 ,
         \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 ,
         \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 ,
         \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 ,
         \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 ,
         \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 ,
         \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 ,
         \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 ,
         \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 ,
         \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 ,
         \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 ,
         \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 ,
         \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 ,
         \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 ,
         \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 ,
         \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 ,
         \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 ,
         \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 ,
         \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 ,
         \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 ,
         \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 ,
         \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 ,
         \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 ,
         \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 ,
         \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 ,
         \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 ,
         \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 ,
         \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 ,
         \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 ,
         \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 ,
         \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 ,
         \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 ,
         \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 ,
         \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 ,
         \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 ,
         \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 ,
         \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 ,
         \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 ,
         \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 ,
         \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 ,
         \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 ,
         \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 ,
         \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 ,
         \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 ,
         \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 ,
         \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 ,
         \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 ,
         \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 ,
         \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 ,
         \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 ,
         \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 ,
         \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 ,
         \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 ,
         \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 ,
         \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 ,
         \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 ,
         \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 ,
         \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 ,
         \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 ,
         \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 ,
         \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 ,
         \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 ,
         \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 ,
         \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 ,
         \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 ,
         \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 ,
         \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 ,
         \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 ,
         \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 ,
         \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 ,
         \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 ,
         \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 ,
         \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 ,
         \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 ,
         \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 ,
         \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 ,
         \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 ,
         \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 ,
         \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 ,
         \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 ,
         \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 ,
         \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 ,
         \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 ,
         \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 ,
         \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 ,
         \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 ,
         \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 ,
         \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 ,
         \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 ,
         \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 ,
         \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 ,
         \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 ,
         \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 ,
         \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 ,
         \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 ,
         \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 ,
         \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 ,
         \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 ,
         \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 ,
         \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 ,
         \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 ,
         \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 ,
         \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 ,
         \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 ,
         \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 ,
         \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 ,
         \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 ,
         \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 ,
         \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 ,
         \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 ,
         \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 ,
         \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 ,
         \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 ,
         \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 ,
         \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 ,
         \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 ,
         \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 ,
         \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 ,
         \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 ,
         \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 ,
         \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 ,
         \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 ,
         \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 ,
         \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 ,
         \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 ,
         \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 ,
         \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 ,
         \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 ,
         \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 ,
         \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 ,
         \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 ,
         \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 ,
         \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 ,
         \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 ,
         \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 ,
         \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 ,
         \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 ,
         \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 ,
         \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 ,
         \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 ,
         \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 ,
         \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 ,
         \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 ,
         \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 ,
         \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 ,
         \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 ,
         \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 ,
         \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 ,
         \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 ,
         \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 ,
         \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 ,
         \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 ,
         \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 ,
         \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 ,
         \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 ,
         \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 ,
         \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 ,
         \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 ,
         \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 ,
         \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 ,
         \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 ,
         \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 ,
         \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 ,
         \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 ,
         \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 ,
         \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 ,
         \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 ,
         \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 ,
         \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 ,
         \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 ,
         \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 ,
         \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 ,
         \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 ,
         \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 ,
         \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 ,
         \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 ,
         \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 ,
         \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 ,
         \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 ,
         \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 ,
         \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 ,
         \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 ,
         \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 ,
         \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 ,
         \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 ,
         \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 ,
         \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 ,
         \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 ,
         \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 ,
         \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 ,
         \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 ,
         \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 ,
         \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 ,
         \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 ,
         \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 ,
         \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 ,
         \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 ,
         \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 ,
         \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 ,
         \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 ,
         \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 ,
         \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 ,
         \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 ,
         \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 ,
         \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 ,
         \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 ,
         \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 ,
         \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 ,
         \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 ,
         \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 ,
         \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 ,
         \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 ,
         \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 ,
         \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 ,
         \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 ,
         \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 ,
         \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 ,
         \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 ,
         \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 ,
         \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 ,
         \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 ,
         \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 ,
         \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 ,
         \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 ,
         \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 ,
         \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 ,
         \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 ,
         \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 ,
         \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 ,
         \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 ,
         \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 ,
         \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 ,
         \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 ,
         \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 ,
         \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 ,
         \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 ,
         \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 ,
         \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 ,
         \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 ,
         \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 ,
         \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 ,
         \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 ,
         \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 ,
         \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 ,
         \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 ,
         \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 ,
         \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 ,
         \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 ,
         \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 ,
         \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 ,
         \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 ,
         \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 ,
         \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 ,
         \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 ,
         \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 ,
         \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 ,
         \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 ,
         \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 ,
         \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 ,
         \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 ,
         \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 ,
         \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 ,
         \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 ,
         \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 ,
         \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 ,
         \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 ,
         \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 ,
         \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 ,
         \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 ,
         \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 ,
         \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 ,
         \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 ,
         \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 ,
         \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 ,
         \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 ,
         \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 ,
         \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 ,
         \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 ,
         \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 ,
         \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 ,
         \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 ,
         \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 ,
         \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 ,
         \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 ,
         \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 ,
         \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 ,
         \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 ,
         \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 ,
         \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 ,
         \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 ,
         \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 ,
         \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 ,
         \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 ,
         \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 ,
         \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 ,
         \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 ,
         \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 ,
         \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 ,
         \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 ,
         \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 ,
         \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 ,
         \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 ,
         \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 ,
         \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 ,
         \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 ,
         \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 ,
         \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 ,
         \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 ,
         \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 ,
         \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 ,
         \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 ,
         \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 ,
         \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 ,
         \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 ,
         \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 ,
         \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 ,
         \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 ,
         \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 ,
         \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 ,
         \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 ,
         \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 ,
         \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 ,
         \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 ,
         \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 ,
         \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 ,
         \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 ,
         \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 ,
         \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 ,
         \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 ,
         \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 ,
         \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 ,
         \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 ,
         \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 ,
         \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 ,
         \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 ,
         \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 ,
         \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 ,
         \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 ,
         \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 ,
         \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 ,
         \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 ,
         \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 ,
         \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 ,
         \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 ,
         \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 ,
         \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 ,
         \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 ,
         \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 ,
         \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 ,
         \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 ,
         \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 ,
         \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 ,
         \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 ,
         \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 ,
         \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 ,
         \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 ,
         \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 ,
         \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 ,
         \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 ,
         \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 ,
         \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 ,
         \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 ,
         \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 ,
         \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 ,
         \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 ,
         \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 ,
         \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 ,
         \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 ,
         \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 ,
         \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 ,
         \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 ,
         \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 ,
         \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 ,
         \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 ,
         \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 ,
         \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 ,
         \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 ,
         \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 ,
         \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 ,
         \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 ,
         \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 ,
         \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 ,
         \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 ,
         \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 ,
         \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 ,
         \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 ,
         \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 ,
         \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 ,
         \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 ,
         \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 ,
         \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 ,
         \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 ,
         \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 ,
         \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 ,
         \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 ,
         \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 ,
         \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 ,
         \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 ,
         \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 ,
         \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 ,
         \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 ,
         \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 ,
         \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 ,
         \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 ,
         \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 ,
         \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 ,
         \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 ,
         \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 ,
         \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 ,
         \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 ,
         \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 ,
         \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 ,
         \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 ,
         \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 ,
         \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 ,
         \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 ,
         \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 ,
         \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 ,
         \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 ,
         \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 ,
         \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 ,
         \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 ,
         \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 ,
         \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 ,
         \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 ,
         \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 ,
         \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 ,
         \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 ,
         \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 ,
         \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 ,
         \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 ,
         \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 ,
         \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 ,
         \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 ,
         \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 ,
         \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 ,
         \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 ,
         \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 ,
         \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 ,
         \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 ,
         \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 ,
         \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 ,
         \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 ,
         \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 ,
         \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 ,
         \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 ,
         \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 ,
         \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 ,
         \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 ,
         \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 ,
         \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 ,
         \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 ,
         \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 ,
         \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 ,
         \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 ,
         \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 ,
         \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 ,
         \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 ,
         \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 ,
         \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 ,
         \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 ,
         \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 ,
         \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 ,
         \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 ,
         \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 ,
         \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 ,
         \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 ,
         \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 ,
         \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 ,
         \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 ,
         \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 ,
         \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 ,
         \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 ,
         \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 ,
         \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 ,
         \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 ,
         \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 ,
         \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 ,
         \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 ,
         \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 ,
         \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 ,
         \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 ,
         \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 ,
         \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 ,
         \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 ,
         \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 ,
         \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 ,
         \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 ,
         \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 ,
         \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 ,
         \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 ,
         \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 ,
         \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 ,
         \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 ,
         \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 ,
         \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 ,
         \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 ,
         \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 ,
         \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 ,
         \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 ,
         \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 ,
         \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 ,
         \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 ,
         \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 ,
         \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 ,
         \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 ,
         \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 ,
         \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 ,
         \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 ,
         \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 ,
         \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 ,
         \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 ,
         \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 ,
         \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 ,
         \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 ,
         \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 ,
         \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 ,
         \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 ,
         \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 ,
         \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 ,
         \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 ,
         \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 ,
         \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 ,
         \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 ,
         \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 ,
         \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 ,
         \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 ,
         \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 ,
         \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 ,
         \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 ,
         \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 ,
         \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 ,
         \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 ,
         \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 ,
         \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 ,
         \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 ,
         \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 ,
         \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 ,
         \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 ,
         \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 ,
         \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 ,
         \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 ,
         \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 ,
         \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 ,
         \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 ,
         \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 ,
         \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 ,
         \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 ,
         \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 ,
         \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 ,
         \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 ,
         \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 ,
         \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 ,
         \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 ,
         \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 ,
         \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 ,
         \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 ,
         \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 ,
         \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 ,
         \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 ,
         \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 ,
         \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 ,
         \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 ,
         \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 ,
         \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 ,
         \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 ,
         \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 ,
         \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 ,
         \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 ,
         \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 ,
         \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 ,
         \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 ,
         \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 ,
         \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 ,
         \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 ,
         \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 ,
         \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 ,
         \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 ,
         \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 ,
         \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 ,
         \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 ,
         \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 ,
         \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 ,
         \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 ,
         \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 ,
         \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 ,
         \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 ,
         \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 ,
         \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 ,
         \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 ,
         \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 ,
         \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 ,
         \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 ,
         \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 ,
         \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 ,
         \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 ,
         \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 ,
         \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 ,
         \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 ,
         \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 ,
         \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 ,
         \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 ,
         \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 ,
         \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 ,
         \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 ,
         \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 ,
         \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 ,
         \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 ,
         \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 ,
         \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 ,
         \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 ,
         \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 ,
         \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 ,
         \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 ,
         \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 ,
         \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 ,
         \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 ,
         \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 ,
         \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 ,
         \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 ,
         \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 ,
         \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 ,
         \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 ,
         \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 ,
         \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 ,
         \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 ,
         \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 ,
         \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 ,
         \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 ,
         \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 ,
         \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 ,
         \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 ,
         \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 ,
         \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 ,
         \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 ,
         \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 ,
         \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 ,
         \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 ,
         \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 ,
         \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 ,
         \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 ,
         \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 ,
         \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 ,
         \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 ,
         \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 ,
         \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 ,
         \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 ,
         \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 ,
         \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 ,
         \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 ,
         \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 ,
         \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 ,
         \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 ,
         \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 ,
         \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 ,
         \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 ,
         \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 ,
         \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 ,
         \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 ,
         \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 ,
         \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 ,
         \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 ,
         \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 ,
         \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 ,
         \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 ,
         \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 ,
         \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 ,
         \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 ,
         \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 ,
         \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 ,
         \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 ,
         \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 ,
         \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 ,
         \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 ,
         \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 ,
         \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 ,
         \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 ,
         \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 ,
         \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 ,
         \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 ,
         \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 ,
         \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 ,
         \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 ,
         \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 ,
         \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 ,
         \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 ,
         \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 ,
         \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 ,
         \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 ,
         \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 ,
         \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 ,
         \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 ,
         \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 ,
         \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 ,
         \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 ,
         \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 ,
         \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 ,
         \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 ,
         \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 ,
         \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 ,
         \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 ,
         \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 ,
         \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 ,
         \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 ,
         \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 ,
         \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 ,
         \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 ,
         \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 ,
         \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 ,
         \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 ,
         \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 ,
         \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 ,
         \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 ,
         \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 ,
         \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 ,
         \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 ,
         \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 ,
         \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 ,
         \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 ,
         \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 ,
         \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 ,
         \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 ,
         \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 ,
         \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 ,
         \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 ,
         \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 ,
         \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 ,
         \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 ,
         \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 ,
         \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 ,
         \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 ,
         \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 ,
         \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 ,
         \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 ,
         \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 ,
         \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 ,
         \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 ,
         \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 ,
         \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 ,
         \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 ,
         \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 ,
         \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 ,
         \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 ,
         \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 ,
         \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 ,
         \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 ,
         \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 ,
         \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 ,
         \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 ,
         \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 ,
         \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 ,
         \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 ,
         \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 ,
         \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 ,
         \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 ,
         \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 ,
         \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 ,
         \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 ,
         \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 ,
         \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 ,
         \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 ,
         \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 ,
         \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 ,
         \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 ,
         \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 ,
         \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 ,
         \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 ,
         \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 ,
         \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 ,
         \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 ,
         \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 ,
         \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 ,
         \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 ,
         \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 ,
         \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 ,
         \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 ,
         \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 ,
         \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 ,
         \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 ,
         \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 ,
         \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 ,
         \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 ,
         \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 ,
         \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 ,
         \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 ,
         \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 ,
         \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 ,
         \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 ,
         \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 ,
         \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 ,
         \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 ,
         \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 ,
         \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 ,
         \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 ,
         \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 ,
         \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 ,
         \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 ,
         \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 ,
         \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 ,
         \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 ,
         \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 ,
         \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 ,
         \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 ,
         \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 ,
         \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 ,
         \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 ,
         \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 ,
         \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 ,
         \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 ,
         \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 ,
         \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 ,
         \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 ,
         \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 ,
         \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 ,
         \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 ,
         \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 ,
         \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 ,
         \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 ,
         \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 ,
         \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 ,
         \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 ,
         \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 ,
         \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 ,
         \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 ,
         \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 ,
         \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 ,
         \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 ,
         \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 ,
         \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 ,
         \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 ,
         \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 ,
         \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 ,
         \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 ,
         \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 ,
         \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 ,
         \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 ,
         \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 ,
         \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 ,
         \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 ,
         \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 ,
         \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 ,
         \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 ,
         \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 ,
         \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 ,
         \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 ,
         \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 ,
         \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 ,
         \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 ,
         \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 ,
         \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 ,
         \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 ,
         \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 ,
         \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 ,
         \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 ,
         \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 ,
         \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 ,
         \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 ,
         \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 ,
         \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 ,
         \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 ,
         \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 ,
         \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 ,
         \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 ,
         \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 ,
         \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 ,
         \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 ,
         \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 ,
         \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 ,
         \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 ,
         \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 ,
         \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 ,
         \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 ,
         \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 ,
         \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 ,
         \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 ,
         \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 ,
         \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 ,
         \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 ,
         \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 ,
         \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 ,
         \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 ,
         \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 ,
         \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 ,
         \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 ,
         \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 ,
         \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 ,
         \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 ,
         \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 ,
         \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 ,
         \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 ,
         \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 ,
         \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 ,
         \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 ,
         \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 ,
         \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 ,
         \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 ,
         \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 ,
         \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 ,
         \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 ,
         \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 ,
         \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 ,
         \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 ,
         \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 ,
         \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 ,
         \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 ,
         \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 ,
         \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 ,
         \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 ,
         \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 ,
         \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 ,
         \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 ,
         \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 ,
         \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 ,
         \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 ,
         \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 ,
         \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 ,
         \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 ,
         \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 ,
         \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 ,
         \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 ,
         \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 ,
         \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 ,
         \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 ,
         \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 ,
         \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 ,
         \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 ,
         \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 ,
         \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 ,
         \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 ,
         \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 ,
         \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 ,
         \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 ,
         \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 ,
         \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 ,
         \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 ,
         \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 ,
         \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 ,
         \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 ,
         \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 ,
         \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 ,
         \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 ,
         \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 ,
         \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 ,
         \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 ,
         \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 ,
         \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 ,
         \16261 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 ,
         \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 ,
         \16281 , \16282 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 ,
         \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 ,
         \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 ,
         \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 ,
         \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 ,
         \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 ,
         \16341 , \16342 , \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 ,
         \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 ,
         \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 ,
         \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 ,
         \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 ,
         \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 ,
         \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 ,
         \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 ,
         \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 ,
         \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 ,
         \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 ,
         \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 ,
         \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 ,
         \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 ,
         \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 ,
         \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 ,
         \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 ,
         \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 ,
         \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 ,
         \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 ,
         \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 ,
         \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 ,
         \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 ,
         \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 ,
         \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 ,
         \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 ,
         \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 ,
         \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 ,
         \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 ,
         \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 ,
         \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 ,
         \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 ,
         \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 ,
         \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 ,
         \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 ,
         \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 ,
         \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 ,
         \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 ,
         \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 ,
         \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 ,
         \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 ,
         \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 ,
         \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 ,
         \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 ,
         \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 ,
         \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 ,
         \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 ,
         \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 ,
         \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 ,
         \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 ,
         \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 ,
         \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 ,
         \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 ,
         \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 ,
         \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 ,
         \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 ,
         \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 ,
         \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 ,
         \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 ,
         \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 ,
         \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 ,
         \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 ,
         \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 ,
         \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 ,
         \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 ,
         \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 ,
         \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 ,
         \17011 , \17012 , \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 ,
         \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 ,
         \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 ,
         \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 ,
         \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 ,
         \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 ,
         \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 ,
         \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 ,
         \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 ,
         \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 ,
         \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 ,
         \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 ,
         \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 ,
         \17141 , \17142 , \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 ,
         \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 ,
         \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 ,
         \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 ,
         \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 ,
         \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 ,
         \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 ,
         \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 ,
         \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 ,
         \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 ,
         \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 ,
         \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 ,
         \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 ,
         \17271 , \17272 , \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 ,
         \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 ,
         \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 ,
         \17301 , \17302 , \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 ,
         \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 ,
         \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 ,
         \17331 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 ,
         \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 ,
         \17351 , \17352 , \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 ,
         \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 ,
         \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 ,
         \17381 , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 ,
         \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 ,
         \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 ,
         \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 ,
         \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 ,
         \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 ,
         \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 ,
         \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 ,
         \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 ,
         \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 ,
         \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 ,
         \17491 , \17492 , \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 ,
         \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 ,
         \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 ,
         \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 ,
         \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 ,
         \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 ,
         \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 ,
         \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 ,
         \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 ,
         \17581 , \17582 , \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 ,
         \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 ,
         \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 ,
         \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 ,
         \17621 , \17622 , \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 ,
         \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 ,
         \17641 , \17642 , \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 ,
         \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 ,
         \17661 , \17662 , \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 ,
         \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 ,
         \17681 , \17682 , \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 ,
         \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 ,
         \17701 , \17702 , \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 ,
         \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 ,
         \17721 , \17722 , \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 ,
         \17731 , \17732 , \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 ,
         \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 ,
         \17751 , \17752 , \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 ,
         \17761 , \17762 , \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 ,
         \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 ,
         \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 ,
         \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 ,
         \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 ,
         \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 ,
         \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 ,
         \17831 , \17832 , \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 ,
         \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 ,
         \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 ,
         \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 ,
         \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 ,
         \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 ,
         \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 ,
         \17901 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 ,
         \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 ,
         \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 ,
         \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 ,
         \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 ,
         \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 ,
         \17961 , \17962 , \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 ,
         \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 ,
         \17981 , \17982 , \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 ,
         \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 ,
         \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 ,
         \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 ,
         \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 ,
         \18031 , \18032 , \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 ,
         \18041 , \18042 , \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 ,
         \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 ,
         \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 ,
         \18071 , \18072 , \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 ,
         \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 ,
         \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 ,
         \18101 , \18102 , \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 ,
         \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 ,
         \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 ,
         \18131 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 ,
         \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 ,
         \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 ,
         \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 ,
         \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 ,
         \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 ,
         \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 ,
         \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 ,
         \18211 , \18212 , \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 ,
         \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 ,
         \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 ,
         \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 ,
         \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 ,
         \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 ,
         \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 ,
         \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 ,
         \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 ,
         \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 ,
         \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 ,
         \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 ,
         \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 ,
         \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 ,
         \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 ,
         \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 ,
         \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 ,
         \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 ,
         \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 ,
         \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 ,
         \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 ,
         \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 ,
         \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 ,
         \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 ,
         \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 ,
         \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 ,
         \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 ,
         \18481 , \18482 , \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 ,
         \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 ,
         \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 ,
         \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 ,
         \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 ,
         \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 ,
         \18541 , \18542 , \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 ,
         \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 ,
         \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 ,
         \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 ,
         \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 ,
         \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 ,
         \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 ,
         \18611 , \18612 , \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 ,
         \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 ,
         \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 ,
         \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 ,
         \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 ,
         \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 ,
         \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 ,
         \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 ,
         \18691 , \18692 , \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 ,
         \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 ,
         \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 ,
         \18721 , \18722 , \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 ,
         \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 ,
         \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 ,
         \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 ,
         \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 ,
         \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 ,
         \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 ,
         \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 ,
         \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 ,
         \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 ,
         \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 ,
         \18831 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 ,
         \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 ,
         \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 ,
         \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 ,
         \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 ,
         \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 ,
         \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 ,
         \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 ,
         \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 ,
         \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 ,
         \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 ,
         \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 ,
         \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 ,
         \18961 , \18962 , \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 ,
         \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 ,
         \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 ,
         \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 ,
         \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 ,
         \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 ,
         \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 ,
         \19031 , \19032 , \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 ,
         \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 ,
         \19051 , \19052 , \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 ,
         \19061 , \19062 , \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 ,
         \19071 , \19072 , \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 ,
         \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 ,
         \19091 , \19092 , \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 ,
         \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 ,
         \19111 , \19112 , \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 ,
         \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 ,
         \19131 , \19132 , \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 ,
         \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 ,
         \19151 , \19152 , \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 ,
         \19161 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 ,
         \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 ,
         \19181 , \19182 , \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 ,
         \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 ,
         \19201 , \19202 , \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 ,
         \19211 , \19212 , \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 ,
         \19221 , \19222 , \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 ,
         \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 ,
         \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 ,
         \19251 , \19252 , \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 ,
         \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 ,
         \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 ,
         \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 ,
         \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 ,
         \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 ,
         \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 ,
         \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 ,
         \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 ,
         \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 ,
         \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 ,
         \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 ,
         \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 ,
         \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 ,
         \19391 , \19392 , \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 ,
         \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 ,
         \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 ,
         \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 ,
         \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 ,
         \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 ,
         \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 ,
         \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 ,
         \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 ,
         \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 ,
         \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 ,
         \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 ,
         \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 ,
         \19521 , \19522 , \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 ,
         \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 ,
         \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 ,
         \19551 , \19552 , \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 ,
         \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 ,
         \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 ,
         \19581 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 ,
         \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 ,
         \19601 , \19602 , \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 ,
         \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 ,
         \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 ,
         \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 ,
         \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 ,
         \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 ,
         \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 ,
         \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 ,
         \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 ,
         \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 ,
         \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 ,
         \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 ,
         \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 ,
         \19731 , \19732 , \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 ,
         \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 ,
         \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 ,
         \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 ,
         \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 ,
         \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 ,
         \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 ,
         \19801 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 ,
         \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 ,
         \19821 , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 ,
         \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 ,
         \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 ,
         \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 ,
         \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 ,
         \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 ,
         \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 ,
         \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 ,
         \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 ,
         \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 ,
         \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 ,
         \19931 , \19932 , \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 ,
         \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 ,
         \19951 , \19952 , \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 ,
         \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 ,
         \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 ,
         \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 ,
         \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 ,
         \20001 , \20002 , \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 ,
         \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 ,
         \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 ,
         \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 ,
         \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 ,
         \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 ,
         \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 ,
         \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 ,
         \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 ,
         \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 ,
         \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 ,
         \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 ,
         \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 ,
         \20131 , \20132 , \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 ,
         \20141 , \20142 , \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 ,
         \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 ,
         \20161 , \20162 , \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 ,
         \20171 , \20172 , \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 ,
         \20181 , \20182 , \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 ,
         \20191 , \20192 , \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 ,
         \20201 , \20202 , \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 ,
         \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 ,
         \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 ,
         \20231 , \20232 , \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 ,
         \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 ,
         \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 ,
         \20261 , \20262 , \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 ,
         \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 ,
         \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 ,
         \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 ,
         \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 ,
         \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 ,
         \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 ,
         \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 ,
         \20341 , \20342 , \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 ,
         \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 ,
         \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 ,
         \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 ,
         \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 ,
         \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 ,
         \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 ,
         \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 ,
         \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 ,
         \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 ,
         \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 ,
         \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 ,
         \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 ,
         \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 ,
         \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 ,
         \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 ,
         \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 ,
         \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 ,
         \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 ,
         \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 ,
         \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 ,
         \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 ,
         \20561 , \20562 , \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 ,
         \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 ,
         \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 ,
         \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 ,
         \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 ,
         \20611 , \20612 , \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 ,
         \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 ,
         \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 ,
         \20641 , \20642 , \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 ,
         \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 ,
         \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 ,
         \20671 , \20672 , \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 ,
         \20681 , \20682 , \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 ,
         \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 ,
         \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 ,
         \20711 , \20712 , \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 ,
         \20721 , \20722 , \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 ,
         \20731 , \20732 , \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 ,
         \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 ,
         \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 ,
         \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 ,
         \20771 , \20772 , \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 ,
         \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 ,
         \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 ,
         \20801 , \20802 , \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 ,
         \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 ,
         \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 ,
         \20831 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 ,
         \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 ,
         \20851 , \20852 , \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 ,
         \20861 , \20862 , \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 ,
         \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 ,
         \20881 , \20882 , \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 ,
         \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 ,
         \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 ,
         \20911 , \20912 , \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 ,
         \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 ,
         \20931 , \20932 , \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 ,
         \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 ,
         \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 ,
         \20961 , \20962 , \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 ,
         \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 ,
         \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 ,
         \20991 , \20992 , \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 ,
         \21001 , \21002 , \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 ,
         \21011 , \21012 , \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 ,
         \21021 , \21022 , \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 ,
         \21031 , \21032 , \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 ,
         \21041 , \21042 , \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 ,
         \21051 , \21052 , \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 ,
         \21061 , \21062 , \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 ,
         \21071 , \21072 , \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 ,
         \21081 , \21082 , \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 ,
         \21091 , \21092 , \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 ,
         \21101 , \21102 , \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 ,
         \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 ,
         \21121 , \21122 , \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 ,
         \21131 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 ,
         \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 ,
         \21151 , \21152 , \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 ,
         \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 ,
         \21171 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 ,
         \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 ,
         \21191 , \21192 , \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 ,
         \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 ,
         \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 ,
         \21221 , \21222 , \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 ,
         \21231 , \21232 , \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 ,
         \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 ,
         \21251 , \21252 , \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 ,
         \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 ,
         \21271 , \21272 , \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 ,
         \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 ,
         \21291 , \21292 , \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 ,
         \21301 , \21302 , \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 ,
         \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 ,
         \21321 , \21322 , \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 ,
         \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 ,
         \21341 , \21342 , \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 ,
         \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 ,
         \21361 , \21362 , \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370 ,
         \21371 , \21372 , \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 ,
         \21381 , \21382 , \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 ,
         \21391 , \21392 , \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 ,
         \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 ,
         \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 ,
         \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 ,
         \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 ,
         \21441 , \21442 , \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 ,
         \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 ,
         \21461 , \21462 , \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 ,
         \21471 , \21472 , \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 ,
         \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 ,
         \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 ,
         \21501 , \21502 , \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 ,
         \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 ,
         \21521 , \21522 , \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 ,
         \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 ,
         \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 ,
         \21551 , \21552 , \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 ,
         \21561 , \21562 , \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 ,
         \21571 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 ,
         \21581 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 ,
         \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 ,
         \21601 , \21602 , \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 ,
         \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 ,
         \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 ,
         \21631 , \21632 , \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 ,
         \21641 , \21642 , \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 ,
         \21651 , \21652 , \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 ,
         \21661 , \21662 , \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 ,
         \21671 , \21672 , \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 ,
         \21681 , \21682 , \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 ,
         \21691 , \21692 , \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 ,
         \21701 , \21702 , \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 ,
         \21711 , \21712 , \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 ,
         \21721 , \21722 , \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 ,
         \21731 , \21732 , \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 ,
         \21741 , \21742 , \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 ,
         \21751 , \21752 , \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 ,
         \21761 , \21762 , \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 ,
         \21771 , \21772 , \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 ,
         \21781 , \21782 , \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 ,
         \21791 , \21792 , \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 ,
         \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 ,
         \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 ,
         \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 ,
         \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 ,
         \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 ,
         \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 ,
         \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 ,
         \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 ,
         \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 ,
         \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 ,
         \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 ,
         \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 ,
         \21921 , \21922 , \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 ,
         \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 ,
         \21941 , \21942 , \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 ,
         \21951 , \21952 , \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 ,
         \21961 , \21962 , \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 ,
         \21971 , \21972 , \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 ,
         \21981 , \21982 , \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 ,
         \21991 , \21992 , \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 ,
         \22001 , \22002 , \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 ,
         \22011 , \22012 , \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 ,
         \22021 , \22022 , \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 ,
         \22031 , \22032 , \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 ,
         \22041 , \22042 , \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 ,
         \22051 , \22052 , \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 ,
         \22061 , \22062 , \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 ,
         \22071 , \22072 , \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 ,
         \22081 , \22082 , \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 ,
         \22091 , \22092 , \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 ,
         \22101 , \22102 , \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 ,
         \22111 , \22112 , \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 ,
         \22121 , \22122 , \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 ,
         \22131 , \22132 , \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 ,
         \22141 , \22142 , \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 ,
         \22151 , \22152 , \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 ,
         \22161 , \22162 , \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 ,
         \22171 , \22172 , \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 ,
         \22181 , \22182 , \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 ,
         \22191 , \22192 , \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 ,
         \22201 , \22202 , \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 ,
         \22211 , \22212 , \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 ,
         \22221 , \22222 , \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 ,
         \22231 , \22232 , \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 ,
         \22241 , \22242 , \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 ,
         \22251 , \22252 , \22253 , \22254 , \22255 , \22256 , \22257 , \22258 , \22259 , \22260 ,
         \22261 , \22262 , \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , \22269 , \22270 ,
         \22271 , \22272 , \22273 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 ,
         \22281 , \22282 , \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 ,
         \22291 , \22292 , \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 ,
         \22301 , \22302 , \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 ,
         \22311 , \22312 , \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 ,
         \22321 , \22322 , \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 ,
         \22331 , \22332 , \22333 , \22334 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 ,
         \22341 , \22342 , \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 ,
         \22351 , \22352 , \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 ,
         \22361 , \22362 , \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 ,
         \22371 , \22372 , \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 ,
         \22381 , \22382 , \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 ,
         \22391 , \22392 , \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 ,
         \22401 , \22402 , \22403 , \22404 , \22405 , \22406 , \22407 , \22408 , \22409 , \22410 ,
         \22411 , \22412 , \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 ,
         \22421 , \22422 , \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 ,
         \22431 , \22432 , \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 ,
         \22441 , \22442 , \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 ,
         \22451 , \22452 , \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 ,
         \22461 , \22462 , \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 , \22470 ,
         \22471 , \22472 , \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 ,
         \22481 , \22482 , \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 ,
         \22491 , \22492 , \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 ,
         \22501 , \22502 , \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 ,
         \22511 , \22512 , \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 ,
         \22521 , \22522 , \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 ,
         \22531 , \22532 , \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 ,
         \22541 , \22542 , \22543 , \22544 , \22545 , \22546 , \22547 , \22548 , \22549 , \22550 ,
         \22551 , \22552 , \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 ,
         \22561 , \22562 , \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 ,
         \22571 , \22572 , \22573 , \22574 , \22575 , \22576 , \22577 , \22578 , \22579 , \22580 ,
         \22581 , \22582 , \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 ,
         \22591 , \22592 , \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 ,
         \22601 , \22602 , \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 ,
         \22611 , \22612 , \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 ,
         \22621 , \22622 , \22623 , \22624 , \22625 , \22626 , \22627 , \22628 , \22629 , \22630 ,
         \22631 , \22632 , \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 ,
         \22641 , \22642 , \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 ,
         \22651 , \22652 , \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 ,
         \22661 , \22662 , \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 ,
         \22671 , \22672 , \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 ,
         \22681 , \22682 , \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 ,
         \22691 , \22692 , \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 ,
         \22701 , \22702 , \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 ,
         \22711 , \22712 , \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 ,
         \22721 , \22722 , \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 ,
         \22731 , \22732 , \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 ,
         \22741 , \22742 , \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 ,
         \22751 , \22752 , \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 ,
         \22761 , \22762 , \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 ,
         \22771 , \22772 , \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 ,
         \22781 , \22782 , \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 ,
         \22791 , \22792 , \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 ,
         \22801 , \22802 , \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 ,
         \22811 , \22812 , \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 ,
         \22821 , \22822 , \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 ,
         \22831 , \22832 , \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 ,
         \22841 , \22842 , \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 ,
         \22851 , \22852 , \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 ,
         \22861 , \22862 , \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 ,
         \22871 , \22872 , \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 ,
         \22881 , \22882 , \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 ,
         \22891 , \22892 , \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 ,
         \22901 , \22902 , \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 ,
         \22911 , \22912 , \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 ,
         \22921 , \22922 , \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 ,
         \22931 , \22932 , \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 ,
         \22941 , \22942 , \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 ,
         \22951 , \22952 , \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 ,
         \22961 , \22962 , \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 ,
         \22971 , \22972 , \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 ,
         \22981 , \22982 , \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 ,
         \22991 , \22992 , \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 ,
         \23001 , \23002 , \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 ,
         \23011 , \23012 , \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 ,
         \23021 , \23022 , \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 ,
         \23031 , \23032 , \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 ,
         \23041 , \23042 , \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 ,
         \23051 , \23052 , \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 ,
         \23061 , \23062 , \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 ,
         \23071 , \23072 , \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 ,
         \23081 , \23082 , \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 ,
         \23091 , \23092 , \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 ,
         \23101 , \23102 , \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 ,
         \23111 , \23112 , \23113 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 ,
         \23121 , \23122 , \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 ,
         \23131 , \23132 , \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 ,
         \23141 , \23142 , \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 ,
         \23151 , \23152 , \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 ,
         \23161 , \23162 , \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 ,
         \23171 , \23172 , \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 ,
         \23181 , \23182 , \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 ,
         \23191 , \23192 , \23193 , \23194 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 ,
         \23201 , \23202 , \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 ,
         \23211 , \23212 , \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 , \23220 ,
         \23221 , \23222 , \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 ,
         \23231 , \23232 , \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 ,
         \23241 , \23242 , \23243 , \23244 , \23245 , \23246 , \23247 , \23248 , \23249 , \23250 ,
         \23251 , \23252 , \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 ,
         \23261 , \23262 , \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 ,
         \23271 , \23272 , \23273 , \23274 , \23275 , \23276 , \23277 , \23278 , \23279 , \23280 ,
         \23281 , \23282 , \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 ,
         \23291 , \23292 , \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 ,
         \23301 , \23302 , \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 ,
         \23311 , \23312 , \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 ,
         \23321 , \23322 , \23323 , \23324 , \23325 , \23326 , \23327 , \23328 , \23329 , \23330 ,
         \23331 , \23332 , \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 ,
         \23341 , \23342 , \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 ,
         \23351 , \23352 , \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 ,
         \23361 , \23362 , \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 ,
         \23371 , \23372 , \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 ,
         \23381 , \23382 , \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 ,
         \23391 , \23392 , \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 ,
         \23401 , \23402 , \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 ,
         \23411 , \23412 , \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 ,
         \23421 , \23422 , \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 ,
         \23431 , \23432 , \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 ,
         \23441 , \23442 , \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 ,
         \23451 , \23452 , \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 ,
         \23461 , \23462 , \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 ,
         \23471 , \23472 , \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 ,
         \23481 , \23482 , \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 ,
         \23491 , \23492 , \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 ,
         \23501 , \23502 , \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 ,
         \23511 , \23512 , \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 ,
         \23521 , \23522 , \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 ,
         \23531 , \23532 , \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 ,
         \23541 , \23542 , \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 ,
         \23551 , \23552 , \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 ,
         \23561 , \23562 , \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 ,
         \23571 , \23572 , \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 ,
         \23581 , \23582 , \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 ,
         \23591 , \23592 , \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 ,
         \23601 , \23602 , \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 ,
         \23611 , \23612 , \23613 , \23614 , \23615 , \23616 , \23617 , \23618 , \23619 , \23620 ,
         \23621 , \23622 , \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 ,
         \23631 , \23632 , \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 ,
         \23641 , \23642 , \23643 , \23644 , \23645 , \23646 , \23647 , \23648 , \23649 , \23650 ,
         \23651 , \23652 , \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 ,
         \23661 , \23662 , \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 ,
         \23671 , \23672 , \23673 , \23674 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 ,
         \23681 , \23682 , \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 ,
         \23691 , \23692 , \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 , \23700 ,
         \23701 , \23702 , \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 ,
         \23711 , \23712 , \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 ,
         \23721 , \23722 , \23723 , \23724 , \23725 , \23726 , \23727 , \23728 , \23729 , \23730 ,
         \23731 , \23732 , \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 ,
         \23741 , \23742 , \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 ,
         \23751 , \23752 , \23753 , \23754 , \23755 , \23756 , \23757 , \23758 , \23759 , \23760 ,
         \23761 , \23762 , \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 ,
         \23771 , \23772 , \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 ,
         \23781 , \23782 , \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 ,
         \23791 , \23792 , \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 ,
         \23801 , \23802 , \23803 , \23804 , \23805 , \23806 , \23807 , \23808 , \23809 , \23810 ,
         \23811 , \23812 , \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 ,
         \23821 , \23822 , \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 ,
         \23831 , \23832 , \23833 , \23834 , \23835 , \23836 , \23837 , \23838 , \23839 , \23840 ,
         \23841 , \23842 , \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 ,
         \23851 , \23852 , \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 ,
         \23861 , \23862 , \23863 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 ,
         \23871 , \23872 , \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 ,
         \23881 , \23882 , \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 ,
         \23891 , \23892 , \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 ,
         \23901 , \23902 , \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 ,
         \23911 , \23912 , \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 ,
         \23921 , \23922 , \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 ,
         \23931 , \23932 , \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 ,
         \23941 , \23942 , \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 ,
         \23951 , \23952 , \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 ,
         \23961 , \23962 , \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 ,
         \23971 , \23972 , \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 ,
         \23981 , \23982 , \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 ,
         \23991 , \23992 , \23993 , \23994 , \23995 , \23996 , \23997 , \23998 , \23999 , \24000 ,
         \24001 , \24002 , \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 ,
         \24011 , \24012 , \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 ,
         \24021 , \24022 , \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 ,
         \24031 , \24032 , \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 ,
         \24041 , \24042 , \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 ,
         \24051 , \24052 , \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 ,
         \24061 , \24062 , \24063 , \24064 , \24065 , \24066 , \24067 , \24068 , \24069 , \24070 ,
         \24071 , \24072 , \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 ,
         \24081 , \24082 , \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 ,
         \24091 , \24092 , \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 ,
         \24101 , \24102 , \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 ,
         \24111 , \24112 , \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 ,
         \24121 , \24122 , \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 ,
         \24131 , \24132 , \24133 , \24134 , \24135 , \24136 , \24137 , \24138 , \24139 , \24140 ,
         \24141 , \24142 , \24143 , \24144 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 ,
         \24151 , \24152 , \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 ,
         \24161 , \24162 , \24163 , \24164 , \24165 , \24166 , \24167 , \24168 , \24169 , \24170 ,
         \24171 , \24172 , \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 ,
         \24181 , \24182 , \24183 , \24184 , \24185 , \24186 , \24187 , \24188 , \24189 , \24190 ,
         \24191 , \24192 , \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 ,
         \24201 , \24202 , \24203 , \24204 , \24205 , \24206 , \24207 , \24208 , \24209 , \24210 ,
         \24211 , \24212 , \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 ,
         \24221 , \24222 , \24223 , \24224 , \24225 , \24226 , \24227 , \24228 , \24229 , \24230 ,
         \24231 , \24232 , \24233 , \24234 , \24235 , \24236 , \24237 , \24238 , \24239 , \24240 ,
         \24241 , \24242 , \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 ,
         \24251 , \24252 , \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 ,
         \24261 , \24262 , \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 ,
         \24271 , \24272 , \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 ,
         \24281 , \24282 , \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 ,
         \24291 , \24292 , \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 ,
         \24301 , \24302 , \24303 , \24304 , \24305 , \24306 , \24307 , \24308 , \24309 , \24310 ,
         \24311 , \24312 , \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 ,
         \24321 , \24322 , \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 ,
         \24331 , \24332 , \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 ,
         \24341 , \24342 , \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 ,
         \24351 , \24352 , \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 ,
         \24361 , \24362 , \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 , \24370 ,
         \24371 , \24372 , \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 ,
         \24381 , \24382 , \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 ,
         \24391 , \24392 , \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 ,
         \24401 , \24402 , \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 ,
         \24411 , \24412 , \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 ,
         \24421 , \24422 , \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 ,
         \24431 , \24432 , \24433 , \24434 , \24435 , \24436 , \24437 , \24438 , \24439 , \24440 ,
         \24441 , \24442 , \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 ,
         \24451 , \24452 , \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 ,
         \24461 , \24462 , \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 ,
         \24471 , \24472 , \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 ,
         \24481 , \24482 , \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 ,
         \24491 , \24492 , \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 ,
         \24501 , \24502 , \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , \24509 , \24510 ,
         \24511 , \24512 , \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 ,
         \24521 , \24522 , \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 ,
         \24531 , \24532 , \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 ,
         \24541 , \24542 , \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 ,
         \24551 , \24552 , \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 ,
         \24561 , \24562 , \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 ,
         \24571 , \24572 , \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 ,
         \24581 , \24582 , \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 ,
         \24591 , \24592 , \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 ,
         \24601 , \24602 , \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 ,
         \24611 , \24612 , \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 ,
         \24621 , \24622 , \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 ,
         \24631 , \24632 , \24633 , \24634 , \24635 , \24636 , \24637 , \24638 , \24639 , \24640 ,
         \24641 , \24642 , \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 ,
         \24651 , \24652 , \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 ,
         \24661 , \24662 , \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 ,
         \24671 , \24672 , \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 ,
         \24681 , \24682 , \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 ,
         \24691 , \24692 , \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 ,
         \24701 , \24702 , \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 ,
         \24711 , \24712 , \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 ,
         \24721 , \24722 , \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 ,
         \24731 , \24732 , \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 ,
         \24741 , \24742 , \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 ,
         \24751 , \24752 , \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 ,
         \24761 , \24762 , \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 ,
         \24771 , \24772 , \24773 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 ,
         \24781 , \24782 , \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 ,
         \24791 , \24792 , \24793 , \24794 , \24795 , \24796 , \24797 , \24798 , \24799 , \24800 ,
         \24801 , \24802 , \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 ,
         \24811 , \24812 , \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 ,
         \24821 , \24822 , \24823 , \24824 , \24825 , \24826 , \24827 , \24828 , \24829 , \24830 ,
         \24831 , \24832 , \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 ,
         \24841 , \24842 , \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 ,
         \24851 , \24852 , \24853 , \24854 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 ,
         \24861 , \24862 , \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 ,
         \24871 , \24872 , \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 , \24880 ,
         \24881 , \24882 , \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 ,
         \24891 , \24892 , \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 ,
         \24901 , \24902 , \24903 , \24904 , \24905 , \24906 , \24907 , \24908 , \24909 , \24910 ,
         \24911 , \24912 , \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 ,
         \24921 , \24922 , \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 ,
         \24931 , \24932 , \24933 , \24934 , \24935 , \24936 , \24937 , \24938 , \24939 , \24940 ,
         \24941 , \24942 , \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 ,
         \24951 , \24952 , \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 ,
         \24961 , \24962 , \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 ,
         \24971 , \24972 , \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 ,
         \24981 , \24982 , \24983 , \24984 , \24985 , \24986 , \24987 , \24988 , \24989 , \24990 ,
         \24991 , \24992 , \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 ,
         \25001 , \25002 , \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 ,
         \25011 , \25012 , \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 ,
         \25021 , \25022 , \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 ,
         \25031 , \25032 , \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 ,
         \25041 , \25042 , \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 ,
         \25051 , \25052 , \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 ,
         \25061 , \25062 , \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 ,
         \25071 , \25072 , \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 ,
         \25081 , \25082 , \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 ,
         \25091 , \25092 , \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 ,
         \25101 , \25102 , \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 ,
         \25111 , \25112 , \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 ,
         \25121 , \25122 , \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 ,
         \25131 , \25132 , \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 ,
         \25141 , \25142 , \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 ,
         \25151 , \25152 , \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 ,
         \25161 , \25162 , \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 ,
         \25171 , \25172 , \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 ,
         \25181 , \25182 , \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 ,
         \25191 , \25192 , \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 ,
         \25201 , \25202 , \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 ,
         \25211 , \25212 , \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 ,
         \25221 , \25222 , \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 ,
         \25231 , \25232 , \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 ,
         \25241 , \25242 , \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 ,
         \25251 , \25252 , \25253 , \25254 , \25255 , \25256 , \25257 , \25258 , \25259 , \25260 ,
         \25261 , \25262 , \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 ,
         \25271 , \25272 , \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 ,
         \25281 , \25282 , \25283 , \25284 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 ,
         \25291 , \25292 , \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 ,
         \25301 , \25302 , \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 , \25310 ,
         \25311 , \25312 , \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 ,
         \25321 , \25322 , \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 ,
         \25331 , \25332 , \25333 , \25334 , \25335 , \25336 , \25337 , \25338 , \25339 , \25340 ,
         \25341 , \25342 , \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 ,
         \25351 , \25352 , \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 ,
         \25361 , \25362 , \25363 , \25364 , \25365 , \25366 , \25367 , \25368 , \25369 , \25370 ,
         \25371 , \25372 , \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 ,
         \25381 , \25382 , \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 ,
         \25391 , \25392 , \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 ,
         \25401 , \25402 , \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 ,
         \25411 , \25412 , \25413 , \25414 , \25415 , \25416 , \25417 , \25418 , \25419 , \25420 ,
         \25421 , \25422 , \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 ,
         \25431 , \25432 , \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 ,
         \25441 , \25442 , \25443 , \25444 , \25445 , \25446 , \25447 , \25448 , \25449 , \25450 ,
         \25451 , \25452 , \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 ,
         \25461 , \25462 , \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 ,
         \25471 , \25472 , \25473 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 ,
         \25481 , \25482 , \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 ,
         \25491 , \25492 , \25493 , \25494 , \25495 , \25496 , \25497 , \25498 , \25499 , \25500 ,
         \25501 , \25502 , \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 ,
         \25511 , \25512 , \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 ,
         \25521 , \25522 , \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 ,
         \25531 , \25532 , \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 ,
         \25541 , \25542 , \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 ,
         \25551 , \25552 , \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 ,
         \25561 , \25562 , \25563 , \25564 , \25565 , \25566 , \25567 , \25568 , \25569 , \25570 ,
         \25571 , \25572 , \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 ,
         \25581 , \25582 , \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 ,
         \25591 , \25592 , \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 ,
         \25601 , \25602 , \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 ,
         \25611 , \25612 , \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 ,
         \25621 , \25622 , \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 ,
         \25631 , \25632 , \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 ,
         \25641 , \25642 , \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 ,
         \25651 , \25652 , \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 ,
         \25661 , \25662 , \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 ,
         \25671 , \25672 , \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 ,
         \25681 , \25682 , \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 ,
         \25691 , \25692 , \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 ,
         \25701 , \25702 , \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 ,
         \25711 , \25712 , \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 ,
         \25721 , \25722 , \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 ,
         \25731 , \25732 , \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 ,
         \25741 , \25742 , \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 ,
         \25751 , \25752 , \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 ,
         \25761 , \25762 , \25763 , \25764 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 ,
         \25771 , \25772 , \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 ,
         \25781 , \25782 , \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 , \25790 ,
         \25791 , \25792 , \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 ,
         \25801 , \25802 , \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 ,
         \25811 , \25812 , \25813 , \25814 , \25815 , \25816 , \25817 , \25818 , \25819 , \25820 ,
         \25821 , \25822 , \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 ,
         \25831 , \25832 , \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 ,
         \25841 , \25842 , \25843 , \25844 , \25845 , \25846 , \25847 , \25848 , \25849 , \25850 ,
         \25851 , \25852 , \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 ,
         \25861 , \25862 , \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 ,
         \25871 , \25872 , \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 ,
         \25881 , \25882 , \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 ,
         \25891 , \25892 , \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 ,
         \25901 , \25902 , \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 ,
         \25911 , \25912 , \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 ,
         \25921 , \25922 , \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 ,
         \25931 , \25932 , \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 ,
         \25941 , \25942 , \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 ,
         \25951 , \25952 , \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 ,
         \25961 , \25962 , \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 ,
         \25971 , \25972 , \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 ,
         \25981 , \25982 , \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 ,
         \25991 , \25992 , \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 ,
         \26001 , \26002 , \26003 , \26004 , \26005 , \26006 , \26007 , \26008 , \26009 , \26010 ,
         \26011 , \26012 , \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 ,
         \26021 , \26022 , \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 ,
         \26031 , \26032 , \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 ,
         \26041 , \26042 , \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 ,
         \26051 , \26052 , \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 ,
         \26061 , \26062 , \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 ,
         \26071 , \26072 , \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 ,
         \26081 , \26082 , \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 ,
         \26091 , \26092 , \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 ,
         \26101 , \26102 , \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 ,
         \26111 , \26112 , \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 ,
         \26121 , \26122 , \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 ,
         \26131 , \26132 , \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 ,
         \26141 , \26142 , \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 ,
         \26151 , \26152 , \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 ,
         \26161 , \26162 , \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 ,
         \26171 , \26172 , \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 ,
         \26181 , \26182 , \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 ,
         \26191 , \26192 , \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 ,
         \26201 , \26202 , \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 ,
         \26211 , \26212 , \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 ,
         \26221 , \26222 , \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 ,
         \26231 , \26232 , \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 ,
         \26241 , \26242 , \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 ,
         \26251 , \26252 , \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 ,
         \26261 , \26262 , \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 ,
         \26271 , \26272 , \26273 , \26274 , \26275 , \26276 , \26277 , \26278 , \26279 , \26280 ,
         \26281 , \26282 , \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 ,
         \26291 , \26292 , \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 ,
         \26301 , \26302 , \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 ,
         \26311 , \26312 , \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 ,
         \26321 , \26322 , \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 ,
         \26331 , \26332 , \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 ,
         \26341 , \26342 , \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 ,
         \26351 , \26352 , \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 ,
         \26361 , \26362 , \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 ,
         \26371 , \26372 , \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 ,
         \26381 , \26382 , \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 ,
         \26391 , \26392 , \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 ,
         \26401 , \26402 , \26403 , \26404 , \26405 , \26406 , \26407 , \26408 , \26409 , \26410 ,
         \26411 , \26412 , \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 ,
         \26421 , \26422 , \26423 , \26424 , \26425 , \26426 , \26427 , \26428 , \26429 , \26430 ,
         \26431 , \26432 , \26433 , \26434 , \26435 , \26436 , \26437 , \26438 , \26439 , \26440 ,
         \26441 , \26442 , \26443 , \26444 , \26445 , \26446 , \26447 , \26448 , \26449 , \26450 ,
         \26451 , \26452 , \26453 , \26454 , \26455 , \26456 , \26457 , \26458 , \26459 , \26460 ,
         \26461 , \26462 , \26463 , \26464 , \26465 , \26466 , \26467 , \26468 , \26469 , \26470 ,
         \26471 , \26472 , \26473 , \26474 , \26475 , \26476 , \26477 , \26478 , \26479 , \26480 ,
         \26481 , \26482 , \26483 , \26484 , \26485 , \26486 , \26487 , \26488 , \26489 , \26490 ,
         \26491 , \26492 , \26493 , \26494 , \26495 , \26496 , \26497 , \26498 , \26499 , \26500 ,
         \26501 , \26502 , \26503 , \26504 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 ,
         \26511 , \26512 , \26513 , \26514 , \26515 , \26516 , \26517 , \26518 , \26519 , \26520 ,
         \26521 , \26522 , \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 ,
         \26531 , \26532 , \26533 , \26534 , \26535 , \26536 , \26537 , \26538 , \26539 , \26540 ,
         \26541 , \26542 , \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 ,
         \26551 , \26552 , \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 ,
         \26561 , \26562 , \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 ,
         \26571 , \26572 , \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 ,
         \26581 , \26582 , \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 ,
         \26591 , \26592 , \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 ,
         \26601 , \26602 , \26603 , \26604 , \26605 , \26606 , \26607 , \26608 , \26609 , \26610 ,
         \26611 , \26612 , \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 ,
         \26621 , \26622 , \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 ,
         \26631 , \26632 , \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 ,
         \26641 , \26642 , \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 ,
         \26651 , \26652 , \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 ,
         \26661 , \26662 , \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 , \26670 ,
         \26671 , \26672 , \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 ,
         \26681 , \26682 , \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 ,
         \26691 , \26692 , \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 ,
         \26701 , \26702 , \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 ,
         \26711 , \26712 , \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 ,
         \26721 , \26722 , \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 ,
         \26731 , \26732 , \26733 , \26734 , \26735 , \26736 , \26737 , \26738 , \26739 , \26740 ,
         \26741 , \26742 , \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 ,
         \26751 , \26752 , \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 ,
         \26761 , \26762 , \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 ,
         \26771 , \26772 , \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 ,
         \26781 , \26782 , \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 ,
         \26791 , \26792 , \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 ,
         \26801 , \26802 , \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 ,
         \26811 , \26812 , \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 , \26820 ,
         \26821 , \26822 , \26823 , \26824 , \26825 , \26826 , \26827 , \26828 , \26829 , \26830 ,
         \26831 , \26832 , \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 ,
         \26841 , \26842 , \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 ,
         \26851 , \26852 , \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 ,
         \26861 , \26862 , \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 ,
         \26871 , \26872 , \26873 , \26874 , \26875 , \26876 , \26877 , \26878 , \26879 , \26880 ,
         \26881 , \26882 , \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 ,
         \26891 , \26892 , \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 ,
         \26901 , \26902 , \26903 , \26904 , \26905 , \26906 , \26907 , \26908 , \26909 , \26910 ,
         \26911 , \26912 , \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 ,
         \26921 , \26922 , \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 ,
         \26931 , \26932 , \26933 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 ,
         \26941 , \26942 , \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 ,
         \26951 , \26952 , \26953 , \26954 , \26955 , \26956 , \26957 , \26958 , \26959 , \26960 ,
         \26961 , \26962 , \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 ,
         \26971 , \26972 , \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 ,
         \26981 , \26982 , \26983 , \26984 , \26985 , \26986 , \26987 , \26988 , \26989 , \26990 ,
         \26991 , \26992 , \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 ,
         \27001 , \27002 , \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 ,
         \27011 , \27012 , \27013 , \27014 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 ,
         \27021 , \27022 , \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 ,
         \27031 , \27032 , \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 ,
         \27041 , \27042 , \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 ,
         \27051 , \27052 , \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 ,
         \27061 , \27062 , \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 ,
         \27071 , \27072 , \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 ,
         \27081 , \27082 , \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 ,
         \27091 , \27092 , \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 ,
         \27101 , \27102 , \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 ,
         \27111 , \27112 , \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 ,
         \27121 , \27122 , \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 ,
         \27131 , \27132 , \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 ,
         \27141 , \27142 , \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 ,
         \27151 , \27152 , \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 ,
         \27161 , \27162 , \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 ,
         \27171 , \27172 , \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 ,
         \27181 , \27182 , \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 ,
         \27191 , \27192 , \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 ,
         \27201 , \27202 , \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 ,
         \27211 , \27212 , \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 ,
         \27221 , \27222 , \27223 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 ,
         \27231 , \27232 , \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 ,
         \27241 , \27242 , \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 ,
         \27251 , \27252 , \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 ,
         \27261 , \27262 , \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 ,
         \27271 , \27272 , \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 ,
         \27281 , \27282 , \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 ,
         \27291 , \27292 , \27293 , \27294 , \27295 , \27296 , \27297 , \27298 , \27299 , \27300 ,
         \27301 , \27302 , \27303 , \27304 , \27305 , \27306 , \27307 , \27308 , \27309 , \27310 ,
         \27311 , \27312 , \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 ,
         \27321 , \27322 , \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 ,
         \27331 , \27332 , \27333 , \27334 , \27335 , \27336 , \27337 , \27338 , \27339 , \27340 ,
         \27341 , \27342 , \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 ,
         \27351 , \27352 , \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 ,
         \27361 , \27362 , \27363 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 ,
         \27371 , \27372 , \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 ,
         \27381 , \27382 , \27383 , \27384 , \27385 , \27386 , \27387 , \27388 , \27389 , \27390 ,
         \27391 , \27392 , \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 ,
         \27401 , \27402 , \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 ,
         \27411 , \27412 , \27413 , \27414 , \27415 , \27416 , \27417 , \27418 , \27419 , \27420 ,
         \27421 , \27422 , \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 ,
         \27431 , \27432 , \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 ,
         \27441 , \27442 , \27443 , \27444 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 ,
         \27451 , \27452 , \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 ,
         \27461 , \27462 , \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 , \27470 ,
         \27471 , \27472 , \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 ,
         \27481 , \27482 , \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 ,
         \27491 , \27492 , \27493 , \27494 , \27495 , \27496 , \27497 , \27498 , \27499 , \27500 ,
         \27501 , \27502 , \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 ,
         \27511 , \27512 , \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 ,
         \27521 , \27522 , \27523 , \27524 , \27525 , \27526 , \27527 , \27528 , \27529 , \27530 ,
         \27531 , \27532 , \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 ,
         \27541 , \27542 , \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 ,
         \27551 , \27552 , \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 ,
         \27561 , \27562 , \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 ,
         \27571 , \27572 , \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 ,
         \27581 , \27582 , \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 ,
         \27591 , \27592 , \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 ,
         \27601 , \27602 , \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 ,
         \27611 , \27612 , \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 ,
         \27621 , \27622 , \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 ,
         \27631 , \27632 , \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 ,
         \27641 , \27642 , \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 ,
         \27651 , \27652 , \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 ,
         \27661 , \27662 , \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 ,
         \27671 , \27672 , \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 ,
         \27681 , \27682 , \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 ,
         \27691 , \27692 , \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 ,
         \27701 , \27702 , \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 ,
         \27711 , \27712 , \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 ,
         \27721 , \27722 , \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 ,
         \27731 , \27732 , \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 ,
         \27741 , \27742 , \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 ,
         \27751 , \27752 , \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 ,
         \27761 , \27762 , \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 ,
         \27771 , \27772 , \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 ,
         \27781 , \27782 , \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 ,
         \27791 , \27792 , \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 ,
         \27801 , \27802 , \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 ,
         \27811 , \27812 , \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 ,
         \27821 , \27822 , \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 ,
         \27831 , \27832 , \27833 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 ,
         \27841 , \27842 , \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 ,
         \27851 , \27852 , \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 ,
         \27861 , \27862 , \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 ,
         \27871 , \27872 , \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 ,
         \27881 , \27882 , \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 ,
         \27891 , \27892 , \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 ,
         \27901 , \27902 , \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 ,
         \27911 , \27912 , \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 ,
         \27921 , \27922 , \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 ,
         \27931 , \27932 , \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 ,
         \27941 , \27942 , \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 ,
         \27951 , \27952 , \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 ,
         \27961 , \27962 , \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 , \27970 ,
         \27971 , \27972 , \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 ,
         \27981 , \27982 , \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 ,
         \27991 , \27992 , \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 ,
         \28001 , \28002 , \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 ,
         \28011 , \28012 , \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 ,
         \28021 , \28022 , \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 ,
         \28031 , \28032 , \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 ,
         \28041 , \28042 , \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 ,
         \28051 , \28052 , \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 ,
         \28061 , \28062 , \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 ,
         \28071 , \28072 , \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 ,
         \28081 , \28082 , \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 ,
         \28091 , \28092 , \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 ,
         \28101 , \28102 , \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 ,
         \28111 , \28112 , \28113 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 ,
         \28121 , \28122 , \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 ,
         \28131 , \28132 , \28133 , \28134 , \28135 , \28136 , \28137 , \28138 , \28139 , \28140 ,
         \28141 , \28142 , \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 ,
         \28151 , \28152 , \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 ,
         \28161 , \28162 , \28163 , \28164 , \28165 , \28166 , \28167 , \28168 , \28169 , \28170 ,
         \28171 , \28172 , \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 ,
         \28181 , \28182 , \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 ,
         \28191 , \28192 , \28193 , \28194 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 ,
         \28201 , \28202 , \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 ,
         \28211 , \28212 , \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 , \28220 ,
         \28221 , \28222 , \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 ,
         \28231 , \28232 , \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 ,
         \28241 , \28242 , \28243 , \28244 , \28245 , \28246 , \28247 , \28248 , \28249 , \28250 ,
         \28251 , \28252 , \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 ,
         \28261 , \28262 , \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 ,
         \28271 , \28272 , \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 ,
         \28281 , \28282 , \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 ,
         \28291 , \28292 , \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 ,
         \28301 , \28302 , \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 ,
         \28311 , \28312 , \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 ,
         \28321 , \28322 , \28323 , \28324 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 ,
         \28331 , \28332 , \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 ,
         \28341 , \28342 , \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 ,
         \28351 , \28352 , \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 ,
         \28361 , \28362 , \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 ,
         \28371 , \28372 , \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 ,
         \28381 , \28382 , \28383 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 ,
         \28391 , \28392 , \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 ,
         \28401 , \28402 , \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 ,
         \28411 , \28412 , \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 ,
         \28421 , \28422 , \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 ,
         \28431 , \28432 , \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 ,
         \28441 , \28442 , \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 ,
         \28451 , \28452 , \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 ,
         \28461 , \28462 , \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 ,
         \28471 , \28472 , \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 ,
         \28481 , \28482 , \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 ,
         \28491 , \28492 , \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 ,
         \28501 , \28502 , \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 ,
         \28511 , \28512 , \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 ,
         \28521 , \28522 , \28523 , \28524 , \28525 , \28526 , \28527 , \28528 , \28529 , \28530 ,
         \28531 , \28532 , \28533 , \28534 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 ,
         \28541 , \28542 , \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 ,
         \28551 , \28552 , \28553 , \28554 , \28555 , \28556 , \28557 , \28558 , \28559 , \28560 ,
         \28561 , \28562 , \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 ,
         \28571 , \28572 , \28573 , \28574 , \28575 , \28576 , \28577 , \28578 , \28579 , \28580 ,
         \28581 , \28582 , \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 ,
         \28591 , \28592 , \28593 , \28594 , \28595 , \28596 , \28597 , \28598 , \28599 , \28600 ,
         \28601 , \28602 , \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 ,
         \28611 , \28612 , \28613 , \28614 , \28615 , \28616 , \28617 , \28618 , \28619 , \28620 ,
         \28621 , \28622 , \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 ,
         \28631 , \28632 , \28633 , \28634 , \28635 , \28636 , \28637 , \28638 , \28639 , \28640 ,
         \28641 , \28642 , \28643 , \28644 , \28645 , \28646 , \28647 , \28648 , \28649 , \28650 ,
         \28651 , \28652 , \28653 , \28654 , \28655 , \28656 , \28657 , \28658 , \28659 , \28660 ,
         \28661 , \28662 , \28663 , \28664 , \28665 , \28666 , \28667 , \28668 , \28669 , \28670 ,
         \28671 , \28672 , \28673 , \28674 , \28675 , \28676 , \28677 , \28678 , \28679 , \28680 ,
         \28681 , \28682 , \28683 , \28684 , \28685 , \28686 , \28687 , \28688 , \28689 , \28690 ,
         \28691 , \28692 , \28693 , \28694 , \28695 , \28696 , \28697 , \28698 , \28699 , \28700 ,
         \28701 , \28702 , \28703 , \28704 , \28705 , \28706 , \28707 , \28708 , \28709 , \28710 ,
         \28711 , \28712 , \28713 , \28714 , \28715 , \28716 , \28717 , \28718 , \28719 , \28720 ,
         \28721 , \28722 , \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 ,
         \28731 , \28732 , \28733 , \28734 , \28735 , \28736 , \28737 , \28738 , \28739 , \28740 ,
         \28741 , \28742 , \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 ,
         \28751 , \28752 , \28753 , \28754 , \28755 , \28756 , \28757 , \28758 , \28759 , \28760 ,
         \28761 , \28762 , \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , \28770 ,
         \28771 , \28772 , \28773 , \28774 , \28775 , \28776 , \28777 , \28778 , \28779 , \28780 ,
         \28781 , \28782 , \28783 , \28784 , \28785 , \28786 , \28787 , \28788 , \28789 , \28790 ,
         \28791 , \28792 , \28793 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 ,
         \28801 , \28802 , \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 ,
         \28811 , \28812 , \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 ,
         \28821 , \28822 , \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 ,
         \28831 , \28832 , \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 ,
         \28841 , \28842 , \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 ,
         \28851 , \28852 , \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 ,
         \28861 , \28862 , \28863 , \28864 , \28865 , \28866 , \28867 , \28868 , \28869 , \28870 ,
         \28871 , \28872 , \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 ,
         \28881 , \28882 , \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 ,
         \28891 , \28892 , \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 ,
         \28901 , \28902 , \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 ,
         \28911 , \28912 , \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 ,
         \28921 , \28922 , \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 ,
         \28931 , \28932 , \28933 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 ,
         \28941 , \28942 , \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 ,
         \28951 , \28952 , \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 ,
         \28961 , \28962 , \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 ,
         \28971 , \28972 , \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 ,
         \28981 , \28982 , \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 ,
         \28991 , \28992 , \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 ,
         \29001 , \29002 , \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 ,
         \29011 , \29012 , \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 ,
         \29021 , \29022 , \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 ,
         \29031 , \29032 , \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 ,
         \29041 , \29042 , \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 ,
         \29051 , \29052 , \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 ,
         \29061 , \29062 , \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 ,
         \29071 , \29072 , \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 ,
         \29081 , \29082 , \29083 , \29084 , \29085 , \29086 , \29087 , \29088 , \29089 , \29090 ,
         \29091 , \29092 , \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 ,
         \29101 , \29102 , \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 ,
         \29111 , \29112 , \29113 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 ,
         \29121 , \29122 , \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 ,
         \29131 , \29132 , \29133 , \29134 , \29135 , \29136 , \29137 , \29138 , \29139 , \29140 ,
         \29141 , \29142 , \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 ,
         \29151 , \29152 , \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 ,
         \29161 , \29162 , \29163 , \29164 , \29165 , \29166 , \29167 , \29168 , \29169 , \29170 ,
         \29171 , \29172 , \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 ,
         \29181 , \29182 , \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 ,
         \29191 , \29192 , \29193 , \29194 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 ,
         \29201 , \29202 , \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 ,
         \29211 , \29212 , \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 , \29220 ,
         \29221 , \29222 , \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 ,
         \29231 , \29232 , \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 ,
         \29241 , \29242 , \29243 , \29244 , \29245 , \29246 , \29247 , \29248 , \29249 , \29250 ,
         \29251 , \29252 , \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 ,
         \29261 , \29262 , \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 ,
         \29271 , \29272 , \29273 , \29274 , \29275 , \29276 , \29277 , \29278 , \29279 , \29280 ,
         \29281 , \29282 , \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 ,
         \29291 , \29292 , \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 ,
         \29301 , \29302 , \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 ,
         \29311 , \29312 , \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 ,
         \29321 , \29322 , \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 ,
         \29331 , \29332 , \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 ,
         \29341 , \29342 , \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 ,
         \29351 , \29352 , \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 ,
         \29361 , \29362 , \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 ,
         \29371 , \29372 , \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 ,
         \29381 , \29382 , \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 ,
         \29391 , \29392 , \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 ,
         \29401 , \29402 , \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 ,
         \29411 , \29412 , \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 ,
         \29421 , \29422 , \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 ,
         \29431 , \29432 , \29433 , \29434 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 ,
         \29441 , \29442 , \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 ,
         \29451 , \29452 , \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 ,
         \29461 , \29462 , \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 ,
         \29471 , \29472 , \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 ,
         \29481 , \29482 , \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 ,
         \29491 , \29492 , \29493 , \29494 , \29495 , \29496 , \29497 , \29498 , \29499 , \29500 ,
         \29501 , \29502 , \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 ,
         \29511 , \29512 , \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 ,
         \29521 , \29522 , \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 ,
         \29531 , \29532 , \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 ,
         \29541 , \29542 , \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 ,
         \29551 , \29552 , \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 ,
         \29561 , \29562 , \29563 , \29564 , \29565 , \29566 , \29567 , \29568 , \29569 , \29570 ,
         \29571 , \29572 , \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 ,
         \29581 , \29582 , \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 ,
         \29591 , \29592 , \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 ,
         \29601 , \29602 , \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 ,
         \29611 , \29612 , \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 ,
         \29621 , \29622 , \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 ,
         \29631 , \29632 , \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 ,
         \29641 , \29642 , \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 ,
         \29651 , \29652 , \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 ,
         \29661 , \29662 , \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 ,
         \29671 , \29672 , \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 ,
         \29681 , \29682 , \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 ,
         \29691 , \29692 , \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 ,
         \29701 , \29702 , \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 ,
         \29711 , \29712 , \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 ,
         \29721 , \29722 , \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 ,
         \29731 , \29732 , \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 ,
         \29741 , \29742 , \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 ,
         \29751 , \29752 , \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 ,
         \29761 , \29762 , \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 ,
         \29771 , \29772 , \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 ,
         \29781 , \29782 , \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 ,
         \29791 , \29792 , \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 ,
         \29801 , \29802 , \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 ,
         \29811 , \29812 , \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 ,
         \29821 , \29822 , \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 ,
         \29831 , \29832 , \29833 , \29834 , \29835 , \29836 , \29837 , \29838 , \29839 , \29840 ,
         \29841 , \29842 , \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 ,
         \29851 , \29852 , \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 ,
         \29861 , \29862 , \29863 , \29864 , \29865 , \29866 , \29867 , \29868 , \29869 , \29870 ,
         \29871 , \29872 , \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 ,
         \29881 , \29882 , \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 ,
         \29891 , \29892 , \29893 , \29894 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 ,
         \29901 , \29902 , \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 ,
         \29911 , \29912 , \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 , \29920 ,
         \29921 , \29922 , \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 ,
         \29931 , \29932 , \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 ,
         \29941 , \29942 , \29943 , \29944 , \29945 , \29946 , \29947 , \29948 , \29949 , \29950 ,
         \29951 , \29952 , \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 ,
         \29961 , \29962 , \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 ,
         \29971 , \29972 , \29973 , \29974 , \29975 , \29976 , \29977 , \29978 , \29979 , \29980 ,
         \29981 , \29982 , \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 ,
         \29991 , \29992 , \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 ,
         \30001 , \30002 , \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 ,
         \30011 , \30012 , \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 ,
         \30021 , \30022 , \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 ,
         \30031 , \30032 , \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 ,
         \30041 , \30042 , \30043 , \30044 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 ,
         \30051 , \30052 , \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 ,
         \30061 , \30062 , \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 ,
         \30071 , \30072 , \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 ,
         \30081 , \30082 , \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 ,
         \30091 , \30092 , \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 ,
         \30101 , \30102 , \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 ,
         \30111 , \30112 , \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 ,
         \30121 , \30122 , \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 ,
         \30131 , \30132 , \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 ,
         \30141 , \30142 , \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 ,
         \30151 , \30152 , \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 ,
         \30161 , \30162 , \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 ,
         \30171 , \30172 , \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 ,
         \30181 , \30182 , \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 ,
         \30191 , \30192 , \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 ,
         \30201 , \30202 , \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 ,
         \30211 , \30212 , \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 ,
         \30221 , \30222 , \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 ,
         \30231 , \30232 , \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 ,
         \30241 , \30242 , \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 ,
         \30251 , \30252 , \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 ,
         \30261 , \30262 , \30263 , \30264 , \30265 , \30266 , \30267 , \30268 , \30269 , \30270 ,
         \30271 , \30272 , \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 ,
         \30281 , \30282 , \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 ,
         \30291 , \30292 , \30293 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 ,
         \30301 , \30302 , \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 ,
         \30311 , \30312 , \30313 , \30314 , \30315 , \30316 , \30317 , \30318 , \30319 , \30320 ,
         \30321 , \30322 , \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 ,
         \30331 , \30332 , \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 ,
         \30341 , \30342 , \30343 , \30344 , \30345 , \30346 , \30347 , \30348 , \30349 , \30350 ,
         \30351 , \30352 , \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 ,
         \30361 , \30362 , \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 ,
         \30371 , \30372 , \30373 , \30374 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 ,
         \30381 , \30382 , \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 ,
         \30391 , \30392 , \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 , \30400 ,
         \30401 , \30402 , \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 ,
         \30411 , \30412 , \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 ,
         \30421 , \30422 , \30423 , \30424 , \30425 , \30426 , \30427 , \30428 , \30429 , \30430 ,
         \30431 , \30432 , \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 ,
         \30441 , \30442 , \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 ,
         \30451 , \30452 , \30453 , \30454 , \30455 , \30456 , \30457 , \30458 , \30459 , \30460 ,
         \30461 , \30462 , \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 ,
         \30471 , \30472 , \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 ,
         \30481 , \30482 , \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 ,
         \30491 , \30492 , \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 ,
         \30501 , \30502 , \30503 , \30504 , \30505 , \30506 , \30507 , \30508 , \30509 , \30510 ,
         \30511 , \30512 , \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 ,
         \30521 , \30522 , \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 ,
         \30531 , \30532 , \30533 , \30534 , \30535 , \30536 , \30537 , \30538 , \30539 , \30540 ,
         \30541 , \30542 , \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 ,
         \30551 , \30552 , \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 ,
         \30561 , \30562 , \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 ,
         \30571 , \30572 , \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 ,
         \30581 , \30582 , \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 ,
         \30591 , \30592 , \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 ,
         \30601 , \30602 , \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 ,
         \30611 , \30612 , \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 ,
         \30621 , \30622 , \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 ,
         \30631 , \30632 , \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 ,
         \30641 , \30642 , \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 ,
         \30651 , \30652 , \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 ,
         \30661 , \30662 , \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 ,
         \30671 , \30672 , \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 ,
         \30681 , \30682 , \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 ,
         \30691 , \30692 , \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 ,
         \30701 , \30702 , \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 ,
         \30711 , \30712 , \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 ,
         \30721 , \30722 , \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 ,
         \30731 , \30732 , \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 ,
         \30741 , \30742 , \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 ,
         \30751 , \30752 , \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 ,
         \30761 , \30762 , \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 ,
         \30771 , \30772 , \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 ,
         \30781 , \30782 , \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 ,
         \30791 , \30792 , \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 ,
         \30801 , \30802 , \30803 , \30804 , \30805 , \30806 , \30807 , \30808 , \30809 , \30810 ,
         \30811 , \30812 , \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 ,
         \30821 , \30822 , \30823 , \30824 , \30825 , \30826 , \30827 , \30828 , \30829 , \30830 ,
         \30831 , \30832 , \30833 , \30834 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 ,
         \30841 , \30842 , \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 ,
         \30851 , \30852 , \30853 , \30854 , \30855 , \30856 , \30857 , \30858 , \30859 , \30860 ,
         \30861 , \30862 , \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 ,
         \30871 , \30872 , \30873 , \30874 , \30875 , \30876 , \30877 , \30878 , \30879 , \30880 ,
         \30881 , \30882 , \30883 , \30884 , \30885 , \30886 , \30887 , \30888 , \30889 , \30890 ,
         \30891 , \30892 , \30893 , \30894 , \30895 , \30896 , \30897 , \30898 , \30899 , \30900 ,
         \30901 , \30902 , \30903 , \30904 , \30905 , \30906 , \30907 , \30908 , \30909 , \30910 ,
         \30911 , \30912 , \30913 , \30914 , \30915 , \30916 , \30917 , \30918 , \30919 , \30920 ,
         \30921 , \30922 , \30923 , \30924 , \30925 , \30926 , \30927 , \30928 , \30929 , \30930 ,
         \30931 , \30932 , \30933 , \30934 , \30935 , \30936 , \30937 , \30938 , \30939 , \30940 ,
         \30941 , \30942 , \30943 , \30944 , \30945 , \30946 , \30947 , \30948 , \30949 , \30950 ,
         \30951 , \30952 , \30953 , \30954 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 ,
         \30961 , \30962 , \30963 , \30964 , \30965 , \30966 , \30967 , \30968 , \30969 , \30970 ,
         \30971 , \30972 , \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 ,
         \30981 , \30982 , \30983 , \30984 , \30985 , \30986 , \30987 , \30988 , \30989 , \30990 ,
         \30991 , \30992 , \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 ,
         \31001 , \31002 , \31003 , \31004 , \31005 , \31006 , \31007 , \31008 , \31009 , \31010 ,
         \31011 , \31012 , \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 ,
         \31021 , \31022 , \31023 , \31024 , \31025 , \31026 , \31027 , \31028 , \31029 , \31030 ,
         \31031 , \31032 , \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 ,
         \31041 , \31042 , \31043 , \31044 , \31045 , \31046 , \31047 , \31048 , \31049 , \31050 ,
         \31051 , \31052 , \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 ,
         \31061 , \31062 , \31063 , \31064 , \31065 , \31066 , \31067 , \31068 , \31069 , \31070 ,
         \31071 , \31072 , \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 ,
         \31081 , \31082 , \31083 , \31084 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 ,
         \31091 , \31092 , \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 ,
         \31101 , \31102 , \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 ,
         \31111 , \31112 , \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 ,
         \31121 , \31122 , \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 ,
         \31131 , \31132 , \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 ,
         \31141 , \31142 , \31143 , \31144 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 ,
         \31151 , \31152 , \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 ,
         \31161 , \31162 , \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 ,
         \31171 , \31172 , \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 ,
         \31181 , \31182 , \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 ,
         \31191 , \31192 , \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 ,
         \31201 , \31202 , \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 ,
         \31211 , \31212 , \31213 , \31214 , \31215 , \31216 , \31217 , \31218 , \31219 , \31220 ,
         \31221 , \31222 , \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 ,
         \31231 , \31232 , \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 ,
         \31241 , \31242 , \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 ,
         \31251 , \31252 , \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 ,
         \31261 , \31262 , \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 ,
         \31271 , \31272 , \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 ,
         \31281 , \31282 , \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 ,
         \31291 , \31292 , \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 ,
         \31301 , \31302 , \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 ,
         \31311 , \31312 , \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 ,
         \31321 , \31322 , \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 ,
         \31331 , \31332 , \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 ,
         \31341 , \31342 , \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 ,
         \31351 , \31352 , \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 ,
         \31361 , \31362 , \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 ,
         \31371 , \31372 , \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 ,
         \31381 , \31382 , \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 ,
         \31391 , \31392 , \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 ,
         \31401 , \31402 , \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 ,
         \31411 , \31412 , \31413 , \31414 , \31415 , \31416 , \31417 , \31418 , \31419 , \31420 ,
         \31421 , \31422 , \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 ,
         \31431 , \31432 , \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 ,
         \31441 , \31442 , \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 ,
         \31451 , \31452 , \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 ,
         \31461 , \31462 , \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 ,
         \31471 , \31472 , \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 ,
         \31481 , \31482 , \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 ,
         \31491 , \31492 , \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 ,
         \31501 , \31502 , \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 ,
         \31511 , \31512 , \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 ,
         \31521 , \31522 , \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 ,
         \31531 , \31532 , \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 ,
         \31541 , \31542 , \31543 , \31544 , \31545 , \31546 , \31547 , \31548 , \31549 , \31550 ,
         \31551 , \31552 , \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 ,
         \31561 , \31562 , \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 ,
         \31571 , \31572 , \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 ,
         \31581 , \31582 , \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 ,
         \31591 , \31592 , \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 ,
         \31601 , \31602 , \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 ,
         \31611 , \31612 , \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 ,
         \31621 , \31622 , \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 , \31630 ,
         \31631 , \31632 , \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 ,
         \31641 , \31642 , \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 ,
         \31651 , \31652 , \31653 , \31654 , \31655 , \31656 , \31657 , \31658 , \31659 , \31660 ,
         \31661 , \31662 , \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 ,
         \31671 , \31672 , \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 ,
         \31681 , \31682 , \31683 , \31684 , \31685 , \31686 , \31687 , \31688 , \31689 , \31690 ,
         \31691 , \31692 , \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 ,
         \31701 , \31702 , \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 ,
         \31711 , \31712 , \31713 , \31714 , \31715 , \31716 , \31717 , \31718 , \31719 , \31720 ,
         \31721 , \31722 , \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 ,
         \31731 , \31732 , \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 ,
         \31741 , \31742 , \31743 , \31744 , \31745 , \31746 , \31747 , \31748 , \31749 , \31750 ,
         \31751 , \31752 , \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 ,
         \31761 , \31762 , \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 ,
         \31771 , \31772 , \31773 , \31774 , \31775 , \31776 , \31777 , \31778 , \31779 , \31780 ,
         \31781 , \31782 , \31783 , \31784 , \31785 , \31786 , \31787 , \31788 , \31789 , \31790 ,
         \31791 , \31792 , \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 ,
         \31801 , \31802 , \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 ,
         \31811 , \31812 , \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 ,
         \31821 , \31822 , \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 ,
         \31831 , \31832 , \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 ,
         \31841 , \31842 , \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 ,
         \31851 , \31852 , \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 ,
         \31861 , \31862 , \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 ,
         \31871 , \31872 , \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 ,
         \31881 , \31882 , \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 ,
         \31891 , \31892 , \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 ,
         \31901 , \31902 , \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 ,
         \31911 , \31912 , \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 ,
         \31921 , \31922 , \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 ,
         \31931 , \31932 , \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 ,
         \31941 , \31942 , \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 ,
         \31951 , \31952 , \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 ,
         \31961 , \31962 , \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 ,
         \31971 , \31972 , \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 ,
         \31981 , \31982 , \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 ,
         \31991 , \31992 , \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 ,
         \32001 , \32002 , \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 ,
         \32011 , \32012 , \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 ,
         \32021 , \32022 , \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 ,
         \32031 , \32032 , \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 ,
         \32041 , \32042 , \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 ,
         \32051 , \32052 , \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 , \32060 ,
         \32061 , \32062 , \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 ,
         \32071 , \32072 , \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 ,
         \32081 , \32082 , \32083 , \32084 , \32085 , \32086 , \32087 , \32088 , \32089 , \32090 ,
         \32091 , \32092 , \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 ,
         \32101 , \32102 , \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 ,
         \32111 , \32112 , \32113 , \32114 , \32115 , \32116 , \32117 , \32118 , \32119 , \32120 ,
         \32121 , \32122 , \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 ,
         \32131 , \32132 , \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 ,
         \32141 , \32142 , \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 ,
         \32151 , \32152 , \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 ,
         \32161 , \32162 , \32163 , \32164 , \32165 , \32166 , \32167 , \32168 , \32169 , \32170 ,
         \32171 , \32172 , \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 ,
         \32181 , \32182 , \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 ,
         \32191 , \32192 , \32193 , \32194 , \32195 , \32196 , \32197 , \32198 , \32199 , \32200 ,
         \32201 , \32202 , \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 ,
         \32211 , \32212 , \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 ,
         \32221 , \32222 , \32223 , \32224 , \32225 , \32226 , \32227 , \32228 , \32229 , \32230 ,
         \32231 , \32232 , \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 ,
         \32241 , \32242 , \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 ,
         \32251 , \32252 , \32253 , \32254 , \32255 , \32256 , \32257 , \32258 , \32259 , \32260 ,
         \32261 , \32262 , \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 ,
         \32271 , \32272 , \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 ,
         \32281 , \32282 , \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32289 , \32290 ,
         \32291 , \32292 , \32293 , \32294 , \32295 , \32296 , \32297 , \32298 , \32299 , \32300 ,
         \32301 , \32302 , \32303 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 ,
         \32311 , \32312 , \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 , \32320 ,
         \32321 , \32322 , \32323 , \32324 , \32325 , \32326 , \32327 , \32328 , \32329 , \32330 ,
         \32331 , \32332 , \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 ,
         \32341 , \32342 , \32343 , \32344 , \32345 , \32346 , \32347 , \32348 , \32349 , \32350 ,
         \32351 , \32352 , \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 ,
         \32361 , \32362 , \32363 , \32364 , \32365 , \32366 , \32367 , \32368 , \32369 , \32370 ,
         \32371 , \32372 , \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 ,
         \32381 , \32382 , \32383 , \32384 , \32385 , \32386 , \32387 , \32388 , \32389 , \32390 ,
         \32391 , \32392 , \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 ,
         \32401 , \32402 , \32403 , \32404 , \32405 , \32406 , \32407 , \32408 , \32409 , \32410 ,
         \32411 , \32412 , \32413 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 ,
         \32421 , \32422 , \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 , \32430 ,
         \32431 , \32432 , \32433 , \32434 , \32435 , \32436 , \32437 , \32438 , \32439 , \32440 ,
         \32441 , \32442 , \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 ,
         \32451 , \32452 , \32453 , \32454 , \32455 , \32456 , \32457 , \32458 , \32459 , \32460 ,
         \32461 , \32462 , \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 ,
         \32471 , \32472 , \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 ,
         \32481 , \32482 , \32483 , \32484 , \32485 , \32486 , \32487 , \32488 , \32489 , \32490 ,
         \32491 , \32492 , \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 ,
         \32501 , \32502 , \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 ,
         \32511 , \32512 , \32513 , \32514 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 ,
         \32521 , \32522 , \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 ,
         \32531 , \32532 , \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 ,
         \32541 , \32542 , \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 ,
         \32551 , \32552 , \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 ,
         \32561 , \32562 , \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 ,
         \32571 , \32572 , \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 ,
         \32581 , \32582 , \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 ,
         \32591 , \32592 , \32593 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 ,
         \32601 , \32602 , \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 ,
         \32611 , \32612 , \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 ,
         \32621 , \32622 , \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 ,
         \32631 , \32632 , \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 ,
         \32641 , \32642 , \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 ,
         \32651 , \32652 , \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 ,
         \32661 , \32662 , \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 ,
         \32671 , \32672 , \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 ,
         \32681 , \32682 , \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 ,
         \32691 , \32692 , \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 ,
         \32701 , \32702 , \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 ,
         \32711 , \32712 , \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 ,
         \32721 , \32722 , \32723 , \32724 , \32725 , \32726 , \32727 , \32728 , \32729 , \32730 ,
         \32731 , \32732 , \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 ,
         \32741 , \32742 , \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 ,
         \32751 , \32752 , \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 ,
         \32761 , \32762 , \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 ,
         \32771 , \32772 , \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 ,
         \32781 , \32782 , \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 ,
         \32791 , \32792 , \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 ,
         \32801 , \32802 , \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 , \32810 ,
         \32811 , \32812 , \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 ,
         \32821 , \32822 , \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 ,
         \32831 , \32832 , \32833 , \32834 , \32835 , \32836 , \32837 , \32838 , \32839 , \32840 ,
         \32841 , \32842 , \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 ,
         \32851 , \32852 , \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 ,
         \32861 , \32862 , \32863 , \32864 , \32865 , \32866 , \32867 , \32868 , \32869 , \32870 ,
         \32871 , \32872 , \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 ,
         \32881 , \32882 , \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 ,
         \32891 , \32892 , \32893 , \32894 , \32895 , \32896 , \32897 , \32898 , \32899 , \32900 ,
         \32901 , \32902 , \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 ,
         \32911 , \32912 , \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 ,
         \32921 , \32922 , \32923 , \32924 , \32925 , \32926 , \32927 , \32928 , \32929 , \32930 ,
         \32931 , \32932 , \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 ,
         \32941 , \32942 , \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 ,
         \32951 , \32952 , \32953 , \32954 , \32955 , \32956 , \32957 , \32958 , \32959 , \32960 ,
         \32961 , \32962 , \32963 , \32964 , \32965 , \32966 , \32967 , \32968 , \32969 , \32970 ,
         \32971 , \32972 , \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 ,
         \32981 , \32982 , \32983 , \32984 , \32985 , \32986 , \32987 , \32988 , \32989 , \32990 ,
         \32991 , \32992 , \32993 , \32994 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 ,
         \33001 , \33002 , \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 ,
         \33011 , \33012 , \33013 , \33014 , \33015 , \33016 , \33017 , \33018 , \33019 , \33020 ,
         \33021 , \33022 , \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 ,
         \33031 , \33032 , \33033 , \33034 , \33035 , \33036 , \33037 , \33038 , \33039 , \33040 ,
         \33041 , \33042 , \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 ,
         \33051 , \33052 , \33053 , \33054 , \33055 , \33056 , \33057 , \33058 , \33059 , \33060 ,
         \33061 , \33062 , \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 ,
         \33071 , \33072 , \33073 , \33074 , \33075 , \33076 , \33077 , \33078 , \33079 , \33080 ,
         \33081 , \33082 , \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 ,
         \33091 , \33092 , \33093 , \33094 , \33095 , \33096 , \33097 , \33098 , \33099 , \33100 ,
         \33101 , \33102 , \33103 , \33104 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 ,
         \33111 , \33112 , \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 ,
         \33121 , \33122 , \33123 , \33124 , \33125 , \33126 , \33127 , \33128 , \33129 , \33130 ,
         \33131 , \33132 , \33133 , \33134 , \33135 , \33136 , \33137 , \33138 , \33139 , \33140 ,
         \33141 , \33142 , \33143 , \33144 , \33145 , \33146 , \33147 , \33148 , \33149 , \33150 ,
         \33151 , \33152 , \33153 , \33154 , \33155 , \33156 , \33157 , \33158 , \33159 , \33160 ,
         \33161 , \33162 , \33163 , \33164 , \33165 , \33166 , \33167 , \33168 , \33169 , \33170 ,
         \33171 , \33172 , \33173 , \33174 , \33175 , \33176 , \33177 , \33178 , \33179 , \33180 ,
         \33181 , \33182 , \33183 , \33184 , \33185 , \33186 , \33187 , \33188 , \33189 , \33190 ,
         \33191 , \33192 , \33193 , \33194 , \33195 , \33196 , \33197 , \33198 , \33199 , \33200 ,
         \33201 , \33202 , \33203 , \33204 , \33205 , \33206 , \33207 , \33208 , \33209 , \33210 ,
         \33211 , \33212 , \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 ,
         \33221 , \33222 , \33223 , \33224 , \33225 , \33226 , \33227 , \33228 , \33229 , \33230 ,
         \33231 , \33232 , \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 ,
         \33241 , \33242 , \33243 , \33244 , \33245 , \33246 , \33247 , \33248 , \33249 , \33250 ,
         \33251 , \33252 , \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 ,
         \33261 , \33262 , \33263 , \33264 , \33265 , \33266 , \33267 , \33268 , \33269 , \33270 ,
         \33271 , \33272 , \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 ,
         \33281 , \33282 , \33283 , \33284 , \33285 , \33286 , \33287 , \33288 , \33289 , \33290 ,
         \33291 , \33292 , \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 ,
         \33301 , \33302 , \33303 , \33304 , \33305 , \33306 , \33307 , \33308 , \33309 , \33310 ,
         \33311 , \33312 , \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 ,
         \33321 , \33322 , \33323 , \33324 , \33325 , \33326 , \33327 , \33328 , \33329 , \33330 ,
         \33331 , \33332 , \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 ,
         \33341 , \33342 , \33343 , \33344 , \33345 , \33346 , \33347 , \33348 , \33349 , \33350 ,
         \33351 , \33352 , \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 ,
         \33361 , \33362 , \33363 , \33364 , \33365 , \33366 , \33367 , \33368 , \33369 , \33370 ,
         \33371 , \33372 , \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 ,
         \33381 , \33382 , \33383 , \33384 , \33385 , \33386 , \33387 , \33388 , \33389 , \33390 ,
         \33391 , \33392 , \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 ,
         \33401 , \33402 , \33403 , \33404 , \33405 , \33406 , \33407 , \33408 , \33409 , \33410 ,
         \33411 , \33412 , \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 ,
         \33421 , \33422 , \33423 , \33424 , \33425 , \33426 , \33427 , \33428 , \33429 , \33430 ,
         \33431 , \33432 , \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 ,
         \33441 , \33442 , \33443 , \33444 , \33445 , \33446 , \33447 , \33448 , \33449 , \33450 ,
         \33451 , \33452 , \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 ,
         \33461 , \33462 , \33463 , \33464 , \33465 , \33466 , \33467 , \33468 , \33469 , \33470 ,
         \33471 , \33472 , \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 ,
         \33481 , \33482 , \33483 , \33484 , \33485 , \33486 , \33487 , \33488 , \33489 , \33490 ,
         \33491 , \33492 , \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 ,
         \33501 , \33502 , \33503 , \33504 , \33505 , \33506 , \33507 , \33508 , \33509 , \33510 ,
         \33511 , \33512 , \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 ,
         \33521 , \33522 , \33523 , \33524 , \33525 , \33526 , \33527 , \33528 , \33529 , \33530 ,
         \33531 , \33532 , \33533 , \33534 , \33535 , \33536 , \33537 , \33538 , \33539 , \33540 ,
         \33541 , \33542 , \33543 , \33544 , \33545 , \33546 , \33547 , \33548 , \33549 , \33550 ,
         \33551 , \33552 , \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 ,
         \33561 , \33562 , \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 ,
         \33571 , \33572 , \33573 , \33574 , \33575 , \33576 , \33577 , \33578 , \33579 , \33580 ,
         \33581 , \33582 , \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 ,
         \33591 , \33592 , \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 ,
         \33601 , \33602 , \33603 , \33604 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 ,
         \33611 , \33612 , \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 ,
         \33621 , \33622 , \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 , \33630 ,
         \33631 , \33632 , \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 ,
         \33641 , \33642 , \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 ,
         \33651 , \33652 , \33653 , \33654 , \33655 , \33656 , \33657 , \33658 , \33659 , \33660 ,
         \33661 , \33662 , \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 ,
         \33671 , \33672 , \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 ,
         \33681 , \33682 , \33683 , \33684 , \33685 , \33686 , \33687 , \33688 , \33689 , \33690 ,
         \33691 , \33692 , \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 ,
         \33701 , \33702 , \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 ,
         \33711 , \33712 , \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 ,
         \33721 , \33722 , \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 ,
         \33731 , \33732 , \33733 , \33734 , \33735 , \33736 , \33737 , \33738 , \33739 , \33740 ,
         \33741 , \33742 , \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 ,
         \33751 , \33752 , \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 ,
         \33761 , \33762 , \33763 , \33764 , \33765 , \33766 , \33767 , \33768 , \33769 , \33770 ,
         \33771 , \33772 , \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 ,
         \33781 , \33782 , \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 ,
         \33791 , \33792 , \33793 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 ,
         \33801 , \33802 , \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 ,
         \33811 , \33812 , \33813 , \33814 , \33815 , \33816 , \33817 , \33818 , \33819 , \33820 ,
         \33821 , \33822 , \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 ,
         \33831 , \33832 , \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 ,
         \33841 , \33842 , \33843 , \33844 , \33845 , \33846 , \33847 , \33848 , \33849 , \33850 ,
         \33851 , \33852 , \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 ,
         \33861 , \33862 , \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 ,
         \33871 , \33872 , \33873 , \33874 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 ,
         \33881 , \33882 , \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 ,
         \33891 , \33892 , \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 , \33900 ,
         \33901 , \33902 , \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 ,
         \33911 , \33912 , \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 ,
         \33921 , \33922 , \33923 , \33924 , \33925 , \33926 , \33927 , \33928 , \33929 , \33930 ,
         \33931 , \33932 , \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 ,
         \33941 , \33942 , \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 ,
         \33951 , \33952 , \33953 , \33954 , \33955 , \33956 , \33957 , \33958 , \33959 , \33960 ,
         \33961 , \33962 , \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 ,
         \33971 , \33972 , \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 ,
         \33981 , \33982 , \33983 , \33984 , \33985 , \33986 , \33987 , \33988 , \33989 , \33990 ,
         \33991 , \33992 , \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 ,
         \34001 , \34002 , \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 ,
         \34011 , \34012 , \34013 , \34014 , \34015 , \34016 , \34017 , \34018 , \34019 , \34020 ,
         \34021 , \34022 , \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 ,
         \34031 , \34032 , \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 ,
         \34041 , \34042 , \34043 , \34044 , \34045 , \34046 , \34047 , \34048 , \34049 , \34050 ,
         \34051 , \34052 , \34053 , \34054 , \34055 , \34056 , \34057 , \34058 , \34059 , \34060 ,
         \34061 , \34062 , \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 ,
         \34071 , \34072 , \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 ,
         \34081 , \34082 , \34083 , \34084 , \34085 , \34086 , \34087 , \34088 , \34089 , \34090 ,
         \34091 , \34092 , \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 ,
         \34101 , \34102 , \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 ,
         \34111 , \34112 , \34113 , \34114 , \34115 , \34116 , \34117 , \34118 , \34119 , \34120 ,
         \34121 , \34122 , \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 ,
         \34131 , \34132 , \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 ,
         \34141 , \34142 , \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 ,
         \34151 , \34152 , \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 ,
         \34161 , \34162 , \34163 , \34164 , \34165 , \34166 , \34167 , \34168 , \34169 , \34170 ,
         \34171 , \34172 , \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 ,
         \34181 , \34182 , \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 ,
         \34191 , \34192 , \34193 , \34194 , \34195 , \34196 , \34197 , \34198 , \34199 , \34200 ,
         \34201 , \34202 , \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 ,
         \34211 , \34212 , \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 ,
         \34221 , \34222 , \34223 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 ,
         \34231 , \34232 , \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 ,
         \34241 , \34242 , \34243 , \34244 , \34245 , \34246 , \34247 , \34248 , \34249 , \34250 ,
         \34251 , \34252 , \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 ,
         \34261 , \34262 , \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 ,
         \34271 , \34272 , \34273 , \34274 , \34275 , \34276 , \34277 , \34278 , \34279 , \34280 ,
         \34281 , \34282 , \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 ,
         \34291 , \34292 , \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 ,
         \34301 , \34302 , \34303 , \34304 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 ,
         \34311 , \34312 , \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 ,
         \34321 , \34322 , \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 , \34330 ,
         \34331 , \34332 , \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 ,
         \34341 , \34342 , \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 ,
         \34351 , \34352 , \34353 , \34354 , \34355 , \34356 , \34357 , \34358 , \34359 , \34360 ,
         \34361 , \34362 , \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 ,
         \34371 , \34372 , \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 ,
         \34381 , \34382 , \34383 , \34384 , \34385 , \34386 , \34387 , \34388 , \34389 , \34390 ,
         \34391 , \34392 , \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 ,
         \34401 , \34402 , \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 ,
         \34411 , \34412 , \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 ,
         \34421 , \34422 , \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 ,
         \34431 , \34432 , \34433 , \34434 , \34435 , \34436 , \34437 , \34438 , \34439 , \34440 ,
         \34441 , \34442 , \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 ,
         \34451 , \34452 , \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 ,
         \34461 , \34462 , \34463 , \34464 , \34465 , \34466 , \34467 , \34468 , \34469 , \34470 ,
         \34471 , \34472 , \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 ,
         \34481 , \34482 , \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 ,
         \34491 , \34492 , \34493 , \34494 , \34495 , \34496 , \34497 , \34498 , \34499 , \34500 ,
         \34501 , \34502 , \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 ,
         \34511 , \34512 , \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 ,
         \34521 , \34522 , \34523 , \34524 , \34525 , \34526 , \34527 , \34528 , \34529 , \34530 ,
         \34531 , \34532 , \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 ,
         \34541 , \34542 , \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 ,
         \34551 , \34552 , \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34559 , \34560 ,
         \34561 , \34562 , \34563 , \34564 , \34565 , \34566 , \34567 , \34568 , \34569 , \34570 ,
         \34571 , \34572 , \34573 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 ,
         \34581 , \34582 , \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 , \34590 ,
         \34591 , \34592 , \34593 , \34594 , \34595 , \34596 , \34597 , \34598 , \34599 , \34600 ,
         \34601 , \34602 , \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 ,
         \34611 , \34612 , \34613 , \34614 , \34615 , \34616 , \34617 , \34618 , \34619 , \34620 ,
         \34621 , \34622 , \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 ,
         \34631 , \34632 , \34633 , \34634 , \34635 , \34636 , \34637 , \34638 , \34639 , \34640 ,
         \34641 , \34642 , \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 ,
         \34651 , \34652 , \34653 , \34654 , \34655 , \34656 , \34657 , \34658 , \34659 , \34660 ,
         \34661 , \34662 , \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 ,
         \34671 , \34672 , \34673 , \34674 , \34675 , \34676 , \34677 , \34678 , \34679 , \34680 ,
         \34681 , \34682 , \34683 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 ,
         \34691 , \34692 , \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 , \34700 ,
         \34701 , \34702 , \34703 , \34704 , \34705 , \34706 , \34707 , \34708 , \34709 , \34710 ,
         \34711 , \34712 , \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 ,
         \34721 , \34722 , \34723 , \34724 , \34725 , \34726 , \34727 , \34728 , \34729 , \34730 ,
         \34731 , \34732 , \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 ,
         \34741 , \34742 , \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 ,
         \34751 , \34752 , \34753 , \34754 , \34755 , \34756 , \34757 , \34758 , \34759 , \34760 ,
         \34761 , \34762 , \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 ,
         \34771 , \34772 , \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 ,
         \34781 , \34782 , \34783 , \34784 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 ,
         \34791 , \34792 , \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 ,
         \34801 , \34802 , \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 , \34810 ,
         \34811 , \34812 , \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 ,
         \34821 , \34822 , \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 ,
         \34831 , \34832 , \34833 , \34834 , \34835 , \34836 , \34837 , \34838 , \34839 , \34840 ,
         \34841 , \34842 , \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 ,
         \34851 , \34852 , \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 ,
         \34861 , \34862 , \34863 , \34864 , \34865 , \34866 , \34867 , \34868 , \34869 , \34870 ,
         \34871 , \34872 , \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 ,
         \34881 , \34882 , \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 ,
         \34891 , \34892 , \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 ,
         \34901 , \34902 , \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 ,
         \34911 , \34912 , \34913 , \34914 , \34915 , \34916 , \34917 , \34918 , \34919 , \34920 ,
         \34921 , \34922 , \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 ,
         \34931 , \34932 , \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 ,
         \34941 , \34942 , \34943 , \34944 , \34945 , \34946 , \34947 , \34948 , \34949 , \34950 ,
         \34951 , \34952 , \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 ,
         \34961 , \34962 , \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 ,
         \34971 , \34972 , \34973 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 ,
         \34981 , \34982 , \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 ,
         \34991 , \34992 , \34993 , \34994 , \34995 , \34996 , \34997 , \34998 , \34999 , \35000 ,
         \35001 , \35002 , \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 ,
         \35011 , \35012 , \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 ,
         \35021 , \35022 , \35023 , \35024 , \35025 , \35026 , \35027 , \35028 , \35029 , \35030 ,
         \35031 , \35032 , \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 ,
         \35041 , \35042 , \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 ,
         \35051 , \35052 , \35053 , \35054 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 ,
         \35061 , \35062 , \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 ,
         \35071 , \35072 , \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 , \35080 ,
         \35081 , \35082 , \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 ,
         \35091 , \35092 , \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 ,
         \35101 , \35102 , \35103 , \35104 , \35105 , \35106 , \35107 , \35108 , \35109 , \35110 ,
         \35111 , \35112 , \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 ,
         \35121 , \35122 , \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 ,
         \35131 , \35132 , \35133 , \35134 , \35135 , \35136 , \35137 , \35138 , \35139 , \35140 ,
         \35141 , \35142 , \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 ,
         \35151 , \35152 , \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 ,
         \35161 , \35162 , \35163 , \35164 , \35165 , \35166 , \35167 , \35168 , \35169 , \35170 ,
         \35171 , \35172 , \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 ,
         \35181 , \35182 , \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 ,
         \35191 , \35192 , \35193 , \35194 , \35195 , \35196 , \35197 , \35198 , \35199 , \35200 ,
         \35201 , \35202 , \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 ,
         \35211 , \35212 , \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 ,
         \35221 , \35222 , \35223 , \35224 , \35225 , \35226 , \35227 , \35228 , \35229 , \35230 ,
         \35231 , \35232 , \35233 , \35234 , \35235 , \35236 , \35237 , \35238 , \35239 , \35240 ,
         \35241 , \35242 , \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 ,
         \35251 , \35252 , \35253 , \35254 , \35255 , \35256 , \35257 , \35258 , \35259 , \35260 ,
         \35261 , \35262 , \35263 , \35264 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 ,
         \35271 , \35272 , \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 ,
         \35281 , \35282 , \35283 , \35284 , \35285 , \35286 , \35287 , \35288 , \35289 , \35290 ,
         \35291 , \35292 , \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 ,
         \35301 , \35302 , \35303 , \35304 , \35305 , \35306 , \35307 , \35308 , \35309 , \35310 ,
         \35311 , \35312 , \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 ,
         \35321 , \35322 , \35323 , \35324 , \35325 , \35326 , \35327 , \35328 , \35329 , \35330 ,
         \35331 , \35332 , \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 ,
         \35341 , \35342 , \35343 , \35344 , \35345 , \35346 , \35347 , \35348 , \35349 , \35350 ,
         \35351 , \35352 , \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 ,
         \35361 , \35362 , \35363 , \35364 , \35365 , \35366 , \35367 , \35368 , \35369 , \35370 ,
         \35371 , \35372 , \35373 , \35374 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 ,
         \35381 , \35382 , \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 ,
         \35391 , \35392 , \35393 , \35394 , \35395 , \35396 , \35397 , \35398 , \35399 , \35400 ,
         \35401 , \35402 , \35403 , \35404 , \35405 , \35406 , \35407 , \35408 , \35409 , \35410 ,
         \35411 , \35412 , \35413 , \35414 , \35415 , \35416 , \35417 , \35418 , \35419 , \35420 ,
         \35421 , \35422 , \35423 , \35424 , \35425 , \35426 , \35427 , \35428 , \35429 , \35430 ,
         \35431 , \35432 , \35433 , \35434 , \35435 , \35436 , \35437 , \35438 , \35439 , \35440 ,
         \35441 , \35442 , \35443 , \35444 , \35445 , \35446 , \35447 , \35448 , \35449 , \35450 ,
         \35451 , \35452 , \35453 , \35454 , \35455 , \35456 , \35457 , \35458 , \35459 , \35460 ,
         \35461 , \35462 , \35463 , \35464 , \35465 , \35466 , \35467 , \35468 , \35469 , \35470 ,
         \35471 , \35472 , \35473 , \35474 , \35475 , \35476 , \35477 , \35478 , \35479 , \35480 ,
         \35481 , \35482 , \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 ,
         \35491 , \35492 , \35493 , \35494 , \35495 , \35496 , \35497 , \35498 , \35499 , \35500 ,
         \35501 , \35502 , \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 ,
         \35511 , \35512 , \35513 , \35514 , \35515 , \35516 , \35517 , \35518 , \35519 , \35520 ,
         \35521 , \35522 , \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 ,
         \35531 , \35532 , \35533 , \35534 , \35535 , \35536 , \35537 , \35538 , \35539 , \35540 ,
         \35541 , \35542 , \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 ,
         \35551 , \35552 , \35553 , \35554 , \35555 , \35556 , \35557 , \35558 , \35559 , \35560 ,
         \35561 , \35562 , \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 ,
         \35571 , \35572 , \35573 , \35574 , \35575 , \35576 , \35577 , \35578 , \35579 , \35580 ,
         \35581 , \35582 , \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 ,
         \35591 , \35592 , \35593 , \35594 , \35595 , \35596 , \35597 , \35598 , \35599 , \35600 ,
         \35601 , \35602 , \35603 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 ,
         \35611 , \35612 , \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , \35619 , \35620 ,
         \35621 , \35622 , \35623 , \35624 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 ,
         \35631 , \35632 , \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , \35640 ,
         \35641 , \35642 , \35643 , \35644 , \35645 , \35646 , \35647 , \35648 , \35649 , \35650 ,
         \35651 , \35652 , \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 ,
         \35661 , \35662 , \35663 , \35664 , \35665 , \35666 , \35667 , \35668 , \35669 , \35670 ,
         \35671 , \35672 , \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 ,
         \35681 , \35682 , \35683 , \35684 , \35685 , \35686 , \35687 , \35688 , \35689 , \35690 ,
         \35691 , \35692 , \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 ,
         \35701 , \35702 , \35703 , \35704 , \35705 , \35706 , \35707 , \35708 , \35709 , \35710 ,
         \35711 , \35712 , \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 ,
         \35721 , \35722 , \35723 , \35724 , \35725 , \35726 , \35727 , \35728 , \35729 , \35730 ,
         \35731 , \35732 , \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 ,
         \35741 , \35742 , \35743 , \35744 , \35745 , \35746 , \35747 , \35748 , \35749 , \35750 ,
         \35751 , \35752 , \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 ,
         \35761 , \35762 , \35763 , \35764 , \35765 , \35766 , \35767 , \35768 , \35769 , \35770 ,
         \35771 , \35772 , \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 ,
         \35781 , \35782 , \35783 , \35784 , \35785 , \35786 , \35787 , \35788 , \35789 , \35790 ,
         \35791 , \35792 , \35793 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 ,
         \35801 , \35802 , \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , \35809 , \35810 ,
         \35811 , \35812 , \35813 , \35814 , \35815 , \35816 , \35817 , \35818 , \35819 , \35820 ,
         \35821 , \35822 , \35823 , \35824 , \35825 , \35826 , \35827 , \35828 , \35829 , \35830 ,
         \35831 , \35832 , \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 ,
         \35841 , \35842 , \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 ,
         \35851 , \35852 , \35853 , \35854 , \35855 , \35856 , \35857 , \35858 , \35859 , \35860 ,
         \35861 , \35862 , \35863 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 ,
         \35871 , \35872 , \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 ,
         \35881 , \35882 , \35883 , \35884 , \35885 , \35886 , \35887 , \35888 , \35889 , \35890 ,
         \35891 , \35892 , \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 ,
         \35901 , \35902 , \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 ,
         \35911 , \35912 , \35913 , \35914 , \35915 , \35916 , \35917 , \35918 , \35919 , \35920 ,
         \35921 , \35922 , \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 ,
         \35931 , \35932 , \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 ,
         \35941 , \35942 , \35943 , \35944 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 ,
         \35951 , \35952 , \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 ,
         \35961 , \35962 , \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 , \35970 ,
         \35971 , \35972 , \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 ,
         \35981 , \35982 , \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 ,
         \35991 , \35992 , \35993 , \35994 , \35995 , \35996 , \35997 , \35998 , \35999 , \36000 ,
         \36001 , \36002 , \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 ,
         \36011 , \36012 , \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 ,
         \36021 , \36022 , \36023 , \36024 , \36025 , \36026 , \36027 , \36028 , \36029 , \36030 ,
         \36031 , \36032 , \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 ,
         \36041 , \36042 , \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 ,
         \36051 , \36052 , \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 ,
         \36061 , \36062 , \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 ,
         \36071 , \36072 , \36073 , \36074 , \36075 , \36076 , \36077 , \36078 , \36079 , \36080 ,
         \36081 , \36082 , \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 ,
         \36091 , \36092 , \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 ,
         \36101 , \36102 , \36103 , \36104 , \36105 , \36106 , \36107 , \36108 , \36109 , \36110 ,
         \36111 , \36112 , \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 ,
         \36121 , \36122 , \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 ,
         \36131 , \36132 , \36133 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 ,
         \36141 , \36142 , \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 ,
         \36151 , \36152 , \36153 , \36154 , \36155 , \36156 , \36157 , \36158 , \36159 , \36160 ,
         \36161 , \36162 , \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 ,
         \36171 , \36172 , \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 ,
         \36181 , \36182 , \36183 , \36184 , \36185 , \36186 , \36187 , \36188 , \36189 , \36190 ,
         \36191 , \36192 , \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 ,
         \36201 , \36202 , \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 ,
         \36211 , \36212 , \36213 , \36214 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 ,
         \36221 , \36222 , \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 ,
         \36231 , \36232 , \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 , \36240 ,
         \36241 , \36242 , \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 ,
         \36251 , \36252 , \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 ,
         \36261 , \36262 , \36263 , \36264 , \36265 , \36266 , \36267 , \36268 , \36269 , \36270 ,
         \36271 , \36272 , \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 ,
         \36281 , \36282 , \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 ,
         \36291 , \36292 , \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 ,
         \36301 , \36302 , \36303 , \36304 , \36305 , \36306 , \36307 , \36308 , \36309 , \36310 ,
         \36311 , \36312 , \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 ,
         \36321 , \36322 , \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 ,
         \36331 , \36332 , \36333 , \36334 , \36335 , \36336 , \36337 , \36338 , \36339 , \36340 ,
         \36341 , \36342 , \36343 , \36344 , \36345 , \36346 , \36347 , \36348 , \36349 , \36350 ,
         \36351 , \36352 , \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 ,
         \36361 , \36362 , \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 ,
         \36371 , \36372 , \36373 , \36374 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 ,
         \36381 , \36382 , \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 ,
         \36391 , \36392 , \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 , \36400 ,
         \36401 , \36402 , \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 ,
         \36411 , \36412 , \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 ,
         \36421 , \36422 , \36423 , \36424 , \36425 , \36426 , \36427 , \36428 , \36429 , \36430 ,
         \36431 , \36432 , \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 ,
         \36441 , \36442 , \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 ,
         \36451 , \36452 , \36453 , \36454 , \36455 , \36456 , \36457 , \36458 , \36459 , \36460 ,
         \36461 , \36462 , \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 ,
         \36471 , \36472 , \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 ,
         \36481 , \36482 , \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 ,
         \36491 , \36492 , \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 ,
         \36501 , \36502 , \36503 , \36504 , \36505 , \36506 , \36507 , \36508 , \36509 , \36510 ,
         \36511 , \36512 , \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 ,
         \36521 , \36522 , \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 ,
         \36531 , \36532 , \36533 , \36534 , \36535 , \36536 , \36537 , \36538 , \36539 , \36540 ,
         \36541 , \36542 , \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 ,
         \36551 , \36552 , \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 ,
         \36561 , \36562 , \36563 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 ,
         \36571 , \36572 , \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 ,
         \36581 , \36582 , \36583 , \36584 , \36585 , \36586 , \36587 , \36588 , \36589 , \36590 ,
         \36591 , \36592 , \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 ,
         \36601 , \36602 , \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 ,
         \36611 , \36612 , \36613 , \36614 , \36615 , \36616 , \36617 , \36618 , \36619 , \36620 ,
         \36621 , \36622 , \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 ,
         \36631 , \36632 , \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 ,
         \36641 , \36642 , \36643 , \36644 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 ,
         \36651 , \36652 , \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 ,
         \36661 , \36662 , \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 , \36670 ,
         \36671 , \36672 , \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 ,
         \36681 , \36682 , \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 ,
         \36691 , \36692 , \36693 , \36694 , \36695 , \36696 , \36697 , \36698 , \36699 , \36700 ,
         \36701 , \36702 , \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 ,
         \36711 , \36712 , \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 ,
         \36721 , \36722 , \36723 , \36724 , \36725 , \36726 , \36727 , \36728 , \36729 , \36730 ,
         \36731 , \36732 , \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 ,
         \36741 , \36742 , \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 ,
         \36751 , \36752 , \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 ,
         \36761 , \36762 , \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 ,
         \36771 , \36772 , \36773 , \36774 , \36775 , \36776 , \36777 , \36778 , \36779 , \36780 ,
         \36781 , \36782 , \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 ,
         \36791 , \36792 , \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 ,
         \36801 , \36802 , \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 ,
         \36811 , \36812 , \36813 , \36814 , \36815 , \36816 , \36817 , \36818 , \36819 , \36820 ,
         \36821 , \36822 , \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 ,
         \36831 , \36832 , \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 ,
         \36841 , \36842 , \36843 , \36844 , \36845 , \36846 , \36847 , \36848 , \36849 , \36850 ,
         \36851 , \36852 , \36853 , \36854 , \36855 , \36856 , \36857 , \36858 , \36859 , \36860 ,
         \36861 , \36862 , \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 ,
         \36871 , \36872 , \36873 , \36874 , \36875 , \36876 , \36877 , \36878 , \36879 , \36880 ,
         \36881 , \36882 , \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 ,
         \36891 , \36892 , \36893 , \36894 , \36895 , \36896 , \36897 , \36898 , \36899 , \36900 ,
         \36901 , \36902 , \36903 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 ,
         \36911 , \36912 , \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 , \36920 ,
         \36921 , \36922 , \36923 , \36924 , \36925 , \36926 , \36927 , \36928 , \36929 , \36930 ,
         \36931 , \36932 , \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 ,
         \36941 , \36942 , \36943 , \36944 , \36945 , \36946 , \36947 , \36948 , \36949 , \36950 ,
         \36951 , \36952 , \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 ,
         \36961 , \36962 , \36963 , \36964 , \36965 , \36966 , \36967 , \36968 , \36969 , \36970 ,
         \36971 , \36972 , \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 ,
         \36981 , \36982 , \36983 , \36984 , \36985 , \36986 , \36987 , \36988 , \36989 , \36990 ,
         \36991 , \36992 , \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 ,
         \37001 , \37002 , \37003 , \37004 , \37005 , \37006 , \37007 , \37008 , \37009 , \37010 ,
         \37011 , \37012 , \37013 , \37014 , \37015 , \37016 , \37017 , \37018 , \37019 , \37020 ,
         \37021 , \37022 , \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 ,
         \37031 , \37032 , \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 ,
         \37041 , \37042 , \37043 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 ,
         \37051 , \37052 , \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 ,
         \37061 , \37062 , \37063 , \37064 , \37065 , \37066 , \37067 , \37068 , \37069 , \37070 ,
         \37071 , \37072 , \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 ,
         \37081 , \37082 , \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 ,
         \37091 , \37092 , \37093 , \37094 , \37095 , \37096 , \37097 , \37098 , \37099 , \37100 ,
         \37101 , \37102 , \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 ,
         \37111 , \37112 , \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 ,
         \37121 , \37122 , \37123 , \37124 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 ,
         \37131 , \37132 , \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 ,
         \37141 , \37142 , \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 , \37150 ,
         \37151 , \37152 , \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 ,
         \37161 , \37162 , \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 ,
         \37171 , \37172 , \37173 , \37174 , \37175 , \37176 , \37177 , \37178 , \37179 , \37180 ,
         \37181 , \37182 , \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 ,
         \37191 , \37192 , \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 ,
         \37201 , \37202 , \37203 , \37204 , \37205 , \37206 , \37207 , \37208 , \37209 , \37210 ,
         \37211 , \37212 , \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 ,
         \37221 , \37222 , \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 ,
         \37231 , \37232 , \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 ,
         \37241 , \37242 , \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 ,
         \37251 , \37252 , \37253 , \37254 , \37255 , \37256 , \37257 , \37258 , \37259 , \37260 ,
         \37261 , \37262 , \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 ,
         \37271 , \37272 , \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 ,
         \37281 , \37282 , \37283 , \37284 , \37285 , \37286 , \37287 , \37288 , \37289 , \37290 ,
         \37291 , \37292 , \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 ,
         \37301 , \37302 , \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 ,
         \37311 , \37312 , \37313 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 ,
         \37321 , \37322 , \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 ,
         \37331 , \37332 , \37333 , \37334 , \37335 , \37336 , \37337 , \37338 , \37339 , \37340 ,
         \37341 , \37342 , \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 ,
         \37351 , \37352 , \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 ,
         \37361 , \37362 , \37363 , \37364 , \37365 , \37366 , \37367 , \37368 , \37369 , \37370 ,
         \37371 , \37372 , \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 ,
         \37381 , \37382 , \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 ,
         \37391 , \37392 , \37393 , \37394 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 ,
         \37401 , \37402 , \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 ,
         \37411 , \37412 , \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 , \37420 ,
         \37421 , \37422 , \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 ,
         \37431 , \37432 , \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 ,
         \37441 , \37442 , \37443 , \37444 , \37445 , \37446 , \37447 , \37448 , \37449 , \37450 ,
         \37451 , \37452 , \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 ,
         \37461 , \37462 , \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 ,
         \37471 , \37472 , \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 ,
         \37481 , \37482 , \37483 , \37484 , \37485 , \37486 , \37487 , \37488 , \37489 , \37490 ,
         \37491 , \37492 , \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 ,
         \37501 , \37502 , \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 ,
         \37511 , \37512 , \37513 , \37514 , \37515 , \37516 , \37517 , \37518 , \37519 , \37520 ,
         \37521 , \37522 , \37523 , \37524 , \37525 , \37526 , \37527 , \37528 , \37529 , \37530 ,
         \37531 , \37532 , \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 ,
         \37541 , \37542 , \37543 , \37544 , \37545 , \37546 , \37547 , \37548 , \37549 , \37550 ,
         \37551 , \37552 , \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 ,
         \37561 , \37562 , \37563 , \37564 , \37565 , \37566 , \37567 , \37568 , \37569 , \37570 ,
         \37571 , \37572 , \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 ,
         \37581 , \37582 , \37583 , \37584 , \37585 , \37586 , \37587 , \37588 , \37589 , \37590 ,
         \37591 , \37592 , \37593 , \37594 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 ,
         \37601 , \37602 , \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 ,
         \37611 , \37612 , \37613 , \37614 , \37615 , \37616 , \37617 , \37618 , \37619 , \37620 ,
         \37621 , \37622 , \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 ,
         \37631 , \37632 , \37633 , \37634 , \37635 , \37636 , \37637 , \37638 , \37639 , \37640 ,
         \37641 , \37642 , \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 ,
         \37651 , \37652 , \37653 , \37654 , \37655 , \37656 , \37657 , \37658 , \37659 , \37660 ,
         \37661 , \37662 , \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 ,
         \37671 , \37672 , \37673 , \37674 , \37675 , \37676 , \37677 , \37678 , \37679 , \37680 ,
         \37681 , \37682 , \37683 , \37684 , \37685 , \37686 , \37687 , \37688 , \37689 , \37690 ,
         \37691 , \37692 , \37693 , \37694 , \37695 , \37696 , \37697 , \37698 , \37699 , \37700 ,
         \37701 , \37702 , \37703 , \37704 , \37705 , \37706 , \37707 , \37708 , \37709 , \37710 ,
         \37711 , \37712 , \37713 , \37714 , \37715 , \37716 , \37717 , \37718 , \37719 , \37720 ,
         \37721 , \37722 , \37723 , \37724 , \37725 , \37726 , \37727 , \37728 , \37729 , \37730 ,
         \37731 , \37732 , \37733 , \37734 , \37735 , \37736 , \37737 , \37738 , \37739 , \37740 ,
         \37741 , \37742 , \37743 , \37744 , \37745 , \37746 , \37747 , \37748 , \37749 , \37750 ,
         \37751 , \37752 , \37753 , \37754 , \37755 , \37756 , \37757 , \37758 , \37759 , \37760 ,
         \37761 , \37762 , \37763 , \37764 , \37765 , \37766 , \37767 , \37768 , \37769 , \37770 ,
         \37771 , \37772 , \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 ,
         \37781 , \37782 , \37783 , \37784 , \37785 , \37786 , \37787 , \37788 , \37789 , \37790 ,
         \37791 , \37792 , \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 ,
         \37801 , \37802 , \37803 , \37804 , \37805 , \37806 , \37807 , \37808 , \37809 , \37810 ,
         \37811 , \37812 , \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 ,
         \37821 , \37822 , \37823 , \37824 , \37825 , \37826 , \37827 , \37828 , \37829 , \37830 ,
         \37831 , \37832 , \37833 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 ,
         \37841 , \37842 , \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 , \37850 ,
         \37851 , \37852 , \37853 , \37854 , \37855 , \37856 , \37857 , \37858 , \37859 , \37860 ,
         \37861 , \37862 , \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 ,
         \37871 , \37872 , \37873 , \37874 , \37875 , \37876 , \37877 , \37878 , \37879 , \37880 ,
         \37881 , \37882 , \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 ,
         \37891 , \37892 , \37893 , \37894 , \37895 , \37896 , \37897 , \37898 , \37899 , \37900 ,
         \37901 , \37902 , \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 ,
         \37911 , \37912 , \37913 , \37914 , \37915 , \37916 , \37917 , \37918 , \37919 , \37920 ,
         \37921 , \37922 , \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 ,
         \37931 , \37932 , \37933 , \37934 , \37935 , \37936 , \37937 , \37938 , \37939 , \37940 ,
         \37941 , \37942 , \37943 , \37944 , \37945 , \37946 , \37947 , \37948 , \37949 , \37950 ,
         \37951 , \37952 , \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 ,
         \37961 , \37962 , \37963 , \37964 , \37965 , \37966 , \37967 , \37968 , \37969 , \37970 ,
         \37971 , \37972 , \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 ,
         \37981 , \37982 , \37983 , \37984 , \37985 , \37986 , \37987 , \37988 , \37989 , \37990 ,
         \37991 , \37992 , \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 ,
         \38001 , \38002 , \38003 , \38004 , \38005 , \38006 , \38007 , \38008 , \38009 , \38010 ,
         \38011 , \38012 , \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 ,
         \38021 , \38022 , \38023 , \38024 , \38025 , \38026 , \38027 , \38028 , \38029 , \38030 ,
         \38031 , \38032 , \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 ,
         \38041 , \38042 , \38043 , \38044 , \38045 , \38046 , \38047 , \38048 , \38049 , \38050 ,
         \38051 , \38052 , \38053 , \38054 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 ,
         \38061 , \38062 , \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 ,
         \38071 , \38072 , \38073 , \38074 , \38075 , \38076 , \38077 , \38078 , \38079 , \38080 ,
         \38081 , \38082 , \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 ,
         \38091 , \38092 , \38093 , \38094 , \38095 , \38096 , \38097 , \38098 , \38099 , \38100 ,
         \38101 , \38102 , \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 ,
         \38111 , \38112 , \38113 , \38114 , \38115 , \38116 , \38117 , \38118 , \38119 , \38120 ,
         \38121 , \38122 , \38123 , \38124 , \38125 , \38126 , \38127 , \38128 , \38129 , \38130 ,
         \38131 , \38132 , \38133 , \38134 , \38135 , \38136 , \38137 , \38138 , \38139 , \38140 ,
         \38141 , \38142 , \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 ,
         \38151 , \38152 , \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 ,
         \38161 , \38162 , \38163 , \38164 , \38165 , \38166 , \38167 , \38168 , \38169 , \38170 ,
         \38171 , \38172 , \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 ,
         \38181 , \38182 , \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 ,
         \38191 , \38192 , \38193 , \38194 , \38195 , \38196 , \38197 , \38198 , \38199 , \38200 ,
         \38201 , \38202 , \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 ,
         \38211 , \38212 , \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 ,
         \38221 , \38222 , \38223 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 ,
         \38231 , \38232 , \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 ,
         \38241 , \38242 , \38243 , \38244 , \38245 , \38246 , \38247 , \38248 , \38249 , \38250 ,
         \38251 , \38252 , \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 ,
         \38261 , \38262 , \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 ,
         \38271 , \38272 , \38273 , \38274 , \38275 , \38276 , \38277 , \38278 , \38279 , \38280 ,
         \38281 , \38282 , \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 ,
         \38291 , \38292 , \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 ,
         \38301 , \38302 , \38303 , \38304 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 ,
         \38311 , \38312 , \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 ,
         \38321 , \38322 , \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 , \38330 ,
         \38331 , \38332 , \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 ,
         \38341 , \38342 , \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 ,
         \38351 , \38352 , \38353 , \38354 , \38355 , \38356 , \38357 , \38358 , \38359 , \38360 ,
         \38361 , \38362 , \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 ,
         \38371 , \38372 , \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 ,
         \38381 , \38382 , \38383 , \38384 , \38385 , \38386 , \38387 , \38388 , \38389 , \38390 ,
         \38391 , \38392 , \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 ,
         \38401 , \38402 , \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 ,
         \38411 , \38412 , \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 ,
         \38421 , \38422 , \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 ,
         \38431 , \38432 , \38433 , \38434 , \38435 , \38436 , \38437 , \38438 , \38439 , \38440 ,
         \38441 , \38442 , \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 ,
         \38451 , \38452 , \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 ,
         \38461 , \38462 , \38463 , \38464 , \38465 , \38466 , \38467 , \38468 , \38469 , \38470 ,
         \38471 , \38472 , \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 ,
         \38481 , \38482 , \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 ,
         \38491 , \38492 , \38493 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 ,
         \38501 , \38502 , \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 ,
         \38511 , \38512 , \38513 , \38514 , \38515 , \38516 , \38517 , \38518 , \38519 , \38520 ,
         \38521 , \38522 , \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 ,
         \38531 , \38532 , \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 ,
         \38541 , \38542 , \38543 , \38544 , \38545 , \38546 , \38547 , \38548 , \38549 , \38550 ,
         \38551 , \38552 , \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 ,
         \38561 , \38562 , \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 ,
         \38571 , \38572 , \38573 , \38574 , \38575 , \38576 , \38577 , \38578 , \38579 , \38580 ,
         \38581 , \38582 , \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 ,
         \38591 , \38592 , \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 ,
         \38601 , \38602 , \38603 , \38604 , \38605 , \38606 , \38607 , \38608 , \38609 , \38610 ,
         \38611 , \38612 , \38613 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 ,
         \38621 , \38622 , \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 ,
         \38631 , \38632 , \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38640 ,
         \38641 , \38642 , \38643 , \38644 , \38645 , \38646 , \38647 , \38648 , \38649 , \38650 ,
         \38651 , \38652 , \38653 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 ,
         \38661 , \38662 , \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 ,
         \38671 , \38672 , \38673 , \38674 , \38675 , \38676 , \38677 , \38678 , \38679 , \38680 ,
         \38681 , \38682 , \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 ,
         \38691 , \38692 , \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 ,
         \38701 , \38702 , \38703 , \38704 , \38705 , \38706 , \38707 , \38708 , \38709 , \38710 ,
         \38711 , \38712 , \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 ,
         \38721 , \38722 , \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 ,
         \38731 , \38732 , \38733 , \38734 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 ,
         \38741 , \38742 , \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 ,
         \38751 , \38752 , \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 , \38760 ,
         \38761 , \38762 , \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 ,
         \38771 , \38772 , \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 ,
         \38781 , \38782 , \38783 , \38784 , \38785 , \38786 , \38787 , \38788 , \38789 , \38790 ,
         \38791 , \38792 , \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 ,
         \38801 , \38802 , \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 ,
         \38811 , \38812 , \38813 , \38814 , \38815 , \38816 , \38817 , \38818 , \38819 , \38820 ,
         \38821 , \38822 , \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 ,
         \38831 , \38832 , \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 ,
         \38841 , \38842 , \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 ,
         \38851 , \38852 , \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 ,
         \38861 , \38862 , \38863 , \38864 , \38865 , \38866 , \38867 , \38868 , \38869 , \38870 ,
         \38871 , \38872 , \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 ,
         \38881 , \38882 , \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 ,
         \38891 , \38892 , \38893 , \38894 , \38895 , \38896 , \38897 , \38898 , \38899 , \38900 ,
         \38901 , \38902 , \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 ,
         \38911 , \38912 , \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 ,
         \38921 , \38922 , \38923 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 ,
         \38931 , \38932 , \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 ,
         \38941 , \38942 , \38943 , \38944 , \38945 , \38946 , \38947 , \38948 , \38949 , \38950 ,
         \38951 , \38952 , \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 ,
         \38961 , \38962 , \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 ,
         \38971 , \38972 , \38973 , \38974 , \38975 , \38976 , \38977 , \38978 , \38979 , \38980 ,
         \38981 , \38982 , \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 ,
         \38991 , \38992 , \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 ,
         \39001 , \39002 , \39003 , \39004 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 ,
         \39011 , \39012 , \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 ,
         \39021 , \39022 , \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 , \39030 ,
         \39031 , \39032 , \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 ,
         \39041 , \39042 , \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 ,
         \39051 , \39052 , \39053 , \39054 , \39055 , \39056 , \39057 , \39058 , \39059 , \39060 ,
         \39061 , \39062 , \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 ,
         \39071 , \39072 , \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 ,
         \39081 , \39082 , \39083 , \39084 , \39085 , \39086 , \39087 , \39088 , \39089 , \39090 ,
         \39091 , \39092 , \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 ,
         \39101 , \39102 , \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 ,
         \39111 , \39112 , \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 , \39120 ,
         \39121 , \39122 , \39123 , \39124 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 ,
         \39131 , \39132 , \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 ,
         \39141 , \39142 , \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 ,
         \39151 , \39152 , \39153 , \39154 , \39155 , \39156 , \39157 , \39158 , \39159 , \39160 ,
         \39161 , \39162 , \39163 , \39164 , \39165 , \39166 , \39167 , \39168 , \39169 , \39170 ,
         \39171 , \39172 , \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 ,
         \39181 , \39182 , \39183 , \39184 , \39185 , \39186 , \39187 , \39188 , \39189 , \39190 ,
         \39191 , \39192 , \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 ,
         \39201 , \39202 , \39203 , \39204 , \39205 , \39206 , \39207 , \39208 , \39209 , \39210 ,
         \39211 , \39212 , \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 ,
         \39221 , \39222 , \39223 , \39224 , \39225 , \39226 , \39227 , \39228 , \39229 , \39230 ,
         \39231 , \39232 , \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 ,
         \39241 , \39242 , \39243 , \39244 , \39245 , \39246 , \39247 , \39248 , \39249 , \39250 ,
         \39251 , \39252 , \39253 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 ,
         \39261 , \39262 , \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 , \39270 ,
         \39271 , \39272 , \39273 , \39274 , \39275 , \39276 , \39277 , \39278 , \39279 , \39280 ,
         \39281 , \39282 , \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 ,
         \39291 , \39292 , \39293 , \39294 , \39295 , \39296 , \39297 , \39298 , \39299 , \39300 ,
         \39301 , \39302 , \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 ,
         \39311 , \39312 , \39313 , \39314 , \39315 , \39316 , \39317 , \39318 , \39319 , \39320 ,
         \39321 , \39322 , \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 ,
         \39331 , \39332 , \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 ,
         \39341 , \39342 , \39343 , \39344 , \39345 , \39346 , \39347 , \39348 , \39349 , \39350 ,
         \39351 , \39352 , \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 ,
         \39361 , \39362 , \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 ,
         \39371 , \39372 , \39373 , \39374 , \39375 , \39376 , \39377 , \39378 , \39379 , \39380 ,
         \39381 , \39382 , \39383 , \39384 , \39385 , \39386 , \39387 , \39388 , \39389 , \39390 ,
         \39391 , \39392 , \39393 , \39394 , \39395 , \39396 , \39397 , \39398 , \39399 , \39400 ,
         \39401 , \39402 , \39403 , \39404 , \39405 , \39406 , \39407 , \39408 , \39409 , \39410 ,
         \39411 , \39412 , \39413 , \39414 , \39415 , \39416 , \39417 , \39418 , \39419 , \39420 ,
         \39421 , \39422 , \39423 , \39424 , \39425 , \39426 , \39427 , \39428 , \39429 , \39430 ,
         \39431 , \39432 , \39433 , \39434 , \39435 , \39436 , \39437 , \39438 , \39439 , \39440 ,
         \39441 , \39442 , \39443 , \39444 , \39445 , \39446 , \39447 , \39448 , \39449 , \39450 ,
         \39451 , \39452 , \39453 , \39454 , \39455 , \39456 , \39457 , \39458 , \39459 , \39460 ,
         \39461 , \39462 , \39463 , \39464 , \39465 , \39466 , \39467 , \39468 , \39469 , \39470 ,
         \39471 , \39472 , \39473 , \39474 , \39475 , \39476 , \39477 , \39478 , \39479 , \39480 ,
         \39481 , \39482 , \39483 , \39484 , \39485 , \39486 , \39487 , \39488 , \39489 , \39490 ,
         \39491 , \39492 , \39493 , \39494 , \39495 , \39496 , \39497 , \39498 , \39499 , \39500 ,
         \39501 , \39502 , \39503 , \39504 , \39505 , \39506 , \39507 , \39508 , \39509 , \39510 ,
         \39511 , \39512 , \39513 , \39514 , \39515 , \39516 , \39517 , \39518 , \39519 , \39520 ,
         \39521 , \39522 , \39523 , \39524 , \39525 , \39526 , \39527 , \39528 , \39529 , \39530 ,
         \39531 , \39532 , \39533 , \39534 , \39535 , \39536 , \39537 , \39538 , \39539 , \39540 ,
         \39541 , \39542 , \39543 , \39544 , \39545 , \39546 , \39547 , \39548 , \39549 , \39550 ,
         \39551 , \39552 , \39553 , \39554 , \39555 , \39556 , \39557 , \39558 , \39559 , \39560 ,
         \39561 , \39562 , \39563 , \39564 , \39565 , \39566 , \39567 , \39568 , \39569 , \39570 ,
         \39571 , \39572 , \39573 , \39574 , \39575 , \39576 , \39577 , \39578 , \39579 , \39580 ,
         \39581 , \39582 , \39583 , \39584 , \39585 , \39586 , \39587 , \39588 , \39589 , \39590 ,
         \39591 , \39592 , \39593 , \39594 , \39595 , \39596 , \39597 , \39598 , \39599 , \39600 ,
         \39601 , \39602 , \39603 , \39604 , \39605 , \39606 , \39607 , \39608 , \39609 , \39610 ,
         \39611 , \39612 , \39613 , \39614 , \39615 , \39616 , \39617 , \39618 , \39619 , \39620 ,
         \39621 , \39622 , \39623 , \39624 , \39625 , \39626 , \39627 , \39628 , \39629 , \39630 ,
         \39631 , \39632 , \39633 , \39634 , \39635 , \39636 , \39637 , \39638 , \39639 , \39640 ,
         \39641 , \39642 , \39643 , \39644 , \39645 , \39646 , \39647 , \39648 , \39649 , \39650 ,
         \39651 , \39652 , \39653 , \39654 , \39655 , \39656 , \39657 , \39658 , \39659 , \39660 ,
         \39661 , \39662 , \39663 , \39664 , \39665 , \39666 , \39667 , \39668 , \39669 , \39670 ,
         \39671 , \39672 , \39673 , \39674 , \39675 , \39676 , \39677 , \39678 , \39679 , \39680 ,
         \39681 , \39682 , \39683 , \39684 , \39685 , \39686 , \39687 , \39688 , \39689 , \39690 ,
         \39691 , \39692 , \39693 , \39694 , \39695 , \39696 , \39697 , \39698 , \39699 , \39700 ,
         \39701 , \39702 , \39703 , \39704 , \39705 , \39706 , \39707 , \39708 , \39709 , \39710 ,
         \39711 , \39712 , \39713 , \39714 , \39715 , \39716 , \39717 , \39718 , \39719 , \39720 ,
         \39721 , \39722 , \39723 , \39724 , \39725 , \39726 , \39727 , \39728 , \39729 , \39730 ,
         \39731 , \39732 , \39733 , \39734 , \39735 , \39736 , \39737 , \39738 , \39739 , \39740 ,
         \39741 , \39742 , \39743 , \39744 , \39745 , \39746 , \39747 , \39748 , \39749 , \39750 ,
         \39751 , \39752 , \39753 , \39754 , \39755 , \39756 , \39757 , \39758 , \39759 , \39760 ,
         \39761 , \39762 , \39763 , \39764 , \39765 , \39766 , \39767 , \39768 , \39769 , \39770 ,
         \39771 , \39772 , \39773 , \39774 , \39775 , \39776 , \39777 , \39778 , \39779 , \39780 ,
         \39781 , \39782 , \39783 , \39784 , \39785 , \39786 , \39787 , \39788 , \39789 , \39790 ,
         \39791 , \39792 , \39793 , \39794 , \39795 , \39796 , \39797 , \39798 , \39799 , \39800 ,
         \39801 , \39802 , \39803 , \39804 , \39805 , \39806 , \39807 , \39808 , \39809 , \39810 ,
         \39811 , \39812 , \39813 , \39814 , \39815 , \39816 , \39817 , \39818 , \39819 , \39820 ,
         \39821 , \39822 , \39823 , \39824 , \39825 , \39826 , \39827 , \39828 , \39829 , \39830 ,
         \39831 , \39832 , \39833 , \39834 , \39835 , \39836 , \39837 , \39838 , \39839 , \39840 ,
         \39841 , \39842 , \39843 , \39844 , \39845 , \39846 , \39847 , \39848 , \39849 , \39850 ,
         \39851 , \39852 , \39853 , \39854 , \39855 , \39856 , \39857 , \39858 , \39859 , \39860 ,
         \39861 , \39862 , \39863 , \39864 , \39865 , \39866 , \39867 , \39868 , \39869 , \39870 ,
         \39871 , \39872 , \39873 , \39874 , \39875 , \39876 , \39877 , \39878 , \39879 , \39880 ,
         \39881 , \39882 , \39883 , \39884 , \39885 , \39886 , \39887 , \39888 , \39889 , \39890 ,
         \39891 , \39892 , \39893 , \39894 , \39895 , \39896 , \39897 , \39898 , \39899 , \39900 ,
         \39901 , \39902 , \39903 , \39904 , \39905 , \39906 , \39907 , \39908 , \39909 , \39910 ,
         \39911 , \39912 , \39913 , \39914 , \39915 , \39916 , \39917 , \39918 , \39919 , \39920 ,
         \39921 , \39922 , \39923 , \39924 , \39925 , \39926 , \39927 , \39928 , \39929 , \39930 ,
         \39931 , \39932 , \39933 , \39934 , \39935 , \39936 , \39937 , \39938 , \39939 , \39940 ,
         \39941 , \39942 , \39943 , \39944 , \39945 , \39946 , \39947 , \39948 , \39949 , \39950 ,
         \39951 , \39952 , \39953 , \39954 , \39955 , \39956 , \39957 , \39958 , \39959 , \39960 ,
         \39961 , \39962 , \39963 , \39964 , \39965 , \39966 , \39967 , \39968 , \39969 , \39970 ,
         \39971 , \39972 , \39973 , \39974 , \39975 , \39976 , \39977 , \39978 , \39979 , \39980 ,
         \39981 , \39982 , \39983 , \39984 , \39985 , \39986 , \39987 , \39988 , \39989 , \39990 ,
         \39991 , \39992 , \39993 , \39994 , \39995 , \39996 , \39997 , \39998 , \39999 , \40000 ,
         \40001 , \40002 , \40003 , \40004 , \40005 , \40006 , \40007 , \40008 , \40009 , \40010 ,
         \40011 , \40012 , \40013 , \40014 , \40015 , \40016 , \40017 , \40018 , \40019 , \40020 ,
         \40021 , \40022 , \40023 , \40024 , \40025 , \40026 , \40027 , \40028 , \40029 , \40030 ,
         \40031 , \40032 , \40033 , \40034 , \40035 , \40036 , \40037 , \40038 , \40039 , \40040 ,
         \40041 , \40042 , \40043 , \40044 , \40045 , \40046 , \40047 , \40048 , \40049 , \40050 ,
         \40051 , \40052 , \40053 , \40054 , \40055 , \40056 , \40057 , \40058 , \40059 , \40060 ,
         \40061 , \40062 , \40063 , \40064 , \40065 , \40066 , \40067 , \40068 , \40069 , \40070 ,
         \40071 , \40072 , \40073 , \40074 , \40075 , \40076 , \40077 , \40078 , \40079 , \40080 ,
         \40081 , \40082 , \40083 , \40084 , \40085 , \40086 , \40087 , \40088 , \40089 , \40090 ,
         \40091 , \40092 , \40093 , \40094 , \40095 , \40096 , \40097 , \40098 , \40099 , \40100 ,
         \40101 , \40102 , \40103 , \40104 , \40105 , \40106 , \40107 , \40108 , \40109 , \40110 ,
         \40111 , \40112 , \40113 , \40114 , \40115 , \40116 , \40117 , \40118 , \40119 , \40120 ,
         \40121 , \40122 , \40123 , \40124 , \40125 , \40126 , \40127 , \40128 , \40129 , \40130 ,
         \40131 , \40132 , \40133 , \40134 , \40135 , \40136 , \40137 , \40138 , \40139 , \40140 ,
         \40141 , \40142 , \40143 , \40144 , \40145 , \40146 , \40147 , \40148 , \40149 , \40150 ,
         \40151 , \40152 , \40153 , \40154 , \40155 , \40156 , \40157 , \40158 , \40159 , \40160 ,
         \40161 , \40162 , \40163 , \40164 , \40165 , \40166 , \40167 , \40168 , \40169 , \40170 ,
         \40171 , \40172 , \40173 , \40174 , \40175 , \40176 , \40177 , \40178 , \40179 , \40180 ,
         \40181 , \40182 , \40183 , \40184 , \40185 , \40186 , \40187 , \40188 , \40189 , \40190 ,
         \40191 , \40192 , \40193 , \40194 , \40195 , \40196 , \40197 , \40198 , \40199 , \40200 ,
         \40201 , \40202 , \40203 , \40204 , \40205 , \40206 , \40207 , \40208 , \40209 , \40210 ,
         \40211 , \40212 , \40213 , \40214 , \40215 , \40216 , \40217 , \40218 , \40219 , \40220 ,
         \40221 , \40222 , \40223 , \40224 , \40225 , \40226 , \40227 , \40228 , \40229 , \40230 ,
         \40231 , \40232 , \40233 , \40234 , \40235 , \40236 , \40237 , \40238 , \40239 , \40240 ,
         \40241 , \40242 , \40243 , \40244 , \40245 , \40246 , \40247 , \40248 , \40249 , \40250 ,
         \40251 , \40252 , \40253 , \40254 , \40255 , \40256 , \40257 , \40258 , \40259 , \40260 ,
         \40261 , \40262 , \40263 , \40264 , \40265 , \40266 , \40267 , \40268 , \40269 , \40270 ,
         \40271 , \40272 , \40273 , \40274 , \40275 , \40276 , \40277 , \40278 , \40279 , \40280 ,
         \40281 , \40282 , \40283 , \40284 , \40285 , \40286 , \40287 , \40288 , \40289 , \40290 ,
         \40291 , \40292 , \40293 , \40294 , \40295 , \40296 , \40297 , \40298 , \40299 , \40300 ,
         \40301 , \40302 , \40303 , \40304 , \40305 , \40306 , \40307 , \40308 , \40309 , \40310 ,
         \40311 , \40312 , \40313 , \40314 , \40315 , \40316 , \40317 , \40318 , \40319 , \40320 ,
         \40321 , \40322 , \40323 , \40324 , \40325 , \40326 , \40327 , \40328 , \40329 , \40330 ,
         \40331 , \40332 , \40333 , \40334 , \40335 , \40336 , \40337 , \40338 , \40339 , \40340 ,
         \40341 , \40342 , \40343 , \40344 , \40345 , \40346 , \40347 , \40348 , \40349 , \40350 ,
         \40351 , \40352 , \40353 , \40354 , \40355 , \40356 , \40357 , \40358 , \40359 , \40360 ,
         \40361 , \40362 , \40363 , \40364 , \40365 , \40366 , \40367 , \40368 , \40369 , \40370 ,
         \40371 , \40372 , \40373 , \40374 , \40375 , \40376 , \40377 , \40378 , \40379 , \40380 ,
         \40381 , \40382 , \40383 , \40384 , \40385 , \40386 , \40387 , \40388 , \40389 , \40390 ,
         \40391 , \40392 , \40393 , \40394 , \40395 , \40396 , \40397 , \40398 , \40399 , \40400 ,
         \40401 , \40402 , \40403 , \40404 , \40405 , \40406 , \40407 , \40408 , \40409 , \40410 ,
         \40411 , \40412 , \40413 , \40414 , \40415 , \40416 , \40417 , \40418 , \40419 , \40420 ,
         \40421 , \40422 , \40423 , \40424 , \40425 , \40426 , \40427 , \40428 , \40429 , \40430 ,
         \40431 , \40432 , \40433 , \40434 , \40435 , \40436 , \40437 , \40438 , \40439 , \40440 ,
         \40441 , \40442 , \40443 , \40444 , \40445 , \40446 , \40447 , \40448 , \40449 , \40450 ,
         \40451 , \40452 , \40453 , \40454 , \40455 , \40456 , \40457 , \40458 , \40459 , \40460 ,
         \40461 , \40462 , \40463 , \40464 , \40465 , \40466 , \40467 , \40468 , \40469 , \40470 ,
         \40471 , \40472 , \40473 , \40474 , \40475 , \40476 , \40477 , \40478 , \40479 , \40480 ,
         \40481 , \40482 , \40483 , \40484 , \40485 , \40486 , \40487 , \40488 , \40489 , \40490 ,
         \40491 , \40492 , \40493 , \40494 , \40495 , \40496 , \40497 , \40498 , \40499 , \40500 ,
         \40501 , \40502 , \40503 , \40504 , \40505 , \40506 , \40507 , \40508 , \40509 , \40510 ,
         \40511 , \40512 , \40513 , \40514 , \40515 , \40516 , \40517 , \40518 , \40519 , \40520 ,
         \40521 , \40522 , \40523 , \40524 , \40525 , \40526 , \40527 , \40528 , \40529 , \40530 ,
         \40531 , \40532 , \40533 , \40534 , \40535 , \40536 , \40537 , \40538 , \40539 , \40540 ,
         \40541 , \40542 , \40543 , \40544 , \40545 , \40546 , \40547 , \40548 , \40549 , \40550 ,
         \40551 , \40552 , \40553 , \40554 , \40555 , \40556 , \40557 , \40558 , \40559 , \40560 ,
         \40561 , \40562 , \40563 , \40564 , \40565 , \40566 , \40567 , \40568 , \40569 , \40570 ,
         \40571 , \40572 , \40573 , \40574 , \40575 , \40576 , \40577 , \40578 , \40579 , \40580 ,
         \40581 , \40582 , \40583 , \40584 , \40585 , \40586 , \40587 , \40588 , \40589 , \40590 ,
         \40591 , \40592 , \40593 , \40594 , \40595 , \40596 , \40597 , \40598 , \40599 , \40600 ,
         \40601 , \40602 , \40603 , \40604 , \40605 , \40606 , \40607 , \40608 , \40609 , \40610 ,
         \40611 , \40612 , \40613 , \40614 , \40615 , \40616 , \40617 , \40618 , \40619 , \40620 ,
         \40621 , \40622 , \40623 , \40624 , \40625 , \40626 , \40627 , \40628 , \40629 , \40630 ,
         \40631 , \40632 , \40633 , \40634 , \40635 , \40636 , \40637 , \40638 , \40639 , \40640 ,
         \40641 , \40642 , \40643 , \40644 , \40645 , \40646 , \40647 , \40648 , \40649 , \40650 ,
         \40651 , \40652 , \40653 , \40654 , \40655 , \40656 , \40657 , \40658 , \40659 , \40660 ,
         \40661 , \40662 , \40663 , \40664 , \40665 , \40666 , \40667 , \40668 , \40669 , \40670 ,
         \40671 , \40672 , \40673 , \40674 , \40675 , \40676 , \40677 , \40678 , \40679 , \40680 ,
         \40681 , \40682 , \40683 , \40684 , \40685 , \40686 , \40687 , \40688 , \40689 , \40690 ,
         \40691 , \40692 , \40693 , \40694 , \40695 , \40696 , \40697 , \40698 , \40699 , \40700 ,
         \40701 , \40702 , \40703 , \40704 , \40705 , \40706 , \40707 , \40708 , \40709 , \40710 ,
         \40711 , \40712 , \40713 , \40714 , \40715 , \40716 , \40717 , \40718 , \40719 , \40720 ,
         \40721 , \40722 , \40723 , \40724 , \40725 , \40726 , \40727 , \40728 , \40729 , \40730 ,
         \40731 , \40732 , \40733 , \40734 , \40735 , \40736 , \40737 , \40738 , \40739 , \40740 ,
         \40741 , \40742 , \40743 , \40744 , \40745 , \40746 , \40747 , \40748 , \40749 , \40750 ,
         \40751 , \40752 , \40753 , \40754 , \40755 , \40756 , \40757 , \40758 , \40759 , \40760 ,
         \40761 , \40762 , \40763 , \40764 , \40765 , \40766 , \40767 , \40768 , \40769 , \40770 ,
         \40771 , \40772 , \40773 , \40774 , \40775 , \40776 , \40777 , \40778 , \40779 , \40780 ,
         \40781 , \40782 , \40783 , \40784 , \40785 , \40786 , \40787 , \40788 , \40789 , \40790 ,
         \40791 , \40792 , \40793 , \40794 , \40795 , \40796 , \40797 , \40798 , \40799 , \40800 ,
         \40801 , \40802 , \40803 , \40804 , \40805 , \40806 , \40807 , \40808 , \40809 , \40810 ,
         \40811 , \40812 , \40813 , \40814 , \40815 , \40816 , \40817 , \40818 , \40819 , \40820 ,
         \40821 , \40822 , \40823 , \40824 , \40825 , \40826 , \40827 , \40828 , \40829 , \40830 ,
         \40831 , \40832 , \40833 , \40834 , \40835 , \40836 , \40837 , \40838 , \40839 , \40840 ,
         \40841 , \40842 , \40843 , \40844 , \40845 , \40846 , \40847 , \40848 , \40849 , \40850 ,
         \40851 , \40852 , \40853 , \40854 , \40855 , \40856 , \40857 , \40858 , \40859 , \40860 ,
         \40861 , \40862 , \40863 , \40864 , \40865 , \40866 , \40867 , \40868 , \40869 , \40870 ,
         \40871 , \40872 , \40873 , \40874 , \40875 , \40876 , \40877 , \40878 , \40879 , \40880 ,
         \40881 , \40882 , \40883 , \40884 , \40885 , \40886 , \40887 , \40888 , \40889 , \40890 ,
         \40891 , \40892 , \40893 , \40894 , \40895 , \40896 , \40897 , \40898 , \40899 , \40900 ,
         \40901 , \40902 , \40903 , \40904 , \40905 , \40906 , \40907 , \40908 , \40909 , \40910 ,
         \40911 , \40912 , \40913 , \40914 , \40915 , \40916 , \40917 , \40918 , \40919 , \40920 ,
         \40921 , \40922 , \40923 , \40924 , \40925 , \40926 , \40927 , \40928 , \40929 , \40930 ,
         \40931 , \40932 , \40933 , \40934 , \40935 , \40936 , \40937 , \40938 , \40939 , \40940 ,
         \40941 , \40942 , \40943 , \40944 , \40945 , \40946 , \40947 , \40948 , \40949 , \40950 ,
         \40951 , \40952 , \40953 , \40954 , \40955 , \40956 , \40957 , \40958 , \40959 , \40960 ,
         \40961 , \40962 , \40963 , \40964 , \40965 , \40966 , \40967 , \40968 , \40969 , \40970 ,
         \40971 , \40972 , \40973 , \40974 , \40975 , \40976 , \40977 , \40978 , \40979 , \40980 ,
         \40981 , \40982 , \40983 , \40984 , \40985 , \40986 , \40987 , \40988 , \40989 , \40990 ,
         \40991 , \40992 , \40993 , \40994 , \40995 , \40996 , \40997 , \40998 , \40999 , \41000 ,
         \41001 , \41002 , \41003 , \41004 , \41005 , \41006 , \41007 , \41008 , \41009 , \41010 ,
         \41011 , \41012 , \41013 , \41014 , \41015 , \41016 , \41017 , \41018 , \41019 , \41020 ,
         \41021 , \41022 , \41023 , \41024 , \41025 , \41026 , \41027 , \41028 , \41029 , \41030 ,
         \41031 , \41032 , \41033 , \41034 , \41035 , \41036 , \41037 , \41038 , \41039 , \41040 ,
         \41041 , \41042 , \41043 , \41044 , \41045 , \41046 , \41047 , \41048 , \41049 , \41050 ,
         \41051 , \41052 , \41053 , \41054 , \41055 , \41056 , \41057 , \41058 , \41059 , \41060 ,
         \41061 , \41062 , \41063 , \41064 , \41065 , \41066 , \41067 , \41068 , \41069 , \41070 ,
         \41071 , \41072 , \41073 , \41074 , \41075 , \41076 , \41077 , \41078 , \41079 , \41080 ,
         \41081 , \41082 , \41083 , \41084 , \41085 , \41086 , \41087 , \41088 , \41089 , \41090 ,
         \41091 , \41092 , \41093 , \41094 , \41095 , \41096 , \41097 , \41098 , \41099 , \41100 ,
         \41101 , \41102 , \41103 , \41104 , \41105 , \41106 , \41107 , \41108 , \41109 , \41110 ,
         \41111 , \41112 , \41113 , \41114 , \41115 , \41116 , \41117 , \41118 , \41119 , \41120 ,
         \41121 , \41122 , \41123 , \41124 , \41125 , \41126 , \41127 , \41128 , \41129 , \41130 ,
         \41131 , \41132 , \41133 , \41134 , \41135 , \41136 , \41137 , \41138 , \41139 , \41140 ,
         \41141 , \41142 , \41143 , \41144 , \41145 , \41146 , \41147 , \41148 , \41149 , \41150 ,
         \41151 , \41152 , \41153 , \41154 , \41155 , \41156 , \41157 , \41158 , \41159 , \41160 ,
         \41161 , \41162 , \41163 , \41164 , \41165 , \41166 , \41167 , \41168 , \41169 , \41170 ,
         \41171 , \41172 , \41173 , \41174 , \41175 , \41176 , \41177 , \41178 , \41179 , \41180 ,
         \41181 , \41182 , \41183 , \41184 , \41185 , \41186 , \41187 , \41188 , \41189 , \41190 ,
         \41191 , \41192 , \41193 , \41194 , \41195 , \41196 , \41197 , \41198 , \41199 , \41200 ,
         \41201 , \41202 , \41203 , \41204 , \41205 , \41206 , \41207 , \41208 , \41209 , \41210 ,
         \41211 , \41212 , \41213 , \41214 , \41215 , \41216 , \41217 , \41218 , \41219 , \41220 ,
         \41221 , \41222 , \41223 , \41224 , \41225 , \41226 , \41227 , \41228 , \41229 , \41230 ,
         \41231 , \41232 , \41233 , \41234 , \41235 , \41236 , \41237 , \41238 , \41239 , \41240 ,
         \41241 , \41242 , \41243 , \41244 , \41245 , \41246 , \41247 , \41248 , \41249 , \41250 ,
         \41251 , \41252 , \41253 , \41254 , \41255 , \41256 , \41257 , \41258 , \41259 , \41260 ,
         \41261 , \41262 , \41263 , \41264 , \41265 , \41266 , \41267 , \41268 , \41269 , \41270 ,
         \41271 , \41272 , \41273 , \41274 , \41275 , \41276 , \41277 , \41278 , \41279 , \41280 ,
         \41281 , \41282 , \41283 , \41284 , \41285 , \41286 , \41287 , \41288 , \41289 , \41290 ,
         \41291 , \41292 , \41293 , \41294 , \41295 , \41296 , \41297 , \41298 , \41299 , \41300 ,
         \41301 , \41302 , \41303 , \41304 , \41305 , \41306 , \41307 , \41308 , \41309 , \41310 ,
         \41311 , \41312 , \41313 , \41314 , \41315 , \41316 , \41317 , \41318 , \41319 , \41320 ,
         \41321 , \41322 , \41323 , \41324 , \41325 , \41326 , \41327 , \41328 , \41329 , \41330 ,
         \41331 , \41332 , \41333 , \41334 , \41335 , \41336 , \41337 , \41338 , \41339 , \41340 ,
         \41341 , \41342 , \41343 , \41344 , \41345 , \41346 , \41347 , \41348 , \41349 , \41350 ,
         \41351 , \41352 , \41353 , \41354 , \41355 , \41356 , \41357 , \41358 , \41359 , \41360 ,
         \41361 , \41362 , \41363 , \41364 , \41365 , \41366 , \41367 , \41368 , \41369 , \41370 ,
         \41371 , \41372 , \41373 , \41374 , \41375 , \41376 , \41377 , \41378 , \41379 , \41380 ,
         \41381 , \41382 , \41383 , \41384 , \41385 , \41386 , \41387 , \41388 , \41389 , \41390 ,
         \41391 , \41392 , \41393 , \41394 , \41395 , \41396 , \41397 , \41398 , \41399 , \41400 ,
         \41401 , \41402 , \41403 , \41404 , \41405 , \41406 , \41407 , \41408 , \41409 , \41410 ,
         \41411 , \41412 , \41413 , \41414 , \41415 , \41416 , \41417 , \41418 , \41419 , \41420 ,
         \41421 , \41422 , \41423 , \41424 , \41425 , \41426 , \41427 , \41428 , \41429 , \41430 ,
         \41431 , \41432 , \41433 , \41434 , \41435 , \41436 , \41437 , \41438 , \41439 , \41440 ,
         \41441 , \41442 , \41443 , \41444 , \41445 , \41446 , \41447 , \41448 , \41449 , \41450 ,
         \41451 , \41452 , \41453 , \41454 , \41455 , \41456 , \41457 , \41458 , \41459 , \41460 ,
         \41461 , \41462 , \41463 , \41464 , \41465 , \41466 , \41467 , \41468 , \41469 , \41470 ,
         \41471 , \41472 , \41473 , \41474 , \41475 , \41476 , \41477 , \41478 , \41479 , \41480 ,
         \41481 , \41482 , \41483 , \41484 , \41485 , \41486 , \41487 , \41488 , \41489 , \41490 ,
         \41491 , \41492 , \41493 , \41494 , \41495 , \41496 , \41497 , \41498 , \41499 , \41500 ,
         \41501 , \41502 , \41503 , \41504 , \41505 , \41506 , \41507 , \41508 , \41509 , \41510 ,
         \41511 , \41512 , \41513 , \41514 , \41515 , \41516 , \41517 , \41518 , \41519 , \41520 ,
         \41521 , \41522 , \41523 , \41524 , \41525 , \41526 , \41527 , \41528 , \41529 , \41530 ,
         \41531 , \41532 , \41533 , \41534 , \41535 , \41536 , \41537 , \41538 , \41539 , \41540 ,
         \41541 , \41542 , \41543 , \41544 , \41545 , \41546 , \41547 , \41548 , \41549 , \41550 ,
         \41551 , \41552 , \41553 , \41554 , \41555 , \41556 , \41557 , \41558 , \41559 , \41560 ,
         \41561 , \41562 , \41563 , \41564 , \41565 , \41566 , \41567 , \41568 , \41569 , \41570 ,
         \41571 , \41572 , \41573 , \41574 , \41575 , \41576 , \41577 , \41578 , \41579 , \41580 ,
         \41581 , \41582 , \41583 , \41584 , \41585 , \41586 , \41587 , \41588 , \41589 , \41590 ,
         \41591 , \41592 , \41593 , \41594 , \41595 , \41596 , \41597 , \41598 , \41599 , \41600 ,
         \41601 , \41602 , \41603 , \41604 , \41605 , \41606 , \41607 , \41608 , \41609 , \41610 ,
         \41611 , \41612 , \41613 , \41614 , \41615 , \41616 , \41617 , \41618 , \41619 , \41620 ,
         \41621 , \41622 , \41623 , \41624 , \41625 , \41626 , \41627 , \41628 , \41629 , \41630 ,
         \41631 , \41632 , \41633 , \41634 , \41635 , \41636 , \41637 , \41638 , \41639 , \41640 ,
         \41641 , \41642 , \41643 , \41644 , \41645 , \41646 , \41647 , \41648 , \41649 , \41650 ,
         \41651 , \41652 , \41653 , \41654 , \41655 , \41656 , \41657 , \41658 , \41659 , \41660 ,
         \41661 , \41662 , \41663 , \41664 , \41665 , \41666 , \41667 , \41668 , \41669 , \41670 ,
         \41671 , \41672 , \41673 , \41674 , \41675 , \41676 , \41677 , \41678 , \41679 , \41680 ,
         \41681 , \41682 , \41683 , \41684 , \41685 , \41686 , \41687 , \41688 , \41689 , \41690 ,
         \41691 , \41692 , \41693 , \41694 , \41695 , \41696 , \41697 , \41698 , \41699 , \41700 ,
         \41701 , \41702 , \41703 , \41704 , \41705 , \41706 , \41707 , \41708 , \41709 , \41710 ,
         \41711 , \41712 , \41713 , \41714 , \41715 , \41716 , \41717 , \41718 , \41719 , \41720 ,
         \41721 , \41722 , \41723 , \41724 , \41725 , \41726 , \41727 , \41728 , \41729 , \41730 ,
         \41731 , \41732 , \41733 , \41734 , \41735 , \41736 , \41737 , \41738 , \41739 , \41740 ,
         \41741 , \41742 , \41743 , \41744 , \41745 , \41746 , \41747 , \41748 , \41749 , \41750 ,
         \41751 , \41752 , \41753 , \41754 , \41755 , \41756 , \41757 , \41758 , \41759 , \41760 ,
         \41761 , \41762 , \41763 , \41764 , \41765 , \41766 , \41767 , \41768 , \41769 , \41770 ,
         \41771 , \41772 , \41773 , \41774 , \41775 , \41776 , \41777 , \41778 , \41779 , \41780 ,
         \41781 , \41782 , \41783 , \41784 , \41785 , \41786 , \41787 , \41788 , \41789 , \41790 ,
         \41791 , \41792 , \41793 , \41794 , \41795 , \41796 , \41797 , \41798 , \41799 , \41800 ,
         \41801 , \41802 , \41803 , \41804 , \41805 , \41806 , \41807 , \41808 , \41809 , \41810 ,
         \41811 , \41812 , \41813 , \41814 , \41815 , \41816 , \41817 , \41818 , \41819 , \41820 ,
         \41821 , \41822 , \41823 , \41824 , \41825 , \41826 , \41827 , \41828 , \41829 , \41830 ,
         \41831 , \41832 , \41833 , \41834 , \41835 , \41836 , \41837 , \41838 , \41839 , \41840 ,
         \41841 , \41842 , \41843 , \41844 , \41845 , \41846 , \41847 , \41848 , \41849 , \41850 ,
         \41851 , \41852 , \41853 , \41854 , \41855 , \41856 , \41857 , \41858 , \41859 , \41860 ,
         \41861 , \41862 , \41863 , \41864 , \41865 , \41866 , \41867 , \41868 , \41869 , \41870 ,
         \41871 , \41872 , \41873 , \41874 , \41875 , \41876 , \41877 , \41878 , \41879 , \41880 ,
         \41881 , \41882 , \41883 , \41884 , \41885 , \41886 , \41887 , \41888 , \41889 , \41890 ,
         \41891 , \41892 , \41893 , \41894 , \41895 , \41896 , \41897 , \41898 , \41899 , \41900 ,
         \41901 , \41902 , \41903 , \41904 , \41905 , \41906 , \41907 , \41908 , \41909 , \41910 ,
         \41911 , \41912 , \41913 , \41914 , \41915 , \41916 , \41917 , \41918 , \41919 , \41920 ,
         \41921 , \41922 , \41923 , \41924 , \41925 , \41926 , \41927 , \41928 , \41929 , \41930 ,
         \41931 , \41932 , \41933 , \41934 , \41935 , \41936 , \41937 , \41938 , \41939 , \41940 ,
         \41941 , \41942 , \41943 , \41944 , \41945 , \41946 , \41947 , \41948 , \41949 , \41950 ,
         \41951 , \41952 , \41953 , \41954 , \41955 , \41956 , \41957 , \41958 , \41959 , \41960 ,
         \41961 , \41962 , \41963 , \41964 , \41965 , \41966 , \41967 , \41968 , \41969 , \41970 ,
         \41971 , \41972 , \41973 , \41974 , \41975 , \41976 , \41977 , \41978 , \41979 , \41980 ,
         \41981 , \41982 , \41983 , \41984 , \41985 , \41986 , \41987 , \41988 , \41989 , \41990 ,
         \41991 , \41992 , \41993 , \41994 , \41995 , \41996 , \41997 , \41998 , \41999 , \42000 ,
         \42001 , \42002 , \42003 , \42004 , \42005 , \42006 , \42007 , \42008 , \42009 , \42010 ,
         \42011 , \42012 , \42013 , \42014 , \42015 , \42016 , \42017 , \42018 , \42019 , \42020 ,
         \42021 , \42022 , \42023 , \42024 , \42025 , \42026 , \42027 , \42028 , \42029 , \42030 ,
         \42031 , \42032 , \42033 , \42034 , \42035 , \42036 , \42037 , \42038 , \42039 , \42040 ,
         \42041 , \42042 , \42043 , \42044 , \42045 , \42046 , \42047 , \42048 , \42049 , \42050 ,
         \42051 , \42052 , \42053 , \42054 , \42055 , \42056 , \42057 , \42058 , \42059 , \42060 ,
         \42061 , \42062 , \42063 , \42064 , \42065 , \42066 , \42067 , \42068 , \42069 , \42070 ,
         \42071 , \42072 , \42073 , \42074 , \42075 , \42076 , \42077 , \42078 , \42079 , \42080 ,
         \42081 , \42082 , \42083 , \42084 , \42085 , \42086 , \42087 , \42088 , \42089 , \42090 ,
         \42091 , \42092 , \42093 , \42094 , \42095 , \42096 , \42097 , \42098 , \42099 , \42100 ,
         \42101 , \42102 , \42103 , \42104 , \42105 , \42106 , \42107 , \42108 , \42109 , \42110 ,
         \42111 , \42112 , \42113 , \42114 , \42115 , \42116 , \42117 , \42118 , \42119 , \42120 ,
         \42121 , \42122 , \42123 , \42124 , \42125 , \42126 , \42127 , \42128 , \42129 , \42130 ,
         \42131 , \42132 , \42133 , \42134 , \42135 , \42136 , \42137 , \42138 , \42139 , \42140 ,
         \42141 , \42142 , \42143 , \42144 , \42145 , \42146 , \42147 , \42148 , \42149 , \42150 ,
         \42151 , \42152 , \42153 , \42154 , \42155 , \42156 , \42157 , \42158 , \42159 , \42160 ,
         \42161 , \42162 , \42163 , \42164 , \42165 , \42166 , \42167 , \42168 , \42169 , \42170 ,
         \42171 , \42172 , \42173 , \42174 , \42175 , \42176 , \42177 , \42178 , \42179 , \42180 ,
         \42181 , \42182 , \42183 , \42184 , \42185 , \42186 , \42187 , \42188 , \42189 , \42190 ,
         \42191 , \42192 , \42193 , \42194 , \42195 , \42196 , \42197 , \42198 , \42199 , \42200 ,
         \42201 , \42202 , \42203 , \42204 , \42205 , \42206 , \42207 , \42208 , \42209 , \42210 ,
         \42211 , \42212 , \42213 , \42214 , \42215 , \42216 , \42217 , \42218 , \42219 , \42220 ,
         \42221 , \42222 , \42223 , \42224 , \42225 , \42226 , \42227 , \42228 , \42229 , \42230 ,
         \42231 , \42232 , \42233 , \42234 , \42235 , \42236 , \42237 , \42238 , \42239 , \42240 ,
         \42241 , \42242 , \42243 , \42244 , \42245 , \42246 , \42247 , \42248 , \42249 , \42250 ,
         \42251 , \42252 , \42253 , \42254 , \42255 , \42256 , \42257 , \42258 , \42259 , \42260 ,
         \42261 , \42262 , \42263 , \42264 , \42265 , \42266 , \42267 , \42268 , \42269 , \42270 ,
         \42271 , \42272 , \42273 , \42274 , \42275 , \42276 , \42277 , \42278 , \42279 , \42280 ,
         \42281 , \42282 , \42283 , \42284 , \42285 , \42286 , \42287 , \42288 , \42289 , \42290 ,
         \42291 , \42292 , \42293 , \42294 , \42295 , \42296 , \42297 , \42298 , \42299 , \42300 ,
         \42301 , \42302 , \42303 , \42304 , \42305 , \42306 , \42307 , \42308 , \42309 , \42310 ,
         \42311 , \42312 , \42313 , \42314 , \42315 , \42316 , \42317 , \42318 , \42319 , \42320 ,
         \42321 , \42322 , \42323 , \42324 , \42325 , \42326 , \42327 , \42328 , \42329 , \42330 ,
         \42331 , \42332 , \42333 , \42334 , \42335 , \42336 , \42337 , \42338 , \42339 , \42340 ,
         \42341 , \42342 , \42343 , \42344 , \42345 , \42346 , \42347 , \42348 , \42349 , \42350 ,
         \42351 , \42352 , \42353 , \42354 , \42355 , \42356 , \42357 , \42358 , \42359 , \42360 ,
         \42361 , \42362 , \42363 , \42364 , \42365 , \42366 , \42367 , \42368 , \42369 , \42370 ,
         \42371 , \42372 , \42373 , \42374 , \42375 , \42376 , \42377 , \42378 , \42379 , \42380 ,
         \42381 , \42382 , \42383 , \42384 , \42385 , \42386 , \42387 , \42388 , \42389 , \42390 ,
         \42391 , \42392 , \42393 , \42394 , \42395 , \42396 , \42397 , \42398 , \42399 , \42400 ,
         \42401 , \42402 , \42403 , \42404 , \42405 , \42406 , \42407 , \42408 , \42409 , \42410 ,
         \42411 , \42412 , \42413 , \42414 , \42415 , \42416 , \42417 , \42418 , \42419 , \42420 ,
         \42421 , \42422 , \42423 , \42424 , \42425 , \42426 , \42427 , \42428 , \42429 , \42430 ,
         \42431 , \42432 , \42433 , \42434 , \42435 , \42436 , \42437 , \42438 , \42439 , \42440 ,
         \42441 , \42442 , \42443 , \42444 , \42445 , \42446 , \42447 , \42448 , \42449 , \42450 ,
         \42451 , \42452 , \42453 , \42454 , \42455 , \42456 , \42457 , \42458 , \42459 , \42460 ,
         \42461 , \42462 , \42463 , \42464 , \42465 , \42466 , \42467 , \42468 , \42469 , \42470 ,
         \42471 , \42472 , \42473 , \42474 , \42475 , \42476 , \42477 , \42478 , \42479 , \42480 ,
         \42481 , \42482 , \42483 , \42484 , \42485 , \42486 , \42487 , \42488 , \42489 , \42490 ,
         \42491 , \42492 , \42493 , \42494 , \42495 , \42496 , \42497 , \42498 , \42499 , \42500 ,
         \42501 , \42502 , \42503 , \42504 , \42505 , \42506 , \42507 , \42508 , \42509 , \42510 ,
         \42511 , \42512 , \42513 , \42514 , \42515 , \42516 , \42517 , \42518 , \42519 , \42520 ,
         \42521 , \42522 , \42523 , \42524 , \42525 , \42526 , \42527 , \42528 , \42529 , \42530 ,
         \42531 , \42532 , \42533 , \42534 , \42535 , \42536 , \42537 , \42538 , \42539 , \42540 ;
buf \U$labaj4295 ( R_109_95e4d78, \41325 );
buf \U$labaj4296 ( R_10a_95e4e20, \41347 );
buf \U$labaj4297 ( R_10c_95e4f70, \41352 );
buf \U$labaj4298 ( R_10f_95e5168, \41362 );
buf \U$labaj4299 ( R_111_95e52b8, \41380 );
buf \U$labaj4300 ( R_119_95e57f8, \41399 );
buf \U$labaj4301 ( R_11c_95e59f0, \41409 );
buf \U$labaj4302 ( R_11d_95e5a98, \41419 );
buf \U$labaj4303 ( R_11f_95e5be8, \41430 );
buf \U$labaj4304 ( R_122_95e5de0, \41455 );
buf \U$labaj4305 ( R_123_95e5e88, \41463 );
buf \U$labaj4306 ( R_124_95e5f30, \41467 );
buf \U$labaj4307 ( R_125_95e5fd8, \41480 );
buf \U$labaj4308 ( R_127_95e6128, \41489 );
buf \U$labaj4309 ( R_128_95e61d0, \41497 );
buf \U$labaj4310 ( R_129_95e6278, \41517 );
buf \U$labaj4311 ( R_12b_95e63c8, \41526 );
buf \U$labaj4312 ( R_12c_95e6470, \41534 );
buf \U$labaj4313 ( R_12e_95e65c0, \41544 );
buf \U$labaj4314 ( R_12f_95e6668, \41554 );
buf \U$labaj4315 ( R_130_95e6710, \41558 );
buf \U$labaj4316 ( R_131_95e67b8, \41599 );
buf \U$labaj4317 ( R_135_95e6a58, \41611 );
buf \U$labaj4318 ( R_136_95e6b00, \41620 );
buf \U$labaj4319 ( R_137_95e6ba8, \41629 );
buf \U$labaj4320 ( R_138_95e6c50, \41636 );
buf \U$labaj4321 ( R_139_95e6cf8, \41657 );
buf \U$labaj4322 ( R_13b_95e6e48, \41668 );
buf \U$labaj4323 ( R_13d_95e6f98, \41684 );
buf \U$labaj4324 ( R_13e_95e7040, \41688 );
buf \U$labaj4325 ( R_13f_95e70e8, \41701 );
buf \U$labaj4326 ( R_140_95e7190, \41710 );
buf \U$labaj4327 ( R_141_95e7238, \41745 );
buf \U$labaj4328 ( R_143_95e7388, \41762 );
buf \U$labaj4329 ( R_144_95e7430, \41769 );
buf \U$labaj4330 ( R_145_95e74d8, \41794 );
buf \U$labaj4331 ( R_146_95e7580, \41806 );
buf \U$labaj4332 ( R_147_95e7628, \41823 );
buf \U$labaj4333 ( R_148_95e76d0, \41835 );
buf \U$labaj4334 ( R_149_95e7778, \41867 );
buf \U$labaj4335 ( R_14a_95e7820, \41880 );
buf \U$labaj4336 ( R_14b_95e78c8, \41897 );
buf \U$labaj4337 ( R_14c_95e7970, \41908 );
buf \U$labaj4338 ( R_14d_95e7a18, \41932 );
buf \U$labaj4339 ( R_14e_95e7ac0, \41944 );
buf \U$labaj4340 ( R_14f_95e7b68, \41957 );
buf \U$labaj4341 ( R_150_95e7c10, \41969 );
buf \U$labaj4342 ( R_151_95e7cb8, \42007 );
buf \U$labaj4343 ( R_152_95e7d60, \42019 );
buf \U$labaj4344 ( R_153_95e7e08, \42038 );
buf \U$labaj4345 ( R_154_95e7eb0, \42050 );
buf \U$labaj4346 ( R_155_95e7f58, \42074 );
buf \U$labaj4347 ( R_156_95e8000, \42086 );
buf \U$labaj4348 ( R_157_95e80a8, \42103 );
buf \U$labaj4349 ( R_158_95e8150, \42116 );
buf \U$labaj4350 ( R_159_95e81f8, \42142 );
buf \U$labaj4351 ( R_15a_95e82a0, \42150 );
buf \U$labaj4352 ( R_15b_95e8348, \42167 );
buf \U$labaj4353 ( R_15c_95e83f0, \42175 );
buf \U$labaj4354 ( R_15d_95e8498, \42195 );
buf \U$labaj4355 ( R_15e_95e8540, \42207 );
buf \U$labaj4356 ( R_15f_95e85e8, \42224 );
buf \U$labaj4357 ( R_160_95e8690, \42236 );
buf \U$labaj4358 ( R_161_95e8738, \42259 );
buf \U$labaj4359 ( R_162_95e87e0, \42271 );
buf \U$labaj4360 ( R_163_95e8888, \42288 );
buf \U$labaj4361 ( R_164_95e8930, \42300 );
buf \U$labaj4362 ( R_165_95e89d8, \42323 );
buf \U$labaj4363 ( R_166_95e8a80, \42335 );
buf \U$labaj4364 ( R_167_95e8b28, \42353 );
buf \U$labaj4365 ( R_168_95e8bd0, \42365 );
buf \U$labaj4366 ( R_169_95e8c78, \42389 );
buf \U$labaj4367 ( R_16a_95e8d20, \42400 );
buf \U$labaj4368 ( R_16b_95e8dc8, \42416 );
buf \U$labaj4369 ( R_16c_95e8e70, \42424 );
buf \U$labaj4370 ( R_16d_95e8f18, \42445 );
buf \U$labaj4371 ( R_16e_95e8fc0, \42457 );
buf \U$labaj4372 ( R_16f_95e9068, \42474 );
buf \U$labaj4373 ( R_170_95e9110, \42485 );
buf \U$labaj4374 ( R_171_95e91b8, \42492 );
buf \U$labaj4375 ( R_172_95e9260, \42499 );
buf \U$labaj4376 ( R_173_95e9308, \42511 );
buf \U$labaj4377 ( R_174_95e93b0, \42519 );
buf \U$labaj4378 ( R_175_95e9458, \42533 );
buf \U$labaj4379 ( R_176_95e9500, \42540 );
nor \U$1 ( \344 , RIbb2d630_69, RIbb317d0_133);
nor \U$2 ( \345 , RIbb2d5b8_70, RIbb31848_134);
nor \U$3 ( \346 , \344 , \345 );
nor \U$4 ( \347 , RIbb2d540_71, RIbb318c0_135);
nor \U$5 ( \348 , RIbb2d4c8_72, RIbb31938_136);
nor \U$6 ( \349 , \347 , \348 );
and \U$7 ( \350 , \346 , \349 );
or \U$8 ( \351 , RIbb2d720_67, RIbb316e0_131);
or \U$9 ( \352 , RIbb2d6a8_68, RIbb31758_132);
nand \U$10 ( \353 , \351 , \352 );
nor \U$11 ( \354 , RIbb2d798_66, RIbb31668_130);
not \U$12 ( \355 , \354 );
or \U$13 ( \356 , RIbb2d810_65, RIbb315f0_129);
nand \U$14 ( \357 , \355 , \356 );
nor \U$15 ( \358 , \353 , \357 );
nand \U$16 ( \359 , \350 , \358 );
not \U$17 ( \360 , \359 );
not \U$18 ( \361 , \360 );
not \U$19 ( \362 , RIbb2cfa0_83);
not \U$20 ( \363 , RIbb31e60_147);
and \U$21 ( \364 , \362 , \363 );
nor \U$22 ( \365 , RIbb2cf28_84, RIbb31ed8_148);
nor \U$23 ( \366 , \364 , \365 );
nor \U$24 ( \367 , RIbb2d090_81, RIbb31d70_145);
nor \U$25 ( \368 , RIbb2d018_82, RIbb31de8_146);
nor \U$26 ( \369 , \367 , \368 );
nand \U$27 ( \370 , \366 , \369 );
not \U$28 ( \371 , \370 );
nor \U$29 ( \372 , RIbb2caf0_93, RIbb32310_157);
nor \U$30 ( \373 , RIbb2ca78_94, RIbb32388_158);
nor \U$31 ( \374 , \372 , \373 );
nor \U$32 ( \375 , RIbb2ca00_95, RIbb32400_159);
nor \U$33 ( \376 , RIbb2c988_96, RIbb32478_160);
nor \U$34 ( \377 , \375 , \376 );
nand \U$35 ( \378 , \374 , \377 );
nor \U$36 ( \379 , RIbb2cc58_90, RIbb321a8_154);
nor \U$37 ( \380 , RIbb2ccd0_89, RIbb32130_153);
nor \U$38 ( \381 , \379 , \380 );
nor \U$39 ( \382 , RIbb2cbe0_91, RIbb32220_155);
nor \U$40 ( \383 , RIbb2cb68_92, RIbb32298_156);
nor \U$41 ( \384 , \382 , \383 );
nand \U$42 ( \385 , \381 , \384 );
nor \U$43 ( \386 , \378 , \385 );
nor \U$44 ( \387 , RIbb2cdc0_87, RIbb32040_151);
nor \U$45 ( \388 , RIbb2cd48_88, RIbb320b8_152);
nor \U$46 ( \389 , \387 , \388 );
or \U$47 ( \390 , RIbb2ceb0_85, RIbb31f50_149);
nor \U$48 ( \391 , RIbb2ce38_86, RIbb31fc8_150);
not \U$49 ( \392 , \391 );
nand \U$50 ( \393 , \389 , \390 , \392 );
not \U$51 ( \394 , \393 );
nand \U$52 ( \395 , \371 , \386 , \394 );
not \U$53 ( \396 , \395 );
not \U$54 ( \397 , \396 );
nor \U$55 ( \398 , RIbb2d360_75, RIbb31aa0_139);
nor \U$56 ( \399 , RIbb2d2e8_76, RIbb31b18_140);
nor \U$57 ( \400 , \398 , \399 );
nor \U$58 ( \401 , RIbb2d3d8_74, RIbb31a28_138);
nor \U$59 ( \402 , RIbb2d450_73, RIbb319b0_137);
nor \U$60 ( \403 , \401 , \402 );
and \U$61 ( \404 , \400 , \403 );
nor \U$62 ( \405 , RIbb2d180_79, RIbb31c80_143);
nor \U$63 ( \406 , RIbb2d108_80, RIbb31cf8_144);
nor \U$64 ( \407 , \405 , \406 );
or \U$65 ( \408 , RIbb2d270_77, RIbb31b90_141);
or \U$66 ( \409 , RIbb2d1f8_78, RIbb31c08_142);
and \U$67 ( \410 , \407 , \408 , \409 );
nand \U$68 ( \411 , \404 , \410 );
buf \U$69 ( \412 , \411 );
nor \U$70 ( \413 , \361 , \397 , \412 );
not \U$71 ( \414 , \413 );
and \U$72 ( \415 , RIbb2be48_120, RIbb32fb8_184);
not \U$73 ( \416 , \415 );
not \U$74 ( \417 , RIbb2bec0_119);
not \U$75 ( \418 , RIbb32f40_183);
nand \U$76 ( \419 , \417 , \418 );
not \U$77 ( \420 , \419 );
or \U$78 ( \421 , \416 , \420 );
nand \U$79 ( \422 , RIbb2bec0_119, RIbb32f40_183);
nand \U$80 ( \423 , \421 , \422 );
not \U$81 ( \424 , \423 );
not \U$82 ( \425 , RIbb2bfb0_117);
not \U$83 ( \426 , RIbb32e50_181);
nand \U$84 ( \427 , \425 , \426 );
not \U$85 ( \428 , \427 );
not \U$86 ( \429 , RIbb2bf38_118);
not \U$87 ( \430 , RIbb32ec8_182);
nand \U$88 ( \431 , \429 , \430 );
not \U$89 ( \432 , \431 );
nor \U$90 ( \433 , \428 , \432 );
not \U$91 ( \434 , \433 );
or \U$92 ( \435 , \424 , \434 );
not \U$93 ( \436 , \428 );
nand \U$94 ( \437 , RIbb2bf38_118, RIbb32ec8_182);
not \U$95 ( \438 , \437 );
and \U$96 ( \439 , \436 , \438 );
nand \U$97 ( \440 , RIbb2bfb0_117, RIbb32e50_181);
not \U$98 ( \441 , \440 );
nor \U$99 ( \442 , \439 , \441 );
nand \U$100 ( \443 , \435 , \442 );
not \U$101 ( \444 , RIbb2c0a0_115);
not \U$102 ( \445 , RIbb32d60_179);
and \U$103 ( \446 , \444 , \445 );
nor \U$104 ( \447 , RIbb2c028_116, RIbb32dd8_180);
nor \U$105 ( \448 , \446 , \447 );
nor \U$106 ( \449 , RIbb2c118_114, RIbb32ce8_178);
nor \U$107 ( \450 , RIbb2c190_113, RIbb32c70_177);
nor \U$108 ( \451 , \449 , \450 );
nand \U$109 ( \452 , \448 , \451 );
not \U$110 ( \453 , \452 );
nand \U$111 ( \454 , \443 , \453 );
not \U$112 ( \455 , \454 );
nor \U$113 ( \456 , RIbb2be48_120, RIbb32fb8_184);
not \U$114 ( \457 , \456 );
nand \U$115 ( \458 , \419 , \457 , \431 , \427 );
nor \U$116 ( \459 , \458 , \452 );
nor \U$117 ( \460 , RIbb2bbf0_125, RIbb33210_189);
nor \U$118 ( \461 , RIbb2bb78_126, RIbb33288_190);
nor \U$119 ( \462 , \460 , \461 );
not \U$120 ( \463 , \462 );
nand \U$121 ( \464 , RIbb31578_128, RIbb33378_192);
nor \U$122 ( \465 , RIbb31500_127, RIbb33300_191);
or \U$123 ( \466 , \464 , \465 );
nand \U$124 ( \467 , RIbb31500_127, RIbb33300_191);
nand \U$125 ( \468 , \466 , \467 );
not \U$126 ( \469 , \468 );
or \U$127 ( \470 , \463 , \469 );
not \U$128 ( \471 , \460 );
nand \U$129 ( \472 , RIbb2bb78_126, RIbb33288_190);
not \U$130 ( \473 , \472 );
and \U$131 ( \474 , \471 , \473 );
nand \U$132 ( \475 , RIbb2bbf0_125, RIbb33210_189);
not \U$133 ( \476 , \475 );
nor \U$134 ( \477 , \474 , \476 );
nand \U$135 ( \478 , \470 , \477 );
not \U$136 ( \479 , RIbb2bce0_123);
not \U$137 ( \480 , RIbb33120_187);
and \U$138 ( \481 , \479 , \480 );
nor \U$139 ( \482 , RIbb2bc68_124, RIbb33198_188);
nor \U$140 ( \483 , \481 , \482 );
not \U$141 ( \484 , RIbb2bdd0_121);
not \U$142 ( \485 , RIbb33030_185);
nand \U$143 ( \486 , \484 , \485 );
not \U$144 ( \487 , RIbb2bd58_122);
not \U$145 ( \488 , RIbb330a8_186);
nand \U$146 ( \489 , \487 , \488 );
and \U$147 ( \490 , \483 , \486 , \489 );
nand \U$148 ( \491 , \459 , \478 , \490 );
not \U$149 ( \492 , \491 );
or \U$150 ( \493 , \455 , \492 );
nor \U$151 ( \494 , RIbb2c370_109, RIbb32a90_173);
not \U$152 ( \495 , \494 );
not \U$153 ( \496 , \495 );
not \U$154 ( \497 , RIbb2c280_111);
not \U$155 ( \498 , RIbb32b80_175);
nand \U$156 ( \499 , \497 , \498 );
not \U$157 ( \500 , \499 );
nor \U$158 ( \501 , \496 , \500 );
nor \U$159 ( \502 , RIbb2c460_107, RIbb329a0_171);
nor \U$160 ( \503 , RIbb2c550_105, RIbb328b0_169);
nor \U$161 ( \504 , \502 , \503 );
not \U$162 ( \505 , RIbb2c2f8_110);
not \U$163 ( \506 , RIbb32b08_174);
nand \U$164 ( \507 , \505 , \506 );
not \U$165 ( \508 , \507 );
nor \U$166 ( \509 , RIbb2c3e8_108, RIbb32a18_172);
nor \U$167 ( \510 , \508 , \509 );
nor \U$168 ( \511 , RIbb2c208_112, RIbb32bf8_176);
nor \U$169 ( \512 , RIbb2c4d8_106, RIbb32928_170);
nor \U$170 ( \513 , \511 , \512 );
and \U$171 ( \514 , \501 , \504 , \510 , \513 );
not \U$172 ( \515 , RIbb2c640_103);
not \U$173 ( \516 , RIbb327c0_167);
and \U$174 ( \517 , \515 , \516 );
nor \U$175 ( \518 , RIbb2c5c8_104, RIbb32838_168);
nor \U$176 ( \519 , \517 , \518 );
nor \U$177 ( \520 , RIbb2c6b8_102, RIbb32748_166);
nor \U$178 ( \521 , RIbb2c730_101, RIbb326d0_165);
nor \U$179 ( \522 , \520 , \521 );
nand \U$180 ( \523 , \519 , \522 );
not \U$181 ( \524 , \523 );
nor \U$182 ( \525 , RIbb2c898_98, RIbb32568_162);
nor \U$183 ( \526 , RIbb2c910_97, RIbb324f0_161);
nor \U$184 ( \527 , \525 , \526 );
nor \U$185 ( \528 , RIbb2c7a8_100, RIbb32658_164);
nor \U$186 ( \529 , RIbb2c820_99, RIbb325e0_163);
nor \U$187 ( \530 , \528 , \529 );
nand \U$188 ( \531 , \527 , \530 );
not \U$189 ( \532 , \531 );
and \U$190 ( \533 , \514 , \524 , \532 );
nand \U$191 ( \534 , \493 , \533 );
and \U$192 ( \535 , RIbb2c208_112, RIbb32bf8_176);
nand \U$193 ( \536 , \499 , \535 );
not \U$194 ( \537 , \536 );
nand \U$195 ( \538 , RIbb2c2f8_110, RIbb32b08_174);
nand \U$196 ( \539 , RIbb2c370_109, RIbb32a90_173);
nand \U$197 ( \540 , RIbb2c280_111, RIbb32b80_175);
and \U$198 ( \541 , \538 , \539 , \540 );
not \U$199 ( \542 , \541 );
or \U$200 ( \543 , \537 , \542 );
not \U$201 ( \544 , \507 );
not \U$202 ( \545 , \495 );
or \U$203 ( \546 , \544 , \545 );
nand \U$204 ( \547 , \546 , \539 );
nand \U$205 ( \548 , \543 , \547 );
not \U$206 ( \549 , \548 );
not \U$207 ( \550 , \451 );
nand \U$208 ( \551 , RIbb2c028_116, RIbb32dd8_180);
not \U$209 ( \552 , \551 );
not \U$210 ( \553 , \552 );
not \U$211 ( \554 , RIbb2c0a0_115);
not \U$212 ( \555 , RIbb32d60_179);
nand \U$213 ( \556 , \554 , \555 );
not \U$214 ( \557 , \556 );
or \U$215 ( \558 , \553 , \557 );
nand \U$216 ( \559 , RIbb2c0a0_115, RIbb32d60_179);
nand \U$217 ( \560 , \558 , \559 );
not \U$218 ( \561 , \560 );
or \U$219 ( \562 , \550 , \561 );
buf \U$220 ( \563 , \450 );
not \U$221 ( \564 , \563 );
nand \U$222 ( \565 , RIbb2c118_114, RIbb32ce8_178);
not \U$223 ( \566 , \565 );
and \U$224 ( \567 , \564 , \566 );
and \U$225 ( \568 , RIbb2c190_113, RIbb32c70_177);
nor \U$226 ( \569 , \567 , \568 );
nand \U$227 ( \570 , \562 , \569 );
nor \U$228 ( \571 , \549 , \570 );
not \U$229 ( \572 , \571 );
nor \U$230 ( \573 , RIbb2bdd0_121, RIbb33030_185);
nor \U$231 ( \574 , RIbb2bd58_122, RIbb330a8_186);
nor \U$232 ( \575 , \573 , \574 );
not \U$233 ( \576 , \575 );
nand \U$234 ( \577 , RIbb2bc68_124, RIbb33198_188);
nor \U$235 ( \578 , RIbb2bce0_123, RIbb33120_187);
or \U$236 ( \579 , \577 , \578 );
nand \U$237 ( \580 , RIbb2bce0_123, RIbb33120_187);
nand \U$238 ( \581 , \579 , \580 );
not \U$239 ( \582 , \581 );
or \U$240 ( \583 , \576 , \582 );
nand \U$241 ( \584 , RIbb2bd58_122, RIbb330a8_186);
not \U$242 ( \585 , \584 );
and \U$243 ( \586 , \486 , \585 );
nand \U$244 ( \587 , RIbb2bdd0_121, RIbb33030_185);
not \U$245 ( \588 , \587 );
nor \U$246 ( \589 , \586 , \588 );
nand \U$247 ( \590 , \583 , \589 );
not \U$248 ( \591 , \458 );
nand \U$249 ( \592 , \590 , \591 , \453 );
not \U$250 ( \593 , \592 );
or \U$251 ( \594 , \572 , \593 );
not \U$252 ( \595 , \500 );
not \U$253 ( \596 , \511 );
nand \U$254 ( \597 , \595 , \495 , \507 , \596 );
nand \U$255 ( \598 , \548 , \597 );
nor \U$256 ( \599 , \523 , \531 );
not \U$257 ( \600 , \502 );
or \U$258 ( \601 , RIbb2c3e8_108, RIbb32a18_172);
nand \U$259 ( \602 , \600 , \601 );
or \U$260 ( \603 , RIbb2c550_105, RIbb328b0_169);
not \U$261 ( \604 , RIbb2c4d8_106);
not \U$262 ( \605 , RIbb32928_170);
nand \U$263 ( \606 , \604 , \605 );
nand \U$264 ( \607 , \603 , \606 );
nor \U$265 ( \608 , \602 , \607 );
and \U$266 ( \609 , \598 , \599 , \608 );
nand \U$267 ( \610 , \594 , \609 );
not \U$268 ( \611 , \532 );
not \U$269 ( \612 , \522 );
nand \U$270 ( \613 , RIbb2c5c8_104, RIbb32838_168);
not \U$271 ( \614 , \613 );
not \U$272 ( \615 , \614 );
or \U$273 ( \616 , RIbb2c640_103, RIbb327c0_167);
not \U$274 ( \617 , \616 );
or \U$275 ( \618 , \615 , \617 );
nand \U$276 ( \619 , RIbb2c640_103, RIbb327c0_167);
nand \U$277 ( \620 , \618 , \619 );
not \U$278 ( \621 , \620 );
or \U$279 ( \622 , \612 , \621 );
not \U$280 ( \623 , \521 );
nand \U$281 ( \624 , RIbb2c6b8_102, RIbb32748_166);
not \U$282 ( \625 , \624 );
and \U$283 ( \626 , \623 , \625 );
and \U$284 ( \627 , RIbb2c730_101, RIbb326d0_165);
nor \U$285 ( \628 , \626 , \627 );
nand \U$286 ( \629 , \622 , \628 );
not \U$287 ( \630 , \629 );
or \U$288 ( \631 , \611 , \630 );
buf \U$289 ( \632 , \529 );
nand \U$290 ( \633 , RIbb2c7a8_100, RIbb32658_164);
or \U$291 ( \634 , \632 , \633 );
nand \U$292 ( \635 , RIbb2c820_99, RIbb325e0_163);
nand \U$293 ( \636 , \634 , \635 );
and \U$294 ( \637 , \636 , \527 );
nand \U$295 ( \638 , RIbb2c898_98, RIbb32568_162);
or \U$296 ( \639 , \526 , \638 );
nand \U$297 ( \640 , RIbb2c910_97, RIbb324f0_161);
nand \U$298 ( \641 , \639 , \640 );
nor \U$299 ( \642 , \637 , \641 );
nand \U$300 ( \643 , \631 , \642 );
not \U$301 ( \644 , \643 );
not \U$302 ( \645 , \607 );
not \U$303 ( \646 , \645 );
nand \U$304 ( \647 , RIbb2c3e8_108, RIbb32a18_172);
not \U$305 ( \648 , \647 );
not \U$306 ( \649 , \648 );
not \U$307 ( \650 , \600 );
or \U$308 ( \651 , \649 , \650 );
nand \U$309 ( \652 , RIbb2c460_107, RIbb329a0_171);
nand \U$310 ( \653 , \651 , \652 );
not \U$311 ( \654 , \653 );
or \U$312 ( \655 , \646 , \654 );
not \U$313 ( \656 , \605 );
nand \U$314 ( \657 , \656 , RIbb2c4d8_106);
not \U$315 ( \658 , \657 );
and \U$316 ( \659 , \603 , \658 );
and \U$317 ( \660 , RIbb2c550_105, RIbb328b0_169);
nor \U$318 ( \661 , \659 , \660 );
nand \U$319 ( \662 , \655 , \661 );
nand \U$320 ( \663 , \599 , \662 );
nand \U$321 ( \664 , \534 , \610 , \644 , \663 );
buf \U$322 ( \665 , \664 );
not \U$323 ( \666 , \665 );
not \U$324 ( \667 , \666 );
not \U$325 ( \668 , \667 );
or \U$326 ( \669 , \414 , \668 );
nand \U$327 ( \670 , RIbb2caf0_93, RIbb32310_157);
nand \U$328 ( \671 , RIbb2ca78_94, RIbb32388_158);
nand \U$329 ( \672 , RIbb2ca00_95, RIbb32400_159);
nand \U$330 ( \673 , \670 , \671 , \672 );
not \U$331 ( \674 , \673 );
not \U$332 ( \675 , \375 );
nand \U$333 ( \676 , \675 , RIbb2c988_96, RIbb32478_160);
nand \U$334 ( \677 , \674 , \676 );
not \U$335 ( \678 , \677 );
not \U$336 ( \679 , \670 );
nor \U$337 ( \680 , \374 , \679 );
nor \U$338 ( \681 , \379 , \383 );
not \U$339 ( \682 , RIbb2cbe0_91);
not \U$340 ( \683 , RIbb32220_155);
and \U$341 ( \684 , \682 , \683 );
nor \U$342 ( \685 , \684 , \380 );
nand \U$343 ( \686 , \681 , \685 );
nor \U$344 ( \687 , \680 , \686 );
not \U$345 ( \688 , \687 );
or \U$346 ( \689 , \678 , \688 );
nand \U$347 ( \690 , RIbb2cb68_92, RIbb32298_156);
or \U$348 ( \691 , \382 , \690 );
nand \U$349 ( \692 , RIbb2cbe0_91, RIbb32220_155);
nand \U$350 ( \693 , \691 , \692 );
and \U$351 ( \694 , \693 , \381 );
nand \U$352 ( \695 , RIbb2cc58_90, RIbb321a8_154);
or \U$353 ( \696 , \380 , \695 );
nand \U$354 ( \697 , RIbb2ccd0_89, RIbb32130_153);
nand \U$355 ( \698 , \696 , \697 );
nor \U$356 ( \699 , \694 , \698 );
nand \U$357 ( \700 , \689 , \699 );
not \U$358 ( \701 , \700 );
nor \U$359 ( \702 , \370 , \393 );
not \U$360 ( \703 , \702 );
or \U$361 ( \704 , \701 , \703 );
nor \U$362 ( \705 , RIbb2ceb0_85, RIbb31f50_149);
nor \U$363 ( \706 , \705 , \391 );
not \U$364 ( \707 , \706 );
nand \U$365 ( \708 , RIbb2cd48_88, RIbb320b8_152);
or \U$366 ( \709 , \387 , \708 );
nand \U$367 ( \710 , RIbb2cdc0_87, RIbb32040_151);
nand \U$368 ( \711 , \709 , \710 );
not \U$369 ( \712 , \711 );
or \U$370 ( \713 , \707 , \712 );
and \U$371 ( \714 , RIbb2ce38_86, RIbb31fc8_150);
and \U$372 ( \715 , \390 , \714 );
and \U$373 ( \716 , RIbb2ceb0_85, RIbb31f50_149);
nor \U$374 ( \717 , \715 , \716 );
nand \U$375 ( \718 , \713 , \717 );
and \U$376 ( \719 , \371 , \718 );
not \U$377 ( \720 , \369 );
and \U$378 ( \721 , RIbb2cf28_84, RIbb31ed8_148);
not \U$379 ( \722 , \721 );
or \U$380 ( \723 , RIbb2cfa0_83, RIbb31e60_147);
not \U$381 ( \724 , \723 );
or \U$382 ( \725 , \722 , \724 );
nand \U$383 ( \726 , RIbb2cfa0_83, RIbb31e60_147);
nand \U$384 ( \727 , \725 , \726 );
not \U$385 ( \728 , \727 );
or \U$386 ( \729 , \720 , \728 );
not \U$387 ( \730 , \367 );
nand \U$388 ( \731 , RIbb2d018_82, RIbb31de8_146);
not \U$389 ( \732 , \731 );
and \U$390 ( \733 , \730 , \732 );
and \U$391 ( \734 , RIbb2d090_81, RIbb31d70_145);
nor \U$392 ( \735 , \733 , \734 );
nand \U$393 ( \736 , \729 , \735 );
nor \U$394 ( \737 , \719 , \736 );
nand \U$395 ( \738 , \704 , \737 );
buf \U$396 ( \739 , \738 );
nor \U$397 ( \740 , \412 , \359 );
and \U$398 ( \741 , \739 , \740 );
not \U$399 ( \742 , \360 );
not \U$400 ( \743 , \404 );
nor \U$401 ( \744 , RIbb2d270_77, RIbb31b90_141);
nor \U$402 ( \745 , RIbb2d1f8_78, RIbb31c08_142);
nor \U$403 ( \746 , \744 , \745 );
not \U$404 ( \747 , \746 );
nand \U$405 ( \748 , RIbb2d108_80, RIbb31cf8_144);
or \U$406 ( \749 , \405 , \748 );
nand \U$407 ( \750 , RIbb2d180_79, RIbb31c80_143);
nand \U$408 ( \751 , \749 , \750 );
not \U$409 ( \752 , \751 );
or \U$410 ( \753 , \747 , \752 );
nand \U$411 ( \754 , RIbb2d1f8_78, RIbb31c08_142);
not \U$412 ( \755 , \754 );
and \U$413 ( \756 , \408 , \755 );
and \U$414 ( \757 , RIbb2d270_77, RIbb31b90_141);
nor \U$415 ( \758 , \756 , \757 );
nand \U$416 ( \759 , \753 , \758 );
not \U$417 ( \760 , \759 );
or \U$418 ( \761 , \743 , \760 );
nand \U$419 ( \762 , RIbb2d2e8_76, RIbb31b18_140);
not \U$420 ( \763 , \762 );
not \U$421 ( \764 , \763 );
not \U$422 ( \765 , \398 );
not \U$423 ( \766 , \765 );
or \U$424 ( \767 , \764 , \766 );
nand \U$425 ( \768 , RIbb2d360_75, RIbb31aa0_139);
nand \U$426 ( \769 , \767 , \768 );
and \U$427 ( \770 , \769 , \403 );
nand \U$428 ( \771 , RIbb2d3d8_74, RIbb31a28_138);
or \U$429 ( \772 , \402 , \771 );
nand \U$430 ( \773 , RIbb2d450_73, RIbb319b0_137);
nand \U$431 ( \774 , \772 , \773 );
nor \U$432 ( \775 , \770 , \774 );
nand \U$433 ( \776 , \761 , \775 );
not \U$434 ( \777 , \776 );
or \U$435 ( \778 , \742 , \777 );
not \U$436 ( \779 , \346 );
nand \U$437 ( \780 , RIbb2d4c8_72, RIbb31938_136);
or \U$438 ( \781 , \780 , \347 );
nand \U$439 ( \782 , RIbb2d540_71, RIbb318c0_135);
nand \U$440 ( \783 , \781 , \782 );
not \U$441 ( \784 , \783 );
or \U$442 ( \785 , \779 , \784 );
not \U$443 ( \786 , \344 );
nand \U$444 ( \787 , RIbb2d5b8_70, RIbb31848_134);
not \U$445 ( \788 , \787 );
and \U$446 ( \789 , \786 , \788 );
and \U$447 ( \790 , RIbb2d630_69, RIbb317d0_133);
nor \U$448 ( \791 , \789 , \790 );
nand \U$449 ( \792 , \785 , \791 );
and \U$450 ( \793 , \358 , \792 );
and \U$451 ( \794 , RIbb2d6a8_68, RIbb31758_132);
not \U$452 ( \795 , \794 );
not \U$453 ( \796 , \351 );
or \U$454 ( \797 , \795 , \796 );
nand \U$455 ( \798 , RIbb2d720_67, RIbb316e0_131);
nand \U$456 ( \799 , \797 , \798 );
not \U$457 ( \800 , \357 );
and \U$458 ( \801 , \799 , \800 );
not \U$459 ( \802 , \356 );
nand \U$460 ( \803 , RIbb2d798_66, RIbb31668_130);
or \U$461 ( \804 , \802 , \803 );
nand \U$462 ( \805 , RIbb2d810_65, RIbb315f0_129);
nand \U$463 ( \806 , \804 , \805 );
nor \U$464 ( \807 , \793 , \801 , \806 );
nand \U$465 ( \808 , \778 , \807 );
nor \U$466 ( \809 , \741 , \808 );
nand \U$467 ( \810 , \669 , \809 );
buf \U$468 ( \811 , \810 );
not \U$469 ( \812 , \811 );
buf \U$470 ( \813 , \812 );
buf \U$471 ( \814 , \813 );
not \U$472 ( \815 , \814 );
not \U$473 ( \816 , RIbb2ee90_17);
or \U$474 ( \817 , \815 , \816 );
or \U$475 ( \818 , \814 , RIbb2ee90_17);
nand \U$476 ( \819 , \817 , \818 );
not \U$477 ( \820 , \819 );
or \U$478 ( \821 , RIbb2ee90_17, RIbb2ee18_18);
not \U$479 ( \822 , RIbb2ee90_17);
not \U$480 ( \823 , RIbb2ee18_18);
or \U$481 ( \824 , \822 , \823 );
and \U$482 ( \825 , RIbb2eda0_19, \823 );
not \U$483 ( \826 , RIbb2eda0_19);
and \U$484 ( \827 , \826 , RIbb2ee18_18);
nor \U$485 ( \828 , \825 , \827 );
nand \U$486 ( \829 , \821 , \824 , \828 );
not \U$487 ( \830 , \829 );
buf \U$488 ( \831 , \830 );
buf \U$489 ( \832 , \831 );
not \U$490 ( \833 , \832 );
or \U$491 ( \834 , \820 , \833 );
not \U$492 ( \835 , \828 );
buf \U$493 ( \836 , \835 );
not \U$494 ( \837 , \836 );
or \U$495 ( \838 , \837 , \822 );
nand \U$496 ( \839 , \834 , \838 );
not \U$497 ( \840 , \839 );
and \U$498 ( \841 , RIbb2ed28_20, RIbb2eda0_19);
not \U$499 ( \842 , RIbb2ed28_20);
not \U$500 ( \843 , RIbb2eda0_19);
and \U$501 ( \844 , \842 , \843 );
nor \U$502 ( \845 , \841 , \844 );
not \U$503 ( \846 , \845 );
and \U$504 ( \847 , RIbb2ed28_20, RIbb2ecb0_21);
not \U$505 ( \848 , RIbb2ed28_20);
not \U$506 ( \849 , RIbb2ecb0_21);
and \U$507 ( \850 , \848 , \849 );
nor \U$508 ( \851 , \847 , \850 );
nor \U$509 ( \852 , \846 , \851 );
buf \U$510 ( \853 , \852 );
buf \U$511 ( \854 , \851 );
buf \U$512 ( \855 , \854 );
or \U$513 ( \856 , \853 , \855 );
nand \U$514 ( \857 , \856 , RIbb2eda0_19);
not \U$515 ( \858 , \832 );
not \U$516 ( \859 , RIbb2ee90_17);
not \U$517 ( \860 , \412 );
nor \U$518 ( \861 , \353 , \354 );
and \U$519 ( \862 , \350 , \861 );
nand \U$520 ( \863 , \860 , \862 );
nor \U$521 ( \864 , \397 , \863 );
not \U$522 ( \865 , \864 );
buf \U$523 ( \866 , \664 );
buf \U$524 ( \867 , \866 );
not \U$525 ( \868 , \867 );
or \U$526 ( \869 , \865 , \868 );
not \U$527 ( \870 , \863 );
not \U$528 ( \871 , \870 );
not \U$529 ( \872 , \739 );
or \U$530 ( \873 , \871 , \872 );
and \U$531 ( \874 , \776 , \862 );
not \U$532 ( \875 , \861 );
not \U$533 ( \876 , \792 );
or \U$534 ( \877 , \875 , \876 );
and \U$535 ( \878 , \799 , \355 );
not \U$536 ( \879 , \803 );
nor \U$537 ( \880 , \878 , \879 );
nand \U$538 ( \881 , \877 , \880 );
nor \U$539 ( \882 , \874 , \881 );
nand \U$540 ( \883 , \873 , \882 );
not \U$541 ( \884 , \883 );
nand \U$542 ( \885 , \869 , \884 );
nand \U$543 ( \886 , \356 , \805 );
not \U$544 ( \887 , \886 );
and \U$545 ( \888 , \885 , \887 );
not \U$546 ( \889 , \885 );
and \U$547 ( \890 , \889 , \886 );
nor \U$548 ( \891 , \888 , \890 );
buf \U$549 ( \892 , \891 );
buf \U$550 ( \893 , \892 );
not \U$551 ( \894 , \893 );
buf \U$552 ( \895 , \894 );
and \U$553 ( \896 , \859 , \895 );
not \U$554 ( \897 , \859 );
not \U$555 ( \898 , \895 );
and \U$556 ( \899 , \897 , \898 );
nor \U$557 ( \900 , \896 , \899 );
not \U$558 ( \901 , \900 );
or \U$559 ( \902 , \858 , \901 );
nand \U$560 ( \903 , \819 , \836 );
nand \U$561 ( \904 , \902 , \903 );
xor \U$562 ( \905 , \857 , \904 );
not \U$563 ( \906 , RIbb2f070_13);
not \U$564 ( \907 , RIbb2eff8_14);
and \U$565 ( \908 , \906 , \907 );
and \U$566 ( \909 , RIbb2f070_13, RIbb2eff8_14);
nor \U$567 ( \910 , \908 , \909 );
and \U$568 ( \911 , RIbb2ef80_15, \907 );
not \U$569 ( \912 , RIbb2ef80_15);
and \U$570 ( \913 , \912 , RIbb2eff8_14);
nor \U$571 ( \914 , \911 , \913 );
and \U$572 ( \915 , \910 , \914 );
buf \U$573 ( \916 , \915 );
not \U$574 ( \917 , \916 );
not \U$575 ( \918 , RIbb2f070_13);
not \U$576 ( \919 , \412 );
not \U$577 ( \920 , \345 );
nand \U$578 ( \921 , \349 , \920 );
not \U$579 ( \922 , \921 );
nand \U$580 ( \923 , \919 , \922 );
nor \U$581 ( \924 , \395 , \923 );
not \U$582 ( \925 , \924 );
not \U$583 ( \926 , \665 );
or \U$584 ( \927 , \925 , \926 );
nor \U$585 ( \928 , \412 , \921 );
not \U$586 ( \929 , \928 );
not \U$587 ( \930 , \739 );
or \U$588 ( \931 , \929 , \930 );
not \U$589 ( \932 , \404 );
not \U$590 ( \933 , \759 );
or \U$591 ( \934 , \932 , \933 );
nand \U$592 ( \935 , \934 , \775 );
and \U$593 ( \936 , \935 , \922 );
not \U$594 ( \937 , \783 );
or \U$595 ( \938 , \937 , \345 );
nand \U$596 ( \939 , \938 , \787 );
nor \U$597 ( \940 , \936 , \939 );
nand \U$598 ( \941 , \931 , \940 );
not \U$599 ( \942 , \941 );
nand \U$600 ( \943 , \927 , \942 );
nor \U$601 ( \944 , \344 , \790 );
and \U$602 ( \945 , \943 , \944 );
not \U$603 ( \946 , \943 );
not \U$604 ( \947 , \944 );
and \U$605 ( \948 , \946 , \947 );
nor \U$606 ( \949 , \945 , \948 );
buf \U$607 ( \950 , \949 );
not \U$608 ( \951 , \950 );
not \U$609 ( \952 , \951 );
not \U$610 ( \953 , \952 );
not \U$611 ( \954 , \953 );
or \U$612 ( \955 , \918 , \954 );
buf \U$613 ( \956 , \950 );
buf \U$614 ( \957 , \956 );
nand \U$615 ( \958 , \957 , \906 );
nand \U$616 ( \959 , \955 , \958 );
not \U$617 ( \960 , \959 );
or \U$618 ( \961 , \917 , \960 );
not \U$619 ( \962 , RIbb2f070_13);
nand \U$620 ( \963 , \919 , \350 );
nor \U$621 ( \964 , \397 , \963 );
not \U$622 ( \965 , \964 );
not \U$623 ( \966 , \866 );
or \U$624 ( \967 , \965 , \966 );
not \U$625 ( \968 , \350 );
nor \U$626 ( \969 , \968 , \412 );
and \U$627 ( \970 , \969 , \739 );
not \U$628 ( \971 , \350 );
not \U$629 ( \972 , \935 );
or \U$630 ( \973 , \971 , \972 );
not \U$631 ( \974 , \792 );
nand \U$632 ( \975 , \973 , \974 );
nor \U$633 ( \976 , \970 , \975 );
nand \U$634 ( \977 , \967 , \976 );
not \U$635 ( \978 , \794 );
nand \U$636 ( \979 , \352 , \978 );
not \U$637 ( \980 , \979 );
and \U$638 ( \981 , \977 , \980 );
not \U$639 ( \982 , \977 );
and \U$640 ( \983 , \982 , \979 );
nor \U$641 ( \984 , \981 , \983 );
not \U$642 ( \985 , \984 );
not \U$643 ( \986 , \985 );
buf \U$644 ( \987 , \986 );
not \U$645 ( \988 , \987 );
buf \U$646 ( \989 , \988 );
not \U$647 ( \990 , \989 );
or \U$648 ( \991 , \962 , \990 );
not \U$649 ( \992 , \986 );
buf \U$650 ( \993 , \992 );
not \U$651 ( \994 , \993 );
nand \U$652 ( \995 , \994 , \906 );
nand \U$653 ( \996 , \991 , \995 );
not \U$654 ( \997 , \914 );
buf \U$655 ( \998 , \997 );
nand \U$656 ( \999 , \996 , \998 );
nand \U$657 ( \1000 , \961 , \999 );
and \U$658 ( \1001 , \905 , \1000 );
and \U$659 ( \1002 , \857 , \904 );
or \U$660 ( \1003 , \1001 , \1002 );
xor \U$661 ( \1004 , \840 , \1003 );
xnor \U$662 ( \1005 , RIbb2f160_11, RIbb2f0e8_12);
and \U$663 ( \1006 , RIbb2f0e8_12, RIbb2f070_13);
not \U$664 ( \1007 , RIbb2f0e8_12);
and \U$665 ( \1008 , \1007 , \906 );
nor \U$666 ( \1009 , \1006 , \1008 );
nor \U$667 ( \1010 , \1005 , \1009 );
buf \U$668 ( \1011 , \1010 );
not \U$669 ( \1012 , \1011 );
not \U$670 ( \1013 , RIbb2f160_11);
not \U$671 ( \1014 , \348 );
nand \U$672 ( \1015 , \919 , \1014 );
nor \U$673 ( \1016 , \397 , \1015 );
not \U$674 ( \1017 , \1016 );
not \U$675 ( \1018 , \866 );
or \U$676 ( \1019 , \1017 , \1018 );
nor \U$677 ( \1020 , \412 , \348 );
not \U$678 ( \1021 , \1020 );
not \U$679 ( \1022 , \739 );
or \U$680 ( \1023 , \1021 , \1022 );
and \U$681 ( \1024 , \935 , \1014 );
not \U$682 ( \1025 , \780 );
nor \U$683 ( \1026 , \1024 , \1025 );
nand \U$684 ( \1027 , \1023 , \1026 );
not \U$685 ( \1028 , \1027 );
nand \U$686 ( \1029 , \1019 , \1028 );
not \U$687 ( \1030 , \782 );
nor \U$688 ( \1031 , \1030 , \347 );
and \U$689 ( \1032 , \1029 , \1031 );
not \U$690 ( \1033 , \1029 );
not \U$691 ( \1034 , \1031 );
and \U$692 ( \1035 , \1033 , \1034 );
nor \U$693 ( \1036 , \1032 , \1035 );
buf \U$694 ( \1037 , \1036 );
buf \U$695 ( \1038 , \1037 );
not \U$696 ( \1039 , \1038 );
not \U$697 ( \1040 , \1039 );
or \U$698 ( \1041 , \1013 , \1040 );
not \U$699 ( \1042 , \1039 );
not \U$700 ( \1043 , RIbb2f160_11);
nand \U$701 ( \1044 , \1042 , \1043 );
nand \U$702 ( \1045 , \1041 , \1044 );
not \U$703 ( \1046 , \1045 );
or \U$704 ( \1047 , \1012 , \1046 );
not \U$705 ( \1048 , RIbb2f160_11);
not \U$706 ( \1049 , \349 );
nor \U$707 ( \1050 , \411 , \1049 );
and \U$708 ( \1051 , \396 , \1050 );
not \U$709 ( \1052 , \1051 );
not \U$710 ( \1053 , \866 );
or \U$711 ( \1054 , \1052 , \1053 );
nor \U$712 ( \1055 , \412 , \1049 );
and \U$713 ( \1056 , \739 , \1055 );
not \U$714 ( \1057 , \349 );
not \U$715 ( \1058 , \935 );
or \U$716 ( \1059 , \1057 , \1058 );
nand \U$717 ( \1060 , \1059 , \937 );
nor \U$718 ( \1061 , \1056 , \1060 );
nand \U$719 ( \1062 , \1054 , \1061 );
nand \U$720 ( \1063 , \920 , \787 );
not \U$721 ( \1064 , \1063 );
and \U$722 ( \1065 , \1062 , \1064 );
not \U$723 ( \1066 , \1062 );
and \U$724 ( \1067 , \1066 , \1063 );
nor \U$725 ( \1068 , \1065 , \1067 );
not \U$726 ( \1069 , \1068 );
buf \U$727 ( \1070 , \1069 );
not \U$728 ( \1071 , \1070 );
not \U$729 ( \1072 , \1071 );
and \U$730 ( \1073 , \1048 , \1072 );
not \U$731 ( \1074 , \1048 );
and \U$732 ( \1075 , \1074 , \1071 );
nor \U$733 ( \1076 , \1073 , \1075 );
buf \U$734 ( \1077 , \1009 );
nand \U$735 ( \1078 , \1076 , \1077 );
nand \U$736 ( \1079 , \1047 , \1078 );
not \U$737 ( \1080 , RIbb2f3b8_6);
and \U$738 ( \1081 , RIbb2f340_7, \1080 );
not \U$739 ( \1082 , RIbb2f340_7);
and \U$740 ( \1083 , \1082 , RIbb2f3b8_6);
nor \U$741 ( \1084 , \1081 , \1083 );
not \U$742 ( \1085 , RIbb2f430_5);
and \U$743 ( \1086 , \1085 , \1080 );
and \U$744 ( \1087 , RIbb2f430_5, RIbb2f3b8_6);
nor \U$745 ( \1088 , \1086 , \1087 );
and \U$746 ( \1089 , \1084 , \1088 );
buf \U$747 ( \1090 , \1089 );
not \U$748 ( \1091 , \1090 );
not \U$749 ( \1092 , \407 );
nor \U$750 ( \1093 , \1092 , \745 );
and \U$751 ( \1094 , \396 , \1093 );
not \U$752 ( \1095 , \1094 );
not \U$753 ( \1096 , \665 );
or \U$754 ( \1097 , \1095 , \1096 );
and \U$755 ( \1098 , \739 , \1093 );
not \U$756 ( \1099 , \751 );
or \U$757 ( \1100 , \1099 , \745 );
nand \U$758 ( \1101 , \1100 , \754 );
nor \U$759 ( \1102 , \1098 , \1101 );
nand \U$760 ( \1103 , \1097 , \1102 );
nor \U$761 ( \1104 , \744 , \757 );
and \U$762 ( \1105 , \1103 , \1104 );
not \U$763 ( \1106 , \1103 );
not \U$764 ( \1107 , \1104 );
and \U$765 ( \1108 , \1106 , \1107 );
nor \U$766 ( \1109 , \1105 , \1108 );
not \U$767 ( \1110 , \1109 );
not \U$768 ( \1111 , \1110 );
not \U$769 ( \1112 , \1111 );
buf \U$770 ( \1113 , \1112 );
not \U$771 ( \1114 , \1113 );
and \U$772 ( \1115 , RIbb2f430_5, \1114 );
not \U$773 ( \1116 , RIbb2f430_5);
and \U$774 ( \1117 , \1116 , \1113 );
nor \U$775 ( \1118 , \1115 , \1117 );
not \U$776 ( \1119 , \1118 );
or \U$777 ( \1120 , \1091 , \1119 );
and \U$778 ( \1121 , \396 , \410 );
not \U$779 ( \1122 , \1121 );
not \U$780 ( \1123 , \866 );
or \U$781 ( \1124 , \1122 , \1123 );
and \U$782 ( \1125 , \739 , \410 );
nor \U$783 ( \1126 , \1125 , \759 );
nand \U$784 ( \1127 , \1124 , \1126 );
not \U$785 ( \1128 , \399 );
nand \U$786 ( \1129 , \1128 , \762 );
not \U$787 ( \1130 , \1129 );
and \U$788 ( \1131 , \1127 , \1130 );
not \U$789 ( \1132 , \1127 );
and \U$790 ( \1133 , \1132 , \1129 );
nor \U$791 ( \1134 , \1131 , \1133 );
not \U$792 ( \1135 , \1134 );
not \U$793 ( \1136 , \1135 );
buf \U$794 ( \1137 , \1136 );
buf \U$795 ( \1138 , \1137 );
buf \U$796 ( \1139 , \1138 );
not \U$797 ( \1140 , \1139 );
and \U$798 ( \1141 , RIbb2f430_5, \1140 );
not \U$799 ( \1142 , RIbb2f430_5);
and \U$800 ( \1143 , \1142 , \1139 );
nor \U$801 ( \1144 , \1141 , \1143 );
not \U$802 ( \1145 , \1144 );
not \U$803 ( \1146 , \1084 );
buf \U$804 ( \1147 , \1146 );
nand \U$805 ( \1148 , \1145 , \1147 );
nand \U$806 ( \1149 , \1120 , \1148 );
xor \U$807 ( \1150 , \1079 , \1149 );
nor \U$808 ( \1151 , \397 , \406 );
not \U$809 ( \1152 , \1151 );
not \U$810 ( \1153 , \866 );
or \U$811 ( \1154 , \1152 , \1153 );
not \U$812 ( \1155 , \406 );
buf \U$813 ( \1156 , \700 );
nand \U$814 ( \1157 , \371 , \1155 , \1156 , \394 );
nand \U$815 ( \1158 , \371 , \718 , \1155 );
nand \U$816 ( \1159 , \736 , \1155 );
and \U$817 ( \1160 , \1157 , \1158 , \1159 , \748 );
nand \U$818 ( \1161 , \1154 , \1160 );
not \U$819 ( \1162 , \750 );
nor \U$820 ( \1163 , \1162 , \405 );
and \U$821 ( \1164 , \1161 , \1163 );
not \U$822 ( \1165 , \1161 );
not \U$823 ( \1166 , \1163 );
and \U$824 ( \1167 , \1165 , \1166 );
nor \U$825 ( \1168 , \1164 , \1167 );
buf \U$826 ( \1169 , \1168 );
not \U$827 ( \1170 , \1169 );
buf \U$828 ( \1171 , \1170 );
not \U$829 ( \1172 , RIbb2bfb0_117);
not \U$830 ( \1173 , RIbb31500_127);
not \U$831 ( \1174 , RIbb31578_128);
nand \U$832 ( \1175 , \1172 , \1173 , \1174 , RIbb2bb78_126);
nor \U$833 ( \1176 , RIbb2c730_101, RIbb2c6b8_102);
nor \U$834 ( \1177 , RIbb2c640_103, RIbb2c5c8_104);
nand \U$835 ( \1178 , \1176 , \1177 );
nor \U$836 ( \1179 , \1175 , \1178 );
nor \U$837 ( \1180 , RIbb2c550_105, RIbb2c4d8_106);
nor \U$838 ( \1181 , RIbb2c460_107, RIbb2c3e8_108);
nand \U$839 ( \1182 , \1180 , \1181 );
nor \U$840 ( \1183 , RIbb2c370_109, RIbb2c2f8_110);
nor \U$841 ( \1184 , RIbb2c280_111, RIbb2c208_112);
nand \U$842 ( \1185 , \1183 , \1184 );
nor \U$843 ( \1186 , \1182 , \1185 );
and \U$844 ( \1187 , \1179 , \1186 );
not \U$845 ( \1188 , \1187 );
nor \U$846 ( \1189 , RIbb2d090_81, RIbb2d018_82);
nor \U$847 ( \1190 , RIbb2cfa0_83, RIbb2cf28_84);
nor \U$848 ( \1191 , RIbb2ceb0_85, RIbb2ce38_86);
nor \U$849 ( \1192 , RIbb2cdc0_87, RIbb2cd48_88);
nand \U$850 ( \1193 , \1189 , \1190 , \1191 , \1192 );
not \U$851 ( \1194 , \1193 );
nor \U$852 ( \1195 , RIbb2d450_73, RIbb2d3d8_74);
nor \U$853 ( \1196 , RIbb2d360_75, RIbb2d2e8_76);
nand \U$854 ( \1197 , \1195 , \1196 );
nor \U$855 ( \1198 , RIbb2ccd0_89, RIbb2cc58_90);
nor \U$856 ( \1199 , RIbb2cbe0_91, RIbb2cb68_92);
nand \U$857 ( \1200 , \1198 , \1199 );
nor \U$858 ( \1201 , \1197 , \1200 );
nand \U$859 ( \1202 , \1194 , \1201 );
nor \U$860 ( \1203 , \1188 , \1202 );
not \U$861 ( \1204 , \1203 );
not \U$862 ( \1205 , RIbb2bc68_124);
not \U$863 ( \1206 , RIbb2bbf0_125);
nand \U$864 ( \1207 , \1205 , \1206 , RIbb2bd58_122, RIbb2bce0_123);
nor \U$865 ( \1208 , RIbb2c910_97, RIbb2c898_98);
nor \U$866 ( \1209 , RIbb2c820_99, RIbb2c7a8_100);
nand \U$867 ( \1210 , \1208 , \1209 );
nor \U$868 ( \1211 , \1207 , \1210 );
nor \U$869 ( \1212 , RIbb2c190_113, RIbb2c118_114);
nor \U$870 ( \1213 , RIbb2c0a0_115, RIbb2c028_116);
nand \U$871 ( \1214 , \1212 , \1213 );
nand \U$872 ( \1215 , RIbb2bf38_118, RIbb2bec0_119, RIbb2be48_120, RIbb2bdd0_121);
nor \U$873 ( \1216 , \1214 , \1215 );
and \U$874 ( \1217 , \1211 , \1216 );
nor \U$875 ( \1218 , RIbb2d810_65, RIbb2d798_66);
nor \U$876 ( \1219 , RIbb2d720_67, RIbb2d6a8_68);
nor \U$877 ( \1220 , RIbb2d630_69, RIbb2d5b8_70);
nor \U$878 ( \1221 , RIbb2d540_71, RIbb2d4c8_72);
and \U$879 ( \1222 , \1218 , \1219 , \1220 , \1221 );
nor \U$880 ( \1223 , RIbb2d270_77, RIbb2d1f8_78);
nor \U$881 ( \1224 , RIbb2d180_79, RIbb2d108_80);
nand \U$882 ( \1225 , \1223 , \1224 );
nor \U$883 ( \1226 , RIbb2caf0_93, RIbb2ca78_94);
nor \U$884 ( \1227 , RIbb2ca00_95, RIbb2c988_96);
nand \U$885 ( \1228 , \1226 , \1227 );
nor \U$886 ( \1229 , \1225 , \1228 );
nand \U$887 ( \1230 , \1222 , \1229 );
not \U$888 ( \1231 , \1230 );
and \U$889 ( \1232 , \1217 , \1231 , RIbb32fb8_184);
not \U$890 ( \1233 , \1232 );
or \U$891 ( \1234 , \1204 , \1233 );
nand \U$892 ( \1235 , \1217 , \1187 );
and \U$893 ( \1236 , \1235 , RIbb2f520_3);
not \U$894 ( \1237 , \1202 );
and \U$895 ( \1238 , \1237 , \1231 );
not \U$896 ( \1239 , RIbb2f520_3);
nor \U$897 ( \1240 , \1238 , \1239 );
nor \U$898 ( \1241 , \1236 , \1240 );
nand \U$899 ( \1242 , \1234 , \1241 );
not \U$900 ( \1243 , \1242 );
buf \U$901 ( \1244 , \1243 );
buf \U$902 ( \1245 , \1244 );
not \U$903 ( \1246 , \1245 );
and \U$904 ( \1247 , \1171 , \1246 );
not \U$905 ( \1248 , \1171 );
and \U$906 ( \1249 , \1248 , \1245 );
nor \U$907 ( \1250 , \1247 , \1249 );
not \U$908 ( \1251 , RIbb2f4a8_4);
not \U$909 ( \1252 , \1242 );
not \U$910 ( \1253 , \1252 );
not \U$911 ( \1254 , \1253 );
or \U$912 ( \1255 , \1251 , \1254 );
not \U$913 ( \1256 , RIbb2f4a8_4);
and \U$914 ( \1257 , \1243 , \1256 );
and \U$915 ( \1258 , RIbb2f430_5, \1256 );
not \U$916 ( \1259 , RIbb2f430_5);
and \U$917 ( \1260 , \1259 , RIbb2f4a8_4);
or \U$918 ( \1261 , \1258 , \1260 );
nor \U$919 ( \1262 , \1257 , \1261 );
nand \U$920 ( \1263 , \1255 , \1262 );
not \U$921 ( \1264 , \1263 );
buf \U$922 ( \1265 , \1264 );
not \U$923 ( \1266 , \1265 );
or \U$924 ( \1267 , \1250 , \1266 );
and \U$925 ( \1268 , \396 , \407 );
not \U$926 ( \1269 , \1268 );
not \U$927 ( \1270 , \866 );
or \U$928 ( \1271 , \1269 , \1270 );
and \U$929 ( \1272 , \739 , \407 );
nor \U$930 ( \1273 , \1272 , \751 );
nand \U$931 ( \1274 , \1271 , \1273 );
nand \U$932 ( \1275 , \409 , \754 );
not \U$933 ( \1276 , \1275 );
and \U$934 ( \1277 , \1274 , \1276 );
not \U$935 ( \1278 , \1274 );
and \U$936 ( \1279 , \1278 , \1275 );
nor \U$937 ( \1280 , \1277 , \1279 );
not \U$938 ( \1281 , \1280 );
not \U$939 ( \1282 , \1281 );
buf \U$940 ( \1283 , \1282 );
not \U$941 ( \1284 , \1283 );
not \U$942 ( \1285 , \1284 );
not \U$943 ( \1286 , \1285 );
and \U$944 ( \1287 , \1286 , \1246 );
not \U$945 ( \1288 , \1244 );
not \U$946 ( \1289 , \1288 );
not \U$947 ( \1290 , \1289 );
not \U$948 ( \1291 , \1290 );
and \U$949 ( \1292 , \1285 , \1291 );
nor \U$950 ( \1293 , \1287 , \1292 );
buf \U$951 ( \1294 , \1261 );
not \U$952 ( \1295 , \1294 );
or \U$953 ( \1296 , \1293 , \1295 );
nand \U$954 ( \1297 , \1267 , \1296 );
and \U$955 ( \1298 , \1150 , \1297 );
and \U$956 ( \1299 , \1079 , \1149 );
or \U$957 ( \1300 , \1298 , \1299 );
and \U$958 ( \1301 , \1004 , \1300 );
and \U$959 ( \1302 , \840 , \1003 );
or \U$960 ( \1303 , \1301 , \1302 );
buf \U$961 ( \1304 , \1217 );
nand \U$962 ( \1305 , \1304 , \1187 , \1237 , \1231 );
not \U$963 ( \1306 , RIbb2f610_1);
and \U$964 ( \1307 , \1305 , \1306 );
not \U$965 ( \1308 , \1305 );
not \U$966 ( \1309 , RIbb2f598_2);
and \U$967 ( \1310 , \1308 , \1309 );
nor \U$968 ( \1311 , \1307 , \1310 );
buf \U$969 ( \1312 , \1311 );
buf \U$970 ( \1313 , \1312 );
nand \U$971 ( \1314 , \394 , \366 );
buf \U$972 ( \1315 , \386 );
not \U$973 ( \1316 , \1315 );
nor \U$974 ( \1317 , \1314 , \1316 );
not \U$975 ( \1318 , \1317 );
not \U$976 ( \1319 , \665 );
or \U$977 ( \1320 , \1318 , \1319 );
not \U$978 ( \1321 , \1314 );
and \U$979 ( \1322 , \1156 , \1321 );
not \U$980 ( \1323 , \366 );
not \U$981 ( \1324 , \718 );
or \U$982 ( \1325 , \1323 , \1324 );
not \U$983 ( \1326 , \727 );
nand \U$984 ( \1327 , \1325 , \1326 );
nor \U$985 ( \1328 , \1322 , \1327 );
nand \U$986 ( \1329 , \1320 , \1328 );
not \U$987 ( \1330 , \368 );
nand \U$988 ( \1331 , \1330 , \731 );
not \U$989 ( \1332 , \1331 );
and \U$990 ( \1333 , \1329 , \1332 );
not \U$991 ( \1334 , \1329 );
and \U$992 ( \1335 , \1334 , \1331 );
nor \U$993 ( \1336 , \1333 , \1335 );
buf \U$994 ( \1337 , \1336 );
buf \U$995 ( \1338 , \1337 );
buf \U$996 ( \1339 , \1338 );
not \U$997 ( \1340 , \1339 );
not \U$998 ( \1341 , \1340 );
and \U$999 ( \1342 , \1313 , \1341 );
nor \U$1000 ( \1343 , \1210 , \1178 );
buf \U$1001 ( \1344 , \1186 );
nand \U$1002 ( \1345 , \1343 , \1344 );
not \U$1003 ( \1346 , \1193 );
nor \U$1004 ( \1347 , \1200 , \1228 );
nand \U$1005 ( \1348 , \1346 , \1347 );
nor \U$1006 ( \1349 , \1345 , \1348 );
not \U$1007 ( \1350 , \1349 );
nor \U$1008 ( \1351 , \1207 , \1175 );
nand \U$1009 ( \1352 , \1216 , \1351 );
nor \U$1010 ( \1353 , \1197 , \1225 );
nand \U$1011 ( \1354 , \1222 , \1353 );
nor \U$1012 ( \1355 , \1352 , \1354 , \1239 );
not \U$1013 ( \1356 , \1355 );
or \U$1014 ( \1357 , \1350 , \1356 );
not \U$1015 ( \1358 , RIbb2f598_2);
not \U$1016 ( \1359 , \1352 );
or \U$1017 ( \1360 , \1358 , \1359 );
nand \U$1018 ( \1361 , \1345 , RIbb2f598_2);
nand \U$1019 ( \1362 , \1360 , \1361 );
not \U$1020 ( \1363 , RIbb2f598_2);
not \U$1021 ( \1364 , \1348 );
or \U$1022 ( \1365 , \1363 , \1364 );
nand \U$1023 ( \1366 , \1354 , RIbb2f598_2);
nand \U$1024 ( \1367 , \1365 , \1366 );
nor \U$1025 ( \1368 , \1362 , \1367 );
nand \U$1026 ( \1369 , \1357 , \1368 );
not \U$1027 ( \1370 , \1369 );
and \U$1028 ( \1371 , \1370 , \1242 );
not \U$1029 ( \1372 , \1370 );
and \U$1030 ( \1373 , \1372 , \1252 );
nor \U$1031 ( \1374 , \1371 , \1373 );
not \U$1032 ( \1375 , \1374 );
buf \U$1033 ( \1376 , \1375 );
not \U$1034 ( \1377 , \1376 );
not \U$1035 ( \1378 , \396 );
not \U$1036 ( \1379 , \665 );
or \U$1037 ( \1380 , \1378 , \1379 );
not \U$1038 ( \1381 , \739 );
nand \U$1039 ( \1382 , \1380 , \1381 );
and \U$1040 ( \1383 , \1155 , \748 );
xor \U$1041 ( \1384 , \1382 , \1383 );
not \U$1042 ( \1385 , \1384 );
not \U$1043 ( \1386 , \1385 );
buf \U$1044 ( \1387 , \1386 );
xor \U$1045 ( \1388 , \1313 , \1387 );
not \U$1046 ( \1389 , \1388 );
or \U$1047 ( \1390 , \1377 , \1389 );
not \U$1048 ( \1391 , \1311 );
buf \U$1049 ( \1392 , \1391 );
not \U$1050 ( \1393 , \1392 );
buf \U$1051 ( \1394 , \1393 );
not \U$1052 ( \1395 , \366 );
nor \U$1053 ( \1396 , \1395 , \368 );
nand \U$1054 ( \1397 , \1396 , \394 );
nor \U$1055 ( \1398 , \1397 , \1316 );
not \U$1056 ( \1399 , \1398 );
not \U$1057 ( \1400 , \866 );
or \U$1058 ( \1401 , \1399 , \1400 );
not \U$1059 ( \1402 , \1397 );
and \U$1060 ( \1403 , \1156 , \1402 );
not \U$1061 ( \1404 , \1396 );
not \U$1062 ( \1405 , \718 );
or \U$1063 ( \1406 , \1404 , \1405 );
and \U$1064 ( \1407 , \727 , \1330 );
not \U$1065 ( \1408 , \731 );
nor \U$1066 ( \1409 , \1407 , \1408 );
nand \U$1067 ( \1410 , \1406 , \1409 );
nor \U$1068 ( \1411 , \1403 , \1410 );
nand \U$1069 ( \1412 , \1401 , \1411 );
nor \U$1070 ( \1413 , \734 , \367 );
and \U$1071 ( \1414 , \1412 , \1413 );
not \U$1072 ( \1415 , \1412 );
not \U$1073 ( \1416 , \1413 );
and \U$1074 ( \1417 , \1415 , \1416 );
nor \U$1075 ( \1418 , \1414 , \1417 );
buf \U$1076 ( \1419 , \1418 );
not \U$1077 ( \1420 , \1419 );
not \U$1078 ( \1421 , \1420 );
buf \U$1079 ( \1422 , \1421 );
xor \U$1080 ( \1423 , \1394 , \1422 );
and \U$1081 ( \1424 , \1311 , \1370 );
not \U$1082 ( \1425 , \1311 );
and \U$1083 ( \1426 , \1425 , \1369 );
or \U$1084 ( \1427 , \1424 , \1426 );
and \U$1085 ( \1428 , \1427 , \1374 );
buf \U$1086 ( \1429 , \1428 );
buf \U$1087 ( \1430 , \1429 );
nand \U$1088 ( \1431 , \1423 , \1430 );
nand \U$1089 ( \1432 , \1390 , \1431 );
xor \U$1090 ( \1433 , \1342 , \1432 );
and \U$1091 ( \1434 , RIbb2ef08_16, RIbb2ee90_17);
not \U$1092 ( \1435 , RIbb2ef08_16);
and \U$1093 ( \1436 , \1435 , \822 );
nor \U$1094 ( \1437 , \1434 , \1436 );
not \U$1095 ( \1438 , \1437 );
and \U$1096 ( \1439 , RIbb2ef80_15, RIbb2ef08_16);
not \U$1097 ( \1440 , RIbb2ef80_15);
not \U$1098 ( \1441 , RIbb2ef08_16);
and \U$1099 ( \1442 , \1440 , \1441 );
nor \U$1100 ( \1443 , \1439 , \1442 );
and \U$1101 ( \1444 , \1438 , \1443 );
buf \U$1102 ( \1445 , \1444 );
not \U$1103 ( \1446 , \1445 );
not \U$1104 ( \1447 , \412 );
and \U$1105 ( \1448 , \350 , \352 );
nand \U$1106 ( \1449 , \1447 , \1448 );
nor \U$1107 ( \1450 , \397 , \1449 );
not \U$1108 ( \1451 , \1450 );
not \U$1109 ( \1452 , \867 );
or \U$1110 ( \1453 , \1451 , \1452 );
not \U$1111 ( \1454 , \1449 );
not \U$1112 ( \1455 , \1454 );
not \U$1113 ( \1456 , \739 );
or \U$1114 ( \1457 , \1455 , \1456 );
and \U$1115 ( \1458 , \776 , \1448 );
not \U$1116 ( \1459 , \352 );
not \U$1117 ( \1460 , \792 );
or \U$1118 ( \1461 , \1459 , \1460 );
nand \U$1119 ( \1462 , \1461 , \978 );
nor \U$1120 ( \1463 , \1458 , \1462 );
nand \U$1121 ( \1464 , \1457 , \1463 );
not \U$1122 ( \1465 , \1464 );
nand \U$1123 ( \1466 , \1453 , \1465 );
nand \U$1124 ( \1467 , \351 , \798 );
not \U$1125 ( \1468 , \1467 );
and \U$1126 ( \1469 , \1466 , \1468 );
not \U$1127 ( \1470 , \1466 );
and \U$1128 ( \1471 , \1470 , \1467 );
nor \U$1129 ( \1472 , \1469 , \1471 );
not \U$1130 ( \1473 , \1472 );
not \U$1131 ( \1474 , \1473 );
not \U$1132 ( \1475 , \1474 );
not \U$1133 ( \1476 , \1475 );
buf \U$1134 ( \1477 , \1476 );
xor \U$1135 ( \1478 , \1477 , RIbb2ef80_15);
not \U$1136 ( \1479 , \1478 );
or \U$1137 ( \1480 , \1446 , \1479 );
not \U$1138 ( \1481 , \353 );
nand \U$1139 ( \1482 , \350 , \1481 );
not \U$1140 ( \1483 , \1482 );
nand \U$1141 ( \1484 , \919 , \1483 );
nor \U$1142 ( \1485 , \395 , \1484 );
not \U$1143 ( \1486 , \1485 );
not \U$1144 ( \1487 , \665 );
or \U$1145 ( \1488 , \1486 , \1487 );
nor \U$1146 ( \1489 , \412 , \1482 );
not \U$1147 ( \1490 , \1489 );
not \U$1148 ( \1491 , \739 );
or \U$1149 ( \1492 , \1490 , \1491 );
and \U$1150 ( \1493 , \776 , \1483 );
not \U$1151 ( \1494 , \1481 );
not \U$1152 ( \1495 , \792 );
or \U$1153 ( \1496 , \1494 , \1495 );
not \U$1154 ( \1497 , \799 );
nand \U$1155 ( \1498 , \1496 , \1497 );
nor \U$1156 ( \1499 , \1493 , \1498 );
nand \U$1157 ( \1500 , \1492 , \1499 );
not \U$1158 ( \1501 , \1500 );
nand \U$1159 ( \1502 , \1488 , \1501 );
nand \U$1160 ( \1503 , \355 , \803 );
not \U$1161 ( \1504 , \1503 );
and \U$1162 ( \1505 , \1502 , \1504 );
not \U$1163 ( \1506 , \1502 );
and \U$1164 ( \1507 , \1506 , \1503 );
nor \U$1165 ( \1508 , \1505 , \1507 );
not \U$1166 ( \1509 , \1508 );
buf \U$1167 ( \1510 , \1509 );
not \U$1168 ( \1511 , \1510 );
and \U$1169 ( \1512 , RIbb2ef80_15, \1511 );
not \U$1170 ( \1513 , RIbb2ef80_15);
not \U$1171 ( \1514 , \1511 );
and \U$1172 ( \1515 , \1513 , \1514 );
nor \U$1173 ( \1516 , \1512 , \1515 );
buf \U$1174 ( \1517 , \1437 );
nand \U$1175 ( \1518 , \1516 , \1517 );
nand \U$1176 ( \1519 , \1480 , \1518 );
and \U$1177 ( \1520 , \1433 , \1519 );
and \U$1178 ( \1521 , \1342 , \1432 );
or \U$1179 ( \1522 , \1520 , \1521 );
and \U$1180 ( \1523 , \1394 , \1422 );
not \U$1181 ( \1524 , RIbb2f250_9);
not \U$1182 ( \1525 , RIbb2f1d8_10);
and \U$1183 ( \1526 , \1524 , \1525 );
and \U$1184 ( \1527 , RIbb2f250_9, RIbb2f1d8_10);
and \U$1185 ( \1528 , RIbb2f1d8_10, RIbb2f160_11);
not \U$1186 ( \1529 , RIbb2f1d8_10);
and \U$1187 ( \1530 , \1529 , \1048 );
nor \U$1188 ( \1531 , \1528 , \1530 );
nor \U$1189 ( \1532 , \1526 , \1527 , \1531 );
buf \U$1190 ( \1533 , \1532 );
not \U$1191 ( \1534 , \1533 );
nor \U$1192 ( \1535 , \395 , \412 );
not \U$1193 ( \1536 , \1535 );
not \U$1194 ( \1537 , \665 );
or \U$1195 ( \1538 , \1536 , \1537 );
and \U$1196 ( \1539 , \919 , \739 );
nor \U$1197 ( \1540 , \1539 , \776 );
nand \U$1198 ( \1541 , \1538 , \1540 );
nand \U$1199 ( \1542 , \1014 , \780 );
not \U$1200 ( \1543 , \1542 );
and \U$1201 ( \1544 , \1541 , \1543 );
not \U$1202 ( \1545 , \1541 );
and \U$1203 ( \1546 , \1545 , \1542 );
nor \U$1204 ( \1547 , \1544 , \1546 );
buf \U$1205 ( \1548 , \1547 );
not \U$1206 ( \1549 , \1548 );
buf \U$1207 ( \1550 , \1549 );
not \U$1208 ( \1551 , \1550 );
and \U$1209 ( \1552 , \1551 , RIbb2f250_9);
not \U$1210 ( \1553 , \1551 );
not \U$1211 ( \1554 , RIbb2f250_9);
and \U$1212 ( \1555 , \1553 , \1554 );
nor \U$1213 ( \1556 , \1552 , \1555 );
not \U$1214 ( \1557 , \1556 );
or \U$1215 ( \1558 , \1534 , \1557 );
not \U$1216 ( \1559 , \1036 );
not \U$1217 ( \1560 , \1559 );
buf \U$1218 ( \1561 , \1560 );
not \U$1219 ( \1562 , \1561 );
not \U$1220 ( \1563 , \1562 );
and \U$1221 ( \1564 , \1563 , RIbb2f250_9);
not \U$1222 ( \1565 , \1563 );
not \U$1223 ( \1566 , RIbb2f250_9);
and \U$1224 ( \1567 , \1565 , \1566 );
nor \U$1225 ( \1568 , \1564 , \1567 );
buf \U$1226 ( \1569 , \1531 );
buf \U$1227 ( \1570 , \1569 );
nand \U$1228 ( \1571 , \1568 , \1570 );
nand \U$1229 ( \1572 , \1558 , \1571 );
xor \U$1230 ( \1573 , \1523 , \1572 );
not \U$1231 ( \1574 , \1516 );
not \U$1232 ( \1575 , \1445 );
or \U$1233 ( \1576 , \1574 , \1575 );
and \U$1234 ( \1577 , RIbb2ef80_15, \895 );
not \U$1235 ( \1578 , RIbb2ef80_15);
not \U$1236 ( \1579 , \892 );
not \U$1237 ( \1580 , \1579 );
buf \U$1238 ( \1581 , \1580 );
and \U$1239 ( \1582 , \1578 , \1581 );
nor \U$1240 ( \1583 , \1577 , \1582 );
not \U$1241 ( \1584 , \1517 );
or \U$1242 ( \1585 , \1583 , \1584 );
nand \U$1243 ( \1586 , \1576 , \1585 );
xor \U$1244 ( \1587 , \1573 , \1586 );
xor \U$1245 ( \1588 , \1522 , \1587 );
not \U$1246 ( \1589 , \1011 );
not \U$1247 ( \1590 , \1076 );
or \U$1248 ( \1591 , \1589 , \1590 );
and \U$1249 ( \1592 , \1043 , \953 );
not \U$1250 ( \1593 , \1043 );
not \U$1251 ( \1594 , \953 );
and \U$1252 ( \1595 , \1593 , \1594 );
nor \U$1253 ( \1596 , \1592 , \1595 );
nand \U$1254 ( \1597 , \1596 , \1077 );
nand \U$1255 ( \1598 , \1591 , \1597 );
not \U$1256 ( \1599 , \1430 );
not \U$1257 ( \1600 , \1388 );
or \U$1258 ( \1601 , \1599 , \1600 );
xor \U$1259 ( \1602 , \1313 , \1248 );
nand \U$1260 ( \1603 , \1602 , \1376 );
nand \U$1261 ( \1604 , \1601 , \1603 );
xor \U$1262 ( \1605 , \1598 , \1604 );
or \U$1263 ( \1606 , \1293 , \1266 );
and \U$1264 ( \1607 , \1113 , \1290 );
and \U$1265 ( \1608 , \1114 , \1245 );
nor \U$1266 ( \1609 , \1607 , \1608 );
or \U$1267 ( \1610 , \1609 , \1295 );
nand \U$1268 ( \1611 , \1606 , \1610 );
xor \U$1269 ( \1612 , \1605 , \1611 );
and \U$1270 ( \1613 , \1588 , \1612 );
and \U$1271 ( \1614 , \1522 , \1587 );
or \U$1272 ( \1615 , \1613 , \1614 );
xor \U$1273 ( \1616 , \1303 , \1615 );
xor \U$1274 ( \1617 , \1523 , \1572 );
and \U$1275 ( \1618 , \1617 , \1586 );
and \U$1276 ( \1619 , \1523 , \1572 );
or \U$1277 ( \1620 , \1618 , \1619 );
not \U$1278 ( \1621 , \1090 );
or \U$1279 ( \1622 , \1621 , \1144 );
and \U$1280 ( \1623 , \410 , \1128 );
and \U$1281 ( \1624 , \396 , \1623 );
not \U$1282 ( \1625 , \1624 );
not \U$1283 ( \1626 , \665 );
or \U$1284 ( \1627 , \1625 , \1626 );
and \U$1285 ( \1628 , \1623 , \739 );
not \U$1286 ( \1629 , \1128 );
not \U$1287 ( \1630 , \759 );
or \U$1288 ( \1631 , \1629 , \1630 );
nand \U$1289 ( \1632 , \1631 , \762 );
nor \U$1290 ( \1633 , \1628 , \1632 );
nand \U$1291 ( \1634 , \1627 , \1633 );
nand \U$1292 ( \1635 , \765 , \768 );
not \U$1293 ( \1636 , \1635 );
and \U$1294 ( \1637 , \1634 , \1636 );
not \U$1295 ( \1638 , \1634 );
and \U$1296 ( \1639 , \1638 , \1635 );
nor \U$1297 ( \1640 , \1637 , \1639 );
not \U$1298 ( \1641 , \1640 );
not \U$1299 ( \1642 , \1641 );
buf \U$1300 ( \1643 , \1642 );
not \U$1301 ( \1644 , \1643 );
and \U$1302 ( \1645 , \1644 , RIbb2f430_5);
not \U$1303 ( \1646 , \1644 );
not \U$1304 ( \1647 , RIbb2f430_5);
and \U$1305 ( \1648 , \1646 , \1647 );
nor \U$1306 ( \1649 , \1645 , \1648 );
not \U$1307 ( \1650 , \1147 );
or \U$1308 ( \1651 , \1649 , \1650 );
nand \U$1309 ( \1652 , \1622 , \1651 );
not \U$1310 ( \1653 , \996 );
not \U$1311 ( \1654 , \916 );
or \U$1312 ( \1655 , \1653 , \1654 );
not \U$1313 ( \1656 , RIbb2f070_13);
and \U$1314 ( \1657 , \1656 , \1477 );
not \U$1315 ( \1658 , \1656 );
not \U$1316 ( \1659 , \1477 );
and \U$1317 ( \1660 , \1658 , \1659 );
nor \U$1318 ( \1661 , \1657 , \1660 );
not \U$1319 ( \1662 , \998 );
or \U$1320 ( \1663 , \1661 , \1662 );
nand \U$1321 ( \1664 , \1655 , \1663 );
xor \U$1322 ( \1665 , \1652 , \1664 );
and \U$1323 ( \1666 , \410 , \400 );
and \U$1324 ( \1667 , \396 , \1666 );
not \U$1325 ( \1668 , \1667 );
not \U$1326 ( \1669 , \866 );
or \U$1327 ( \1670 , \1668 , \1669 );
and \U$1328 ( \1671 , \739 , \1666 );
not \U$1329 ( \1672 , \400 );
not \U$1330 ( \1673 , \759 );
or \U$1331 ( \1674 , \1672 , \1673 );
not \U$1332 ( \1675 , \769 );
nand \U$1333 ( \1676 , \1674 , \1675 );
nor \U$1334 ( \1677 , \1671 , \1676 );
nand \U$1335 ( \1678 , \1670 , \1677 );
not \U$1336 ( \1679 , \401 );
nand \U$1337 ( \1680 , \1679 , \771 );
not \U$1338 ( \1681 , \1680 );
and \U$1339 ( \1682 , \1678 , \1681 );
not \U$1340 ( \1683 , \1678 );
and \U$1341 ( \1684 , \1683 , \1680 );
nor \U$1342 ( \1685 , \1682 , \1684 );
not \U$1343 ( \1686 , \1685 );
not \U$1344 ( \1687 , \1686 );
not \U$1345 ( \1688 , \1687 );
buf \U$1346 ( \1689 , \1688 );
and \U$1347 ( \1690 , \1689 , RIbb2f340_7);
not \U$1348 ( \1691 , \1689 );
not \U$1349 ( \1692 , RIbb2f340_7);
and \U$1350 ( \1693 , \1691 , \1692 );
nor \U$1351 ( \1694 , \1690 , \1693 );
xor \U$1352 ( \1695 , RIbb2f340_7, RIbb2f2c8_8);
not \U$1353 ( \1696 , \1695 );
and \U$1354 ( \1697 , RIbb2f2c8_8, RIbb2f250_9);
not \U$1355 ( \1698 , RIbb2f2c8_8);
and \U$1356 ( \1699 , \1698 , \1566 );
nor \U$1357 ( \1700 , \1697 , \1699 );
nor \U$1358 ( \1701 , \1696 , \1700 );
buf \U$1359 ( \1702 , \1701 );
not \U$1360 ( \1703 , \1702 );
or \U$1361 ( \1704 , \1694 , \1703 );
not \U$1362 ( \1705 , \400 );
nor \U$1363 ( \1706 , \1705 , \401 );
and \U$1364 ( \1707 , \1706 , \410 );
and \U$1365 ( \1708 , \396 , \1707 );
not \U$1366 ( \1709 , \1708 );
not \U$1367 ( \1710 , \866 );
or \U$1368 ( \1711 , \1709 , \1710 );
and \U$1369 ( \1712 , \739 , \1707 );
not \U$1370 ( \1713 , \1706 );
not \U$1371 ( \1714 , \759 );
or \U$1372 ( \1715 , \1713 , \1714 );
and \U$1373 ( \1716 , \769 , \1679 );
not \U$1374 ( \1717 , \771 );
nor \U$1375 ( \1718 , \1716 , \1717 );
nand \U$1376 ( \1719 , \1715 , \1718 );
nor \U$1377 ( \1720 , \1712 , \1719 );
nand \U$1378 ( \1721 , \1711 , \1720 );
not \U$1379 ( \1722 , \773 );
nor \U$1380 ( \1723 , \1722 , \402 );
and \U$1381 ( \1724 , \1721 , \1723 );
not \U$1382 ( \1725 , \1721 );
not \U$1383 ( \1726 , \1723 );
and \U$1384 ( \1727 , \1725 , \1726 );
nor \U$1385 ( \1728 , \1724 , \1727 );
not \U$1386 ( \1729 , \1728 );
not \U$1387 ( \1730 , \1729 );
not \U$1388 ( \1731 , \1730 );
and \U$1389 ( \1732 , \1731 , RIbb2f340_7);
not \U$1390 ( \1733 , \1731 );
not \U$1391 ( \1734 , RIbb2f340_7);
and \U$1392 ( \1735 , \1733 , \1734 );
nor \U$1393 ( \1736 , \1732 , \1735 );
buf \U$1394 ( \1737 , \1700 );
not \U$1395 ( \1738 , \1737 );
or \U$1396 ( \1739 , \1736 , \1738 );
nand \U$1397 ( \1740 , \1704 , \1739 );
and \U$1398 ( \1741 , \1665 , \1740 );
and \U$1399 ( \1742 , \1652 , \1664 );
or \U$1400 ( \1743 , \1741 , \1742 );
xor \U$1401 ( \1744 , \1620 , \1743 );
and \U$1402 ( \1745 , \1313 , \1387 );
or \U$1403 ( \1746 , \1661 , \1654 );
and \U$1404 ( \1747 , \1514 , RIbb2f070_13);
and \U$1405 ( \1748 , \1511 , \1656 );
nor \U$1406 ( \1749 , \1747 , \1748 );
or \U$1407 ( \1750 , \1749 , \1662 );
nand \U$1408 ( \1751 , \1746 , \1750 );
xor \U$1409 ( \1752 , \1745 , \1751 );
or \U$1410 ( \1753 , \1736 , \1703 );
and \U$1411 ( \1754 , \1551 , \1734 );
not \U$1412 ( \1755 , \1551 );
and \U$1413 ( \1756 , \1755 , RIbb2f340_7);
nor \U$1414 ( \1757 , \1754 , \1756 );
or \U$1415 ( \1758 , \1757 , \1738 );
nand \U$1416 ( \1759 , \1753 , \1758 );
xor \U$1417 ( \1760 , \1752 , \1759 );
xor \U$1418 ( \1761 , \1744 , \1760 );
xor \U$1419 ( \1762 , \1616 , \1761 );
not \U$1420 ( \1763 , \1570 );
not \U$1421 ( \1764 , \1556 );
or \U$1422 ( \1765 , \1763 , \1764 );
not \U$1423 ( \1766 , \1730 );
not \U$1424 ( \1767 , \1524 );
and \U$1425 ( \1768 , \1766 , \1767 );
and \U$1426 ( \1769 , \1733 , \1554 );
nor \U$1427 ( \1770 , \1768 , \1769 );
not \U$1428 ( \1771 , \1533 );
or \U$1429 ( \1772 , \1770 , \1771 );
nand \U$1430 ( \1773 , \1765 , \1772 );
and \U$1431 ( \1774 , \814 , RIbb2eda0_19);
not \U$1432 ( \1775 , \814 );
not \U$1433 ( \1776 , RIbb2eda0_19);
and \U$1434 ( \1777 , \1775 , \1776 );
nor \U$1435 ( \1778 , \1774 , \1777 );
not \U$1436 ( \1779 , \853 );
or \U$1437 ( \1780 , \1778 , \1779 );
not \U$1438 ( \1781 , \855 );
or \U$1439 ( \1782 , \1781 , \1776 );
nand \U$1440 ( \1783 , \1780 , \1782 );
xor \U$1441 ( \1784 , \1773 , \1783 );
not \U$1442 ( \1785 , \1702 );
or \U$1443 ( \1786 , \1646 , \1692 );
or \U$1444 ( \1787 , \1644 , RIbb2f340_7);
nand \U$1445 ( \1788 , \1786 , \1787 );
not \U$1446 ( \1789 , \1788 );
or \U$1447 ( \1790 , \1785 , \1789 );
or \U$1448 ( \1791 , \1694 , \1738 );
nand \U$1449 ( \1792 , \1790 , \1791 );
and \U$1450 ( \1793 , \1784 , \1792 );
and \U$1451 ( \1794 , \1773 , \1783 );
or \U$1452 ( \1795 , \1793 , \1794 );
xor \U$1453 ( \1796 , \1652 , \1664 );
xor \U$1454 ( \1797 , \1796 , \1740 );
and \U$1455 ( \1798 , \1795 , \1797 );
not \U$1456 ( \1799 , \1077 );
not \U$1457 ( \1800 , \1045 );
or \U$1458 ( \1801 , \1799 , \1800 );
not \U$1459 ( \1802 , RIbb2f160_11);
not \U$1460 ( \1803 , \1550 );
or \U$1461 ( \1804 , \1802 , \1803 );
not \U$1462 ( \1805 , RIbb2f160_11);
nand \U$1463 ( \1806 , \1551 , \1805 );
nand \U$1464 ( \1807 , \1804 , \1806 );
nand \U$1465 ( \1808 , \1807 , \1011 );
nand \U$1466 ( \1809 , \1801 , \1808 );
not \U$1467 ( \1810 , \1376 );
not \U$1468 ( \1811 , \1423 );
or \U$1469 ( \1812 , \1810 , \1811 );
xor \U$1470 ( \1813 , \1313 , \1341 );
nand \U$1471 ( \1814 , \1813 , \1430 );
nand \U$1472 ( \1815 , \1812 , \1814 );
xor \U$1473 ( \1816 , \1809 , \1815 );
not \U$1474 ( \1817 , \1265 );
and \U$1475 ( \1818 , \1246 , \1387 );
not \U$1476 ( \1819 , \1246 );
not \U$1477 ( \1820 , \1387 );
and \U$1478 ( \1821 , \1819 , \1820 );
nor \U$1479 ( \1822 , \1818 , \1821 );
not \U$1480 ( \1823 , \1822 );
or \U$1481 ( \1824 , \1817 , \1823 );
or \U$1482 ( \1825 , \1250 , \1295 );
nand \U$1483 ( \1826 , \1824 , \1825 );
and \U$1484 ( \1827 , \1816 , \1826 );
and \U$1485 ( \1828 , \1809 , \1815 );
or \U$1486 ( \1829 , \1827 , \1828 );
not \U$1487 ( \1830 , \365 );
nand \U$1488 ( \1831 , \394 , \1830 );
nor \U$1489 ( \1832 , \1831 , \1316 );
not \U$1490 ( \1833 , \1832 );
not \U$1491 ( \1834 , \665 );
or \U$1492 ( \1835 , \1833 , \1834 );
not \U$1493 ( \1836 , \1831 );
and \U$1494 ( \1837 , \1156 , \1836 );
not \U$1495 ( \1838 , \1830 );
not \U$1496 ( \1839 , \718 );
or \U$1497 ( \1840 , \1838 , \1839 );
nand \U$1498 ( \1841 , RIbb2cf28_84, RIbb31ed8_148);
nand \U$1499 ( \1842 , \1840 , \1841 );
nor \U$1500 ( \1843 , \1837 , \1842 );
nand \U$1501 ( \1844 , \1835 , \1843 );
nand \U$1502 ( \1845 , \723 , \726 );
not \U$1503 ( \1846 , \1845 );
and \U$1504 ( \1847 , \1844 , \1846 );
not \U$1505 ( \1848 , \1844 );
and \U$1506 ( \1849 , \1848 , \1845 );
nor \U$1507 ( \1850 , \1847 , \1849 );
buf \U$1508 ( \1851 , \1850 );
buf \U$1509 ( \1852 , \1851 );
not \U$1510 ( \1853 , \1852 );
buf \U$1511 ( \1854 , \1853 );
not \U$1512 ( \1855 , \1854 );
and \U$1513 ( \1856 , \1394 , \1855 );
not \U$1514 ( \1857 , \1570 );
not \U$1515 ( \1858 , \1770 );
not \U$1516 ( \1859 , \1858 );
or \U$1517 ( \1860 , \1857 , \1859 );
not \U$1518 ( \1861 , RIbb2f250_9);
not \U$1519 ( \1862 , \1689 );
or \U$1520 ( \1863 , \1861 , \1862 );
nand \U$1521 ( \1864 , \1691 , \1524 );
nand \U$1522 ( \1865 , \1863 , \1864 );
nand \U$1523 ( \1866 , \1865 , \1533 );
nand \U$1524 ( \1867 , \1860 , \1866 );
xor \U$1525 ( \1868 , \1856 , \1867 );
not \U$1526 ( \1869 , \1517 );
not \U$1527 ( \1870 , \1478 );
or \U$1528 ( \1871 , \1869 , \1870 );
and \U$1529 ( \1872 , RIbb2ef80_15, \994 );
not \U$1530 ( \1873 , RIbb2ef80_15);
and \U$1531 ( \1874 , \1873 , \989 );
nor \U$1532 ( \1875 , \1872 , \1874 );
nand \U$1533 ( \1876 , \1875 , \1445 );
nand \U$1534 ( \1877 , \1871 , \1876 );
and \U$1535 ( \1878 , \1868 , \1877 );
and \U$1536 ( \1879 , \1856 , \1867 );
or \U$1537 ( \1880 , \1878 , \1879 );
xor \U$1538 ( \1881 , \1829 , \1880 );
not \U$1539 ( \1882 , \998 );
not \U$1540 ( \1883 , \959 );
or \U$1541 ( \1884 , \1882 , \1883 );
and \U$1542 ( \1885 , \1072 , RIbb2f070_13);
buf \U$1543 ( \1886 , \1068 );
not \U$1544 ( \1887 , \1886 );
not \U$1545 ( \1888 , \1887 );
and \U$1546 ( \1889 , \1888 , \906 );
nor \U$1547 ( \1890 , \1885 , \1889 );
or \U$1548 ( \1891 , \1890 , \1654 );
nand \U$1549 ( \1892 , \1884 , \1891 );
not \U$1550 ( \1893 , \1147 );
not \U$1551 ( \1894 , \1118 );
or \U$1552 ( \1895 , \1893 , \1894 );
and \U$1553 ( \1896 , \1285 , RIbb2f430_5);
not \U$1554 ( \1897 , \1285 );
not \U$1555 ( \1898 , RIbb2f430_5);
and \U$1556 ( \1899 , \1897 , \1898 );
nor \U$1557 ( \1900 , \1896 , \1899 );
nand \U$1558 ( \1901 , \1900 , \1090 );
nand \U$1559 ( \1902 , \1895 , \1901 );
xor \U$1560 ( \1903 , \1892 , \1902 );
not \U$1561 ( \1904 , \836 );
not \U$1562 ( \1905 , \900 );
or \U$1563 ( \1906 , \1904 , \1905 );
and \U$1564 ( \1907 , \1511 , RIbb2ee90_17);
not \U$1565 ( \1908 , \1511 );
and \U$1566 ( \1909 , \1908 , \816 );
nor \U$1567 ( \1910 , \1907 , \1909 );
not \U$1568 ( \1911 , \1910 );
or \U$1569 ( \1912 , \1911 , \833 );
nand \U$1570 ( \1913 , \1906 , \1912 );
and \U$1571 ( \1914 , \1903 , \1913 );
and \U$1572 ( \1915 , \1892 , \1902 );
or \U$1573 ( \1916 , \1914 , \1915 );
and \U$1574 ( \1917 , \1881 , \1916 );
and \U$1575 ( \1918 , \1829 , \1880 );
or \U$1576 ( \1919 , \1917 , \1918 );
xor \U$1577 ( \1920 , \1652 , \1664 );
xor \U$1578 ( \1921 , \1920 , \1740 );
and \U$1579 ( \1922 , \1919 , \1921 );
and \U$1580 ( \1923 , \1795 , \1919 );
or \U$1581 ( \1924 , \1798 , \1922 , \1923 );
or \U$1582 ( \1925 , \1583 , \1575 );
and \U$1583 ( \1926 , RIbb2ef80_15, \814 );
not \U$1584 ( \1927 , RIbb2ef80_15);
and \U$1585 ( \1928 , \1927 , \1775 );
nor \U$1586 ( \1929 , \1926 , \1928 );
or \U$1587 ( \1930 , \1929 , \1584 );
nand \U$1588 ( \1931 , \1925 , \1930 );
or \U$1589 ( \1932 , \832 , \836 );
nand \U$1590 ( \1933 , \1932 , RIbb2ee90_17);
xor \U$1591 ( \1934 , \1931 , \1933 );
not \U$1592 ( \1935 , \1011 );
not \U$1593 ( \1936 , \1596 );
or \U$1594 ( \1937 , \1935 , \1936 );
and \U$1595 ( \1938 , \993 , RIbb2f160_11);
not \U$1596 ( \1939 , \989 );
buf \U$1597 ( \1940 , \1939 );
and \U$1598 ( \1941 , \1940 , \1805 );
nor \U$1599 ( \1942 , \1938 , \1941 );
not \U$1600 ( \1943 , \1077 );
or \U$1601 ( \1944 , \1942 , \1943 );
nand \U$1602 ( \1945 , \1937 , \1944 );
xor \U$1603 ( \1946 , \1934 , \1945 );
not \U$1604 ( \1947 , \1602 );
not \U$1605 ( \1948 , \1430 );
or \U$1606 ( \1949 , \1947 , \1948 );
and \U$1607 ( \1950 , \1286 , \1394 );
not \U$1608 ( \1951 , \1313 );
and \U$1609 ( \1952 , \1285 , \1951 );
nor \U$1610 ( \1953 , \1950 , \1952 );
not \U$1611 ( \1954 , \1376 );
or \U$1612 ( \1955 , \1953 , \1954 );
nand \U$1613 ( \1956 , \1949 , \1955 );
not \U$1614 ( \1957 , \1570 );
and \U$1615 ( \1958 , RIbb2f250_9, \1888 );
not \U$1616 ( \1959 , RIbb2f250_9);
and \U$1617 ( \1960 , \1959 , \1887 );
nor \U$1618 ( \1961 , \1958 , \1960 );
not \U$1619 ( \1962 , \1961 );
or \U$1620 ( \1963 , \1957 , \1962 );
not \U$1621 ( \1964 , \1568 );
or \U$1622 ( \1965 , \1964 , \1771 );
nand \U$1623 ( \1966 , \1963 , \1965 );
xor \U$1624 ( \1967 , \1956 , \1966 );
not \U$1625 ( \1968 , \1294 );
and \U$1626 ( \1969 , \1139 , \1246 );
not \U$1627 ( \1970 , \1139 );
and \U$1628 ( \1971 , \1970 , \1289 );
nor \U$1629 ( \1972 , \1969 , \1971 );
not \U$1630 ( \1973 , \1972 );
or \U$1631 ( \1974 , \1968 , \1973 );
or \U$1632 ( \1975 , \1609 , \1266 );
nand \U$1633 ( \1976 , \1974 , \1975 );
xor \U$1634 ( \1977 , \1967 , \1976 );
xor \U$1635 ( \1978 , \1946 , \1977 );
not \U$1636 ( \1979 , \1147 );
not \U$1637 ( \1980 , RIbb2f430_5);
and \U$1638 ( \1981 , \1689 , \1980 );
not \U$1639 ( \1982 , \1689 );
and \U$1640 ( \1983 , \1982 , RIbb2f430_5);
nor \U$1641 ( \1984 , \1981 , \1983 );
not \U$1642 ( \1985 , \1984 );
or \U$1643 ( \1986 , \1979 , \1985 );
or \U$1644 ( \1987 , \1649 , \1621 );
nand \U$1645 ( \1988 , \1986 , \1987 );
xor \U$1646 ( \1989 , \1988 , \839 );
xor \U$1647 ( \1990 , \1598 , \1604 );
and \U$1648 ( \1991 , \1990 , \1611 );
and \U$1649 ( \1992 , \1598 , \1604 );
or \U$1650 ( \1993 , \1991 , \1992 );
xor \U$1651 ( \1994 , \1989 , \1993 );
xor \U$1652 ( \1995 , \1978 , \1994 );
xor \U$1653 ( \1996 , \1924 , \1995 );
xor \U$1654 ( \1997 , \840 , \1003 );
xor \U$1655 ( \1998 , \1997 , \1300 );
xor \U$1656 ( \1999 , \857 , \904 );
xor \U$1657 ( \2000 , \1999 , \1000 );
xor \U$1658 ( \2001 , \1342 , \1432 );
xor \U$1659 ( \2002 , \2001 , \1519 );
xor \U$1660 ( \2003 , \2000 , \2002 );
xor \U$1661 ( \2004 , \1079 , \1149 );
xor \U$1662 ( \2005 , \2004 , \1297 );
and \U$1663 ( \2006 , \2003 , \2005 );
and \U$1664 ( \2007 , \2000 , \2002 );
or \U$1665 ( \2008 , \2006 , \2007 );
xor \U$1666 ( \2009 , \1998 , \2008 );
xor \U$1667 ( \2010 , \1522 , \1587 );
xor \U$1668 ( \2011 , \2010 , \1612 );
and \U$1669 ( \2012 , \2009 , \2011 );
and \U$1670 ( \2013 , \1998 , \2008 );
or \U$1671 ( \2014 , \2012 , \2013 );
xor \U$1672 ( \2015 , \1996 , \2014 );
xor \U$1673 ( \2016 , \1762 , \2015 );
xor \U$1674 ( \2017 , \1652 , \1664 );
xor \U$1675 ( \2018 , \2017 , \1740 );
xor \U$1676 ( \2019 , \1795 , \1919 );
xor \U$1677 ( \2020 , \2018 , \2019 );
xor \U$1678 ( \2021 , \1773 , \1783 );
xor \U$1679 ( \2022 , \2021 , \1792 );
not \U$1680 ( \2023 , \1737 );
not \U$1681 ( \2024 , \1788 );
or \U$1682 ( \2025 , \2023 , \2024 );
and \U$1683 ( \2026 , \1140 , RIbb2f340_7);
and \U$1684 ( \2027 , \1139 , \1734 );
nor \U$1685 ( \2028 , \2026 , \2027 );
or \U$1686 ( \2029 , \2028 , \1703 );
nand \U$1687 ( \2030 , \2025 , \2029 );
not \U$1688 ( \2031 , \1783 );
xor \U$1689 ( \2032 , \2030 , \2031 );
not \U$1690 ( \2033 , \1430 );
xor \U$1691 ( \2034 , \1394 , \1855 );
not \U$1692 ( \2035 , \2034 );
or \U$1693 ( \2036 , \2033 , \2035 );
nand \U$1694 ( \2037 , \1813 , \1376 );
nand \U$1695 ( \2038 , \2036 , \2037 );
not \U$1696 ( \2039 , \832 );
and \U$1697 ( \2040 , RIbb2ee90_17, \1477 );
not \U$1698 ( \2041 , RIbb2ee90_17);
and \U$1699 ( \2042 , \2041 , \1659 );
nor \U$1700 ( \2043 , \2040 , \2042 );
not \U$1701 ( \2044 , \2043 );
or \U$1702 ( \2045 , \2039 , \2044 );
nand \U$1703 ( \2046 , \1910 , \836 );
nand \U$1704 ( \2047 , \2045 , \2046 );
xor \U$1705 ( \2048 , \2038 , \2047 );
not \U$1706 ( \2049 , \1294 );
not \U$1707 ( \2050 , \1822 );
or \U$1708 ( \2051 , \2049 , \2050 );
not \U$1709 ( \2052 , \1422 );
and \U$1710 ( \2053 , \2052 , \1290 );
and \U$1711 ( \2054 , \1422 , \1291 );
nor \U$1712 ( \2055 , \2053 , \2054 );
or \U$1713 ( \2056 , \2055 , \1266 );
nand \U$1714 ( \2057 , \2051 , \2056 );
and \U$1715 ( \2058 , \2048 , \2057 );
and \U$1716 ( \2059 , \2038 , \2047 );
or \U$1717 ( \2060 , \2058 , \2059 );
and \U$1718 ( \2061 , \2032 , \2060 );
and \U$1719 ( \2062 , \2030 , \2031 );
or \U$1720 ( \2063 , \2061 , \2062 );
xor \U$1721 ( \2064 , \2022 , \2063 );
and \U$1722 ( \2065 , RIbb2ec38_22, RIbb2ecb0_21);
not \U$1723 ( \2066 , RIbb2ec38_22);
not \U$1724 ( \2067 , RIbb2ecb0_21);
and \U$1725 ( \2068 , \2066 , \2067 );
nor \U$1726 ( \2069 , \2065 , \2068 );
not \U$1727 ( \2070 , \2069 );
and \U$1728 ( \2071 , RIbb2ec38_22, RIbb2ebc0_23);
not \U$1729 ( \2072 , RIbb2ec38_22);
not \U$1730 ( \2073 , RIbb2ebc0_23);
and \U$1731 ( \2074 , \2072 , \2073 );
nor \U$1732 ( \2075 , \2071 , \2074 );
nor \U$1733 ( \2076 , \2070 , \2075 );
buf \U$1734 ( \2077 , \2076 );
buf \U$1735 ( \2078 , \2075 );
or \U$1736 ( \2079 , \2077 , \2078 );
nand \U$1737 ( \2080 , \2079 , RIbb2ecb0_21);
not \U$1738 ( \2081 , \1581 );
and \U$1739 ( \2082 , \2081 , RIbb2eda0_19);
and \U$1740 ( \2083 , \1581 , \1776 );
nor \U$1741 ( \2084 , \2082 , \2083 );
or \U$1742 ( \2085 , \2084 , \1779 );
or \U$1743 ( \2086 , \1778 , \1781 );
nand \U$1744 ( \2087 , \2085 , \2086 );
xor \U$1745 ( \2088 , \2080 , \2087 );
and \U$1746 ( \2089 , RIbb2ef80_15, \953 );
not \U$1747 ( \2090 , RIbb2ef80_15);
and \U$1748 ( \2091 , \2090 , \1594 );
nor \U$1749 ( \2092 , \2089 , \2091 );
or \U$1750 ( \2093 , \2092 , \1575 );
not \U$1751 ( \2094 , \1875 );
or \U$1752 ( \2095 , \2094 , \1584 );
nand \U$1753 ( \2096 , \2093 , \2095 );
and \U$1754 ( \2097 , \2088 , \2096 );
and \U$1755 ( \2098 , \2080 , \2087 );
or \U$1756 ( \2099 , \2097 , \2098 );
and \U$1757 ( \2100 , \1315 , \394 );
not \U$1758 ( \2101 , \2100 );
not \U$1759 ( \2102 , \665 );
or \U$1760 ( \2103 , \2101 , \2102 );
nand \U$1761 ( \2104 , \1156 , \394 );
not \U$1762 ( \2105 , \2104 );
nor \U$1763 ( \2106 , \2105 , \718 );
nand \U$1764 ( \2107 , \2103 , \2106 );
nand \U$1765 ( \2108 , \1830 , \1841 );
not \U$1766 ( \2109 , \2108 );
and \U$1767 ( \2110 , \2107 , \2109 );
not \U$1768 ( \2111 , \2107 );
and \U$1769 ( \2112 , \2111 , \2108 );
nor \U$1770 ( \2113 , \2110 , \2112 );
buf \U$1771 ( \2114 , \2113 );
not \U$1772 ( \2115 , \2114 );
buf \U$1773 ( \2116 , \2115 );
not \U$1774 ( \2117 , \2116 );
and \U$1775 ( \2118 , \1394 , \2117 );
and \U$1776 ( \2119 , \1731 , RIbb2f160_11);
and \U$1777 ( \2120 , \1733 , \1043 );
nor \U$1778 ( \2121 , \2119 , \2120 );
not \U$1779 ( \2122 , \1011 );
or \U$1780 ( \2123 , \2121 , \2122 );
not \U$1781 ( \2124 , \1807 );
or \U$1782 ( \2125 , \2124 , \1943 );
nand \U$1783 ( \2126 , \2123 , \2125 );
xor \U$1784 ( \2127 , \2118 , \2126 );
and \U$1785 ( \2128 , \1644 , RIbb2f250_9);
and \U$1786 ( \2129 , \1646 , \1566 );
nor \U$1787 ( \2130 , \2128 , \2129 );
or \U$1788 ( \2131 , \2130 , \1771 );
not \U$1789 ( \2132 , \1865 );
not \U$1790 ( \2133 , \1570 );
or \U$1791 ( \2134 , \2132 , \2133 );
nand \U$1792 ( \2135 , \2131 , \2134 );
and \U$1793 ( \2136 , \2127 , \2135 );
and \U$1794 ( \2137 , \2118 , \2126 );
or \U$1795 ( \2138 , \2136 , \2137 );
xor \U$1796 ( \2139 , \2099 , \2138 );
and \U$1797 ( \2140 , \1113 , RIbb2f340_7);
and \U$1798 ( \2141 , \1114 , \1734 );
nor \U$1799 ( \2142 , \2140 , \2141 );
or \U$1800 ( \2143 , \2142 , \1703 );
or \U$1801 ( \2144 , \2028 , \1738 );
nand \U$1802 ( \2145 , \2143 , \2144 );
not \U$1803 ( \2146 , \1563 );
and \U$1804 ( \2147 , \2146 , RIbb2f070_13);
and \U$1805 ( \2148 , \1563 , \906 );
nor \U$1806 ( \2149 , \2147 , \2148 );
or \U$1807 ( \2150 , \2149 , \1654 );
or \U$1808 ( \2151 , \1890 , \1662 );
nand \U$1809 ( \2152 , \2150 , \2151 );
xor \U$1810 ( \2153 , \2145 , \2152 );
and \U$1811 ( \2154 , \1171 , RIbb2f430_5);
and \U$1812 ( \2155 , \1248 , \1647 );
nor \U$1813 ( \2156 , \2154 , \2155 );
or \U$1814 ( \2157 , \2156 , \1621 );
not \U$1815 ( \2158 , \1900 );
or \U$1816 ( \2159 , \2158 , \1650 );
nand \U$1817 ( \2160 , \2157 , \2159 );
and \U$1818 ( \2161 , \2153 , \2160 );
and \U$1819 ( \2162 , \2145 , \2152 );
or \U$1820 ( \2163 , \2161 , \2162 );
and \U$1821 ( \2164 , \2139 , \2163 );
and \U$1822 ( \2165 , \2099 , \2138 );
or \U$1823 ( \2166 , \2164 , \2165 );
and \U$1824 ( \2167 , \2064 , \2166 );
and \U$1825 ( \2168 , \2022 , \2063 );
or \U$1826 ( \2169 , \2167 , \2168 );
xor \U$1827 ( \2170 , \2020 , \2169 );
xor \U$1828 ( \2171 , \1856 , \1867 );
xor \U$1829 ( \2172 , \2171 , \1877 );
xor \U$1830 ( \2173 , \1809 , \1815 );
xor \U$1831 ( \2174 , \2173 , \1826 );
xor \U$1832 ( \2175 , \2172 , \2174 );
xor \U$1833 ( \2176 , \1892 , \1902 );
xor \U$1834 ( \2177 , \2176 , \1913 );
and \U$1835 ( \2178 , \2175 , \2177 );
and \U$1836 ( \2179 , \2172 , \2174 );
or \U$1837 ( \2180 , \2178 , \2179 );
xor \U$1838 ( \2181 , \1829 , \1880 );
xor \U$1839 ( \2182 , \2181 , \1916 );
xor \U$1840 ( \2183 , \2180 , \2182 );
xor \U$1841 ( \2184 , \2000 , \2002 );
xor \U$1842 ( \2185 , \2184 , \2005 );
and \U$1843 ( \2186 , \2183 , \2185 );
and \U$1844 ( \2187 , \2180 , \2182 );
or \U$1845 ( \2188 , \2186 , \2187 );
and \U$1846 ( \2189 , \2170 , \2188 );
and \U$1847 ( \2190 , \2020 , \2169 );
or \U$1848 ( \2191 , \2189 , \2190 );
xor \U$1849 ( \2192 , \2016 , \2191 );
xor \U$1850 ( \2193 , \1998 , \2008 );
xor \U$1851 ( \2194 , \2193 , \2011 );
xor \U$1852 ( \2195 , \2020 , \2169 );
xor \U$1853 ( \2196 , \2195 , \2188 );
xor \U$1854 ( \2197 , \2194 , \2196 );
xor \U$1855 ( \2198 , \2022 , \2063 );
xor \U$1856 ( \2199 , \2198 , \2166 );
xor \U$1857 ( \2200 , \2030 , \2031 );
xor \U$1858 ( \2201 , \2200 , \2060 );
buf \U$1859 ( \2202 , \389 );
and \U$1860 ( \2203 , \2202 , \392 );
and \U$1861 ( \2204 , \1315 , \2203 );
not \U$1862 ( \2205 , \2204 );
not \U$1863 ( \2206 , \665 );
or \U$1864 ( \2207 , \2205 , \2206 );
not \U$1865 ( \2208 , \2203 );
not \U$1866 ( \2209 , \1156 );
or \U$1867 ( \2210 , \2208 , \2209 );
and \U$1868 ( \2211 , \711 , \392 );
nor \U$1869 ( \2212 , \2211 , \714 );
nand \U$1870 ( \2213 , \2210 , \2212 );
not \U$1871 ( \2214 , \2213 );
nand \U$1872 ( \2215 , \2207 , \2214 );
nor \U$1873 ( \2216 , \705 , \716 );
and \U$1874 ( \2217 , \2215 , \2216 );
not \U$1875 ( \2218 , \2215 );
not \U$1876 ( \2219 , \2216 );
and \U$1877 ( \2220 , \2218 , \2219 );
nor \U$1878 ( \2221 , \2217 , \2220 );
buf \U$1879 ( \2222 , \2221 );
not \U$1880 ( \2223 , \2222 );
buf \U$1881 ( \2224 , \2223 );
not \U$1882 ( \2225 , \2224 );
and \U$1883 ( \2226 , \1313 , \2225 );
not \U$1884 ( \2227 , \1376 );
not \U$1885 ( \2228 , \2034 );
or \U$1886 ( \2229 , \2227 , \2228 );
xor \U$1887 ( \2230 , \1394 , \2117 );
nand \U$1888 ( \2231 , \2230 , \1430 );
nand \U$1889 ( \2232 , \2229 , \2231 );
xor \U$1890 ( \2233 , \2226 , \2232 );
not \U$1891 ( \2234 , \836 );
not \U$1892 ( \2235 , \2043 );
or \U$1893 ( \2236 , \2234 , \2235 );
not \U$1894 ( \2237 , RIbb2ee90_17);
not \U$1895 ( \2238 , \989 );
or \U$1896 ( \2239 , \2237 , \2238 );
not \U$1897 ( \2240 , RIbb2ee90_17);
nand \U$1898 ( \2241 , \1940 , \2240 );
nand \U$1899 ( \2242 , \2239 , \2241 );
not \U$1900 ( \2243 , \2242 );
or \U$1901 ( \2244 , \2243 , \833 );
nand \U$1902 ( \2245 , \2236 , \2244 );
and \U$1903 ( \2246 , \2233 , \2245 );
and \U$1904 ( \2247 , \2226 , \2232 );
or \U$1905 ( \2248 , \2246 , \2247 );
not \U$1906 ( \2249 , RIbb2ecb0_21);
not \U$1907 ( \2250 , \2249 );
buf \U$1908 ( \2251 , \811 );
not \U$1909 ( \2252 , \2251 );
or \U$1910 ( \2253 , \2250 , \2252 );
not \U$1911 ( \2254 , RIbb2ecb0_21);
or \U$1912 ( \2255 , \1775 , \2254 );
nand \U$1913 ( \2256 , \2253 , \2255 );
and \U$1914 ( \2257 , \2256 , \2077 );
and \U$1915 ( \2258 , \2078 , RIbb2ecb0_21);
nor \U$1916 ( \2259 , \2257 , \2258 );
not \U$1917 ( \2260 , \2259 );
xor \U$1918 ( \2261 , \2248 , \2260 );
and \U$1919 ( \2262 , RIbb2ef80_15, \1072 );
not \U$1920 ( \2263 , RIbb2ef80_15);
and \U$1921 ( \2264 , \2263 , \1888 );
nor \U$1922 ( \2265 , \2262 , \2264 );
or \U$1923 ( \2266 , \2265 , \1575 );
or \U$1924 ( \2267 , \2092 , \1584 );
nand \U$1925 ( \2268 , \2266 , \2267 );
not \U$1926 ( \2269 , \853 );
and \U$1927 ( \2270 , \1511 , RIbb2eda0_19);
not \U$1928 ( \2271 , \1511 );
and \U$1929 ( \2272 , \2271 , \843 );
nor \U$1930 ( \2273 , \2270 , \2272 );
not \U$1931 ( \2274 , \2273 );
or \U$1932 ( \2275 , \2269 , \2274 );
or \U$1933 ( \2276 , \2084 , \1781 );
nand \U$1934 ( \2277 , \2275 , \2276 );
xor \U$1935 ( \2278 , \2268 , \2277 );
not \U$1936 ( \2279 , \1702 );
and \U$1937 ( \2280 , \1285 , RIbb2f340_7);
not \U$1938 ( \2281 , \1285 );
and \U$1939 ( \2282 , \2281 , \1734 );
nor \U$1940 ( \2283 , \2280 , \2282 );
not \U$1941 ( \2284 , \2283 );
or \U$1942 ( \2285 , \2279 , \2284 );
or \U$1943 ( \2286 , \2142 , \1738 );
nand \U$1944 ( \2287 , \2285 , \2286 );
and \U$1945 ( \2288 , \2278 , \2287 );
and \U$1946 ( \2289 , \2268 , \2277 );
or \U$1947 ( \2290 , \2288 , \2289 );
and \U$1948 ( \2291 , \2261 , \2290 );
and \U$1949 ( \2292 , \2248 , \2260 );
or \U$1950 ( \2293 , \2291 , \2292 );
xor \U$1951 ( \2294 , \2201 , \2293 );
xor \U$1952 ( \2295 , \2080 , \2087 );
xor \U$1953 ( \2296 , \2295 , \2096 );
xor \U$1954 ( \2297 , \2145 , \2152 );
xor \U$1955 ( \2298 , \2297 , \2160 );
xor \U$1956 ( \2299 , \2296 , \2298 );
xor \U$1957 ( \2300 , \2038 , \2047 );
xor \U$1958 ( \2301 , \2300 , \2057 );
and \U$1959 ( \2302 , \2299 , \2301 );
and \U$1960 ( \2303 , \2296 , \2298 );
or \U$1961 ( \2304 , \2302 , \2303 );
and \U$1962 ( \2305 , \2294 , \2304 );
and \U$1963 ( \2306 , \2201 , \2293 );
or \U$1964 ( \2307 , \2305 , \2306 );
xor \U$1965 ( \2308 , \2199 , \2307 );
xor \U$1966 ( \2309 , \2180 , \2182 );
xor \U$1967 ( \2310 , \2309 , \2185 );
and \U$1968 ( \2311 , \2308 , \2310 );
and \U$1969 ( \2312 , \2199 , \2307 );
or \U$1970 ( \2313 , \2311 , \2312 );
and \U$1971 ( \2314 , \2197 , \2313 );
and \U$1972 ( \2315 , \2194 , \2196 );
or \U$1973 ( \2316 , \2314 , \2315 );
nor \U$1974 ( \2317 , \2192 , \2316 );
xor \U$1975 ( \2318 , \1988 , \839 );
and \U$1976 ( \2319 , \2318 , \1993 );
and \U$1977 ( \2320 , \1988 , \839 );
or \U$1978 ( \2321 , \2319 , \2320 );
xor \U$1979 ( \2322 , \1620 , \1743 );
and \U$1980 ( \2323 , \2322 , \1760 );
and \U$1981 ( \2324 , \1620 , \1743 );
or \U$1982 ( \2325 , \2323 , \2324 );
xor \U$1983 ( \2326 , \2321 , \2325 );
xor \U$1984 ( \2327 , \1931 , \1933 );
and \U$1985 ( \2328 , \2327 , \1945 );
and \U$1986 ( \2329 , \1931 , \1933 );
or \U$1987 ( \2330 , \2328 , \2329 );
xor \U$1988 ( \2331 , \1745 , \1751 );
and \U$1989 ( \2332 , \2331 , \1759 );
and \U$1990 ( \2333 , \1745 , \1751 );
or \U$1991 ( \2334 , \2332 , \2333 );
xor \U$1992 ( \2335 , \2330 , \2334 );
xor \U$1993 ( \2336 , \1956 , \1966 );
and \U$1994 ( \2337 , \2336 , \1976 );
and \U$1995 ( \2338 , \1956 , \1966 );
or \U$1996 ( \2339 , \2337 , \2338 );
xor \U$1997 ( \2340 , \2335 , \2339 );
xor \U$1998 ( \2341 , \2326 , \2340 );
xor \U$1999 ( \2342 , \1924 , \1995 );
and \U$2000 ( \2343 , \2342 , \2014 );
and \U$2001 ( \2344 , \1924 , \1995 );
or \U$2002 ( \2345 , \2343 , \2344 );
xor \U$2003 ( \2346 , \2341 , \2345 );
not \U$2004 ( \2347 , \1265 );
not \U$2005 ( \2348 , \1972 );
or \U$2006 ( \2349 , \2347 , \2348 );
and \U$2007 ( \2350 , \1644 , \1290 );
and \U$2008 ( \2351 , \1646 , \1289 );
nor \U$2009 ( \2352 , \2350 , \2351 );
or \U$2010 ( \2353 , \2352 , \1295 );
nand \U$2011 ( \2354 , \2349 , \2353 );
or \U$2012 ( \2355 , \1929 , \1575 );
not \U$2013 ( \2356 , RIbb2ef80_15);
or \U$2014 ( \2357 , \1584 , \2356 );
nand \U$2015 ( \2358 , \2355 , \2357 );
not \U$2016 ( \2359 , \2358 );
xor \U$2017 ( \2360 , \2354 , \2359 );
not \U$2018 ( \2361 , \1090 );
not \U$2019 ( \2362 , \1984 );
or \U$2020 ( \2363 , \2361 , \2362 );
and \U$2021 ( \2364 , \1731 , RIbb2f430_5);
and \U$2022 ( \2365 , \1733 , \1898 );
nor \U$2023 ( \2366 , \2364 , \2365 );
or \U$2024 ( \2367 , \2366 , \1650 );
nand \U$2025 ( \2368 , \2363 , \2367 );
xor \U$2026 ( \2369 , \2360 , \2368 );
or \U$2027 ( \2370 , \1749 , \1654 );
and \U$2028 ( \2371 , RIbb2f070_13, \2081 );
not \U$2029 ( \2372 , RIbb2f070_13);
and \U$2030 ( \2373 , \2372 , \1581 );
nor \U$2031 ( \2374 , \2371 , \2373 );
or \U$2032 ( \2375 , \2374 , \1662 );
nand \U$2033 ( \2376 , \2370 , \2375 );
not \U$2034 ( \2377 , \1077 );
and \U$2035 ( \2378 , \1477 , RIbb2f160_11);
not \U$2036 ( \2379 , \1477 );
and \U$2037 ( \2380 , \2379 , \1048 );
nor \U$2038 ( \2381 , \2378 , \2380 );
not \U$2039 ( \2382 , \2381 );
or \U$2040 ( \2383 , \2377 , \2382 );
or \U$2041 ( \2384 , \1942 , \2122 );
nand \U$2042 ( \2385 , \2383 , \2384 );
xor \U$2043 ( \2386 , \2376 , \2385 );
or \U$2044 ( \2387 , \1757 , \1703 );
and \U$2045 ( \2388 , \2146 , RIbb2f340_7);
and \U$2046 ( \2389 , \1042 , \1734 );
nor \U$2047 ( \2390 , \2388 , \2389 );
or \U$2048 ( \2391 , \2390 , \1738 );
nand \U$2049 ( \2392 , \2387 , \2391 );
xor \U$2050 ( \2393 , \2386 , \2392 );
xor \U$2051 ( \2394 , \2369 , \2393 );
and \U$2052 ( \2395 , \1313 , \1248 );
not \U$2053 ( \2396 , \1533 );
not \U$2054 ( \2397 , \1961 );
or \U$2055 ( \2398 , \2396 , \2397 );
not \U$2056 ( \2399 , \957 );
and \U$2057 ( \2400 , \1554 , \2399 );
not \U$2058 ( \2401 , \1554 );
and \U$2059 ( \2402 , \2401 , \1594 );
nor \U$2060 ( \2403 , \2400 , \2402 );
nand \U$2061 ( \2404 , \2403 , \1570 );
nand \U$2062 ( \2405 , \2398 , \2404 );
xor \U$2063 ( \2406 , \2395 , \2405 );
or \U$2064 ( \2407 , \1953 , \1948 );
and \U$2065 ( \2408 , \1113 , \1394 );
not \U$2066 ( \2409 , \1394 );
and \U$2067 ( \2410 , \1114 , \2409 );
nor \U$2068 ( \2411 , \2408 , \2410 );
or \U$2069 ( \2412 , \2411 , \1954 );
nand \U$2070 ( \2413 , \2407 , \2412 );
xor \U$2071 ( \2414 , \2406 , \2413 );
xor \U$2072 ( \2415 , \2394 , \2414 );
xor \U$2073 ( \2416 , \1946 , \1977 );
and \U$2074 ( \2417 , \2416 , \1994 );
and \U$2075 ( \2418 , \1946 , \1977 );
or \U$2076 ( \2419 , \2417 , \2418 );
xor \U$2077 ( \2420 , \1303 , \1615 );
and \U$2078 ( \2421 , \2420 , \1761 );
and \U$2079 ( \2422 , \1303 , \1615 );
or \U$2080 ( \2423 , \2421 , \2422 );
xor \U$2081 ( \2424 , \2419 , \2423 );
xor \U$2082 ( \2425 , \2415 , \2424 );
xor \U$2083 ( \2426 , \2346 , \2425 );
xor \U$2084 ( \2427 , \1762 , \2015 );
and \U$2085 ( \2428 , \2427 , \2191 );
and \U$2086 ( \2429 , \1762 , \2015 );
or \U$2087 ( \2430 , \2428 , \2429 );
nor \U$2088 ( \2431 , \2426 , \2430 );
nor \U$2089 ( \2432 , \2317 , \2431 );
and \U$2090 ( \2433 , \1285 , \1394 );
or \U$2091 ( \2434 , \2390 , \1703 );
and \U$2092 ( \2435 , RIbb2f340_7, \1072 );
not \U$2093 ( \2436 , RIbb2f340_7);
and \U$2094 ( \2437 , \2436 , \1071 );
nor \U$2095 ( \2438 , \2435 , \2437 );
or \U$2096 ( \2439 , \2438 , \1738 );
nand \U$2097 ( \2440 , \2434 , \2439 );
xor \U$2098 ( \2441 , \2433 , \2440 );
or \U$2099 ( \2442 , \2411 , \1948 );
and \U$2100 ( \2443 , \1140 , \1313 );
and \U$2101 ( \2444 , \1139 , \2409 );
nor \U$2102 ( \2445 , \2443 , \2444 );
or \U$2103 ( \2446 , \2445 , \1954 );
nand \U$2104 ( \2447 , \2442 , \2446 );
xor \U$2105 ( \2448 , \2441 , \2447 );
xor \U$2106 ( \2449 , \2395 , \2405 );
and \U$2107 ( \2450 , \2449 , \2413 );
and \U$2108 ( \2451 , \2395 , \2405 );
or \U$2109 ( \2452 , \2450 , \2451 );
xor \U$2110 ( \2453 , \2358 , \2452 );
xor \U$2111 ( \2454 , \2376 , \2385 );
and \U$2112 ( \2455 , \2454 , \2392 );
and \U$2113 ( \2456 , \2376 , \2385 );
or \U$2114 ( \2457 , \2455 , \2456 );
xor \U$2115 ( \2458 , \2453 , \2457 );
and \U$2116 ( \2459 , \2448 , \2458 );
xor \U$2117 ( \2460 , \2330 , \2334 );
and \U$2118 ( \2461 , \2460 , \2339 );
and \U$2119 ( \2462 , \2330 , \2334 );
or \U$2120 ( \2463 , \2461 , \2462 );
xor \U$2121 ( \2464 , \2358 , \2452 );
xor \U$2122 ( \2465 , \2464 , \2457 );
and \U$2123 ( \2466 , \2463 , \2465 );
and \U$2124 ( \2467 , \2448 , \2463 );
or \U$2125 ( \2468 , \2459 , \2466 , \2467 );
not \U$2126 ( \2469 , \1147 );
and \U$2127 ( \2470 , \1551 , RIbb2f430_5);
not \U$2128 ( \2471 , \1551 );
and \U$2129 ( \2472 , \2471 , \1980 );
nor \U$2130 ( \2473 , \2470 , \2472 );
not \U$2131 ( \2474 , \2473 );
or \U$2132 ( \2475 , \2469 , \2474 );
or \U$2133 ( \2476 , \2366 , \1621 );
nand \U$2134 ( \2477 , \2475 , \2476 );
not \U$2135 ( \2478 , \1011 );
not \U$2136 ( \2479 , \2381 );
or \U$2137 ( \2480 , \2478 , \2479 );
and \U$2138 ( \2481 , \1514 , RIbb2f160_11);
and \U$2139 ( \2482 , \1511 , \1805 );
nor \U$2140 ( \2483 , \2481 , \2482 );
or \U$2141 ( \2484 , \2483 , \1943 );
nand \U$2142 ( \2485 , \2480 , \2484 );
xor \U$2143 ( \2486 , \2477 , \2485 );
not \U$2144 ( \2487 , \1294 );
or \U$2145 ( \2488 , \1691 , \1245 );
or \U$2146 ( \2489 , \1689 , \1290 );
nand \U$2147 ( \2490 , \2488 , \2489 );
not \U$2148 ( \2491 , \2490 );
or \U$2149 ( \2492 , \2487 , \2491 );
or \U$2150 ( \2493 , \2352 , \1266 );
nand \U$2151 ( \2494 , \2492 , \2493 );
and \U$2152 ( \2495 , \2486 , \2494 );
and \U$2153 ( \2496 , \2477 , \2485 );
or \U$2154 ( \2497 , \2495 , \2496 );
xor \U$2155 ( \2498 , \2433 , \2440 );
and \U$2156 ( \2499 , \2498 , \2447 );
and \U$2157 ( \2500 , \2433 , \2440 );
or \U$2158 ( \2501 , \2499 , \2500 );
xor \U$2159 ( \2502 , \2497 , \2501 );
and \U$2160 ( \2503 , \993 , RIbb2f250_9);
and \U$2161 ( \2504 , \1940 , \1554 );
nor \U$2162 ( \2505 , \2503 , \2504 );
or \U$2163 ( \2506 , \2505 , \1771 );
and \U$2164 ( \2507 , \1659 , RIbb2f250_9);
and \U$2165 ( \2508 , \1477 , \1566 );
nor \U$2166 ( \2509 , \2507 , \2508 );
or \U$2167 ( \2510 , \2509 , \2133 );
nand \U$2168 ( \2511 , \2506 , \2510 );
not \U$2169 ( \2512 , \2473 );
or \U$2170 ( \2513 , \2512 , \1621 );
not \U$2171 ( \2514 , RIbb2f430_5);
not \U$2172 ( \2515 , \1039 );
or \U$2173 ( \2516 , \2514 , \2515 );
nand \U$2174 ( \2517 , \1042 , \1980 );
nand \U$2175 ( \2518 , \2516 , \2517 );
not \U$2176 ( \2519 , \2518 );
or \U$2177 ( \2520 , \2519 , \1650 );
nand \U$2178 ( \2521 , \2513 , \2520 );
xor \U$2179 ( \2522 , \2511 , \2521 );
not \U$2180 ( \2523 , \1265 );
not \U$2181 ( \2524 , \2490 );
or \U$2182 ( \2525 , \2523 , \2524 );
and \U$2183 ( \2526 , \1731 , \1246 );
and \U$2184 ( \2527 , \1733 , \1291 );
nor \U$2185 ( \2528 , \2526 , \2527 );
or \U$2186 ( \2529 , \2528 , \1295 );
nand \U$2187 ( \2530 , \2525 , \2529 );
xor \U$2188 ( \2531 , \2522 , \2530 );
xor \U$2189 ( \2532 , \2502 , \2531 );
xor \U$2190 ( \2533 , \2354 , \2359 );
and \U$2191 ( \2534 , \2533 , \2368 );
and \U$2192 ( \2535 , \2354 , \2359 );
or \U$2193 ( \2536 , \2534 , \2535 );
or \U$2194 ( \2537 , \1445 , \1517 );
nand \U$2195 ( \2538 , \2537 , RIbb2ef80_15);
or \U$2196 ( \2539 , \2374 , \1654 );
and \U$2197 ( \2540 , \814 , RIbb2f070_13);
and \U$2198 ( \2541 , \815 , \906 );
nor \U$2199 ( \2542 , \2540 , \2541 );
or \U$2200 ( \2543 , \2542 , \1662 );
nand \U$2201 ( \2544 , \2539 , \2543 );
xor \U$2202 ( \2545 , \2538 , \2544 );
not \U$2203 ( \2546 , \2403 );
or \U$2204 ( \2547 , \2546 , \1771 );
or \U$2205 ( \2548 , \2505 , \2133 );
nand \U$2206 ( \2549 , \2547 , \2548 );
xor \U$2207 ( \2550 , \2545 , \2549 );
xor \U$2208 ( \2551 , \2536 , \2550 );
xor \U$2209 ( \2552 , \2477 , \2485 );
xor \U$2210 ( \2553 , \2552 , \2494 );
and \U$2211 ( \2554 , \2551 , \2553 );
and \U$2212 ( \2555 , \2536 , \2550 );
or \U$2213 ( \2556 , \2554 , \2555 );
xor \U$2214 ( \2557 , \2532 , \2556 );
not \U$2215 ( \2558 , \1394 );
nor \U$2216 ( \2559 , \2558 , \1113 );
or \U$2217 ( \2560 , \2438 , \1703 );
and \U$2218 ( \2561 , \953 , RIbb2f340_7);
and \U$2219 ( \2562 , \1594 , \1692 );
nor \U$2220 ( \2563 , \2561 , \2562 );
or \U$2221 ( \2564 , \2563 , \1738 );
nand \U$2222 ( \2565 , \2560 , \2564 );
xor \U$2223 ( \2566 , \2559 , \2565 );
not \U$2224 ( \2567 , \1077 );
and \U$2225 ( \2568 , \1581 , RIbb2f160_11);
not \U$2226 ( \2569 , \1581 );
and \U$2227 ( \2570 , \2569 , \1048 );
nor \U$2228 ( \2571 , \2568 , \2570 );
not \U$2229 ( \2572 , \2571 );
or \U$2230 ( \2573 , \2567 , \2572 );
or \U$2231 ( \2574 , \2483 , \2122 );
nand \U$2232 ( \2575 , \2573 , \2574 );
xor \U$2233 ( \2576 , \2566 , \2575 );
or \U$2234 ( \2577 , \2445 , \1948 );
and \U$2235 ( \2578 , \1644 , \1313 );
and \U$2236 ( \2579 , \1646 , \1951 );
nor \U$2237 ( \2580 , \2578 , \2579 );
or \U$2238 ( \2581 , \2580 , \1954 );
nand \U$2239 ( \2582 , \2577 , \2581 );
or \U$2240 ( \2583 , \2542 , \1654 );
or \U$2241 ( \2584 , \1662 , \1656 );
nand \U$2242 ( \2585 , \2583 , \2584 );
not \U$2243 ( \2586 , \2585 );
xor \U$2244 ( \2587 , \2582 , \2586 );
xor \U$2245 ( \2588 , \2538 , \2544 );
and \U$2246 ( \2589 , \2588 , \2549 );
and \U$2247 ( \2590 , \2538 , \2544 );
or \U$2248 ( \2591 , \2589 , \2590 );
xor \U$2249 ( \2592 , \2587 , \2591 );
xor \U$2250 ( \2593 , \2576 , \2592 );
xor \U$2251 ( \2594 , \2358 , \2452 );
and \U$2252 ( \2595 , \2594 , \2457 );
and \U$2253 ( \2596 , \2358 , \2452 );
or \U$2254 ( \2597 , \2595 , \2596 );
xor \U$2255 ( \2598 , \2593 , \2597 );
xor \U$2256 ( \2599 , \2557 , \2598 );
xor \U$2257 ( \2600 , \2468 , \2599 );
xor \U$2258 ( \2601 , \2369 , \2393 );
and \U$2259 ( \2602 , \2601 , \2414 );
and \U$2260 ( \2603 , \2369 , \2393 );
or \U$2261 ( \2604 , \2602 , \2603 );
xor \U$2262 ( \2605 , \2536 , \2550 );
xor \U$2263 ( \2606 , \2605 , \2553 );
xor \U$2264 ( \2607 , \2604 , \2606 );
xor \U$2265 ( \2608 , \2321 , \2325 );
and \U$2266 ( \2609 , \2608 , \2340 );
and \U$2267 ( \2610 , \2321 , \2325 );
or \U$2268 ( \2611 , \2609 , \2610 );
and \U$2269 ( \2612 , \2607 , \2611 );
and \U$2270 ( \2613 , \2604 , \2606 );
or \U$2271 ( \2614 , \2612 , \2613 );
xor \U$2272 ( \2615 , \2600 , \2614 );
xor \U$2273 ( \2616 , \2358 , \2452 );
xor \U$2274 ( \2617 , \2616 , \2457 );
xor \U$2275 ( \2618 , \2448 , \2463 );
xor \U$2276 ( \2619 , \2617 , \2618 );
xor \U$2277 ( \2620 , \2369 , \2393 );
xor \U$2278 ( \2621 , \2620 , \2414 );
and \U$2279 ( \2622 , \2419 , \2621 );
xor \U$2280 ( \2623 , \2369 , \2393 );
xor \U$2281 ( \2624 , \2623 , \2414 );
and \U$2282 ( \2625 , \2423 , \2624 );
and \U$2283 ( \2626 , \2419 , \2423 );
or \U$2284 ( \2627 , \2622 , \2625 , \2626 );
xor \U$2285 ( \2628 , \2619 , \2627 );
xor \U$2286 ( \2629 , \2604 , \2606 );
xor \U$2287 ( \2630 , \2629 , \2611 );
and \U$2288 ( \2631 , \2628 , \2630 );
and \U$2289 ( \2632 , \2619 , \2627 );
or \U$2290 ( \2633 , \2631 , \2632 );
or \U$2291 ( \2634 , \2615 , \2633 );
xor \U$2292 ( \2635 , \2619 , \2627 );
xor \U$2293 ( \2636 , \2635 , \2630 );
xor \U$2294 ( \2637 , \2341 , \2345 );
and \U$2295 ( \2638 , \2637 , \2425 );
and \U$2296 ( \2639 , \2341 , \2345 );
or \U$2297 ( \2640 , \2638 , \2639 );
or \U$2298 ( \2641 , \2636 , \2640 );
and \U$2299 ( \2642 , \2432 , \2634 , \2641 );
or \U$2300 ( \2643 , \2580 , \1948 );
and \U$2301 ( \2644 , \1689 , \1313 );
and \U$2302 ( \2645 , \1691 , \2409 );
nor \U$2303 ( \2646 , \2644 , \2645 );
or \U$2304 ( \2647 , \2646 , \1954 );
nand \U$2305 ( \2648 , \2643 , \2647 );
xor \U$2306 ( \2649 , \2585 , \2648 );
or \U$2307 ( \2650 , \2528 , \1266 );
and \U$2308 ( \2651 , \1550 , \1290 );
not \U$2309 ( \2652 , \1550 );
and \U$2310 ( \2653 , \2652 , \1289 );
nor \U$2311 ( \2654 , \2651 , \2653 );
or \U$2312 ( \2655 , \2654 , \1295 );
nand \U$2313 ( \2656 , \2650 , \2655 );
xor \U$2314 ( \2657 , \2649 , \2656 );
nor \U$2315 ( \2658 , \1140 , \2409 );
not \U$2316 ( \2659 , \1147 );
and \U$2317 ( \2660 , RIbb2f430_5, \1888 );
not \U$2318 ( \2661 , RIbb2f430_5);
and \U$2319 ( \2662 , \2661 , \1072 );
nor \U$2320 ( \2663 , \2660 , \2662 );
not \U$2321 ( \2664 , \2663 );
or \U$2322 ( \2665 , \2659 , \2664 );
nand \U$2323 ( \2666 , \2518 , \1090 );
nand \U$2324 ( \2667 , \2665 , \2666 );
xor \U$2325 ( \2668 , \2658 , \2667 );
or \U$2326 ( \2669 , \2509 , \1771 );
and \U$2327 ( \2670 , \1514 , RIbb2f250_9);
and \U$2328 ( \2671 , \1511 , \1566 );
nor \U$2329 ( \2672 , \2670 , \2671 );
or \U$2330 ( \2673 , \2672 , \2133 );
nand \U$2331 ( \2674 , \2669 , \2673 );
xor \U$2332 ( \2675 , \2668 , \2674 );
xor \U$2333 ( \2676 , \2582 , \2586 );
and \U$2334 ( \2677 , \2676 , \2591 );
and \U$2335 ( \2678 , \2582 , \2586 );
or \U$2336 ( \2679 , \2677 , \2678 );
xor \U$2337 ( \2680 , \2675 , \2679 );
xor \U$2338 ( \2681 , \2657 , \2680 );
xor \U$2339 ( \2682 , \2497 , \2501 );
and \U$2340 ( \2683 , \2682 , \2531 );
and \U$2341 ( \2684 , \2497 , \2501 );
or \U$2342 ( \2685 , \2683 , \2684 );
or \U$2343 ( \2686 , \916 , \998 );
nand \U$2344 ( \2687 , \2686 , RIbb2f070_13);
not \U$2345 ( \2688 , \1011 );
not \U$2346 ( \2689 , \2571 );
or \U$2347 ( \2690 , \2688 , \2689 );
and \U$2348 ( \2691 , \814 , RIbb2f160_11);
and \U$2349 ( \2692 , \815 , \1805 );
nor \U$2350 ( \2693 , \2691 , \2692 );
or \U$2351 ( \2694 , \2693 , \1943 );
nand \U$2352 ( \2695 , \2690 , \2694 );
xor \U$2353 ( \2696 , \2687 , \2695 );
not \U$2354 ( \2697 , \1737 );
and \U$2355 ( \2698 , \994 , RIbb2f340_7);
not \U$2356 ( \2699 , \994 );
not \U$2357 ( \2700 , RIbb2f340_7);
and \U$2358 ( \2701 , \2699 , \2700 );
nor \U$2359 ( \2702 , \2698 , \2701 );
not \U$2360 ( \2703 , \2702 );
or \U$2361 ( \2704 , \2697 , \2703 );
or \U$2362 ( \2705 , \2563 , \1703 );
nand \U$2363 ( \2706 , \2704 , \2705 );
xor \U$2364 ( \2707 , \2696 , \2706 );
xor \U$2365 ( \2708 , \2559 , \2565 );
and \U$2366 ( \2709 , \2708 , \2575 );
and \U$2367 ( \2710 , \2559 , \2565 );
or \U$2368 ( \2711 , \2709 , \2710 );
xor \U$2369 ( \2712 , \2511 , \2521 );
and \U$2370 ( \2713 , \2712 , \2530 );
and \U$2371 ( \2714 , \2511 , \2521 );
or \U$2372 ( \2715 , \2713 , \2714 );
xor \U$2373 ( \2716 , \2711 , \2715 );
xor \U$2374 ( \2717 , \2707 , \2716 );
xor \U$2375 ( \2718 , \2685 , \2717 );
xor \U$2376 ( \2719 , \2576 , \2592 );
and \U$2377 ( \2720 , \2719 , \2597 );
and \U$2378 ( \2721 , \2576 , \2592 );
or \U$2379 ( \2722 , \2720 , \2721 );
xor \U$2380 ( \2723 , \2718 , \2722 );
xor \U$2381 ( \2724 , \2681 , \2723 );
xor \U$2382 ( \2725 , \2532 , \2556 );
and \U$2383 ( \2726 , \2725 , \2598 );
and \U$2384 ( \2727 , \2532 , \2556 );
or \U$2385 ( \2728 , \2726 , \2727 );
xor \U$2386 ( \2729 , \2724 , \2728 );
xor \U$2387 ( \2730 , \2468 , \2599 );
and \U$2388 ( \2731 , \2730 , \2614 );
and \U$2389 ( \2732 , \2468 , \2599 );
or \U$2390 ( \2733 , \2731 , \2732 );
nor \U$2391 ( \2734 , \2729 , \2733 );
xor \U$2392 ( \2735 , \2681 , \2723 );
and \U$2393 ( \2736 , \2735 , \2728 );
and \U$2394 ( \2737 , \2681 , \2723 );
or \U$2395 ( \2738 , \2736 , \2737 );
xor \U$2396 ( \2739 , \2585 , \2648 );
xor \U$2397 ( \2740 , \2739 , \2656 );
and \U$2398 ( \2741 , \2675 , \2740 );
xor \U$2399 ( \2742 , \2585 , \2648 );
xor \U$2400 ( \2743 , \2742 , \2656 );
and \U$2401 ( \2744 , \2679 , \2743 );
and \U$2402 ( \2745 , \2675 , \2679 );
or \U$2403 ( \2746 , \2741 , \2744 , \2745 );
xor \U$2404 ( \2747 , \2658 , \2667 );
and \U$2405 ( \2748 , \2747 , \2674 );
and \U$2406 ( \2749 , \2658 , \2667 );
or \U$2407 ( \2750 , \2748 , \2749 );
or \U$2408 ( \2751 , \2693 , \2122 );
or \U$2409 ( \2752 , \1943 , \1043 );
nand \U$2410 ( \2753 , \2751 , \2752 );
not \U$2411 ( \2754 , \2753 );
xor \U$2412 ( \2755 , \2750 , \2754 );
xor \U$2413 ( \2756 , \2687 , \2695 );
and \U$2414 ( \2757 , \2756 , \2706 );
and \U$2415 ( \2758 , \2687 , \2695 );
or \U$2416 ( \2759 , \2757 , \2758 );
xor \U$2417 ( \2760 , \2755 , \2759 );
xor \U$2418 ( \2761 , \2687 , \2695 );
xor \U$2419 ( \2762 , \2761 , \2706 );
and \U$2420 ( \2763 , \2711 , \2762 );
xor \U$2421 ( \2764 , \2687 , \2695 );
xor \U$2422 ( \2765 , \2764 , \2706 );
and \U$2423 ( \2766 , \2715 , \2765 );
and \U$2424 ( \2767 , \2711 , \2715 );
or \U$2425 ( \2768 , \2763 , \2766 , \2767 );
xor \U$2426 ( \2769 , \2760 , \2768 );
not \U$2427 ( \2770 , \1090 );
not \U$2428 ( \2771 , \2663 );
or \U$2429 ( \2772 , \2770 , \2771 );
and \U$2430 ( \2773 , RIbb2f430_5, \953 );
not \U$2431 ( \2774 , RIbb2f430_5);
and \U$2432 ( \2775 , \2774 , \957 );
nor \U$2433 ( \2776 , \2773 , \2775 );
or \U$2434 ( \2777 , \2776 , \1650 );
nand \U$2435 ( \2778 , \2772 , \2777 );
or \U$2436 ( \2779 , \2654 , \1266 );
and \U$2437 ( \2780 , \1562 , \1246 );
and \U$2438 ( \2781 , \1563 , \1291 );
nor \U$2439 ( \2782 , \2780 , \2781 );
or \U$2440 ( \2783 , \2782 , \1295 );
nand \U$2441 ( \2784 , \2779 , \2783 );
xor \U$2442 ( \2785 , \2778 , \2784 );
or \U$2443 ( \2786 , \2672 , \1771 );
and \U$2444 ( \2787 , \2081 , RIbb2f250_9);
and \U$2445 ( \2788 , \1581 , \1524 );
nor \U$2446 ( \2789 , \2787 , \2788 );
or \U$2447 ( \2790 , \2789 , \2133 );
nand \U$2448 ( \2791 , \2786 , \2790 );
xor \U$2449 ( \2792 , \2785 , \2791 );
xor \U$2450 ( \2793 , \2585 , \2648 );
and \U$2451 ( \2794 , \2793 , \2656 );
and \U$2452 ( \2795 , \2585 , \2648 );
or \U$2453 ( \2796 , \2794 , \2795 );
xor \U$2454 ( \2797 , \2792 , \2796 );
and \U$2455 ( \2798 , \1646 , \1394 );
not \U$2456 ( \2799 , \1702 );
not \U$2457 ( \2800 , \2702 );
or \U$2458 ( \2801 , \2799 , \2800 );
and \U$2459 ( \2802 , \1734 , \1659 );
not \U$2460 ( \2803 , \1734 );
and \U$2461 ( \2804 , \2803 , \1477 );
nor \U$2462 ( \2805 , \2802 , \2804 );
nand \U$2463 ( \2806 , \2805 , \1737 );
nand \U$2464 ( \2807 , \2801 , \2806 );
xor \U$2465 ( \2808 , \2798 , \2807 );
or \U$2466 ( \2809 , \2646 , \1948 );
and \U$2467 ( \2810 , \1731 , \1313 );
and \U$2468 ( \2811 , \1733 , \1951 );
nor \U$2469 ( \2812 , \2810 , \2811 );
or \U$2470 ( \2813 , \2812 , \1954 );
nand \U$2471 ( \2814 , \2809 , \2813 );
xor \U$2472 ( \2815 , \2808 , \2814 );
xor \U$2473 ( \2816 , \2797 , \2815 );
xor \U$2474 ( \2817 , \2769 , \2816 );
xor \U$2475 ( \2818 , \2746 , \2817 );
xor \U$2476 ( \2819 , \2685 , \2717 );
and \U$2477 ( \2820 , \2819 , \2722 );
and \U$2478 ( \2821 , \2685 , \2717 );
or \U$2479 ( \2822 , \2820 , \2821 );
xor \U$2480 ( \2823 , \2818 , \2822 );
nor \U$2481 ( \2824 , \2738 , \2823 );
nor \U$2482 ( \2825 , \2734 , \2824 );
xor \U$2483 ( \2826 , \2746 , \2817 );
and \U$2484 ( \2827 , \2826 , \2822 );
and \U$2485 ( \2828 , \2746 , \2817 );
or \U$2486 ( \2829 , \2827 , \2828 );
xor \U$2487 ( \2830 , \2760 , \2768 );
and \U$2488 ( \2831 , \2830 , \2816 );
and \U$2489 ( \2832 , \2760 , \2768 );
or \U$2490 ( \2833 , \2831 , \2832 );
xor \U$2491 ( \2834 , \2798 , \2807 );
and \U$2492 ( \2835 , \2834 , \2814 );
and \U$2493 ( \2836 , \2798 , \2807 );
or \U$2494 ( \2837 , \2835 , \2836 );
or \U$2495 ( \2838 , \1011 , \1077 );
nand \U$2496 ( \2839 , \2838 , RIbb2f160_11);
or \U$2497 ( \2840 , \2789 , \1771 );
and \U$2498 ( \2841 , \814 , RIbb2f250_9);
and \U$2499 ( \2842 , \2251 , \1524 );
nor \U$2500 ( \2843 , \2841 , \2842 );
or \U$2501 ( \2844 , \2843 , \2133 );
nand \U$2502 ( \2845 , \2840 , \2844 );
xor \U$2503 ( \2846 , \2839 , \2845 );
not \U$2504 ( \2847 , \1147 );
and \U$2505 ( \2848 , \1940 , RIbb2f430_5);
not \U$2506 ( \2849 , \1940 );
and \U$2507 ( \2850 , \2849 , \1647 );
nor \U$2508 ( \2851 , \2848 , \2850 );
not \U$2509 ( \2852 , \2851 );
or \U$2510 ( \2853 , \2847 , \2852 );
or \U$2511 ( \2854 , \2776 , \1621 );
nand \U$2512 ( \2855 , \2853 , \2854 );
xor \U$2513 ( \2856 , \2846 , \2855 );
xor \U$2514 ( \2857 , \2837 , \2856 );
not \U$2515 ( \2858 , \1376 );
xor \U$2516 ( \2859 , \1313 , \1551 );
not \U$2517 ( \2860 , \2859 );
or \U$2518 ( \2861 , \2858 , \2860 );
or \U$2519 ( \2862 , \2812 , \1948 );
nand \U$2520 ( \2863 , \2861 , \2862 );
not \U$2521 ( \2864 , \1702 );
not \U$2522 ( \2865 , \2805 );
or \U$2523 ( \2866 , \2864 , \2865 );
and \U$2524 ( \2867 , \1514 , RIbb2f340_7);
and \U$2525 ( \2868 , \1511 , \1692 );
nor \U$2526 ( \2869 , \2867 , \2868 );
or \U$2527 ( \2870 , \2869 , \1738 );
nand \U$2528 ( \2871 , \2866 , \2870 );
xor \U$2529 ( \2872 , \2863 , \2871 );
or \U$2530 ( \2873 , \2782 , \1266 );
not \U$2531 ( \2874 , \1246 );
not \U$2532 ( \2875 , \1887 );
or \U$2533 ( \2876 , \2874 , \2875 );
nand \U$2534 ( \2877 , \1071 , \1291 );
nand \U$2535 ( \2878 , \2876 , \2877 );
not \U$2536 ( \2879 , \2878 );
or \U$2537 ( \2880 , \2879 , \1295 );
nand \U$2538 ( \2881 , \2873 , \2880 );
xor \U$2539 ( \2882 , \2872 , \2881 );
xor \U$2540 ( \2883 , \2857 , \2882 );
xor \U$2541 ( \2884 , \2833 , \2883 );
not \U$2542 ( \2885 , \1394 );
nor \U$2543 ( \2886 , \2885 , \1689 );
xor \U$2544 ( \2887 , \2753 , \2886 );
xor \U$2545 ( \2888 , \2778 , \2784 );
and \U$2546 ( \2889 , \2888 , \2791 );
and \U$2547 ( \2890 , \2778 , \2784 );
or \U$2548 ( \2891 , \2889 , \2890 );
xor \U$2549 ( \2892 , \2887 , \2891 );
xor \U$2550 ( \2893 , \2750 , \2754 );
and \U$2551 ( \2894 , \2893 , \2759 );
and \U$2552 ( \2895 , \2750 , \2754 );
or \U$2553 ( \2896 , \2894 , \2895 );
xor \U$2554 ( \2897 , \2792 , \2796 );
and \U$2555 ( \2898 , \2897 , \2815 );
and \U$2556 ( \2899 , \2792 , \2796 );
or \U$2557 ( \2900 , \2898 , \2899 );
xor \U$2558 ( \2901 , \2896 , \2900 );
xor \U$2559 ( \2902 , \2892 , \2901 );
xor \U$2560 ( \2903 , \2884 , \2902 );
or \U$2561 ( \2904 , \2829 , \2903 );
and \U$2562 ( \2905 , \2825 , \2904 );
and \U$2563 ( \2906 , \2642 , \2905 );
not \U$2564 ( \2907 , \2906 );
not \U$2565 ( \2908 , RIbb2e8f0_29);
not \U$2566 ( \2909 , \814 );
or \U$2567 ( \2910 , \2908 , \2909 );
not \U$2568 ( \2911 , RIbb2e8f0_29);
nand \U$2569 ( \2912 , \815 , \2911 );
nand \U$2570 ( \2913 , \2910 , \2912 );
and \U$2571 ( \2914 , RIbb2e8f0_29, RIbb2e878_30);
and \U$2572 ( \2915 , RIbb2e878_30, RIbb2e800_31);
not \U$2573 ( \2916 , RIbb2e878_30);
not \U$2574 ( \2917 , RIbb2e800_31);
and \U$2575 ( \2918 , \2916 , \2917 );
nor \U$2576 ( \2919 , \2915 , \2918 );
nor \U$2577 ( \2920 , RIbb2e8f0_29, RIbb2e878_30);
nor \U$2578 ( \2921 , \2914 , \2919 , \2920 );
buf \U$2579 ( \2922 , \2921 );
and \U$2580 ( \2923 , \2913 , \2922 );
buf \U$2581 ( \2924 , \2919 );
buf \U$2582 ( \2925 , \2924 );
and \U$2583 ( \2926 , \2925 , RIbb2e8f0_29);
nor \U$2584 ( \2927 , \2923 , \2926 );
and \U$2585 ( \2928 , RIbb2e788_32, RIbb2e800_31);
not \U$2586 ( \2929 , RIbb2e788_32);
and \U$2587 ( \2930 , \2929 , \2917 );
nor \U$2588 ( \2931 , \2928 , \2930 );
not \U$2589 ( \2932 , \2931 );
and \U$2590 ( \2933 , RIbb2e788_32, RIbb2e710_33);
not \U$2591 ( \2934 , RIbb2e788_32);
not \U$2592 ( \2935 , RIbb2e710_33);
and \U$2593 ( \2936 , \2934 , \2935 );
nor \U$2594 ( \2937 , \2933 , \2936 );
nor \U$2595 ( \2938 , \2932 , \2937 );
buf \U$2596 ( \2939 , \2938 );
buf \U$2597 ( \2940 , \2939 );
buf \U$2598 ( \2941 , \2937 );
or \U$2599 ( \2942 , \2940 , \2941 );
nand \U$2600 ( \2943 , \2942 , RIbb2e800_31);
not \U$2601 ( \2944 , \2922 );
not \U$2602 ( \2945 , RIbb2e8f0_29);
not \U$2603 ( \2946 , \893 );
not \U$2604 ( \2947 , \2946 );
or \U$2605 ( \2948 , \2945 , \2947 );
not \U$2606 ( \2949 , RIbb2e8f0_29);
nand \U$2607 ( \2950 , \1580 , \2949 );
nand \U$2608 ( \2951 , \2948 , \2950 );
not \U$2609 ( \2952 , \2951 );
or \U$2610 ( \2953 , \2944 , \2952 );
nand \U$2611 ( \2954 , \2913 , \2925 );
nand \U$2612 ( \2955 , \2953 , \2954 );
xor \U$2613 ( \2956 , \2943 , \2955 );
not \U$2614 ( \2957 , RIbb2ea58_26);
and \U$2615 ( \2958 , RIbb2e9e0_27, \2957 );
not \U$2616 ( \2959 , RIbb2e9e0_27);
and \U$2617 ( \2960 , \2959 , RIbb2ea58_26);
nor \U$2618 ( \2961 , \2958 , \2960 );
not \U$2619 ( \2962 , \2961 );
buf \U$2620 ( \2963 , \2962 );
not \U$2621 ( \2964 , \2963 );
and \U$2622 ( \2965 , RIbb2ead0_25, \988 );
not \U$2623 ( \2966 , RIbb2ead0_25);
and \U$2624 ( \2967 , \2966 , \987 );
or \U$2625 ( \2968 , \2965 , \2967 );
not \U$2626 ( \2969 , \2968 );
or \U$2627 ( \2970 , \2964 , \2969 );
and \U$2628 ( \2971 , RIbb2ead0_25, \953 );
not \U$2629 ( \2972 , RIbb2ead0_25);
and \U$2630 ( \2973 , \2972 , \957 );
or \U$2631 ( \2974 , \2971 , \2973 );
and \U$2632 ( \2975 , RIbb2ead0_25, RIbb2ea58_26);
not \U$2633 ( \2976 , RIbb2ead0_25);
and \U$2634 ( \2977 , \2976 , \2957 );
nor \U$2635 ( \2978 , \2975 , \2977 );
and \U$2636 ( \2979 , \2961 , \2978 );
buf \U$2637 ( \2980 , \2979 );
nand \U$2638 ( \2981 , \2974 , \2980 );
nand \U$2639 ( \2982 , \2970 , \2981 );
and \U$2640 ( \2983 , \2956 , \2982 );
and \U$2641 ( \2984 , \2943 , \2955 );
or \U$2642 ( \2985 , \2983 , \2984 );
xor \U$2643 ( \2986 , \2927 , \2985 );
not \U$2644 ( \2987 , \377 );
not \U$2645 ( \2988 , \665 );
or \U$2646 ( \2989 , \2987 , \2988 );
not \U$2647 ( \2990 , \676 );
and \U$2648 ( \2991 , RIbb2ca00_95, RIbb32400_159);
nor \U$2649 ( \2992 , \2990 , \2991 );
nand \U$2650 ( \2993 , \2989 , \2992 );
not \U$2651 ( \2994 , \671 );
nor \U$2652 ( \2995 , \2994 , \373 );
and \U$2653 ( \2996 , \2993 , \2995 );
not \U$2654 ( \2997 , \2993 );
not \U$2655 ( \2998 , \2995 );
and \U$2656 ( \2999 , \2997 , \2998 );
nor \U$2657 ( \3000 , \2996 , \2999 );
not \U$2658 ( \3001 , \3000 );
not \U$2659 ( \3002 , \3001 );
buf \U$2660 ( \3003 , \3002 );
and \U$2661 ( \3004 , \3003 , \1313 );
not \U$2662 ( \3005 , \1376 );
buf \U$2663 ( \3006 , \378 );
not \U$2664 ( \3007 , \3006 );
not \U$2665 ( \3008 , \3007 );
not \U$2666 ( \3009 , \866 );
or \U$2667 ( \3010 , \3008 , \3009 );
not \U$2668 ( \3011 , \680 );
nand \U$2669 ( \3012 , \3011 , \677 );
nand \U$2670 ( \3013 , \3010 , \3012 );
not \U$2671 ( \3014 , \383 );
nand \U$2672 ( \3015 , \3014 , \690 );
not \U$2673 ( \3016 , \3015 );
and \U$2674 ( \3017 , \3013 , \3016 );
not \U$2675 ( \3018 , \3013 );
and \U$2676 ( \3019 , \3018 , \3015 );
nor \U$2677 ( \3020 , \3017 , \3019 );
not \U$2678 ( \3021 , \3020 );
not \U$2679 ( \3022 , \3021 );
not \U$2680 ( \3023 , \3022 );
not \U$2681 ( \3024 , \3023 );
xor \U$2682 ( \3025 , \1393 , \3024 );
not \U$2683 ( \3026 , \3025 );
or \U$2684 ( \3027 , \3005 , \3026 );
not \U$2685 ( \3028 , \377 );
nor \U$2686 ( \3029 , \3028 , \373 );
not \U$2687 ( \3030 , \3029 );
not \U$2688 ( \3031 , \665 );
or \U$2689 ( \3032 , \3030 , \3031 );
not \U$2690 ( \3033 , \2992 );
not \U$2691 ( \3034 , \373 );
and \U$2692 ( \3035 , \3033 , \3034 );
nor \U$2693 ( \3036 , \3035 , \2994 );
nand \U$2694 ( \3037 , \3032 , \3036 );
nor \U$2695 ( \3038 , \679 , \372 );
and \U$2696 ( \3039 , \3037 , \3038 );
not \U$2697 ( \3040 , \3037 );
not \U$2698 ( \3041 , \3038 );
and \U$2699 ( \3042 , \3040 , \3041 );
nor \U$2700 ( \3043 , \3039 , \3042 );
buf \U$2701 ( \3044 , \3043 );
not \U$2702 ( \3045 , \3044 );
not \U$2703 ( \3046 , \3045 );
xor \U$2704 ( \3047 , \1393 , \3046 );
nand \U$2705 ( \3048 , \3047 , \1430 );
nand \U$2706 ( \3049 , \3027 , \3048 );
xor \U$2707 ( \3050 , \3004 , \3049 );
not \U$2708 ( \3051 , \836 );
not \U$2709 ( \3052 , RIbb2ee90_17);
not \U$2710 ( \3053 , \1135 );
not \U$2711 ( \3054 , \3053 );
not \U$2712 ( \3055 , \3054 );
or \U$2713 ( \3056 , \3052 , \3055 );
not \U$2714 ( \3057 , RIbb2ee90_17);
nand \U$2715 ( \3058 , \1139 , \3057 );
nand \U$2716 ( \3059 , \3056 , \3058 );
not \U$2717 ( \3060 , \3059 );
or \U$2718 ( \3061 , \3051 , \3060 );
not \U$2719 ( \3062 , RIbb2ee90_17);
not \U$2720 ( \3063 , \1113 );
or \U$2721 ( \3064 , \3062 , \3063 );
buf \U$2722 ( \3065 , \1110 );
buf \U$2723 ( \3066 , \3065 );
not \U$2724 ( \3067 , \3066 );
nand \U$2725 ( \3068 , \3067 , \816 );
nand \U$2726 ( \3069 , \3064 , \3068 );
nand \U$2727 ( \3070 , \3069 , \832 );
nand \U$2728 ( \3071 , \3061 , \3070 );
and \U$2729 ( \3072 , \3050 , \3071 );
and \U$2730 ( \3073 , \3004 , \3049 );
or \U$2731 ( \3074 , \3072 , \3073 );
xor \U$2732 ( \3075 , \2986 , \3074 );
not \U$2733 ( \3076 , \376 );
not \U$2734 ( \3077 , \3076 );
not \U$2735 ( \3078 , \665 );
or \U$2736 ( \3079 , \3077 , \3078 );
nand \U$2737 ( \3080 , RIbb2c988_96, RIbb32478_160);
buf \U$2738 ( \3081 , \3080 );
nand \U$2739 ( \3082 , \3079 , \3081 );
nor \U$2740 ( \3083 , \2991 , \375 );
and \U$2741 ( \3084 , \3082 , \3083 );
not \U$2742 ( \3085 , \3082 );
not \U$2743 ( \3086 , \3083 );
and \U$2744 ( \3087 , \3085 , \3086 );
nor \U$2745 ( \3088 , \3084 , \3087 );
buf \U$2746 ( \3089 , \3088 );
not \U$2747 ( \3090 , \3089 );
not \U$2748 ( \3091 , \3090 );
buf \U$2749 ( \3092 , \3091 );
and \U$2750 ( \3093 , \3092 , \1394 );
not \U$2751 ( \3094 , \2963 );
not \U$2752 ( \3095 , \2974 );
or \U$2753 ( \3096 , \3094 , \3095 );
and \U$2754 ( \3097 , RIbb2ead0_25, \1887 );
not \U$2755 ( \3098 , RIbb2ead0_25);
not \U$2756 ( \3099 , \1887 );
and \U$2757 ( \3100 , \3098 , \3099 );
or \U$2758 ( \3101 , \3097 , \3100 );
nand \U$2759 ( \3102 , \3101 , \2980 );
nand \U$2760 ( \3103 , \3096 , \3102 );
xor \U$2761 ( \3104 , \3093 , \3103 );
buf \U$2762 ( \3105 , \1517 );
not \U$2763 ( \3106 , \3105 );
and \U$2764 ( \3107 , RIbb2ef80_15, \1170 );
not \U$2765 ( \3108 , RIbb2ef80_15);
buf \U$2766 ( \3109 , \1169 );
and \U$2767 ( \3110 , \3108 , \3109 );
or \U$2768 ( \3111 , \3107 , \3110 );
not \U$2769 ( \3112 , \3111 );
or \U$2770 ( \3113 , \3106 , \3112 );
and \U$2771 ( \3114 , RIbb2ef80_15, \1820 );
not \U$2772 ( \3115 , RIbb2ef80_15);
not \U$2773 ( \3116 , \1386 );
not \U$2774 ( \3117 , \3116 );
and \U$2775 ( \3118 , \3115 , \3117 );
or \U$2776 ( \3119 , \3114 , \3118 );
nand \U$2777 ( \3120 , \3119 , \1445 );
nand \U$2778 ( \3121 , \3113 , \3120 );
and \U$2779 ( \3122 , \3104 , \3121 );
and \U$2780 ( \3123 , \3093 , \3103 );
or \U$2781 ( \3124 , \3122 , \3123 );
not \U$2782 ( \3125 , \1702 );
not \U$2783 ( \3126 , RIbb2f340_7);
not \U$2784 ( \3127 , \1315 );
not \U$2785 ( \3128 , \665 );
or \U$2786 ( \3129 , \3127 , \3128 );
not \U$2787 ( \3130 , \1156 );
nand \U$2788 ( \3131 , \3129 , \3130 );
not \U$2789 ( \3132 , \388 );
nand \U$2790 ( \3133 , \3132 , \708 );
not \U$2791 ( \3134 , \3133 );
and \U$2792 ( \3135 , \3131 , \3134 );
not \U$2793 ( \3136 , \3131 );
and \U$2794 ( \3137 , \3136 , \3133 );
nor \U$2795 ( \3138 , \3135 , \3137 );
buf \U$2796 ( \3139 , \3138 );
not \U$2797 ( \3140 , \3139 );
buf \U$2798 ( \3141 , \3140 );
not \U$2799 ( \3142 , \3141 );
not \U$2800 ( \3143 , \3142 );
not \U$2801 ( \3144 , \3143 );
or \U$2802 ( \3145 , \3126 , \3144 );
buf \U$2803 ( \3146 , \3139 );
nand \U$2804 ( \3147 , \3146 , \2700 );
nand \U$2805 ( \3148 , \3145 , \3147 );
not \U$2806 ( \3149 , \3148 );
or \U$2807 ( \3150 , \3125 , \3149 );
not \U$2808 ( \3151 , RIbb2f340_7);
and \U$2809 ( \3152 , \1315 , \3132 );
not \U$2810 ( \3153 , \3152 );
not \U$2811 ( \3154 , \665 );
or \U$2812 ( \3155 , \3153 , \3154 );
nand \U$2813 ( \3156 , \1156 , \3132 );
and \U$2814 ( \3157 , \3156 , \708 );
nand \U$2815 ( \3158 , \3155 , \3157 );
not \U$2816 ( \3159 , \710 );
nor \U$2817 ( \3160 , \3159 , \387 );
and \U$2818 ( \3161 , \3158 , \3160 );
not \U$2819 ( \3162 , \3158 );
not \U$2820 ( \3163 , \3160 );
and \U$2821 ( \3164 , \3162 , \3163 );
nor \U$2822 ( \3165 , \3161 , \3164 );
buf \U$2823 ( \3166 , \3165 );
buf \U$2824 ( \3167 , \3166 );
not \U$2825 ( \3168 , \3167 );
not \U$2826 ( \3169 , \3168 );
or \U$2827 ( \3170 , \3151 , \3169 );
nand \U$2828 ( \3171 , \3167 , \1692 );
nand \U$2829 ( \3172 , \3170 , \3171 );
nand \U$2830 ( \3173 , \3172 , \1737 );
nand \U$2831 ( \3174 , \3150 , \3173 );
not \U$2832 ( \3175 , \3174 );
not \U$2833 ( \3176 , \1147 );
not \U$2834 ( \3177 , RIbb2f430_5);
not \U$2835 ( \3178 , \379 );
nand \U$2836 ( \3179 , \384 , \3178 );
nor \U$2837 ( \3180 , \3179 , \3006 );
not \U$2838 ( \3181 , \3180 );
not \U$2839 ( \3182 , \866 );
or \U$2840 ( \3183 , \3181 , \3182 );
not \U$2841 ( \3184 , \3012 );
not \U$2842 ( \3185 , \3179 );
and \U$2843 ( \3186 , \3184 , \3185 );
not \U$2844 ( \3187 , \3178 );
not \U$2845 ( \3188 , \693 );
or \U$2846 ( \3189 , \3187 , \3188 );
nand \U$2847 ( \3190 , \3189 , \695 );
nor \U$2848 ( \3191 , \3186 , \3190 );
nand \U$2849 ( \3192 , \3183 , \3191 );
not \U$2850 ( \3193 , \697 );
nor \U$2851 ( \3194 , \3193 , \380 );
and \U$2852 ( \3195 , \3192 , \3194 );
not \U$2853 ( \3196 , \3192 );
not \U$2854 ( \3197 , \3194 );
and \U$2855 ( \3198 , \3196 , \3197 );
nor \U$2856 ( \3199 , \3195 , \3198 );
not \U$2857 ( \3200 , \3199 );
not \U$2858 ( \3201 , \3200 );
buf \U$2859 ( \3202 , \3201 );
not \U$2860 ( \3203 , \3202 );
not \U$2861 ( \3204 , \3203 );
or \U$2862 ( \3205 , \3177 , \3204 );
nand \U$2863 ( \3206 , \3202 , \1085 );
nand \U$2864 ( \3207 , \3205 , \3206 );
not \U$2865 ( \3208 , \3207 );
or \U$2866 ( \3209 , \3176 , \3208 );
not \U$2867 ( \3210 , \384 );
nor \U$2868 ( \3211 , \3210 , \3006 );
not \U$2869 ( \3212 , \3211 );
not \U$2870 ( \3213 , \665 );
or \U$2871 ( \3214 , \3212 , \3213 );
and \U$2872 ( \3215 , \3184 , \384 );
nor \U$2873 ( \3216 , \3215 , \693 );
nand \U$2874 ( \3217 , \3214 , \3216 );
nand \U$2875 ( \3218 , \3178 , \695 );
not \U$2876 ( \3219 , \3218 );
and \U$2877 ( \3220 , \3217 , \3219 );
not \U$2878 ( \3221 , \3217 );
and \U$2879 ( \3222 , \3221 , \3218 );
nor \U$2880 ( \3223 , \3220 , \3222 );
buf \U$2881 ( \3224 , \3223 );
not \U$2882 ( \3225 , \3224 );
buf \U$2883 ( \3226 , \3225 );
nand \U$2884 ( \3227 , RIbb2f430_5, \3226 );
buf \U$2885 ( \3228 , \3224 );
nand \U$2886 ( \3229 , \3228 , \1980 );
nand \U$2887 ( \3230 , \3227 , \3229 );
nand \U$2888 ( \3231 , \3230 , \1090 );
nand \U$2889 ( \3232 , \3209 , \3231 );
not \U$2890 ( \3233 , \3232 );
or \U$2891 ( \3234 , \3175 , \3233 );
or \U$2892 ( \3235 , \3232 , \3174 );
not \U$2893 ( \3236 , \855 );
not \U$2894 ( \3237 , RIbb2eda0_19);
not \U$2895 ( \3238 , \1640 );
buf \U$2896 ( \3239 , \3238 );
not \U$2897 ( \3240 , \3239 );
or \U$2898 ( \3241 , \3237 , \3240 );
buf \U$2899 ( \3242 , \1641 );
not \U$2900 ( \3243 , \3242 );
nand \U$2901 ( \3244 , \3243 , \1776 );
nand \U$2902 ( \3245 , \3241 , \3244 );
not \U$2903 ( \3246 , \3245 );
or \U$2904 ( \3247 , \3236 , \3246 );
not \U$2905 ( \3248 , RIbb2eda0_19);
not \U$2906 ( \3249 , \3054 );
or \U$2907 ( \3250 , \3248 , \3249 );
not \U$2908 ( \3251 , RIbb2eda0_19);
nand \U$2909 ( \3252 , \1138 , \3251 );
nand \U$2910 ( \3253 , \3250 , \3252 );
nand \U$2911 ( \3254 , \3253 , \853 );
nand \U$2912 ( \3255 , \3247 , \3254 );
nand \U$2913 ( \3256 , \3235 , \3255 );
nand \U$2914 ( \3257 , \3234 , \3256 );
xor \U$2915 ( \3258 , \3124 , \3257 );
not \U$2916 ( \3259 , \2922 );
not \U$2917 ( \3260 , RIbb2e8f0_29);
buf \U$2918 ( \3261 , \1508 );
not \U$2919 ( \3262 , \3261 );
not \U$2920 ( \3263 , \3262 );
or \U$2921 ( \3264 , \3260 , \3263 );
not \U$2922 ( \3265 , RIbb2e8f0_29);
nand \U$2923 ( \3266 , \3261 , \3265 );
nand \U$2924 ( \3267 , \3264 , \3266 );
not \U$2925 ( \3268 , \3267 );
or \U$2926 ( \3269 , \3259 , \3268 );
nand \U$2927 ( \3270 , \2951 , \2925 );
nand \U$2928 ( \3271 , \3269 , \3270 );
not \U$2929 ( \3272 , \1430 );
not \U$2930 ( \3273 , \1394 );
buf \U$2931 ( \3274 , \3000 );
buf \U$2932 ( \3275 , \3274 );
not \U$2933 ( \3276 , \3275 );
not \U$2934 ( \3277 , \3276 );
or \U$2935 ( \3278 , \3273 , \3277 );
nand \U$2936 ( \3279 , \3003 , \1951 );
nand \U$2937 ( \3280 , \3278 , \3279 );
not \U$2938 ( \3281 , \3280 );
or \U$2939 ( \3282 , \3272 , \3281 );
nand \U$2940 ( \3283 , \3047 , \1376 );
nand \U$2941 ( \3284 , \3282 , \3283 );
xor \U$2942 ( \3285 , \3271 , \3284 );
not \U$2943 ( \3286 , \832 );
not \U$2944 ( \3287 , RIbb2ee90_17);
not \U$2945 ( \3288 , \1284 );
or \U$2946 ( \3289 , \3287 , \3288 );
not \U$2947 ( \3290 , \1282 );
not \U$2948 ( \3291 , \3290 );
nand \U$2949 ( \3292 , \3291 , \2240 );
nand \U$2950 ( \3293 , \3289 , \3292 );
not \U$2951 ( \3294 , \3293 );
or \U$2952 ( \3295 , \3286 , \3294 );
nand \U$2953 ( \3296 , \3069 , \836 );
nand \U$2954 ( \3297 , \3295 , \3296 );
and \U$2955 ( \3298 , \3285 , \3297 );
and \U$2956 ( \3299 , \3271 , \3284 );
or \U$2957 ( \3300 , \3298 , \3299 );
and \U$2958 ( \3301 , \3258 , \3300 );
and \U$2959 ( \3302 , \3124 , \3257 );
or \U$2960 ( \3303 , \3301 , \3302 );
xor \U$2961 ( \3304 , \3075 , \3303 );
not \U$2962 ( \3305 , \1570 );
not \U$2963 ( \3306 , RIbb2f250_9);
not \U$2964 ( \3307 , \2116 );
or \U$2965 ( \3308 , \3306 , \3307 );
buf \U$2966 ( \3309 , \2113 );
not \U$2967 ( \3310 , \3309 );
not \U$2968 ( \3311 , \3310 );
nand \U$2969 ( \3312 , \3311 , \1566 );
nand \U$2970 ( \3313 , \3308 , \3312 );
not \U$2971 ( \3314 , \3313 );
or \U$2972 ( \3315 , \3305 , \3314 );
not \U$2973 ( \3316 , RIbb2f250_9);
not \U$2974 ( \3317 , \2224 );
or \U$2975 ( \3318 , \3316 , \3317 );
not \U$2976 ( \3319 , \2222 );
not \U$2977 ( \3320 , \3319 );
nand \U$2978 ( \3321 , \3320 , \1554 );
nand \U$2979 ( \3322 , \3318 , \3321 );
nand \U$2980 ( \3323 , \3322 , \1533 );
nand \U$2981 ( \3324 , \3315 , \3323 );
not \U$2982 ( \3325 , \3324 );
not \U$2983 ( \3326 , \1737 );
not \U$2984 ( \3327 , RIbb2f340_7);
and \U$2985 ( \3328 , \1315 , \2202 );
not \U$2986 ( \3329 , \3328 );
not \U$2987 ( \3330 , \866 );
or \U$2988 ( \3331 , \3329 , \3330 );
and \U$2989 ( \3332 , \1156 , \2202 );
nor \U$2990 ( \3333 , \3332 , \711 );
nand \U$2991 ( \3334 , \3331 , \3333 );
nor \U$2992 ( \3335 , \714 , \391 );
and \U$2993 ( \3336 , \3334 , \3335 );
not \U$2994 ( \3337 , \3334 );
not \U$2995 ( \3338 , \3335 );
and \U$2996 ( \3339 , \3337 , \3338 );
nor \U$2997 ( \3340 , \3336 , \3339 );
buf \U$2998 ( \3341 , \3340 );
not \U$2999 ( \3342 , \3341 );
not \U$3000 ( \3343 , \3342 );
not \U$3001 ( \3344 , \3343 );
not \U$3002 ( \3345 , \3344 );
or \U$3003 ( \3346 , \3327 , \3345 );
not \U$3004 ( \3347 , \3344 );
nand \U$3005 ( \3348 , \3347 , \1692 );
nand \U$3006 ( \3349 , \3346 , \3348 );
not \U$3007 ( \3350 , \3349 );
or \U$3008 ( \3351 , \3326 , \3350 );
nand \U$3009 ( \3352 , \3172 , \1702 );
nand \U$3010 ( \3353 , \3351 , \3352 );
not \U$3011 ( \3354 , \3353 );
or \U$3012 ( \3355 , \3325 , \3354 );
not \U$3013 ( \3356 , \3353 );
not \U$3014 ( \3357 , \3356 );
not \U$3015 ( \3358 , \3324 );
not \U$3016 ( \3359 , \3358 );
or \U$3017 ( \3360 , \3357 , \3359 );
not \U$3018 ( \3361 , \855 );
not \U$3019 ( \3362 , RIbb2eda0_19);
buf \U$3020 ( \3363 , \1685 );
buf \U$3021 ( \3364 , \3363 );
not \U$3022 ( \3365 , \3364 );
not \U$3023 ( \3366 , \3365 );
or \U$3024 ( \3367 , \3362 , \3366 );
not \U$3025 ( \3368 , \1685 );
not \U$3026 ( \3369 , \3368 );
not \U$3027 ( \3370 , \3369 );
not \U$3028 ( \3371 , \3370 );
nand \U$3029 ( \3372 , \3371 , \1776 );
nand \U$3030 ( \3373 , \3367 , \3372 );
not \U$3031 ( \3374 , \3373 );
or \U$3032 ( \3375 , \3361 , \3374 );
nand \U$3033 ( \3376 , \3245 , \853 );
nand \U$3034 ( \3377 , \3375 , \3376 );
nand \U$3035 ( \3378 , \3360 , \3377 );
nand \U$3036 ( \3379 , \3355 , \3378 );
xor \U$3037 ( \3380 , RIbb2eb48_24, RIbb2ead0_25);
buf \U$3038 ( \3381 , \3380 );
buf \U$3039 ( \3382 , \3381 );
buf \U$3040 ( \3383 , \3382 );
not \U$3041 ( \3384 , \3383 );
not \U$3042 ( \3385 , RIbb2ebc0_23);
not \U$3043 ( \3386 , \1072 );
or \U$3044 ( \3387 , \3385 , \3386 );
not \U$3045 ( \3388 , RIbb2ebc0_23);
nand \U$3046 ( \3389 , \3099 , \3388 );
nand \U$3047 ( \3390 , \3387 , \3389 );
not \U$3048 ( \3391 , \3390 );
or \U$3049 ( \3392 , \3384 , \3391 );
not \U$3050 ( \3393 , RIbb2ebc0_23);
not \U$3051 ( \3394 , \1562 );
or \U$3052 ( \3395 , \3393 , \3394 );
not \U$3053 ( \3396 , RIbb2ebc0_23);
nand \U$3054 ( \3397 , \1042 , \3396 );
nand \U$3055 ( \3398 , \3395 , \3397 );
and \U$3056 ( \3399 , RIbb2eb48_24, RIbb2ebc0_23);
not \U$3057 ( \3400 , RIbb2eb48_24);
not \U$3058 ( \3401 , RIbb2ebc0_23);
and \U$3059 ( \3402 , \3400 , \3401 );
nor \U$3060 ( \3403 , \3399 , \3402 );
not \U$3061 ( \3404 , \3403 );
nor \U$3062 ( \3405 , \3404 , \3380 );
buf \U$3063 ( \3406 , \3405 );
buf \U$3064 ( \3407 , \3406 );
nand \U$3065 ( \3408 , \3398 , \3407 );
nand \U$3066 ( \3409 , \3392 , \3408 );
not \U$3067 ( \3410 , \1445 );
not \U$3068 ( \3411 , \3111 );
or \U$3069 ( \3412 , \3410 , \3411 );
xnor \U$3070 ( \3413 , RIbb2ef80_15, \1284 );
nand \U$3071 ( \3414 , \3413 , \3105 );
nand \U$3072 ( \3415 , \3412 , \3414 );
xor \U$3073 ( \3416 , \3409 , \3415 );
not \U$3074 ( \3417 , \998 );
not \U$3075 ( \3418 , RIbb2f070_13);
not \U$3076 ( \3419 , \1820 );
or \U$3077 ( \3420 , \3418 , \3419 );
not \U$3078 ( \3421 , RIbb2f070_13);
nand \U$3079 ( \3422 , \1387 , \3421 );
nand \U$3080 ( \3423 , \3420 , \3422 );
not \U$3081 ( \3424 , \3423 );
or \U$3082 ( \3425 , \3417 , \3424 );
not \U$3083 ( \3426 , RIbb2f070_13);
not \U$3084 ( \3427 , \2052 );
or \U$3085 ( \3428 , \3426 , \3427 );
nand \U$3086 ( \3429 , \1422 , \906 );
nand \U$3087 ( \3430 , \3428 , \3429 );
nand \U$3088 ( \3431 , \3430 , \916 );
nand \U$3089 ( \3432 , \3425 , \3431 );
and \U$3090 ( \3433 , \3416 , \3432 );
and \U$3091 ( \3434 , \3409 , \3415 );
or \U$3092 ( \3435 , \3433 , \3434 );
xor \U$3093 ( \3436 , \3379 , \3435 );
and \U$3094 ( \3437 , RIbb2e9e0_27, RIbb2e968_28);
and \U$3095 ( \3438 , RIbb2e968_28, RIbb2e8f0_29);
not \U$3096 ( \3439 , RIbb2e968_28);
not \U$3097 ( \3440 , RIbb2e8f0_29);
and \U$3098 ( \3441 , \3439 , \3440 );
nor \U$3099 ( \3442 , \3438 , \3441 );
nor \U$3100 ( \3443 , RIbb2e9e0_27, RIbb2e968_28);
nor \U$3101 ( \3444 , \3437 , \3442 , \3443 );
buf \U$3102 ( \3445 , \3444 );
not \U$3103 ( \3446 , \3445 );
not \U$3104 ( \3447 , RIbb2e9e0_27);
not \U$3105 ( \3448 , \1475 );
or \U$3106 ( \3449 , \3447 , \3448 );
buf \U$3107 ( \3450 , \1472 );
not \U$3108 ( \3451 , \3450 );
buf \U$3109 ( \3452 , \3451 );
not \U$3110 ( \3453 , \3452 );
not \U$3111 ( \3454 , RIbb2e9e0_27);
nand \U$3112 ( \3455 , \3453 , \3454 );
nand \U$3113 ( \3456 , \3449 , \3455 );
not \U$3114 ( \3457 , \3456 );
or \U$3115 ( \3458 , \3446 , \3457 );
not \U$3116 ( \3459 , RIbb2e9e0_27);
not \U$3117 ( \3460 , \1509 );
or \U$3118 ( \3461 , \3459 , \3460 );
not \U$3119 ( \3462 , RIbb2e9e0_27);
nand \U$3120 ( \3463 , \3261 , \3462 );
nand \U$3121 ( \3464 , \3461 , \3463 );
buf \U$3122 ( \3465 , \3442 );
nand \U$3123 ( \3466 , \3464 , \3465 );
nand \U$3124 ( \3467 , \3458 , \3466 );
not \U$3125 ( \3468 , \2078 );
not \U$3126 ( \3469 , RIbb2ecb0_21);
not \U$3127 ( \3470 , \1550 );
or \U$3128 ( \3471 , \3469 , \3470 );
not \U$3129 ( \3472 , \1550 );
nand \U$3130 ( \3473 , \3472 , \849 );
nand \U$3131 ( \3474 , \3471 , \3473 );
not \U$3132 ( \3475 , \3474 );
or \U$3133 ( \3476 , \3468 , \3475 );
not \U$3134 ( \3477 , RIbb2ecb0_21);
buf \U$3135 ( \3478 , \1728 );
not \U$3136 ( \3479 , \3478 );
not \U$3137 ( \3480 , \3479 );
not \U$3138 ( \3481 , \3480 );
not \U$3139 ( \3482 , \3481 );
or \U$3140 ( \3483 , \3477 , \3482 );
buf \U$3141 ( \3484 , \3478 );
nand \U$3142 ( \3485 , \3484 , \2254 );
nand \U$3143 ( \3486 , \3483 , \3485 );
nand \U$3144 ( \3487 , \2077 , \3486 );
nand \U$3145 ( \3488 , \3476 , \3487 );
xor \U$3146 ( \3489 , \3467 , \3488 );
not \U$3147 ( \3490 , \1077 );
not \U$3148 ( \3491 , RIbb2f160_11);
not \U$3149 ( \3492 , \1340 );
or \U$3150 ( \3493 , \3491 , \3492 );
not \U$3151 ( \3494 , \1337 );
not \U$3152 ( \3495 , \3494 );
nand \U$3153 ( \3496 , \3495 , \1805 );
nand \U$3154 ( \3497 , \3493 , \3496 );
not \U$3155 ( \3498 , \3497 );
or \U$3156 ( \3499 , \3490 , \3498 );
not \U$3157 ( \3500 , RIbb2f160_11);
not \U$3158 ( \3501 , \1854 );
or \U$3159 ( \3502 , \3500 , \3501 );
not \U$3160 ( \3503 , \1854 );
nand \U$3161 ( \3504 , \3503 , \1805 );
nand \U$3162 ( \3505 , \3502 , \3504 );
nand \U$3163 ( \3506 , \3505 , \1011 );
nand \U$3164 ( \3507 , \3499 , \3506 );
and \U$3165 ( \3508 , \3489 , \3507 );
and \U$3166 ( \3509 , \3467 , \3488 );
or \U$3167 ( \3510 , \3508 , \3509 );
xor \U$3168 ( \3511 , \3436 , \3510 );
xnor \U$3169 ( \3512 , \3304 , \3511 );
not \U$3170 ( \3513 , \3512 );
not \U$3171 ( \3514 , \1533 );
not \U$3172 ( \3515 , RIbb2f250_9);
not \U$3173 ( \3516 , \3341 );
buf \U$3174 ( \3517 , \3516 );
not \U$3175 ( \3518 , \3517 );
or \U$3176 ( \3519 , \3515 , \3518 );
not \U$3177 ( \3520 , \3341 );
not \U$3178 ( \3521 , \3520 );
nand \U$3179 ( \3522 , \3521 , \1566 );
nand \U$3180 ( \3523 , \3519 , \3522 );
not \U$3181 ( \3524 , \3523 );
or \U$3182 ( \3525 , \3514 , \3524 );
nand \U$3183 ( \3526 , \3322 , \1570 );
nand \U$3184 ( \3527 , \3525 , \3526 );
not \U$3185 ( \3528 , \3527 );
not \U$3186 ( \3529 , \3465 );
not \U$3187 ( \3530 , \3456 );
or \U$3188 ( \3531 , \3529 , \3530 );
not \U$3189 ( \3532 , RIbb2e9e0_27);
not \U$3190 ( \3533 , \992 );
or \U$3191 ( \3534 , \3532 , \3533 );
nand \U$3192 ( \3535 , \994 , \3462 );
nand \U$3193 ( \3536 , \3534 , \3535 );
nand \U$3194 ( \3537 , \3536 , \3445 );
nand \U$3195 ( \3538 , \3531 , \3537 );
not \U$3196 ( \3539 , \3538 );
or \U$3197 ( \3540 , \3528 , \3539 );
not \U$3198 ( \3541 , \3538 );
not \U$3199 ( \3542 , \3541 );
not \U$3200 ( \3543 , \3527 );
not \U$3201 ( \3544 , \3543 );
or \U$3202 ( \3545 , \3542 , \3544 );
not \U$3203 ( \3546 , \2078 );
not \U$3204 ( \3547 , \3486 );
or \U$3205 ( \3548 , \3546 , \3547 );
not \U$3206 ( \3549 , RIbb2ecb0_21);
not \U$3207 ( \3550 , \1689 );
or \U$3208 ( \3551 , \3549 , \3550 );
buf \U$3209 ( \3552 , \1687 );
nand \U$3210 ( \3553 , \3552 , \849 );
nand \U$3211 ( \3554 , \3551 , \3553 );
nand \U$3212 ( \3555 , \3554 , \2077 );
nand \U$3213 ( \3556 , \3548 , \3555 );
nand \U$3214 ( \3557 , \3545 , \3556 );
nand \U$3215 ( \3558 , \3540 , \3557 );
not \U$3216 ( \3559 , \1011 );
not \U$3217 ( \3560 , RIbb2f160_11);
not \U$3218 ( \3561 , \3310 );
or \U$3219 ( \3562 , \3560 , \3561 );
not \U$3220 ( \3563 , \2114 );
not \U$3221 ( \3564 , \3563 );
nand \U$3222 ( \3565 , \3564 , \1805 );
nand \U$3223 ( \3566 , \3562 , \3565 );
not \U$3224 ( \3567 , \3566 );
or \U$3225 ( \3568 , \3559 , \3567 );
nand \U$3226 ( \3569 , \3505 , \1077 );
nand \U$3227 ( \3570 , \3568 , \3569 );
not \U$3228 ( \3571 , \998 );
not \U$3229 ( \3572 , \3430 );
or \U$3230 ( \3573 , \3571 , \3572 );
not \U$3231 ( \3574 , RIbb2f070_13);
not \U$3232 ( \3575 , \3495 );
not \U$3233 ( \3576 , \3575 );
or \U$3234 ( \3577 , \3574 , \3576 );
nand \U$3235 ( \3578 , \1339 , \906 );
nand \U$3236 ( \3579 , \3577 , \3578 );
nand \U$3237 ( \3580 , \3579 , \916 );
nand \U$3238 ( \3581 , \3573 , \3580 );
xor \U$3239 ( \3582 , \3570 , \3581 );
not \U$3240 ( \3583 , \3407 );
not \U$3241 ( \3584 , RIbb2ebc0_23);
not \U$3242 ( \3585 , \1550 );
or \U$3243 ( \3586 , \3584 , \3585 );
nand \U$3244 ( \3587 , \1551 , \2073 );
nand \U$3245 ( \3588 , \3586 , \3587 );
not \U$3246 ( \3589 , \3588 );
or \U$3247 ( \3590 , \3583 , \3589 );
nand \U$3248 ( \3591 , \3398 , \3383 );
nand \U$3249 ( \3592 , \3590 , \3591 );
and \U$3250 ( \3593 , \3582 , \3592 );
and \U$3251 ( \3594 , \3570 , \3581 );
or \U$3252 ( \3595 , \3593 , \3594 );
xor \U$3253 ( \3596 , \3558 , \3595 );
xor \U$3254 ( \3597 , \3004 , \3049 );
xor \U$3255 ( \3598 , \3597 , \3071 );
and \U$3256 ( \3599 , \3596 , \3598 );
and \U$3257 ( \3600 , \3558 , \3595 );
or \U$3258 ( \3601 , \3599 , \3600 );
xor \U$3259 ( \3602 , \2943 , \2955 );
xor \U$3260 ( \3603 , \3602 , \2982 );
not \U$3261 ( \3604 , \2940 );
not \U$3262 ( \3605 , RIbb2e800_31);
not \U$3263 ( \3606 , \814 );
or \U$3264 ( \3607 , \3605 , \3606 );
not \U$3265 ( \3608 , RIbb2e800_31);
nand \U$3266 ( \3609 , \2251 , \3608 );
nand \U$3267 ( \3610 , \3607 , \3609 );
not \U$3268 ( \3611 , \3610 );
or \U$3269 ( \3612 , \3604 , \3611 );
buf \U$3270 ( \3613 , \2941 );
nand \U$3271 ( \3614 , \3613 , RIbb2e800_31);
nand \U$3272 ( \3615 , \3612 , \3614 );
not \U$3273 ( \3616 , \1147 );
not \U$3274 ( \3617 , RIbb2f430_5);
not \U$3275 ( \3618 , \3143 );
or \U$3276 ( \3619 , \3617 , \3618 );
buf \U$3277 ( \3620 , \3146 );
nand \U$3278 ( \3621 , \3620 , \1980 );
nand \U$3279 ( \3622 , \3619 , \3621 );
not \U$3280 ( \3623 , \3622 );
or \U$3281 ( \3624 , \3616 , \3623 );
nand \U$3282 ( \3625 , \3207 , \1090 );
nand \U$3283 ( \3626 , \3624 , \3625 );
xor \U$3284 ( \3627 , \3615 , \3626 );
not \U$3285 ( \3628 , \1294 );
not \U$3286 ( \3629 , \1246 );
not \U$3287 ( \3630 , \3226 );
or \U$3288 ( \3631 , \3629 , \3630 );
not \U$3289 ( \3632 , \3226 );
nand \U$3290 ( \3633 , \3632 , \1245 );
nand \U$3291 ( \3634 , \3631 , \3633 );
not \U$3292 ( \3635 , \3634 );
or \U$3293 ( \3636 , \3628 , \3635 );
not \U$3294 ( \3637 , \1246 );
nor \U$3295 ( \3638 , \3006 , \383 );
not \U$3296 ( \3639 , \3638 );
not \U$3297 ( \3640 , \866 );
or \U$3298 ( \3641 , \3639 , \3640 );
and \U$3299 ( \3642 , \3184 , \3014 );
not \U$3300 ( \3643 , \690 );
nor \U$3301 ( \3644 , \3642 , \3643 );
nand \U$3302 ( \3645 , \3641 , \3644 );
not \U$3303 ( \3646 , \692 );
nor \U$3304 ( \3647 , \3646 , \382 );
and \U$3305 ( \3648 , \3645 , \3647 );
not \U$3306 ( \3649 , \3645 );
not \U$3307 ( \3650 , \3647 );
and \U$3308 ( \3651 , \3649 , \3650 );
nor \U$3309 ( \3652 , \3648 , \3651 );
buf \U$3310 ( \3653 , \3652 );
buf \U$3311 ( \3654 , \3653 );
not \U$3312 ( \3655 , \3654 );
not \U$3313 ( \3656 , \3655 );
or \U$3314 ( \3657 , \3637 , \3656 );
nand \U$3315 ( \3658 , \3654 , \1245 );
nand \U$3316 ( \3659 , \3657 , \3658 );
nand \U$3317 ( \3660 , \3659 , \1265 );
nand \U$3318 ( \3661 , \3636 , \3660 );
xor \U$3319 ( \3662 , \3627 , \3661 );
xor \U$3320 ( \3663 , \3603 , \3662 );
xor \U$3321 ( \3664 , \3409 , \3415 );
xor \U$3322 ( \3665 , \3664 , \3432 );
and \U$3323 ( \3666 , \3663 , \3665 );
and \U$3324 ( \3667 , \3603 , \3662 );
or \U$3325 ( \3668 , \3666 , \3667 );
xor \U$3326 ( \3669 , \3601 , \3668 );
and \U$3327 ( \3670 , \1393 , \3046 );
not \U$3328 ( \3671 , \3465 );
not \U$3329 ( \3672 , RIbb2e9e0_27);
not \U$3330 ( \3673 , \894 );
or \U$3331 ( \3674 , \3672 , \3673 );
nand \U$3332 ( \3675 , \893 , \3454 );
nand \U$3333 ( \3676 , \3674 , \3675 );
not \U$3334 ( \3677 , \3676 );
or \U$3335 ( \3678 , \3671 , \3677 );
nand \U$3336 ( \3679 , \3464 , \3445 );
nand \U$3337 ( \3680 , \3678 , \3679 );
xor \U$3338 ( \3681 , \3670 , \3680 );
not \U$3339 ( \3682 , \3383 );
not \U$3340 ( \3683 , RIbb2ebc0_23);
not \U$3341 ( \3684 , \953 );
or \U$3342 ( \3685 , \3683 , \3684 );
nand \U$3343 ( \3686 , \957 , \3388 );
nand \U$3344 ( \3687 , \3685 , \3686 );
not \U$3345 ( \3688 , \3687 );
or \U$3346 ( \3689 , \3682 , \3688 );
nand \U$3347 ( \3690 , \3390 , \3407 );
nand \U$3348 ( \3691 , \3689 , \3690 );
xor \U$3349 ( \3692 , \3681 , \3691 );
not \U$3350 ( \3693 , \832 );
not \U$3351 ( \3694 , \3059 );
or \U$3352 ( \3695 , \3693 , \3694 );
not \U$3353 ( \3696 , RIbb2ee90_17);
not \U$3354 ( \3697 , \1644 );
or \U$3355 ( \3698 , \3696 , \3697 );
not \U$3356 ( \3699 , RIbb2ee90_17);
nand \U$3357 ( \3700 , \1643 , \3699 );
nand \U$3358 ( \3701 , \3698 , \3700 );
nand \U$3359 ( \3702 , \3701 , \836 );
nand \U$3360 ( \3703 , \3695 , \3702 );
not \U$3361 ( \3704 , \1294 );
not \U$3362 ( \3705 , \1290 );
not \U$3363 ( \3706 , \3203 );
or \U$3364 ( \3707 , \3705 , \3706 );
nand \U$3365 ( \3708 , \3202 , \1289 );
nand \U$3366 ( \3709 , \3707 , \3708 );
not \U$3367 ( \3710 , \3709 );
or \U$3368 ( \3711 , \3704 , \3710 );
nand \U$3369 ( \3712 , \3634 , \1265 );
nand \U$3370 ( \3713 , \3711 , \3712 );
xor \U$3371 ( \3714 , \3703 , \3713 );
not \U$3372 ( \3715 , \1376 );
xor \U$3373 ( \3716 , \1313 , \3654 );
not \U$3374 ( \3717 , \3716 );
or \U$3375 ( \3718 , \3715 , \3717 );
nand \U$3376 ( \3719 , \3025 , \1430 );
nand \U$3377 ( \3720 , \3718 , \3719 );
xor \U$3378 ( \3721 , \3714 , \3720 );
xor \U$3379 ( \3722 , \3692 , \3721 );
not \U$3380 ( \3723 , \2078 );
not \U$3381 ( \3724 , RIbb2ecb0_21);
not \U$3382 ( \3725 , \1039 );
or \U$3383 ( \3726 , \3724 , \3725 );
nand \U$3384 ( \3727 , \1563 , \2254 );
nand \U$3385 ( \3728 , \3726 , \3727 );
not \U$3386 ( \3729 , \3728 );
or \U$3387 ( \3730 , \3723 , \3729 );
nand \U$3388 ( \3731 , \3474 , \2077 );
nand \U$3389 ( \3732 , \3730 , \3731 );
not \U$3390 ( \3733 , \916 );
not \U$3391 ( \3734 , \3423 );
or \U$3392 ( \3735 , \3733 , \3734 );
not \U$3393 ( \3736 , \1170 );
and \U$3394 ( \3737 , \3736 , \1656 );
not \U$3395 ( \3738 , \3736 );
and \U$3396 ( \3739 , \3738 , RIbb2f070_13);
or \U$3397 ( \3740 , \3737 , \3739 );
nand \U$3398 ( \3741 , \3740 , \998 );
nand \U$3399 ( \3742 , \3735 , \3741 );
xor \U$3400 ( \3743 , \3732 , \3742 );
not \U$3401 ( \3744 , \1445 );
not \U$3402 ( \3745 , \3413 );
or \U$3403 ( \3746 , \3744 , \3745 );
not \U$3404 ( \3747 , \3067 );
not \U$3405 ( \3748 , \2356 );
and \U$3406 ( \3749 , \3747 , \3748 );
and \U$3407 ( \3750 , \1114 , \2356 );
nor \U$3408 ( \3751 , \3749 , \3750 );
not \U$3409 ( \3752 , \3751 );
nand \U$3410 ( \3753 , \3752 , \1517 );
nand \U$3411 ( \3754 , \3746 , \3753 );
xor \U$3412 ( \3755 , \3743 , \3754 );
xor \U$3413 ( \3756 , \3722 , \3755 );
xor \U$3414 ( \3757 , \3669 , \3756 );
not \U$3415 ( \3758 , \1090 );
not \U$3416 ( \3759 , RIbb2f430_5);
not \U$3417 ( \3760 , \3655 );
or \U$3418 ( \3761 , \3759 , \3760 );
buf \U$3419 ( \3762 , \3653 );
nand \U$3420 ( \3763 , \3762 , \1980 );
nand \U$3421 ( \3764 , \3761 , \3763 );
not \U$3422 ( \3765 , \3764 );
or \U$3423 ( \3766 , \3758 , \3765 );
nand \U$3424 ( \3767 , \3230 , \1147 );
nand \U$3425 ( \3768 , \3766 , \3767 );
not \U$3426 ( \3769 , \2078 );
not \U$3427 ( \3770 , \3554 );
or \U$3428 ( \3771 , \3769 , \3770 );
not \U$3429 ( \3772 , RIbb2ecb0_21);
buf \U$3430 ( \3773 , \3242 );
not \U$3431 ( \3774 , \3773 );
or \U$3432 ( \3775 , \3772 , \3774 );
nand \U$3433 ( \3776 , \1643 , \849 );
nand \U$3434 ( \3777 , \3775 , \3776 );
nand \U$3435 ( \3778 , \3777 , \2077 );
nand \U$3436 ( \3779 , \3771 , \3778 );
xor \U$3437 ( \3780 , \3768 , \3779 );
not \U$3438 ( \3781 , \1737 );
not \U$3439 ( \3782 , \3148 );
or \U$3440 ( \3783 , \3781 , \3782 );
not \U$3441 ( \3784 , RIbb2f340_7);
not \U$3442 ( \3785 , \3203 );
or \U$3443 ( \3786 , \3784 , \3785 );
nand \U$3444 ( \3787 , \3202 , \1692 );
nand \U$3445 ( \3788 , \3786 , \3787 );
nand \U$3446 ( \3789 , \3788 , \1702 );
nand \U$3447 ( \3790 , \3783 , \3789 );
and \U$3448 ( \3791 , \3780 , \3790 );
and \U$3449 ( \3792 , \3768 , \3779 );
or \U$3450 ( \3793 , \3791 , \3792 );
not \U$3451 ( \3794 , \2925 );
not \U$3452 ( \3795 , \3267 );
or \U$3453 ( \3796 , \3794 , \3795 );
not \U$3454 ( \3797 , RIbb2e8f0_29);
not \U$3455 ( \3798 , \3452 );
or \U$3456 ( \3799 , \3797 , \3798 );
not \U$3457 ( \3800 , RIbb2e8f0_29);
nand \U$3458 ( \3801 , \1476 , \3800 );
nand \U$3459 ( \3802 , \3799 , \3801 );
nand \U$3460 ( \3803 , \3802 , \2922 );
nand \U$3461 ( \3804 , \3796 , \3803 );
not \U$3462 ( \3805 , \916 );
not \U$3463 ( \3806 , RIbb2f070_13);
not \U$3464 ( \3807 , \1851 );
not \U$3465 ( \3808 , \3807 );
or \U$3466 ( \3809 , \3806 , \3808 );
not \U$3467 ( \3810 , \3807 );
nand \U$3468 ( \3811 , \3810 , \906 );
nand \U$3469 ( \3812 , \3809 , \3811 );
not \U$3470 ( \3813 , \3812 );
or \U$3471 ( \3814 , \3805 , \3813 );
nand \U$3472 ( \3815 , \3579 , \998 );
nand \U$3473 ( \3816 , \3814 , \3815 );
xor \U$3474 ( \3817 , \3804 , \3816 );
not \U$3475 ( \3818 , \1517 );
not \U$3476 ( \3819 , \3119 );
or \U$3477 ( \3820 , \3818 , \3819 );
buf \U$3478 ( \3821 , \1419 );
not \U$3479 ( \3822 , \3821 );
and \U$3480 ( \3823 , RIbb2ef80_15, \3822 );
not \U$3481 ( \3824 , RIbb2ef80_15);
and \U$3482 ( \3825 , \3824 , \3821 );
or \U$3483 ( \3826 , \3823 , \3825 );
nand \U$3484 ( \3827 , \3826 , \1445 );
nand \U$3485 ( \3828 , \3820 , \3827 );
and \U$3486 ( \3829 , \3817 , \3828 );
and \U$3487 ( \3830 , \3804 , \3816 );
or \U$3488 ( \3831 , \3829 , \3830 );
xor \U$3489 ( \3832 , \3793 , \3831 );
xor \U$3490 ( \3833 , \3271 , \3284 );
xor \U$3491 ( \3834 , \3833 , \3297 );
and \U$3492 ( \3835 , \3832 , \3834 );
and \U$3493 ( \3836 , \3793 , \3831 );
or \U$3494 ( \3837 , \3835 , \3836 );
not \U$3495 ( \3838 , \3837 );
not \U$3496 ( \3839 , \3838 );
not \U$3497 ( \3840 , \3839 );
xor \U$3498 ( \3841 , \3603 , \3662 );
xor \U$3499 ( \3842 , \3841 , \3665 );
not \U$3500 ( \3843 , \3842 );
or \U$3501 ( \3844 , \3840 , \3843 );
or \U$3502 ( \3845 , \3839 , \3842 );
xor \U$3503 ( \3846 , \3093 , \3103 );
xor \U$3504 ( \3847 , \3846 , \3121 );
xor \U$3505 ( \3848 , \3570 , \3581 );
xor \U$3506 ( \3849 , \3848 , \3592 );
xor \U$3507 ( \3850 , \3847 , \3849 );
xor \U$3508 ( \3851 , \3174 , \3255 );
xor \U$3509 ( \3852 , \3851 , \3232 );
and \U$3510 ( \3853 , \3850 , \3852 );
and \U$3511 ( \3854 , \3847 , \3849 );
or \U$3512 ( \3855 , \3853 , \3854 );
nand \U$3513 ( \3856 , \3845 , \3855 );
nand \U$3514 ( \3857 , \3844 , \3856 );
not \U$3515 ( \3858 , \3857 );
and \U$3516 ( \3859 , \3757 , \3858 );
not \U$3517 ( \3860 , \3757 );
and \U$3518 ( \3861 , \3860 , \3857 );
nor \U$3519 ( \3862 , \3859 , \3861 );
xnor \U$3520 ( \3863 , \3513 , \3862 );
not \U$3521 ( \3864 , RIbb2e710_33);
not \U$3522 ( \3865 , \3864 );
not \U$3523 ( \3866 , RIbb2e620_35);
and \U$3524 ( \3867 , RIbb2e698_34, \3866 );
not \U$3525 ( \3868 , RIbb2e698_34);
and \U$3526 ( \3869 , \3868 , RIbb2e620_35);
nor \U$3527 ( \3870 , \3867 , \3869 );
buf \U$3528 ( \3871 , \3870 );
not \U$3529 ( \3872 , \3871 );
and \U$3530 ( \3873 , \3865 , \3872 );
not \U$3531 ( \3874 , RIbb2e710_33);
not \U$3532 ( \3875 , \813 );
or \U$3533 ( \3876 , \3874 , \3875 );
not \U$3534 ( \3877 , RIbb2e710_33);
nand \U$3535 ( \3878 , \2251 , \3877 );
nand \U$3536 ( \3879 , \3876 , \3878 );
and \U$3537 ( \3880 , RIbb2e698_34, RIbb2e710_33);
not \U$3538 ( \3881 , RIbb2e698_34);
not \U$3539 ( \3882 , RIbb2e710_33);
and \U$3540 ( \3883 , \3881 , \3882 );
nor \U$3541 ( \3884 , \3880 , \3883 );
and \U$3542 ( \3885 , \3870 , \3884 );
buf \U$3543 ( \3886 , \3885 );
buf \U$3544 ( \3887 , \3886 );
and \U$3545 ( \3888 , \3879 , \3887 );
nor \U$3546 ( \3889 , \3873 , \3888 );
not \U$3547 ( \3890 , \1147 );
not \U$3548 ( \3891 , \3764 );
or \U$3549 ( \3892 , \3890 , \3891 );
not \U$3550 ( \3893 , RIbb2f430_5);
not \U$3551 ( \3894 , \3023 );
or \U$3552 ( \3895 , \3893 , \3894 );
nand \U$3553 ( \3896 , \3022 , \1647 );
nand \U$3554 ( \3897 , \3895 , \3896 );
nand \U$3555 ( \3898 , \3897 , \1090 );
nand \U$3556 ( \3899 , \3892 , \3898 );
xor \U$3557 ( \3900 , \3889 , \3899 );
not \U$3558 ( \3901 , \1737 );
not \U$3559 ( \3902 , \3788 );
or \U$3560 ( \3903 , \3901 , \3902 );
not \U$3561 ( \3904 , RIbb2f340_7);
not \U$3562 ( \3905 , \3228 );
not \U$3563 ( \3906 , \3905 );
or \U$3564 ( \3907 , \3904 , \3906 );
nand \U$3565 ( \3908 , \3228 , \1692 );
nand \U$3566 ( \3909 , \3907 , \3908 );
nand \U$3567 ( \3910 , \3909 , \1702 );
nand \U$3568 ( \3911 , \3903 , \3910 );
and \U$3569 ( \3912 , \3900 , \3911 );
and \U$3570 ( \3913 , \3889 , \3899 );
or \U$3571 ( \3914 , \3912 , \3913 );
xor \U$3572 ( \3915 , \3804 , \3816 );
xor \U$3573 ( \3916 , \3915 , \3828 );
xor \U$3574 ( \3917 , \3914 , \3916 );
xor \U$3575 ( \3918 , \3768 , \3779 );
xor \U$3576 ( \3919 , \3918 , \3790 );
and \U$3577 ( \3920 , \3917 , \3919 );
and \U$3578 ( \3921 , \3914 , \3916 );
or \U$3579 ( \3922 , \3920 , \3921 );
not \U$3580 ( \3923 , \1077 );
not \U$3581 ( \3924 , RIbb2f160_11);
not \U$3582 ( \3925 , \2224 );
or \U$3583 ( \3926 , \3924 , \3925 );
nand \U$3584 ( \3927 , \3320 , \1805 );
nand \U$3585 ( \3928 , \3926 , \3927 );
not \U$3586 ( \3929 , \3928 );
or \U$3587 ( \3930 , \3923 , \3929 );
not \U$3588 ( \3931 , RIbb2f160_11);
not \U$3589 ( \3932 , \3342 );
or \U$3590 ( \3933 , \3931 , \3932 );
nand \U$3591 ( \3934 , \3343 , \1805 );
nand \U$3592 ( \3935 , \3933 , \3934 );
nand \U$3593 ( \3936 , \3935 , \1011 );
nand \U$3594 ( \3937 , \3930 , \3936 );
not \U$3595 ( \3938 , \2077 );
not \U$3596 ( \3939 , RIbb2ecb0_21);
not \U$3597 ( \3940 , \3054 );
or \U$3598 ( \3941 , \3939 , \3940 );
nand \U$3599 ( \3942 , \1138 , \2067 );
nand \U$3600 ( \3943 , \3941 , \3942 );
not \U$3601 ( \3944 , \3943 );
or \U$3602 ( \3945 , \3938 , \3944 );
nand \U$3603 ( \3946 , \3777 , \2078 );
nand \U$3604 ( \3947 , \3945 , \3946 );
xor \U$3605 ( \3948 , \3937 , \3947 );
not \U$3606 ( \3949 , \1570 );
not \U$3607 ( \3950 , RIbb2f250_9);
buf \U$3608 ( \3951 , \3166 );
not \U$3609 ( \3952 , \3951 );
not \U$3610 ( \3953 , \3952 );
or \U$3611 ( \3954 , \3950 , \3953 );
nand \U$3612 ( \3955 , \3167 , \1566 );
nand \U$3613 ( \3956 , \3954 , \3955 );
not \U$3614 ( \3957 , \3956 );
or \U$3615 ( \3958 , \3949 , \3957 );
not \U$3616 ( \3959 , RIbb2f250_9);
not \U$3617 ( \3960 , \3143 );
or \U$3618 ( \3961 , \3959 , \3960 );
nand \U$3619 ( \3962 , \3620 , \1554 );
nand \U$3620 ( \3963 , \3961 , \3962 );
nand \U$3621 ( \3964 , \3963 , \1533 );
nand \U$3622 ( \3965 , \3958 , \3964 );
and \U$3623 ( \3966 , \3948 , \3965 );
and \U$3624 ( \3967 , \3937 , \3947 );
or \U$3625 ( \3968 , \3966 , \3967 );
not \U$3626 ( \3969 , \2980 );
and \U$3627 ( \3970 , RIbb2ead0_25, \1562 );
not \U$3628 ( \3971 , RIbb2ead0_25);
and \U$3629 ( \3972 , \3971 , \1038 );
or \U$3630 ( \3973 , \3970 , \3972 );
not \U$3631 ( \3974 , \3973 );
or \U$3632 ( \3975 , \3969 , \3974 );
nand \U$3633 ( \3976 , \3101 , \2963 );
nand \U$3634 ( \3977 , \3975 , \3976 );
not \U$3635 ( \3978 , \3465 );
not \U$3636 ( \3979 , \3536 );
or \U$3637 ( \3980 , \3978 , \3979 );
buf \U$3638 ( \3981 , \951 );
and \U$3639 ( \3982 , \3981 , RIbb2e9e0_27);
not \U$3640 ( \3983 , \3981 );
and \U$3641 ( \3984 , \3983 , \3454 );
or \U$3642 ( \3985 , \3982 , \3984 );
nand \U$3643 ( \3986 , \3985 , \3445 );
nand \U$3644 ( \3987 , \3980 , \3986 );
xor \U$3645 ( \3988 , \3977 , \3987 );
not \U$3646 ( \3989 , \832 );
not \U$3647 ( \3990 , \1169 );
buf \U$3648 ( \3991 , \3990 );
and \U$3649 ( \3992 , \3991 , RIbb2ee90_17);
not \U$3650 ( \3993 , \3991 );
and \U$3651 ( \3994 , \3993 , \3057 );
or \U$3652 ( \3995 , \3992 , \3994 );
not \U$3653 ( \3996 , \3995 );
or \U$3654 ( \3997 , \3989 , \3996 );
nand \U$3655 ( \3998 , \3293 , \836 );
nand \U$3656 ( \3999 , \3997 , \3998 );
xor \U$3657 ( \4000 , \3988 , \3999 );
xor \U$3658 ( \4001 , \3968 , \4000 );
not \U$3659 ( \4002 , \853 );
not \U$3660 ( \4003 , RIbb2eda0_19);
not \U$3661 ( \4004 , \1113 );
or \U$3662 ( \4005 , \4003 , \4004 );
not \U$3663 ( \4006 , \3065 );
nand \U$3664 ( \4007 , \4006 , \1776 );
nand \U$3665 ( \4008 , \4005 , \4007 );
not \U$3666 ( \4009 , \4008 );
or \U$3667 ( \4010 , \4002 , \4009 );
nand \U$3668 ( \4011 , \3253 , \855 );
nand \U$3669 ( \4012 , \4010 , \4011 );
not \U$3670 ( \4013 , \1294 );
not \U$3671 ( \4014 , \1246 );
not \U$3672 ( \4015 , \3022 );
not \U$3673 ( \4016 , \4015 );
not \U$3674 ( \4017 , \4016 );
not \U$3675 ( \4018 , \4017 );
or \U$3676 ( \4019 , \4014 , \4018 );
buf \U$3677 ( \4020 , \3020 );
not \U$3678 ( \4021 , \4020 );
not \U$3679 ( \4022 , \4021 );
nand \U$3680 ( \4023 , \4022 , \1245 );
nand \U$3681 ( \4024 , \4019 , \4023 );
not \U$3682 ( \4025 , \4024 );
or \U$3683 ( \4026 , \4013 , \4025 );
not \U$3684 ( \4027 , \1246 );
not \U$3685 ( \4028 , \3044 );
buf \U$3686 ( \4029 , \4028 );
not \U$3687 ( \4030 , \4029 );
not \U$3688 ( \4031 , \4030 );
not \U$3689 ( \4032 , \4031 );
or \U$3690 ( \4033 , \4027 , \4032 );
nand \U$3691 ( \4034 , \4030 , \1289 );
nand \U$3692 ( \4035 , \4033 , \4034 );
nand \U$3693 ( \4036 , \1265 , \4035 );
nand \U$3694 ( \4037 , \4026 , \4036 );
xor \U$3695 ( \4038 , \4012 , \4037 );
not \U$3696 ( \4039 , \1430 );
not \U$3697 ( \4040 , \3092 );
and \U$3698 ( \4041 , \1394 , \4040 );
not \U$3699 ( \4042 , \1394 );
and \U$3700 ( \4043 , \4042 , \3092 );
or \U$3701 ( \4044 , \4041 , \4043 );
not \U$3702 ( \4045 , \4044 );
or \U$3703 ( \4046 , \4039 , \4045 );
nand \U$3704 ( \4047 , \3280 , \1376 );
nand \U$3705 ( \4048 , \4046 , \4047 );
xor \U$3706 ( \4049 , \4038 , \4048 );
and \U$3707 ( \4050 , \4001 , \4049 );
and \U$3708 ( \4051 , \3968 , \4000 );
or \U$3709 ( \4052 , \4050 , \4051 );
xor \U$3710 ( \4053 , \3922 , \4052 );
xor \U$3711 ( \4054 , \3847 , \3849 );
xor \U$3712 ( \4055 , \4054 , \3852 );
and \U$3713 ( \4056 , \4053 , \4055 );
and \U$3714 ( \4057 , \3922 , \4052 );
or \U$3715 ( \4058 , \4056 , \4057 );
not \U$3716 ( \4059 , \4058 );
not \U$3717 ( \4060 , \4059 );
not \U$3718 ( \4061 , \3838 );
not \U$3719 ( \4062 , \3855 );
or \U$3720 ( \4063 , \4061 , \4062 );
or \U$3721 ( \4064 , \3855 , \3838 );
nand \U$3722 ( \4065 , \4063 , \4064 );
not \U$3723 ( \4066 , \3842 );
and \U$3724 ( \4067 , \4065 , \4066 );
not \U$3725 ( \4068 , \4065 );
and \U$3726 ( \4069 , \4068 , \3842 );
nor \U$3727 ( \4070 , \4067 , \4069 );
not \U$3728 ( \4071 , \4070 );
or \U$3729 ( \4072 , \4060 , \4071 );
xor \U$3730 ( \4073 , \3558 , \3595 );
xor \U$3731 ( \4074 , \4073 , \3598 );
not \U$3732 ( \4075 , \3871 );
or \U$3733 ( \4076 , \3887 , \4075 );
nand \U$3734 ( \4077 , \4076 , RIbb2e710_33);
nand \U$3735 ( \4078 , \3076 , \3080 );
not \U$3736 ( \4079 , \4078 );
not \U$3737 ( \4080 , \4079 );
not \U$3738 ( \4081 , \666 );
or \U$3739 ( \4082 , \4080 , \4081 );
nand \U$3740 ( \4083 , \867 , \4078 );
nand \U$3741 ( \4084 , \4082 , \4083 );
buf \U$3742 ( \4085 , \4084 );
buf \U$3743 ( \4086 , \4085 );
not \U$3744 ( \4087 , \4086 );
buf \U$3745 ( \4088 , \4087 );
not \U$3746 ( \4089 , \4088 );
and \U$3747 ( \4090 , \4089 , \1313 );
xor \U$3748 ( \4091 , \4077 , \4090 );
not \U$3749 ( \4092 , \2940 );
not \U$3750 ( \4093 , RIbb2e800_31);
not \U$3751 ( \4094 , \2946 );
or \U$3752 ( \4095 , \4093 , \4094 );
not \U$3753 ( \4096 , RIbb2e800_31);
nand \U$3754 ( \4097 , \893 , \4096 );
nand \U$3755 ( \4098 , \4095 , \4097 );
not \U$3756 ( \4099 , \4098 );
or \U$3757 ( \4100 , \4092 , \4099 );
nand \U$3758 ( \4101 , \3610 , \3613 );
nand \U$3759 ( \4102 , \4100 , \4101 );
and \U$3760 ( \4103 , \4091 , \4102 );
and \U$3761 ( \4104 , \4077 , \4090 );
or \U$3762 ( \4105 , \4103 , \4104 );
xor \U$3763 ( \4106 , \3977 , \3987 );
and \U$3764 ( \4107 , \4106 , \3999 );
and \U$3765 ( \4108 , \3977 , \3987 );
or \U$3766 ( \4109 , \4107 , \4108 );
xor \U$3767 ( \4110 , \4105 , \4109 );
xor \U$3768 ( \4111 , \4012 , \4037 );
and \U$3769 ( \4112 , \4111 , \4048 );
and \U$3770 ( \4113 , \4012 , \4037 );
or \U$3771 ( \4114 , \4112 , \4113 );
and \U$3772 ( \4115 , \4110 , \4114 );
and \U$3773 ( \4116 , \4105 , \4109 );
or \U$3774 ( \4117 , \4115 , \4116 );
xor \U$3775 ( \4118 , \4074 , \4117 );
xor \U$3776 ( \4119 , \3124 , \3257 );
xor \U$3777 ( \4120 , \4119 , \3300 );
xor \U$3778 ( \4121 , \4118 , \4120 );
nand \U$3779 ( \4122 , \4072 , \4121 );
not \U$3780 ( \4123 , \4070 );
nand \U$3781 ( \4124 , \4123 , \4058 );
nand \U$3782 ( \4125 , \4122 , \4124 );
not \U$3783 ( \4126 , \4125 );
not \U$3784 ( \4127 , \1294 );
not \U$3785 ( \4128 , \3659 );
or \U$3786 ( \4129 , \4127 , \4128 );
nand \U$3787 ( \4130 , \4024 , \1265 );
nand \U$3788 ( \4131 , \4129 , \4130 );
not \U$3789 ( \4132 , \4131 );
nand \U$3790 ( \4133 , \4132 , \3615 );
not \U$3791 ( \4134 , \4133 );
not \U$3792 ( \4135 , \1077 );
not \U$3793 ( \4136 , \3566 );
or \U$3794 ( \4137 , \4135 , \4136 );
nand \U$3795 ( \4138 , \3928 , \1011 );
nand \U$3796 ( \4139 , \4137 , \4138 );
not \U$3797 ( \4140 , \4139 );
not \U$3798 ( \4141 , \1570 );
not \U$3799 ( \4142 , \3523 );
or \U$3800 ( \4143 , \4141 , \4142 );
nand \U$3801 ( \4144 , \3956 , \1533 );
nand \U$3802 ( \4145 , \4143 , \4144 );
not \U$3803 ( \4146 , \4145 );
or \U$3804 ( \4147 , \4140 , \4146 );
not \U$3805 ( \4148 , \4139 );
not \U$3806 ( \4149 , \4148 );
not \U$3807 ( \4150 , \4145 );
not \U$3808 ( \4151 , \4150 );
or \U$3809 ( \4152 , \4149 , \4151 );
not \U$3810 ( \4153 , \3383 );
not \U$3811 ( \4154 , \3588 );
or \U$3812 ( \4155 , \4153 , \4154 );
not \U$3813 ( \4156 , RIbb2ebc0_23);
not \U$3814 ( \4157 , \3481 );
or \U$3815 ( \4158 , \4156 , \4157 );
nand \U$3816 ( \4159 , \3484 , \3388 );
nand \U$3817 ( \4160 , \4158 , \4159 );
nand \U$3818 ( \4161 , \4160 , \3407 );
nand \U$3819 ( \4162 , \4155 , \4161 );
nand \U$3820 ( \4163 , \4152 , \4162 );
nand \U$3821 ( \4164 , \4147 , \4163 );
not \U$3822 ( \4165 , \4164 );
or \U$3823 ( \4166 , \4134 , \4165 );
not \U$3824 ( \4167 , \3615 );
nand \U$3825 ( \4168 , \4167 , \4131 );
nand \U$3826 ( \4169 , \4166 , \4168 );
not \U$3827 ( \4170 , \4169 );
xor \U$3828 ( \4171 , \3467 , \3488 );
xor \U$3829 ( \4172 , \4171 , \3507 );
not \U$3830 ( \4173 , \4172 );
and \U$3831 ( \4174 , \3377 , \3358 );
not \U$3832 ( \4175 , \3377 );
and \U$3833 ( \4176 , \4175 , \3324 );
or \U$3834 ( \4177 , \4174 , \4176 );
and \U$3835 ( \4178 , \4177 , \3356 );
not \U$3836 ( \4179 , \4177 );
and \U$3837 ( \4180 , \4179 , \3353 );
nor \U$3838 ( \4181 , \4178 , \4180 );
nand \U$3839 ( \4182 , \4173 , \4181 );
not \U$3840 ( \4183 , \4182 );
or \U$3841 ( \4184 , \4170 , \4183 );
or \U$3842 ( \4185 , \4181 , \4173 );
nand \U$3843 ( \4186 , \4184 , \4185 );
xor \U$3844 ( \4187 , \3615 , \3626 );
and \U$3845 ( \4188 , \4187 , \3661 );
and \U$3846 ( \4189 , \3615 , \3626 );
or \U$3847 ( \4190 , \4188 , \4189 );
not \U$3848 ( \4191 , \853 );
not \U$3849 ( \4192 , \3373 );
or \U$3850 ( \4193 , \4191 , \4192 );
not \U$3851 ( \4194 , RIbb2eda0_19);
not \U$3852 ( \4195 , \1731 );
or \U$3853 ( \4196 , \4194 , \4195 );
nand \U$3854 ( \4197 , \1730 , \1776 );
nand \U$3855 ( \4198 , \4196 , \4197 );
nand \U$3856 ( \4199 , \4198 , \855 );
nand \U$3857 ( \4200 , \4193 , \4199 );
not \U$3858 ( \4201 , \1702 );
not \U$3859 ( \4202 , \3349 );
or \U$3860 ( \4203 , \4201 , \4202 );
not \U$3861 ( \4204 , RIbb2f340_7);
not \U$3862 ( \4205 , \2224 );
or \U$3863 ( \4206 , \4204 , \4205 );
nand \U$3864 ( \4207 , \2225 , \1692 );
nand \U$3865 ( \4208 , \4206 , \4207 );
nand \U$3866 ( \4209 , \4208 , \1737 );
nand \U$3867 ( \4210 , \4203 , \4209 );
xor \U$3868 ( \4211 , \4200 , \4210 );
not \U$3869 ( \4212 , \1090 );
not \U$3870 ( \4213 , \3622 );
or \U$3871 ( \4214 , \4212 , \4213 );
not \U$3872 ( \4215 , RIbb2f430_5);
buf \U$3873 ( \4216 , \3952 );
not \U$3874 ( \4217 , \4216 );
or \U$3875 ( \4218 , \4215 , \4217 );
not \U$3876 ( \4219 , \3166 );
not \U$3877 ( \4220 , \4219 );
nand \U$3878 ( \4221 , \4220 , \1085 );
nand \U$3879 ( \4222 , \4218 , \4221 );
nand \U$3880 ( \4223 , \4222 , \1147 );
nand \U$3881 ( \4224 , \4214 , \4223 );
xor \U$3882 ( \4225 , \4211 , \4224 );
xor \U$3883 ( \4226 , \4190 , \4225 );
not \U$3884 ( \4227 , \1077 );
not \U$3885 ( \4228 , RIbb2f160_11);
not \U$3886 ( \4229 , \2052 );
or \U$3887 ( \4230 , \4228 , \4229 );
nand \U$3888 ( \4231 , \1421 , \1048 );
nand \U$3889 ( \4232 , \4230 , \4231 );
not \U$3890 ( \4233 , \4232 );
or \U$3891 ( \4234 , \4227 , \4233 );
nand \U$3892 ( \4235 , \3497 , \1011 );
nand \U$3893 ( \4236 , \4234 , \4235 );
not \U$3894 ( \4237 , \2963 );
and \U$3895 ( \4238 , RIbb2ead0_25, \1475 );
not \U$3896 ( \4239 , RIbb2ead0_25);
and \U$3897 ( \4240 , \4239 , \1476 );
or \U$3898 ( \4241 , \4238 , \4240 );
not \U$3899 ( \4242 , \4241 );
or \U$3900 ( \4243 , \4237 , \4242 );
nand \U$3901 ( \4244 , \2968 , \2980 );
nand \U$3902 ( \4245 , \4243 , \4244 );
xor \U$3903 ( \4246 , \4236 , \4245 );
not \U$3904 ( \4247 , \1533 );
not \U$3905 ( \4248 , \3313 );
or \U$3906 ( \4249 , \4247 , \4248 );
not \U$3907 ( \4250 , RIbb2f250_9);
not \U$3908 ( \4251 , \1854 );
or \U$3909 ( \4252 , \4250 , \4251 );
nand \U$3910 ( \4253 , \3503 , \1566 );
nand \U$3911 ( \4254 , \4252 , \4253 );
nand \U$3912 ( \4255 , \4254 , \1570 );
nand \U$3913 ( \4256 , \4249 , \4255 );
xor \U$3914 ( \4257 , \4246 , \4256 );
xor \U$3915 ( \4258 , \4226 , \4257 );
not \U$3916 ( \4259 , \4258 );
and \U$3917 ( \4260 , \4186 , \4259 );
not \U$3918 ( \4261 , \4186 );
and \U$3919 ( \4262 , \4261 , \4258 );
or \U$3920 ( \4263 , \4260 , \4262 );
not \U$3921 ( \4264 , \4117 );
not \U$3922 ( \4265 , \4120 );
or \U$3923 ( \4266 , \4264 , \4265 );
or \U$3924 ( \4267 , \4120 , \4117 );
nand \U$3925 ( \4268 , \4267 , \4074 );
nand \U$3926 ( \4269 , \4266 , \4268 );
xnor \U$3927 ( \4270 , \4263 , \4269 );
not \U$3928 ( \4271 , \4270 );
not \U$3929 ( \4272 , \1517 );
not \U$3930 ( \4273 , \3826 );
or \U$3931 ( \4274 , \4272 , \4273 );
and \U$3932 ( \4275 , RIbb2ef80_15, \1340 );
not \U$3933 ( \4276 , RIbb2ef80_15);
and \U$3934 ( \4277 , \4276 , \1339 );
or \U$3935 ( \4278 , \4275 , \4277 );
nand \U$3936 ( \4279 , \4278 , \1445 );
nand \U$3937 ( \4280 , \4274 , \4279 );
not \U$3938 ( \4281 , \4280 );
not \U$3939 ( \4282 , \4281 );
not \U$3940 ( \4283 , \3445 );
not \U$3941 ( \4284 , \1886 );
and \U$3942 ( \4285 , \4284 , RIbb2e9e0_27);
not \U$3943 ( \4286 , \4284 );
and \U$3944 ( \4287 , \4286 , \3462 );
or \U$3945 ( \4288 , \4285 , \4287 );
not \U$3946 ( \4289 , \4288 );
or \U$3947 ( \4290 , \4283 , \4289 );
nand \U$3948 ( \4291 , \3985 , \3465 );
nand \U$3949 ( \4292 , \4290 , \4291 );
not \U$3950 ( \4293 , \4292 );
not \U$3951 ( \4294 , \4293 );
or \U$3952 ( \4295 , \4282 , \4294 );
not \U$3953 ( \4296 , \2963 );
not \U$3954 ( \4297 , \3973 );
or \U$3955 ( \4298 , \4296 , \4297 );
not \U$3956 ( \4299 , \1548 );
and \U$3957 ( \4300 , RIbb2ead0_25, \4299 );
not \U$3958 ( \4301 , RIbb2ead0_25);
and \U$3959 ( \4302 , \4301 , \1548 );
or \U$3960 ( \4303 , \4300 , \4302 );
nand \U$3961 ( \4304 , \4303 , \2980 );
nand \U$3962 ( \4305 , \4298 , \4304 );
nand \U$3963 ( \4306 , \4295 , \4305 );
nand \U$3964 ( \4307 , \4280 , \4292 );
nand \U$3965 ( \4308 , \4306 , \4307 );
not \U$3966 ( \4309 , \3613 );
not \U$3967 ( \4310 , \4098 );
or \U$3968 ( \4311 , \4309 , \4310 );
not \U$3969 ( \4312 , RIbb2e800_31);
not \U$3970 ( \4313 , \3262 );
or \U$3971 ( \4314 , \4312 , \4313 );
not \U$3972 ( \4315 , \1509 );
nand \U$3973 ( \4316 , \4315 , \3608 );
nand \U$3974 ( \4317 , \4314 , \4316 );
nand \U$3975 ( \4318 , \4317 , \2940 );
nand \U$3976 ( \4319 , \4311 , \4318 );
not \U$3977 ( \4320 , \1376 );
not \U$3978 ( \4321 , \4044 );
or \U$3979 ( \4322 , \4320 , \4321 );
not \U$3980 ( \4323 , \1394 );
buf \U$3981 ( \4324 , \4084 );
not \U$3982 ( \4325 , \4324 );
not \U$3983 ( \4326 , \4325 );
or \U$3984 ( \4327 , \4323 , \4326 );
nand \U$3985 ( \4328 , \4089 , \1951 );
nand \U$3986 ( \4329 , \4327 , \4328 );
nand \U$3987 ( \4330 , \4329 , \1430 );
nand \U$3988 ( \4331 , \4322 , \4330 );
xor \U$3989 ( \4332 , \4319 , \4331 );
not \U$3990 ( \4333 , \836 );
not \U$3991 ( \4334 , \3995 );
or \U$3992 ( \4335 , \4333 , \4334 );
not \U$3993 ( \4336 , RIbb2ee90_17);
not \U$3994 ( \4337 , \1820 );
or \U$3995 ( \4338 , \4336 , \4337 );
not \U$3996 ( \4339 , \1384 );
not \U$3997 ( \4340 , \4339 );
not \U$3998 ( \4341 , \4340 );
not \U$3999 ( \4342 , \4341 );
nand \U$4000 ( \4343 , \4342 , \859 );
nand \U$4001 ( \4344 , \4338 , \4343 );
nand \U$4002 ( \4345 , \4344 , \832 );
nand \U$4003 ( \4346 , \4335 , \4345 );
and \U$4004 ( \4347 , \4332 , \4346 );
and \U$4005 ( \4348 , \4319 , \4331 );
or \U$4006 ( \4349 , \4347 , \4348 );
or \U$4007 ( \4350 , \4308 , \4349 );
not \U$4008 ( \4351 , \525 );
and \U$4009 ( \4352 , \530 , \4351 );
nand \U$4010 ( \4353 , \524 , \4352 );
buf \U$4011 ( \4354 , \514 );
not \U$4012 ( \4355 , \4354 );
nor \U$4013 ( \4356 , \4353 , \4355 );
not \U$4014 ( \4357 , \4356 );
buf \U$4015 ( \4358 , \592 );
not \U$4016 ( \4359 , \570 );
nand \U$4017 ( \4360 , \4358 , \491 , \454 , \4359 );
buf \U$4018 ( \4361 , \4360 );
not \U$4019 ( \4362 , \4361 );
or \U$4020 ( \4363 , \4357 , \4362 );
buf \U$4021 ( \4364 , \548 );
not \U$4022 ( \4365 , \4364 );
buf \U$4023 ( \4366 , \608 );
nand \U$4024 ( \4367 , \4365 , \4366 );
not \U$4025 ( \4368 , \662 );
nand \U$4026 ( \4369 , \4367 , \4368 );
buf \U$4027 ( \4370 , \4369 );
not \U$4028 ( \4371 , \4353 );
and \U$4029 ( \4372 , \4370 , \4371 );
not \U$4030 ( \4373 , \4352 );
buf \U$4031 ( \4374 , \629 );
not \U$4032 ( \4375 , \4374 );
or \U$4033 ( \4376 , \4373 , \4375 );
and \U$4034 ( \4377 , \636 , \4351 );
not \U$4035 ( \4378 , \638 );
nor \U$4036 ( \4379 , \4377 , \4378 );
nand \U$4037 ( \4380 , \4376 , \4379 );
nor \U$4038 ( \4381 , \4372 , \4380 );
nand \U$4039 ( \4382 , \4363 , \4381 );
not \U$4040 ( \4383 , \640 );
nor \U$4041 ( \4384 , \4383 , \526 );
and \U$4042 ( \4385 , \4382 , \4384 );
not \U$4043 ( \4386 , \4382 );
not \U$4044 ( \4387 , \4384 );
and \U$4045 ( \4388 , \4386 , \4387 );
nor \U$4046 ( \4389 , \4385 , \4388 );
buf \U$4047 ( \4390 , \4389 );
buf \U$4048 ( \4391 , \4390 );
not \U$4049 ( \4392 , \4391 );
buf \U$4050 ( \4393 , \4392 );
not \U$4051 ( \4394 , \4393 );
and \U$4052 ( \4395 , \4394 , \1313 );
not \U$4053 ( \4396 , \853 );
not \U$4054 ( \4397 , RIbb2eda0_19);
not \U$4055 ( \4398 , \1284 );
or \U$4056 ( \4399 , \4397 , \4398 );
nand \U$4057 ( \4400 , \1283 , \1776 );
nand \U$4058 ( \4401 , \4399 , \4400 );
not \U$4059 ( \4402 , \4401 );
or \U$4060 ( \4403 , \4396 , \4402 );
nand \U$4061 ( \4404 , \4008 , \855 );
nand \U$4062 ( \4405 , \4403 , \4404 );
xor \U$4063 ( \4406 , \4395 , \4405 );
not \U$4064 ( \4407 , \1294 );
not \U$4065 ( \4408 , \4035 );
or \U$4066 ( \4409 , \4407 , \4408 );
not \U$4067 ( \4410 , \1246 );
not \U$4068 ( \4411 , \3003 );
not \U$4069 ( \4412 , \4411 );
or \U$4070 ( \4413 , \4410 , \4412 );
nand \U$4071 ( \4414 , \3003 , \1245 );
nand \U$4072 ( \4415 , \4413 , \4414 );
nand \U$4073 ( \4416 , \4415 , \1265 );
nand \U$4074 ( \4417 , \4409 , \4416 );
and \U$4075 ( \4418 , \4406 , \4417 );
and \U$4076 ( \4419 , \4395 , \4405 );
or \U$4077 ( \4420 , \4418 , \4419 );
nand \U$4078 ( \4421 , \4350 , \4420 );
nand \U$4079 ( \4422 , \4308 , \4349 );
nand \U$4080 ( \4423 , \4421 , \4422 );
xor \U$4081 ( \4424 , \4105 , \4109 );
xor \U$4082 ( \4425 , \4424 , \4114 );
xor \U$4083 ( \4426 , \4423 , \4425 );
xor \U$4084 ( \4427 , \3793 , \3831 );
xor \U$4085 ( \4428 , \4427 , \3834 );
and \U$4086 ( \4429 , \4426 , \4428 );
and \U$4087 ( \4430 , \4423 , \4425 );
or \U$4088 ( \4431 , \4429 , \4430 );
not \U$4089 ( \4432 , \4431 );
xor \U$4090 ( \4433 , \4131 , \3615 );
xor \U$4091 ( \4434 , \4164 , \4433 );
not \U$4092 ( \4435 , \4434 );
xor \U$4093 ( \4436 , \3556 , \3543 );
not \U$4094 ( \4437 , \3541 );
xor \U$4095 ( \4438 , \4436 , \4437 );
not \U$4096 ( \4439 , \4438 );
or \U$4097 ( \4440 , \4435 , \4439 );
not \U$4098 ( \4441 , \3889 );
xor \U$4099 ( \4442 , \4077 , \4090 );
xor \U$4100 ( \4443 , \4442 , \4102 );
xor \U$4101 ( \4444 , \4441 , \4443 );
not \U$4102 ( \4445 , \916 );
not \U$4103 ( \4446 , RIbb2f070_13);
not \U$4104 ( \4447 , \3310 );
or \U$4105 ( \4448 , \4446 , \4447 );
not \U$4106 ( \4449 , \3309 );
not \U$4107 ( \4450 , \4449 );
nand \U$4108 ( \4451 , \4450 , \1656 );
nand \U$4109 ( \4452 , \4448 , \4451 );
not \U$4110 ( \4453 , \4452 );
or \U$4111 ( \4454 , \4445 , \4453 );
nand \U$4112 ( \4455 , \3812 , \998 );
nand \U$4113 ( \4456 , \4454 , \4455 );
not \U$4114 ( \4457 , \4456 );
not \U$4115 ( \4458 , \3802 );
not \U$4116 ( \4459 , \4458 );
not \U$4117 ( \4460 , \2925 );
not \U$4118 ( \4461 , \4460 );
and \U$4119 ( \4462 , \4459 , \4461 );
not \U$4120 ( \4463 , RIbb2e8f0_29);
not \U$4121 ( \4464 , \992 );
or \U$4122 ( \4465 , \4463 , \4464 );
nand \U$4123 ( \4466 , \994 , \3800 );
nand \U$4124 ( \4467 , \4465 , \4466 );
and \U$4125 ( \4468 , \4467 , \2922 );
nor \U$4126 ( \4469 , \4462 , \4468 );
not \U$4127 ( \4470 , \4469 );
not \U$4128 ( \4471 , \4470 );
or \U$4129 ( \4472 , \4457 , \4471 );
not \U$4130 ( \4473 , \4456 );
not \U$4131 ( \4474 , \4473 );
not \U$4132 ( \4475 , \4469 );
or \U$4133 ( \4476 , \4474 , \4475 );
not \U$4134 ( \4477 , \3407 );
not \U$4135 ( \4478 , RIbb2ebc0_23);
not \U$4136 ( \4479 , \3365 );
or \U$4137 ( \4480 , \4478 , \4479 );
nand \U$4138 ( \4481 , \3364 , \3401 );
nand \U$4139 ( \4482 , \4480 , \4481 );
not \U$4140 ( \4483 , \4482 );
or \U$4141 ( \4484 , \4477 , \4483 );
nand \U$4142 ( \4485 , \4160 , \3383 );
nand \U$4143 ( \4486 , \4484 , \4485 );
nand \U$4144 ( \4487 , \4476 , \4486 );
nand \U$4145 ( \4488 , \4472 , \4487 );
and \U$4146 ( \4489 , \4444 , \4488 );
and \U$4147 ( \4490 , \4441 , \4443 );
or \U$4148 ( \4491 , \4489 , \4490 );
nand \U$4149 ( \4492 , \4440 , \4491 );
not \U$4150 ( \4493 , \4438 );
not \U$4151 ( \4494 , \4434 );
nand \U$4152 ( \4495 , \4493 , \4494 );
nand \U$4153 ( \4496 , \4492 , \4495 );
not \U$4154 ( \4497 , \4496 );
xor \U$4155 ( \4498 , \4181 , \4172 );
xor \U$4156 ( \4499 , \4498 , \4169 );
nand \U$4157 ( \4500 , \4497 , \4499 );
not \U$4158 ( \4501 , \4500 );
or \U$4159 ( \4502 , \4432 , \4501 );
not \U$4160 ( \4503 , \4499 );
nand \U$4161 ( \4504 , \4503 , \4496 );
nand \U$4162 ( \4505 , \4502 , \4504 );
not \U$4163 ( \4506 , \4505 );
and \U$4164 ( \4507 , \4271 , \4506 );
and \U$4165 ( \4508 , \4270 , \4505 );
nor \U$4166 ( \4509 , \4507 , \4508 );
not \U$4167 ( \4510 , \4509 );
or \U$4168 ( \4511 , \4126 , \4510 );
or \U$4169 ( \4512 , \4125 , \4509 );
nand \U$4170 ( \4513 , \4511 , \4512 );
xor \U$4171 ( \4514 , \3863 , \4513 );
xor \U$4172 ( \4515 , \4496 , \4499 );
xor \U$4173 ( \4516 , \4515 , \4431 );
not \U$4174 ( \4517 , \4516 );
not \U$4175 ( \4518 , \4517 );
xor \U$4176 ( \4519 , \3914 , \3916 );
xor \U$4177 ( \4520 , \4519 , \3919 );
xor \U$4178 ( \4521 , \3889 , \3899 );
xor \U$4179 ( \4522 , \4521 , \3911 );
xor \U$4180 ( \4523 , \4395 , \4405 );
xor \U$4181 ( \4524 , \4523 , \4417 );
xor \U$4182 ( \4525 , \4522 , \4524 );
xor \U$4183 ( \4526 , \4319 , \4331 );
xor \U$4184 ( \4527 , \4526 , \4346 );
and \U$4185 ( \4528 , \4525 , \4527 );
and \U$4186 ( \4529 , \4522 , \4524 );
or \U$4187 ( \4530 , \4528 , \4529 );
or \U$4188 ( \4531 , \4520 , \4530 );
xor \U$4189 ( \4532 , \3968 , \4000 );
xor \U$4190 ( \4533 , \4532 , \4049 );
nand \U$4191 ( \4534 , \4531 , \4533 );
nand \U$4192 ( \4535 , \4520 , \4530 );
nand \U$4193 ( \4536 , \4534 , \4535 );
xor \U$4194 ( \4537 , \4423 , \4425 );
xor \U$4195 ( \4538 , \4537 , \4428 );
xor \U$4196 ( \4539 , \4536 , \4538 );
xor \U$4197 ( \4540 , \3922 , \4052 );
xor \U$4198 ( \4541 , \4540 , \4055 );
and \U$4199 ( \4542 , \4539 , \4541 );
and \U$4200 ( \4543 , \4536 , \4538 );
or \U$4201 ( \4544 , \4542 , \4543 );
not \U$4202 ( \4545 , \4544 );
or \U$4203 ( \4546 , \4518 , \4545 );
or \U$4204 ( \4547 , \4544 , \4517 );
not \U$4205 ( \4548 , \4139 );
not \U$4206 ( \4549 , \4150 );
or \U$4207 ( \4550 , \4548 , \4549 );
or \U$4208 ( \4551 , \4150 , \4139 );
nand \U$4209 ( \4552 , \4550 , \4551 );
xor \U$4210 ( \4553 , \4162 , \4552 );
not \U$4211 ( \4554 , \2940 );
not \U$4212 ( \4555 , RIbb2e800_31);
not \U$4213 ( \4556 , \1475 );
or \U$4214 ( \4557 , \4555 , \4556 );
buf \U$4215 ( \4558 , \1474 );
nand \U$4216 ( \4559 , \4558 , \2917 );
nand \U$4217 ( \4560 , \4557 , \4559 );
not \U$4218 ( \4561 , \4560 );
or \U$4219 ( \4562 , \4554 , \4561 );
nand \U$4220 ( \4563 , \4317 , \2941 );
nand \U$4221 ( \4564 , \4562 , \4563 );
not \U$4222 ( \4565 , \4564 );
not \U$4223 ( \4566 , \998 );
not \U$4224 ( \4567 , \4452 );
or \U$4225 ( \4568 , \4566 , \4567 );
not \U$4226 ( \4569 , RIbb2f070_13);
not \U$4227 ( \4570 , \3319 );
or \U$4228 ( \4571 , \4569 , \4570 );
nand \U$4229 ( \4572 , \2225 , \3421 );
nand \U$4230 ( \4573 , \4571 , \4572 );
nand \U$4231 ( \4574 , \4573 , \916 );
nand \U$4232 ( \4575 , \4568 , \4574 );
not \U$4233 ( \4576 , \4575 );
or \U$4234 ( \4577 , \4565 , \4576 );
or \U$4235 ( \4578 , \4575 , \4564 );
not \U$4236 ( \4579 , \2980 );
not \U$4237 ( \4580 , \3480 );
and \U$4238 ( \4581 , RIbb2ead0_25, \4580 );
not \U$4239 ( \4582 , RIbb2ead0_25);
and \U$4240 ( \4583 , \4582 , \3480 );
or \U$4241 ( \4584 , \4581 , \4583 );
not \U$4242 ( \4585 , \4584 );
or \U$4243 ( \4586 , \4579 , \4585 );
nand \U$4244 ( \4587 , \4303 , \2963 );
nand \U$4245 ( \4588 , \4586 , \4587 );
nand \U$4246 ( \4589 , \4578 , \4588 );
nand \U$4247 ( \4590 , \4577 , \4589 );
not \U$4248 ( \4591 , \3465 );
not \U$4249 ( \4592 , \4288 );
or \U$4250 ( \4593 , \4591 , \4592 );
not \U$4251 ( \4594 , RIbb2e9e0_27);
not \U$4252 ( \4595 , \1038 );
not \U$4253 ( \4596 , \4595 );
or \U$4254 ( \4597 , \4594 , \4596 );
not \U$4255 ( \4598 , RIbb2e9e0_27);
nand \U$4256 ( \4599 , \1561 , \4598 );
nand \U$4257 ( \4600 , \4597 , \4599 );
nand \U$4258 ( \4601 , \4600 , \3445 );
nand \U$4259 ( \4602 , \4593 , \4601 );
not \U$4260 ( \4603 , \4602 );
not \U$4261 ( \4604 , \1517 );
not \U$4262 ( \4605 , \4278 );
or \U$4263 ( \4606 , \4604 , \4605 );
and \U$4264 ( \4607 , RIbb2ef80_15, \1853 );
not \U$4265 ( \4608 , RIbb2ef80_15);
not \U$4266 ( \4609 , \1851 );
not \U$4267 ( \4610 , \4609 );
and \U$4268 ( \4611 , \4608 , \4610 );
or \U$4269 ( \4612 , \4607 , \4611 );
nand \U$4270 ( \4613 , \4612 , \1445 );
nand \U$4271 ( \4614 , \4606 , \4613 );
not \U$4272 ( \4615 , \4614 );
or \U$4273 ( \4616 , \4603 , \4615 );
or \U$4274 ( \4617 , \4614 , \4602 );
not \U$4275 ( \4618 , \836 );
not \U$4276 ( \4619 , \4344 );
or \U$4277 ( \4620 , \4618 , \4619 );
not \U$4278 ( \4621 , RIbb2ee90_17);
not \U$4279 ( \4622 , \1420 );
or \U$4280 ( \4623 , \4621 , \4622 );
nand \U$4281 ( \4624 , \1421 , \859 );
nand \U$4282 ( \4625 , \4623 , \4624 );
nand \U$4283 ( \4626 , \4625 , \832 );
nand \U$4284 ( \4627 , \4620 , \4626 );
nand \U$4285 ( \4628 , \4617 , \4627 );
nand \U$4286 ( \4629 , \4616 , \4628 );
or \U$4287 ( \4630 , \4590 , \4629 );
not \U$4288 ( \4631 , \1570 );
not \U$4289 ( \4632 , \3963 );
or \U$4290 ( \4633 , \4631 , \4632 );
not \U$4291 ( \4634 , RIbb2f250_9);
not \U$4292 ( \4635 , \3203 );
or \U$4293 ( \4636 , \4634 , \4635 );
buf \U$4294 ( \4637 , \3199 );
not \U$4295 ( \4638 , \4637 );
buf \U$4296 ( \4639 , \4638 );
not \U$4297 ( \4640 , \4639 );
nand \U$4298 ( \4641 , \4640 , \1554 );
nand \U$4299 ( \4642 , \4636 , \4641 );
nand \U$4300 ( \4643 , \4642 , \1533 );
nand \U$4301 ( \4644 , \4633 , \4643 );
not \U$4302 ( \4645 , \4644 );
not \U$4303 ( \4646 , \1077 );
not \U$4304 ( \4647 , \3935 );
or \U$4305 ( \4648 , \4646 , \4647 );
not \U$4306 ( \4649 , RIbb2f160_11);
not \U$4307 ( \4650 , \4219 );
or \U$4308 ( \4651 , \4649 , \4650 );
nand \U$4309 ( \4652 , \3951 , \1048 );
nand \U$4310 ( \4653 , \4651 , \4652 );
nand \U$4311 ( \4654 , \4653 , \1011 );
nand \U$4312 ( \4655 , \4648 , \4654 );
not \U$4313 ( \4656 , \4655 );
or \U$4314 ( \4657 , \4645 , \4656 );
or \U$4315 ( \4658 , \4655 , \4644 );
not \U$4316 ( \4659 , \3383 );
not \U$4317 ( \4660 , \4482 );
or \U$4318 ( \4661 , \4659 , \4660 );
not \U$4319 ( \4662 , RIbb2ebc0_23);
not \U$4320 ( \4663 , \3239 );
or \U$4321 ( \4664 , \4662 , \4663 );
nand \U$4322 ( \4665 , \1643 , \3401 );
nand \U$4323 ( \4666 , \4664 , \4665 );
nand \U$4324 ( \4667 , \4666 , \3407 );
nand \U$4325 ( \4668 , \4661 , \4667 );
nand \U$4326 ( \4669 , \4658 , \4668 );
nand \U$4327 ( \4670 , \4657 , \4669 );
nand \U$4328 ( \4671 , \4630 , \4670 );
nand \U$4329 ( \4672 , \4629 , \4590 );
nand \U$4330 ( \4673 , \4671 , \4672 );
xor \U$4331 ( \4674 , \4553 , \4673 );
nand \U$4332 ( \4675 , \524 , \530 );
nor \U$4333 ( \4676 , \4675 , \4355 );
not \U$4334 ( \4677 , \4676 );
not \U$4335 ( \4678 , \4361 );
or \U$4336 ( \4679 , \4677 , \4678 );
not \U$4337 ( \4680 , \4675 );
nand \U$4338 ( \4681 , \4367 , \4368 );
and \U$4339 ( \4682 , \4680 , \4681 );
not \U$4340 ( \4683 , \530 );
not \U$4341 ( \4684 , \4374 );
or \U$4342 ( \4685 , \4683 , \4684 );
not \U$4343 ( \4686 , \636 );
nand \U$4344 ( \4687 , \4685 , \4686 );
nor \U$4345 ( \4688 , \4682 , \4687 );
nand \U$4346 ( \4689 , \4679 , \4688 );
nand \U$4347 ( \4690 , \4351 , \638 );
not \U$4348 ( \4691 , \4690 );
and \U$4349 ( \4692 , \4689 , \4691 );
not \U$4350 ( \4693 , \4689 );
and \U$4351 ( \4694 , \4693 , \4690 );
nor \U$4352 ( \4695 , \4692 , \4694 );
not \U$4353 ( \4696 , \4695 );
not \U$4354 ( \4697 , \4696 );
not \U$4355 ( \4698 , \4697 );
not \U$4356 ( \4699 , \4698 );
nand \U$4357 ( \4700 , \4699 , \1394 );
and \U$4358 ( \4701 , RIbb2e5a8_36, RIbb2e620_35);
not \U$4359 ( \4702 , RIbb2e5a8_36);
and \U$4360 ( \4703 , \4702 , \3866 );
nor \U$4361 ( \4704 , \4701 , \4703 );
not \U$4362 ( \4705 , \4704 );
and \U$4363 ( \4706 , RIbb2e5a8_36, RIbb2e530_37);
not \U$4364 ( \4707 , RIbb2e5a8_36);
not \U$4365 ( \4708 , RIbb2e530_37);
and \U$4366 ( \4709 , \4707 , \4708 );
nor \U$4367 ( \4710 , \4706 , \4709 );
nor \U$4368 ( \4711 , \4705 , \4710 );
buf \U$4369 ( \4712 , \4711 );
not \U$4370 ( \4713 , \4712 );
buf \U$4371 ( \4714 , \4710 );
not \U$4372 ( \4715 , \4714 );
and \U$4373 ( \4716 , \4713 , \4715 );
nor \U$4374 ( \4717 , \4716 , \3866 );
nand \U$4375 ( \4718 , \4700 , \4717 );
not \U$4376 ( \4719 , \4718 );
not \U$4377 ( \4720 , \1376 );
not \U$4378 ( \4721 , \4329 );
or \U$4379 ( \4722 , \4720 , \4721 );
not \U$4380 ( \4723 , \1394 );
not \U$4381 ( \4724 , \4393 );
or \U$4382 ( \4725 , \4723 , \4724 );
nand \U$4383 ( \4726 , \1392 , \4394 );
nand \U$4384 ( \4727 , \4725 , \4726 );
nand \U$4385 ( \4728 , \4727 , \1429 );
nand \U$4386 ( \4729 , \4722 , \4728 );
not \U$4387 ( \4730 , \4729 );
or \U$4388 ( \4731 , \4719 , \4730 );
nor \U$4389 ( \4732 , \4700 , \4717 );
not \U$4390 ( \4733 , \4732 );
nand \U$4391 ( \4734 , \4731 , \4733 );
not \U$4392 ( \4735 , \1147 );
not \U$4393 ( \4736 , \3897 );
or \U$4394 ( \4737 , \4735 , \4736 );
not \U$4395 ( \4738 , RIbb2f430_5);
not \U$4396 ( \4739 , \4029 );
or \U$4397 ( \4740 , \4738 , \4739 );
nand \U$4398 ( \4741 , \4030 , \1085 );
nand \U$4399 ( \4742 , \4740 , \4741 );
nand \U$4400 ( \4743 , \1090 , \4742 );
nand \U$4401 ( \4744 , \4737 , \4743 );
not \U$4402 ( \4745 , \4744 );
not \U$4403 ( \4746 , \1265 );
not \U$4404 ( \4747 , \1246 );
not \U$4405 ( \4748 , \3089 );
buf \U$4406 ( \4749 , \4748 );
not \U$4407 ( \4750 , \4749 );
or \U$4408 ( \4751 , \4747 , \4750 );
not \U$4409 ( \4752 , \3089 );
not \U$4410 ( \4753 , \4752 );
nand \U$4411 ( \4754 , \4753 , \1245 );
nand \U$4412 ( \4755 , \4751 , \4754 );
not \U$4413 ( \4756 , \4755 );
or \U$4414 ( \4757 , \4746 , \4756 );
nand \U$4415 ( \4758 , \4415 , \1294 );
nand \U$4416 ( \4759 , \4757 , \4758 );
not \U$4417 ( \4760 , \4759 );
or \U$4418 ( \4761 , \4745 , \4760 );
or \U$4419 ( \4762 , \4744 , \4759 );
not \U$4420 ( \4763 , \2077 );
not \U$4421 ( \4764 , RIbb2ecb0_21);
buf \U$4422 ( \4765 , \1109 );
not \U$4423 ( \4766 , \4765 );
not \U$4424 ( \4767 , \4766 );
or \U$4425 ( \4768 , \4764 , \4767 );
buf \U$4426 ( \4769 , \1111 );
buf \U$4427 ( \4770 , \4769 );
nand \U$4428 ( \4771 , \4770 , \2254 );
nand \U$4429 ( \4772 , \4768 , \4771 );
not \U$4430 ( \4773 , \4772 );
or \U$4431 ( \4774 , \4763 , \4773 );
nand \U$4432 ( \4775 , \3943 , \2078 );
nand \U$4433 ( \4776 , \4774 , \4775 );
nand \U$4434 ( \4777 , \4762 , \4776 );
nand \U$4435 ( \4778 , \4761 , \4777 );
xor \U$4436 ( \4779 , \4734 , \4778 );
not \U$4437 ( \4780 , \3887 );
not \U$4438 ( \4781 , RIbb2e710_33);
not \U$4439 ( \4782 , \1579 );
or \U$4440 ( \4783 , \4781 , \4782 );
not \U$4441 ( \4784 , \894 );
not \U$4442 ( \4785 , RIbb2e710_33);
nand \U$4443 ( \4786 , \4784 , \4785 );
nand \U$4444 ( \4787 , \4783 , \4786 );
not \U$4445 ( \4788 , \4787 );
or \U$4446 ( \4789 , \4780 , \4788 );
buf \U$4447 ( \4790 , \4075 );
buf \U$4448 ( \4791 , \4790 );
nand \U$4449 ( \4792 , \3879 , \4791 );
nand \U$4450 ( \4793 , \4789 , \4792 );
not \U$4451 ( \4794 , \2925 );
not \U$4452 ( \4795 , \4467 );
or \U$4453 ( \4796 , \4794 , \4795 );
not \U$4454 ( \4797 , RIbb2e8f0_29);
not \U$4455 ( \4798 , \953 );
or \U$4456 ( \4799 , \4797 , \4798 );
not \U$4457 ( \4800 , RIbb2e8f0_29);
nand \U$4458 ( \4801 , \956 , \4800 );
nand \U$4459 ( \4802 , \4799 , \4801 );
nand \U$4460 ( \4803 , \4802 , \2922 );
nand \U$4461 ( \4804 , \4796 , \4803 );
xor \U$4462 ( \4805 , \4793 , \4804 );
not \U$4463 ( \4806 , \855 );
not \U$4464 ( \4807 , \4401 );
or \U$4465 ( \4808 , \4806 , \4807 );
not \U$4466 ( \4809 , RIbb2eda0_19);
not \U$4467 ( \4810 , \1170 );
or \U$4468 ( \4811 , \4809 , \4810 );
nand \U$4469 ( \4812 , \3736 , \843 );
nand \U$4470 ( \4813 , \4811 , \4812 );
nand \U$4471 ( \4814 , \4813 , \853 );
nand \U$4472 ( \4815 , \4808 , \4814 );
and \U$4473 ( \4816 , \4805 , \4815 );
and \U$4474 ( \4817 , \4793 , \4804 );
or \U$4475 ( \4818 , \4816 , \4817 );
and \U$4476 ( \4819 , \4779 , \4818 );
and \U$4477 ( \4820 , \4734 , \4778 );
or \U$4478 ( \4821 , \4819 , \4820 );
and \U$4479 ( \4822 , \4674 , \4821 );
and \U$4480 ( \4823 , \4553 , \4673 );
or \U$4481 ( \4824 , \4822 , \4823 );
xor \U$4482 ( \4825 , \4438 , \4491 );
xnor \U$4483 ( \4826 , \4825 , \4494 );
xor \U$4484 ( \4827 , \4824 , \4826 );
xor \U$4485 ( \4828 , \4441 , \4443 );
xor \U$4486 ( \4829 , \4828 , \4488 );
xor \U$4487 ( \4830 , \4305 , \4281 );
xnor \U$4488 ( \4831 , \4830 , \4293 );
not \U$4489 ( \4832 , \4831 );
xnor \U$4490 ( \4833 , \4486 , \4473 );
and \U$4491 ( \4834 , \4833 , \4469 );
not \U$4492 ( \4835 , \4833 );
and \U$4493 ( \4836 , \4835 , \4470 );
nor \U$4494 ( \4837 , \4834 , \4836 );
not \U$4495 ( \4838 , \4837 );
or \U$4496 ( \4839 , \4832 , \4838 );
xor \U$4497 ( \4840 , \3937 , \3947 );
xor \U$4498 ( \4841 , \4840 , \3965 );
nand \U$4499 ( \4842 , \4839 , \4841 );
not \U$4500 ( \4843 , \4837 );
not \U$4501 ( \4844 , \4831 );
nand \U$4502 ( \4845 , \4843 , \4844 );
nand \U$4503 ( \4846 , \4842 , \4845 );
xor \U$4504 ( \4847 , \4829 , \4846 );
not \U$4505 ( \4848 , \4308 );
not \U$4506 ( \4849 , \4420 );
not \U$4507 ( \4850 , \4849 );
or \U$4508 ( \4851 , \4848 , \4850 );
or \U$4509 ( \4852 , \4308 , \4849 );
nand \U$4510 ( \4853 , \4851 , \4852 );
xor \U$4511 ( \4854 , \4349 , \4853 );
and \U$4512 ( \4855 , \4847 , \4854 );
and \U$4513 ( \4856 , \4829 , \4846 );
or \U$4514 ( \4857 , \4855 , \4856 );
and \U$4515 ( \4858 , \4827 , \4857 );
and \U$4516 ( \4859 , \4824 , \4826 );
or \U$4517 ( \4860 , \4858 , \4859 );
nand \U$4518 ( \4861 , \4547 , \4860 );
nand \U$4519 ( \4862 , \4546 , \4861 );
and \U$4520 ( \4863 , \4514 , \4862 );
and \U$4521 ( \4864 , \3863 , \4513 );
or \U$4522 ( \4865 , \4863 , \4864 );
xor \U$4523 ( \4866 , \2927 , \2985 );
and \U$4524 ( \4867 , \4866 , \3074 );
and \U$4525 ( \4868 , \2927 , \2985 );
or \U$4526 ( \4869 , \4867 , \4868 );
not \U$4527 ( \4870 , \2927 );
not \U$4528 ( \4871 , \1430 );
not \U$4529 ( \4872 , \3716 );
or \U$4530 ( \4873 , \4871 , \4872 );
xor \U$4531 ( \4874 , \1313 , \3632 );
nand \U$4532 ( \4875 , \4874 , \1376 );
nand \U$4533 ( \4876 , \4873 , \4875 );
xor \U$4534 ( \4877 , \4870 , \4876 );
xor \U$4535 ( \4878 , \3670 , \3680 );
and \U$4536 ( \4879 , \4878 , \3691 );
and \U$4537 ( \4880 , \3670 , \3680 );
or \U$4538 ( \4881 , \4879 , \4880 );
xor \U$4539 ( \4882 , \4877 , \4881 );
xor \U$4540 ( \4883 , \4869 , \4882 );
xor \U$4541 ( \4884 , \3379 , \3435 );
and \U$4542 ( \4885 , \4884 , \3510 );
and \U$4543 ( \4886 , \3379 , \3435 );
or \U$4544 ( \4887 , \4885 , \4886 );
xor \U$4545 ( \4888 , \4883 , \4887 );
xor \U$4546 ( \4889 , \3601 , \3668 );
and \U$4547 ( \4890 , \4889 , \3756 );
and \U$4548 ( \4891 , \3601 , \3668 );
or \U$4549 ( \4892 , \4890 , \4891 );
xor \U$4550 ( \4893 , \4888 , \4892 );
xor \U$4551 ( \4894 , \4190 , \4225 );
and \U$4552 ( \4895 , \4894 , \4257 );
and \U$4553 ( \4896 , \4190 , \4225 );
or \U$4554 ( \4897 , \4895 , \4896 );
xor \U$4555 ( \4898 , \3732 , \3742 );
and \U$4556 ( \4899 , \4898 , \3754 );
and \U$4557 ( \4900 , \3732 , \3742 );
or \U$4558 ( \4901 , \4899 , \4900 );
xor \U$4559 ( \4902 , \4236 , \4245 );
and \U$4560 ( \4903 , \4902 , \4256 );
and \U$4561 ( \4904 , \4236 , \4245 );
or \U$4562 ( \4905 , \4903 , \4904 );
xor \U$4563 ( \4906 , \4901 , \4905 );
xor \U$4564 ( \4907 , \4200 , \4210 );
and \U$4565 ( \4908 , \4907 , \4224 );
and \U$4566 ( \4909 , \4200 , \4210 );
or \U$4567 ( \4910 , \4908 , \4909 );
xor \U$4568 ( \4911 , \4906 , \4910 );
xor \U$4569 ( \4912 , \4897 , \4911 );
xor \U$4570 ( \4913 , \3692 , \3721 );
and \U$4571 ( \4914 , \4913 , \3755 );
and \U$4572 ( \4915 , \3692 , \3721 );
or \U$4573 ( \4916 , \4914 , \4915 );
xor \U$4574 ( \4917 , \4912 , \4916 );
xor \U$4575 ( \4918 , \4893 , \4917 );
not \U$4576 ( \4919 , \4186 );
not \U$4577 ( \4920 , \4258 );
or \U$4578 ( \4921 , \4919 , \4920 );
not \U$4579 ( \4922 , \4186 );
nand \U$4580 ( \4923 , \4922 , \4259 );
nand \U$4581 ( \4924 , \4269 , \4923 );
nand \U$4582 ( \4925 , \4921 , \4924 );
xor \U$4583 ( \4926 , \3703 , \3713 );
and \U$4584 ( \4927 , \4926 , \3720 );
and \U$4585 ( \4928 , \3703 , \3713 );
or \U$4586 ( \4929 , \4927 , \4928 );
or \U$4587 ( \4930 , \2922 , \2925 );
nand \U$4588 ( \4931 , \4930 , RIbb2e8f0_29);
not \U$4589 ( \4932 , \3445 );
not \U$4590 ( \4933 , \3676 );
or \U$4591 ( \4934 , \4932 , \4933 );
not \U$4592 ( \4935 , RIbb2e9e0_27);
not \U$4593 ( \4936 , \814 );
or \U$4594 ( \4937 , \4935 , \4936 );
nand \U$4595 ( \4938 , \2251 , \3462 );
nand \U$4596 ( \4939 , \4937 , \4938 );
nand \U$4597 ( \4940 , \4939 , \3465 );
nand \U$4598 ( \4941 , \4934 , \4940 );
xor \U$4599 ( \4942 , \4931 , \4941 );
not \U$4600 ( \4943 , \3383 );
not \U$4601 ( \4944 , RIbb2ebc0_23);
not \U$4602 ( \4945 , \989 );
or \U$4603 ( \4946 , \4944 , \4945 );
nand \U$4604 ( \4947 , \987 , \3396 );
nand \U$4605 ( \4948 , \4946 , \4947 );
not \U$4606 ( \4949 , \4948 );
or \U$4607 ( \4950 , \4943 , \4949 );
nand \U$4608 ( \4951 , \3687 , \3407 );
nand \U$4609 ( \4952 , \4950 , \4951 );
xor \U$4610 ( \4953 , \4942 , \4952 );
xor \U$4611 ( \4954 , \4929 , \4953 );
and \U$4612 ( \4955 , \1393 , \3024 );
not \U$4613 ( \4956 , \998 );
and \U$4614 ( \4957 , \1283 , \906 );
not \U$4615 ( \4958 , \1283 );
and \U$4616 ( \4959 , \4958 , RIbb2f070_13);
or \U$4617 ( \4960 , \4957 , \4959 );
not \U$4618 ( \4961 , \4960 );
or \U$4619 ( \4962 , \4956 , \4961 );
nand \U$4620 ( \4963 , \3740 , \916 );
nand \U$4621 ( \4964 , \4962 , \4963 );
xor \U$4622 ( \4965 , \4955 , \4964 );
or \U$4623 ( \4966 , \3751 , \1575 );
not \U$4624 ( \4967 , RIbb2ef80_15);
nand \U$4625 ( \4968 , \4967 , \1139 );
not \U$4626 ( \4969 , \4968 );
not \U$4627 ( \4970 , RIbb2ef80_15);
nor \U$4628 ( \4971 , \4970 , \1139 );
nor \U$4629 ( \4972 , \4969 , \4971 );
or \U$4630 ( \4973 , \4972 , \1584 );
nand \U$4631 ( \4974 , \4966 , \4973 );
xor \U$4632 ( \4975 , \4965 , \4974 );
xor \U$4633 ( \4976 , \4954 , \4975 );
not \U$4634 ( \4977 , \1737 );
not \U$4635 ( \4978 , RIbb2f340_7);
not \U$4636 ( \4979 , \2116 );
or \U$4637 ( \4980 , \4978 , \4979 );
nand \U$4638 ( \4981 , \4450 , \2700 );
nand \U$4639 ( \4982 , \4980 , \4981 );
not \U$4640 ( \4983 , \4982 );
or \U$4641 ( \4984 , \4977 , \4983 );
nand \U$4642 ( \4985 , \4208 , \1702 );
nand \U$4643 ( \4986 , \4984 , \4985 );
not \U$4644 ( \4987 , \2980 );
not \U$4645 ( \4988 , \4241 );
or \U$4646 ( \4989 , \4987 , \4988 );
and \U$4647 ( \4990 , RIbb2ead0_25, \1509 );
not \U$4648 ( \4991 , RIbb2ead0_25);
and \U$4649 ( \4992 , \4991 , \4315 );
or \U$4650 ( \4993 , \4990 , \4992 );
nand \U$4651 ( \4994 , \4993 , \2963 );
nand \U$4652 ( \4995 , \4989 , \4994 );
xor \U$4653 ( \4996 , \4986 , \4995 );
not \U$4654 ( \4997 , \853 );
not \U$4655 ( \4998 , \4198 );
or \U$4656 ( \4999 , \4997 , \4998 );
not \U$4657 ( \5000 , RIbb2eda0_19);
not \U$4658 ( \5001 , \1550 );
or \U$4659 ( \5002 , \5000 , \5001 );
not \U$4660 ( \5003 , \1547 );
not \U$4661 ( \5004 , \5003 );
nand \U$4662 ( \5005 , \5004 , \1776 );
nand \U$4663 ( \5006 , \5002 , \5005 );
nand \U$4664 ( \5007 , \5006 , \855 );
nand \U$4665 ( \5008 , \4999 , \5007 );
not \U$4666 ( \5009 , \5008 );
and \U$4667 ( \5010 , \4996 , \5009 );
not \U$4668 ( \5011 , \4996 );
and \U$4669 ( \5012 , \5011 , \5008 );
nor \U$4670 ( \5013 , \5010 , \5012 );
not \U$4671 ( \5014 , \1090 );
not \U$4672 ( \5015 , \4222 );
or \U$4673 ( \5016 , \5014 , \5015 );
not \U$4674 ( \5017 , RIbb2f430_5);
not \U$4675 ( \5018 , \3517 );
or \U$4676 ( \5019 , \5017 , \5018 );
nand \U$4677 ( \5020 , \3347 , \1647 );
nand \U$4678 ( \5021 , \5019 , \5020 );
nand \U$4679 ( \5022 , \5021 , \1147 );
nand \U$4680 ( \5023 , \5016 , \5022 );
not \U$4681 ( \5024 , \1294 );
not \U$4682 ( \5025 , \1290 );
not \U$4683 ( \5026 , \3143 );
or \U$4684 ( \5027 , \5025 , \5026 );
not \U$4685 ( \5028 , \3143 );
nand \U$4686 ( \5029 , \5028 , \1289 );
nand \U$4687 ( \5030 , \5027 , \5029 );
not \U$4688 ( \5031 , \5030 );
or \U$4689 ( \5032 , \5024 , \5031 );
nand \U$4690 ( \5033 , \3709 , \1265 );
nand \U$4691 ( \5034 , \5032 , \5033 );
xor \U$4692 ( \5035 , \5023 , \5034 );
not \U$4693 ( \5036 , \836 );
not \U$4694 ( \5037 , RIbb2ee90_17);
not \U$4695 ( \5038 , \1689 );
or \U$4696 ( \5039 , \5037 , \5038 );
nand \U$4697 ( \5040 , \1691 , \816 );
nand \U$4698 ( \5041 , \5039 , \5040 );
not \U$4699 ( \5042 , \5041 );
or \U$4700 ( \5043 , \5036 , \5042 );
nand \U$4701 ( \5044 , \3701 , \832 );
nand \U$4702 ( \5045 , \5043 , \5044 );
xor \U$4703 ( \5046 , \5035 , \5045 );
xor \U$4704 ( \5047 , \5013 , \5046 );
not \U$4705 ( \5048 , \1077 );
not \U$4706 ( \5049 , RIbb2f160_11);
not \U$4707 ( \5050 , \1820 );
or \U$4708 ( \5051 , \5049 , \5050 );
nand \U$4709 ( \5052 , \1387 , \1048 );
nand \U$4710 ( \5053 , \5051 , \5052 );
not \U$4711 ( \5054 , \5053 );
or \U$4712 ( \5055 , \5048 , \5054 );
nand \U$4713 ( \5056 , \4232 , \1011 );
nand \U$4714 ( \5057 , \5055 , \5056 );
not \U$4715 ( \5058 , \1533 );
not \U$4716 ( \5059 , \4254 );
or \U$4717 ( \5060 , \5058 , \5059 );
not \U$4718 ( \5061 , RIbb2f250_9);
not \U$4719 ( \5062 , \1340 );
or \U$4720 ( \5063 , \5061 , \5062 );
not \U$4721 ( \5064 , RIbb2f250_9);
nand \U$4722 ( \5065 , \3495 , \5064 );
nand \U$4723 ( \5066 , \5063 , \5065 );
nand \U$4724 ( \5067 , \5066 , \1570 );
nand \U$4725 ( \5068 , \5060 , \5067 );
not \U$4726 ( \5069 , \2078 );
not \U$4727 ( \5070 , RIbb2ecb0_21);
not \U$4728 ( \5071 , \1072 );
or \U$4729 ( \5072 , \5070 , \5071 );
nand \U$4730 ( \5073 , \1888 , \2067 );
nand \U$4731 ( \5074 , \5072 , \5073 );
not \U$4732 ( \5075 , \5074 );
or \U$4733 ( \5076 , \5069 , \5075 );
nand \U$4734 ( \5077 , \3728 , \2077 );
nand \U$4735 ( \5078 , \5076 , \5077 );
xor \U$4736 ( \5079 , \5068 , \5078 );
xor \U$4737 ( \5080 , \5057 , \5079 );
xnor \U$4738 ( \5081 , \5047 , \5080 );
xor \U$4739 ( \5082 , \4976 , \5081 );
not \U$4740 ( \5083 , \3075 );
not \U$4741 ( \5084 , \3303 );
or \U$4742 ( \5085 , \5083 , \5084 );
or \U$4743 ( \5086 , \3303 , \3075 );
nand \U$4744 ( \5087 , \5086 , \3511 );
nand \U$4745 ( \5088 , \5085 , \5087 );
xor \U$4746 ( \5089 , \5082 , \5088 );
xor \U$4747 ( \5090 , \4925 , \5089 );
not \U$4748 ( \5091 , \3513 );
not \U$4749 ( \5092 , \3857 );
or \U$4750 ( \5093 , \5091 , \5092 );
not \U$4751 ( \5094 , \3858 );
not \U$4752 ( \5095 , \3512 );
or \U$4753 ( \5096 , \5094 , \5095 );
nand \U$4754 ( \5097 , \5096 , \3757 );
nand \U$4755 ( \5098 , \5093 , \5097 );
xor \U$4756 ( \5099 , \5090 , \5098 );
xor \U$4757 ( \5100 , \4918 , \5099 );
not \U$4758 ( \5101 , \4505 );
nand \U$4759 ( \5102 , \5101 , \4270 );
not \U$4760 ( \5103 , \5102 );
not \U$4761 ( \5104 , \4125 );
or \U$4762 ( \5105 , \5103 , \5104 );
not \U$4763 ( \5106 , \4270 );
nand \U$4764 ( \5107 , \5106 , \4505 );
nand \U$4765 ( \5108 , \5105 , \5107 );
xor \U$4766 ( \5109 , \5100 , \5108 );
or \U$4767 ( \5110 , \4865 , \5109 );
xor \U$4768 ( \5111 , \4918 , \5099 );
and \U$4769 ( \5112 , \5111 , \5108 );
and \U$4770 ( \5113 , \4918 , \5099 );
or \U$4771 ( \5114 , \5112 , \5113 );
not \U$4772 ( \5115 , \5114 );
not \U$4773 ( \5116 , \1702 );
not \U$4774 ( \5117 , \4982 );
or \U$4775 ( \5118 , \5116 , \5117 );
not \U$4776 ( \5119 , RIbb2f340_7);
not \U$4777 ( \5120 , \1854 );
or \U$4778 ( \5121 , \5119 , \5120 );
nand \U$4779 ( \5122 , \3503 , \1734 );
nand \U$4780 ( \5123 , \5121 , \5122 );
nand \U$4781 ( \5124 , \5123 , \1737 );
nand \U$4782 ( \5125 , \5118 , \5124 );
not \U$4783 ( \5126 , \832 );
not \U$4784 ( \5127 , \5041 );
or \U$4785 ( \5128 , \5126 , \5127 );
not \U$4786 ( \5129 , RIbb2ee90_17);
not \U$4787 ( \5130 , \1730 );
not \U$4788 ( \5131 , \5130 );
or \U$4789 ( \5132 , \5129 , \5131 );
nand \U$4790 ( \5133 , \1733 , \816 );
nand \U$4791 ( \5134 , \5132 , \5133 );
nand \U$4792 ( \5135 , \5134 , \836 );
nand \U$4793 ( \5136 , \5128 , \5135 );
xor \U$4794 ( \5137 , \5125 , \5136 );
not \U$4795 ( \5138 , \3383 );
not \U$4796 ( \5139 , RIbb2ebc0_23);
not \U$4797 ( \5140 , \1659 );
or \U$4798 ( \5141 , \5139 , \5140 );
nand \U$4799 ( \5142 , \1477 , \3401 );
nand \U$4800 ( \5143 , \5141 , \5142 );
not \U$4801 ( \5144 , \5143 );
or \U$4802 ( \5145 , \5138 , \5144 );
nand \U$4803 ( \5146 , \4948 , \3407 );
nand \U$4804 ( \5147 , \5145 , \5146 );
xor \U$4805 ( \5148 , \5137 , \5147 );
xor \U$4806 ( \5149 , \4870 , \4876 );
and \U$4807 ( \5150 , \5149 , \4881 );
and \U$4808 ( \5151 , \4870 , \4876 );
or \U$4809 ( \5152 , \5150 , \5151 );
xor \U$4810 ( \5153 , \5148 , \5152 );
xor \U$4811 ( \5154 , \4901 , \4905 );
and \U$4812 ( \5155 , \5154 , \4910 );
and \U$4813 ( \5156 , \4901 , \4905 );
or \U$4814 ( \5157 , \5155 , \5156 );
xor \U$4815 ( \5158 , \5153 , \5157 );
xor \U$4816 ( \5159 , \4897 , \4911 );
and \U$4817 ( \5160 , \5159 , \4916 );
and \U$4818 ( \5161 , \4897 , \4911 );
or \U$4819 ( \5162 , \5160 , \5161 );
xor \U$4820 ( \5163 , \5158 , \5162 );
not \U$4821 ( \5164 , \5013 );
not \U$4822 ( \5165 , \5164 );
not \U$4823 ( \5166 , \5080 );
or \U$4824 ( \5167 , \5165 , \5166 );
or \U$4825 ( \5168 , \5080 , \5164 );
nand \U$4826 ( \5169 , \5168 , \5046 );
nand \U$4827 ( \5170 , \5167 , \5169 );
xor \U$4828 ( \5171 , \4955 , \4964 );
and \U$4829 ( \5172 , \5171 , \4974 );
and \U$4830 ( \5173 , \4955 , \4964 );
or \U$4831 ( \5174 , \5172 , \5173 );
xor \U$4832 ( \5175 , \4931 , \4941 );
and \U$4833 ( \5176 , \5175 , \4952 );
and \U$4834 ( \5177 , \4931 , \4941 );
or \U$4835 ( \5178 , \5176 , \5177 );
not \U$4836 ( \5179 , \5178 );
and \U$4837 ( \5180 , \5174 , \5179 );
not \U$4838 ( \5181 , \5174 );
and \U$4839 ( \5182 , \5181 , \5178 );
or \U$4840 ( \5183 , \5180 , \5182 );
or \U$4841 ( \5184 , \5057 , \5068 );
nand \U$4842 ( \5185 , \5184 , \5078 );
nand \U$4843 ( \5186 , \5068 , \5057 );
nand \U$4844 ( \5187 , \5185 , \5186 );
not \U$4845 ( \5188 , \5187 );
and \U$4846 ( \5189 , \5183 , \5188 );
not \U$4847 ( \5190 , \5183 );
and \U$4848 ( \5191 , \5190 , \5187 );
nor \U$4849 ( \5192 , \5189 , \5191 );
xnor \U$4850 ( \5193 , \5170 , \5192 );
xor \U$4851 ( \5194 , \5023 , \5034 );
and \U$4852 ( \5195 , \5194 , \5045 );
and \U$4853 ( \5196 , \5023 , \5034 );
or \U$4854 ( \5197 , \5195 , \5196 );
not \U$4855 ( \5198 , \4995 );
buf \U$4856 ( \5199 , \4986 );
not \U$4857 ( \5200 , \5199 );
or \U$4858 ( \5201 , \5198 , \5200 );
or \U$4859 ( \5202 , \5199 , \4995 );
nand \U$4860 ( \5203 , \5202 , \5008 );
nand \U$4861 ( \5204 , \5201 , \5203 );
xor \U$4862 ( \5205 , \5197 , \5204 );
and \U$4863 ( \5206 , \1313 , \3654 );
nand \U$4864 ( \5207 , \4939 , \3445 );
nand \U$4865 ( \5208 , \3465 , RIbb2e9e0_27);
and \U$4866 ( \5209 , \5207 , \5208 );
xor \U$4867 ( \5210 , \5206 , \5209 );
not \U$4868 ( \5211 , \1430 );
not \U$4869 ( \5212 , \4874 );
or \U$4870 ( \5213 , \5211 , \5212 );
xor \U$4871 ( \5214 , \1394 , \3202 );
nand \U$4872 ( \5215 , \5214 , \1376 );
nand \U$4873 ( \5216 , \5213 , \5215 );
xor \U$4874 ( \5217 , \5210 , \5216 );
xor \U$4875 ( \5218 , \5205 , \5217 );
xnor \U$4876 ( \5219 , \5193 , \5218 );
not \U$4877 ( \5220 , \5219 );
xnor \U$4878 ( \5221 , \5163 , \5220 );
xor \U$4879 ( \5222 , \4925 , \5089 );
and \U$4880 ( \5223 , \5222 , \5098 );
and \U$4881 ( \5224 , \4925 , \5089 );
or \U$4882 ( \5225 , \5223 , \5224 );
not \U$4883 ( \5226 , \5225 );
xor \U$4884 ( \5227 , \5221 , \5226 );
xor \U$4885 ( \5228 , \4888 , \4892 );
and \U$4886 ( \5229 , \5228 , \4917 );
and \U$4887 ( \5230 , \4888 , \4892 );
or \U$4888 ( \5231 , \5229 , \5230 );
xor \U$4889 ( \5232 , \4976 , \5081 );
and \U$4890 ( \5233 , \5232 , \5088 );
and \U$4891 ( \5234 , \4976 , \5081 );
or \U$4892 ( \5235 , \5233 , \5234 );
xor \U$4893 ( \5236 , \4929 , \4953 );
and \U$4894 ( \5237 , \5236 , \4975 );
and \U$4895 ( \5238 , \4929 , \4953 );
or \U$4896 ( \5239 , \5237 , \5238 );
not \U$4897 ( \5240 , \5239 );
not \U$4898 ( \5241 , \5240 );
not \U$4899 ( \5242 , \2963 );
and \U$4900 ( \5243 , RIbb2ead0_25, \1579 );
not \U$4901 ( \5244 , RIbb2ead0_25);
and \U$4902 ( \5245 , \5244 , \1580 );
or \U$4903 ( \5246 , \5243 , \5245 );
not \U$4904 ( \5247 , \5246 );
or \U$4905 ( \5248 , \5242 , \5247 );
nand \U$4906 ( \5249 , \4993 , \2980 );
nand \U$4907 ( \5250 , \5248 , \5249 );
not \U$4908 ( \5251 , \2078 );
not \U$4909 ( \5252 , RIbb2ecb0_21);
not \U$4910 ( \5253 , \2399 );
or \U$4911 ( \5254 , \5252 , \5253 );
nand \U$4912 ( \5255 , \957 , \849 );
nand \U$4913 ( \5256 , \5254 , \5255 );
not \U$4914 ( \5257 , \5256 );
or \U$4915 ( \5258 , \5251 , \5257 );
nand \U$4916 ( \5259 , \5074 , \2077 );
nand \U$4917 ( \5260 , \5258 , \5259 );
xor \U$4918 ( \5261 , \5250 , \5260 );
not \U$4919 ( \5262 , \998 );
not \U$4920 ( \5263 , RIbb2f070_13);
not \U$4921 ( \5264 , \3066 );
or \U$4922 ( \5265 , \5263 , \5264 );
nand \U$4923 ( \5266 , \3067 , \1656 );
nand \U$4924 ( \5267 , \5265 , \5266 );
not \U$4925 ( \5268 , \5267 );
or \U$4926 ( \5269 , \5262 , \5268 );
nand \U$4927 ( \5270 , \4960 , \916 );
nand \U$4928 ( \5271 , \5269 , \5270 );
xor \U$4929 ( \5272 , \5261 , \5271 );
not \U$4930 ( \5273 , \855 );
not \U$4931 ( \5274 , RIbb2eda0_19);
not \U$4932 ( \5275 , \1039 );
or \U$4933 ( \5276 , \5274 , \5275 );
not \U$4934 ( \5277 , RIbb2eda0_19);
nand \U$4935 ( \5278 , \1038 , \5277 );
nand \U$4936 ( \5279 , \5276 , \5278 );
not \U$4937 ( \5280 , \5279 );
or \U$4938 ( \5281 , \5273 , \5280 );
nand \U$4939 ( \5282 , \5006 , \853 );
nand \U$4940 ( \5283 , \5281 , \5282 );
not \U$4941 ( \5284 , \5283 );
not \U$4942 ( \5285 , \1570 );
not \U$4943 ( \5286 , RIbb2f250_9);
not \U$4944 ( \5287 , \2052 );
or \U$4945 ( \5288 , \5286 , \5287 );
nand \U$4946 ( \5289 , \1421 , \1566 );
nand \U$4947 ( \5290 , \5288 , \5289 );
not \U$4948 ( \5291 , \5290 );
or \U$4949 ( \5292 , \5285 , \5291 );
nand \U$4950 ( \5293 , \5066 , \1533 );
nand \U$4951 ( \5294 , \5292 , \5293 );
not \U$4952 ( \5295 , \5294 );
not \U$4953 ( \5296 , \5295 );
or \U$4954 ( \5297 , \5284 , \5296 );
or \U$4955 ( \5298 , \5295 , \5283 );
nand \U$4956 ( \5299 , \5297 , \5298 );
not \U$4957 ( \5300 , \1011 );
not \U$4958 ( \5301 , \5053 );
or \U$4959 ( \5302 , \5300 , \5301 );
not \U$4960 ( \5303 , RIbb2f160_11);
not \U$4961 ( \5304 , \3991 );
or \U$4962 ( \5305 , \5303 , \5304 );
nand \U$4963 ( \5306 , \3109 , \1805 );
nand \U$4964 ( \5307 , \5305 , \5306 );
nand \U$4965 ( \5308 , \5307 , \1077 );
nand \U$4966 ( \5309 , \5302 , \5308 );
not \U$4967 ( \5310 , \5309 );
and \U$4968 ( \5311 , \5299 , \5310 );
not \U$4969 ( \5312 , \5299 );
and \U$4970 ( \5313 , \5312 , \5309 );
nor \U$4971 ( \5314 , \5311 , \5313 );
xor \U$4972 ( \5315 , \5272 , \5314 );
not \U$4973 ( \5316 , \1147 );
not \U$4974 ( \5317 , RIbb2f430_5);
not \U$4975 ( \5318 , \2224 );
or \U$4976 ( \5319 , \5317 , \5318 );
nand \U$4977 ( \5320 , \2225 , \1980 );
nand \U$4978 ( \5321 , \5319 , \5320 );
not \U$4979 ( \5322 , \5321 );
or \U$4980 ( \5323 , \5316 , \5322 );
nand \U$4981 ( \5324 , \5021 , \1090 );
nand \U$4982 ( \5325 , \5323 , \5324 );
not \U$4983 ( \5326 , \1265 );
not \U$4984 ( \5327 , \5030 );
or \U$4985 ( \5328 , \5326 , \5327 );
not \U$4986 ( \5329 , \1290 );
not \U$4987 ( \5330 , \4216 );
or \U$4988 ( \5331 , \5329 , \5330 );
nand \U$4989 ( \5332 , \4220 , \1289 );
nand \U$4990 ( \5333 , \5331 , \5332 );
nand \U$4991 ( \5334 , \5333 , \1294 );
nand \U$4992 ( \5335 , \5328 , \5334 );
xor \U$4993 ( \5336 , \5325 , \5335 );
not \U$4994 ( \5337 , \3105 );
and \U$4995 ( \5338 , RIbb2ef80_15, \1644 );
not \U$4996 ( \5339 , RIbb2ef80_15);
and \U$4997 ( \5340 , \5339 , \1643 );
or \U$4998 ( \5341 , \5338 , \5340 );
not \U$4999 ( \5342 , \5341 );
or \U$5000 ( \5343 , \5337 , \5342 );
not \U$5001 ( \5344 , RIbb2ef80_15);
not \U$5002 ( \5345 , \1140 );
or \U$5003 ( \5346 , \5344 , \5345 );
nand \U$5004 ( \5347 , \5346 , \4968 );
nand \U$5005 ( \5348 , \5347 , \1445 );
nand \U$5006 ( \5349 , \5343 , \5348 );
xor \U$5007 ( \5350 , \5336 , \5349 );
xor \U$5008 ( \5351 , \5315 , \5350 );
not \U$5009 ( \5352 , \5351 );
not \U$5010 ( \5353 , \5352 );
or \U$5011 ( \5354 , \5241 , \5353 );
nand \U$5012 ( \5355 , \5351 , \5239 );
nand \U$5013 ( \5356 , \5354 , \5355 );
xor \U$5014 ( \5357 , \4869 , \4882 );
and \U$5015 ( \5358 , \5357 , \4887 );
and \U$5016 ( \5359 , \4869 , \4882 );
or \U$5017 ( \5360 , \5358 , \5359 );
not \U$5018 ( \5361 , \5360 );
and \U$5019 ( \5362 , \5356 , \5361 );
not \U$5020 ( \5363 , \5356 );
and \U$5021 ( \5364 , \5363 , \5360 );
nor \U$5022 ( \5365 , \5362 , \5364 );
xnor \U$5023 ( \5366 , \5235 , \5365 );
not \U$5024 ( \5367 , \5366 );
xor \U$5025 ( \5368 , \5231 , \5367 );
xor \U$5026 ( \5369 , \5227 , \5368 );
nand \U$5027 ( \5370 , \5115 , \5369 );
nand \U$5028 ( \5371 , \5110 , \5370 );
xor \U$5029 ( \5372 , \5148 , \5152 );
and \U$5030 ( \5373 , \5372 , \5157 );
and \U$5031 ( \5374 , \5148 , \5152 );
or \U$5032 ( \5375 , \5373 , \5374 );
xor \U$5033 ( \5376 , \5197 , \5204 );
and \U$5034 ( \5377 , \5376 , \5217 );
and \U$5035 ( \5378 , \5197 , \5204 );
or \U$5036 ( \5379 , \5377 , \5378 );
not \U$5037 ( \5380 , \5209 );
not \U$5038 ( \5381 , \5295 );
not \U$5039 ( \5382 , \5310 );
or \U$5040 ( \5383 , \5381 , \5382 );
nand \U$5041 ( \5384 , \5383 , \5283 );
nand \U$5042 ( \5385 , \5294 , \5309 );
nand \U$5043 ( \5386 , \5384 , \5385 );
xor \U$5044 ( \5387 , \5380 , \5386 );
xor \U$5045 ( \5388 , \5250 , \5260 );
and \U$5046 ( \5389 , \5388 , \5271 );
and \U$5047 ( \5390 , \5250 , \5260 );
or \U$5048 ( \5391 , \5389 , \5390 );
xor \U$5049 ( \5392 , \5387 , \5391 );
xor \U$5050 ( \5393 , \5379 , \5392 );
not \U$5051 ( \5394 , \5136 );
not \U$5052 ( \5395 , \5125 );
or \U$5053 ( \5396 , \5394 , \5395 );
or \U$5054 ( \5397 , \5125 , \5136 );
nand \U$5055 ( \5398 , \5397 , \5147 );
nand \U$5056 ( \5399 , \5396 , \5398 );
xor \U$5057 ( \5400 , \5325 , \5335 );
and \U$5058 ( \5401 , \5400 , \5349 );
and \U$5059 ( \5402 , \5325 , \5335 );
or \U$5060 ( \5403 , \5401 , \5402 );
xor \U$5061 ( \5404 , \5399 , \5403 );
not \U$5062 ( \5405 , \1077 );
not \U$5063 ( \5406 , RIbb2f160_11);
not \U$5064 ( \5407 , \1283 );
not \U$5065 ( \5408 , \5407 );
or \U$5066 ( \5409 , \5406 , \5408 );
nand \U$5067 ( \5410 , \3291 , \1043 );
nand \U$5068 ( \5411 , \5409 , \5410 );
not \U$5069 ( \5412 , \5411 );
or \U$5070 ( \5413 , \5405 , \5412 );
nand \U$5071 ( \5414 , \5307 , \1011 );
nand \U$5072 ( \5415 , \5413 , \5414 );
and \U$5073 ( \5416 , \1656 , \3053 );
not \U$5074 ( \5417 , \1656 );
and \U$5075 ( \5418 , \5417 , \1140 );
nor \U$5076 ( \5419 , \5416 , \5418 );
not \U$5077 ( \5420 , \5419 );
not \U$5078 ( \5421 , \1662 );
and \U$5079 ( \5422 , \5420 , \5421 );
and \U$5080 ( \5423 , \5267 , \916 );
nor \U$5081 ( \5424 , \5422 , \5423 );
xor \U$5082 ( \5425 , \5415 , \5424 );
not \U$5083 ( \5426 , \855 );
not \U$5084 ( \5427 , RIbb2eda0_19);
not \U$5085 ( \5428 , \1072 );
or \U$5086 ( \5429 , \5427 , \5428 );
nand \U$5087 ( \5430 , \1888 , \1776 );
nand \U$5088 ( \5431 , \5429 , \5430 );
not \U$5089 ( \5432 , \5431 );
or \U$5090 ( \5433 , \5426 , \5432 );
nand \U$5091 ( \5434 , \5279 , \853 );
nand \U$5092 ( \5435 , \5433 , \5434 );
xnor \U$5093 ( \5436 , \5425 , \5435 );
xor \U$5094 ( \5437 , \5404 , \5436 );
xor \U$5095 ( \5438 , \5393 , \5437 );
xor \U$5096 ( \5439 , \5375 , \5438 );
not \U$5097 ( \5440 , \5192 );
or \U$5098 ( \5441 , \5440 , \5218 );
nand \U$5099 ( \5442 , \5441 , \5170 );
nand \U$5100 ( \5443 , \5218 , \5440 );
nand \U$5101 ( \5444 , \5442 , \5443 );
and \U$5102 ( \5445 , \5439 , \5444 );
and \U$5103 ( \5446 , \5375 , \5438 );
or \U$5104 ( \5447 , \5445 , \5446 );
xor \U$5105 ( \5448 , \5399 , \5403 );
and \U$5106 ( \5449 , \5448 , \5436 );
and \U$5107 ( \5450 , \5399 , \5403 );
or \U$5108 ( \5451 , \5449 , \5450 );
and \U$5109 ( \5452 , \1313 , \3632 );
not \U$5110 ( \5453 , \1376 );
xor \U$5111 ( \5454 , \1313 , \5028 );
not \U$5112 ( \5455 , \5454 );
or \U$5113 ( \5456 , \5453 , \5455 );
nand \U$5114 ( \5457 , \5214 , \1430 );
nand \U$5115 ( \5458 , \5456 , \5457 );
xor \U$5116 ( \5459 , \5452 , \5458 );
not \U$5117 ( \5460 , \1517 );
xor \U$5118 ( \5461 , RIbb2ef80_15, \1691 );
not \U$5119 ( \5462 , \5461 );
or \U$5120 ( \5463 , \5460 , \5462 );
nand \U$5121 ( \5464 , \5341 , \1445 );
nand \U$5122 ( \5465 , \5463 , \5464 );
and \U$5123 ( \5466 , \5459 , \5465 );
and \U$5124 ( \5467 , \5452 , \5458 );
or \U$5125 ( \5468 , \5466 , \5467 );
and \U$5126 ( \5469 , \1394 , \3202 );
not \U$5127 ( \5470 , \1430 );
not \U$5128 ( \5471 , \5454 );
or \U$5129 ( \5472 , \5470 , \5471 );
xor \U$5130 ( \5473 , \1394 , \4220 );
nand \U$5131 ( \5474 , \5473 , \1376 );
nand \U$5132 ( \5475 , \5472 , \5474 );
xor \U$5133 ( \5476 , \5469 , \5475 );
not \U$5134 ( \5477 , \2077 );
not \U$5135 ( \5478 , RIbb2ecb0_21);
not \U$5136 ( \5479 , \993 );
or \U$5137 ( \5480 , \5478 , \5479 );
not \U$5138 ( \5481 , RIbb2ecb0_21);
nand \U$5139 ( \5482 , \1939 , \5481 );
nand \U$5140 ( \5483 , \5480 , \5482 );
not \U$5141 ( \5484 , \5483 );
or \U$5142 ( \5485 , \5477 , \5484 );
and \U$5143 ( \5486 , \2249 , \1659 );
not \U$5144 ( \5487 , \2249 );
and \U$5145 ( \5488 , \5487 , \1477 );
nor \U$5146 ( \5489 , \5486 , \5488 );
nand \U$5147 ( \5490 , \5489 , \2078 );
nand \U$5148 ( \5491 , \5485 , \5490 );
xor \U$5149 ( \5492 , \5476 , \5491 );
xor \U$5150 ( \5493 , \5468 , \5492 );
not \U$5151 ( \5494 , \855 );
not \U$5152 ( \5495 , RIbb2eda0_19);
not \U$5153 ( \5496 , \2399 );
or \U$5154 ( \5497 , \5495 , \5496 );
nand \U$5155 ( \5498 , \957 , \1776 );
nand \U$5156 ( \5499 , \5497 , \5498 );
not \U$5157 ( \5500 , \5499 );
or \U$5158 ( \5501 , \5494 , \5500 );
nand \U$5159 ( \5502 , \5431 , \853 );
nand \U$5160 ( \5503 , \5501 , \5502 );
not \U$5161 ( \5504 , \3383 );
not \U$5162 ( \5505 , RIbb2ebc0_23);
not \U$5163 ( \5506 , \895 );
or \U$5164 ( \5507 , \5505 , \5506 );
nand \U$5165 ( \5508 , \1581 , \3388 );
nand \U$5166 ( \5509 , \5507 , \5508 );
not \U$5167 ( \5510 , \5509 );
or \U$5168 ( \5511 , \5504 , \5510 );
not \U$5169 ( \5512 , RIbb2ebc0_23);
not \U$5170 ( \5513 , \1510 );
or \U$5171 ( \5514 , \5512 , \5513 );
nand \U$5172 ( \5515 , \1511 , \3396 );
nand \U$5173 ( \5516 , \5514 , \5515 );
nand \U$5174 ( \5517 , \5516 , \3407 );
nand \U$5175 ( \5518 , \5511 , \5517 );
xor \U$5176 ( \5519 , \5503 , \5518 );
not \U$5177 ( \5520 , \1077 );
not \U$5178 ( \5521 , RIbb2f160_11);
not \U$5179 ( \5522 , \1113 );
or \U$5180 ( \5523 , \5521 , \5522 );
nand \U$5181 ( \5524 , \1114 , \1048 );
nand \U$5182 ( \5525 , \5523 , \5524 );
not \U$5183 ( \5526 , \5525 );
or \U$5184 ( \5527 , \5520 , \5526 );
nand \U$5185 ( \5528 , \5411 , \1011 );
nand \U$5186 ( \5529 , \5527 , \5528 );
xor \U$5187 ( \5530 , \5519 , \5529 );
xor \U$5188 ( \5531 , \5493 , \5530 );
xor \U$5189 ( \5532 , \5451 , \5531 );
not \U$5190 ( \5533 , \1294 );
not \U$5191 ( \5534 , \1290 );
not \U$5192 ( \5535 , \2224 );
or \U$5193 ( \5536 , \5534 , \5535 );
not \U$5194 ( \5537 , \1246 );
nand \U$5195 ( \5538 , \5537 , \2225 );
nand \U$5196 ( \5539 , \5536 , \5538 );
not \U$5197 ( \5540 , \5539 );
or \U$5198 ( \5541 , \5533 , \5540 );
and \U$5199 ( \5542 , \3517 , \1246 );
not \U$5200 ( \5543 , \3517 );
and \U$5201 ( \5544 , \5543 , \1289 );
or \U$5202 ( \5545 , \5542 , \5544 );
nand \U$5203 ( \5546 , \5545 , \1265 );
nand \U$5204 ( \5547 , \5541 , \5546 );
not \U$5205 ( \5548 , \1090 );
not \U$5206 ( \5549 , RIbb2f430_5);
not \U$5207 ( \5550 , \4450 );
not \U$5208 ( \5551 , \5550 );
or \U$5209 ( \5552 , \5549 , \5551 );
nand \U$5210 ( \5553 , \4450 , \1980 );
nand \U$5211 ( \5554 , \5552 , \5553 );
not \U$5212 ( \5555 , \5554 );
or \U$5213 ( \5556 , \5548 , \5555 );
not \U$5214 ( \5557 , RIbb2f430_5);
not \U$5215 ( \5558 , \1854 );
or \U$5216 ( \5559 , \5557 , \5558 );
nand \U$5217 ( \5560 , \3503 , \1085 );
nand \U$5218 ( \5561 , \5559 , \5560 );
nand \U$5219 ( \5562 , \5561 , \1147 );
nand \U$5220 ( \5563 , \5556 , \5562 );
xor \U$5221 ( \5564 , \5547 , \5563 );
not \U$5222 ( \5565 , \1445 );
not \U$5223 ( \5566 , \5461 );
or \U$5224 ( \5567 , \5565 , \5566 );
and \U$5225 ( \5568 , RIbb2ef80_15, \5130 );
not \U$5226 ( \5569 , RIbb2ef80_15);
and \U$5227 ( \5570 , \5569 , \1730 );
or \U$5228 ( \5571 , \5568 , \5570 );
nand \U$5229 ( \5572 , \5571 , \1517 );
nand \U$5230 ( \5573 , \5567 , \5572 );
xor \U$5231 ( \5574 , \5564 , \5573 );
not \U$5232 ( \5575 , \836 );
not \U$5233 ( \5576 , RIbb2ee90_17);
not \U$5234 ( \5577 , \1562 );
or \U$5235 ( \5578 , \5576 , \5577 );
nand \U$5236 ( \5579 , \1042 , \816 );
nand \U$5237 ( \5580 , \5578 , \5579 );
not \U$5238 ( \5581 , \5580 );
or \U$5239 ( \5582 , \5575 , \5581 );
and \U$5240 ( \5583 , \1550 , RIbb2ee90_17);
not \U$5241 ( \5584 , \1550 );
and \U$5242 ( \5585 , \5584 , \816 );
or \U$5243 ( \5586 , \5583 , \5585 );
nand \U$5244 ( \5587 , \5586 , \832 );
nand \U$5245 ( \5588 , \5582 , \5587 );
not \U$5246 ( \5589 , \1702 );
not \U$5247 ( \5590 , RIbb2f340_7);
not \U$5248 ( \5591 , \1340 );
or \U$5249 ( \5592 , \5590 , \5591 );
nand \U$5250 ( \5593 , \1339 , \2700 );
nand \U$5251 ( \5594 , \5592 , \5593 );
not \U$5252 ( \5595 , \5594 );
or \U$5253 ( \5596 , \5589 , \5595 );
not \U$5254 ( \5597 , RIbb2f340_7);
not \U$5255 ( \5598 , \2052 );
or \U$5256 ( \5599 , \5597 , \5598 );
nand \U$5257 ( \5600 , \1422 , \1692 );
nand \U$5258 ( \5601 , \5599 , \5600 );
nand \U$5259 ( \5602 , \5601 , \1737 );
nand \U$5260 ( \5603 , \5596 , \5602 );
xor \U$5261 ( \5604 , \5588 , \5603 );
not \U$5262 ( \5605 , \1533 );
not \U$5263 ( \5606 , RIbb2f250_9);
not \U$5264 ( \5607 , \1820 );
or \U$5265 ( \5608 , \5606 , \5607 );
nand \U$5266 ( \5609 , \1387 , \1566 );
nand \U$5267 ( \5610 , \5608 , \5609 );
not \U$5268 ( \5611 , \5610 );
or \U$5269 ( \5612 , \5605 , \5611 );
not \U$5270 ( \5613 , RIbb2f250_9);
not \U$5271 ( \5614 , \1171 );
or \U$5272 ( \5615 , \5613 , \5614 );
nand \U$5273 ( \5616 , \1248 , \1566 );
nand \U$5274 ( \5617 , \5615 , \5616 );
nand \U$5275 ( \5618 , \5617 , \1570 );
nand \U$5276 ( \5619 , \5612 , \5618 );
xor \U$5277 ( \5620 , \5604 , \5619 );
xor \U$5278 ( \5621 , \5574 , \5620 );
xor \U$5279 ( \5622 , \5380 , \5386 );
and \U$5280 ( \5623 , \5622 , \5391 );
and \U$5281 ( \5624 , \5380 , \5386 );
or \U$5282 ( \5625 , \5623 , \5624 );
xor \U$5283 ( \5626 , \5621 , \5625 );
xor \U$5284 ( \5627 , \5532 , \5626 );
not \U$5285 ( \5628 , \5314 );
or \U$5286 ( \5629 , \5628 , \5350 );
nand \U$5287 ( \5630 , \5629 , \5272 );
nand \U$5288 ( \5631 , \5350 , \5628 );
nand \U$5289 ( \5632 , \5630 , \5631 );
or \U$5290 ( \5633 , \3445 , \3465 );
nand \U$5291 ( \5634 , \5633 , RIbb2e9e0_27);
not \U$5292 ( \5635 , \2980 );
not \U$5293 ( \5636 , \5246 );
or \U$5294 ( \5637 , \5635 , \5636 );
not \U$5295 ( \5638 , \2251 );
and \U$5296 ( \5639 , RIbb2ead0_25, \5638 );
not \U$5297 ( \5640 , RIbb2ead0_25);
and \U$5298 ( \5641 , \5640 , \1775 );
or \U$5299 ( \5642 , \5639 , \5641 );
nand \U$5300 ( \5643 , \5642 , \2963 );
nand \U$5301 ( \5644 , \5637 , \5643 );
xor \U$5302 ( \5645 , \5634 , \5644 );
not \U$5303 ( \5646 , \2078 );
not \U$5304 ( \5647 , \5483 );
or \U$5305 ( \5648 , \5646 , \5647 );
nand \U$5306 ( \5649 , \5256 , \2077 );
nand \U$5307 ( \5650 , \5648 , \5649 );
xor \U$5308 ( \5651 , \5645 , \5650 );
not \U$5309 ( \5652 , \1090 );
not \U$5310 ( \5653 , \5321 );
or \U$5311 ( \5654 , \5652 , \5653 );
nand \U$5312 ( \5655 , \5554 , \1147 );
nand \U$5313 ( \5656 , \5654 , \5655 );
not \U$5314 ( \5657 , \1265 );
not \U$5315 ( \5658 , \5333 );
or \U$5316 ( \5659 , \5657 , \5658 );
nand \U$5317 ( \5660 , \5545 , \1294 );
nand \U$5318 ( \5661 , \5659 , \5660 );
xor \U$5319 ( \5662 , \5656 , \5661 );
not \U$5320 ( \5663 , \832 );
not \U$5321 ( \5664 , \5134 );
or \U$5322 ( \5665 , \5663 , \5664 );
nand \U$5323 ( \5666 , \5586 , \836 );
nand \U$5324 ( \5667 , \5665 , \5666 );
xor \U$5325 ( \5668 , \5662 , \5667 );
xor \U$5326 ( \5669 , \5651 , \5668 );
xor \U$5327 ( \5670 , \5452 , \5458 );
xor \U$5328 ( \5671 , \5670 , \5465 );
xor \U$5329 ( \5672 , \5669 , \5671 );
xor \U$5330 ( \5673 , \5632 , \5672 );
xor \U$5331 ( \5674 , \5206 , \5209 );
and \U$5332 ( \5675 , \5674 , \5216 );
and \U$5333 ( \5676 , \5206 , \5209 );
or \U$5334 ( \5677 , \5675 , \5676 );
not \U$5335 ( \5678 , \1737 );
not \U$5336 ( \5679 , \5594 );
or \U$5337 ( \5680 , \5678 , \5679 );
nand \U$5338 ( \5681 , \5123 , \1702 );
nand \U$5339 ( \5682 , \5680 , \5681 );
not \U$5340 ( \5683 , \3407 );
not \U$5341 ( \5684 , \5143 );
or \U$5342 ( \5685 , \5683 , \5684 );
nand \U$5343 ( \5686 , \5516 , \3383 );
nand \U$5344 ( \5687 , \5685 , \5686 );
xor \U$5345 ( \5688 , \5682 , \5687 );
not \U$5346 ( \5689 , \1570 );
not \U$5347 ( \5690 , \5610 );
or \U$5348 ( \5691 , \5689 , \5690 );
nand \U$5349 ( \5692 , \5290 , \1533 );
nand \U$5350 ( \5693 , \5691 , \5692 );
xor \U$5351 ( \5694 , \5688 , \5693 );
xor \U$5352 ( \5695 , \5677 , \5694 );
not \U$5353 ( \5696 , \5179 );
not \U$5354 ( \5697 , \5188 );
or \U$5355 ( \5698 , \5696 , \5697 );
nand \U$5356 ( \5699 , \5698 , \5174 );
nand \U$5357 ( \5700 , \5178 , \5187 );
nand \U$5358 ( \5701 , \5699 , \5700 );
xor \U$5359 ( \5702 , \5695 , \5701 );
and \U$5360 ( \5703 , \5673 , \5702 );
and \U$5361 ( \5704 , \5632 , \5672 );
or \U$5362 ( \5705 , \5703 , \5704 );
xor \U$5363 ( \5706 , \5627 , \5705 );
xor \U$5364 ( \5707 , \5677 , \5694 );
and \U$5365 ( \5708 , \5707 , \5701 );
and \U$5366 ( \5709 , \5677 , \5694 );
or \U$5367 ( \5710 , \5708 , \5709 );
not \U$5368 ( \5711 , \2980 );
not \U$5369 ( \5712 , \5642 );
or \U$5370 ( \5713 , \5711 , \5712 );
nand \U$5371 ( \5714 , \2963 , RIbb2ead0_25);
nand \U$5372 ( \5715 , \5713 , \5714 );
not \U$5373 ( \5716 , \5715 );
not \U$5374 ( \5717 , \998 );
not \U$5375 ( \5718 , RIbb2f070_13);
not \U$5376 ( \5719 , \1644 );
or \U$5377 ( \5720 , \5718 , \5719 );
nand \U$5378 ( \5721 , \1646 , \906 );
nand \U$5379 ( \5722 , \5720 , \5721 );
not \U$5380 ( \5723 , \5722 );
or \U$5381 ( \5724 , \5717 , \5723 );
not \U$5382 ( \5725 , \5419 );
nand \U$5383 ( \5726 , \5725 , \916 );
nand \U$5384 ( \5727 , \5724 , \5726 );
xor \U$5385 ( \5728 , \5716 , \5727 );
not \U$5386 ( \5729 , \5661 );
not \U$5387 ( \5730 , \5656 );
or \U$5388 ( \5731 , \5729 , \5730 );
or \U$5389 ( \5732 , \5656 , \5661 );
nand \U$5390 ( \5733 , \5732 , \5667 );
nand \U$5391 ( \5734 , \5731 , \5733 );
xor \U$5392 ( \5735 , \5728 , \5734 );
xor \U$5393 ( \5736 , \5634 , \5644 );
and \U$5394 ( \5737 , \5736 , \5650 );
and \U$5395 ( \5738 , \5634 , \5644 );
or \U$5396 ( \5739 , \5737 , \5738 );
not \U$5397 ( \5740 , \5693 );
not \U$5398 ( \5741 , \5682 );
or \U$5399 ( \5742 , \5740 , \5741 );
or \U$5400 ( \5743 , \5682 , \5693 );
nand \U$5401 ( \5744 , \5743 , \5687 );
nand \U$5402 ( \5745 , \5742 , \5744 );
xor \U$5403 ( \5746 , \5739 , \5745 );
not \U$5404 ( \5747 , \5424 );
not \U$5405 ( \5748 , \5747 );
not \U$5406 ( \5749 , \5415 );
or \U$5407 ( \5750 , \5748 , \5749 );
or \U$5408 ( \5751 , \5747 , \5415 );
nand \U$5409 ( \5752 , \5751 , \5435 );
nand \U$5410 ( \5753 , \5750 , \5752 );
xor \U$5411 ( \5754 , \5746 , \5753 );
xor \U$5412 ( \5755 , \5735 , \5754 );
xor \U$5413 ( \5756 , \5651 , \5668 );
and \U$5414 ( \5757 , \5756 , \5671 );
and \U$5415 ( \5758 , \5651 , \5668 );
or \U$5416 ( \5759 , \5757 , \5758 );
xor \U$5417 ( \5760 , \5755 , \5759 );
xor \U$5418 ( \5761 , \5710 , \5760 );
xor \U$5419 ( \5762 , \5379 , \5392 );
and \U$5420 ( \5763 , \5762 , \5437 );
and \U$5421 ( \5764 , \5379 , \5392 );
or \U$5422 ( \5765 , \5763 , \5764 );
xor \U$5423 ( \5766 , \5761 , \5765 );
xor \U$5424 ( \5767 , \5706 , \5766 );
xor \U$5425 ( \5768 , \5447 , \5767 );
not \U$5426 ( \5769 , \5158 );
not \U$5427 ( \5770 , \5220 );
or \U$5428 ( \5771 , \5769 , \5770 );
not \U$5429 ( \5772 , \5158 );
nand \U$5430 ( \5773 , \5772 , \5219 );
nand \U$5431 ( \5774 , \5773 , \5162 );
nand \U$5432 ( \5775 , \5771 , \5774 );
xor \U$5433 ( \5776 , \5632 , \5672 );
xor \U$5434 ( \5777 , \5776 , \5702 );
nand \U$5435 ( \5778 , \5775 , \5777 );
or \U$5436 ( \5779 , \5775 , \5777 );
not \U$5437 ( \5780 , \5239 );
not \U$5438 ( \5781 , \5352 );
or \U$5439 ( \5782 , \5780 , \5781 );
nand \U$5440 ( \5783 , \5351 , \5240 );
nand \U$5441 ( \5784 , \5783 , \5360 );
nand \U$5442 ( \5785 , \5782 , \5784 );
nand \U$5443 ( \5786 , \5779 , \5785 );
nand \U$5444 ( \5787 , \5778 , \5786 );
xor \U$5445 ( \5788 , \5768 , \5787 );
not \U$5446 ( \5789 , \5777 );
and \U$5447 ( \5790 , \5785 , \5789 );
not \U$5448 ( \5791 , \5785 );
and \U$5449 ( \5792 , \5791 , \5777 );
nor \U$5450 ( \5793 , \5790 , \5792 );
not \U$5451 ( \5794 , \5793 );
not \U$5452 ( \5795 , \5775 );
and \U$5453 ( \5796 , \5794 , \5795 );
and \U$5454 ( \5797 , \5775 , \5793 );
nor \U$5455 ( \5798 , \5796 , \5797 );
not \U$5456 ( \5799 , \5798 );
xor \U$5457 ( \5800 , \5375 , \5438 );
xor \U$5458 ( \5801 , \5800 , \5444 );
or \U$5459 ( \5802 , \5799 , \5801 );
not \U$5460 ( \5803 , \5235 );
nand \U$5461 ( \5804 , \5803 , \5365 );
not \U$5462 ( \5805 , \5804 );
not \U$5463 ( \5806 , \5231 );
or \U$5464 ( \5807 , \5805 , \5806 );
not \U$5465 ( \5808 , \5365 );
nand \U$5466 ( \5809 , \5808 , \5235 );
nand \U$5467 ( \5810 , \5807 , \5809 );
nand \U$5468 ( \5811 , \5802 , \5810 );
nand \U$5469 ( \5812 , \5799 , \5801 );
nand \U$5470 ( \5813 , \5811 , \5812 );
or \U$5471 ( \5814 , \5788 , \5813 );
xor \U$5472 ( \5815 , \5801 , \5798 );
xor \U$5473 ( \5816 , \5815 , \5810 );
xor \U$5474 ( \5817 , \5221 , \5226 );
and \U$5475 ( \5818 , \5817 , \5368 );
and \U$5476 ( \5819 , \5221 , \5226 );
or \U$5477 ( \5820 , \5818 , \5819 );
nand \U$5478 ( \5821 , \5816 , \5820 );
nand \U$5479 ( \5822 , \5814 , \5821 );
nor \U$5480 ( \5823 , \5371 , \5822 );
not \U$5481 ( \5824 , \5823 );
xor \U$5482 ( \5825 , \4829 , \4846 );
xor \U$5483 ( \5826 , \5825 , \4854 );
xor \U$5484 ( \5827 , \4533 , \4520 );
xor \U$5485 ( \5828 , \5827 , \4530 );
xor \U$5486 ( \5829 , \5826 , \5828 );
xor \U$5487 ( \5830 , \4614 , \4602 );
xor \U$5488 ( \5831 , \5830 , \4627 );
xor \U$5489 ( \5832 , \4575 , \4564 );
xnor \U$5490 ( \5833 , \5832 , \4588 );
not \U$5491 ( \5834 , \5833 );
or \U$5492 ( \5835 , \5831 , \5834 );
not \U$5493 ( \5836 , \4712 );
not \U$5494 ( \5837 , RIbb2e620_35);
not \U$5495 ( \5838 , \814 );
or \U$5496 ( \5839 , \5837 , \5838 );
not \U$5497 ( \5840 , RIbb2e620_35);
nand \U$5498 ( \5841 , \2251 , \5840 );
nand \U$5499 ( \5842 , \5839 , \5841 );
not \U$5500 ( \5843 , \5842 );
or \U$5501 ( \5844 , \5836 , \5843 );
buf \U$5502 ( \5845 , \4714 );
nand \U$5503 ( \5846 , \5845 , RIbb2e620_35);
nand \U$5504 ( \5847 , \5844 , \5846 );
not \U$5505 ( \5848 , \1737 );
not \U$5506 ( \5849 , \3909 );
or \U$5507 ( \5850 , \5848 , \5849 );
not \U$5508 ( \5851 , RIbb2f340_7);
not \U$5509 ( \5852 , \3655 );
or \U$5510 ( \5853 , \5851 , \5852 );
nand \U$5511 ( \5854 , \3654 , \1734 );
nand \U$5512 ( \5855 , \5853 , \5854 );
nand \U$5513 ( \5856 , \5855 , \1702 );
nand \U$5514 ( \5857 , \5850 , \5856 );
xor \U$5515 ( \5858 , \5847 , \5857 );
not \U$5516 ( \5859 , \4718 );
nor \U$5517 ( \5860 , \5859 , \4732 );
not \U$5518 ( \5861 , \5860 );
not \U$5519 ( \5862 , \4729 );
and \U$5520 ( \5863 , \5861 , \5862 );
and \U$5521 ( \5864 , \5860 , \4729 );
nor \U$5522 ( \5865 , \5863 , \5864 );
xor \U$5523 ( \5866 , \5858 , \5865 );
nand \U$5524 ( \5867 , \5835 , \5866 );
nand \U$5525 ( \5868 , \5831 , \5834 );
nand \U$5526 ( \5869 , \5867 , \5868 );
xor \U$5527 ( \5870 , \4522 , \4524 );
xor \U$5528 ( \5871 , \5870 , \4527 );
xor \U$5529 ( \5872 , \5869 , \5871 );
not \U$5530 ( \5873 , \4837 );
not \U$5531 ( \5874 , \4841 );
or \U$5532 ( \5875 , \5873 , \5874 );
or \U$5533 ( \5876 , \4837 , \4841 );
nand \U$5534 ( \5877 , \5875 , \5876 );
and \U$5535 ( \5878 , \5877 , \4844 );
not \U$5536 ( \5879 , \5877 );
and \U$5537 ( \5880 , \5879 , \4831 );
nor \U$5538 ( \5881 , \5878 , \5880 );
and \U$5539 ( \5882 , \5872 , \5881 );
and \U$5540 ( \5883 , \5869 , \5871 );
or \U$5541 ( \5884 , \5882 , \5883 );
and \U$5542 ( \5885 , \5829 , \5884 );
and \U$5543 ( \5886 , \5826 , \5828 );
or \U$5544 ( \5887 , \5885 , \5886 );
not \U$5545 ( \5888 , \2922 );
not \U$5546 ( \5889 , RIbb2e8f0_29);
not \U$5547 ( \5890 , \4595 );
or \U$5548 ( \5891 , \5889 , \5890 );
nand \U$5549 ( \5892 , \1563 , \3265 );
nand \U$5550 ( \5893 , \5891 , \5892 );
not \U$5551 ( \5894 , \5893 );
or \U$5552 ( \5895 , \5888 , \5894 );
not \U$5553 ( \5896 , RIbb2e8f0_29);
not \U$5554 ( \5897 , \4284 );
or \U$5555 ( \5898 , \5896 , \5897 );
nand \U$5556 ( \5899 , \1071 , \3440 );
nand \U$5557 ( \5900 , \5898 , \5899 );
nand \U$5558 ( \5901 , \5900 , \2925 );
nand \U$5559 ( \5902 , \5895 , \5901 );
not \U$5560 ( \5903 , \5902 );
not \U$5561 ( \5904 , \2940 );
not \U$5562 ( \5905 , RIbb2e800_31);
not \U$5563 ( \5906 , \2399 );
or \U$5564 ( \5907 , \5905 , \5906 );
nand \U$5565 ( \5908 , \957 , \2917 );
nand \U$5566 ( \5909 , \5907 , \5908 );
not \U$5567 ( \5910 , \5909 );
or \U$5568 ( \5911 , \5904 , \5910 );
not \U$5569 ( \5912 , RIbb2e800_31);
not \U$5570 ( \5913 , \988 );
or \U$5571 ( \5914 , \5912 , \5913 );
nand \U$5572 ( \5915 , \987 , \2917 );
nand \U$5573 ( \5916 , \5914 , \5915 );
nand \U$5574 ( \5917 , \5916 , \2941 );
nand \U$5575 ( \5918 , \5911 , \5917 );
not \U$5576 ( \5919 , \5918 );
or \U$5577 ( \5920 , \5903 , \5919 );
or \U$5578 ( \5921 , \5918 , \5902 );
not \U$5579 ( \5922 , \853 );
not \U$5580 ( \5923 , RIbb2eda0_19);
not \U$5581 ( \5924 , \3822 );
or \U$5582 ( \5925 , \5923 , \5924 );
nand \U$5583 ( \5926 , \1422 , \1776 );
nand \U$5584 ( \5927 , \5925 , \5926 );
not \U$5585 ( \5928 , \5927 );
or \U$5586 ( \5929 , \5922 , \5928 );
not \U$5587 ( \5930 , RIbb2eda0_19);
not \U$5588 ( \5931 , \3116 );
or \U$5589 ( \5932 , \5930 , \5931 );
nand \U$5590 ( \5933 , \4340 , \1776 );
nand \U$5591 ( \5934 , \5932 , \5933 );
nand \U$5592 ( \5935 , \5934 , \855 );
nand \U$5593 ( \5936 , \5929 , \5935 );
nand \U$5594 ( \5937 , \5921 , \5936 );
nand \U$5595 ( \5938 , \5920 , \5937 );
nor \U$5596 ( \5939 , \4355 , \523 );
not \U$5597 ( \5940 , \5939 );
buf \U$5598 ( \5941 , \4360 );
not \U$5599 ( \5942 , \5941 );
or \U$5600 ( \5943 , \5940 , \5942 );
and \U$5601 ( \5944 , \4370 , \524 );
nor \U$5602 ( \5945 , \5944 , \4374 );
nand \U$5603 ( \5946 , \5943 , \5945 );
not \U$5604 ( \5947 , \528 );
nand \U$5605 ( \5948 , \5947 , \633 );
not \U$5606 ( \5949 , \5948 );
and \U$5607 ( \5950 , \5946 , \5949 );
not \U$5608 ( \5951 , \5946 );
and \U$5609 ( \5952 , \5951 , \5948 );
nor \U$5610 ( \5953 , \5950 , \5952 );
buf \U$5611 ( \5954 , \5953 );
buf \U$5612 ( \5955 , \5954 );
not \U$5613 ( \5956 , \5955 );
not \U$5614 ( \5957 , \5956 );
and \U$5615 ( \5958 , \1313 , \5957 );
not \U$5616 ( \5959 , \5958 );
not \U$5617 ( \5960 , \1737 );
not \U$5618 ( \5961 , RIbb2f340_7);
not \U$5619 ( \5962 , \4020 );
not \U$5620 ( \5963 , \5962 );
or \U$5621 ( \5964 , \5961 , \5963 );
nand \U$5622 ( \5965 , \3024 , \1734 );
nand \U$5623 ( \5966 , \5964 , \5965 );
not \U$5624 ( \5967 , \5966 );
or \U$5625 ( \5968 , \5960 , \5967 );
not \U$5626 ( \5969 , RIbb2f340_7);
not \U$5627 ( \5970 , \3045 );
or \U$5628 ( \5971 , \5969 , \5970 );
nand \U$5629 ( \5972 , \4030 , \1734 );
nand \U$5630 ( \5973 , \5971 , \5972 );
nand \U$5631 ( \5974 , \5973 , \1702 );
nand \U$5632 ( \5975 , \5968 , \5974 );
not \U$5633 ( \5976 , \5975 );
or \U$5634 ( \5977 , \5959 , \5976 );
or \U$5635 ( \5978 , \5975 , \5958 );
not \U$5636 ( \5979 , \3407 );
not \U$5637 ( \5980 , RIbb2ebc0_23);
not \U$5638 ( \5981 , \3066 );
or \U$5639 ( \5982 , \5980 , \5981 );
nand \U$5640 ( \5983 , \1114 , \2073 );
nand \U$5641 ( \5984 , \5982 , \5983 );
not \U$5642 ( \5985 , \5984 );
or \U$5643 ( \5986 , \5979 , \5985 );
not \U$5644 ( \5987 , RIbb2ebc0_23);
not \U$5645 ( \5988 , \1138 );
not \U$5646 ( \5989 , \5988 );
or \U$5647 ( \5990 , \5987 , \5989 );
nand \U$5648 ( \5991 , \1138 , \3388 );
nand \U$5649 ( \5992 , \5990 , \5991 );
nand \U$5650 ( \5993 , \5992 , \3383 );
nand \U$5651 ( \5994 , \5986 , \5993 );
nand \U$5652 ( \5995 , \5978 , \5994 );
nand \U$5653 ( \5996 , \5977 , \5995 );
nor \U$5654 ( \5997 , \5938 , \5996 );
not \U$5655 ( \5998 , \4712 );
not \U$5656 ( \5999 , RIbb2e620_35);
not \U$5657 ( \6000 , \1579 );
or \U$5658 ( \6001 , \5999 , \6000 );
not \U$5659 ( \6002 , RIbb2e620_35);
nand \U$5660 ( \6003 , \1580 , \6002 );
nand \U$5661 ( \6004 , \6001 , \6003 );
not \U$5662 ( \6005 , \6004 );
or \U$5663 ( \6006 , \5998 , \6005 );
nand \U$5664 ( \6007 , \5842 , \5845 );
nand \U$5665 ( \6008 , \6006 , \6007 );
not \U$5666 ( \6009 , \1090 );
not \U$5667 ( \6010 , RIbb2f430_5);
not \U$5668 ( \6011 , \4040 );
or \U$5669 ( \6012 , \6010 , \6011 );
not \U$5670 ( \6013 , \4749 );
nand \U$5671 ( \6014 , \6013 , \1980 );
nand \U$5672 ( \6015 , \6012 , \6014 );
not \U$5673 ( \6016 , \6015 );
or \U$5674 ( \6017 , \6009 , \6016 );
not \U$5675 ( \6018 , RIbb2f430_5);
not \U$5676 ( \6019 , \4411 );
or \U$5677 ( \6020 , \6018 , \6019 );
not \U$5678 ( \6021 , \3276 );
nand \U$5679 ( \6022 , \6021 , \1647 );
nand \U$5680 ( \6023 , \6020 , \6022 );
nand \U$5681 ( \6024 , \6023 , \1147 );
nand \U$5682 ( \6025 , \6017 , \6024 );
or \U$5683 ( \6026 , \6008 , \6025 );
not \U$5684 ( \6027 , \2077 );
not \U$5685 ( \6028 , RIbb2ecb0_21);
not \U$5686 ( \6029 , \1170 );
or \U$5687 ( \6030 , \6028 , \6029 );
nand \U$5688 ( \6031 , \3736 , \5481 );
nand \U$5689 ( \6032 , \6030 , \6031 );
not \U$5690 ( \6033 , \6032 );
or \U$5691 ( \6034 , \6027 , \6033 );
not \U$5692 ( \6035 , RIbb2ecb0_21);
not \U$5693 ( \6036 , \1284 );
or \U$5694 ( \6037 , \6035 , \6036 );
nand \U$5695 ( \6038 , \1283 , \2249 );
nand \U$5696 ( \6039 , \6037 , \6038 );
nand \U$5697 ( \6040 , \6039 , \2078 );
nand \U$5698 ( \6041 , \6034 , \6040 );
nand \U$5699 ( \6042 , \6026 , \6041 );
nand \U$5700 ( \6043 , \6008 , \6025 );
nand \U$5701 ( \6044 , \6042 , \6043 );
not \U$5702 ( \6045 , \6044 );
or \U$5703 ( \6046 , \5997 , \6045 );
nand \U$5704 ( \6047 , \5938 , \5996 );
nand \U$5705 ( \6048 , \6046 , \6047 );
not \U$5706 ( \6049 , \6048 );
and \U$5707 ( \6050 , \1476 , \3864 );
not \U$5708 ( \6051 , \1476 );
and \U$5709 ( \6052 , \6051 , RIbb2e710_33);
or \U$5710 ( \6053 , \6050 , \6052 );
and \U$5711 ( \6054 , \6053 , \3887 );
not \U$5712 ( \6055 , RIbb2e710_33);
not \U$5713 ( \6056 , \3262 );
or \U$5714 ( \6057 , \6055 , \6056 );
not \U$5715 ( \6058 , RIbb2e710_33);
nand \U$5716 ( \6059 , \4315 , \6058 );
nand \U$5717 ( \6060 , \6057 , \6059 );
and \U$5718 ( \6061 , \6060 , \4791 );
nor \U$5719 ( \6062 , \6054 , \6061 );
not \U$5720 ( \6063 , \6062 );
not \U$5721 ( \6064 , \6063 );
not \U$5722 ( \6065 , RIbb2e9e0_27);
and \U$5723 ( \6066 , \6065 , \3480 );
not \U$5724 ( \6067 , \6065 );
and \U$5725 ( \6068 , \6067 , \5130 );
nor \U$5726 ( \6069 , \6066 , \6068 );
not \U$5727 ( \6070 , \6069 );
not \U$5728 ( \6071 , \3445 );
not \U$5729 ( \6072 , \6071 );
and \U$5730 ( \6073 , \6070 , \6072 );
not \U$5731 ( \6074 , \3465 );
and \U$5732 ( \6075 , \4598 , \1548 );
not \U$5733 ( \6076 , \4598 );
and \U$5734 ( \6077 , \6076 , \5003 );
nor \U$5735 ( \6078 , \6075 , \6077 );
nor \U$5736 ( \6079 , \6074 , \6078 );
nor \U$5737 ( \6080 , \6073 , \6079 );
not \U$5738 ( \6081 , \6080 );
not \U$5739 ( \6082 , \6081 );
or \U$5740 ( \6083 , \6064 , \6082 );
not \U$5741 ( \6084 , \6062 );
not \U$5742 ( \6085 , \6080 );
or \U$5743 ( \6086 , \6084 , \6085 );
not \U$5744 ( \6087 , \832 );
not \U$5745 ( \6088 , RIbb2ee90_17);
not \U$5746 ( \6089 , \3807 );
or \U$5747 ( \6090 , \6088 , \6089 );
nand \U$5748 ( \6091 , \3503 , \822 );
nand \U$5749 ( \6092 , \6090 , \6091 );
not \U$5750 ( \6093 , \6092 );
or \U$5751 ( \6094 , \6087 , \6093 );
not \U$5752 ( \6095 , \1337 );
not \U$5753 ( \6096 , \6095 );
not \U$5754 ( \6097 , \6096 );
and \U$5755 ( \6098 , \6097 , RIbb2ee90_17);
not \U$5756 ( \6099 , \6097 );
and \U$5757 ( \6100 , \6099 , \3057 );
or \U$5758 ( \6101 , \6098 , \6100 );
nand \U$5759 ( \6102 , \6101 , \836 );
nand \U$5760 ( \6103 , \6094 , \6102 );
nand \U$5761 ( \6104 , \6086 , \6103 );
nand \U$5762 ( \6105 , \6083 , \6104 );
not \U$5763 ( \6106 , \6105 );
not \U$5764 ( \6107 , \3166 );
not \U$5765 ( \6108 , \6107 );
not \U$5766 ( \6109 , \6108 );
not \U$5767 ( \6110 , \906 );
and \U$5768 ( \6111 , \6109 , \6110 );
and \U$5769 ( \6112 , \3167 , \1656 );
nor \U$5770 ( \6113 , \6111 , \6112 );
not \U$5771 ( \6114 , \6113 );
not \U$5772 ( \6115 , \1654 );
and \U$5773 ( \6116 , \6114 , \6115 );
not \U$5774 ( \6117 , RIbb2f070_13);
not \U$5775 ( \6118 , \3342 );
or \U$5776 ( \6119 , \6117 , \6118 );
not \U$5777 ( \6120 , \3517 );
nand \U$5778 ( \6121 , \6120 , \3421 );
nand \U$5779 ( \6122 , \6119 , \6121 );
and \U$5780 ( \6123 , \6122 , \998 );
nor \U$5781 ( \6124 , \6116 , \6123 );
not \U$5782 ( \6125 , \6124 );
and \U$5783 ( \6126 , RIbb2ead0_25, \3243 );
not \U$5784 ( \6127 , RIbb2ead0_25);
and \U$5785 ( \6128 , \6127 , \3239 );
or \U$5786 ( \6129 , \6126 , \6128 );
not \U$5787 ( \6130 , \6129 );
not \U$5788 ( \6131 , \2980 );
not \U$5789 ( \6132 , \6131 );
and \U$5790 ( \6133 , \6130 , \6132 );
xor \U$5791 ( \6134 , RIbb2ead0_25, \3364 );
and \U$5792 ( \6135 , \6134 , \2963 );
nor \U$5793 ( \6136 , \6133 , \6135 );
not \U$5794 ( \6137 , \6136 );
or \U$5795 ( \6138 , \6125 , \6137 );
not \U$5796 ( \6139 , \3105 );
and \U$5797 ( \6140 , RIbb2ef80_15, \5550 );
not \U$5798 ( \6141 , RIbb2ef80_15);
and \U$5799 ( \6142 , \6141 , \4450 );
or \U$5800 ( \6143 , \6140 , \6142 );
not \U$5801 ( \6144 , \6143 );
or \U$5802 ( \6145 , \6139 , \6144 );
and \U$5803 ( \6146 , RIbb2ef80_15, \2224 );
not \U$5804 ( \6147 , RIbb2ef80_15);
and \U$5805 ( \6148 , \6147 , \2225 );
or \U$5806 ( \6149 , \6146 , \6148 );
nand \U$5807 ( \6150 , \6149 , \1445 );
nand \U$5808 ( \6151 , \6145 , \6150 );
nand \U$5809 ( \6152 , \6138 , \6151 );
not \U$5810 ( \6153 , \6136 );
not \U$5811 ( \6154 , \6124 );
nand \U$5812 ( \6155 , \6153 , \6154 );
nand \U$5813 ( \6156 , \6152 , \6155 );
not \U$5814 ( \6157 , \6156 );
nand \U$5815 ( \6158 , \6106 , \6157 );
not \U$5816 ( \6159 , \6158 );
not \U$5817 ( \6160 , \1702 );
not \U$5818 ( \6161 , \5966 );
or \U$5819 ( \6162 , \6160 , \6161 );
nand \U$5820 ( \6163 , \5855 , \1737 );
nand \U$5821 ( \6164 , \6162 , \6163 );
not \U$5822 ( \6165 , \1570 );
not \U$5823 ( \6166 , \4642 );
or \U$5824 ( \6167 , \6165 , \6166 );
not \U$5825 ( \6168 , RIbb2f250_9);
not \U$5826 ( \6169 , \3226 );
or \U$5827 ( \6170 , \6168 , \6169 );
buf \U$5828 ( \6171 , \3223 );
not \U$5829 ( \6172 , \6171 );
buf \U$5830 ( \6173 , \6172 );
not \U$5831 ( \6174 , \6173 );
nand \U$5832 ( \6175 , \6174 , \5064 );
nand \U$5833 ( \6176 , \6170 , \6175 );
nand \U$5834 ( \6177 , \6176 , \1533 );
nand \U$5835 ( \6178 , \6167 , \6177 );
xor \U$5836 ( \6179 , \6164 , \6178 );
not \U$5837 ( \6180 , \3406 );
not \U$5838 ( \6181 , \5992 );
or \U$5839 ( \6182 , \6180 , \6181 );
nand \U$5840 ( \6183 , \4666 , \3383 );
nand \U$5841 ( \6184 , \6182 , \6183 );
not \U$5842 ( \6185 , \6184 );
xnor \U$5843 ( \6186 , \6179 , \6185 );
not \U$5844 ( \6187 , \6186 );
or \U$5845 ( \6188 , \6159 , \6187 );
nand \U$5846 ( \6189 , \6156 , \6105 );
nand \U$5847 ( \6190 , \6188 , \6189 );
not \U$5848 ( \6191 , \6190 );
or \U$5849 ( \6192 , \6049 , \6191 );
or \U$5850 ( \6193 , \6048 , \6190 );
not \U$5851 ( \6194 , \5847 );
not \U$5852 ( \6195 , \1376 );
not \U$5853 ( \6196 , \1394 );
not \U$5854 ( \6197 , \4695 );
not \U$5855 ( \6198 , \6197 );
not \U$5856 ( \6199 , \6198 );
not \U$5857 ( \6200 , \6199 );
or \U$5858 ( \6201 , \6196 , \6200 );
buf \U$5859 ( \6202 , \6198 );
nand \U$5860 ( \6203 , \6202 , \1392 );
nand \U$5861 ( \6204 , \6201 , \6203 );
not \U$5862 ( \6205 , \6204 );
or \U$5863 ( \6206 , \6195 , \6205 );
not \U$5864 ( \6207 , \1429 );
not \U$5865 ( \6208 , \6207 );
nand \U$5866 ( \6209 , \524 , \5947 );
nor \U$5867 ( \6210 , \6209 , \4355 );
not \U$5868 ( \6211 , \6210 );
not \U$5869 ( \6212 , \5941 );
or \U$5870 ( \6213 , \6211 , \6212 );
not \U$5871 ( \6214 , \6209 );
and \U$5872 ( \6215 , \4370 , \6214 );
not \U$5873 ( \6216 , \5947 );
not \U$5874 ( \6217 , \4374 );
or \U$5875 ( \6218 , \6216 , \6217 );
nand \U$5876 ( \6219 , \6218 , \633 );
nor \U$5877 ( \6220 , \6215 , \6219 );
nand \U$5878 ( \6221 , \6213 , \6220 );
not \U$5879 ( \6222 , \635 );
nor \U$5880 ( \6223 , \6222 , \632 );
and \U$5881 ( \6224 , \6221 , \6223 );
not \U$5882 ( \6225 , \6221 );
not \U$5883 ( \6226 , \6223 );
and \U$5884 ( \6227 , \6225 , \6226 );
nor \U$5885 ( \6228 , \6224 , \6227 );
buf \U$5886 ( \6229 , \6228 );
not \U$5887 ( \6230 , \6229 );
buf \U$5888 ( \6231 , \6230 );
not \U$5889 ( \6232 , \6231 );
xor \U$5890 ( \6233 , \1393 , \6232 );
nand \U$5891 ( \6234 , \6208 , \6233 );
nand \U$5892 ( \6235 , \6206 , \6234 );
and \U$5893 ( \6236 , RIbb2e440_39, RIbb2e4b8_38);
not \U$5894 ( \6237 , RIbb2e440_39);
not \U$5895 ( \6238 , RIbb2e4b8_38);
and \U$5896 ( \6239 , \6237 , \6238 );
nor \U$5897 ( \6240 , \6236 , \6239 );
buf \U$5898 ( \6241 , \6240 );
buf \U$5899 ( \6242 , \6241 );
not \U$5900 ( \6243 , \6242 );
not \U$5901 ( \6244 , \6243 );
not \U$5902 ( \6245 , \6240 );
not \U$5903 ( \6246 , RIbb2e530_37);
and \U$5904 ( \6247 , \6246 , \6238 );
and \U$5905 ( \6248 , RIbb2e530_37, RIbb2e4b8_38);
nor \U$5906 ( \6249 , \6247 , \6248 );
and \U$5907 ( \6250 , \6245 , \6249 );
buf \U$5908 ( \6251 , \6250 );
not \U$5909 ( \6252 , \6251 );
not \U$5910 ( \6253 , \6252 );
or \U$5911 ( \6254 , \6244 , \6253 );
nand \U$5912 ( \6255 , \6254 , RIbb2e530_37);
or \U$5913 ( \6256 , \6235 , \6255 );
not \U$5914 ( \6257 , \1294 );
not \U$5915 ( \6258 , \1246 );
not \U$5916 ( \6259 , \4325 );
or \U$5917 ( \6260 , \6258 , \6259 );
nand \U$5918 ( \6261 , \4089 , \1245 );
nand \U$5919 ( \6262 , \6260 , \6261 );
not \U$5920 ( \6263 , \6262 );
or \U$5921 ( \6264 , \6257 , \6263 );
not \U$5922 ( \6265 , \1290 );
not \U$5923 ( \6266 , \4393 );
or \U$5924 ( \6267 , \6265 , \6266 );
not \U$5925 ( \6268 , \4390 );
not \U$5926 ( \6269 , \6268 );
nand \U$5927 ( \6270 , \6269 , \1245 );
nand \U$5928 ( \6271 , \6267 , \6270 );
nand \U$5929 ( \6272 , \6271 , \1265 );
nand \U$5930 ( \6273 , \6264 , \6272 );
nand \U$5931 ( \6274 , \6256 , \6273 );
nand \U$5932 ( \6275 , \6235 , \6255 );
nand \U$5933 ( \6276 , \6274 , \6275 );
xor \U$5934 ( \6277 , \6194 , \6276 );
and \U$5935 ( \6278 , \1393 , \6232 );
not \U$5936 ( \6279 , \1429 );
not \U$5937 ( \6280 , \6204 );
or \U$5938 ( \6281 , \6279 , \6280 );
nand \U$5939 ( \6282 , \4727 , \1376 );
nand \U$5940 ( \6283 , \6281 , \6282 );
xor \U$5941 ( \6284 , \6278 , \6283 );
not \U$5942 ( \6285 , \2077 );
not \U$5943 ( \6286 , \6039 );
or \U$5944 ( \6287 , \6285 , \6286 );
nand \U$5945 ( \6288 , \4772 , \2078 );
nand \U$5946 ( \6289 , \6287 , \6288 );
xor \U$5947 ( \6290 , \6284 , \6289 );
and \U$5948 ( \6291 , \6277 , \6290 );
and \U$5949 ( \6292 , \6194 , \6276 );
or \U$5950 ( \6293 , \6291 , \6292 );
nand \U$5951 ( \6294 , \6193 , \6293 );
nand \U$5952 ( \6295 , \6192 , \6294 );
and \U$5953 ( \6296 , \6134 , \2980 );
and \U$5954 ( \6297 , \4584 , \2963 );
nor \U$5955 ( \6298 , \6296 , \6297 );
not \U$5956 ( \6299 , \1011 );
not \U$5957 ( \6300 , RIbb2f160_11);
not \U$5958 ( \6301 , \3146 );
not \U$5959 ( \6302 , \6301 );
or \U$5960 ( \6303 , \6300 , \6302 );
nand \U$5961 ( \6304 , \3142 , \1805 );
nand \U$5962 ( \6305 , \6303 , \6304 );
not \U$5963 ( \6306 , \6305 );
or \U$5964 ( \6307 , \6299 , \6306 );
nand \U$5965 ( \6308 , \4653 , \1077 );
nand \U$5966 ( \6309 , \6307 , \6308 );
not \U$5967 ( \6310 , \916 );
not \U$5968 ( \6311 , \6122 );
or \U$5969 ( \6312 , \6310 , \6311 );
nand \U$5970 ( \6313 , \4573 , \998 );
nand \U$5971 ( \6314 , \6312 , \6313 );
nor \U$5972 ( \6315 , \6309 , \6314 );
or \U$5973 ( \6316 , \6298 , \6315 );
nand \U$5974 ( \6317 , \6309 , \6314 );
nand \U$5975 ( \6318 , \6316 , \6317 );
not \U$5976 ( \6319 , \836 );
not \U$5977 ( \6320 , \4625 );
or \U$5978 ( \6321 , \6319 , \6320 );
nand \U$5979 ( \6322 , \6101 , \832 );
nand \U$5980 ( \6323 , \6321 , \6322 );
not \U$5981 ( \6324 , \2940 );
not \U$5982 ( \6325 , \5916 );
or \U$5983 ( \6326 , \6324 , \6325 );
nand \U$5984 ( \6327 , \4560 , \2941 );
nand \U$5985 ( \6328 , \6326 , \6327 );
or \U$5986 ( \6329 , \6323 , \6328 );
not \U$5987 ( \6330 , \1445 );
not \U$5988 ( \6331 , \6143 );
or \U$5989 ( \6332 , \6330 , \6331 );
nand \U$5990 ( \6333 , \4612 , \1517 );
nand \U$5991 ( \6334 , \6332 , \6333 );
nand \U$5992 ( \6335 , \6329 , \6334 );
nand \U$5993 ( \6336 , \6323 , \6328 );
nand \U$5994 ( \6337 , \6335 , \6336 );
xor \U$5995 ( \6338 , \6318 , \6337 );
nor \U$5996 ( \6339 , \6178 , \6164 );
or \U$5997 ( \6340 , \6339 , \6185 );
nand \U$5998 ( \6341 , \6178 , \6164 );
nand \U$5999 ( \6342 , \6340 , \6341 );
xor \U$6000 ( \6343 , \6338 , \6342 );
not \U$6001 ( \6344 , \6343 );
not \U$6002 ( \6345 , \855 );
not \U$6003 ( \6346 , \4813 );
or \U$6004 ( \6347 , \6345 , \6346 );
nand \U$6005 ( \6348 , \5934 , \853 );
nand \U$6006 ( \6349 , \6347 , \6348 );
not \U$6007 ( \6350 , \2922 );
not \U$6008 ( \6351 , \5900 );
or \U$6009 ( \6352 , \6350 , \6351 );
nand \U$6010 ( \6353 , \4802 , \2925 );
nand \U$6011 ( \6354 , \6352 , \6353 );
not \U$6012 ( \6355 , \6354 );
xor \U$6013 ( \6356 , \6349 , \6355 );
not \U$6014 ( \6357 , \3445 );
not \U$6015 ( \6358 , \6078 );
not \U$6016 ( \6359 , \6358 );
or \U$6017 ( \6360 , \6357 , \6359 );
nand \U$6018 ( \6361 , \4600 , \3465 );
nand \U$6019 ( \6362 , \6360 , \6361 );
xor \U$6020 ( \6363 , \6356 , \6362 );
not \U$6021 ( \6364 , \6363 );
not \U$6022 ( \6365 , \6364 );
not \U$6023 ( \6366 , \1294 );
not \U$6024 ( \6367 , \4755 );
or \U$6025 ( \6368 , \6366 , \6367 );
nand \U$6026 ( \6369 , \6262 , \1265 );
nand \U$6027 ( \6370 , \6368 , \6369 );
not \U$6028 ( \6371 , \6370 );
not \U$6029 ( \6372 , \3887 );
not \U$6030 ( \6373 , \6060 );
or \U$6031 ( \6374 , \6372 , \6373 );
nand \U$6032 ( \6375 , \4787 , \4791 );
nand \U$6033 ( \6376 , \6374 , \6375 );
not \U$6034 ( \6377 , \6376 );
not \U$6035 ( \6378 , \6377 );
or \U$6036 ( \6379 , \6371 , \6378 );
or \U$6037 ( \6380 , \6370 , \6377 );
nand \U$6038 ( \6381 , \6379 , \6380 );
and \U$6039 ( \6382 , \4742 , \1147 );
and \U$6040 ( \6383 , \6023 , \1090 );
nor \U$6041 ( \6384 , \6382 , \6383 );
and \U$6042 ( \6385 , \6381 , \6384 );
not \U$6043 ( \6386 , \6381 );
not \U$6044 ( \6387 , \6384 );
and \U$6045 ( \6388 , \6386 , \6387 );
nor \U$6046 ( \6389 , \6385 , \6388 );
not \U$6047 ( \6390 , \6389 );
not \U$6048 ( \6391 , \6390 );
or \U$6049 ( \6392 , \6365 , \6391 );
not \U$6050 ( \6393 , \6363 );
not \U$6051 ( \6394 , \6389 );
or \U$6052 ( \6395 , \6393 , \6394 );
xor \U$6053 ( \6396 , \6328 , \6323 );
xor \U$6054 ( \6397 , \6396 , \6334 );
nand \U$6055 ( \6398 , \6395 , \6397 );
nand \U$6056 ( \6399 , \6392 , \6398 );
not \U$6057 ( \6400 , \6399 );
or \U$6058 ( \6401 , \6344 , \6400 );
or \U$6059 ( \6402 , \6343 , \6399 );
xor \U$6060 ( \6403 , \6278 , \6283 );
and \U$6061 ( \6404 , \6403 , \6289 );
and \U$6062 ( \6405 , \6278 , \6283 );
or \U$6063 ( \6406 , \6404 , \6405 );
not \U$6064 ( \6407 , \6362 );
nand \U$6065 ( \6408 , \6407 , \6355 );
not \U$6066 ( \6409 , \6408 );
not \U$6067 ( \6410 , \6349 );
or \U$6068 ( \6411 , \6409 , \6410 );
nand \U$6069 ( \6412 , \6354 , \6362 );
nand \U$6070 ( \6413 , \6411 , \6412 );
xor \U$6071 ( \6414 , \6406 , \6413 );
not \U$6072 ( \6415 , \6377 );
not \U$6073 ( \6416 , \6384 );
or \U$6074 ( \6417 , \6415 , \6416 );
nand \U$6075 ( \6418 , \6417 , \6370 );
nand \U$6076 ( \6419 , \6387 , \6376 );
nand \U$6077 ( \6420 , \6418 , \6419 );
xor \U$6078 ( \6421 , \6414 , \6420 );
nand \U$6079 ( \6422 , \6402 , \6421 );
nand \U$6080 ( \6423 , \6401 , \6422 );
or \U$6081 ( \6424 , \6295 , \6423 );
xor \U$6082 ( \6425 , \5847 , \5857 );
and \U$6083 ( \6426 , \6425 , \5865 );
and \U$6084 ( \6427 , \5847 , \5857 );
or \U$6085 ( \6428 , \6426 , \6427 );
xor \U$6086 ( \6429 , \6318 , \6337 );
and \U$6087 ( \6430 , \6429 , \6342 );
and \U$6088 ( \6431 , \6318 , \6337 );
or \U$6089 ( \6432 , \6430 , \6431 );
xor \U$6090 ( \6433 , \6428 , \6432 );
xor \U$6091 ( \6434 , \6406 , \6413 );
and \U$6092 ( \6435 , \6434 , \6420 );
and \U$6093 ( \6436 , \6406 , \6413 );
or \U$6094 ( \6437 , \6435 , \6436 );
xor \U$6095 ( \6438 , \6433 , \6437 );
nand \U$6096 ( \6439 , \6424 , \6438 );
nand \U$6097 ( \6440 , \6295 , \6423 );
nand \U$6098 ( \6441 , \6439 , \6440 );
xor \U$6099 ( \6442 , \6428 , \6432 );
and \U$6100 ( \6443 , \6442 , \6437 );
and \U$6101 ( \6444 , \6428 , \6432 );
or \U$6102 ( \6445 , \6443 , \6444 );
xor \U$6103 ( \6446 , \4553 , \4673 );
xor \U$6104 ( \6447 , \6446 , \4821 );
xor \U$6105 ( \6448 , \6445 , \6447 );
xor \U$6106 ( \6449 , \4734 , \4778 );
xor \U$6107 ( \6450 , \6449 , \4818 );
xor \U$6108 ( \6451 , \4590 , \4670 );
xor \U$6109 ( \6452 , \6451 , \4629 );
xor \U$6110 ( \6453 , \6450 , \6452 );
xor \U$6111 ( \6454 , \4759 , \4776 );
xor \U$6112 ( \6455 , \6454 , \4744 );
xor \U$6113 ( \6456 , \4793 , \4804 );
xor \U$6114 ( \6457 , \6456 , \4815 );
xor \U$6115 ( \6458 , \6455 , \6457 );
xor \U$6116 ( \6459 , \4655 , \4668 );
xor \U$6117 ( \6460 , \6459 , \4644 );
and \U$6118 ( \6461 , \6458 , \6460 );
and \U$6119 ( \6462 , \6455 , \6457 );
or \U$6120 ( \6463 , \6461 , \6462 );
and \U$6121 ( \6464 , \6453 , \6463 );
and \U$6122 ( \6465 , \6450 , \6452 );
or \U$6123 ( \6466 , \6464 , \6465 );
xor \U$6124 ( \6467 , \6448 , \6466 );
xor \U$6125 ( \6468 , \6441 , \6467 );
xor \U$6126 ( \6469 , \6455 , \6457 );
xor \U$6127 ( \6470 , \6469 , \6460 );
not \U$6128 ( \6471 , \1011 );
not \U$6129 ( \6472 , RIbb2f160_11);
not \U$6130 ( \6473 , \4639 );
or \U$6131 ( \6474 , \6472 , \6473 );
nand \U$6132 ( \6475 , \3202 , \1805 );
nand \U$6133 ( \6476 , \6474 , \6475 );
not \U$6134 ( \6477 , \6476 );
or \U$6135 ( \6478 , \6471 , \6477 );
nand \U$6136 ( \6479 , \1077 , \6305 );
nand \U$6137 ( \6480 , \6478 , \6479 );
not \U$6138 ( \6481 , \1533 );
not \U$6139 ( \6482 , RIbb2f250_9);
not \U$6140 ( \6483 , \3655 );
or \U$6141 ( \6484 , \6482 , \6483 );
nand \U$6142 ( \6485 , \3654 , \1566 );
nand \U$6143 ( \6486 , \6484 , \6485 );
not \U$6144 ( \6487 , \6486 );
or \U$6145 ( \6488 , \6481 , \6487 );
nand \U$6146 ( \6489 , \6176 , \1570 );
nand \U$6147 ( \6490 , \6488 , \6489 );
or \U$6148 ( \6491 , \6480 , \6490 );
not \U$6149 ( \6492 , \6251 );
not \U$6150 ( \6493 , RIbb2e530_37);
not \U$6151 ( \6494 , \814 );
or \U$6152 ( \6495 , \6493 , \6494 );
nand \U$6153 ( \6496 , \2251 , \6246 );
nand \U$6154 ( \6497 , \6495 , \6496 );
not \U$6155 ( \6498 , \6497 );
or \U$6156 ( \6499 , \6492 , \6498 );
nand \U$6157 ( \6500 , \6242 , RIbb2e530_37);
nand \U$6158 ( \6501 , \6499 , \6500 );
nand \U$6159 ( \6502 , \6491 , \6501 );
nand \U$6160 ( \6503 , \6480 , \6490 );
nand \U$6161 ( \6504 , \6502 , \6503 );
not \U$6162 ( \6505 , \6504 );
xor \U$6163 ( \6506 , \6314 , \6309 );
xor \U$6164 ( \6507 , \6506 , \6298 );
nand \U$6165 ( \6508 , \6505 , \6507 );
not \U$6166 ( \6509 , \6508 );
xor \U$6167 ( \6510 , \6194 , \6276 );
xor \U$6168 ( \6511 , \6510 , \6290 );
not \U$6169 ( \6512 , \6511 );
or \U$6170 ( \6513 , \6509 , \6512 );
not \U$6171 ( \6514 , \6507 );
nand \U$6172 ( \6515 , \6504 , \6514 );
nand \U$6173 ( \6516 , \6513 , \6515 );
nor \U$6174 ( \6517 , \6470 , \6516 );
and \U$6175 ( \6518 , \5831 , \5833 );
not \U$6176 ( \6519 , \5831 );
and \U$6177 ( \6520 , \6519 , \5834 );
or \U$6178 ( \6521 , \6518 , \6520 );
xnor \U$6179 ( \6522 , \6521 , \5866 );
or \U$6180 ( \6523 , \6517 , \6522 );
nand \U$6181 ( \6524 , \6470 , \6516 );
nand \U$6182 ( \6525 , \6523 , \6524 );
xor \U$6183 ( \6526 , \6450 , \6452 );
xor \U$6184 ( \6527 , \6526 , \6463 );
xor \U$6185 ( \6528 , \6525 , \6527 );
xor \U$6186 ( \6529 , \5869 , \5871 );
xor \U$6187 ( \6530 , \6529 , \5881 );
and \U$6188 ( \6531 , \6528 , \6530 );
and \U$6189 ( \6532 , \6525 , \6527 );
or \U$6190 ( \6533 , \6531 , \6532 );
and \U$6191 ( \6534 , \6468 , \6533 );
and \U$6192 ( \6535 , \6441 , \6467 );
or \U$6193 ( \6536 , \6534 , \6535 );
xor \U$6194 ( \6537 , \5887 , \6536 );
xor \U$6195 ( \6538 , \6445 , \6447 );
and \U$6196 ( \6539 , \6538 , \6466 );
and \U$6197 ( \6540 , \6445 , \6447 );
or \U$6198 ( \6541 , \6539 , \6540 );
xor \U$6199 ( \6542 , \4824 , \4826 );
xor \U$6200 ( \6543 , \6542 , \4857 );
xor \U$6201 ( \6544 , \6541 , \6543 );
xor \U$6202 ( \6545 , \4536 , \4538 );
xor \U$6203 ( \6546 , \6545 , \4541 );
xor \U$6204 ( \6547 , \6544 , \6546 );
and \U$6205 ( \6548 , \6537 , \6547 );
and \U$6206 ( \6549 , \5887 , \6536 );
or \U$6207 ( \6550 , \6548 , \6549 );
not \U$6208 ( \6551 , \6550 );
and \U$6209 ( \6552 , \4121 , \4070 );
not \U$6210 ( \6553 , \4121 );
and \U$6211 ( \6554 , \6553 , \4123 );
or \U$6212 ( \6555 , \6552 , \6554 );
and \U$6213 ( \6556 , \6555 , \4058 );
not \U$6214 ( \6557 , \6555 );
and \U$6215 ( \6558 , \6557 , \4059 );
nor \U$6216 ( \6559 , \6556 , \6558 );
not \U$6217 ( \6560 , \6559 );
xor \U$6218 ( \6561 , \4860 , \4516 );
xor \U$6219 ( \6562 , \6561 , \4544 );
not \U$6220 ( \6563 , \6562 );
or \U$6221 ( \6564 , \6560 , \6563 );
or \U$6222 ( \6565 , \6559 , \6562 );
nand \U$6223 ( \6566 , \6564 , \6565 );
xor \U$6224 ( \6567 , \6541 , \6543 );
and \U$6225 ( \6568 , \6567 , \6546 );
and \U$6226 ( \6569 , \6541 , \6543 );
or \U$6227 ( \6570 , \6568 , \6569 );
xnor \U$6228 ( \6571 , \6566 , \6570 );
nand \U$6229 ( \6572 , \6551 , \6571 );
not \U$6230 ( \6573 , \6572 );
xor \U$6231 ( \6574 , \5887 , \6536 );
xor \U$6232 ( \6575 , \6574 , \6547 );
not \U$6233 ( \6576 , \6575 );
xor \U$6234 ( \6577 , \5826 , \5828 );
xor \U$6235 ( \6578 , \6577 , \5884 );
xor \U$6236 ( \6579 , \6293 , \6190 );
xnor \U$6237 ( \6580 , \6579 , \6048 );
not \U$6238 ( \6581 , \6580 );
not \U$6239 ( \6582 , \6581 );
not \U$6240 ( \6583 , \520 );
nand \U$6241 ( \6584 , \519 , \6583 );
nor \U$6242 ( \6585 , \4355 , \6584 );
not \U$6243 ( \6586 , \6585 );
not \U$6244 ( \6587 , \5941 );
or \U$6245 ( \6588 , \6586 , \6587 );
not \U$6246 ( \6589 , \6584 );
and \U$6247 ( \6590 , \4370 , \6589 );
not \U$6248 ( \6591 , \6583 );
not \U$6249 ( \6592 , \620 );
or \U$6250 ( \6593 , \6591 , \6592 );
nand \U$6251 ( \6594 , \6593 , \624 );
nor \U$6252 ( \6595 , \6590 , \6594 );
nand \U$6253 ( \6596 , \6588 , \6595 );
nor \U$6254 ( \6597 , \627 , \521 );
and \U$6255 ( \6598 , \6596 , \6597 );
not \U$6256 ( \6599 , \6596 );
not \U$6257 ( \6600 , \6597 );
and \U$6258 ( \6601 , \6599 , \6600 );
nor \U$6259 ( \6602 , \6598 , \6601 );
buf \U$6260 ( \6603 , \6602 );
buf \U$6261 ( \6604 , \6603 );
and \U$6262 ( \6605 , \6604 , \1393 );
not \U$6263 ( \6606 , \1376 );
not \U$6264 ( \6607 , \6233 );
or \U$6265 ( \6608 , \6606 , \6607 );
xor \U$6266 ( \6609 , \1313 , \5957 );
nand \U$6267 ( \6610 , \6609 , \1429 );
nand \U$6268 ( \6611 , \6608 , \6610 );
xor \U$6269 ( \6612 , \6605 , \6611 );
not \U$6270 ( \6613 , \1294 );
not \U$6271 ( \6614 , \6271 );
or \U$6272 ( \6615 , \6613 , \6614 );
not \U$6273 ( \6616 , \1246 );
not \U$6274 ( \6617 , \4698 );
or \U$6275 ( \6618 , \6616 , \6617 );
nand \U$6276 ( \6619 , \4699 , \1245 );
nand \U$6277 ( \6620 , \6618 , \6619 );
nand \U$6278 ( \6621 , \6620 , \1265 );
nand \U$6279 ( \6622 , \6615 , \6621 );
and \U$6280 ( \6623 , \6612 , \6622 );
and \U$6281 ( \6624 , \6605 , \6611 );
or \U$6282 ( \6625 , \6623 , \6624 );
not \U$6283 ( \6626 , \6625 );
xor \U$6284 ( \6627 , \6255 , \6235 );
xnor \U$6285 ( \6628 , \6627 , \6273 );
nand \U$6286 ( \6629 , \6626 , \6628 );
not \U$6287 ( \6630 , \6629 );
not \U$6288 ( \6631 , \1077 );
not \U$6289 ( \6632 , \6476 );
or \U$6290 ( \6633 , \6631 , \6632 );
not \U$6291 ( \6634 , RIbb2f160_11);
not \U$6292 ( \6635 , \3905 );
or \U$6293 ( \6636 , \6634 , \6635 );
nand \U$6294 ( \6637 , \3632 , \1805 );
nand \U$6295 ( \6638 , \6636 , \6637 );
nand \U$6296 ( \6639 , \6638 , \1011 );
nand \U$6297 ( \6640 , \6633 , \6639 );
not \U$6298 ( \6641 , \916 );
not \U$6299 ( \6642 , RIbb2f070_13);
not \U$6300 ( \6643 , \6301 );
or \U$6301 ( \6644 , \6642 , \6643 );
nand \U$6302 ( \6645 , \3620 , \1656 );
nand \U$6303 ( \6646 , \6644 , \6645 );
not \U$6304 ( \6647 , \6646 );
or \U$6305 ( \6648 , \6641 , \6647 );
not \U$6306 ( \6649 , \6113 );
nand \U$6307 ( \6650 , \6649 , \998 );
nand \U$6308 ( \6651 , \6648 , \6650 );
or \U$6309 ( \6652 , \6640 , \6651 );
not \U$6310 ( \6653 , \2980 );
and \U$6311 ( \6654 , RIbb2ead0_25, \1140 );
not \U$6312 ( \6655 , RIbb2ead0_25);
and \U$6313 ( \6656 , \6655 , \1139 );
or \U$6314 ( \6657 , \6654 , \6656 );
not \U$6315 ( \6658 , \6657 );
or \U$6316 ( \6659 , \6653 , \6658 );
not \U$6317 ( \6660 , \6129 );
nand \U$6318 ( \6661 , \6660 , \2963 );
nand \U$6319 ( \6662 , \6659 , \6661 );
nand \U$6320 ( \6663 , \6652 , \6662 );
nand \U$6321 ( \6664 , \6640 , \6651 );
nand \U$6322 ( \6665 , \6663 , \6664 );
not \U$6323 ( \6666 , \6665 );
or \U$6324 ( \6667 , \6630 , \6666 );
not \U$6325 ( \6668 , \6628 );
nand \U$6326 ( \6669 , \6668 , \6625 );
nand \U$6327 ( \6670 , \6667 , \6669 );
not \U$6328 ( \6671 , \2941 );
not \U$6329 ( \6672 , \5909 );
or \U$6330 ( \6673 , \6671 , \6672 );
not \U$6331 ( \6674 , RIbb2e800_31);
not \U$6332 ( \6675 , \1887 );
or \U$6333 ( \6676 , \6674 , \6675 );
nand \U$6334 ( \6677 , \1071 , \2917 );
nand \U$6335 ( \6678 , \6676 , \6677 );
nand \U$6336 ( \6679 , \6678 , \2940 );
nand \U$6337 ( \6680 , \6673 , \6679 );
not \U$6338 ( \6681 , \6680 );
not \U$6339 ( \6682 , \5845 );
not \U$6340 ( \6683 , \6004 );
or \U$6341 ( \6684 , \6682 , \6683 );
not \U$6342 ( \6685 , RIbb2e620_35);
not \U$6343 ( \6686 , \3262 );
or \U$6344 ( \6687 , \6685 , \6686 );
not \U$6345 ( \6688 , RIbb2e620_35);
nand \U$6346 ( \6689 , \3261 , \6688 );
nand \U$6347 ( \6690 , \6687 , \6689 );
nand \U$6348 ( \6691 , \6690 , \4712 );
nand \U$6349 ( \6692 , \6684 , \6691 );
not \U$6350 ( \6693 , \6692 );
or \U$6351 ( \6694 , \6681 , \6693 );
not \U$6352 ( \6695 , \6692 );
not \U$6353 ( \6696 , \6695 );
not \U$6354 ( \6697 , \6680 );
not \U$6355 ( \6698 , \6697 );
or \U$6356 ( \6699 , \6696 , \6698 );
not \U$6357 ( \6700 , \2078 );
not \U$6358 ( \6701 , \6032 );
or \U$6359 ( \6702 , \6700 , \6701 );
not \U$6360 ( \6703 , RIbb2ecb0_21);
not \U$6361 ( \6704 , \3116 );
or \U$6362 ( \6705 , \6703 , \6704 );
nand \U$6363 ( \6706 , \3117 , \849 );
nand \U$6364 ( \6707 , \6705 , \6706 );
nand \U$6365 ( \6708 , \6707 , \2077 );
nand \U$6366 ( \6709 , \6702 , \6708 );
nand \U$6367 ( \6710 , \6699 , \6709 );
nand \U$6368 ( \6711 , \6694 , \6710 );
not \U$6369 ( \6712 , \6711 );
not \U$6370 ( \6713 , \1147 );
not \U$6371 ( \6714 , \6015 );
or \U$6372 ( \6715 , \6713 , \6714 );
not \U$6373 ( \6716 , RIbb2f430_5);
not \U$6374 ( \6717 , \4088 );
or \U$6375 ( \6718 , \6716 , \6717 );
nand \U$6376 ( \6719 , \4089 , \1980 );
nand \U$6377 ( \6720 , \6718 , \6719 );
nand \U$6378 ( \6721 , \6720 , \1090 );
nand \U$6379 ( \6722 , \6715 , \6721 );
not \U$6380 ( \6723 , \6722 );
not \U$6381 ( \6724 , \1702 );
not \U$6382 ( \6725 , RIbb2f340_7);
not \U$6383 ( \6726 , \4411 );
or \U$6384 ( \6727 , \6725 , \6726 );
nand \U$6385 ( \6728 , \3003 , \2700 );
nand \U$6386 ( \6729 , \6727 , \6728 );
not \U$6387 ( \6730 , \6729 );
or \U$6388 ( \6731 , \6724 , \6730 );
nand \U$6389 ( \6732 , \5973 , \1737 );
nand \U$6390 ( \6733 , \6731 , \6732 );
not \U$6391 ( \6734 , \6733 );
nand \U$6392 ( \6735 , \6723 , \6734 );
not \U$6393 ( \6736 , \3407 );
not \U$6394 ( \6737 , RIbb2ebc0_23);
not \U$6395 ( \6738 , \1284 );
or \U$6396 ( \6739 , \6737 , \6738 );
not \U$6397 ( \6740 , \5407 );
nand \U$6398 ( \6741 , \6740 , \2073 );
nand \U$6399 ( \6742 , \6739 , \6741 );
not \U$6400 ( \6743 , \6742 );
or \U$6401 ( \6744 , \6736 , \6743 );
nand \U$6402 ( \6745 , \5984 , \3383 );
nand \U$6403 ( \6746 , \6744 , \6745 );
and \U$6404 ( \6747 , \6735 , \6746 );
nor \U$6405 ( \6748 , \6723 , \6734 );
nor \U$6406 ( \6749 , \6747 , \6748 );
nand \U$6407 ( \6750 , \6712 , \6749 );
not \U$6408 ( \6751 , \6750 );
not \U$6409 ( \6752 , \2922 );
not \U$6410 ( \6753 , RIbb2e8f0_29);
not \U$6411 ( \6754 , \1550 );
or \U$6412 ( \6755 , \6753 , \6754 );
nand \U$6413 ( \6756 , \5004 , \2911 );
nand \U$6414 ( \6757 , \6755 , \6756 );
not \U$6415 ( \6758 , \6757 );
or \U$6416 ( \6759 , \6752 , \6758 );
nand \U$6417 ( \6760 , \5893 , \2925 );
nand \U$6418 ( \6761 , \6759 , \6760 );
not \U$6419 ( \6762 , \6761 );
not \U$6420 ( \6763 , \832 );
not \U$6421 ( \6764 , RIbb2ee90_17);
not \U$6422 ( \6765 , \2116 );
or \U$6423 ( \6766 , \6764 , \6765 );
nand \U$6424 ( \6767 , \4450 , \3699 );
nand \U$6425 ( \6768 , \6766 , \6767 );
not \U$6426 ( \6769 , \6768 );
or \U$6427 ( \6770 , \6763 , \6769 );
nand \U$6428 ( \6771 , \6092 , \836 );
nand \U$6429 ( \6772 , \6770 , \6771 );
not \U$6430 ( \6773 , \6772 );
or \U$6431 ( \6774 , \6762 , \6773 );
or \U$6432 ( \6775 , \6772 , \6761 );
not \U$6433 ( \6776 , \855 );
not \U$6434 ( \6777 , \5927 );
or \U$6435 ( \6778 , \6776 , \6777 );
not \U$6436 ( \6779 , RIbb2eda0_19);
not \U$6437 ( \6780 , \6097 );
or \U$6438 ( \6781 , \6779 , \6780 );
nand \U$6439 ( \6782 , \1339 , \1776 );
nand \U$6440 ( \6783 , \6781 , \6782 );
nand \U$6441 ( \6784 , \6783 , \853 );
nand \U$6442 ( \6785 , \6778 , \6784 );
nand \U$6443 ( \6786 , \6775 , \6785 );
nand \U$6444 ( \6787 , \6774 , \6786 );
not \U$6445 ( \6788 , \6787 );
or \U$6446 ( \6789 , \6751 , \6788 );
not \U$6447 ( \6790 , \6749 );
nand \U$6448 ( \6791 , \6711 , \6790 );
nand \U$6449 ( \6792 , \6789 , \6791 );
xor \U$6450 ( \6793 , \6670 , \6792 );
not \U$6451 ( \6794 , \6105 );
not \U$6452 ( \6795 , \6157 );
or \U$6453 ( \6796 , \6794 , \6795 );
or \U$6454 ( \6797 , \6105 , \6157 );
nand \U$6455 ( \6798 , \6796 , \6797 );
xor \U$6456 ( \6799 , \6186 , \6798 );
and \U$6457 ( \6800 , \6793 , \6799 );
and \U$6458 ( \6801 , \6670 , \6792 );
or \U$6459 ( \6802 , \6800 , \6801 );
not \U$6460 ( \6803 , \6802 );
or \U$6461 ( \6804 , \6582 , \6803 );
not \U$6462 ( \6805 , \6580 );
not \U$6463 ( \6806 , \6802 );
not \U$6464 ( \6807 , \6806 );
or \U$6465 ( \6808 , \6805 , \6807 );
and \U$6466 ( \6809 , \5938 , \6044 );
not \U$6467 ( \6810 , \5938 );
and \U$6468 ( \6811 , \6810 , \6045 );
nor \U$6469 ( \6812 , \6809 , \6811 );
xor \U$6470 ( \6813 , \6812 , \5996 );
not \U$6471 ( \6814 , \6813 );
not \U$6472 ( \6815 , \6501 );
xor \U$6473 ( \6816 , \6815 , \6480 );
xor \U$6474 ( \6817 , \6816 , \6490 );
not \U$6475 ( \6818 , \6817 );
not \U$6476 ( \6819 , \6818 );
xnor \U$6477 ( \6820 , \6103 , \6080 );
and \U$6478 ( \6821 , \6820 , \6063 );
not \U$6479 ( \6822 , \6820 );
and \U$6480 ( \6823 , \6822 , \6062 );
or \U$6481 ( \6824 , \6821 , \6823 );
not \U$6482 ( \6825 , \6824 );
not \U$6483 ( \6826 , \6825 );
or \U$6484 ( \6827 , \6819 , \6826 );
not \U$6485 ( \6828 , \6817 );
not \U$6486 ( \6829 , \6824 );
or \U$6487 ( \6830 , \6828 , \6829 );
xor \U$6488 ( \6831 , \5975 , \5994 );
xor \U$6489 ( \6832 , \6831 , \5958 );
nand \U$6490 ( \6833 , \6830 , \6832 );
nand \U$6491 ( \6834 , \6827 , \6833 );
not \U$6492 ( \6835 , \6834 );
or \U$6493 ( \6836 , \6814 , \6835 );
or \U$6494 ( \6837 , \6834 , \6813 );
not \U$6495 ( \6838 , \4791 );
not \U$6496 ( \6839 , \6053 );
or \U$6497 ( \6840 , \6838 , \6839 );
not \U$6498 ( \6841 , RIbb2e710_33);
not \U$6499 ( \6842 , \993 );
or \U$6500 ( \6843 , \6841 , \6842 );
not \U$6501 ( \6844 , RIbb2e710_33);
nand \U$6502 ( \6845 , \987 , \6844 );
nand \U$6503 ( \6846 , \6843 , \6845 );
nand \U$6504 ( \6847 , \6846 , \3887 );
nand \U$6505 ( \6848 , \6840 , \6847 );
not \U$6506 ( \6849 , \3445 );
not \U$6507 ( \6850 , RIbb2e9e0_27);
not \U$6508 ( \6851 , \1689 );
or \U$6509 ( \6852 , \6850 , \6851 );
nand \U$6510 ( \6853 , \1691 , \3462 );
nand \U$6511 ( \6854 , \6852 , \6853 );
not \U$6512 ( \6855 , \6854 );
or \U$6513 ( \6856 , \6849 , \6855 );
not \U$6514 ( \6857 , \6069 );
nand \U$6515 ( \6858 , \6857 , \3465 );
nand \U$6516 ( \6859 , \6856 , \6858 );
xor \U$6517 ( \6860 , \6848 , \6859 );
not \U$6518 ( \6861 , \1445 );
and \U$6519 ( \6862 , RIbb2ef80_15, \3344 );
not \U$6520 ( \6863 , RIbb2ef80_15);
and \U$6521 ( \6864 , \6863 , \3343 );
or \U$6522 ( \6865 , \6862 , \6864 );
not \U$6523 ( \6866 , \6865 );
or \U$6524 ( \6867 , \6861 , \6866 );
nand \U$6525 ( \6868 , \6149 , \1517 );
nand \U$6526 ( \6869 , \6867 , \6868 );
and \U$6527 ( \6870 , \6860 , \6869 );
and \U$6528 ( \6871 , \6848 , \6859 );
or \U$6529 ( \6872 , \6870 , \6871 );
xor \U$6530 ( \6873 , \5918 , \5902 );
xor \U$6531 ( \6874 , \6873 , \5936 );
xor \U$6532 ( \6875 , \6872 , \6874 );
xor \U$6533 ( \6876 , \6041 , \6008 );
xor \U$6534 ( \6877 , \6876 , \6025 );
and \U$6535 ( \6878 , \6875 , \6877 );
and \U$6536 ( \6879 , \6872 , \6874 );
or \U$6537 ( \6880 , \6878 , \6879 );
nand \U$6538 ( \6881 , \6837 , \6880 );
nand \U$6539 ( \6882 , \6836 , \6881 );
nand \U$6540 ( \6883 , \6808 , \6882 );
nand \U$6541 ( \6884 , \6804 , \6883 );
xor \U$6542 ( \6885 , \6295 , \6423 );
xor \U$6543 ( \6886 , \6885 , \6438 );
or \U$6544 ( \6887 , \6884 , \6886 );
xor \U$6545 ( \6888 , \6525 , \6527 );
xor \U$6546 ( \6889 , \6888 , \6530 );
nand \U$6547 ( \6890 , \6887 , \6889 );
nand \U$6548 ( \6891 , \6886 , \6884 );
nand \U$6549 ( \6892 , \6890 , \6891 );
xor \U$6550 ( \6893 , \6578 , \6892 );
xor \U$6551 ( \6894 , \6441 , \6467 );
xor \U$6552 ( \6895 , \6894 , \6533 );
and \U$6553 ( \6896 , \6893 , \6895 );
and \U$6554 ( \6897 , \6578 , \6892 );
or \U$6555 ( \6898 , \6896 , \6897 );
not \U$6556 ( \6899 , \6898 );
nand \U$6557 ( \6900 , \6576 , \6899 );
buf \U$6558 ( \6901 , \6900 );
xor \U$6559 ( \6902 , \6578 , \6892 );
xor \U$6560 ( \6903 , \6902 , \6895 );
xor \U$6561 ( \6904 , \6625 , \6668 );
xnor \U$6562 ( \6905 , \6904 , \6665 );
not \U$6563 ( \6906 , \6905 );
not \U$6564 ( \6907 , \6906 );
xor \U$6565 ( \6908 , \6787 , \6790 );
xnor \U$6566 ( \6909 , \6908 , \6711 );
not \U$6567 ( \6910 , \6909 );
not \U$6568 ( \6911 , \6910 );
or \U$6569 ( \6912 , \6907 , \6911 );
xor \U$6570 ( \6913 , \6872 , \6874 );
xor \U$6571 ( \6914 , \6913 , \6877 );
nand \U$6572 ( \6915 , \6909 , \6905 );
nand \U$6573 ( \6916 , \6914 , \6915 );
nand \U$6574 ( \6917 , \6912 , \6916 );
xor \U$6575 ( \6918 , \6670 , \6792 );
xor \U$6576 ( \6919 , \6918 , \6799 );
xor \U$6577 ( \6920 , \6917 , \6919 );
xor \U$6578 ( \6921 , \6605 , \6611 );
xor \U$6579 ( \6922 , \6921 , \6622 );
not \U$6580 ( \6923 , \519 );
nor \U$6581 ( \6924 , \6923 , \4355 );
not \U$6582 ( \6925 , \6924 );
not \U$6583 ( \6926 , \5941 );
or \U$6584 ( \6927 , \6925 , \6926 );
and \U$6585 ( \6928 , \4370 , \519 );
nor \U$6586 ( \6929 , \6928 , \620 );
nand \U$6587 ( \6930 , \6927 , \6929 );
nand \U$6588 ( \6931 , \6583 , \624 );
not \U$6589 ( \6932 , \6931 );
and \U$6590 ( \6933 , \6930 , \6932 );
not \U$6591 ( \6934 , \6930 );
and \U$6592 ( \6935 , \6934 , \6931 );
nor \U$6593 ( \6936 , \6933 , \6935 );
buf \U$6594 ( \6937 , \6936 );
not \U$6595 ( \6938 , \6937 );
not \U$6596 ( \6939 , \6938 );
and \U$6597 ( \6940 , \1313 , \6939 );
not \U$6598 ( \6941 , \1430 );
not \U$6599 ( \6942 , \1313 );
not \U$6600 ( \6943 , \6604 );
not \U$6601 ( \6944 , \6943 );
or \U$6602 ( \6945 , \6942 , \6944 );
nand \U$6603 ( \6946 , \6604 , \1951 );
nand \U$6604 ( \6947 , \6945 , \6946 );
not \U$6605 ( \6948 , \6947 );
or \U$6606 ( \6949 , \6941 , \6948 );
nand \U$6607 ( \6950 , \6609 , \1376 );
nand \U$6608 ( \6951 , \6949 , \6950 );
xor \U$6609 ( \6952 , \6940 , \6951 );
not \U$6610 ( \6953 , \2963 );
not \U$6611 ( \6954 , \6657 );
or \U$6612 ( \6955 , \6953 , \6954 );
and \U$6613 ( \6956 , RIbb2ead0_25, \3066 );
not \U$6614 ( \6957 , RIbb2ead0_25);
and \U$6615 ( \6958 , \6957 , \1114 );
or \U$6616 ( \6959 , \6956 , \6958 );
nand \U$6617 ( \6960 , \6959 , \2980 );
nand \U$6618 ( \6961 , \6955 , \6960 );
and \U$6619 ( \6962 , \6952 , \6961 );
and \U$6620 ( \6963 , \6940 , \6951 );
or \U$6621 ( \6964 , \6962 , \6963 );
xor \U$6622 ( \6965 , \6922 , \6964 );
not \U$6623 ( \6966 , \2922 );
not \U$6624 ( \6967 , RIbb2e8f0_29);
not \U$6625 ( \6968 , \4580 );
or \U$6626 ( \6969 , \6967 , \6968 );
not \U$6627 ( \6970 , RIbb2e8f0_29);
nand \U$6628 ( \6971 , \3484 , \6970 );
nand \U$6629 ( \6972 , \6969 , \6971 );
not \U$6630 ( \6973 , \6972 );
or \U$6631 ( \6974 , \6966 , \6973 );
nand \U$6632 ( \6975 , \6757 , \2925 );
nand \U$6633 ( \6976 , \6974 , \6975 );
not \U$6634 ( \6977 , \3105 );
not \U$6635 ( \6978 , \6865 );
or \U$6636 ( \6979 , \6977 , \6978 );
and \U$6637 ( \6980 , RIbb2ef80_15, \4216 );
not \U$6638 ( \6981 , RIbb2ef80_15);
and \U$6639 ( \6982 , \6981 , \3167 );
or \U$6640 ( \6983 , \6980 , \6982 );
nand \U$6641 ( \6984 , \6983 , \1445 );
nand \U$6642 ( \6985 , \6979 , \6984 );
xor \U$6643 ( \6986 , \6976 , \6985 );
not \U$6644 ( \6987 , \836 );
not \U$6645 ( \6988 , \6768 );
or \U$6646 ( \6989 , \6987 , \6988 );
not \U$6647 ( \6990 , RIbb2ee90_17);
not \U$6648 ( \6991 , \3319 );
or \U$6649 ( \6992 , \6990 , \6991 );
nand \U$6650 ( \6993 , \2225 , \3057 );
nand \U$6651 ( \6994 , \6992 , \6993 );
nand \U$6652 ( \6995 , \6994 , \832 );
nand \U$6653 ( \6996 , \6989 , \6995 );
and \U$6654 ( \6997 , \6986 , \6996 );
and \U$6655 ( \6998 , \6976 , \6985 );
or \U$6656 ( \6999 , \6997 , \6998 );
and \U$6657 ( \7000 , \6965 , \6999 );
and \U$6658 ( \7001 , \6922 , \6964 );
or \U$6659 ( \7002 , \7000 , \7001 );
not \U$6660 ( \7003 , \998 );
not \U$6661 ( \7004 , \6646 );
or \U$6662 ( \7005 , \7003 , \7004 );
not \U$6663 ( \7006 , RIbb2f070_13);
not \U$6664 ( \7007 , \4639 );
or \U$6665 ( \7008 , \7006 , \7007 );
not \U$6666 ( \7009 , \4639 );
nand \U$6667 ( \7010 , \7009 , \1656 );
nand \U$6668 ( \7011 , \7008 , \7010 );
nand \U$6669 ( \7012 , \7011 , \916 );
nand \U$6670 ( \7013 , \7005 , \7012 );
not \U$6671 ( \7014 , \1077 );
not \U$6672 ( \7015 , \6638 );
or \U$6673 ( \7016 , \7014 , \7015 );
not \U$6674 ( \7017 , RIbb2f160_11);
not \U$6675 ( \7018 , \3653 );
not \U$6676 ( \7019 , \7018 );
or \U$6677 ( \7020 , \7017 , \7019 );
not \U$6678 ( \7021 , \7018 );
nand \U$6679 ( \7022 , \7021 , \1805 );
nand \U$6680 ( \7023 , \7020 , \7022 );
nand \U$6681 ( \7024 , \7023 , \1011 );
nand \U$6682 ( \7025 , \7016 , \7024 );
or \U$6683 ( \7026 , \7013 , \7025 );
not \U$6684 ( \7027 , \3465 );
not \U$6685 ( \7028 , \6854 );
or \U$6686 ( \7029 , \7027 , \7028 );
not \U$6687 ( \7030 , RIbb2e9e0_27);
not \U$6688 ( \7031 , \3773 );
or \U$6689 ( \7032 , \7030 , \7031 );
not \U$6690 ( \7033 , \3773 );
nand \U$6691 ( \7034 , \7033 , \3462 );
nand \U$6692 ( \7035 , \7032 , \7034 );
nand \U$6693 ( \7036 , \7035 , \3445 );
nand \U$6694 ( \7037 , \7029 , \7036 );
nand \U$6695 ( \7038 , \7026 , \7037 );
nand \U$6696 ( \7039 , \7025 , \7013 );
nand \U$6697 ( \7040 , \7038 , \7039 );
not \U$6698 ( \7041 , \6761 );
xor \U$6699 ( \7042 , \6772 , \6785 );
xnor \U$6700 ( \7043 , \7041 , \7042 );
xor \U$6701 ( \7044 , \7040 , \7043 );
xor \U$6702 ( \7045 , \6709 , \6692 );
xnor \U$6703 ( \7046 , \7045 , \6697 );
and \U$6704 ( \7047 , \7044 , \7046 );
and \U$6705 ( \7048 , \7040 , \7043 );
or \U$6706 ( \7049 , \7047 , \7048 );
xor \U$6707 ( \7050 , \7002 , \7049 );
xor \U$6708 ( \7051 , \6848 , \6859 );
xor \U$6709 ( \7052 , \7051 , \6869 );
xnor \U$6710 ( \7053 , \6746 , \6723 );
and \U$6711 ( \7054 , \7053 , \6733 );
not \U$6712 ( \7055 , \7053 );
and \U$6713 ( \7056 , \7055 , \6734 );
nor \U$6714 ( \7057 , \7054 , \7056 );
or \U$6715 ( \7058 , \7052 , \7057 );
xor \U$6716 ( \7059 , \6651 , \6640 );
xnor \U$6717 ( \7060 , \7059 , \6662 );
not \U$6718 ( \7061 , \7060 );
nand \U$6719 ( \7062 , \7058 , \7061 );
nand \U$6720 ( \7063 , \7057 , \7052 );
nand \U$6721 ( \7064 , \7062 , \7063 );
and \U$6722 ( \7065 , \7050 , \7064 );
and \U$6723 ( \7066 , \7002 , \7049 );
or \U$6724 ( \7067 , \7065 , \7066 );
and \U$6725 ( \7068 , \6920 , \7067 );
and \U$6726 ( \7069 , \6917 , \6919 );
or \U$6727 ( \7070 , \7068 , \7069 );
not \U$6728 ( \7071 , \7070 );
not \U$6729 ( \7072 , \6882 );
not \U$6730 ( \7073 , \6806 );
or \U$6731 ( \7074 , \7072 , \7073 );
or \U$6732 ( \7075 , \6882 , \6806 );
nand \U$6733 ( \7076 , \7074 , \7075 );
and \U$6734 ( \7077 , \7076 , \6581 );
not \U$6735 ( \7078 , \7076 );
and \U$6736 ( \7079 , \7078 , \6580 );
nor \U$6737 ( \7080 , \7077 , \7079 );
not \U$6738 ( \7081 , \7080 );
or \U$6739 ( \7082 , \7071 , \7081 );
or \U$6740 ( \7083 , \7080 , \7070 );
not \U$6741 ( \7084 , \1570 );
not \U$6742 ( \7085 , \6486 );
or \U$6743 ( \7086 , \7084 , \7085 );
not \U$6744 ( \7087 , RIbb2f250_9);
not \U$6745 ( \7088 , \4017 );
or \U$6746 ( \7089 , \7087 , \7088 );
nand \U$6747 ( \7090 , \4022 , \1554 );
nand \U$6748 ( \7091 , \7089 , \7090 );
nand \U$6749 ( \7092 , \7091 , \1533 );
nand \U$6750 ( \7093 , \7086 , \7092 );
xor \U$6751 ( \7094 , \6815 , \7093 );
and \U$6752 ( \7095 , RIbb2e3c8_40, RIbb2e350_41);
not \U$6753 ( \7096 , RIbb2e3c8_40);
not \U$6754 ( \7097 , RIbb2e350_41);
and \U$6755 ( \7098 , \7096 , \7097 );
nor \U$6756 ( \7099 , \7095 , \7098 );
not \U$6757 ( \7100 , \7099 );
xor \U$6758 ( \7101 , RIbb2e440_39, RIbb2e3c8_40);
and \U$6759 ( \7102 , \7100 , \7101 );
buf \U$6760 ( \7103 , \7102 );
buf \U$6761 ( \7104 , \7099 );
or \U$6762 ( \7105 , \7103 , \7104 );
nand \U$6763 ( \7106 , \7105 , RIbb2e440_39);
not \U$6764 ( \7107 , \1265 );
not \U$6765 ( \7108 , \1246 );
not \U$6766 ( \7109 , \6231 );
or \U$6767 ( \7110 , \7108 , \7109 );
buf \U$6768 ( \7111 , \6229 );
nand \U$6769 ( \7112 , \7111 , \1245 );
nand \U$6770 ( \7113 , \7110 , \7112 );
not \U$6771 ( \7114 , \7113 );
or \U$6772 ( \7115 , \7107 , \7114 );
nand \U$6773 ( \7116 , \6620 , \1294 );
nand \U$6774 ( \7117 , \7115 , \7116 );
xor \U$6775 ( \7118 , \7106 , \7117 );
not \U$6776 ( \7119 , \1147 );
not \U$6777 ( \7120 , \6720 );
or \U$6778 ( \7121 , \7119 , \7120 );
not \U$6779 ( \7122 , RIbb2f430_5);
not \U$6780 ( \7123 , \4393 );
or \U$6781 ( \7124 , \7122 , \7123 );
nand \U$6782 ( \7125 , \4394 , \1980 );
nand \U$6783 ( \7126 , \7124 , \7125 );
nand \U$6784 ( \7127 , \7126 , \1090 );
nand \U$6785 ( \7128 , \7121 , \7127 );
and \U$6786 ( \7129 , \7118 , \7128 );
and \U$6787 ( \7130 , \7106 , \7117 );
or \U$6788 ( \7131 , \7129 , \7130 );
and \U$6789 ( \7132 , \7094 , \7131 );
and \U$6790 ( \7133 , \6815 , \7093 );
or \U$6791 ( \7134 , \7132 , \7133 );
xor \U$6792 ( \7135 , \6151 , \6136 );
and \U$6793 ( \7136 , \7135 , \6124 );
not \U$6794 ( \7137 , \7135 );
and \U$6795 ( \7138 , \7137 , \6154 );
nor \U$6796 ( \7139 , \7136 , \7138 );
xor \U$6797 ( \7140 , \7134 , \7139 );
not \U$6798 ( \7141 , \4712 );
not \U$6799 ( \7142 , RIbb2e620_35);
not \U$6800 ( \7143 , \4558 );
not \U$6801 ( \7144 , \7143 );
or \U$6802 ( \7145 , \7142 , \7144 );
nand \U$6803 ( \7146 , \3453 , \3866 );
nand \U$6804 ( \7147 , \7145 , \7146 );
not \U$6805 ( \7148 , \7147 );
or \U$6806 ( \7149 , \7141 , \7148 );
nand \U$6807 ( \7150 , \6690 , \5845 );
nand \U$6808 ( \7151 , \7149 , \7150 );
not \U$6809 ( \7152 , \7151 );
not \U$6810 ( \7153 , \3613 );
not \U$6811 ( \7154 , \6678 );
or \U$6812 ( \7155 , \7153 , \7154 );
not \U$6813 ( \7156 , RIbb2e800_31);
not \U$6814 ( \7157 , \4595 );
or \U$6815 ( \7158 , \7156 , \7157 );
nand \U$6816 ( \7159 , \1038 , \2917 );
nand \U$6817 ( \7160 , \7158 , \7159 );
nand \U$6818 ( \7161 , \7160 , \2940 );
nand \U$6819 ( \7162 , \7155 , \7161 );
not \U$6820 ( \7163 , \7162 );
or \U$6821 ( \7164 , \7152 , \7163 );
or \U$6822 ( \7165 , \7151 , \7162 );
not \U$6823 ( \7166 , \853 );
not \U$6824 ( \7167 , RIbb2eda0_19);
not \U$6825 ( \7168 , \3807 );
or \U$6826 ( \7169 , \7167 , \7168 );
nand \U$6827 ( \7170 , \3810 , \1776 );
nand \U$6828 ( \7171 , \7169 , \7170 );
not \U$6829 ( \7172 , \7171 );
or \U$6830 ( \7173 , \7166 , \7172 );
nand \U$6831 ( \7174 , \6783 , \855 );
nand \U$6832 ( \7175 , \7173 , \7174 );
nand \U$6833 ( \7176 , \7165 , \7175 );
nand \U$6834 ( \7177 , \7164 , \7176 );
not \U$6835 ( \7178 , \7177 );
not \U$6836 ( \7179 , \2078 );
not \U$6837 ( \7180 , \6707 );
or \U$6838 ( \7181 , \7179 , \7180 );
not \U$6839 ( \7182 , RIbb2ecb0_21);
not \U$6840 ( \7183 , \1420 );
or \U$6841 ( \7184 , \7182 , \7183 );
nand \U$6842 ( \7185 , \1422 , \2067 );
nand \U$6843 ( \7186 , \7184 , \7185 );
nand \U$6844 ( \7187 , \7186 , \2077 );
nand \U$6845 ( \7188 , \7181 , \7187 );
not \U$6846 ( \7189 , \7188 );
not \U$6847 ( \7190 , \4791 );
not \U$6848 ( \7191 , \6846 );
or \U$6849 ( \7192 , \7190 , \7191 );
not \U$6850 ( \7193 , RIbb2e710_33);
not \U$6851 ( \7194 , \2399 );
or \U$6852 ( \7195 , \7193 , \7194 );
nand \U$6853 ( \7196 , \957 , \3864 );
nand \U$6854 ( \7197 , \7195 , \7196 );
nand \U$6855 ( \7198 , \7197 , \3887 );
nand \U$6856 ( \7199 , \7192 , \7198 );
not \U$6857 ( \7200 , \7199 );
or \U$6858 ( \7201 , \7189 , \7200 );
or \U$6859 ( \7202 , \7199 , \7188 );
not \U$6860 ( \7203 , \3383 );
not \U$6861 ( \7204 , \6742 );
or \U$6862 ( \7205 , \7203 , \7204 );
not \U$6863 ( \7206 , RIbb2ebc0_23);
not \U$6864 ( \7207 , \1170 );
or \U$6865 ( \7208 , \7206 , \7207 );
nand \U$6866 ( \7209 , \3736 , \3401 );
nand \U$6867 ( \7210 , \7208 , \7209 );
nand \U$6868 ( \7211 , \7210 , \3407 );
nand \U$6869 ( \7212 , \7205 , \7211 );
nand \U$6870 ( \7213 , \7202 , \7212 );
nand \U$6871 ( \7214 , \7201 , \7213 );
not \U$6872 ( \7215 , \7214 );
or \U$6873 ( \7216 , \7178 , \7215 );
or \U$6874 ( \7217 , \7214 , \7177 );
not \U$6875 ( \7218 , \1702 );
not \U$6876 ( \7219 , RIbb2f340_7);
not \U$6877 ( \7220 , \4040 );
or \U$6878 ( \7221 , \7219 , \7220 );
nand \U$6879 ( \7222 , \3092 , \1692 );
nand \U$6880 ( \7223 , \7221 , \7222 );
not \U$6881 ( \7224 , \7223 );
or \U$6882 ( \7225 , \7218 , \7224 );
nand \U$6883 ( \7226 , \6729 , \1737 );
nand \U$6884 ( \7227 , \7225 , \7226 );
not \U$6885 ( \7228 , \1533 );
not \U$6886 ( \7229 , RIbb2f250_9);
not \U$6887 ( \7230 , \4031 );
or \U$6888 ( \7231 , \7229 , \7230 );
nand \U$6889 ( \7232 , \4030 , \1566 );
nand \U$6890 ( \7233 , \7231 , \7232 );
not \U$6891 ( \7234 , \7233 );
or \U$6892 ( \7235 , \7228 , \7234 );
nand \U$6893 ( \7236 , \7091 , \1570 );
nand \U$6894 ( \7237 , \7235 , \7236 );
or \U$6895 ( \7238 , \7227 , \7237 );
not \U$6896 ( \7239 , \6251 );
not \U$6897 ( \7240 , RIbb2e530_37);
not \U$6898 ( \7241 , \894 );
or \U$6899 ( \7242 , \7240 , \7241 );
not \U$6900 ( \7243 , RIbb2e530_37);
nand \U$6901 ( \7244 , \893 , \7243 );
nand \U$6902 ( \7245 , \7242 , \7244 );
not \U$6903 ( \7246 , \7245 );
or \U$6904 ( \7247 , \7239 , \7246 );
nand \U$6905 ( \7248 , \6497 , \6242 );
nand \U$6906 ( \7249 , \7247 , \7248 );
nand \U$6907 ( \7250 , \7238 , \7249 );
nand \U$6908 ( \7251 , \7227 , \7237 );
nand \U$6909 ( \7252 , \7250 , \7251 );
nand \U$6910 ( \7253 , \7217 , \7252 );
nand \U$6911 ( \7254 , \7216 , \7253 );
xor \U$6912 ( \7255 , \7140 , \7254 );
not \U$6913 ( \7256 , \7255 );
not \U$6914 ( \7257 , \6817 );
not \U$6915 ( \7258 , \6825 );
or \U$6916 ( \7259 , \7257 , \7258 );
nand \U$6917 ( \7260 , \6824 , \6818 );
nand \U$6918 ( \7261 , \7259 , \7260 );
xor \U$6919 ( \7262 , \7261 , \6832 );
not \U$6920 ( \7263 , \7262 );
or \U$6921 ( \7264 , \7256 , \7263 );
or \U$6922 ( \7265 , \7255 , \7262 );
xor \U$6923 ( \7266 , \6815 , \7093 );
xor \U$6924 ( \7267 , \7266 , \7131 );
not \U$6925 ( \7268 , \7103 );
not \U$6926 ( \7269 , RIbb2e440_39);
not \U$6927 ( \7270 , \814 );
or \U$6928 ( \7271 , \7269 , \7270 );
not \U$6929 ( \7272 , RIbb2e440_39);
nand \U$6930 ( \7273 , \7272 , \2251 );
nand \U$6931 ( \7274 , \7271 , \7273 );
not \U$6932 ( \7275 , \7274 );
or \U$6933 ( \7276 , \7268 , \7275 );
nand \U$6934 ( \7277 , \7104 , RIbb2e440_39);
nand \U$6935 ( \7278 , \7276 , \7277 );
nor \U$6936 ( \7279 , \4355 , \518 );
not \U$6937 ( \7280 , \7279 );
not \U$6938 ( \7281 , \5941 );
or \U$6939 ( \7282 , \7280 , \7281 );
not \U$6940 ( \7283 , \518 );
not \U$6941 ( \7284 , \7283 );
not \U$6942 ( \7285 , \4369 );
or \U$6943 ( \7286 , \7284 , \7285 );
nand \U$6944 ( \7287 , \7286 , \613 );
not \U$6945 ( \7288 , \7287 );
nand \U$6946 ( \7289 , \7282 , \7288 );
nand \U$6947 ( \7290 , \616 , \619 );
not \U$6948 ( \7291 , \7290 );
and \U$6949 ( \7292 , \7289 , \7291 );
not \U$6950 ( \7293 , \7289 );
and \U$6951 ( \7294 , \7293 , \7290 );
nor \U$6952 ( \7295 , \7292 , \7294 );
buf \U$6953 ( \7296 , \7295 );
not \U$6954 ( \7297 , \7296 );
buf \U$6955 ( \7298 , \7297 );
not \U$6956 ( \7299 , \7298 );
buf \U$6957 ( \7300 , \7299 );
and \U$6958 ( \7301 , \1313 , \7300 );
not \U$6959 ( \7302 , \1294 );
not \U$6960 ( \7303 , \7113 );
or \U$6961 ( \7304 , \7302 , \7303 );
not \U$6962 ( \7305 , \1246 );
not \U$6963 ( \7306 , \5956 );
or \U$6964 ( \7307 , \7305 , \7306 );
buf \U$6965 ( \7308 , \5954 );
nand \U$6966 ( \7309 , \7308 , \1245 );
nand \U$6967 ( \7310 , \7307 , \7309 );
nand \U$6968 ( \7311 , \7310 , \1265 );
nand \U$6969 ( \7312 , \7304 , \7311 );
xor \U$6970 ( \7313 , \7301 , \7312 );
not \U$6971 ( \7314 , \1147 );
not \U$6972 ( \7315 , \7126 );
or \U$6973 ( \7316 , \7314 , \7315 );
not \U$6974 ( \7317 , RIbb2f430_5);
not \U$6975 ( \7318 , \4698 );
or \U$6976 ( \7319 , \7317 , \7318 );
nand \U$6977 ( \7320 , \4699 , \1898 );
nand \U$6978 ( \7321 , \7319 , \7320 );
nand \U$6979 ( \7322 , \7321 , \1090 );
nand \U$6980 ( \7323 , \7316 , \7322 );
and \U$6981 ( \7324 , \7313 , \7323 );
and \U$6982 ( \7325 , \7301 , \7312 );
or \U$6983 ( \7326 , \7324 , \7325 );
xor \U$6984 ( \7327 , \7278 , \7326 );
not \U$6985 ( \7328 , \2925 );
not \U$6986 ( \7329 , \6972 );
or \U$6987 ( \7330 , \7328 , \7329 );
not \U$6988 ( \7331 , RIbb2e8f0_29);
not \U$6989 ( \7332 , \1688 );
or \U$6990 ( \7333 , \7331 , \7332 );
nand \U$6991 ( \7334 , \3364 , \3440 );
nand \U$6992 ( \7335 , \7333 , \7334 );
nand \U$6993 ( \7336 , \7335 , \2922 );
nand \U$6994 ( \7337 , \7330 , \7336 );
not \U$6995 ( \7338 , \7337 );
not \U$6996 ( \7339 , \5845 );
not \U$6997 ( \7340 , \7147 );
or \U$6998 ( \7341 , \7339 , \7340 );
not \U$6999 ( \7342 , RIbb2e620_35);
not \U$7000 ( \7343 , \989 );
or \U$7001 ( \7344 , \7342 , \7343 );
not \U$7002 ( \7345 , \992 );
nand \U$7003 ( \7346 , \7345 , \6002 );
nand \U$7004 ( \7347 , \7344 , \7346 );
nand \U$7005 ( \7348 , \7347 , \4712 );
nand \U$7006 ( \7349 , \7341 , \7348 );
not \U$7007 ( \7350 , \7349 );
or \U$7008 ( \7351 , \7338 , \7350 );
not \U$7009 ( \7352 , \7349 );
not \U$7010 ( \7353 , \7352 );
not \U$7011 ( \7354 , \7337 );
not \U$7012 ( \7355 , \7354 );
or \U$7013 ( \7356 , \7353 , \7355 );
not \U$7014 ( \7357 , \855 );
not \U$7015 ( \7358 , \7171 );
or \U$7016 ( \7359 , \7357 , \7358 );
not \U$7017 ( \7360 , RIbb2eda0_19);
not \U$7018 ( \7361 , \5550 );
or \U$7019 ( \7362 , \7360 , \7361 );
not \U$7020 ( \7363 , \2116 );
nand \U$7021 ( \7364 , \7363 , \843 );
nand \U$7022 ( \7365 , \7362 , \7364 );
nand \U$7023 ( \7366 , \7365 , \853 );
nand \U$7024 ( \7367 , \7359 , \7366 );
nand \U$7025 ( \7368 , \7356 , \7367 );
nand \U$7026 ( \7369 , \7351 , \7368 );
and \U$7027 ( \7370 , \7327 , \7369 );
and \U$7028 ( \7371 , \7278 , \7326 );
or \U$7029 ( \7372 , \7370 , \7371 );
xor \U$7030 ( \7373 , \7267 , \7372 );
not \U$7031 ( \7374 , \3613 );
not \U$7032 ( \7375 , \7160 );
or \U$7033 ( \7376 , \7374 , \7375 );
not \U$7034 ( \7377 , RIbb2e800_31);
not \U$7035 ( \7378 , \1550 );
or \U$7036 ( \7379 , \7377 , \7378 );
nand \U$7037 ( \7380 , \1548 , \4096 );
nand \U$7038 ( \7381 , \7379 , \7380 );
nand \U$7039 ( \7382 , \7381 , \2940 );
nand \U$7040 ( \7383 , \7376 , \7382 );
not \U$7041 ( \7384 , \4791 );
not \U$7042 ( \7385 , \7197 );
or \U$7043 ( \7386 , \7384 , \7385 );
not \U$7044 ( \7387 , RIbb2e710_33);
not \U$7045 ( \7388 , \1070 );
or \U$7046 ( \7389 , \7387 , \7388 );
not \U$7047 ( \7390 , RIbb2e710_33);
nand \U$7048 ( \7391 , \1886 , \7390 );
nand \U$7049 ( \7392 , \7389 , \7391 );
nand \U$7050 ( \7393 , \7392 , \3887 );
nand \U$7051 ( \7394 , \7386 , \7393 );
xor \U$7052 ( \7395 , \7383 , \7394 );
not \U$7053 ( \7396 , \2077 );
not \U$7054 ( \7397 , RIbb2ecb0_21);
not \U$7055 ( \7398 , \1340 );
or \U$7056 ( \7399 , \7397 , \7398 );
nand \U$7057 ( \7400 , \6096 , \2249 );
nand \U$7058 ( \7401 , \7399 , \7400 );
not \U$7059 ( \7402 , \7401 );
or \U$7060 ( \7403 , \7396 , \7402 );
nand \U$7061 ( \7404 , \7186 , \2078 );
nand \U$7062 ( \7405 , \7403 , \7404 );
and \U$7063 ( \7406 , \7395 , \7405 );
and \U$7064 ( \7407 , \7383 , \7394 );
or \U$7065 ( \7408 , \7406 , \7407 );
not \U$7066 ( \7409 , \836 );
not \U$7067 ( \7410 , \6994 );
or \U$7068 ( \7411 , \7409 , \7410 );
not \U$7069 ( \7412 , RIbb2ee90_17);
not \U$7070 ( \7413 , \3520 );
or \U$7071 ( \7414 , \7412 , \7413 );
nand \U$7072 ( \7415 , \3343 , \2240 );
nand \U$7073 ( \7416 , \7414 , \7415 );
nand \U$7074 ( \7417 , \7416 , \832 );
nand \U$7075 ( \7418 , \7411 , \7417 );
not \U$7076 ( \7419 , \3465 );
not \U$7077 ( \7420 , \7035 );
or \U$7078 ( \7421 , \7419 , \7420 );
not \U$7079 ( \7422 , RIbb2e9e0_27);
not \U$7080 ( \7423 , \1134 );
buf \U$7081 ( \7424 , \7423 );
not \U$7082 ( \7425 , \7424 );
or \U$7083 ( \7426 , \7422 , \7425 );
not \U$7084 ( \7427 , \7424 );
nand \U$7085 ( \7428 , \7427 , \3454 );
nand \U$7086 ( \7429 , \7426 , \7428 );
nand \U$7087 ( \7430 , \7429 , \3445 );
nand \U$7088 ( \7431 , \7421 , \7430 );
xor \U$7089 ( \7432 , \7418 , \7431 );
not \U$7090 ( \7433 , \1517 );
not \U$7091 ( \7434 , \6983 );
or \U$7092 ( \7435 , \7433 , \7434 );
and \U$7093 ( \7436 , RIbb2ef80_15, \3143 );
not \U$7094 ( \7437 , RIbb2ef80_15);
and \U$7095 ( \7438 , \7437 , \3146 );
or \U$7096 ( \7439 , \7436 , \7438 );
nand \U$7097 ( \7440 , \7439 , \1445 );
nand \U$7098 ( \7441 , \7435 , \7440 );
and \U$7099 ( \7442 , \7432 , \7441 );
and \U$7100 ( \7443 , \7418 , \7431 );
or \U$7101 ( \7444 , \7442 , \7443 );
xor \U$7102 ( \7445 , \7408 , \7444 );
not \U$7103 ( \7446 , \1737 );
not \U$7104 ( \7447 , \7223 );
or \U$7105 ( \7448 , \7446 , \7447 );
not \U$7106 ( \7449 , RIbb2f340_7);
not \U$7107 ( \7450 , \4325 );
or \U$7108 ( \7451 , \7449 , \7450 );
nand \U$7109 ( \7452 , \4324 , \1734 );
nand \U$7110 ( \7453 , \7451 , \7452 );
nand \U$7111 ( \7454 , \7453 , \1702 );
nand \U$7112 ( \7455 , \7448 , \7454 );
not \U$7113 ( \7456 , \3406 );
not \U$7114 ( \7457 , RIbb2ebc0_23);
not \U$7115 ( \7458 , \3116 );
or \U$7116 ( \7459 , \7457 , \7458 );
nand \U$7117 ( \7460 , \1387 , \3401 );
nand \U$7118 ( \7461 , \7459 , \7460 );
not \U$7119 ( \7462 , \7461 );
or \U$7120 ( \7463 , \7456 , \7462 );
nand \U$7121 ( \7464 , \7210 , \3383 );
nand \U$7122 ( \7465 , \7463 , \7464 );
or \U$7123 ( \7466 , \7455 , \7465 );
not \U$7124 ( \7467 , \6242 );
not \U$7125 ( \7468 , \7245 );
or \U$7126 ( \7469 , \7467 , \7468 );
not \U$7127 ( \7470 , RIbb2e530_37);
not \U$7128 ( \7471 , \1509 );
or \U$7129 ( \7472 , \7470 , \7471 );
not \U$7130 ( \7473 , RIbb2e530_37);
nand \U$7131 ( \7474 , \4315 , \7473 );
nand \U$7132 ( \7475 , \7472 , \7474 );
nand \U$7133 ( \7476 , \7475 , \6251 );
nand \U$7134 ( \7477 , \7469 , \7476 );
nand \U$7135 ( \7478 , \7466 , \7477 );
nand \U$7136 ( \7479 , \7455 , \7465 );
nand \U$7137 ( \7480 , \7478 , \7479 );
and \U$7138 ( \7481 , \7445 , \7480 );
and \U$7139 ( \7482 , \7408 , \7444 );
or \U$7140 ( \7483 , \7481 , \7482 );
and \U$7141 ( \7484 , \7373 , \7483 );
and \U$7142 ( \7485 , \7267 , \7372 );
or \U$7143 ( \7486 , \7484 , \7485 );
nand \U$7144 ( \7487 , \7265 , \7486 );
nand \U$7145 ( \7488 , \7264 , \7487 );
not \U$7146 ( \7489 , \7488 );
not \U$7147 ( \7490 , \7489 );
xor \U$7148 ( \7491 , \6813 , \6834 );
not \U$7149 ( \7492 , \6880 );
and \U$7150 ( \7493 , \7491 , \7492 );
not \U$7151 ( \7494 , \7491 );
and \U$7152 ( \7495 , \7494 , \6880 );
nor \U$7153 ( \7496 , \7493 , \7495 );
not \U$7154 ( \7497 , \7496 );
or \U$7155 ( \7498 , \7490 , \7497 );
xor \U$7156 ( \7499 , \6389 , \6397 );
xnor \U$7157 ( \7500 , \7499 , \6364 );
xor \U$7158 ( \7501 , \6514 , \6505 );
xnor \U$7159 ( \7502 , \7501 , \6511 );
xor \U$7160 ( \7503 , \7500 , \7502 );
xor \U$7161 ( \7504 , \7134 , \7139 );
and \U$7162 ( \7505 , \7504 , \7254 );
and \U$7163 ( \7506 , \7134 , \7139 );
or \U$7164 ( \7507 , \7505 , \7506 );
xor \U$7165 ( \7508 , \7503 , \7507 );
nand \U$7166 ( \7509 , \7498 , \7508 );
not \U$7167 ( \7510 , \7496 );
nand \U$7168 ( \7511 , \7510 , \7488 );
nand \U$7169 ( \7512 , \7509 , \7511 );
nand \U$7170 ( \7513 , \7083 , \7512 );
nand \U$7171 ( \7514 , \7082 , \7513 );
xor \U$7172 ( \7515 , \6421 , \6399 );
xor \U$7173 ( \7516 , \7515 , \6343 );
xor \U$7174 ( \7517 , \6516 , \6470 );
xnor \U$7175 ( \7518 , \7517 , \6522 );
xor \U$7176 ( \7519 , \7516 , \7518 );
xor \U$7177 ( \7520 , \7500 , \7502 );
and \U$7178 ( \7521 , \7520 , \7507 );
and \U$7179 ( \7522 , \7500 , \7502 );
or \U$7180 ( \7523 , \7521 , \7522 );
and \U$7181 ( \7524 , \7519 , \7523 );
and \U$7182 ( \7525 , \7516 , \7518 );
or \U$7183 ( \7526 , \7524 , \7525 );
or \U$7184 ( \7527 , \7514 , \7526 );
xor \U$7185 ( \7528 , \6884 , \6886 );
xor \U$7186 ( \7529 , \7528 , \6889 );
nand \U$7187 ( \7530 , \7527 , \7529 );
nand \U$7188 ( \7531 , \7514 , \7526 );
nand \U$7189 ( \7532 , \7530 , \7531 );
or \U$7190 ( \7533 , \6903 , \7532 );
nand \U$7191 ( \7534 , \6901 , \7533 );
nor \U$7192 ( \7535 , \6573 , \7534 );
not \U$7193 ( \7536 , \6562 );
not \U$7194 ( \7537 , \7536 );
not \U$7195 ( \7538 , \6559 );
or \U$7196 ( \7539 , \7537 , \7538 );
or \U$7197 ( \7540 , \7536 , \6559 );
nand \U$7198 ( \7541 , \7540 , \6570 );
nand \U$7199 ( \7542 , \7539 , \7541 );
xor \U$7200 ( \7543 , \3863 , \4513 );
xor \U$7201 ( \7544 , \7543 , \4862 );
or \U$7202 ( \7545 , \7542 , \7544 );
nand \U$7203 ( \7546 , \7535 , \7545 );
nor \U$7204 ( \7547 , \5824 , \7546 );
not \U$7205 ( \7548 , \1570 );
and \U$7206 ( \7549 , \1139 , RIbb2f250_9);
not \U$7207 ( \7550 , \1139 );
and \U$7208 ( \7551 , \7550 , \1554 );
nor \U$7209 ( \7552 , \7549 , \7551 );
not \U$7210 ( \7553 , \7552 );
or \U$7211 ( \7554 , \7548 , \7553 );
and \U$7212 ( \7555 , RIbb2f250_9, \1114 );
not \U$7213 ( \7556 , RIbb2f250_9);
and \U$7214 ( \7557 , \7556 , \1113 );
nor \U$7215 ( \7558 , \7555 , \7557 );
nand \U$7216 ( \7559 , \7558 , \1533 );
nand \U$7217 ( \7560 , \7554 , \7559 );
and \U$7218 ( \7561 , RIbb2ef80_15, \1562 );
not \U$7219 ( \7562 , RIbb2ef80_15);
and \U$7220 ( \7563 , \7562 , \1563 );
nor \U$7221 ( \7564 , \7561 , \7563 );
or \U$7222 ( \7565 , \7564 , \1575 );
or \U$7223 ( \7566 , \2265 , \1584 );
nand \U$7224 ( \7567 , \7565 , \7566 );
xor \U$7225 ( \7568 , \7560 , \7567 );
not \U$7226 ( \7569 , \1737 );
not \U$7227 ( \7570 , \2283 );
or \U$7228 ( \7571 , \7569 , \7570 );
not \U$7229 ( \7572 , RIbb2f340_7);
not \U$7230 ( \7573 , \1171 );
or \U$7231 ( \7574 , \7572 , \7573 );
nand \U$7232 ( \7575 , \1248 , \2700 );
nand \U$7233 ( \7576 , \7574 , \7575 );
not \U$7234 ( \7577 , \7576 );
or \U$7235 ( \7578 , \7577 , \1703 );
nand \U$7236 ( \7579 , \7571 , \7578 );
and \U$7237 ( \7580 , \7568 , \7579 );
and \U$7238 ( \7581 , \7560 , \7567 );
or \U$7239 ( \7582 , \7580 , \7581 );
xor \U$7240 ( \7583 , \2226 , \2232 );
xor \U$7241 ( \7584 , \7583 , \2245 );
xor \U$7242 ( \7585 , \7582 , \7584 );
and \U$7243 ( \7586 , \1689 , RIbb2f160_11);
and \U$7244 ( \7587 , \1691 , \1043 );
nor \U$7245 ( \7588 , \7586 , \7587 );
or \U$7246 ( \7589 , \7588 , \2122 );
or \U$7247 ( \7590 , \2121 , \1943 );
nand \U$7248 ( \7591 , \7589 , \7590 );
xor \U$7249 ( \7592 , \7591 , \2259 );
not \U$7250 ( \7593 , \1533 );
not \U$7251 ( \7594 , \7552 );
or \U$7252 ( \7595 , \7593 , \7594 );
or \U$7253 ( \7596 , \2130 , \2133 );
nand \U$7254 ( \7597 , \7595 , \7596 );
xor \U$7255 ( \7598 , \7592 , \7597 );
xor \U$7256 ( \7599 , \7585 , \7598 );
xor \U$7257 ( \7600 , \2268 , \2277 );
xor \U$7258 ( \7601 , \7600 , \2287 );
not \U$7259 ( \7602 , \916 );
and \U$7260 ( \7603 , \1551 , RIbb2f070_13);
not \U$7261 ( \7604 , \1551 );
and \U$7262 ( \7605 , \7604 , \1656 );
nor \U$7263 ( \7606 , \7603 , \7605 );
not \U$7264 ( \7607 , \7606 );
or \U$7265 ( \7608 , \7602 , \7607 );
or \U$7266 ( \7609 , \2149 , \1662 );
nand \U$7267 ( \7610 , \7608 , \7609 );
not \U$7268 ( \7611 , \1090 );
and \U$7269 ( \7612 , \1387 , RIbb2f430_5);
not \U$7270 ( \7613 , \1387 );
and \U$7271 ( \7614 , \7613 , \1898 );
nor \U$7272 ( \7615 , \7612 , \7614 );
not \U$7273 ( \7616 , \7615 );
or \U$7274 ( \7617 , \7611 , \7616 );
or \U$7275 ( \7618 , \2156 , \1650 );
nand \U$7276 ( \7619 , \7617 , \7618 );
xor \U$7277 ( \7620 , \7610 , \7619 );
and \U$7278 ( \7621 , \1340 , \1290 );
and \U$7279 ( \7622 , \1341 , \1289 );
nor \U$7280 ( \7623 , \7621 , \7622 );
or \U$7281 ( \7624 , \7623 , \1266 );
or \U$7282 ( \7625 , \2055 , \1295 );
nand \U$7283 ( \7626 , \7624 , \7625 );
xor \U$7284 ( \7627 , \7620 , \7626 );
not \U$7285 ( \7628 , \3407 );
and \U$7286 ( \7629 , RIbb2ebc0_23, \815 );
not \U$7287 ( \7630 , RIbb2ebc0_23);
and \U$7288 ( \7631 , \7630 , \814 );
nor \U$7289 ( \7632 , \7629 , \7631 );
not \U$7290 ( \7633 , \7632 );
or \U$7291 ( \7634 , \7628 , \7633 );
not \U$7292 ( \7635 , \3383 );
or \U$7293 ( \7636 , \7635 , \3401 );
nand \U$7294 ( \7637 , \7634 , \7636 );
not \U$7295 ( \7638 , RIbb2f160_11);
not \U$7296 ( \7639 , \1644 );
or \U$7297 ( \7640 , \7638 , \7639 );
nand \U$7298 ( \7641 , \1646 , \1805 );
nand \U$7299 ( \7642 , \7640 , \7641 );
not \U$7300 ( \7643 , \7642 );
or \U$7301 ( \7644 , \7643 , \2122 );
or \U$7302 ( \7645 , \7588 , \1943 );
nand \U$7303 ( \7646 , \7644 , \7645 );
xor \U$7304 ( \7647 , \7637 , \7646 );
not \U$7305 ( \7648 , \1090 );
and \U$7306 ( \7649 , \1647 , \1340 );
not \U$7307 ( \7650 , \1647 );
and \U$7308 ( \7651 , \7650 , \1341 );
nor \U$7309 ( \7652 , \7649 , \7651 );
not \U$7310 ( \7653 , \7652 );
or \U$7311 ( \7654 , \7648 , \7653 );
not \U$7312 ( \7655 , RIbb2f430_5);
not \U$7313 ( \7656 , \2052 );
or \U$7314 ( \7657 , \7655 , \7656 );
nand \U$7315 ( \7658 , \1422 , \1898 );
nand \U$7316 ( \7659 , \7657 , \7658 );
nand \U$7317 ( \7660 , \7659 , \1147 );
nand \U$7318 ( \7661 , \7654 , \7660 );
not \U$7319 ( \7662 , \1702 );
not \U$7320 ( \7663 , RIbb2f340_7);
not \U$7321 ( \7664 , \1820 );
or \U$7322 ( \7665 , \7663 , \7664 );
nand \U$7323 ( \7666 , \1387 , \1734 );
nand \U$7324 ( \7667 , \7665 , \7666 );
not \U$7325 ( \7668 , \7667 );
or \U$7326 ( \7669 , \7662 , \7668 );
nand \U$7327 ( \7670 , \7576 , \1737 );
nand \U$7328 ( \7671 , \7669 , \7670 );
xor \U$7329 ( \7672 , \7661 , \7671 );
and \U$7330 ( \7673 , RIbb2ef80_15, \1551 );
not \U$7331 ( \7674 , RIbb2ef80_15);
and \U$7332 ( \7675 , \7674 , \1550 );
nor \U$7333 ( \7676 , \7673 , \7675 );
not \U$7334 ( \7677 , \7676 );
not \U$7335 ( \7678 , \1445 );
or \U$7336 ( \7679 , \7677 , \7678 );
or \U$7337 ( \7680 , \7564 , \1584 );
nand \U$7338 ( \7681 , \7679 , \7680 );
and \U$7339 ( \7682 , \7672 , \7681 );
and \U$7340 ( \7683 , \7661 , \7671 );
or \U$7341 ( \7684 , \7682 , \7683 );
and \U$7342 ( \7685 , \7647 , \7684 );
and \U$7343 ( \7686 , \7637 , \7646 );
or \U$7344 ( \7687 , \7685 , \7686 );
xor \U$7345 ( \7688 , \7627 , \7687 );
xor \U$7346 ( \7689 , \7601 , \7688 );
xor \U$7347 ( \7690 , \7599 , \7689 );
and \U$7348 ( \7691 , \1313 , \3347 );
not \U$7349 ( \7692 , \998 );
not \U$7350 ( \7693 , \7606 );
or \U$7351 ( \7694 , \7692 , \7693 );
not \U$7352 ( \7695 , RIbb2f070_13);
not \U$7353 ( \7696 , \1731 );
or \U$7354 ( \7697 , \7695 , \7696 );
nand \U$7355 ( \7698 , \1733 , \1656 );
nand \U$7356 ( \7699 , \7697 , \7698 );
nand \U$7357 ( \7700 , \7699 , \916 );
nand \U$7358 ( \7701 , \7694 , \7700 );
xor \U$7359 ( \7702 , \7691 , \7701 );
not \U$7360 ( \7703 , \1430 );
xor \U$7361 ( \7704 , \1313 , \2225 );
not \U$7362 ( \7705 , \7704 );
or \U$7363 ( \7706 , \7703 , \7705 );
not \U$7364 ( \7707 , \2230 );
or \U$7365 ( \7708 , \7707 , \1954 );
nand \U$7366 ( \7709 , \7706 , \7708 );
xor \U$7367 ( \7710 , \7702 , \7709 );
xor \U$7368 ( \7711 , \7637 , \7646 );
xor \U$7369 ( \7712 , \7711 , \7684 );
xor \U$7370 ( \7713 , \7710 , \7712 );
not \U$7371 ( \7714 , \7637 );
not \U$7372 ( \7715 , \1570 );
and \U$7373 ( \7716 , RIbb2f250_9, \1285 );
not \U$7374 ( \7717 , RIbb2f250_9);
and \U$7375 ( \7718 , \7717 , \1284 );
nor \U$7376 ( \7719 , \7716 , \7718 );
not \U$7377 ( \7720 , \7719 );
or \U$7378 ( \7721 , \7715 , \7720 );
not \U$7379 ( \7722 , \5617 );
or \U$7380 ( \7723 , \7722 , \1771 );
nand \U$7381 ( \7724 , \7721 , \7723 );
not \U$7382 ( \7725 , \836 );
not \U$7383 ( \7726 , RIbb2ee90_17);
not \U$7384 ( \7727 , \1072 );
or \U$7385 ( \7728 , \7726 , \7727 );
nand \U$7386 ( \7729 , \1888 , \816 );
nand \U$7387 ( \7730 , \7728 , \7729 );
not \U$7388 ( \7731 , \7730 );
or \U$7389 ( \7732 , \7725 , \7731 );
nand \U$7390 ( \7733 , \5580 , \832 );
nand \U$7391 ( \7734 , \7732 , \7733 );
xor \U$7392 ( \7735 , \7724 , \7734 );
not \U$7393 ( \7736 , \1011 );
not \U$7394 ( \7737 , \5525 );
or \U$7395 ( \7738 , \7736 , \7737 );
not \U$7396 ( \7739 , RIbb2f160_11);
not \U$7397 ( \7740 , \1140 );
or \U$7398 ( \7741 , \7739 , \7740 );
nand \U$7399 ( \7742 , \1139 , \1048 );
nand \U$7400 ( \7743 , \7741 , \7742 );
nand \U$7401 ( \7744 , \7743 , \1077 );
nand \U$7402 ( \7745 , \7738 , \7744 );
and \U$7403 ( \7746 , \7735 , \7745 );
and \U$7404 ( \7747 , \7724 , \7734 );
or \U$7405 ( \7748 , \7746 , \7747 );
xor \U$7406 ( \7749 , \7714 , \7748 );
not \U$7407 ( \7750 , \1737 );
not \U$7408 ( \7751 , \7667 );
or \U$7409 ( \7752 , \7750 , \7751 );
nand \U$7410 ( \7753 , \5601 , \1702 );
nand \U$7411 ( \7754 , \7752 , \7753 );
not \U$7412 ( \7755 , \1147 );
not \U$7413 ( \7756 , \7652 );
or \U$7414 ( \7757 , \7755 , \7756 );
not \U$7415 ( \7758 , \5561 );
or \U$7416 ( \7759 , \7758 , \1621 );
nand \U$7417 ( \7760 , \7757 , \7759 );
xor \U$7418 ( \7761 , \7754 , \7760 );
not \U$7419 ( \7762 , \5489 );
not \U$7420 ( \7763 , \2077 );
or \U$7421 ( \7764 , \7762 , \7763 );
and \U$7422 ( \7765 , \1514 , RIbb2ecb0_21);
and \U$7423 ( \7766 , \1511 , \5481 );
nor \U$7424 ( \7767 , \7765 , \7766 );
not \U$7425 ( \7768 , \2078 );
or \U$7426 ( \7769 , \7767 , \7768 );
nand \U$7427 ( \7770 , \7764 , \7769 );
and \U$7428 ( \7771 , \7761 , \7770 );
and \U$7429 ( \7772 , \7754 , \7760 );
or \U$7430 ( \7773 , \7771 , \7772 );
and \U$7431 ( \7774 , \7749 , \7773 );
and \U$7432 ( \7775 , \7714 , \7748 );
or \U$7433 ( \7776 , \7774 , \7775 );
and \U$7434 ( \7777 , \7713 , \7776 );
and \U$7435 ( \7778 , \7710 , \7712 );
or \U$7436 ( \7779 , \7777 , \7778 );
xor \U$7437 ( \7780 , \7690 , \7779 );
xor \U$7438 ( \7781 , \7710 , \7712 );
xor \U$7439 ( \7782 , \7781 , \7776 );
or \U$7440 ( \7783 , \2980 , \2963 );
nand \U$7441 ( \7784 , \7783 , RIbb2ead0_25);
not \U$7442 ( \7785 , \3407 );
not \U$7443 ( \7786 , \5509 );
or \U$7444 ( \7787 , \7785 , \7786 );
nand \U$7445 ( \7788 , \7632 , \3383 );
nand \U$7446 ( \7789 , \7787 , \7788 );
xor \U$7447 ( \7790 , \7784 , \7789 );
not \U$7448 ( \7791 , \855 );
and \U$7449 ( \7792 , RIbb2eda0_19, \1940 );
not \U$7450 ( \7793 , RIbb2eda0_19);
and \U$7451 ( \7794 , \7793 , \989 );
nor \U$7452 ( \7795 , \7792 , \7794 );
not \U$7453 ( \7796 , \7795 );
or \U$7454 ( \7797 , \7791 , \7796 );
nand \U$7455 ( \7798 , \5499 , \853 );
nand \U$7456 ( \7799 , \7797 , \7798 );
and \U$7457 ( \7800 , \7790 , \7799 );
and \U$7458 ( \7801 , \7784 , \7789 );
or \U$7459 ( \7802 , \7800 , \7801 );
not \U$7460 ( \7803 , \1376 );
xor \U$7461 ( \7804 , \1313 , \3347 );
not \U$7462 ( \7805 , \7804 );
or \U$7463 ( \7806 , \7803 , \7805 );
nand \U$7464 ( \7807 , \5473 , \1430 );
nand \U$7465 ( \7808 , \7806 , \7807 );
not \U$7466 ( \7809 , \1294 );
not \U$7467 ( \7810 , \1290 );
not \U$7468 ( \7811 , \2116 );
or \U$7469 ( \7812 , \7810 , \7811 );
nand \U$7470 ( \7813 , \2117 , \1291 );
nand \U$7471 ( \7814 , \7812 , \7813 );
not \U$7472 ( \7815 , \7814 );
or \U$7473 ( \7816 , \7809 , \7815 );
nand \U$7474 ( \7817 , \5539 , \1265 );
nand \U$7475 ( \7818 , \7816 , \7817 );
xor \U$7476 ( \7819 , \7808 , \7818 );
not \U$7477 ( \7820 , \1517 );
not \U$7478 ( \7821 , \7676 );
or \U$7479 ( \7822 , \7820 , \7821 );
nand \U$7480 ( \7823 , \5571 , \1445 );
nand \U$7481 ( \7824 , \7822 , \7823 );
and \U$7482 ( \7825 , \7819 , \7824 );
and \U$7483 ( \7826 , \7808 , \7818 );
or \U$7484 ( \7827 , \7825 , \7826 );
xor \U$7485 ( \7828 , \7802 , \7827 );
and \U$7486 ( \7829 , \1394 , \4220 );
not \U$7487 ( \7830 , \1011 );
not \U$7488 ( \7831 , \7743 );
or \U$7489 ( \7832 , \7830 , \7831 );
nand \U$7490 ( \7833 , \7642 , \1077 );
nand \U$7491 ( \7834 , \7832 , \7833 );
xor \U$7492 ( \7835 , \7829 , \7834 );
not \U$7493 ( \7836 , \853 );
not \U$7494 ( \7837 , \7795 );
or \U$7495 ( \7838 , \7836 , \7837 );
not \U$7496 ( \7839 , RIbb2eda0_19);
not \U$7497 ( \7840 , \1659 );
or \U$7498 ( \7841 , \7839 , \7840 );
nand \U$7499 ( \7842 , \1477 , \1776 );
nand \U$7500 ( \7843 , \7841 , \7842 );
not \U$7501 ( \7844 , \7843 );
or \U$7502 ( \7845 , \7844 , \1781 );
nand \U$7503 ( \7846 , \7838 , \7845 );
xor \U$7504 ( \7847 , \7835 , \7846 );
and \U$7505 ( \7848 , \7828 , \7847 );
and \U$7506 ( \7849 , \7802 , \7827 );
or \U$7507 ( \7850 , \7848 , \7849 );
not \U$7508 ( \7851 , \916 );
not \U$7509 ( \7852 , RIbb2f070_13);
not \U$7510 ( \7853 , \1689 );
or \U$7511 ( \7854 , \7852 , \7853 );
nand \U$7512 ( \7855 , \1691 , \3421 );
nand \U$7513 ( \7856 , \7854 , \7855 );
not \U$7514 ( \7857 , \7856 );
or \U$7515 ( \7858 , \7851 , \7857 );
nand \U$7516 ( \7859 , \7699 , \998 );
nand \U$7517 ( \7860 , \7858 , \7859 );
not \U$7518 ( \7861 , \1430 );
not \U$7519 ( \7862 , \7804 );
or \U$7520 ( \7863 , \7861 , \7862 );
nand \U$7521 ( \7864 , \7704 , \1376 );
nand \U$7522 ( \7865 , \7863 , \7864 );
xor \U$7523 ( \7866 , \7860 , \7865 );
not \U$7524 ( \7867 , \1265 );
not \U$7525 ( \7868 , \7814 );
or \U$7526 ( \7869 , \7867 , \7868 );
not \U$7527 ( \7870 , \1290 );
not \U$7528 ( \7871 , \1854 );
or \U$7529 ( \7872 , \7870 , \7871 );
nand \U$7530 ( \7873 , \1855 , \1291 );
nand \U$7531 ( \7874 , \7872 , \7873 );
nand \U$7532 ( \7875 , \7874 , \1294 );
nand \U$7533 ( \7876 , \7869 , \7875 );
xor \U$7534 ( \7877 , \7866 , \7876 );
xor \U$7535 ( \7878 , \7661 , \7671 );
xor \U$7536 ( \7879 , \7878 , \7681 );
xor \U$7537 ( \7880 , \7877 , \7879 );
not \U$7538 ( \7881 , \836 );
not \U$7539 ( \7882 , RIbb2ee90_17);
not \U$7540 ( \7883 , \953 );
or \U$7541 ( \7884 , \7882 , \7883 );
nand \U$7542 ( \7885 , \957 , \816 );
nand \U$7543 ( \7886 , \7884 , \7885 );
not \U$7544 ( \7887 , \7886 );
or \U$7545 ( \7888 , \7881 , \7887 );
nand \U$7546 ( \7889 , \7730 , \832 );
nand \U$7547 ( \7890 , \7888 , \7889 );
not \U$7548 ( \7891 , \1533 );
not \U$7549 ( \7892 , \7719 );
or \U$7550 ( \7893 , \7891 , \7892 );
nand \U$7551 ( \7894 , \7558 , \1570 );
nand \U$7552 ( \7895 , \7893 , \7894 );
xor \U$7553 ( \7896 , \7890 , \7895 );
or \U$7554 ( \7897 , \7767 , \7763 );
and \U$7555 ( \7898 , \2067 , \2081 );
not \U$7556 ( \7899 , \2067 );
and \U$7557 ( \7900 , \7899 , \898 );
nor \U$7558 ( \7901 , \7898 , \7900 );
not \U$7559 ( \7902 , \7901 );
or \U$7560 ( \7903 , \7902 , \7768 );
nand \U$7561 ( \7904 , \7897 , \7903 );
xor \U$7562 ( \7905 , \7896 , \7904 );
and \U$7563 ( \7906 , \7880 , \7905 );
and \U$7564 ( \7907 , \7877 , \7879 );
or \U$7565 ( \7908 , \7906 , \7907 );
xor \U$7566 ( \7909 , \7850 , \7908 );
xor \U$7567 ( \7910 , \7860 , \7865 );
and \U$7568 ( \7911 , \7910 , \7876 );
and \U$7569 ( \7912 , \7860 , \7865 );
or \U$7570 ( \7913 , \7911 , \7912 );
xor \U$7571 ( \7914 , \7890 , \7895 );
and \U$7572 ( \7915 , \7914 , \7904 );
and \U$7573 ( \7916 , \7890 , \7895 );
or \U$7574 ( \7917 , \7915 , \7916 );
xor \U$7575 ( \7918 , \7913 , \7917 );
xor \U$7576 ( \7919 , \7829 , \7834 );
and \U$7577 ( \7920 , \7919 , \7846 );
and \U$7578 ( \7921 , \7829 , \7834 );
or \U$7579 ( \7922 , \7920 , \7921 );
xor \U$7580 ( \7923 , \7918 , \7922 );
xor \U$7581 ( \7924 , \7909 , \7923 );
xor \U$7582 ( \7925 , \7782 , \7924 );
xor \U$7583 ( \7926 , \7877 , \7879 );
xor \U$7584 ( \7927 , \7926 , \7905 );
not \U$7585 ( \7928 , \5753 );
not \U$7586 ( \7929 , \5739 );
or \U$7587 ( \7930 , \7928 , \7929 );
or \U$7588 ( \7931 , \5739 , \5753 );
nand \U$7589 ( \7932 , \7931 , \5745 );
nand \U$7590 ( \7933 , \7930 , \7932 );
xor \U$7591 ( \7934 , \5716 , \5727 );
and \U$7592 ( \7935 , \7934 , \5734 );
and \U$7593 ( \7936 , \5716 , \5727 );
or \U$7594 ( \7937 , \7935 , \7936 );
xor \U$7595 ( \7938 , \7933 , \7937 );
not \U$7596 ( \7939 , \5547 );
not \U$7597 ( \7940 , \5563 );
or \U$7598 ( \7941 , \7939 , \7940 );
or \U$7599 ( \7942 , \5563 , \5547 );
nand \U$7600 ( \7943 , \7942 , \5573 );
nand \U$7601 ( \7944 , \7941 , \7943 );
xor \U$7602 ( \7945 , \5588 , \5603 );
and \U$7603 ( \7946 , \7945 , \5619 );
and \U$7604 ( \7947 , \5588 , \5603 );
or \U$7605 ( \7948 , \7946 , \7947 );
xor \U$7606 ( \7949 , \7944 , \7948 );
xor \U$7607 ( \7950 , \5503 , \5518 );
and \U$7608 ( \7951 , \7950 , \5529 );
and \U$7609 ( \7952 , \5503 , \5518 );
or \U$7610 ( \7953 , \7951 , \7952 );
xor \U$7611 ( \7954 , \7949 , \7953 );
and \U$7612 ( \7955 , \7938 , \7954 );
and \U$7613 ( \7956 , \7933 , \7937 );
or \U$7614 ( \7957 , \7955 , \7956 );
xor \U$7615 ( \7958 , \7927 , \7957 );
and \U$7616 ( \7959 , \1313 , \5028 );
xor \U$7617 ( \7960 , \7959 , \5715 );
not \U$7618 ( \7961 , \998 );
not \U$7619 ( \7962 , \7856 );
or \U$7620 ( \7963 , \7961 , \7962 );
nand \U$7621 ( \7964 , \5722 , \916 );
nand \U$7622 ( \7965 , \7963 , \7964 );
and \U$7623 ( \7966 , \7960 , \7965 );
and \U$7624 ( \7967 , \7959 , \5715 );
or \U$7625 ( \7968 , \7966 , \7967 );
xor \U$7626 ( \7969 , \7944 , \7948 );
and \U$7627 ( \7970 , \7969 , \7953 );
and \U$7628 ( \7971 , \7944 , \7948 );
or \U$7629 ( \7972 , \7970 , \7971 );
xor \U$7630 ( \7973 , \7968 , \7972 );
xor \U$7631 ( \7974 , \7714 , \7748 );
xor \U$7632 ( \7975 , \7974 , \7773 );
xor \U$7633 ( \7976 , \7973 , \7975 );
and \U$7634 ( \7977 , \7958 , \7976 );
and \U$7635 ( \7978 , \7927 , \7957 );
or \U$7636 ( \7979 , \7977 , \7978 );
and \U$7637 ( \7980 , \7925 , \7979 );
and \U$7638 ( \7981 , \7782 , \7924 );
or \U$7639 ( \7982 , \7980 , \7981 );
xor \U$7640 ( \7983 , \7780 , \7982 );
xor \U$7641 ( \7984 , \7913 , \7917 );
and \U$7642 ( \7985 , \7984 , \7922 );
and \U$7643 ( \7986 , \7913 , \7917 );
or \U$7644 ( \7987 , \7985 , \7986 );
or \U$7645 ( \7988 , \3407 , \3383 );
nand \U$7646 ( \7989 , \7988 , RIbb2ebc0_23);
not \U$7647 ( \7990 , \2077 );
not \U$7648 ( \7991 , \7901 );
or \U$7649 ( \7992 , \7990 , \7991 );
nand \U$7650 ( \7993 , \2256 , \2078 );
nand \U$7651 ( \7994 , \7992 , \7993 );
xor \U$7652 ( \7995 , \7989 , \7994 );
not \U$7653 ( \7996 , \832 );
not \U$7654 ( \7997 , \7886 );
or \U$7655 ( \7998 , \7996 , \7997 );
nand \U$7656 ( \7999 , \2242 , \836 );
nand \U$7657 ( \8000 , \7998 , \7999 );
xor \U$7658 ( \8001 , \7995 , \8000 );
not \U$7659 ( \8002 , \855 );
not \U$7660 ( \8003 , \2273 );
or \U$7661 ( \8004 , \8002 , \8003 );
nand \U$7662 ( \8005 , \7843 , \853 );
nand \U$7663 ( \8006 , \8004 , \8005 );
not \U$7664 ( \8007 , \1147 );
not \U$7665 ( \8008 , \7615 );
or \U$7666 ( \8009 , \8007 , \8008 );
nand \U$7667 ( \8010 , \7659 , \1090 );
nand \U$7668 ( \8011 , \8009 , \8010 );
xor \U$7669 ( \8012 , \8006 , \8011 );
not \U$7670 ( \8013 , \1265 );
not \U$7671 ( \8014 , \7874 );
or \U$7672 ( \8015 , \8013 , \8014 );
or \U$7673 ( \8016 , \7623 , \1295 );
nand \U$7674 ( \8017 , \8015 , \8016 );
xor \U$7675 ( \8018 , \8012 , \8017 );
xor \U$7676 ( \8019 , \8001 , \8018 );
xor \U$7677 ( \8020 , \7560 , \7567 );
xor \U$7678 ( \8021 , \8020 , \7579 );
and \U$7679 ( \8022 , \8019 , \8021 );
and \U$7680 ( \8023 , \8001 , \8018 );
or \U$7681 ( \8024 , \8022 , \8023 );
xor \U$7682 ( \8025 , \7987 , \8024 );
xor \U$7683 ( \8026 , \7691 , \7701 );
and \U$7684 ( \8027 , \8026 , \7709 );
and \U$7685 ( \8028 , \7691 , \7701 );
or \U$7686 ( \8029 , \8027 , \8028 );
xor \U$7687 ( \8030 , \7989 , \7994 );
and \U$7688 ( \8031 , \8030 , \8000 );
and \U$7689 ( \8032 , \7989 , \7994 );
or \U$7690 ( \8033 , \8031 , \8032 );
xor \U$7691 ( \8034 , \8029 , \8033 );
xor \U$7692 ( \8035 , \8006 , \8011 );
and \U$7693 ( \8036 , \8035 , \8017 );
and \U$7694 ( \8037 , \8006 , \8011 );
or \U$7695 ( \8038 , \8036 , \8037 );
xor \U$7696 ( \8039 , \8034 , \8038 );
xor \U$7697 ( \8040 , \8025 , \8039 );
xor \U$7698 ( \8041 , \7850 , \7908 );
and \U$7699 ( \8042 , \8041 , \7923 );
and \U$7700 ( \8043 , \7850 , \7908 );
or \U$7701 ( \8044 , \8042 , \8043 );
xor \U$7702 ( \8045 , \8040 , \8044 );
xor \U$7703 ( \8046 , \8001 , \8018 );
xor \U$7704 ( \8047 , \8046 , \8021 );
xor \U$7705 ( \8048 , \7968 , \7972 );
and \U$7706 ( \8049 , \8048 , \7975 );
and \U$7707 ( \8050 , \7968 , \7972 );
or \U$7708 ( \8051 , \8049 , \8050 );
xor \U$7709 ( \8052 , \8047 , \8051 );
xor \U$7710 ( \8053 , \5469 , \5475 );
and \U$7711 ( \8054 , \8053 , \5491 );
and \U$7712 ( \8055 , \5469 , \5475 );
or \U$7713 ( \8056 , \8054 , \8055 );
xor \U$7714 ( \8057 , \7959 , \5715 );
xor \U$7715 ( \8058 , \8057 , \7965 );
xor \U$7716 ( \8059 , \8056 , \8058 );
xor \U$7717 ( \8060 , \7724 , \7734 );
xor \U$7718 ( \8061 , \8060 , \7745 );
and \U$7719 ( \8062 , \8059 , \8061 );
and \U$7720 ( \8063 , \8056 , \8058 );
or \U$7721 ( \8064 , \8062 , \8063 );
xor \U$7722 ( \8065 , \7802 , \7827 );
xor \U$7723 ( \8066 , \8065 , \7847 );
xor \U$7724 ( \8067 , \8064 , \8066 );
xor \U$7725 ( \8068 , \7784 , \7789 );
xor \U$7726 ( \8069 , \8068 , \7799 );
xor \U$7727 ( \8070 , \7808 , \7818 );
xor \U$7728 ( \8071 , \8070 , \7824 );
xor \U$7729 ( \8072 , \8069 , \8071 );
xor \U$7730 ( \8073 , \7754 , \7760 );
xor \U$7731 ( \8074 , \8073 , \7770 );
and \U$7732 ( \8075 , \8072 , \8074 );
and \U$7733 ( \8076 , \8069 , \8071 );
or \U$7734 ( \8077 , \8075 , \8076 );
and \U$7735 ( \8078 , \8067 , \8077 );
and \U$7736 ( \8079 , \8064 , \8066 );
or \U$7737 ( \8080 , \8078 , \8079 );
and \U$7738 ( \8081 , \8052 , \8080 );
and \U$7739 ( \8082 , \8047 , \8051 );
or \U$7740 ( \8083 , \8081 , \8082 );
xor \U$7741 ( \8084 , \8045 , \8083 );
xor \U$7742 ( \8085 , \7983 , \8084 );
xor \U$7743 ( \8086 , \8047 , \8051 );
xor \U$7744 ( \8087 , \8086 , \8080 );
xor \U$7745 ( \8088 , \7782 , \7924 );
xor \U$7746 ( \8089 , \8088 , \7979 );
or \U$7747 ( \8090 , \8087 , \8089 );
xor \U$7748 ( \8091 , \5468 , \5492 );
and \U$7749 ( \8092 , \8091 , \5530 );
and \U$7750 ( \8093 , \5468 , \5492 );
or \U$7751 ( \8094 , \8092 , \8093 );
xor \U$7752 ( \8095 , \8056 , \8058 );
xor \U$7753 ( \8096 , \8095 , \8061 );
xor \U$7754 ( \8097 , \8094 , \8096 );
xor \U$7755 ( \8098 , \8069 , \8071 );
xor \U$7756 ( \8099 , \8098 , \8074 );
and \U$7757 ( \8100 , \8097 , \8099 );
and \U$7758 ( \8101 , \8094 , \8096 );
or \U$7759 ( \8102 , \8100 , \8101 );
xor \U$7760 ( \8103 , \8064 , \8066 );
xor \U$7761 ( \8104 , \8103 , \8077 );
xor \U$7762 ( \8105 , \8102 , \8104 );
xor \U$7763 ( \8106 , \5574 , \5620 );
and \U$7764 ( \8107 , \8106 , \5625 );
and \U$7765 ( \8108 , \5574 , \5620 );
or \U$7766 ( \8109 , \8107 , \8108 );
xor \U$7767 ( \8110 , \5735 , \5754 );
and \U$7768 ( \8111 , \8110 , \5759 );
and \U$7769 ( \8112 , \5735 , \5754 );
or \U$7770 ( \8113 , \8111 , \8112 );
xor \U$7771 ( \8114 , \8109 , \8113 );
xor \U$7772 ( \8115 , \7933 , \7937 );
xor \U$7773 ( \8116 , \8115 , \7954 );
and \U$7774 ( \8117 , \8114 , \8116 );
and \U$7775 ( \8118 , \8109 , \8113 );
or \U$7776 ( \8119 , \8117 , \8118 );
and \U$7777 ( \8120 , \8105 , \8119 );
and \U$7778 ( \8121 , \8102 , \8104 );
or \U$7779 ( \8122 , \8120 , \8121 );
nand \U$7780 ( \8123 , \8090 , \8122 );
nand \U$7781 ( \8124 , \8089 , \8087 );
nand \U$7782 ( \8125 , \8123 , \8124 );
or \U$7783 ( \8126 , \8085 , \8125 );
xor \U$7784 ( \8127 , \7927 , \7957 );
xor \U$7785 ( \8128 , \8127 , \7976 );
xor \U$7786 ( \8129 , \5451 , \5531 );
and \U$7787 ( \8130 , \8129 , \5626 );
and \U$7788 ( \8131 , \5451 , \5531 );
or \U$7789 ( \8132 , \8130 , \8131 );
xor \U$7790 ( \8133 , \8094 , \8096 );
xor \U$7791 ( \8134 , \8133 , \8099 );
xor \U$7792 ( \8135 , \8132 , \8134 );
xor \U$7793 ( \8136 , \8109 , \8113 );
xor \U$7794 ( \8137 , \8136 , \8116 );
and \U$7795 ( \8138 , \8135 , \8137 );
and \U$7796 ( \8139 , \8132 , \8134 );
or \U$7797 ( \8140 , \8138 , \8139 );
xor \U$7798 ( \8141 , \8128 , \8140 );
xor \U$7799 ( \8142 , \8102 , \8104 );
xor \U$7800 ( \8143 , \8142 , \8119 );
and \U$7801 ( \8144 , \8141 , \8143 );
and \U$7802 ( \8145 , \8128 , \8140 );
or \U$7803 ( \8146 , \8144 , \8145 );
not \U$7804 ( \8147 , \8146 );
xor \U$7805 ( \8148 , \8087 , \8122 );
xnor \U$7806 ( \8149 , \8148 , \8089 );
nand \U$7807 ( \8150 , \8147 , \8149 );
nand \U$7808 ( \8151 , \8126 , \8150 );
xor \U$7809 ( \8152 , \5710 , \5760 );
and \U$7810 ( \8153 , \8152 , \5765 );
and \U$7811 ( \8154 , \5710 , \5760 );
or \U$7812 ( \8155 , \8153 , \8154 );
xor \U$7813 ( \8156 , \5627 , \5705 );
and \U$7814 ( \8157 , \8156 , \5766 );
and \U$7815 ( \8158 , \5627 , \5705 );
or \U$7816 ( \8159 , \8157 , \8158 );
xor \U$7817 ( \8160 , \8155 , \8159 );
xor \U$7818 ( \8161 , \8132 , \8134 );
xor \U$7819 ( \8162 , \8161 , \8137 );
and \U$7820 ( \8163 , \8160 , \8162 );
and \U$7821 ( \8164 , \8155 , \8159 );
or \U$7822 ( \8165 , \8163 , \8164 );
xor \U$7823 ( \8166 , \8128 , \8140 );
xor \U$7824 ( \8167 , \8166 , \8143 );
nor \U$7825 ( \8168 , \8165 , \8167 );
not \U$7826 ( \8169 , \8168 );
xor \U$7827 ( \8170 , \8155 , \8159 );
xor \U$7828 ( \8171 , \8170 , \8162 );
xor \U$7829 ( \8172 , \5447 , \5767 );
and \U$7830 ( \8173 , \8172 , \5787 );
and \U$7831 ( \8174 , \5447 , \5767 );
or \U$7832 ( \8175 , \8173 , \8174 );
or \U$7833 ( \8176 , \8171 , \8175 );
nand \U$7834 ( \8177 , \8169 , \8176 );
nor \U$7835 ( \8178 , \8151 , \8177 );
xor \U$7836 ( \8179 , \2118 , \2126 );
xor \U$7837 ( \8180 , \8179 , \2135 );
xor \U$7838 ( \8181 , \7610 , \7619 );
and \U$7839 ( \8182 , \8181 , \7626 );
and \U$7840 ( \8183 , \7610 , \7619 );
or \U$7841 ( \8184 , \8182 , \8183 );
xor \U$7842 ( \8185 , \8180 , \8184 );
xor \U$7843 ( \8186 , \7591 , \2259 );
and \U$7844 ( \8187 , \8186 , \7597 );
and \U$7845 ( \8188 , \7591 , \2259 );
or \U$7846 ( \8189 , \8187 , \8188 );
xor \U$7847 ( \8190 , \8185 , \8189 );
xor \U$7848 ( \8191 , \2268 , \2277 );
xor \U$7849 ( \8192 , \8191 , \2287 );
and \U$7850 ( \8193 , \7627 , \8192 );
xor \U$7851 ( \8194 , \2268 , \2277 );
xor \U$7852 ( \8195 , \8194 , \2287 );
and \U$7853 ( \8196 , \7687 , \8195 );
and \U$7854 ( \8197 , \7627 , \7687 );
or \U$7855 ( \8198 , \8193 , \8196 , \8197 );
xor \U$7856 ( \8199 , \8190 , \8198 );
xor \U$7857 ( \8200 , \2296 , \2298 );
xor \U$7858 ( \8201 , \8200 , \2301 );
and \U$7859 ( \8202 , \8199 , \8201 );
and \U$7860 ( \8203 , \8190 , \8198 );
or \U$7861 ( \8204 , \8202 , \8203 );
xor \U$7862 ( \8205 , \8029 , \8033 );
and \U$7863 ( \8206 , \8205 , \8038 );
and \U$7864 ( \8207 , \8029 , \8033 );
or \U$7865 ( \8208 , \8206 , \8207 );
xor \U$7866 ( \8209 , \7582 , \7584 );
and \U$7867 ( \8210 , \8209 , \7598 );
and \U$7868 ( \8211 , \7582 , \7584 );
or \U$7869 ( \8212 , \8210 , \8211 );
xor \U$7870 ( \8213 , \8208 , \8212 );
xor \U$7871 ( \8214 , \2248 , \2260 );
xor \U$7872 ( \8215 , \8214 , \2290 );
and \U$7873 ( \8216 , \8213 , \8215 );
and \U$7874 ( \8217 , \8208 , \8212 );
or \U$7875 ( \8218 , \8216 , \8217 );
xor \U$7876 ( \8219 , \2201 , \2293 );
xor \U$7877 ( \8220 , \8219 , \2304 );
xor \U$7878 ( \8221 , \8218 , \8220 );
xor \U$7879 ( \8222 , \8180 , \8184 );
and \U$7880 ( \8223 , \8222 , \8189 );
and \U$7881 ( \8224 , \8180 , \8184 );
or \U$7882 ( \8225 , \8223 , \8224 );
xor \U$7883 ( \8226 , \2099 , \2138 );
xor \U$7884 ( \8227 , \8226 , \2163 );
xor \U$7885 ( \8228 , \8225 , \8227 );
xor \U$7886 ( \8229 , \2172 , \2174 );
xor \U$7887 ( \8230 , \8229 , \2177 );
xor \U$7888 ( \8231 , \8228 , \8230 );
xor \U$7889 ( \8232 , \8221 , \8231 );
xor \U$7890 ( \8233 , \8204 , \8232 );
xor \U$7891 ( \8234 , \8208 , \8212 );
xor \U$7892 ( \8235 , \8234 , \8215 );
xor \U$7893 ( \8236 , \7987 , \8024 );
and \U$7894 ( \8237 , \8236 , \8039 );
and \U$7895 ( \8238 , \7987 , \8024 );
or \U$7896 ( \8239 , \8237 , \8238 );
xor \U$7897 ( \8240 , \8235 , \8239 );
xor \U$7898 ( \8241 , \8190 , \8198 );
xor \U$7899 ( \8242 , \8241 , \8201 );
and \U$7900 ( \8243 , \8240 , \8242 );
and \U$7901 ( \8244 , \8235 , \8239 );
or \U$7902 ( \8245 , \8243 , \8244 );
xor \U$7903 ( \8246 , \8233 , \8245 );
xor \U$7904 ( \8247 , \7599 , \7689 );
and \U$7905 ( \8248 , \8247 , \7779 );
and \U$7906 ( \8249 , \7599 , \7689 );
or \U$7907 ( \8250 , \8248 , \8249 );
xor \U$7908 ( \8251 , \8235 , \8239 );
xor \U$7909 ( \8252 , \8251 , \8242 );
xor \U$7910 ( \8253 , \8250 , \8252 );
xor \U$7911 ( \8254 , \8040 , \8044 );
and \U$7912 ( \8255 , \8254 , \8083 );
and \U$7913 ( \8256 , \8040 , \8044 );
or \U$7914 ( \8257 , \8255 , \8256 );
and \U$7915 ( \8258 , \8253 , \8257 );
and \U$7916 ( \8259 , \8250 , \8252 );
or \U$7917 ( \8260 , \8258 , \8259 );
nor \U$7918 ( \8261 , \8246 , \8260 );
not \U$7919 ( \8262 , \8261 );
xor \U$7920 ( \8263 , \7780 , \7982 );
and \U$7921 ( \8264 , \8263 , \8084 );
and \U$7922 ( \8265 , \7780 , \7982 );
or \U$7923 ( \8266 , \8264 , \8265 );
not \U$7924 ( \8267 , \8266 );
xor \U$7925 ( \8268 , \8250 , \8252 );
xor \U$7926 ( \8269 , \8268 , \8257 );
not \U$7927 ( \8270 , \8269 );
nand \U$7928 ( \8271 , \8267 , \8270 );
nand \U$7929 ( \8272 , \8262 , \8271 );
xor \U$7930 ( \8273 , \8225 , \8227 );
and \U$7931 ( \8274 , \8273 , \8230 );
and \U$7932 ( \8275 , \8225 , \8227 );
or \U$7933 ( \8276 , \8274 , \8275 );
xor \U$7934 ( \8277 , \2199 , \2307 );
xor \U$7935 ( \8278 , \8277 , \2310 );
xor \U$7936 ( \8279 , \8276 , \8278 );
xor \U$7937 ( \8280 , \8218 , \8220 );
and \U$7938 ( \8281 , \8280 , \8231 );
and \U$7939 ( \8282 , \8218 , \8220 );
or \U$7940 ( \8283 , \8281 , \8282 );
xor \U$7941 ( \8284 , \8279 , \8283 );
xor \U$7942 ( \8285 , \8204 , \8232 );
and \U$7943 ( \8286 , \8285 , \8245 );
and \U$7944 ( \8287 , \8204 , \8232 );
or \U$7945 ( \8288 , \8286 , \8287 );
nor \U$7946 ( \8289 , \8284 , \8288 );
nor \U$7947 ( \8290 , \8272 , \8289 );
nand \U$7948 ( \8291 , \8178 , \8290 );
xor \U$7949 ( \8292 , \8276 , \8278 );
and \U$7950 ( \8293 , \8292 , \8283 );
and \U$7951 ( \8294 , \8276 , \8278 );
or \U$7952 ( \8295 , \8293 , \8294 );
xor \U$7953 ( \8296 , \2194 , \2196 );
xor \U$7954 ( \8297 , \8296 , \2313 );
nor \U$7955 ( \8298 , \8295 , \8297 );
nor \U$7956 ( \8299 , \8291 , \8298 );
and \U$7957 ( \8300 , \7547 , \8299 );
not \U$7958 ( \8301 , \8300 );
xor \U$7959 ( \8302 , \7040 , \7043 );
xor \U$7960 ( \8303 , \8302 , \7046 );
xor \U$7961 ( \8304 , \7267 , \7372 );
xor \U$7962 ( \8305 , \8304 , \7483 );
xor \U$7963 ( \8306 , \8303 , \8305 );
not \U$7964 ( \8307 , \4354 );
not \U$7965 ( \8308 , \5941 );
or \U$7966 ( \8309 , \8307 , \8308 );
not \U$7967 ( \8310 , \4370 );
nand \U$7968 ( \8311 , \8309 , \8310 );
nand \U$7969 ( \8312 , \7283 , \613 );
not \U$7970 ( \8313 , \8312 );
and \U$7971 ( \8314 , \8311 , \8313 );
not \U$7972 ( \8315 , \8311 );
and \U$7973 ( \8316 , \8315 , \8312 );
nor \U$7974 ( \8317 , \8314 , \8316 );
buf \U$7975 ( \8318 , \8317 );
not \U$7976 ( \8319 , \8318 );
buf \U$7977 ( \8320 , \8319 );
not \U$7978 ( \8321 , \8320 );
and \U$7979 ( \8322 , \1393 , \8321 );
not \U$7980 ( \8323 , \1376 );
xor \U$7981 ( \8324 , \1313 , \6939 );
not \U$7982 ( \8325 , \8324 );
or \U$7983 ( \8326 , \8323 , \8325 );
xor \U$7984 ( \8327 , \1313 , \7300 );
nand \U$7985 ( \8328 , \8327 , \1429 );
nand \U$7986 ( \8329 , \8326 , \8328 );
xor \U$7987 ( \8330 , \8322 , \8329 );
not \U$7988 ( \8331 , \1294 );
not \U$7989 ( \8332 , \7310 );
or \U$7990 ( \8333 , \8331 , \8332 );
not \U$7991 ( \8334 , \1288 );
not \U$7992 ( \8335 , \6943 );
or \U$7993 ( \8336 , \8334 , \8335 );
not \U$7994 ( \8337 , \6602 );
buf \U$7995 ( \8338 , \8337 );
not \U$7996 ( \8339 , \8338 );
nand \U$7997 ( \8340 , \8339 , \1245 );
nand \U$7998 ( \8341 , \8336 , \8340 );
nand \U$7999 ( \8342 , \8341 , \1265 );
nand \U$8000 ( \8343 , \8333 , \8342 );
and \U$8001 ( \8344 , \8330 , \8343 );
and \U$8002 ( \8345 , \8322 , \8329 );
or \U$8003 ( \8346 , \8344 , \8345 );
not \U$8004 ( \8347 , RIbb2e260_43);
and \U$8005 ( \8348 , \8347 , RIbb2e2d8_42);
not \U$8006 ( \8349 , RIbb2e2d8_42);
and \U$8007 ( \8350 , RIbb2e260_43, \8349 );
nor \U$8008 ( \8351 , \8348 , \8350 );
buf \U$8009 ( \8352 , \8351 );
not \U$8010 ( \8353 , \8352 );
buf \U$8011 ( \8354 , \8353 );
not \U$8012 ( \8355 , \8354 );
not \U$8013 ( \8356 , \8355 );
not \U$8014 ( \8357 , RIbb2e350_41);
and \U$8015 ( \8358 , \8357 , \8349 );
and \U$8016 ( \8359 , RIbb2e350_41, RIbb2e2d8_42);
nor \U$8017 ( \8360 , \8358 , \8359 );
and \U$8018 ( \8361 , \8360 , \8351 );
buf \U$8019 ( \8362 , \8361 );
not \U$8020 ( \8363 , \8362 );
not \U$8021 ( \8364 , \8363 );
or \U$8022 ( \8365 , \8356 , \8364 );
nand \U$8023 ( \8366 , \8365 , RIbb2e350_41);
not \U$8024 ( \8367 , \8366 );
not \U$8025 ( \8368 , \1737 );
not \U$8026 ( \8369 , \7453 );
or \U$8027 ( \8370 , \8368 , \8369 );
not \U$8028 ( \8371 , \1703 );
not \U$8029 ( \8372 , RIbb2f340_7);
not \U$8030 ( \8373 , \4393 );
or \U$8031 ( \8374 , \8372 , \8373 );
buf \U$8032 ( \8375 , \4390 );
nand \U$8033 ( \8376 , \8375 , \2700 );
nand \U$8034 ( \8377 , \8374 , \8376 );
nand \U$8035 ( \8378 , \8371 , \8377 );
nand \U$8036 ( \8379 , \8370 , \8378 );
not \U$8037 ( \8380 , \8379 );
or \U$8038 ( \8381 , \8367 , \8380 );
or \U$8039 ( \8382 , \8379 , \8366 );
not \U$8040 ( \8383 , \1147 );
not \U$8041 ( \8384 , \7321 );
or \U$8042 ( \8385 , \8383 , \8384 );
not \U$8043 ( \8386 , RIbb2f430_5);
buf \U$8044 ( \8387 , \6229 );
not \U$8045 ( \8388 , \8387 );
not \U$8046 ( \8389 , \8388 );
or \U$8047 ( \8390 , \8386 , \8389 );
nand \U$8048 ( \8391 , \7111 , \1085 );
nand \U$8049 ( \8392 , \8390 , \8391 );
nand \U$8050 ( \8393 , \8392 , \1090 );
nand \U$8051 ( \8394 , \8385 , \8393 );
nand \U$8052 ( \8395 , \8382 , \8394 );
nand \U$8053 ( \8396 , \8381 , \8395 );
xor \U$8054 ( \8397 , \8346 , \8396 );
xor \U$8055 ( \8398 , \7301 , \7312 );
xor \U$8056 ( \8399 , \8398 , \7323 );
and \U$8057 ( \8400 , \8397 , \8399 );
and \U$8058 ( \8401 , \8346 , \8396 );
or \U$8059 ( \8402 , \8400 , \8401 );
xor \U$8060 ( \8403 , \7278 , \7326 );
xor \U$8061 ( \8404 , \8403 , \7369 );
xor \U$8062 ( \8405 , \8402 , \8404 );
not \U$8063 ( \8406 , \4791 );
not \U$8064 ( \8407 , \7392 );
or \U$8065 ( \8408 , \8406 , \8407 );
not \U$8066 ( \8409 , RIbb2e710_33);
not \U$8067 ( \8410 , \4595 );
or \U$8068 ( \8411 , \8409 , \8410 );
nand \U$8069 ( \8412 , \1038 , \2935 );
nand \U$8070 ( \8413 , \8411 , \8412 );
nand \U$8071 ( \8414 , \8413 , \3887 );
nand \U$8072 ( \8415 , \8408 , \8414 );
not \U$8073 ( \8416 , \8415 );
not \U$8074 ( \8417 , \8416 );
not \U$8075 ( \8418 , \2078 );
not \U$8076 ( \8419 , \7401 );
or \U$8077 ( \8420 , \8418 , \8419 );
not \U$8078 ( \8421 , RIbb2ecb0_21);
not \U$8079 ( \8422 , \1853 );
or \U$8080 ( \8423 , \8421 , \8422 );
nand \U$8081 ( \8424 , \1852 , \2249 );
nand \U$8082 ( \8425 , \8423 , \8424 );
nand \U$8083 ( \8426 , \8425 , \2077 );
nand \U$8084 ( \8427 , \8420 , \8426 );
not \U$8085 ( \8428 , \8427 );
not \U$8086 ( \8429 , \8428 );
or \U$8087 ( \8430 , \8417 , \8429 );
not \U$8088 ( \8431 , \3383 );
not \U$8089 ( \8432 , \7461 );
or \U$8090 ( \8433 , \8431 , \8432 );
not \U$8091 ( \8434 , RIbb2ebc0_23);
not \U$8092 ( \8435 , \3822 );
or \U$8093 ( \8436 , \8434 , \8435 );
nand \U$8094 ( \8437 , \3821 , \3388 );
nand \U$8095 ( \8438 , \8436 , \8437 );
nand \U$8096 ( \8439 , \8438 , \3406 );
nand \U$8097 ( \8440 , \8433 , \8439 );
nand \U$8098 ( \8441 , \8430 , \8440 );
nand \U$8099 ( \8442 , \8427 , \8415 );
nand \U$8100 ( \8443 , \8441 , \8442 );
not \U$8101 ( \8444 , \7102 );
not \U$8102 ( \8445 , \8444 );
not \U$8103 ( \8446 , \8445 );
xnor \U$8104 ( \8447 , RIbb2e440_39, \894 );
not \U$8105 ( \8448 , \8447 );
or \U$8106 ( \8449 , \8446 , \8448 );
buf \U$8107 ( \8450 , \7104 );
nand \U$8108 ( \8451 , \7274 , \8450 );
nand \U$8109 ( \8452 , \8449 , \8451 );
not \U$8110 ( \8453 , \5845 );
not \U$8111 ( \8454 , \7347 );
or \U$8112 ( \8455 , \8453 , \8454 );
not \U$8113 ( \8456 , RIbb2e620_35);
not \U$8114 ( \8457 , \3981 );
or \U$8115 ( \8458 , \8456 , \8457 );
nand \U$8116 ( \8459 , \952 , \5840 );
nand \U$8117 ( \8460 , \8458 , \8459 );
nand \U$8118 ( \8461 , \8460 , \4712 );
nand \U$8119 ( \8462 , \8455 , \8461 );
xor \U$8120 ( \8463 , \8452 , \8462 );
not \U$8121 ( \8464 , \2963 );
and \U$8122 ( \8465 , RIbb2ead0_25, \5407 );
not \U$8123 ( \8466 , RIbb2ead0_25);
and \U$8124 ( \8467 , \8466 , \3291 );
or \U$8125 ( \8468 , \8465 , \8467 );
not \U$8126 ( \8469 , \8468 );
or \U$8127 ( \8470 , \8464 , \8469 );
and \U$8128 ( \8471 , RIbb2ead0_25, \1170 );
not \U$8129 ( \8472 , RIbb2ead0_25);
and \U$8130 ( \8473 , \8472 , \3736 );
or \U$8131 ( \8474 , \8471 , \8473 );
nand \U$8132 ( \8475 , \8474 , \2980 );
nand \U$8133 ( \8476 , \8470 , \8475 );
and \U$8134 ( \8477 , \8463 , \8476 );
and \U$8135 ( \8478 , \8452 , \8462 );
or \U$8136 ( \8479 , \8477 , \8478 );
xor \U$8137 ( \8480 , \8443 , \8479 );
not \U$8138 ( \8481 , \1011 );
not \U$8139 ( \8482 , RIbb2f160_11);
not \U$8140 ( \8483 , \3044 );
not \U$8141 ( \8484 , \8483 );
or \U$8142 ( \8485 , \8482 , \8484 );
nand \U$8143 ( \8486 , \3046 , \1043 );
nand \U$8144 ( \8487 , \8485 , \8486 );
not \U$8145 ( \8488 , \8487 );
or \U$8146 ( \8489 , \8481 , \8488 );
not \U$8147 ( \8490 , RIbb2f160_11);
buf \U$8148 ( \8491 , \4020 );
not \U$8149 ( \8492 , \8491 );
not \U$8150 ( \8493 , \8492 );
or \U$8151 ( \8494 , \8490 , \8493 );
nand \U$8152 ( \8495 , \3022 , \1048 );
nand \U$8153 ( \8496 , \8494 , \8495 );
nand \U$8154 ( \8497 , \8496 , \1077 );
nand \U$8155 ( \8498 , \8489 , \8497 );
not \U$8156 ( \8499 , \3445 );
not \U$8157 ( \8500 , RIbb2e9e0_27);
not \U$8158 ( \8501 , \4006 );
not \U$8159 ( \8502 , \8501 );
or \U$8160 ( \8503 , \8500 , \8502 );
nand \U$8161 ( \8504 , \4006 , \3454 );
nand \U$8162 ( \8505 , \8503 , \8504 );
not \U$8163 ( \8506 , \8505 );
or \U$8164 ( \8507 , \8499 , \8506 );
nand \U$8165 ( \8508 , \7429 , \3465 );
nand \U$8166 ( \8509 , \8507 , \8508 );
xor \U$8167 ( \8510 , \8498 , \8509 );
not \U$8168 ( \8511 , \1533 );
not \U$8169 ( \8512 , RIbb2f250_9);
not \U$8170 ( \8513 , \4749 );
or \U$8171 ( \8514 , \8512 , \8513 );
nand \U$8172 ( \8515 , \3092 , \1566 );
nand \U$8173 ( \8516 , \8514 , \8515 );
not \U$8174 ( \8517 , \8516 );
or \U$8175 ( \8518 , \8511 , \8517 );
not \U$8176 ( \8519 , RIbb2f250_9);
not \U$8177 ( \8520 , \3276 );
or \U$8178 ( \8521 , \8519 , \8520 );
nand \U$8179 ( \8522 , \3003 , \1566 );
nand \U$8180 ( \8523 , \8521 , \8522 );
nand \U$8181 ( \8524 , \8523 , \1570 );
nand \U$8182 ( \8525 , \8518 , \8524 );
and \U$8183 ( \8526 , \8510 , \8525 );
and \U$8184 ( \8527 , \8498 , \8509 );
or \U$8185 ( \8528 , \8526 , \8527 );
and \U$8186 ( \8529 , \8480 , \8528 );
and \U$8187 ( \8530 , \8443 , \8479 );
or \U$8188 ( \8531 , \8529 , \8530 );
and \U$8189 ( \8532 , \8405 , \8531 );
and \U$8190 ( \8533 , \8402 , \8404 );
or \U$8191 ( \8534 , \8532 , \8533 );
xor \U$8192 ( \8535 , \8306 , \8534 );
not \U$8193 ( \8536 , \7278 );
not \U$8194 ( \8537 , \1011 );
not \U$8195 ( \8538 , \8496 );
or \U$8196 ( \8539 , \8537 , \8538 );
nand \U$8197 ( \8540 , \7023 , \1077 );
nand \U$8198 ( \8541 , \8539 , \8540 );
xor \U$8199 ( \8542 , \8536 , \8541 );
not \U$8200 ( \8543 , \998 );
not \U$8201 ( \8544 , \7011 );
or \U$8202 ( \8545 , \8543 , \8544 );
not \U$8203 ( \8546 , RIbb2f070_13);
not \U$8204 ( \8547 , \3226 );
or \U$8205 ( \8548 , \8546 , \8547 );
nand \U$8206 ( \8549 , \3228 , \1656 );
nand \U$8207 ( \8550 , \8548 , \8549 );
nand \U$8208 ( \8551 , \8550 , \916 );
nand \U$8209 ( \8552 , \8545 , \8551 );
and \U$8210 ( \8553 , \8542 , \8552 );
and \U$8211 ( \8554 , \8536 , \8541 );
or \U$8212 ( \8555 , \8553 , \8554 );
xor \U$8213 ( \8556 , \6976 , \6985 );
xor \U$8214 ( \8557 , \8556 , \6996 );
xor \U$8215 ( \8558 , \8555 , \8557 );
xor \U$8216 ( \8559 , \7227 , \7249 );
xor \U$8217 ( \8560 , \8559 , \7237 );
and \U$8218 ( \8561 , \8558 , \8560 );
and \U$8219 ( \8562 , \8555 , \8557 );
or \U$8220 ( \8563 , \8561 , \8562 );
xor \U$8221 ( \8564 , \7106 , \7117 );
xor \U$8222 ( \8565 , \8564 , \7128 );
nand \U$8223 ( \8566 , \1376 , \6947 );
nand \U$8224 ( \8567 , \8324 , \1430 );
nand \U$8225 ( \8568 , \8566 , \8567 );
not \U$8226 ( \8569 , \1570 );
not \U$8227 ( \8570 , \7233 );
or \U$8228 ( \8571 , \8569 , \8570 );
nand \U$8229 ( \8572 , \8523 , \1533 );
nand \U$8230 ( \8573 , \8571 , \8572 );
xor \U$8231 ( \8574 , \8568 , \8573 );
not \U$8232 ( \8575 , \2963 );
not \U$8233 ( \8576 , \6959 );
or \U$8234 ( \8577 , \8575 , \8576 );
nand \U$8235 ( \8578 , \8468 , \2980 );
nand \U$8236 ( \8579 , \8577 , \8578 );
and \U$8237 ( \8580 , \8574 , \8579 );
and \U$8238 ( \8581 , \8568 , \8573 );
or \U$8239 ( \8582 , \8580 , \8581 );
xor \U$8240 ( \8583 , \8565 , \8582 );
xor \U$8241 ( \8584 , \6940 , \6951 );
xor \U$8242 ( \8585 , \8584 , \6961 );
and \U$8243 ( \8586 , \8583 , \8585 );
and \U$8244 ( \8587 , \8565 , \8582 );
or \U$8245 ( \8588 , \8586 , \8587 );
xnor \U$8246 ( \8589 , \8563 , \8588 );
xor \U$8247 ( \8590 , \7162 , \7175 );
xor \U$8248 ( \8591 , \8590 , \7151 );
xor \U$8249 ( \8592 , \7199 , \7188 );
xor \U$8250 ( \8593 , \8592 , \7212 );
xor \U$8251 ( \8594 , \8591 , \8593 );
xor \U$8252 ( \8595 , \7025 , \7013 );
xor \U$8253 ( \8596 , \7037 , \8595 );
and \U$8254 ( \8597 , \8594 , \8596 );
and \U$8255 ( \8598 , \8591 , \8593 );
or \U$8256 ( \8599 , \8597 , \8598 );
buf \U$8257 ( \8600 , \8599 );
xnor \U$8258 ( \8601 , \8589 , \8600 );
xor \U$8259 ( \8602 , \8535 , \8601 );
xor \U$8260 ( \8603 , \8591 , \8593 );
xor \U$8261 ( \8604 , \8603 , \8596 );
xor \U$8262 ( \8605 , \8322 , \8329 );
xor \U$8263 ( \8606 , \8605 , \8343 );
not \U$8264 ( \8607 , \8606 );
buf \U$8265 ( \8608 , \597 );
not \U$8266 ( \8609 , \602 );
nand \U$8267 ( \8610 , \8609 , \606 );
nor \U$8268 ( \8611 , \8608 , \8610 );
not \U$8269 ( \8612 , \8611 );
not \U$8270 ( \8613 , \4361 );
or \U$8271 ( \8614 , \8612 , \8613 );
not \U$8272 ( \8615 , \4364 );
not \U$8273 ( \8616 , \8610 );
and \U$8274 ( \8617 , \8615 , \8616 );
not \U$8275 ( \8618 , \606 );
not \U$8276 ( \8619 , \653 );
or \U$8277 ( \8620 , \8618 , \8619 );
nand \U$8278 ( \8621 , \8620 , \657 );
nor \U$8279 ( \8622 , \8617 , \8621 );
nand \U$8280 ( \8623 , \8614 , \8622 );
nor \U$8281 ( \8624 , \660 , \503 );
and \U$8282 ( \8625 , \8623 , \8624 );
not \U$8283 ( \8626 , \8623 );
not \U$8284 ( \8627 , \8624 );
and \U$8285 ( \8628 , \8626 , \8627 );
nor \U$8286 ( \8629 , \8625 , \8628 );
buf \U$8287 ( \8630 , \8629 );
buf \U$8288 ( \8631 , \8630 );
and \U$8289 ( \8632 , \1313 , \8631 );
not \U$8290 ( \8633 , \1265 );
not \U$8291 ( \8634 , \1246 );
not \U$8292 ( \8635 , \6938 );
or \U$8293 ( \8636 , \8634 , \8635 );
buf \U$8294 ( \8637 , \6936 );
buf \U$8295 ( \8638 , \8637 );
not \U$8296 ( \8639 , \8638 );
not \U$8297 ( \8640 , \8639 );
nand \U$8298 ( \8641 , \8640 , \1289 );
nand \U$8299 ( \8642 , \8636 , \8641 );
not \U$8300 ( \8643 , \8642 );
or \U$8301 ( \8644 , \8633 , \8643 );
nand \U$8302 ( \8645 , \8341 , \1294 );
nand \U$8303 ( \8646 , \8644 , \8645 );
xor \U$8304 ( \8647 , \8632 , \8646 );
not \U$8305 ( \8648 , \3445 );
not \U$8306 ( \8649 , RIbb2e9e0_27);
not \U$8307 ( \8650 , \3290 );
or \U$8308 ( \8651 , \8649 , \8650 );
nand \U$8309 ( \8652 , \1283 , \3454 );
nand \U$8310 ( \8653 , \8651 , \8652 );
not \U$8311 ( \8654 , \8653 );
or \U$8312 ( \8655 , \8648 , \8654 );
nand \U$8313 ( \8656 , \8505 , \3465 );
nand \U$8314 ( \8657 , \8655 , \8656 );
and \U$8315 ( \8658 , \8647 , \8657 );
and \U$8316 ( \8659 , \8632 , \8646 );
or \U$8317 ( \8660 , \8658 , \8659 );
not \U$8318 ( \8661 , \8660 );
xor \U$8319 ( \8662 , \8366 , \8379 );
xnor \U$8320 ( \8663 , \8662 , \8394 );
nand \U$8321 ( \8664 , \8661 , \8663 );
not \U$8322 ( \8665 , \8664 );
or \U$8323 ( \8666 , \8607 , \8665 );
not \U$8324 ( \8667 , \8663 );
nand \U$8325 ( \8668 , \8667 , \8660 );
nand \U$8326 ( \8669 , \8666 , \8668 );
xor \U$8327 ( \8670 , \8346 , \8396 );
xor \U$8328 ( \8671 , \8670 , \8399 );
xor \U$8329 ( \8672 , \8669 , \8671 );
not \U$8330 ( \8673 , \4791 );
not \U$8331 ( \8674 , \8413 );
or \U$8332 ( \8675 , \8673 , \8674 );
not \U$8333 ( \8676 , RIbb2e710_33);
not \U$8334 ( \8677 , \5003 );
or \U$8335 ( \8678 , \8676 , \8677 );
nand \U$8336 ( \8679 , \1548 , \3877 );
nand \U$8337 ( \8680 , \8678 , \8679 );
nand \U$8338 ( \8681 , \8680 , \3887 );
nand \U$8339 ( \8682 , \8675 , \8681 );
not \U$8340 ( \8683 , \8682 );
not \U$8341 ( \8684 , \2077 );
not \U$8342 ( \8685 , RIbb2ecb0_21);
not \U$8343 ( \8686 , \5550 );
or \U$8344 ( \8687 , \8685 , \8686 );
nand \U$8345 ( \8688 , \3564 , \2249 );
nand \U$8346 ( \8689 , \8687 , \8688 );
not \U$8347 ( \8690 , \8689 );
or \U$8348 ( \8691 , \8684 , \8690 );
nand \U$8349 ( \8692 , \8425 , \2078 );
nand \U$8350 ( \8693 , \8691 , \8692 );
not \U$8351 ( \8694 , \8693 );
or \U$8352 ( \8695 , \8683 , \8694 );
or \U$8353 ( \8696 , \8693 , \8682 );
not \U$8354 ( \8697 , \6242 );
not \U$8355 ( \8698 , RIbb2e530_37);
not \U$8356 ( \8699 , \1475 );
or \U$8357 ( \8700 , \8698 , \8699 );
not \U$8358 ( \8701 , RIbb2e530_37);
nand \U$8359 ( \8702 , \4558 , \8701 );
nand \U$8360 ( \8703 , \8700 , \8702 );
not \U$8361 ( \8704 , \8703 );
or \U$8362 ( \8705 , \8697 , \8704 );
not \U$8363 ( \8706 , RIbb2e530_37);
not \U$8364 ( \8707 , \988 );
or \U$8365 ( \8708 , \8706 , \8707 );
nand \U$8366 ( \8709 , \7345 , \7243 );
nand \U$8367 ( \8710 , \8708 , \8709 );
nand \U$8368 ( \8711 , \8710 , \6251 );
nand \U$8369 ( \8712 , \8705 , \8711 );
nand \U$8370 ( \8713 , \8696 , \8712 );
nand \U$8371 ( \8714 , \8695 , \8713 );
not \U$8372 ( \8715 , \5845 );
not \U$8373 ( \8716 , \8460 );
or \U$8374 ( \8717 , \8715 , \8716 );
not \U$8375 ( \8718 , RIbb2e620_35);
not \U$8376 ( \8719 , \1070 );
or \U$8377 ( \8720 , \8718 , \8719 );
nand \U$8378 ( \8721 , \3099 , \6002 );
nand \U$8379 ( \8722 , \8720 , \8721 );
nand \U$8380 ( \8723 , \8722 , \4712 );
nand \U$8381 ( \8724 , \8717 , \8723 );
not \U$8382 ( \8725 , \3383 );
not \U$8383 ( \8726 , \8438 );
or \U$8384 ( \8727 , \8725 , \8726 );
not \U$8385 ( \8728 , RIbb2ebc0_23);
not \U$8386 ( \8729 , \3575 );
or \U$8387 ( \8730 , \8728 , \8729 );
nand \U$8388 ( \8731 , \1339 , \3388 );
nand \U$8389 ( \8732 , \8730 , \8731 );
nand \U$8390 ( \8733 , \3407 , \8732 );
nand \U$8391 ( \8734 , \8727 , \8733 );
xor \U$8392 ( \8735 , \8724 , \8734 );
not \U$8393 ( \8736 , \2963 );
not \U$8394 ( \8737 , \8474 );
or \U$8395 ( \8738 , \8736 , \8737 );
and \U$8396 ( \8739 , RIbb2ead0_25, \3116 );
not \U$8397 ( \8740 , RIbb2ead0_25);
and \U$8398 ( \8741 , \8740 , \4340 );
or \U$8399 ( \8742 , \8739 , \8741 );
nand \U$8400 ( \8743 , \8742 , \2980 );
nand \U$8401 ( \8744 , \8738 , \8743 );
and \U$8402 ( \8745 , \8735 , \8744 );
and \U$8403 ( \8746 , \8724 , \8734 );
or \U$8404 ( \8747 , \8745 , \8746 );
xor \U$8405 ( \8748 , \8714 , \8747 );
not \U$8406 ( \8749 , \8450 );
not \U$8407 ( \8750 , \8447 );
or \U$8408 ( \8751 , \8749 , \8750 );
and \U$8409 ( \8752 , RIbb2e440_39, \3262 );
not \U$8410 ( \8753 , RIbb2e440_39);
not \U$8411 ( \8754 , \1508 );
not \U$8412 ( \8755 , \8754 );
and \U$8413 ( \8756 , \8753 , \8755 );
or \U$8414 ( \8757 , \8752 , \8756 );
nand \U$8415 ( \8758 , \8757 , \8445 );
nand \U$8416 ( \8759 , \8751 , \8758 );
not \U$8417 ( \8760 , \1570 );
not \U$8418 ( \8761 , \8516 );
or \U$8419 ( \8762 , \8760 , \8761 );
not \U$8420 ( \8763 , RIbb2f250_9);
not \U$8421 ( \8764 , \4088 );
or \U$8422 ( \8765 , \8763 , \8764 );
nand \U$8423 ( \8766 , \4089 , \1566 );
nand \U$8424 ( \8767 , \8765 , \8766 );
nand \U$8425 ( \8768 , \8767 , \1533 );
nand \U$8426 ( \8769 , \8762 , \8768 );
xor \U$8427 ( \8770 , \8759 , \8769 );
not \U$8428 ( \8771 , \1077 );
not \U$8429 ( \8772 , \8487 );
or \U$8430 ( \8773 , \8771 , \8772 );
not \U$8431 ( \8774 , RIbb2f160_11);
not \U$8432 ( \8775 , \4411 );
or \U$8433 ( \8776 , \8774 , \8775 );
nand \U$8434 ( \8777 , \3275 , \1805 );
nand \U$8435 ( \8778 , \8776 , \8777 );
nand \U$8436 ( \8779 , \8778 , \1011 );
nand \U$8437 ( \8780 , \8773 , \8779 );
and \U$8438 ( \8781 , \8770 , \8780 );
and \U$8439 ( \8782 , \8759 , \8769 );
or \U$8440 ( \8783 , \8781 , \8782 );
and \U$8441 ( \8784 , \8748 , \8783 );
and \U$8442 ( \8785 , \8714 , \8747 );
or \U$8443 ( \8786 , \8784 , \8785 );
and \U$8444 ( \8787 , \8672 , \8786 );
and \U$8445 ( \8788 , \8669 , \8671 );
or \U$8446 ( \8789 , \8787 , \8788 );
xor \U$8447 ( \8790 , \8604 , \8789 );
xor \U$8448 ( \8791 , \8402 , \8404 );
xor \U$8449 ( \8792 , \8791 , \8531 );
and \U$8450 ( \8793 , \8790 , \8792 );
and \U$8451 ( \8794 , \8604 , \8789 );
or \U$8452 ( \8795 , \8793 , \8794 );
xor \U$8453 ( \8796 , \8602 , \8795 );
xor \U$8454 ( \8797 , \8498 , \8509 );
xor \U$8455 ( \8798 , \8797 , \8525 );
not \U$8456 ( \8799 , \2940 );
not \U$8457 ( \8800 , RIbb2e800_31);
not \U$8458 ( \8801 , \1688 );
or \U$8459 ( \8802 , \8800 , \8801 );
nand \U$8460 ( \8803 , \3371 , \4096 );
nand \U$8461 ( \8804 , \8802 , \8803 );
not \U$8462 ( \8805 , \8804 );
or \U$8463 ( \8806 , \8799 , \8805 );
not \U$8464 ( \8807 , RIbb2e800_31);
not \U$8465 ( \8808 , \3481 );
or \U$8466 ( \8809 , \8807 , \8808 );
not \U$8467 ( \8810 , RIbb2e800_31);
nand \U$8468 ( \8811 , \3480 , \8810 );
nand \U$8469 ( \8812 , \8809 , \8811 );
nand \U$8470 ( \8813 , \8812 , \3613 );
nand \U$8471 ( \8814 , \8806 , \8813 );
not \U$8472 ( \8815 , \8814 );
not \U$8473 ( \8816 , \853 );
not \U$8474 ( \8817 , RIbb2eda0_19);
not \U$8475 ( \8818 , \3517 );
or \U$8476 ( \8819 , \8817 , \8818 );
nand \U$8477 ( \8820 , \3521 , \1776 );
nand \U$8478 ( \8821 , \8819 , \8820 );
not \U$8479 ( \8822 , \8821 );
or \U$8480 ( \8823 , \8816 , \8822 );
not \U$8481 ( \8824 , RIbb2eda0_19);
not \U$8482 ( \8825 , \3319 );
or \U$8483 ( \8826 , \8824 , \8825 );
nand \U$8484 ( \8827 , \2225 , \3251 );
nand \U$8485 ( \8828 , \8826 , \8827 );
nand \U$8486 ( \8829 , \8828 , \855 );
nand \U$8487 ( \8830 , \8823 , \8829 );
not \U$8488 ( \8831 , \8830 );
or \U$8489 ( \8832 , \8815 , \8831 );
or \U$8490 ( \8833 , \8830 , \8814 );
not \U$8491 ( \8834 , \832 );
not \U$8492 ( \8835 , RIbb2ee90_17);
not \U$8493 ( \8836 , \3141 );
or \U$8494 ( \8837 , \8835 , \8836 );
nand \U$8495 ( \8838 , \3146 , \816 );
nand \U$8496 ( \8839 , \8837 , \8838 );
not \U$8497 ( \8840 , \8839 );
or \U$8498 ( \8841 , \8834 , \8840 );
not \U$8499 ( \8842 , RIbb2ee90_17);
not \U$8500 ( \8843 , \3952 );
or \U$8501 ( \8844 , \8842 , \8843 );
nand \U$8502 ( \8845 , \6108 , \859 );
nand \U$8503 ( \8846 , \8844 , \8845 );
nand \U$8504 ( \8847 , \8846 , \836 );
nand \U$8505 ( \8848 , \8841 , \8847 );
nand \U$8506 ( \8849 , \8833 , \8848 );
nand \U$8507 ( \8850 , \8832 , \8849 );
or \U$8508 ( \8851 , \8798 , \8850 );
not \U$8509 ( \8852 , \2925 );
not \U$8510 ( \8853 , RIbb2e8f0_29);
not \U$8511 ( \8854 , \3242 );
or \U$8512 ( \8855 , \8853 , \8854 );
not \U$8513 ( \8856 , \3238 );
nand \U$8514 ( \8857 , \8856 , \3265 );
nand \U$8515 ( \8858 , \8855 , \8857 );
not \U$8516 ( \8859 , \8858 );
or \U$8517 ( \8860 , \8852 , \8859 );
not \U$8518 ( \8861 , RIbb2e8f0_29);
buf \U$8519 ( \8862 , \1135 );
not \U$8520 ( \8863 , \8862 );
or \U$8521 ( \8864 , \8861 , \8863 );
nand \U$8522 ( \8865 , \7427 , \3800 );
nand \U$8523 ( \8866 , \8864 , \8865 );
nand \U$8524 ( \8867 , \2922 , \8866 );
nand \U$8525 ( \8868 , \8860 , \8867 );
not \U$8526 ( \8869 , \8868 );
not \U$8527 ( \8870 , \916 );
not \U$8528 ( \8871 , RIbb2f070_13);
not \U$8529 ( \8872 , \4021 );
or \U$8530 ( \8873 , \8871 , \8872 );
not \U$8531 ( \8874 , \5962 );
nand \U$8532 ( \8875 , \8874 , \3421 );
nand \U$8533 ( \8876 , \8873 , \8875 );
not \U$8534 ( \8877 , \8876 );
or \U$8535 ( \8878 , \8870 , \8877 );
and \U$8536 ( \8879 , RIbb2f070_13, \7018 );
not \U$8537 ( \8880 , RIbb2f070_13);
and \U$8538 ( \8881 , \8880 , \3654 );
or \U$8539 ( \8882 , \8879 , \8881 );
nand \U$8540 ( \8883 , \8882 , \998 );
nand \U$8541 ( \8884 , \8878 , \8883 );
not \U$8542 ( \8885 , \8884 );
or \U$8543 ( \8886 , \8869 , \8885 );
or \U$8544 ( \8887 , \8884 , \8868 );
not \U$8545 ( \8888 , \1445 );
and \U$8546 ( \8889 , RIbb2ef80_15, \3905 );
not \U$8547 ( \8890 , RIbb2ef80_15);
and \U$8548 ( \8891 , \8890 , \3632 );
or \U$8549 ( \8892 , \8889 , \8891 );
not \U$8550 ( \8893 , \8892 );
or \U$8551 ( \8894 , \8888 , \8893 );
not \U$8552 ( \8895 , \1584 );
and \U$8553 ( \8896 , RIbb2ef80_15, \4639 );
not \U$8554 ( \8897 , RIbb2ef80_15);
and \U$8555 ( \8898 , \8897 , \4640 );
or \U$8556 ( \8899 , \8896 , \8898 );
nand \U$8557 ( \8900 , \8895 , \8899 );
nand \U$8558 ( \8901 , \8894 , \8900 );
nand \U$8559 ( \8902 , \8887 , \8901 );
nand \U$8560 ( \8903 , \8886 , \8902 );
nand \U$8561 ( \8904 , \8851 , \8903 );
nand \U$8562 ( \8905 , \8798 , \8850 );
nand \U$8563 ( \8906 , \8904 , \8905 );
xor \U$8564 ( \8907 , \8452 , \8462 );
xor \U$8565 ( \8908 , \8907 , \8476 );
not \U$8566 ( \8909 , \8908 );
not \U$8567 ( \8910 , \3613 );
not \U$8568 ( \8911 , \7381 );
or \U$8569 ( \8912 , \8910 , \8911 );
nand \U$8570 ( \8913 , \8812 , \2940 );
nand \U$8571 ( \8914 , \8912 , \8913 );
not \U$8572 ( \8915 , \855 );
not \U$8573 ( \8916 , \7365 );
or \U$8574 ( \8917 , \8915 , \8916 );
nand \U$8575 ( \8918 , \8828 , \853 );
nand \U$8576 ( \8919 , \8917 , \8918 );
xor \U$8577 ( \8920 , \8914 , \8919 );
not \U$8578 ( \8921 , \6251 );
not \U$8579 ( \8922 , \8703 );
or \U$8580 ( \8923 , \8921 , \8922 );
nand \U$8581 ( \8924 , \7475 , \6242 );
nand \U$8582 ( \8925 , \8923 , \8924 );
xor \U$8583 ( \8926 , \8920 , \8925 );
not \U$8584 ( \8927 , \8926 );
or \U$8585 ( \8928 , \8909 , \8927 );
or \U$8586 ( \8929 , \8926 , \8908 );
and \U$8587 ( \8930 , \8428 , \8416 );
not \U$8588 ( \8931 , \8428 );
and \U$8589 ( \8932 , \8931 , \8415 );
nor \U$8590 ( \8933 , \8930 , \8932 );
not \U$8591 ( \8934 , \8440 );
and \U$8592 ( \8935 , \8933 , \8934 );
not \U$8593 ( \8936 , \8933 );
and \U$8594 ( \8937 , \8936 , \8440 );
nor \U$8595 ( \8938 , \8935 , \8937 );
not \U$8596 ( \8939 , \8938 );
nand \U$8597 ( \8940 , \8929 , \8939 );
nand \U$8598 ( \8941 , \8928 , \8940 );
xor \U$8599 ( \8942 , \8906 , \8941 );
not \U$8600 ( \8943 , \2925 );
not \U$8601 ( \8944 , \7335 );
or \U$8602 ( \8945 , \8943 , \8944 );
nand \U$8603 ( \8946 , \8858 , \2922 );
nand \U$8604 ( \8947 , \8945 , \8946 );
not \U$8605 ( \8948 , \1517 );
not \U$8606 ( \8949 , \7439 );
or \U$8607 ( \8950 , \8948 , \8949 );
nand \U$8608 ( \8951 , \8899 , \1445 );
nand \U$8609 ( \8952 , \8950 , \8951 );
xor \U$8610 ( \8953 , \8947 , \8952 );
not \U$8611 ( \8954 , \836 );
not \U$8612 ( \8955 , \7416 );
or \U$8613 ( \8956 , \8954 , \8955 );
nand \U$8614 ( \8957 , \8846 , \832 );
nand \U$8615 ( \8958 , \8956 , \8957 );
and \U$8616 ( \8959 , \8953 , \8958 );
and \U$8617 ( \8960 , \8947 , \8952 );
or \U$8618 ( \8961 , \8959 , \8960 );
xor \U$8619 ( \8962 , \8914 , \8919 );
and \U$8620 ( \8963 , \8962 , \8925 );
and \U$8621 ( \8964 , \8914 , \8919 );
or \U$8622 ( \8965 , \8963 , \8964 );
xor \U$8623 ( \8966 , \8961 , \8965 );
xor \U$8624 ( \8967 , \8536 , \8541 );
xor \U$8625 ( \8968 , \8967 , \8552 );
xor \U$8626 ( \8969 , \8966 , \8968 );
and \U$8627 ( \8970 , \8942 , \8969 );
and \U$8628 ( \8971 , \8906 , \8941 );
or \U$8629 ( \8972 , \8970 , \8971 );
xor \U$8630 ( \8973 , \8961 , \8965 );
and \U$8631 ( \8974 , \8973 , \8968 );
and \U$8632 ( \8975 , \8961 , \8965 );
or \U$8633 ( \8976 , \8974 , \8975 );
xor \U$8634 ( \8977 , \8565 , \8582 );
xor \U$8635 ( \8978 , \8977 , \8585 );
xor \U$8636 ( \8979 , \8976 , \8978 );
xor \U$8637 ( \8980 , \7408 , \7444 );
xor \U$8638 ( \8981 , \8980 , \7480 );
xor \U$8639 ( \8982 , \8979 , \8981 );
xor \U$8640 ( \8983 , \8972 , \8982 );
xor \U$8641 ( \8984 , \8443 , \8479 );
xor \U$8642 ( \8985 , \8984 , \8528 );
xor \U$8643 ( \8986 , \8947 , \8952 );
xor \U$8644 ( \8987 , \8986 , \8958 );
not \U$8645 ( \8988 , \8362 );
and \U$8646 ( \8989 , \813 , RIbb2e350_41);
not \U$8647 ( \8990 , \813 );
and \U$8648 ( \8991 , \8990 , \7097 );
or \U$8649 ( \8992 , \8989 , \8991 );
not \U$8650 ( \8993 , \8992 );
or \U$8651 ( \8994 , \8988 , \8993 );
buf \U$8652 ( \8995 , \8354 );
nand \U$8653 ( \8996 , \8995 , RIbb2e350_41);
nand \U$8654 ( \8997 , \8994 , \8996 );
not \U$8655 ( \8998 , \998 );
not \U$8656 ( \8999 , \8550 );
or \U$8657 ( \9000 , \8998 , \8999 );
nand \U$8658 ( \9001 , \8882 , \916 );
nand \U$8659 ( \9002 , \9000 , \9001 );
xor \U$8660 ( \9003 , \8997 , \9002 );
not \U$8661 ( \9004 , \1147 );
not \U$8662 ( \9005 , \8392 );
or \U$8663 ( \9006 , \9004 , \9005 );
not \U$8664 ( \9007 , RIbb2f430_5);
not \U$8665 ( \9008 , \5956 );
or \U$8666 ( \9009 , \9007 , \9008 );
not \U$8667 ( \9010 , \7308 );
not \U$8668 ( \9011 , \9010 );
nand \U$8669 ( \9012 , \9011 , \1085 );
nand \U$8670 ( \9013 , \9009 , \9012 );
nand \U$8671 ( \9014 , \9013 , \1090 );
nand \U$8672 ( \9015 , \9006 , \9014 );
not \U$8673 ( \9016 , \1737 );
not \U$8674 ( \9017 , \8377 );
or \U$8675 ( \9018 , \9016 , \9017 );
not \U$8676 ( \9019 , RIbb2f340_7);
buf \U$8677 ( \9020 , \4695 );
not \U$8678 ( \9021 , \9020 );
not \U$8679 ( \9022 , \9021 );
not \U$8680 ( \9023 , \9022 );
not \U$8681 ( \9024 , \9023 );
or \U$8682 ( \9025 , \9019 , \9024 );
nand \U$8683 ( \9026 , \6198 , \1692 );
nand \U$8684 ( \9027 , \9025 , \9026 );
nand \U$8685 ( \9028 , \9027 , \1702 );
nand \U$8686 ( \9029 , \9018 , \9028 );
or \U$8687 ( \9030 , \9015 , \9029 );
not \U$8688 ( \9031 , \1376 );
not \U$8689 ( \9032 , \8327 );
or \U$8690 ( \9033 , \9031 , \9032 );
not \U$8691 ( \9034 , \6207 );
xor \U$8692 ( \9035 , \1393 , \8321 );
nand \U$8693 ( \9036 , \9034 , \9035 );
nand \U$8694 ( \9037 , \9033 , \9036 );
nand \U$8695 ( \9038 , \9030 , \9037 );
nand \U$8696 ( \9039 , \9015 , \9029 );
nand \U$8697 ( \9040 , \9038 , \9039 );
xor \U$8698 ( \9041 , \9003 , \9040 );
xor \U$8699 ( \9042 , \8987 , \9041 );
not \U$8700 ( \9043 , \8997 );
not \U$8701 ( \9044 , \1429 );
xor \U$8702 ( \9045 , \1313 , \8631 );
not \U$8703 ( \9046 , \9045 );
or \U$8704 ( \9047 , \9044 , \9046 );
nand \U$8705 ( \9048 , \9035 , \1376 );
nand \U$8706 ( \9049 , \9047 , \9048 );
not \U$8707 ( \9050 , \9049 );
not \U$8708 ( \9051 , \9050 );
not \U$8709 ( \9052 , \1147 );
not \U$8710 ( \9053 , \9013 );
or \U$8711 ( \9054 , \9052 , \9053 );
not \U$8712 ( \9055 , RIbb2f430_5);
not \U$8713 ( \9056 , \8338 );
not \U$8714 ( \9057 , \9056 );
not \U$8715 ( \9058 , \9057 );
or \U$8716 ( \9059 , \9055 , \9058 );
not \U$8717 ( \9060 , \6943 );
nand \U$8718 ( \9061 , \9060 , \1647 );
nand \U$8719 ( \9062 , \9059 , \9061 );
nand \U$8720 ( \9063 , \9062 , \1090 );
nand \U$8721 ( \9064 , \9054 , \9063 );
not \U$8722 ( \9065 , \9064 );
not \U$8723 ( \9066 , \9065 );
or \U$8724 ( \9067 , \9051 , \9066 );
not \U$8725 ( \9068 , \1265 );
not \U$8726 ( \9069 , \1246 );
not \U$8727 ( \9070 , \7296 );
buf \U$8728 ( \9071 , \9070 );
not \U$8729 ( \9072 , \9071 );
or \U$8730 ( \9073 , \9069 , \9072 );
not \U$8731 ( \9074 , \9071 );
nand \U$8732 ( \9075 , \9074 , \1289 );
nand \U$8733 ( \9076 , \9073 , \9075 );
not \U$8734 ( \9077 , \9076 );
or \U$8735 ( \9078 , \9068 , \9077 );
nand \U$8736 ( \9079 , \8642 , \1294 );
nand \U$8737 ( \9080 , \9078 , \9079 );
not \U$8738 ( \9081 , \9080 );
not \U$8739 ( \9082 , \9081 );
nand \U$8740 ( \9083 , \9067 , \9082 );
nand \U$8741 ( \9084 , \9049 , \9064 );
nand \U$8742 ( \9085 , \9083 , \9084 );
xor \U$8743 ( \9086 , \9043 , \9085 );
and \U$8744 ( \9087 , RIbb2e1e8_44, RIbb2e260_43);
not \U$8745 ( \9088 , RIbb2e1e8_44);
and \U$8746 ( \9089 , \9088 , \8347 );
nor \U$8747 ( \9090 , \9087 , \9089 );
not \U$8748 ( \9091 , \9090 );
and \U$8749 ( \9092 , RIbb2e1e8_44, RIbb2e170_45);
not \U$8750 ( \9093 , RIbb2e1e8_44);
not \U$8751 ( \9094 , RIbb2e170_45);
and \U$8752 ( \9095 , \9093 , \9094 );
nor \U$8753 ( \9096 , \9092 , \9095 );
nor \U$8754 ( \9097 , \9091 , \9096 );
buf \U$8755 ( \9098 , \9097 );
buf \U$8756 ( \9099 , \9096 );
or \U$8757 ( \9100 , \9098 , \9099 );
nand \U$8758 ( \9101 , \9100 , RIbb2e260_43);
not \U$8759 ( \9102 , \1737 );
not \U$8760 ( \9103 , \9027 );
or \U$8761 ( \9104 , \9102 , \9103 );
not \U$8762 ( \9105 , RIbb2f340_7);
not \U$8763 ( \9106 , \8388 );
or \U$8764 ( \9107 , \9105 , \9106 );
not \U$8765 ( \9108 , \6229 );
buf \U$8766 ( \9109 , \9108 );
not \U$8767 ( \9110 , \9109 );
nand \U$8768 ( \9111 , \9110 , \2700 );
nand \U$8769 ( \9112 , \9107 , \9111 );
nand \U$8770 ( \9113 , \9112 , \1702 );
nand \U$8771 ( \9114 , \9104 , \9113 );
xor \U$8772 ( \9115 , \9101 , \9114 );
not \U$8773 ( \9116 , \1570 );
not \U$8774 ( \9117 , \8767 );
or \U$8775 ( \9118 , \9116 , \9117 );
not \U$8776 ( \9119 , RIbb2f250_9);
not \U$8777 ( \9120 , \6268 );
or \U$8778 ( \9121 , \9119 , \9120 );
nand \U$8779 ( \9122 , \6269 , \1554 );
nand \U$8780 ( \9123 , \9121 , \9122 );
nand \U$8781 ( \9124 , \9123 , \1533 );
nand \U$8782 ( \9125 , \9118 , \9124 );
and \U$8783 ( \9126 , \9115 , \9125 );
and \U$8784 ( \9127 , \9101 , \9114 );
or \U$8785 ( \9128 , \9126 , \9127 );
and \U$8786 ( \9129 , \9086 , \9128 );
and \U$8787 ( \9130 , \9043 , \9085 );
or \U$8788 ( \9131 , \9129 , \9130 );
and \U$8789 ( \9132 , \9042 , \9131 );
and \U$8790 ( \9133 , \8987 , \9041 );
or \U$8791 ( \9134 , \9132 , \9133 );
xor \U$8792 ( \9135 , \8985 , \9134 );
xor \U$8793 ( \9136 , \7418 , \7431 );
xor \U$8794 ( \9137 , \9136 , \7441 );
not \U$8795 ( \9138 , \9137 );
not \U$8796 ( \9139 , \9138 );
xor \U$8797 ( \9140 , \7477 , \7465 );
xnor \U$8798 ( \9141 , \9140 , \7455 );
not \U$8799 ( \9142 , \9141 );
not \U$8800 ( \9143 , \9142 );
or \U$8801 ( \9144 , \9139 , \9143 );
nand \U$8802 ( \9145 , \9137 , \9141 );
nand \U$8803 ( \9146 , \9144 , \9145 );
xor \U$8804 ( \9147 , \8997 , \9002 );
and \U$8805 ( \9148 , \9147 , \9040 );
and \U$8806 ( \9149 , \8997 , \9002 );
or \U$8807 ( \9150 , \9148 , \9149 );
xor \U$8808 ( \9151 , \9146 , \9150 );
and \U$8809 ( \9152 , \9135 , \9151 );
and \U$8810 ( \9153 , \8985 , \9134 );
or \U$8811 ( \9154 , \9152 , \9153 );
xor \U$8812 ( \9155 , \8983 , \9154 );
xor \U$8813 ( \9156 , \8985 , \9134 );
xor \U$8814 ( \9157 , \9156 , \9151 );
not \U$8815 ( \9158 , \9157 );
xor \U$8816 ( \9159 , \8906 , \8941 );
xor \U$8817 ( \9160 , \9159 , \8969 );
buf \U$8818 ( \9161 , \9160 );
not \U$8819 ( \9162 , \9161 );
or \U$8820 ( \9163 , \9158 , \9162 );
or \U$8821 ( \9164 , \9157 , \9161 );
not \U$8822 ( \9165 , \2940 );
not \U$8823 ( \9166 , RIbb2e800_31);
not \U$8824 ( \9167 , \3773 );
or \U$8825 ( \9168 , \9166 , \9167 );
not \U$8826 ( \9169 , RIbb2e800_31);
nand \U$8827 ( \9170 , \1643 , \9169 );
nand \U$8828 ( \9171 , \9168 , \9170 );
not \U$8829 ( \9172 , \9171 );
or \U$8830 ( \9173 , \9165 , \9172 );
nand \U$8831 ( \9174 , \8804 , \3613 );
nand \U$8832 ( \9175 , \9173 , \9174 );
not \U$8833 ( \9176 , \9175 );
not \U$8834 ( \9177 , \9176 );
not \U$8835 ( \9178 , \2077 );
not \U$8836 ( \9179 , RIbb2ecb0_21);
not \U$8837 ( \9180 , \2224 );
or \U$8838 ( \9181 , \9179 , \9180 );
nand \U$8839 ( \9182 , \3320 , \849 );
nand \U$8840 ( \9183 , \9181 , \9182 );
not \U$8841 ( \9184 , \9183 );
or \U$8842 ( \9185 , \9178 , \9184 );
nand \U$8843 ( \9186 , \8689 , \2078 );
nand \U$8844 ( \9187 , \9185 , \9186 );
not \U$8845 ( \9188 , \9187 );
not \U$8846 ( \9189 , \9188 );
or \U$8847 ( \9190 , \9177 , \9189 );
not \U$8848 ( \9191 , \855 );
not \U$8849 ( \9192 , \8821 );
or \U$8850 ( \9193 , \9191 , \9192 );
not \U$8851 ( \9194 , RIbb2eda0_19);
not \U$8852 ( \9195 , \3168 );
or \U$8853 ( \9196 , \9194 , \9195 );
nand \U$8854 ( \9197 , \3167 , \1776 );
nand \U$8855 ( \9198 , \9196 , \9197 );
nand \U$8856 ( \9199 , \9198 , \853 );
nand \U$8857 ( \9200 , \9193 , \9199 );
nand \U$8858 ( \9201 , \9190 , \9200 );
nand \U$8859 ( \9202 , \9187 , \9175 );
nand \U$8860 ( \9203 , \9201 , \9202 );
not \U$8861 ( \9204 , \9203 );
xor \U$8862 ( \9205 , \8759 , \8769 );
xor \U$8863 ( \9206 , \9205 , \8780 );
not \U$8864 ( \9207 , \9206 );
or \U$8865 ( \9208 , \9204 , \9207 );
or \U$8866 ( \9209 , \9206 , \9203 );
xor \U$8867 ( \9210 , \8693 , \8712 );
xor \U$8868 ( \9211 , \9210 , \8682 );
nand \U$8869 ( \9212 , \9209 , \9211 );
nand \U$8870 ( \9213 , \9208 , \9212 );
xor \U$8871 ( \9214 , \8850 , \8903 );
xnor \U$8872 ( \9215 , \9214 , \8798 );
not \U$8873 ( \9216 , \9215 );
or \U$8874 ( \9217 , \9213 , \9216 );
xor \U$8875 ( \9218 , \8714 , \8747 );
xor \U$8876 ( \9219 , \9218 , \8783 );
nand \U$8877 ( \9220 , \9217 , \9219 );
nand \U$8878 ( \9221 , \9216 , \9213 );
nand \U$8879 ( \9222 , \9220 , \9221 );
nand \U$8880 ( \9223 , \9164 , \9222 );
nand \U$8881 ( \9224 , \9163 , \9223 );
xor \U$8882 ( \9225 , \9155 , \9224 );
xor \U$8883 ( \9226 , \7367 , \7354 );
and \U$8884 ( \9227 , \9226 , \7349 );
not \U$8885 ( \9228 , \9226 );
and \U$8886 ( \9229 , \9228 , \7352 );
nor \U$8887 ( \9230 , \9227 , \9229 );
not \U$8888 ( \9231 , \9230 );
xor \U$8889 ( \9232 , \7383 , \7394 );
xor \U$8890 ( \9233 , \9232 , \7405 );
not \U$8891 ( \9234 , \9233 );
not \U$8892 ( \9235 , \9234 );
or \U$8893 ( \9236 , \9231 , \9235 );
xor \U$8894 ( \9237 , \8568 , \8573 );
xor \U$8895 ( \9238 , \9237 , \8579 );
nand \U$8896 ( \9239 , \9236 , \9238 );
not \U$8897 ( \9240 , \9230 );
nand \U$8898 ( \9241 , \9240 , \9233 );
nand \U$8899 ( \9242 , \9239 , \9241 );
not \U$8900 ( \9243 , \9142 );
not \U$8901 ( \9244 , \9137 );
or \U$8902 ( \9245 , \9243 , \9244 );
or \U$8903 ( \9246 , \9137 , \9142 );
nand \U$8904 ( \9247 , \9246 , \9150 );
nand \U$8905 ( \9248 , \9245 , \9247 );
xor \U$8906 ( \9249 , \9242 , \9248 );
xor \U$8907 ( \9250 , \8555 , \8557 );
xor \U$8908 ( \9251 , \9250 , \8560 );
xor \U$8909 ( \9252 , \9249 , \9251 );
not \U$8910 ( \9253 , \9240 );
not \U$8911 ( \9254 , \9234 );
or \U$8912 ( \9255 , \9253 , \9254 );
nand \U$8913 ( \9256 , \9233 , \9230 );
nand \U$8914 ( \9257 , \9255 , \9256 );
xor \U$8915 ( \9258 , \9257 , \9238 );
xor \U$8916 ( \9259 , \8632 , \8646 );
xor \U$8917 ( \9260 , \9259 , \8657 );
xor \U$8918 ( \9261 , \9015 , \9029 );
xor \U$8919 ( \9262 , \9261 , \9037 );
or \U$8920 ( \9263 , \9260 , \9262 );
nor \U$8921 ( \9264 , \8608 , \602 );
not \U$8922 ( \9265 , \9264 );
not \U$8923 ( \9266 , \5941 );
or \U$8924 ( \9267 , \9265 , \9266 );
nor \U$8925 ( \9268 , \4364 , \602 );
nor \U$8926 ( \9269 , \9268 , \653 );
nand \U$8927 ( \9270 , \9267 , \9269 );
nand \U$8928 ( \9271 , \606 , \657 );
not \U$8929 ( \9272 , \9271 );
and \U$8930 ( \9273 , \9270 , \9272 );
not \U$8931 ( \9274 , \9270 );
and \U$8932 ( \9275 , \9274 , \9271 );
nor \U$8933 ( \9276 , \9273 , \9275 );
buf \U$8934 ( \9277 , \9276 );
buf \U$8935 ( \9278 , \9277 );
not \U$8936 ( \9279 , \9278 );
not \U$8937 ( \9280 , \9279 );
nand \U$8938 ( \9281 , \9280 , \1393 );
not \U$8939 ( \9282 , \9281 );
not \U$8940 ( \9283 , \9282 );
not \U$8941 ( \9284 , \2922 );
not \U$8942 ( \9285 , RIbb2e8f0_29);
not \U$8943 ( \9286 , \4766 );
or \U$8944 ( \9287 , \9285 , \9286 );
nand \U$8945 ( \9288 , \4770 , \3440 );
nand \U$8946 ( \9289 , \9287 , \9288 );
not \U$8947 ( \9290 , \9289 );
or \U$8948 ( \9291 , \9284 , \9290 );
not \U$8949 ( \9292 , \4460 );
nand \U$8950 ( \9293 , \9292 , \8866 );
nand \U$8951 ( \9294 , \9291 , \9293 );
not \U$8952 ( \9295 , \9294 );
or \U$8953 ( \9296 , \9283 , \9295 );
or \U$8954 ( \9297 , \9294 , \9282 );
not \U$8955 ( \9298 , \916 );
not \U$8956 ( \9299 , RIbb2f070_13);
not \U$8957 ( \9300 , \4029 );
or \U$8958 ( \9301 , \9299 , \9300 );
nand \U$8959 ( \9302 , \3046 , \3421 );
nand \U$8960 ( \9303 , \9301 , \9302 );
not \U$8961 ( \9304 , \9303 );
or \U$8962 ( \9305 , \9298 , \9304 );
nand \U$8963 ( \9306 , \8876 , \998 );
nand \U$8964 ( \9307 , \9305 , \9306 );
nand \U$8965 ( \9308 , \9297 , \9307 );
nand \U$8966 ( \9309 , \9296 , \9308 );
nand \U$8967 ( \9310 , \9263 , \9309 );
nand \U$8968 ( \9311 , \9260 , \9262 );
nand \U$8969 ( \9312 , \9310 , \9311 );
not \U$8970 ( \9313 , \9312 );
not \U$8971 ( \9314 , \9313 );
not \U$8972 ( \9315 , \1533 );
and \U$8973 ( \9316 , \6199 , RIbb2f250_9);
not \U$8974 ( \9317 , \6199 );
and \U$8975 ( \9318 , \9317 , \1554 );
or \U$8976 ( \9319 , \9316 , \9318 );
not \U$8977 ( \9320 , \9319 );
or \U$8978 ( \9321 , \9315 , \9320 );
nand \U$8979 ( \9322 , \9123 , \1570 );
nand \U$8980 ( \9323 , \9321 , \9322 );
not \U$8981 ( \9324 , \836 );
not \U$8982 ( \9325 , \8839 );
or \U$8983 ( \9326 , \9324 , \9325 );
not \U$8984 ( \9327 , RIbb2ee90_17);
not \U$8985 ( \9328 , \3203 );
or \U$8986 ( \9329 , \9327 , \9328 );
nand \U$8987 ( \9330 , \4640 , \3699 );
nand \U$8988 ( \9331 , \9329 , \9330 );
nand \U$8989 ( \9332 , \9331 , \832 );
nand \U$8990 ( \9333 , \9326 , \9332 );
xor \U$8991 ( \9334 , \9323 , \9333 );
not \U$8992 ( \9335 , \1445 );
and \U$8993 ( \9336 , RIbb2ef80_15, \3655 );
not \U$8994 ( \9337 , RIbb2ef80_15);
and \U$8995 ( \9338 , \9337 , \3654 );
or \U$8996 ( \9339 , \9336 , \9338 );
not \U$8997 ( \9340 , \9339 );
or \U$8998 ( \9341 , \9335 , \9340 );
nand \U$8999 ( \9342 , \8892 , \1517 );
nand \U$9000 ( \9343 , \9341 , \9342 );
and \U$9001 ( \9344 , \9334 , \9343 );
and \U$9002 ( \9345 , \9323 , \9333 );
or \U$9003 ( \9346 , \9344 , \9345 );
not \U$9004 ( \9347 , \9346 );
xor \U$9005 ( \9348 , \8724 , \8734 );
xor \U$9006 ( \9349 , \9348 , \8744 );
not \U$9007 ( \9350 , \9349 );
or \U$9008 ( \9351 , \9347 , \9350 );
or \U$9009 ( \9352 , \9349 , \9346 );
xor \U$9010 ( \9353 , \8848 , \8830 );
not \U$9011 ( \9354 , \8814 );
and \U$9012 ( \9355 , \9353 , \9354 );
not \U$9013 ( \9356 , \9353 );
and \U$9014 ( \9357 , \9356 , \8814 );
nor \U$9015 ( \9358 , \9355 , \9357 );
not \U$9016 ( \9359 , \9358 );
nand \U$9017 ( \9360 , \9352 , \9359 );
nand \U$9018 ( \9361 , \9351 , \9360 );
not \U$9019 ( \9362 , \9361 );
not \U$9020 ( \9363 , \9362 );
or \U$9021 ( \9364 , \9314 , \9363 );
not \U$9022 ( \9365 , \5845 );
not \U$9023 ( \9366 , \8722 );
or \U$9024 ( \9367 , \9365 , \9366 );
not \U$9025 ( \9368 , RIbb2e620_35);
not \U$9026 ( \9369 , \1562 );
or \U$9027 ( \9370 , \9368 , \9369 );
nand \U$9028 ( \9371 , \1038 , \6002 );
nand \U$9029 ( \9372 , \9370 , \9371 );
nand \U$9030 ( \9373 , \9372 , \4712 );
nand \U$9031 ( \9374 , \9367 , \9373 );
not \U$9032 ( \9375 , \6242 );
not \U$9033 ( \9376 , \8710 );
or \U$9034 ( \9377 , \9375 , \9376 );
not \U$9035 ( \9378 , \6252 );
not \U$9036 ( \9379 , RIbb2e530_37);
not \U$9037 ( \9380 , \951 );
or \U$9038 ( \9381 , \9379 , \9380 );
nand \U$9039 ( \9382 , \952 , \4708 );
nand \U$9040 ( \9383 , \9381 , \9382 );
nand \U$9041 ( \9384 , \9378 , \9383 );
nand \U$9042 ( \9385 , \9377 , \9384 );
or \U$9043 ( \9386 , \9374 , \9385 );
not \U$9044 ( \9387 , \2980 );
xor \U$9045 ( \9388 , RIbb2ead0_25, \3821 );
not \U$9046 ( \9389 , \9388 );
or \U$9047 ( \9390 , \9387 , \9389 );
nand \U$9048 ( \9391 , \8742 , \2963 );
nand \U$9049 ( \9392 , \9390 , \9391 );
nand \U$9050 ( \9393 , \9386 , \9392 );
nand \U$9051 ( \9394 , \9374 , \9385 );
nand \U$9052 ( \9395 , \9393 , \9394 );
not \U$9053 ( \9396 , \9395 );
not \U$9054 ( \9397 , \9396 );
not \U$9055 ( \9398 , \8362 );
not \U$9056 ( \9399 , RIbb2e350_41);
not \U$9057 ( \9400 , \894 );
or \U$9058 ( \9401 , \9399 , \9400 );
not \U$9059 ( \9402 , RIbb2e350_41);
nand \U$9060 ( \9403 , \893 , \9402 );
nand \U$9061 ( \9404 , \9401 , \9403 );
not \U$9062 ( \9405 , \9404 );
or \U$9063 ( \9406 , \9398 , \9405 );
nand \U$9064 ( \9407 , \8992 , \8995 );
nand \U$9065 ( \9408 , \9406 , \9407 );
not \U$9066 ( \9409 , \9408 );
not \U$9067 ( \9410 , \1011 );
not \U$9068 ( \9411 , RIbb2f160_11);
not \U$9069 ( \9412 , \4749 );
or \U$9070 ( \9413 , \9411 , \9412 );
nand \U$9071 ( \9414 , \4753 , \1805 );
nand \U$9072 ( \9415 , \9413 , \9414 );
not \U$9073 ( \9416 , \9415 );
or \U$9074 ( \9417 , \9410 , \9416 );
nand \U$9075 ( \9418 , \8778 , \1077 );
nand \U$9076 ( \9419 , \9417 , \9418 );
not \U$9077 ( \9420 , \9419 );
or \U$9078 ( \9421 , \9409 , \9420 );
or \U$9079 ( \9422 , \9408 , \9419 );
not \U$9080 ( \9423 , \3465 );
not \U$9081 ( \9424 , \8653 );
or \U$9082 ( \9425 , \9423 , \9424 );
not \U$9083 ( \9426 , \6071 );
not \U$9084 ( \9427 , RIbb2e9e0_27);
not \U$9085 ( \9428 , \3991 );
or \U$9086 ( \9429 , \9427 , \9428 );
nand \U$9087 ( \9430 , \3736 , \4598 );
nand \U$9088 ( \9431 , \9429 , \9430 );
nand \U$9089 ( \9432 , \9426 , \9431 );
nand \U$9090 ( \9433 , \9425 , \9432 );
nand \U$9091 ( \9434 , \9422 , \9433 );
nand \U$9092 ( \9435 , \9421 , \9434 );
not \U$9093 ( \9436 , \9435 );
not \U$9094 ( \9437 , \9436 );
or \U$9095 ( \9438 , \9397 , \9437 );
not \U$9096 ( \9439 , \8445 );
and \U$9097 ( \9440 , RIbb2e440_39, \1475 );
not \U$9098 ( \9441 , RIbb2e440_39);
and \U$9099 ( \9442 , \9441 , \1474 );
or \U$9100 ( \9443 , \9440 , \9442 );
not \U$9101 ( \9444 , \9443 );
or \U$9102 ( \9445 , \9439 , \9444 );
nand \U$9103 ( \9446 , \8757 , \7104 );
nand \U$9104 ( \9447 , \9445 , \9446 );
not \U$9105 ( \9448 , \3887 );
not \U$9106 ( \9449 , RIbb2e710_33);
not \U$9107 ( \9450 , \3479 );
or \U$9108 ( \9451 , \9449 , \9450 );
nand \U$9109 ( \9452 , \3484 , \2935 );
nand \U$9110 ( \9453 , \9451 , \9452 );
not \U$9111 ( \9454 , \9453 );
or \U$9112 ( \9455 , \9448 , \9454 );
nand \U$9113 ( \9456 , \8680 , \4791 );
nand \U$9114 ( \9457 , \9455 , \9456 );
or \U$9115 ( \9458 , \9447 , \9457 );
not \U$9116 ( \9459 , \3406 );
not \U$9117 ( \9460 , RIbb2ebc0_23);
not \U$9118 ( \9461 , \4609 );
or \U$9119 ( \9462 , \9460 , \9461 );
nand \U$9120 ( \9463 , \3810 , \3396 );
nand \U$9121 ( \9464 , \9462 , \9463 );
not \U$9122 ( \9465 , \9464 );
or \U$9123 ( \9466 , \9459 , \9465 );
nand \U$9124 ( \9467 , \3383 , \8732 );
nand \U$9125 ( \9468 , \9466 , \9467 );
nand \U$9126 ( \9469 , \9458 , \9468 );
nand \U$9127 ( \9470 , \9457 , \9447 );
nand \U$9128 ( \9471 , \9469 , \9470 );
nand \U$9129 ( \9472 , \9438 , \9471 );
nand \U$9130 ( \9473 , \9435 , \9395 );
nand \U$9131 ( \9474 , \9472 , \9473 );
nand \U$9132 ( \9475 , \9364 , \9474 );
not \U$9133 ( \9476 , \9313 );
nand \U$9134 ( \9477 , \9476 , \9361 );
nand \U$9135 ( \9478 , \9475 , \9477 );
xor \U$9136 ( \9479 , \9258 , \9478 );
xor \U$9137 ( \9480 , \8669 , \8671 );
xor \U$9138 ( \9481 , \9480 , \8786 );
and \U$9139 ( \9482 , \9479 , \9481 );
and \U$9140 ( \9483 , \9258 , \9478 );
or \U$9141 ( \9484 , \9482 , \9483 );
xor \U$9142 ( \9485 , \9252 , \9484 );
xor \U$9143 ( \9486 , \8604 , \8789 );
xor \U$9144 ( \9487 , \9486 , \8792 );
xor \U$9145 ( \9488 , \9485 , \9487 );
and \U$9146 ( \9489 , \9225 , \9488 );
and \U$9147 ( \9490 , \9155 , \9224 );
or \U$9148 ( \9491 , \9489 , \9490 );
xor \U$9149 ( \9492 , \8796 , \9491 );
xor \U$9150 ( \9493 , \8972 , \8982 );
and \U$9151 ( \9494 , \9493 , \9154 );
and \U$9152 ( \9495 , \8972 , \8982 );
or \U$9153 ( \9496 , \9494 , \9495 );
xor \U$9154 ( \9497 , \8976 , \8978 );
and \U$9155 ( \9498 , \9497 , \8981 );
and \U$9156 ( \9499 , \8976 , \8978 );
or \U$9157 ( \9500 , \9498 , \9499 );
xor \U$9158 ( \9501 , \9242 , \9248 );
and \U$9159 ( \9502 , \9501 , \9251 );
and \U$9160 ( \9503 , \9242 , \9248 );
or \U$9161 ( \9504 , \9502 , \9503 );
xor \U$9162 ( \9505 , \9500 , \9504 );
xor \U$9163 ( \9506 , \7214 , \7177 );
xor \U$9164 ( \9507 , \9506 , \7252 );
xor \U$9165 ( \9508 , \6922 , \6964 );
xor \U$9166 ( \9509 , \9508 , \6999 );
xor \U$9167 ( \9510 , \9507 , \9509 );
not \U$9168 ( \9511 , \7052 );
not \U$9169 ( \9512 , \9511 );
not \U$9170 ( \9513 , \7061 );
or \U$9171 ( \9514 , \9512 , \9513 );
nand \U$9172 ( \9515 , \7060 , \7052 );
nand \U$9173 ( \9516 , \9514 , \9515 );
xor \U$9174 ( \9517 , \7057 , \9516 );
xor \U$9175 ( \9518 , \9510 , \9517 );
xor \U$9176 ( \9519 , \9505 , \9518 );
xor \U$9177 ( \9520 , \9496 , \9519 );
xor \U$9178 ( \9521 , \9252 , \9484 );
and \U$9179 ( \9522 , \9521 , \9487 );
and \U$9180 ( \9523 , \9252 , \9484 );
or \U$9181 ( \9524 , \9522 , \9523 );
xor \U$9182 ( \9525 , \9520 , \9524 );
and \U$9183 ( \9526 , \9492 , \9525 );
and \U$9184 ( \9527 , \8796 , \9491 );
or \U$9185 ( \9528 , \9526 , \9527 );
not \U$9186 ( \9529 , \9528 );
and \U$9187 ( \9530 , \6910 , \6906 );
not \U$9188 ( \9531 , \6910 );
and \U$9189 ( \9532 , \9531 , \6905 );
nor \U$9190 ( \9533 , \9530 , \9532 );
xor \U$9191 ( \9534 , \9533 , \6914 );
xor \U$9192 ( \9535 , \7255 , \7486 );
xor \U$9193 ( \9536 , \9535 , \7262 );
xor \U$9194 ( \9537 , \9534 , \9536 );
xor \U$9195 ( \9538 , \8303 , \8305 );
and \U$9196 ( \9539 , \9538 , \8534 );
and \U$9197 ( \9540 , \8303 , \8305 );
or \U$9198 ( \9541 , \9539 , \9540 );
xor \U$9199 ( \9542 , \9537 , \9541 );
not \U$9200 ( \9543 , \9542 );
not \U$9201 ( \9544 , \9500 );
not \U$9202 ( \9545 , \9504 );
or \U$9203 ( \9546 , \9544 , \9545 );
or \U$9204 ( \9547 , \9504 , \9500 );
nand \U$9205 ( \9548 , \9547 , \9518 );
nand \U$9206 ( \9549 , \9546 , \9548 );
or \U$9207 ( \9550 , \8599 , \8588 );
nand \U$9208 ( \9551 , \9550 , \8563 );
nand \U$9209 ( \9552 , \8599 , \8588 );
nand \U$9210 ( \9553 , \9551 , \9552 );
xor \U$9211 ( \9554 , \7002 , \7049 );
xor \U$9212 ( \9555 , \9554 , \7064 );
xor \U$9213 ( \9556 , \9553 , \9555 );
xor \U$9214 ( \9557 , \9507 , \9509 );
and \U$9215 ( \9558 , \9557 , \9517 );
and \U$9216 ( \9559 , \9507 , \9509 );
or \U$9217 ( \9560 , \9558 , \9559 );
xor \U$9218 ( \9561 , \9556 , \9560 );
xor \U$9219 ( \9562 , \9549 , \9561 );
not \U$9220 ( \9563 , \8601 );
not \U$9221 ( \9564 , \8535 );
or \U$9222 ( \9565 , \9563 , \9564 );
or \U$9223 ( \9566 , \8535 , \8601 );
nand \U$9224 ( \9567 , \9566 , \8795 );
nand \U$9225 ( \9568 , \9565 , \9567 );
xnor \U$9226 ( \9569 , \9562 , \9568 );
not \U$9227 ( \9570 , \9569 );
or \U$9228 ( \9571 , \9543 , \9570 );
or \U$9229 ( \9572 , \9569 , \9542 );
nand \U$9230 ( \9573 , \9571 , \9572 );
xor \U$9231 ( \9574 , \9496 , \9519 );
and \U$9232 ( \9575 , \9574 , \9524 );
and \U$9233 ( \9576 , \9496 , \9519 );
or \U$9234 ( \9577 , \9575 , \9576 );
not \U$9235 ( \9578 , \9577 );
and \U$9236 ( \9579 , \9573 , \9578 );
not \U$9237 ( \9580 , \9573 );
and \U$9238 ( \9581 , \9580 , \9577 );
nor \U$9239 ( \9582 , \9579 , \9581 );
nand \U$9240 ( \9583 , \9529 , \9582 );
not \U$9241 ( \9584 , \9542 );
not \U$9242 ( \9585 , \9584 );
not \U$9243 ( \9586 , \9569 );
or \U$9244 ( \9587 , \9585 , \9586 );
nand \U$9245 ( \9588 , \9587 , \9577 );
not \U$9246 ( \9589 , \9569 );
nand \U$9247 ( \9590 , \9589 , \9542 );
nand \U$9248 ( \9591 , \9588 , \9590 );
not \U$9249 ( \9592 , \9591 );
xor \U$9250 ( \9593 , \9534 , \9536 );
and \U$9251 ( \9594 , \9593 , \9541 );
and \U$9252 ( \9595 , \9534 , \9536 );
or \U$9253 ( \9596 , \9594 , \9595 );
not \U$9254 ( \9597 , \9596 );
not \U$9255 ( \9598 , \9597 );
xor \U$9256 ( \9599 , \9553 , \9555 );
and \U$9257 ( \9600 , \9599 , \9560 );
and \U$9258 ( \9601 , \9553 , \9555 );
or \U$9259 ( \9602 , \9600 , \9601 );
xor \U$9260 ( \9603 , \6917 , \6919 );
xor \U$9261 ( \9604 , \9603 , \7067 );
not \U$9262 ( \9605 , \9604 );
and \U$9263 ( \9606 , \9602 , \9605 );
not \U$9264 ( \9607 , \9602 );
and \U$9265 ( \9608 , \9607 , \9604 );
or \U$9266 ( \9609 , \9606 , \9608 );
not \U$9267 ( \9610 , \7488 );
not \U$9268 ( \9611 , \7496 );
or \U$9269 ( \9612 , \9610 , \9611 );
or \U$9270 ( \9613 , \7496 , \7488 );
nand \U$9271 ( \9614 , \9612 , \9613 );
xor \U$9272 ( \9615 , \9614 , \7508 );
not \U$9273 ( \9616 , \9615 );
and \U$9274 ( \9617 , \9609 , \9616 );
not \U$9275 ( \9618 , \9609 );
and \U$9276 ( \9619 , \9618 , \9615 );
nor \U$9277 ( \9620 , \9617 , \9619 );
not \U$9278 ( \9621 , \9620 );
not \U$9279 ( \9622 , \9621 );
or \U$9280 ( \9623 , \9598 , \9622 );
nand \U$9281 ( \9624 , \9620 , \9596 );
nand \U$9282 ( \9625 , \9623 , \9624 );
not \U$9283 ( \9626 , \9561 );
not \U$9284 ( \9627 , \9568 );
or \U$9285 ( \9628 , \9626 , \9627 );
or \U$9286 ( \9629 , \9561 , \9568 );
nand \U$9287 ( \9630 , \9629 , \9549 );
nand \U$9288 ( \9631 , \9628 , \9630 );
not \U$9289 ( \9632 , \9631 );
and \U$9290 ( \9633 , \9625 , \9632 );
not \U$9291 ( \9634 , \9625 );
and \U$9292 ( \9635 , \9634 , \9631 );
nor \U$9293 ( \9636 , \9633 , \9635 );
nand \U$9294 ( \9637 , \9592 , \9636 );
not \U$9295 ( \9638 , \9597 );
not \U$9296 ( \9639 , \9620 );
or \U$9297 ( \9640 , \9638 , \9639 );
nand \U$9298 ( \9641 , \9640 , \9631 );
nand \U$9299 ( \9642 , \9621 , \9596 );
nand \U$9300 ( \9643 , \9641 , \9642 );
not \U$9301 ( \9644 , \9643 );
xor \U$9302 ( \9645 , \7516 , \7518 );
xor \U$9303 ( \9646 , \9645 , \7523 );
not \U$9304 ( \9647 , \9646 );
not \U$9305 ( \9648 , \9647 );
and \U$9306 ( \9649 , \7080 , \7070 );
not \U$9307 ( \9650 , \7080 );
not \U$9308 ( \9651 , \7070 );
and \U$9309 ( \9652 , \9650 , \9651 );
nor \U$9310 ( \9653 , \9649 , \9652 );
buf \U$9311 ( \9654 , \7512 );
not \U$9312 ( \9655 , \9654 );
and \U$9313 ( \9656 , \9653 , \9655 );
not \U$9314 ( \9657 , \9653 );
and \U$9315 ( \9658 , \9657 , \9654 );
nor \U$9316 ( \9659 , \9656 , \9658 );
not \U$9317 ( \9660 , \9659 );
not \U$9318 ( \9661 , \9660 );
or \U$9319 ( \9662 , \9648 , \9661 );
nand \U$9320 ( \9663 , \9659 , \9646 );
nand \U$9321 ( \9664 , \9662 , \9663 );
not \U$9322 ( \9665 , \9604 );
not \U$9323 ( \9666 , \9615 );
or \U$9324 ( \9667 , \9665 , \9666 );
not \U$9325 ( \9668 , \9605 );
not \U$9326 ( \9669 , \9616 );
or \U$9327 ( \9670 , \9668 , \9669 );
nand \U$9328 ( \9671 , \9670 , \9602 );
nand \U$9329 ( \9672 , \9667 , \9671 );
xnor \U$9330 ( \9673 , \9664 , \9672 );
nand \U$9331 ( \9674 , \9644 , \9673 );
and \U$9332 ( \9675 , \9583 , \9637 , \9674 );
nand \U$9333 ( \9676 , \8664 , \8668 );
xnor \U$9334 ( \9677 , \9676 , \8606 );
not \U$9335 ( \9678 , \8926 );
not \U$9336 ( \9679 , \9678 );
not \U$9337 ( \9680 , \8939 );
or \U$9338 ( \9681 , \9679 , \9680 );
nand \U$9339 ( \9682 , \8938 , \8926 );
nand \U$9340 ( \9683 , \9681 , \9682 );
buf \U$9341 ( \9684 , \8908 );
xor \U$9342 ( \9685 , \9683 , \9684 );
xor \U$9343 ( \9686 , \9677 , \9685 );
xor \U$9344 ( \9687 , \8868 , \8901 );
xor \U$9345 ( \9688 , \9687 , \8884 );
xor \U$9346 ( \9689 , \9043 , \9085 );
xor \U$9347 ( \9690 , \9689 , \9128 );
xor \U$9348 ( \9691 , \9688 , \9690 );
not \U$9349 ( \9692 , \2940 );
not \U$9350 ( \9693 , RIbb2e800_31);
not \U$9351 ( \9694 , \3054 );
or \U$9352 ( \9695 , \9693 , \9694 );
nand \U$9353 ( \9696 , \1138 , \2917 );
nand \U$9354 ( \9697 , \9695 , \9696 );
not \U$9355 ( \9698 , \9697 );
or \U$9356 ( \9699 , \9692 , \9698 );
nand \U$9357 ( \9700 , \9171 , \3613 );
nand \U$9358 ( \9701 , \9699 , \9700 );
not \U$9359 ( \9702 , \9701 );
not \U$9360 ( \9703 , \853 );
not \U$9361 ( \9704 , RIbb2eda0_19);
not \U$9362 ( \9705 , \3141 );
or \U$9363 ( \9706 , \9704 , \9705 );
not \U$9364 ( \9707 , \3141 );
nand \U$9365 ( \9708 , \9707 , \3251 );
nand \U$9366 ( \9709 , \9706 , \9708 );
not \U$9367 ( \9710 , \9709 );
or \U$9368 ( \9711 , \9703 , \9710 );
nand \U$9369 ( \9712 , \9198 , \855 );
nand \U$9370 ( \9713 , \9711 , \9712 );
not \U$9371 ( \9714 , \9713 );
or \U$9372 ( \9715 , \9702 , \9714 );
or \U$9373 ( \9716 , \9713 , \9701 );
not \U$9374 ( \9717 , \832 );
not \U$9375 ( \9718 , RIbb2ee90_17);
not \U$9376 ( \9719 , \3226 );
or \U$9377 ( \9720 , \9718 , \9719 );
nand \U$9378 ( \9721 , \3228 , \816 );
nand \U$9379 ( \9722 , \9720 , \9721 );
not \U$9380 ( \9723 , \9722 );
or \U$9381 ( \9724 , \9717 , \9723 );
nand \U$9382 ( \9725 , \9331 , \836 );
nand \U$9383 ( \9726 , \9724 , \9725 );
nand \U$9384 ( \9727 , \9716 , \9726 );
nand \U$9385 ( \9728 , \9715 , \9727 );
xor \U$9386 ( \9729 , \9101 , \9114 );
xor \U$9387 ( \9730 , \9729 , \9125 );
nor \U$9388 ( \9731 , \9728 , \9730 );
not \U$9389 ( \9732 , \1077 );
not \U$9390 ( \9733 , \9415 );
or \U$9391 ( \9734 , \9732 , \9733 );
not \U$9392 ( \9735 , RIbb2f160_11);
not \U$9393 ( \9736 , \4325 );
or \U$9394 ( \9737 , \9735 , \9736 );
nand \U$9395 ( \9738 , \4324 , \1043 );
nand \U$9396 ( \9739 , \9737 , \9738 );
nand \U$9397 ( \9740 , \9739 , \1011 );
nand \U$9398 ( \9741 , \9734 , \9740 );
not \U$9399 ( \9742 , \2922 );
not \U$9400 ( \9743 , RIbb2e8f0_29);
not \U$9401 ( \9744 , \3290 );
or \U$9402 ( \9745 , \9743 , \9744 );
nand \U$9403 ( \9746 , \1283 , \3440 );
nand \U$9404 ( \9747 , \9745 , \9746 );
not \U$9405 ( \9748 , \9747 );
or \U$9406 ( \9749 , \9742 , \9748 );
nand \U$9407 ( \9750 , \9289 , \2925 );
nand \U$9408 ( \9751 , \9749 , \9750 );
xor \U$9409 ( \9752 , \9741 , \9751 );
not \U$9410 ( \9753 , \916 );
not \U$9411 ( \9754 , \906 );
not \U$9412 ( \9755 , \3003 );
or \U$9413 ( \9756 , \9754 , \9755 );
not \U$9414 ( \9757 , \3275 );
nand \U$9415 ( \9758 , \9757 , RIbb2f070_13);
nand \U$9416 ( \9759 , \9756 , \9758 );
not \U$9417 ( \9760 , \9759 );
or \U$9418 ( \9761 , \9753 , \9760 );
nand \U$9419 ( \9762 , \9303 , \998 );
nand \U$9420 ( \9763 , \9761 , \9762 );
and \U$9421 ( \9764 , \9752 , \9763 );
and \U$9422 ( \9765 , \9741 , \9751 );
or \U$9423 ( \9766 , \9764 , \9765 );
not \U$9424 ( \9767 , \9766 );
or \U$9425 ( \9768 , \9731 , \9767 );
nand \U$9426 ( \9769 , \9728 , \9730 );
nand \U$9427 ( \9770 , \9768 , \9769 );
and \U$9428 ( \9771 , \9691 , \9770 );
and \U$9429 ( \9772 , \9688 , \9690 );
or \U$9430 ( \9773 , \9771 , \9772 );
and \U$9431 ( \9774 , \9686 , \9773 );
and \U$9432 ( \9775 , \9677 , \9685 );
or \U$9433 ( \9776 , \9774 , \9775 );
xor \U$9434 ( \9777 , \8987 , \9041 );
xor \U$9435 ( \9778 , \9777 , \9131 );
not \U$9436 ( \9779 , \9778 );
xor \U$9437 ( \9780 , \9474 , \9313 );
xnor \U$9438 ( \9781 , \9780 , \9362 );
not \U$9439 ( \9782 , \9781 );
not \U$9440 ( \9783 , \9782 );
or \U$9441 ( \9784 , \9779 , \9783 );
not \U$9442 ( \9785 , \9778 );
not \U$9443 ( \9786 , \9785 );
not \U$9444 ( \9787 , \9781 );
or \U$9445 ( \9788 , \9786 , \9787 );
not \U$9446 ( \9789 , \1090 );
not \U$9447 ( \9790 , RIbb2f430_5);
not \U$9448 ( \9791 , \8638 );
not \U$9449 ( \9792 , \9791 );
or \U$9450 ( \9793 , \9790 , \9792 );
nand \U$9451 ( \9794 , \8638 , \1085 );
nand \U$9452 ( \9795 , \9793 , \9794 );
not \U$9453 ( \9796 , \9795 );
or \U$9454 ( \9797 , \9789 , \9796 );
nand \U$9455 ( \9798 , \9062 , \1147 );
nand \U$9456 ( \9799 , \9797 , \9798 );
not \U$9457 ( \9800 , \1702 );
not \U$9458 ( \9801 , RIbb2f340_7);
not \U$9459 ( \9802 , \5956 );
or \U$9460 ( \9803 , \9801 , \9802 );
nand \U$9461 ( \9804 , \5955 , \1734 );
nand \U$9462 ( \9805 , \9803 , \9804 );
not \U$9463 ( \9806 , \9805 );
or \U$9464 ( \9807 , \9800 , \9806 );
nand \U$9465 ( \9808 , \9112 , \1737 );
nand \U$9466 ( \9809 , \9807 , \9808 );
nand \U$9467 ( \9810 , \9799 , \9809 );
not \U$9468 ( \9811 , \9810 );
not \U$9469 ( \9812 , \9799 );
not \U$9470 ( \9813 , \9809 );
and \U$9471 ( \9814 , \9812 , \9813 );
not \U$9472 ( \9815 , \8321 );
not \U$9473 ( \9816 , \1245 );
and \U$9474 ( \9817 , \9815 , \9816 );
buf \U$9475 ( \9818 , \8318 );
buf \U$9476 ( \9819 , \9818 );
and \U$9477 ( \9820 , \9819 , \1245 );
nor \U$9478 ( \9821 , \9817 , \9820 );
not \U$9479 ( \9822 , \9821 );
not \U$9480 ( \9823 , \1266 );
and \U$9481 ( \9824 , \9822 , \9823 );
and \U$9482 ( \9825 , \9076 , \1294 );
nor \U$9483 ( \9826 , \9824 , \9825 );
nor \U$9484 ( \9827 , \9814 , \9826 );
nor \U$9485 ( \9828 , \9811 , \9827 );
not \U$9486 ( \9829 , \9828 );
not \U$9487 ( \9830 , \9829 );
nor \U$9488 ( \9831 , \8608 , \509 );
not \U$9489 ( \9832 , \9831 );
not \U$9490 ( \9833 , \4360 );
or \U$9491 ( \9834 , \9832 , \9833 );
nor \U$9492 ( \9835 , \4364 , \509 );
nor \U$9493 ( \9836 , \9835 , \648 );
nand \U$9494 ( \9837 , \9834 , \9836 );
nand \U$9495 ( \9838 , \600 , \652 );
xnor \U$9496 ( \9839 , \9837 , \9838 );
buf \U$9497 ( \9840 , \9839 );
buf \U$9498 ( \9841 , \9840 );
nand \U$9499 ( \9842 , \9841 , \1313 );
not \U$9500 ( \9843 , \9098 );
not \U$9501 ( \9844 , RIbb2e260_43);
not \U$9502 ( \9845 , \5638 );
or \U$9503 ( \9846 , \9844 , \9845 );
not \U$9504 ( \9847 , RIbb2e260_43);
nand \U$9505 ( \9848 , \2251 , \9847 );
nand \U$9506 ( \9849 , \9846 , \9848 );
not \U$9507 ( \9850 , \9849 );
or \U$9508 ( \9851 , \9843 , \9850 );
nand \U$9509 ( \9852 , \9099 , RIbb2e260_43);
nand \U$9510 ( \9853 , \9851 , \9852 );
not \U$9511 ( \9854 , \9853 );
xor \U$9512 ( \9855 , \9842 , \9854 );
not \U$9513 ( \9856 , \1313 );
not \U$9514 ( \9857 , \9278 );
not \U$9515 ( \9858 , \9857 );
or \U$9516 ( \9859 , \9856 , \9858 );
not \U$9517 ( \9860 , \9857 );
nand \U$9518 ( \9861 , \9860 , \1951 );
nand \U$9519 ( \9862 , \9859 , \9861 );
and \U$9520 ( \9863 , \9862 , \1429 );
and \U$9521 ( \9864 , \9045 , \1376 );
nor \U$9522 ( \9865 , \9863 , \9864 );
and \U$9523 ( \9866 , \9855 , \9865 );
and \U$9524 ( \9867 , \9842 , \9854 );
or \U$9525 ( \9868 , \9866 , \9867 );
not \U$9526 ( \9869 , \9868 );
not \U$9527 ( \9870 , \9869 );
or \U$9528 ( \9871 , \9830 , \9870 );
not \U$9529 ( \9872 , \9868 );
not \U$9530 ( \9873 , \9828 );
or \U$9531 ( \9874 , \9872 , \9873 );
not \U$9532 ( \9875 , \9064 );
not \U$9533 ( \9876 , \9081 );
or \U$9534 ( \9877 , \9875 , \9876 );
or \U$9535 ( \9878 , \9081 , \9064 );
nand \U$9536 ( \9879 , \9877 , \9878 );
and \U$9537 ( \9880 , \9879 , \9049 );
not \U$9538 ( \9881 , \9879 );
and \U$9539 ( \9882 , \9881 , \9050 );
nor \U$9540 ( \9883 , \9880 , \9882 );
nand \U$9541 ( \9884 , \9874 , \9883 );
nand \U$9542 ( \9885 , \9871 , \9884 );
not \U$9543 ( \9886 , \6242 );
not \U$9544 ( \9887 , \9383 );
or \U$9545 ( \9888 , \9886 , \9887 );
not \U$9546 ( \9889 , RIbb2e530_37);
not \U$9547 ( \9890 , \1887 );
or \U$9548 ( \9891 , \9889 , \9890 );
nand \U$9549 ( \9892 , \1071 , \6246 );
nand \U$9550 ( \9893 , \9891 , \9892 );
nand \U$9551 ( \9894 , \9893 , \6251 );
nand \U$9552 ( \9895 , \9888 , \9894 );
not \U$9553 ( \9896 , \8995 );
not \U$9554 ( \9897 , \9404 );
or \U$9555 ( \9898 , \9896 , \9897 );
not \U$9556 ( \9899 , RIbb2e350_41);
not \U$9557 ( \9900 , \3262 );
or \U$9558 ( \9901 , \9899 , \9900 );
nand \U$9559 ( \9902 , \4315 , \9402 );
nand \U$9560 ( \9903 , \9901 , \9902 );
nand \U$9561 ( \9904 , \9903 , \8362 );
nand \U$9562 ( \9905 , \9898 , \9904 );
nor \U$9563 ( \9906 , \9895 , \9905 );
and \U$9564 ( \9907 , \9431 , \3465 );
not \U$9565 ( \9908 , RIbb2e9e0_27);
not \U$9566 ( \9909 , \4341 );
or \U$9567 ( \9910 , \9908 , \9909 );
nand \U$9568 ( \9911 , \1387 , \6065 );
nand \U$9569 ( \9912 , \9910 , \9911 );
not \U$9570 ( \9913 , \9912 );
nor \U$9571 ( \9914 , \9913 , \6071 );
nor \U$9572 ( \9915 , \9907 , \9914 );
or \U$9573 ( \9916 , \9906 , \9915 );
nand \U$9574 ( \9917 , \9905 , \9895 );
nand \U$9575 ( \9918 , \9916 , \9917 );
not \U$9576 ( \9919 , \9918 );
not \U$9577 ( \9920 , \8445 );
and \U$9578 ( \9921 , RIbb2e440_39, \993 );
not \U$9579 ( \9922 , RIbb2e440_39);
and \U$9580 ( \9923 , \9922 , \7345 );
or \U$9581 ( \9924 , \9921 , \9923 );
not \U$9582 ( \9925 , \9924 );
or \U$9583 ( \9926 , \9920 , \9925 );
nand \U$9584 ( \9927 , \9443 , \8450 );
nand \U$9585 ( \9928 , \9926 , \9927 );
not \U$9586 ( \9929 , \9928 );
not \U$9587 ( \9930 , \3887 );
not \U$9588 ( \9931 , RIbb2e710_33);
not \U$9589 ( \9932 , \1688 );
or \U$9590 ( \9933 , \9931 , \9932 );
not \U$9591 ( \9934 , \3370 );
nand \U$9592 ( \9935 , \9934 , \2935 );
nand \U$9593 ( \9936 , \9933 , \9935 );
not \U$9594 ( \9937 , \9936 );
or \U$9595 ( \9938 , \9930 , \9937 );
nand \U$9596 ( \9939 , \9453 , \4791 );
nand \U$9597 ( \9940 , \9938 , \9939 );
not \U$9598 ( \9941 , \9940 );
or \U$9599 ( \9942 , \9929 , \9941 );
or \U$9600 ( \9943 , \9928 , \9940 );
not \U$9601 ( \9944 , \2078 );
not \U$9602 ( \9945 , \9183 );
or \U$9603 ( \9946 , \9944 , \9945 );
not \U$9604 ( \9947 , RIbb2ecb0_21);
not \U$9605 ( \9948 , \3342 );
or \U$9606 ( \9949 , \9947 , \9948 );
nand \U$9607 ( \9950 , \3521 , \2249 );
nand \U$9608 ( \9951 , \9949 , \9950 );
nand \U$9609 ( \9952 , \9951 , \2077 );
nand \U$9610 ( \9953 , \9946 , \9952 );
nand \U$9611 ( \9954 , \9943 , \9953 );
nand \U$9612 ( \9955 , \9942 , \9954 );
not \U$9613 ( \9956 , \9955 );
or \U$9614 ( \9957 , \9919 , \9956 );
or \U$9615 ( \9958 , \9955 , \9918 );
and \U$9616 ( \9959 , \9372 , \5845 );
not \U$9617 ( \9960 , RIbb2e620_35);
not \U$9618 ( \9961 , \4299 );
or \U$9619 ( \9962 , \9960 , \9961 );
nand \U$9620 ( \9963 , \1548 , \6002 );
nand \U$9621 ( \9964 , \9962 , \9963 );
and \U$9622 ( \9965 , \9964 , \4712 );
nor \U$9623 ( \9966 , \9959 , \9965 );
not \U$9624 ( \9967 , \9966 );
not \U$9625 ( \9968 , \9967 );
xor \U$9626 ( \9969 , RIbb2ead0_25, \1339 );
and \U$9627 ( \9970 , \9969 , \2980 );
and \U$9628 ( \9971 , \9388 , \2963 );
nor \U$9629 ( \9972 , \9970 , \9971 );
not \U$9630 ( \9973 , \9972 );
not \U$9631 ( \9974 , \9973 );
or \U$9632 ( \9975 , \9968 , \9974 );
not \U$9633 ( \9976 , \9966 );
not \U$9634 ( \9977 , \9972 );
or \U$9635 ( \9978 , \9976 , \9977 );
not \U$9636 ( \9979 , \3407 );
not \U$9637 ( \9980 , RIbb2ebc0_23);
not \U$9638 ( \9981 , \3563 );
or \U$9639 ( \9982 , \9980 , \9981 );
not \U$9640 ( \9983 , \2114 );
not \U$9641 ( \9984 , \9983 );
nand \U$9642 ( \9985 , \9984 , \3396 );
nand \U$9643 ( \9986 , \9982 , \9985 );
not \U$9644 ( \9987 , \9986 );
or \U$9645 ( \9988 , \9979 , \9987 );
nand \U$9646 ( \9989 , \9464 , \3383 );
nand \U$9647 ( \9990 , \9988 , \9989 );
nand \U$9648 ( \9991 , \9978 , \9990 );
nand \U$9649 ( \9992 , \9975 , \9991 );
nand \U$9650 ( \9993 , \9958 , \9992 );
nand \U$9651 ( \9994 , \9957 , \9993 );
xor \U$9652 ( \9995 , \9885 , \9994 );
not \U$9653 ( \9996 , \9471 );
not \U$9654 ( \9997 , \9396 );
or \U$9655 ( \9998 , \9996 , \9997 );
or \U$9656 ( \9999 , \9471 , \9396 );
nand \U$9657 ( \10000 , \9998 , \9999 );
xor \U$9658 ( \10001 , \9435 , \10000 );
and \U$9659 ( \10002 , \9995 , \10001 );
and \U$9660 ( \10003 , \9885 , \9994 );
or \U$9661 ( \10004 , \10002 , \10003 );
nand \U$9662 ( \10005 , \9788 , \10004 );
nand \U$9663 ( \10006 , \9784 , \10005 );
xor \U$9664 ( \10007 , \9776 , \10006 );
xor \U$9665 ( \10008 , \9258 , \9478 );
xor \U$9666 ( \10009 , \10008 , \9481 );
xnor \U$9667 ( \10010 , \10007 , \10009 );
xor \U$9668 ( \10011 , \9677 , \9685 );
xor \U$9669 ( \10012 , \10011 , \9773 );
not \U$9670 ( \10013 , \10012 );
xor \U$9671 ( \10014 , \9385 , \9374 );
buf \U$9672 ( \10015 , \9392 );
not \U$9673 ( \10016 , \10015 );
and \U$9674 ( \10017 , \10014 , \10016 );
not \U$9675 ( \10018 , \10014 );
and \U$9676 ( \10019 , \10018 , \10015 );
nor \U$9677 ( \10020 , \10017 , \10019 );
not \U$9678 ( \10021 , \10020 );
xor \U$9679 ( \10022 , \9323 , \9333 );
xor \U$9680 ( \10023 , \10022 , \9343 );
not \U$9681 ( \10024 , \10023 );
not \U$9682 ( \10025 , \10024 );
or \U$9683 ( \10026 , \10021 , \10025 );
xor \U$9684 ( \10027 , \9281 , \9294 );
xor \U$9685 ( \10028 , \10027 , \9307 );
not \U$9686 ( \10029 , \10028 );
nand \U$9687 ( \10030 , \10026 , \10029 );
not \U$9688 ( \10031 , \10020 );
nand \U$9689 ( \10032 , \10031 , \10023 );
nand \U$9690 ( \10033 , \10030 , \10032 );
xor \U$9691 ( \10034 , \9309 , \9260 );
xor \U$9692 ( \10035 , \10034 , \9262 );
xor \U$9693 ( \10036 , \10033 , \10035 );
and \U$9694 ( \10037 , \9468 , \9457 );
not \U$9695 ( \10038 , \9468 );
not \U$9696 ( \10039 , \9457 );
and \U$9697 ( \10040 , \10038 , \10039 );
nor \U$9698 ( \10041 , \10037 , \10040 );
xor \U$9699 ( \10042 , \9447 , \10041 );
xor \U$9700 ( \10043 , \9408 , \9433 );
xor \U$9701 ( \10044 , \10043 , \9419 );
xor \U$9702 ( \10045 , \10042 , \10044 );
not \U$9703 ( \10046 , \9200 );
not \U$9704 ( \10047 , \9188 );
or \U$9705 ( \10048 , \10046 , \10047 );
or \U$9706 ( \10049 , \9188 , \9200 );
nand \U$9707 ( \10050 , \10048 , \10049 );
and \U$9708 ( \10051 , \10050 , \9175 );
not \U$9709 ( \10052 , \10050 );
and \U$9710 ( \10053 , \10052 , \9176 );
nor \U$9711 ( \10054 , \10051 , \10053 );
and \U$9712 ( \10055 , \10045 , \10054 );
and \U$9713 ( \10056 , \10042 , \10044 );
or \U$9714 ( \10057 , \10055 , \10056 );
and \U$9715 ( \10058 , \10036 , \10057 );
and \U$9716 ( \10059 , \10033 , \10035 );
or \U$9717 ( \10060 , \10058 , \10059 );
not \U$9718 ( \10061 , \10060 );
not \U$9719 ( \10062 , \9219 );
not \U$9720 ( \10063 , \10062 );
not \U$9721 ( \10064 , \9216 );
or \U$9722 ( \10065 , \10063 , \10064 );
nand \U$9723 ( \10066 , \9215 , \9219 );
nand \U$9724 ( \10067 , \10065 , \10066 );
not \U$9725 ( \10068 , \9213 );
and \U$9726 ( \10069 , \10067 , \10068 );
not \U$9727 ( \10070 , \10067 );
and \U$9728 ( \10071 , \10070 , \9213 );
nor \U$9729 ( \10072 , \10069 , \10071 );
nand \U$9730 ( \10073 , \10061 , \10072 );
not \U$9731 ( \10074 , \10073 );
or \U$9732 ( \10075 , \10013 , \10074 );
not \U$9733 ( \10076 , \10072 );
buf \U$9734 ( \10077 , \10060 );
nand \U$9735 ( \10078 , \10076 , \10077 );
nand \U$9736 ( \10079 , \10075 , \10078 );
not \U$9737 ( \10080 , \10079 );
xor \U$9738 ( \10081 , \9222 , \9160 );
not \U$9739 ( \10082 , \9157 );
and \U$9740 ( \10083 , \10081 , \10082 );
not \U$9741 ( \10084 , \10081 );
and \U$9742 ( \10085 , \10084 , \9157 );
nor \U$9743 ( \10086 , \10083 , \10085 );
not \U$9744 ( \10087 , \10086 );
and \U$9745 ( \10088 , \10080 , \10087 );
not \U$9746 ( \10089 , \10080 );
and \U$9747 ( \10090 , \10089 , \10086 );
nor \U$9748 ( \10091 , \10088 , \10090 );
not \U$9749 ( \10092 , \10091 );
not \U$9750 ( \10093 , \9323 );
not \U$9751 ( \10094 , \1445 );
not \U$9752 ( \10095 , \3021 );
not \U$9753 ( \10096 , \10095 );
and \U$9754 ( \10097 , RIbb2ef80_15, \10096 );
not \U$9755 ( \10098 , RIbb2ef80_15);
and \U$9756 ( \10099 , \10098 , \10095 );
or \U$9757 ( \10100 , \10097 , \10099 );
not \U$9758 ( \10101 , \10100 );
or \U$9759 ( \10102 , \10094 , \10101 );
nand \U$9760 ( \10103 , \9339 , \1517 );
nand \U$9761 ( \10104 , \10102 , \10103 );
xor \U$9762 ( \10105 , \10093 , \10104 );
and \U$9763 ( \10106 , RIbb2e0f8_46, RIbb2e170_45);
not \U$9764 ( \10107 , RIbb2e0f8_46);
and \U$9765 ( \10108 , \10107 , \9094 );
nor \U$9766 ( \10109 , \10106 , \10108 );
not \U$9767 ( \10110 , \10109 );
and \U$9768 ( \10111 , RIbb2e0f8_46, RIbb2e080_47);
not \U$9769 ( \10112 , RIbb2e0f8_46);
not \U$9770 ( \10113 , RIbb2e080_47);
and \U$9771 ( \10114 , \10112 , \10113 );
nor \U$9772 ( \10115 , \10111 , \10114 );
nor \U$9773 ( \10116 , \10110 , \10115 );
buf \U$9774 ( \10117 , \10116 );
buf \U$9775 ( \10118 , \10115 );
buf \U$9776 ( \10119 , \10118 );
or \U$9777 ( \10120 , \10117 , \10119 );
nand \U$9778 ( \10121 , \10120 , RIbb2e170_45);
not \U$9779 ( \10122 , \1570 );
not \U$9780 ( \10123 , \9319 );
or \U$9781 ( \10124 , \10122 , \10123 );
not \U$9782 ( \10125 , RIbb2f250_9);
not \U$9783 ( \10126 , \7111 );
not \U$9784 ( \10127 , \10126 );
or \U$9785 ( \10128 , \10125 , \10127 );
nand \U$9786 ( \10129 , \6232 , \1554 );
nand \U$9787 ( \10130 , \10128 , \10129 );
nand \U$9788 ( \10131 , \1533 , \10130 );
nand \U$9789 ( \10132 , \10124 , \10131 );
xor \U$9790 ( \10133 , \10121 , \10132 );
not \U$9791 ( \10134 , \1077 );
not \U$9792 ( \10135 , \9739 );
or \U$9793 ( \10136 , \10134 , \10135 );
and \U$9794 ( \10137 , RIbb2f160_11, \6268 );
not \U$9795 ( \10138 , RIbb2f160_11);
and \U$9796 ( \10139 , \10138 , \4394 );
nor \U$9797 ( \10140 , \10137 , \10139 );
not \U$9798 ( \10141 , \10140 );
nand \U$9799 ( \10142 , \10141 , \1011 );
nand \U$9800 ( \10143 , \10136 , \10142 );
and \U$9801 ( \10144 , \10133 , \10143 );
and \U$9802 ( \10145 , \10121 , \10132 );
or \U$9803 ( \10146 , \10144 , \10145 );
and \U$9804 ( \10147 , \10105 , \10146 );
and \U$9805 ( \10148 , \10093 , \10104 );
or \U$9806 ( \10149 , \10147 , \10148 );
not \U$9807 ( \10150 , \1737 );
not \U$9808 ( \10151 , \9805 );
or \U$9809 ( \10152 , \10150 , \10151 );
not \U$9810 ( \10153 , RIbb2f340_7);
not \U$9811 ( \10154 , \8338 );
or \U$9812 ( \10155 , \10153 , \10154 );
buf \U$9813 ( \10156 , \9056 );
nand \U$9814 ( \10157 , \10156 , \2700 );
nand \U$9815 ( \10158 , \10155 , \10157 );
nand \U$9816 ( \10159 , \10158 , \1702 );
nand \U$9817 ( \10160 , \10152 , \10159 );
not \U$9818 ( \10161 , \1147 );
not \U$9819 ( \10162 , \9795 );
or \U$9820 ( \10163 , \10161 , \10162 );
not \U$9821 ( \10164 , RIbb2f430_5);
not \U$9822 ( \10165 , \7300 );
not \U$9823 ( \10166 , \10165 );
or \U$9824 ( \10167 , \10164 , \10166 );
nand \U$9825 ( \10168 , \7300 , \1980 );
nand \U$9826 ( \10169 , \10167 , \10168 );
nand \U$9827 ( \10170 , \10169 , \1090 );
nand \U$9828 ( \10171 , \10163 , \10170 );
xor \U$9829 ( \10172 , \10160 , \10171 );
not \U$9830 ( \10173 , \1265 );
not \U$9831 ( \10174 , \1246 );
not \U$9832 ( \10175 , \8630 );
not \U$9833 ( \10176 , \10175 );
or \U$9834 ( \10177 , \10174 , \10176 );
not \U$9835 ( \10178 , \10175 );
nand \U$9836 ( \10179 , \10178 , \1245 );
nand \U$9837 ( \10180 , \10177 , \10179 );
not \U$9838 ( \10181 , \10180 );
or \U$9839 ( \10182 , \10173 , \10181 );
not \U$9840 ( \10183 , \9821 );
nand \U$9841 ( \10184 , \10183 , \1294 );
nand \U$9842 ( \10185 , \10182 , \10184 );
and \U$9843 ( \10186 , \10172 , \10185 );
and \U$9844 ( \10187 , \10160 , \10171 );
or \U$9845 ( \10188 , \10186 , \10187 );
not \U$9846 ( \10189 , \10188 );
xor \U$9847 ( \10190 , \9842 , \9854 );
xor \U$9848 ( \10191 , \10190 , \9865 );
nand \U$9849 ( \10192 , \10189 , \10191 );
not \U$9850 ( \10193 , \10192 );
not \U$9851 ( \10194 , \3887 );
not \U$9852 ( \10195 , RIbb2e710_33);
not \U$9853 ( \10196 , \3773 );
or \U$9854 ( \10197 , \10195 , \10196 );
nand \U$9855 ( \10198 , \3243 , \3877 );
nand \U$9856 ( \10199 , \10197 , \10198 );
not \U$9857 ( \10200 , \10199 );
or \U$9858 ( \10201 , \10194 , \10200 );
nand \U$9859 ( \10202 , \9936 , \4791 );
nand \U$9860 ( \10203 , \10201 , \10202 );
not \U$9861 ( \10204 , \836 );
not \U$9862 ( \10205 , \9722 );
or \U$9863 ( \10206 , \10204 , \10205 );
not \U$9864 ( \10207 , RIbb2ee90_17);
not \U$9865 ( \10208 , \3655 );
or \U$9866 ( \10209 , \10207 , \10208 );
nand \U$9867 ( \10210 , \7021 , \3057 );
nand \U$9868 ( \10211 , \10209 , \10210 );
nand \U$9869 ( \10212 , \10211 , \832 );
nand \U$9870 ( \10213 , \10206 , \10212 );
xor \U$9871 ( \10214 , \10203 , \10213 );
not \U$9872 ( \10215 , \855 );
not \U$9873 ( \10216 , \9709 );
or \U$9874 ( \10217 , \10215 , \10216 );
not \U$9875 ( \10218 , RIbb2eda0_19);
not \U$9876 ( \10219 , \3203 );
or \U$9877 ( \10220 , \10218 , \10219 );
nand \U$9878 ( \10221 , \3202 , \1776 );
nand \U$9879 ( \10222 , \10220 , \10221 );
nand \U$9880 ( \10223 , \10222 , \853 );
nand \U$9881 ( \10224 , \10217 , \10223 );
and \U$9882 ( \10225 , \10214 , \10224 );
and \U$9883 ( \10226 , \10203 , \10213 );
or \U$9884 ( \10227 , \10225 , \10226 );
not \U$9885 ( \10228 , \10227 );
or \U$9886 ( \10229 , \10193 , \10228 );
not \U$9887 ( \10230 , \10191 );
nand \U$9888 ( \10231 , \10230 , \10188 );
nand \U$9889 ( \10232 , \10229 , \10231 );
xor \U$9890 ( \10233 , \10149 , \10232 );
xor \U$9891 ( \10234 , \9809 , \9799 );
not \U$9892 ( \10235 , \9826 );
and \U$9893 ( \10236 , \10234 , \10235 );
not \U$9894 ( \10237 , \10234 );
and \U$9895 ( \10238 , \10237 , \9826 );
nor \U$9896 ( \10239 , \10236 , \10238 );
not \U$9897 ( \10240 , \10239 );
not \U$9898 ( \10241 , \5845 );
not \U$9899 ( \10242 , \9964 );
or \U$9900 ( \10243 , \10241 , \10242 );
not \U$9901 ( \10244 , RIbb2e620_35);
not \U$9902 ( \10245 , \3479 );
or \U$9903 ( \10246 , \10244 , \10245 );
nand \U$9904 ( \10247 , \3480 , \6002 );
nand \U$9905 ( \10248 , \10246 , \10247 );
nand \U$9906 ( \10249 , \10248 , \4712 );
nand \U$9907 ( \10250 , \10243 , \10249 );
not \U$9908 ( \10251 , \10250 );
not \U$9909 ( \10252 , \3406 );
not \U$9910 ( \10253 , RIbb2ebc0_23);
not \U$9911 ( \10254 , \2224 );
or \U$9912 ( \10255 , \10253 , \10254 );
nand \U$9913 ( \10256 , \3320 , \3396 );
nand \U$9914 ( \10257 , \10255 , \10256 );
not \U$9915 ( \10258 , \10257 );
or \U$9916 ( \10259 , \10252 , \10258 );
nand \U$9917 ( \10260 , \9986 , \3383 );
nand \U$9918 ( \10261 , \10259 , \10260 );
not \U$9919 ( \10262 , \10261 );
nand \U$9920 ( \10263 , \10251 , \10262 );
not \U$9921 ( \10264 , \10263 );
not \U$9922 ( \10265 , \2078 );
not \U$9923 ( \10266 , \9951 );
or \U$9924 ( \10267 , \10265 , \10266 );
not \U$9925 ( \10268 , RIbb2ecb0_21);
not \U$9926 ( \10269 , \3168 );
or \U$9927 ( \10270 , \10268 , \10269 );
nand \U$9928 ( \10271 , \3167 , \849 );
nand \U$9929 ( \10272 , \10270 , \10271 );
nand \U$9930 ( \10273 , \10272 , \2077 );
nand \U$9931 ( \10274 , \10267 , \10273 );
not \U$9932 ( \10275 , \10274 );
or \U$9933 ( \10276 , \10264 , \10275 );
nand \U$9934 ( \10277 , \10250 , \10261 );
nand \U$9935 ( \10278 , \10276 , \10277 );
not \U$9936 ( \10279 , \10278 );
or \U$9937 ( \10280 , \10240 , \10279 );
or \U$9938 ( \10281 , \10278 , \10239 );
not \U$9939 ( \10282 , \3613 );
not \U$9940 ( \10283 , \9697 );
or \U$9941 ( \10284 , \10282 , \10283 );
not \U$9942 ( \10285 , RIbb2e800_31);
not \U$9943 ( \10286 , \1113 );
or \U$9944 ( \10287 , \10285 , \10286 );
not \U$9945 ( \10288 , \4766 );
nand \U$9946 ( \10289 , \10288 , \2917 );
nand \U$9947 ( \10290 , \10287 , \10289 );
nand \U$9948 ( \10291 , \10290 , \2940 );
nand \U$9949 ( \10292 , \10284 , \10291 );
not \U$9950 ( \10293 , \8608 );
not \U$9951 ( \10294 , \10293 );
not \U$9952 ( \10295 , \4360 );
or \U$9953 ( \10296 , \10294 , \10295 );
nand \U$9954 ( \10297 , \10296 , \4364 );
nand \U$9955 ( \10298 , \601 , \647 );
xnor \U$9956 ( \10299 , \10297 , \10298 );
buf \U$9957 ( \10300 , \10299 );
buf \U$9958 ( \10301 , \10300 );
and \U$9959 ( \10302 , \1313 , \10301 );
or \U$9960 ( \10303 , \10292 , \10302 );
not \U$9961 ( \10304 , \1429 );
not \U$9962 ( \10305 , \1313 );
not \U$9963 ( \10306 , \9841 );
not \U$9964 ( \10307 , \10306 );
or \U$9965 ( \10308 , \10305 , \10307 );
nand \U$9966 ( \10309 , \9841 , \1951 );
nand \U$9967 ( \10310 , \10308 , \10309 );
not \U$9968 ( \10311 , \10310 );
or \U$9969 ( \10312 , \10304 , \10311 );
nand \U$9970 ( \10313 , \9862 , \1376 );
nand \U$9971 ( \10314 , \10312 , \10313 );
nand \U$9972 ( \10315 , \10303 , \10314 );
nand \U$9973 ( \10316 , \10292 , \10302 );
nand \U$9974 ( \10317 , \10315 , \10316 );
nand \U$9975 ( \10318 , \10281 , \10317 );
nand \U$9976 ( \10319 , \10280 , \10318 );
and \U$9977 ( \10320 , \10233 , \10319 );
and \U$9978 ( \10321 , \10149 , \10232 );
or \U$9979 ( \10322 , \10320 , \10321 );
not \U$9980 ( \10323 , \10322 );
xor \U$9981 ( \10324 , \9203 , \9206 );
xnor \U$9982 ( \10325 , \10324 , \9211 );
not \U$9983 ( \10326 , \9359 );
not \U$9984 ( \10327 , \9346 );
not \U$9985 ( \10328 , \10327 );
or \U$9986 ( \10329 , \10326 , \10328 );
nand \U$9987 ( \10330 , \9358 , \9346 );
nand \U$9988 ( \10331 , \10329 , \10330 );
buf \U$9989 ( \10332 , \9349 );
not \U$9990 ( \10333 , \10332 );
and \U$9991 ( \10334 , \10331 , \10333 );
not \U$9992 ( \10335 , \10331 );
and \U$9993 ( \10336 , \10335 , \10332 );
nor \U$9994 ( \10337 , \10334 , \10336 );
nand \U$9995 ( \10338 , \10325 , \10337 );
not \U$9996 ( \10339 , \10338 );
or \U$9997 ( \10340 , \10323 , \10339 );
not \U$9998 ( \10341 , \10325 );
not \U$9999 ( \10342 , \10337 );
nand \U$10000 ( \10343 , \10341 , \10342 );
nand \U$10001 ( \10344 , \10340 , \10343 );
not \U$10002 ( \10345 , \10344 );
xor \U$10003 ( \10346 , \9778 , \10004 );
xor \U$10004 ( \10347 , \10346 , \9781 );
buf \U$10005 ( \10348 , \10347 );
not \U$10006 ( \10349 , \10348 );
not \U$10007 ( \10350 , \10349 );
or \U$10008 ( \10351 , \10345 , \10350 );
not \U$10009 ( \10352 , \10344 );
not \U$10010 ( \10353 , \10352 );
not \U$10011 ( \10354 , \10348 );
or \U$10012 ( \10355 , \10353 , \10354 );
xor \U$10013 ( \10356 , \9885 , \9994 );
xor \U$10014 ( \10357 , \10356 , \10001 );
not \U$10015 ( \10358 , \9869 );
not \U$10016 ( \10359 , \9828 );
or \U$10017 ( \10360 , \10358 , \10359 );
nand \U$10018 ( \10361 , \9829 , \9868 );
nand \U$10019 ( \10362 , \10360 , \10361 );
and \U$10020 ( \10363 , \10362 , \9883 );
not \U$10021 ( \10364 , \10362 );
not \U$10022 ( \10365 , \9883 );
and \U$10023 ( \10366 , \10364 , \10365 );
nor \U$10024 ( \10367 , \10363 , \10366 );
not \U$10025 ( \10368 , \10367 );
not \U$10026 ( \10369 , \10368 );
not \U$10027 ( \10370 , \8362 );
not \U$10028 ( \10371 , RIbb2e350_41);
not \U$10029 ( \10372 , \3452 );
or \U$10030 ( \10373 , \10371 , \10372 );
nand \U$10031 ( \10374 , \4558 , \8357 );
nand \U$10032 ( \10375 , \10373 , \10374 );
not \U$10033 ( \10376 , \10375 );
or \U$10034 ( \10377 , \10370 , \10376 );
nand \U$10035 ( \10378 , \9903 , \8995 );
nand \U$10036 ( \10379 , \10377 , \10378 );
not \U$10037 ( \10380 , \10379 );
not \U$10038 ( \10381 , \2963 );
not \U$10039 ( \10382 , \9969 );
or \U$10040 ( \10383 , \10381 , \10382 );
and \U$10041 ( \10384 , RIbb2ead0_25, \3807 );
not \U$10042 ( \10385 , RIbb2ead0_25);
and \U$10043 ( \10386 , \10385 , \3810 );
or \U$10044 ( \10387 , \10384 , \10386 );
nand \U$10045 ( \10388 , \10387 , \2980 );
nand \U$10046 ( \10389 , \10383 , \10388 );
not \U$10047 ( \10390 , \10389 );
or \U$10048 ( \10391 , \10380 , \10390 );
or \U$10049 ( \10392 , \10389 , \10379 );
not \U$10050 ( \10393 , \6251 );
not \U$10051 ( \10394 , RIbb2e530_37);
not \U$10052 ( \10395 , \4595 );
or \U$10053 ( \10396 , \10394 , \10395 );
nand \U$10054 ( \10397 , \1563 , \8701 );
nand \U$10055 ( \10398 , \10396 , \10397 );
not \U$10056 ( \10399 , \10398 );
or \U$10057 ( \10400 , \10393 , \10399 );
nand \U$10058 ( \10401 , \9893 , \6242 );
nand \U$10059 ( \10402 , \10400 , \10401 );
nand \U$10060 ( \10403 , \10392 , \10402 );
nand \U$10061 ( \10404 , \10391 , \10403 );
not \U$10062 ( \10405 , \2925 );
not \U$10063 ( \10406 , \9747 );
or \U$10064 ( \10407 , \10405 , \10406 );
not \U$10065 ( \10408 , \3800 );
not \U$10066 ( \10409 , \3109 );
or \U$10067 ( \10410 , \10408 , \10409 );
not \U$10068 ( \10411 , \3736 );
nand \U$10069 ( \10412 , \10411 , RIbb2e8f0_29);
nand \U$10070 ( \10413 , \10410 , \10412 );
nand \U$10071 ( \10414 , \10413 , \2922 );
nand \U$10072 ( \10415 , \10407 , \10414 );
not \U$10073 ( \10416 , \10415 );
not \U$10074 ( \10417 , \8445 );
not \U$10075 ( \10418 , RIbb2e440_39);
not \U$10076 ( \10419 , \3981 );
or \U$10077 ( \10420 , \10418 , \10419 );
not \U$10078 ( \10421 , \956 );
or \U$10079 ( \10422 , \10421 , RIbb2e440_39);
nand \U$10080 ( \10423 , \10420 , \10422 );
not \U$10081 ( \10424 , \10423 );
or \U$10082 ( \10425 , \10417 , \10424 );
nand \U$10083 ( \10426 , \9924 , \8450 );
nand \U$10084 ( \10427 , \10425 , \10426 );
not \U$10085 ( \10428 , \10427 );
or \U$10086 ( \10429 , \10416 , \10428 );
or \U$10087 ( \10430 , \10427 , \10415 );
not \U$10088 ( \10431 , \3445 );
not \U$10089 ( \10432 , RIbb2e9e0_27);
not \U$10090 ( \10433 , \1420 );
or \U$10091 ( \10434 , \10432 , \10433 );
nand \U$10092 ( \10435 , \1422 , \3454 );
nand \U$10093 ( \10436 , \10434 , \10435 );
not \U$10094 ( \10437 , \10436 );
or \U$10095 ( \10438 , \10431 , \10437 );
nand \U$10096 ( \10439 , \9912 , \3465 );
nand \U$10097 ( \10440 , \10438 , \10439 );
nand \U$10098 ( \10441 , \10430 , \10440 );
nand \U$10099 ( \10442 , \10429 , \10441 );
xor \U$10100 ( \10443 , \10404 , \10442 );
not \U$10101 ( \10444 , RIbb2e260_43);
and \U$10102 ( \10445 , \1580 , \10444 );
not \U$10103 ( \10446 , \1580 );
and \U$10104 ( \10447 , \10446 , RIbb2e260_43);
or \U$10105 ( \10448 , \10445 , \10447 );
buf \U$10106 ( \10449 , \9097 );
and \U$10107 ( \10450 , \10448 , \10449 );
buf \U$10108 ( \10451 , \9099 );
and \U$10109 ( \10452 , \9849 , \10451 );
nor \U$10110 ( \10453 , \10450 , \10452 );
not \U$10111 ( \10454 , \10453 );
not \U$10112 ( \10455 , RIbb2f070_13);
not \U$10113 ( \10456 , \4040 );
or \U$10114 ( \10457 , \10455 , \10456 );
buf \U$10115 ( \10458 , \3089 );
nand \U$10116 ( \10459 , \10458 , \3421 );
nand \U$10117 ( \10460 , \10457 , \10459 );
and \U$10118 ( \10461 , \10460 , \916 );
and \U$10119 ( \10462 , \9759 , \998 );
nor \U$10120 ( \10463 , \10461 , \10462 );
not \U$10121 ( \10464 , \10463 );
or \U$10122 ( \10465 , \10454 , \10464 );
not \U$10123 ( \10466 , \1445 );
and \U$10124 ( \10467 , RIbb2ef80_15, \4031 );
not \U$10125 ( \10468 , RIbb2ef80_15);
and \U$10126 ( \10469 , \10468 , \4030 );
or \U$10127 ( \10470 , \10467 , \10469 );
not \U$10128 ( \10471 , \10470 );
or \U$10129 ( \10472 , \10466 , \10471 );
nand \U$10130 ( \10473 , \10100 , \1517 );
nand \U$10131 ( \10474 , \10472 , \10473 );
nand \U$10132 ( \10475 , \10465 , \10474 );
not \U$10133 ( \10476 , \10463 );
not \U$10134 ( \10477 , \10453 );
nand \U$10135 ( \10478 , \10476 , \10477 );
nand \U$10136 ( \10479 , \10475 , \10478 );
and \U$10137 ( \10480 , \10443 , \10479 );
and \U$10138 ( \10481 , \10404 , \10442 );
or \U$10139 ( \10482 , \10480 , \10481 );
not \U$10140 ( \10483 , \10482 );
not \U$10141 ( \10484 , \10483 );
or \U$10142 ( \10485 , \10369 , \10484 );
xor \U$10143 ( \10486 , \9905 , \9895 );
and \U$10144 ( \10487 , \10486 , \9915 );
not \U$10145 ( \10488 , \10486 );
not \U$10146 ( \10489 , \9915 );
and \U$10147 ( \10490 , \10488 , \10489 );
nor \U$10148 ( \10491 , \10487 , \10490 );
not \U$10149 ( \10492 , \10491 );
xor \U$10150 ( \10493 , \9953 , \9940 );
xnor \U$10151 ( \10494 , \10493 , \9928 );
not \U$10152 ( \10495 , \10494 );
or \U$10153 ( \10496 , \10492 , \10495 );
xor \U$10154 ( \10497 , \9726 , \9713 );
xor \U$10155 ( \10498 , \10497 , \9701 );
nand \U$10156 ( \10499 , \10496 , \10498 );
not \U$10157 ( \10500 , \10494 );
not \U$10158 ( \10501 , \10491 );
nand \U$10159 ( \10502 , \10500 , \10501 );
nand \U$10160 ( \10503 , \10499 , \10502 );
nand \U$10161 ( \10504 , \10485 , \10503 );
nand \U$10162 ( \10505 , \10482 , \10367 );
nand \U$10163 ( \10506 , \10504 , \10505 );
or \U$10164 ( \10507 , \10357 , \10506 );
xor \U$10165 ( \10508 , \9688 , \9690 );
xor \U$10166 ( \10509 , \10508 , \9770 );
nand \U$10167 ( \10510 , \10507 , \10509 );
nand \U$10168 ( \10511 , \10506 , \10357 );
nand \U$10169 ( \10512 , \10510 , \10511 );
nand \U$10170 ( \10513 , \10355 , \10512 );
nand \U$10171 ( \10514 , \10351 , \10513 );
not \U$10172 ( \10515 , \10514 );
and \U$10173 ( \10516 , \10092 , \10515 );
and \U$10174 ( \10517 , \10091 , \10514 );
nor \U$10175 ( \10518 , \10516 , \10517 );
xor \U$10176 ( \10519 , \10010 , \10518 );
xor \U$10177 ( \10520 , \10033 , \10035 );
xor \U$10178 ( \10521 , \10520 , \10057 );
xor \U$10179 ( \10522 , \9992 , \9955 );
xnor \U$10180 ( \10523 , \10522 , \9918 );
not \U$10181 ( \10524 , \10523 );
not \U$10182 ( \10525 , \10524 );
xor \U$10183 ( \10526 , \9730 , \9728 );
xnor \U$10184 ( \10527 , \10526 , \9766 );
not \U$10185 ( \10528 , \10527 );
not \U$10186 ( \10529 , \10528 );
or \U$10187 ( \10530 , \10525 , \10529 );
not \U$10188 ( \10531 , \10523 );
not \U$10189 ( \10532 , \10527 );
or \U$10190 ( \10533 , \10531 , \10532 );
xor \U$10191 ( \10534 , \9741 , \9751 );
xor \U$10192 ( \10535 , \10534 , \9763 );
not \U$10193 ( \10536 , \10535 );
and \U$10194 ( \10537 , \9990 , \9972 );
not \U$10195 ( \10538 , \9990 );
and \U$10196 ( \10539 , \10538 , \9973 );
or \U$10197 ( \10540 , \10537 , \10539 );
and \U$10198 ( \10541 , \10540 , \9967 );
not \U$10199 ( \10542 , \10540 );
and \U$10200 ( \10543 , \10542 , \9966 );
nor \U$10201 ( \10544 , \10541 , \10543 );
not \U$10202 ( \10545 , \10544 );
or \U$10203 ( \10546 , \10536 , \10545 );
or \U$10204 ( \10547 , \10544 , \10535 );
not \U$10205 ( \10548 , \10140 );
not \U$10206 ( \10549 , \1943 );
and \U$10207 ( \10550 , \10548 , \10549 );
not \U$10208 ( \10551 , RIbb2f160_11);
not \U$10209 ( \10552 , \6202 );
not \U$10210 ( \10553 , \10552 );
or \U$10211 ( \10554 , \10551 , \10553 );
buf \U$10212 ( \10555 , \4696 );
buf \U$10213 ( \10556 , \10555 );
not \U$10214 ( \10557 , \10556 );
nand \U$10215 ( \10558 , \10557 , \1048 );
nand \U$10216 ( \10559 , \10554 , \10558 );
and \U$10217 ( \10560 , \10559 , \1011 );
nor \U$10218 ( \10561 , \10550 , \10560 );
not \U$10219 ( \10562 , \10561 );
not \U$10220 ( \10563 , \1702 );
not \U$10221 ( \10564 , RIbb2f340_7);
not \U$10222 ( \10565 , \8639 );
or \U$10223 ( \10566 , \10564 , \10565 );
nand \U$10224 ( \10567 , \6939 , \1692 );
nand \U$10225 ( \10568 , \10566 , \10567 );
not \U$10226 ( \10569 , \10568 );
or \U$10227 ( \10570 , \10563 , \10569 );
nand \U$10228 ( \10571 , \10158 , \1737 );
nand \U$10229 ( \10572 , \10570 , \10571 );
not \U$10230 ( \10573 , \1570 );
not \U$10231 ( \10574 , \10130 );
or \U$10232 ( \10575 , \10573 , \10574 );
not \U$10233 ( \10576 , RIbb2f250_9);
not \U$10234 ( \10577 , \7308 );
not \U$10235 ( \10578 , \10577 );
or \U$10236 ( \10579 , \10576 , \10578 );
nand \U$10237 ( \10580 , \5955 , \5064 );
nand \U$10238 ( \10581 , \10579 , \10580 );
nand \U$10239 ( \10582 , \10581 , \1533 );
nand \U$10240 ( \10583 , \10575 , \10582 );
xor \U$10241 ( \10584 , \10572 , \10583 );
not \U$10242 ( \10585 , \1090 );
not \U$10243 ( \10586 , RIbb2f430_5);
not \U$10244 ( \10587 , \8320 );
or \U$10245 ( \10588 , \10586 , \10587 );
nand \U$10246 ( \10589 , \9819 , \1898 );
nand \U$10247 ( \10590 , \10588 , \10589 );
not \U$10248 ( \10591 , \10590 );
or \U$10249 ( \10592 , \10585 , \10591 );
nand \U$10250 ( \10593 , \10169 , \1147 );
nand \U$10251 ( \10594 , \10592 , \10593 );
and \U$10252 ( \10595 , \10584 , \10594 );
and \U$10253 ( \10596 , \10572 , \10583 );
or \U$10254 ( \10597 , \10595 , \10596 );
xor \U$10255 ( \10598 , \10562 , \10597 );
buf \U$10256 ( \10599 , \10117 );
not \U$10257 ( \10600 , \10599 );
not \U$10258 ( \10601 , RIbb2e170_45);
not \U$10259 ( \10602 , \813 );
or \U$10260 ( \10603 , \10601 , \10602 );
not \U$10261 ( \10604 , \813 );
nand \U$10262 ( \10605 , \10604 , \9094 );
nand \U$10263 ( \10606 , \10603 , \10605 );
not \U$10264 ( \10607 , \10606 );
or \U$10265 ( \10608 , \10600 , \10607 );
nand \U$10266 ( \10609 , \10119 , RIbb2e170_45);
nand \U$10267 ( \10610 , \10608 , \10609 );
not \U$10268 ( \10611 , \1376 );
not \U$10269 ( \10612 , \10310 );
or \U$10270 ( \10613 , \10611 , \10612 );
xor \U$10271 ( \10614 , \1313 , \10301 );
nand \U$10272 ( \10615 , \10614 , \1429 );
nand \U$10273 ( \10616 , \10613 , \10615 );
xor \U$10274 ( \10617 , \10610 , \10616 );
not \U$10275 ( \10618 , \1294 );
not \U$10276 ( \10619 , \10180 );
or \U$10277 ( \10620 , \10618 , \10619 );
not \U$10278 ( \10621 , \1290 );
not \U$10279 ( \10622 , \9279 );
or \U$10280 ( \10623 , \10621 , \10622 );
nand \U$10281 ( \10624 , \9280 , \1245 );
nand \U$10282 ( \10625 , \10623 , \10624 );
nand \U$10283 ( \10626 , \10625 , \1265 );
nand \U$10284 ( \10627 , \10620 , \10626 );
and \U$10285 ( \10628 , \10617 , \10627 );
and \U$10286 ( \10629 , \10610 , \10616 );
or \U$10287 ( \10630 , \10628 , \10629 );
and \U$10288 ( \10631 , \10598 , \10630 );
and \U$10289 ( \10632 , \10562 , \10597 );
or \U$10290 ( \10633 , \10631 , \10632 );
nand \U$10291 ( \10634 , \10547 , \10633 );
nand \U$10292 ( \10635 , \10546 , \10634 );
nand \U$10293 ( \10636 , \10533 , \10635 );
nand \U$10294 ( \10637 , \10530 , \10636 );
or \U$10295 ( \10638 , \10521 , \10637 );
not \U$10296 ( \10639 , \10029 );
not \U$10297 ( \10640 , \10024 );
or \U$10298 ( \10641 , \10639 , \10640 );
nand \U$10299 ( \10642 , \10023 , \10028 );
nand \U$10300 ( \10643 , \10641 , \10642 );
buf \U$10301 ( \10644 , \10020 );
not \U$10302 ( \10645 , \10644 );
and \U$10303 ( \10646 , \10643 , \10645 );
not \U$10304 ( \10647 , \10643 );
and \U$10305 ( \10648 , \10647 , \10644 );
nor \U$10306 ( \10649 , \10646 , \10648 );
xor \U$10307 ( \10650 , \10042 , \10044 );
xor \U$10308 ( \10651 , \10650 , \10054 );
xor \U$10309 ( \10652 , \10649 , \10651 );
xor \U$10310 ( \10653 , \10093 , \10104 );
xor \U$10311 ( \10654 , \10653 , \10146 );
not \U$10312 ( \10655 , \4712 );
not \U$10313 ( \10656 , RIbb2e620_35);
not \U$10314 ( \10657 , \1688 );
or \U$10315 ( \10658 , \10656 , \10657 );
nand \U$10316 ( \10659 , \3552 , \5840 );
nand \U$10317 ( \10660 , \10658 , \10659 );
not \U$10318 ( \10661 , \10660 );
or \U$10319 ( \10662 , \10655 , \10661 );
nand \U$10320 ( \10663 , \10248 , \5845 );
nand \U$10321 ( \10664 , \10662 , \10663 );
not \U$10322 ( \10665 , \10664 );
not \U$10323 ( \10666 , \10665 );
not \U$10324 ( \10667 , \4791 );
not \U$10325 ( \10668 , \10199 );
or \U$10326 ( \10669 , \10667 , \10668 );
not \U$10327 ( \10670 , RIbb2e710_33);
not \U$10328 ( \10671 , \7424 );
or \U$10329 ( \10672 , \10670 , \10671 );
not \U$10330 ( \10673 , \8862 );
nand \U$10331 ( \10674 , \10673 , \4785 );
nand \U$10332 ( \10675 , \10672 , \10674 );
nand \U$10333 ( \10676 , \10675 , \3887 );
nand \U$10334 ( \10677 , \10669 , \10676 );
not \U$10335 ( \10678 , \10677 );
not \U$10336 ( \10679 , \10678 );
or \U$10337 ( \10680 , \10666 , \10679 );
not \U$10338 ( \10681 , \2077 );
not \U$10339 ( \10682 , RIbb2ecb0_21);
not \U$10340 ( \10683 , \3143 );
or \U$10341 ( \10684 , \10682 , \10683 );
nand \U$10342 ( \10685 , \3146 , \2254 );
nand \U$10343 ( \10686 , \10684 , \10685 );
not \U$10344 ( \10687 , \10686 );
or \U$10345 ( \10688 , \10681 , \10687 );
nand \U$10346 ( \10689 , \10272 , \2078 );
nand \U$10347 ( \10690 , \10688 , \10689 );
nand \U$10348 ( \10691 , \10680 , \10690 );
nand \U$10349 ( \10692 , \10677 , \10664 );
nand \U$10350 ( \10693 , \10691 , \10692 );
not \U$10351 ( \10694 , \10693 );
xor \U$10352 ( \10695 , \10302 , \10314 );
xnor \U$10353 ( \10696 , \10695 , \10292 );
not \U$10354 ( \10697 , \10696 );
not \U$10355 ( \10698 , \10697 );
or \U$10356 ( \10699 , \10694 , \10698 );
not \U$10357 ( \10700 , \10696 );
not \U$10358 ( \10701 , \10693 );
not \U$10359 ( \10702 , \10701 );
or \U$10360 ( \10703 , \10700 , \10702 );
xor \U$10361 ( \10704 , \10160 , \10171 );
xor \U$10362 ( \10705 , \10704 , \10185 );
nand \U$10363 ( \10706 , \10703 , \10705 );
nand \U$10364 ( \10707 , \10699 , \10706 );
or \U$10365 ( \10708 , \10654 , \10707 );
not \U$10366 ( \10709 , \8995 );
not \U$10367 ( \10710 , \10375 );
or \U$10368 ( \10711 , \10709 , \10710 );
not \U$10369 ( \10712 , RIbb2e350_41);
not \U$10370 ( \10713 , \989 );
or \U$10371 ( \10714 , \10712 , \10713 );
nand \U$10372 ( \10715 , \7345 , \7097 );
nand \U$10373 ( \10716 , \10714 , \10715 );
nand \U$10374 ( \10717 , \10716 , \8362 );
nand \U$10375 ( \10718 , \10711 , \10717 );
not \U$10376 ( \10719 , \10718 );
not \U$10377 ( \10720 , \2980 );
and \U$10378 ( \10721 , RIbb2ead0_25, \5550 );
not \U$10379 ( \10722 , RIbb2ead0_25);
and \U$10380 ( \10723 , \10722 , \3311 );
or \U$10381 ( \10724 , \10721 , \10723 );
not \U$10382 ( \10725 , \10724 );
or \U$10383 ( \10726 , \10720 , \10725 );
nand \U$10384 ( \10727 , \10387 , \2963 );
nand \U$10385 ( \10728 , \10726 , \10727 );
not \U$10386 ( \10729 , \10728 );
or \U$10387 ( \10730 , \10719 , \10729 );
or \U$10388 ( \10731 , \10728 , \10718 );
not \U$10389 ( \10732 , \3407 );
not \U$10390 ( \10733 , RIbb2ebc0_23);
not \U$10391 ( \10734 , \3517 );
or \U$10392 ( \10735 , \10733 , \10734 );
nand \U$10393 ( \10736 , \3521 , \3388 );
nand \U$10394 ( \10737 , \10735 , \10736 );
not \U$10395 ( \10738 , \10737 );
or \U$10396 ( \10739 , \10732 , \10738 );
nand \U$10397 ( \10740 , \10257 , \3383 );
nand \U$10398 ( \10741 , \10739 , \10740 );
nand \U$10399 ( \10742 , \10731 , \10741 );
nand \U$10400 ( \10743 , \10730 , \10742 );
xor \U$10401 ( \10744 , \10121 , \10132 );
xor \U$10402 ( \10745 , \10744 , \10143 );
or \U$10403 ( \10746 , \10743 , \10745 );
buf \U$10404 ( \10747 , \507 );
not \U$10405 ( \10748 , \10747 );
nand \U$10406 ( \10749 , \595 , \596 );
nor \U$10407 ( \10750 , \10748 , \10749 );
not \U$10408 ( \10751 , \10750 );
not \U$10409 ( \10752 , \4360 );
or \U$10410 ( \10753 , \10751 , \10752 );
not \U$10411 ( \10754 , \10747 );
nand \U$10412 ( \10755 , \536 , \540 );
not \U$10413 ( \10756 , \10755 );
or \U$10414 ( \10757 , \10754 , \10756 );
nand \U$10415 ( \10758 , RIbb2c2f8_110, RIbb32b08_174);
nand \U$10416 ( \10759 , \10757 , \10758 );
not \U$10417 ( \10760 , \10759 );
nand \U$10418 ( \10761 , \10753 , \10760 );
nand \U$10419 ( \10762 , \495 , \539 );
xnor \U$10420 ( \10763 , \10761 , \10762 );
buf \U$10421 ( \10764 , \10763 );
and \U$10422 ( \10765 , \1313 , \10764 );
not \U$10423 ( \10766 , \2940 );
not \U$10424 ( \10767 , RIbb2e800_31);
not \U$10425 ( \10768 , \1284 );
or \U$10426 ( \10769 , \10767 , \10768 );
nand \U$10427 ( \10770 , \1283 , \4096 );
nand \U$10428 ( \10771 , \10769 , \10770 );
not \U$10429 ( \10772 , \10771 );
or \U$10430 ( \10773 , \10766 , \10772 );
nand \U$10431 ( \10774 , \10290 , \3613 );
nand \U$10432 ( \10775 , \10773 , \10774 );
xor \U$10433 ( \10776 , \10765 , \10775 );
not \U$10434 ( \10777 , \1517 );
not \U$10435 ( \10778 , \10470 );
or \U$10436 ( \10779 , \10777 , \10778 );
and \U$10437 ( \10780 , RIbb2ef80_15, \3276 );
not \U$10438 ( \10781 , RIbb2ef80_15);
and \U$10439 ( \10782 , \10781 , \3275 );
or \U$10440 ( \10783 , \10780 , \10782 );
nand \U$10441 ( \10784 , \10783 , \1445 );
nand \U$10442 ( \10785 , \10779 , \10784 );
and \U$10443 ( \10786 , \10776 , \10785 );
and \U$10444 ( \10787 , \10765 , \10775 );
or \U$10445 ( \10788 , \10786 , \10787 );
nand \U$10446 ( \10789 , \10746 , \10788 );
nand \U$10447 ( \10790 , \10743 , \10745 );
nand \U$10448 ( \10791 , \10789 , \10790 );
nand \U$10449 ( \10792 , \10708 , \10791 );
nand \U$10450 ( \10793 , \10654 , \10707 );
nand \U$10451 ( \10794 , \10792 , \10793 );
and \U$10452 ( \10795 , \10652 , \10794 );
and \U$10453 ( \10796 , \10649 , \10651 );
or \U$10454 ( \10797 , \10795 , \10796 );
nand \U$10455 ( \10798 , \10638 , \10797 );
nand \U$10456 ( \10799 , \10521 , \10637 );
and \U$10457 ( \10800 , \10798 , \10799 );
xor \U$10458 ( \10801 , \10060 , \10076 );
xnor \U$10459 ( \10802 , \10801 , \10012 );
xor \U$10460 ( \10803 , \10800 , \10802 );
xor \U$10461 ( \10804 , \10344 , \10347 );
xor \U$10462 ( \10805 , \10804 , \10512 );
and \U$10463 ( \10806 , \10803 , \10805 );
and \U$10464 ( \10807 , \10800 , \10802 );
or \U$10465 ( \10808 , \10806 , \10807 );
xor \U$10466 ( \10809 , \10519 , \10808 );
and \U$10467 ( \10810 , \10341 , \10342 );
not \U$10468 ( \10811 , \10341 );
and \U$10469 ( \10812 , \10811 , \10337 );
nor \U$10470 ( \10813 , \10810 , \10812 );
xor \U$10471 ( \10814 , \10322 , \10813 );
not \U$10472 ( \10815 , \10814 );
xor \U$10473 ( \10816 , \10149 , \10232 );
xor \U$10474 ( \10817 , \10816 , \10319 );
not \U$10475 ( \10818 , \10483 );
not \U$10476 ( \10819 , \10367 );
or \U$10477 ( \10820 , \10818 , \10819 );
or \U$10478 ( \10821 , \10483 , \10367 );
nand \U$10479 ( \10822 , \10820 , \10821 );
and \U$10480 ( \10823 , \10822 , \10503 );
not \U$10481 ( \10824 , \10822 );
not \U$10482 ( \10825 , \10503 );
and \U$10483 ( \10826 , \10824 , \10825 );
nor \U$10484 ( \10827 , \10823 , \10826 );
xor \U$10485 ( \10828 , \10817 , \10827 );
xor \U$10486 ( \10829 , \10191 , \10188 );
xor \U$10487 ( \10830 , \10829 , \10227 );
not \U$10488 ( \10831 , \10830 );
xor \U$10489 ( \10832 , \10404 , \10442 );
xor \U$10490 ( \10833 , \10832 , \10479 );
not \U$10491 ( \10834 , \10833 );
not \U$10492 ( \10835 , \10834 );
or \U$10493 ( \10836 , \10831 , \10835 );
not \U$10494 ( \10837 , RIbb2e8f0_29);
not \U$10495 ( \10838 , \4341 );
or \U$10496 ( \10839 , \10837 , \10838 );
nand \U$10497 ( \10840 , \4340 , \3440 );
nand \U$10498 ( \10841 , \10839 , \10840 );
and \U$10499 ( \10842 , \10841 , \2922 );
and \U$10500 ( \10843 , \10413 , \2925 );
nor \U$10501 ( \10844 , \10842 , \10843 );
not \U$10502 ( \10845 , \10844 );
not \U$10503 ( \10846 , \10845 );
not \U$10504 ( \10847 , \998 );
not \U$10505 ( \10848 , \10460 );
or \U$10506 ( \10849 , \10847 , \10848 );
not \U$10507 ( \10850 , RIbb2f070_13);
not \U$10508 ( \10851 , \4088 );
or \U$10509 ( \10852 , \10850 , \10851 );
nand \U$10510 ( \10853 , \4324 , \1656 );
nand \U$10511 ( \10854 , \10852 , \10853 );
nand \U$10512 ( \10855 , \10854 , \916 );
nand \U$10513 ( \10856 , \10849 , \10855 );
not \U$10514 ( \10857 , \10856 );
or \U$10515 ( \10858 , \10846 , \10857 );
not \U$10516 ( \10859 , \10856 );
not \U$10517 ( \10860 , \10859 );
not \U$10518 ( \10861 , \10844 );
or \U$10519 ( \10862 , \10860 , \10861 );
not \U$10520 ( \10863 , \10451 );
not \U$10521 ( \10864 , \10448 );
or \U$10522 ( \10865 , \10863 , \10864 );
not \U$10523 ( \10866 , RIbb2e260_43);
not \U$10524 ( \10867 , \1509 );
or \U$10525 ( \10868 , \10866 , \10867 );
nand \U$10526 ( \10869 , \4315 , \8347 );
nand \U$10527 ( \10870 , \10868 , \10869 );
nand \U$10528 ( \10871 , \10870 , \10449 );
nand \U$10529 ( \10872 , \10865 , \10871 );
nand \U$10530 ( \10873 , \10862 , \10872 );
nand \U$10531 ( \10874 , \10858 , \10873 );
not \U$10532 ( \10875 , \10874 );
not \U$10533 ( \10876 , \10875 );
not \U$10534 ( \10877 , \832 );
and \U$10535 ( \10878 , \5962 , RIbb2ee90_17);
not \U$10536 ( \10879 , \5962 );
and \U$10537 ( \10880 , \10879 , \2240 );
or \U$10538 ( \10881 , \10878 , \10880 );
not \U$10539 ( \10882 , \10881 );
or \U$10540 ( \10883 , \10877 , \10882 );
nand \U$10541 ( \10884 , \10211 , \836 );
nand \U$10542 ( \10885 , \10883 , \10884 );
xor \U$10543 ( \10886 , \10561 , \10885 );
not \U$10544 ( \10887 , \855 );
not \U$10545 ( \10888 , \10222 );
or \U$10546 ( \10889 , \10887 , \10888 );
and \U$10547 ( \10890 , \3228 , \5277 );
not \U$10548 ( \10891 , \3228 );
and \U$10549 ( \10892 , \10891 , RIbb2eda0_19);
or \U$10550 ( \10893 , \10890 , \10892 );
nand \U$10551 ( \10894 , \10893 , \853 );
nand \U$10552 ( \10895 , \10889 , \10894 );
and \U$10553 ( \10896 , \10886 , \10895 );
and \U$10554 ( \10897 , \10561 , \10885 );
or \U$10555 ( \10898 , \10896 , \10897 );
not \U$10556 ( \10899 , \10898 );
not \U$10557 ( \10900 , \10899 );
or \U$10558 ( \10901 , \10876 , \10900 );
not \U$10559 ( \10902 , \8450 );
not \U$10560 ( \10903 , \10423 );
or \U$10561 ( \10904 , \10902 , \10903 );
not \U$10562 ( \10905 , RIbb2e440_39);
not \U$10563 ( \10906 , \4284 );
or \U$10564 ( \10907 , \10905 , \10906 );
not \U$10565 ( \10908 , RIbb2e440_39);
nand \U$10566 ( \10909 , \3099 , \10908 );
nand \U$10567 ( \10910 , \10907 , \10909 );
nand \U$10568 ( \10911 , \10910 , \8445 );
nand \U$10569 ( \10912 , \10904 , \10911 );
not \U$10570 ( \10913 , \6242 );
not \U$10571 ( \10914 , \10398 );
or \U$10572 ( \10915 , \10913 , \10914 );
not \U$10573 ( \10916 , RIbb2e530_37);
not \U$10574 ( \10917 , \4299 );
or \U$10575 ( \10918 , \10916 , \10917 );
nand \U$10576 ( \10919 , \3472 , \6246 );
nand \U$10577 ( \10920 , \10918 , \10919 );
nand \U$10578 ( \10921 , \10920 , \6251 );
nand \U$10579 ( \10922 , \10915 , \10921 );
xor \U$10580 ( \10923 , \10912 , \10922 );
not \U$10581 ( \10924 , \3465 );
not \U$10582 ( \10925 , \10436 );
or \U$10583 ( \10926 , \10924 , \10925 );
not \U$10584 ( \10927 , RIbb2e9e0_27);
not \U$10585 ( \10928 , \1340 );
or \U$10586 ( \10929 , \10927 , \10928 );
nand \U$10587 ( \10930 , \1339 , \6065 );
nand \U$10588 ( \10931 , \10929 , \10930 );
nand \U$10589 ( \10932 , \10931 , \3445 );
nand \U$10590 ( \10933 , \10926 , \10932 );
and \U$10591 ( \10934 , \10923 , \10933 );
and \U$10592 ( \10935 , \10912 , \10922 );
or \U$10593 ( \10936 , \10934 , \10935 );
nand \U$10594 ( \10937 , \10901 , \10936 );
nand \U$10595 ( \10938 , \10898 , \10874 );
nand \U$10596 ( \10939 , \10937 , \10938 );
nand \U$10597 ( \10940 , \10836 , \10939 );
not \U$10598 ( \10941 , \10830 );
nand \U$10599 ( \10942 , \10833 , \10941 );
nand \U$10600 ( \10943 , \10940 , \10942 );
and \U$10601 ( \10944 , \10828 , \10943 );
and \U$10602 ( \10945 , \10817 , \10827 );
or \U$10603 ( \10946 , \10944 , \10945 );
not \U$10604 ( \10947 , \10946 );
nand \U$10605 ( \10948 , \10815 , \10947 );
xor \U$10606 ( \10949 , \10357 , \10509 );
buf \U$10607 ( \10950 , \10506 );
xor \U$10608 ( \10951 , \10949 , \10950 );
and \U$10609 ( \10952 , \10948 , \10951 );
not \U$10610 ( \10953 , \10814 );
nor \U$10611 ( \10954 , \10953 , \10947 );
nor \U$10612 ( \10955 , \10952 , \10954 );
xor \U$10613 ( \10956 , \10637 , \10521 );
xnor \U$10614 ( \10957 , \10956 , \10797 );
not \U$10615 ( \10958 , \10957 );
xor \U$10616 ( \10959 , \10649 , \10651 );
xor \U$10617 ( \10960 , \10959 , \10794 );
and \U$10618 ( \10961 , \10278 , \10239 );
not \U$10619 ( \10962 , \10278 );
not \U$10620 ( \10963 , \10239 );
and \U$10621 ( \10964 , \10962 , \10963 );
nor \U$10622 ( \10965 , \10961 , \10964 );
not \U$10623 ( \10966 , \10965 );
not \U$10624 ( \10967 , \10317 );
not \U$10625 ( \10968 , \10967 );
and \U$10626 ( \10969 , \10966 , \10968 );
and \U$10627 ( \10970 , \10965 , \10967 );
nor \U$10628 ( \10971 , \10969 , \10970 );
not \U$10629 ( \10972 , \10971 );
not \U$10630 ( \10973 , \10972 );
not \U$10631 ( \10974 , \10494 );
not \U$10632 ( \10975 , \10498 );
or \U$10633 ( \10976 , \10974 , \10975 );
or \U$10634 ( \10977 , \10498 , \10494 );
nand \U$10635 ( \10978 , \10976 , \10977 );
and \U$10636 ( \10979 , \10978 , \10491 );
not \U$10637 ( \10980 , \10978 );
and \U$10638 ( \10981 , \10980 , \10501 );
nor \U$10639 ( \10982 , \10979 , \10981 );
not \U$10640 ( \10983 , \10982 );
not \U$10641 ( \10984 , \10983 );
or \U$10642 ( \10985 , \10973 , \10984 );
not \U$10643 ( \10986 , \10971 );
not \U$10644 ( \10987 , \10982 );
or \U$10645 ( \10988 , \10986 , \10987 );
xor \U$10646 ( \10989 , \10427 , \10440 );
xor \U$10647 ( \10990 , \10989 , \10415 );
not \U$10648 ( \10991 , \10990 );
xor \U$10649 ( \10992 , \10203 , \10213 );
xor \U$10650 ( \10993 , \10992 , \10224 );
not \U$10651 ( \10994 , \10993 );
or \U$10652 ( \10995 , \10991 , \10994 );
or \U$10653 ( \10996 , \10990 , \10993 );
xor \U$10654 ( \10997 , \10274 , \10262 );
xnor \U$10655 ( \10998 , \10997 , \10250 );
nand \U$10656 ( \10999 , \10996 , \10998 );
nand \U$10657 ( \11000 , \10995 , \10999 );
nand \U$10658 ( \11001 , \10988 , \11000 );
nand \U$10659 ( \11002 , \10985 , \11001 );
or \U$10660 ( \11003 , \10960 , \11002 );
not \U$10661 ( \11004 , \10524 );
not \U$10662 ( \11005 , \10527 );
or \U$10663 ( \11006 , \11004 , \11005 );
nand \U$10664 ( \11007 , \10528 , \10523 );
nand \U$10665 ( \11008 , \11006 , \11007 );
not \U$10666 ( \11009 , \10635 );
and \U$10667 ( \11010 , \11008 , \11009 );
not \U$10668 ( \11011 , \11008 );
and \U$10669 ( \11012 , \11011 , \10635 );
nor \U$10670 ( \11013 , \11010 , \11012 );
not \U$10671 ( \11014 , \11013 );
nand \U$10672 ( \11015 , \11003 , \11014 );
nand \U$10673 ( \11016 , \10960 , \11002 );
nand \U$10674 ( \11017 , \11015 , \11016 );
not \U$10675 ( \11018 , \11017 );
not \U$10676 ( \11019 , \11018 );
or \U$10677 ( \11020 , \10958 , \11019 );
and \U$10678 ( \11021 , \10936 , \10875 );
not \U$10679 ( \11022 , \10936 );
and \U$10680 ( \11023 , \11022 , \10874 );
or \U$10681 ( \11024 , \11021 , \11023 );
and \U$10682 ( \11025 , \11024 , \10898 );
not \U$10683 ( \11026 , \11024 );
and \U$10684 ( \11027 , \11026 , \10899 );
nor \U$10685 ( \11028 , \11025 , \11027 );
xnor \U$10686 ( \11029 , \10701 , \10705 );
and \U$10687 ( \11030 , \11029 , \10697 );
not \U$10688 ( \11031 , \11029 );
and \U$10689 ( \11032 , \11031 , \10696 );
nor \U$10690 ( \11033 , \11030 , \11032 );
or \U$10691 ( \11034 , \11028 , \11033 );
xor \U$10692 ( \11035 , \10998 , \10993 );
xor \U$10693 ( \11036 , \11035 , \10990 );
nand \U$10694 ( \11037 , \11034 , \11036 );
nand \U$10695 ( \11038 , \11033 , \11028 );
nand \U$10696 ( \11039 , \11037 , \11038 );
not \U$10697 ( \11040 , \11039 );
xor \U$10698 ( \11041 , \10654 , \10707 );
xnor \U$10699 ( \11042 , \11041 , \10791 );
not \U$10700 ( \11043 , \11042 );
not \U$10701 ( \11044 , \11043 );
or \U$10702 ( \11045 , \11040 , \11044 );
not \U$10703 ( \11046 , \11042 );
not \U$10704 ( \11047 , \11039 );
not \U$10705 ( \11048 , \11047 );
or \U$10706 ( \11049 , \11046 , \11048 );
not \U$10707 ( \11050 , \2941 );
not \U$10708 ( \11051 , \10771 );
or \U$10709 ( \11052 , \11050 , \11051 );
not \U$10710 ( \11053 , RIbb2e800_31);
not \U$10711 ( \11054 , \3109 );
not \U$10712 ( \11055 , \11054 );
or \U$10713 ( \11056 , \11053 , \11055 );
nand \U$10714 ( \11057 , \3109 , \2917 );
nand \U$10715 ( \11058 , \11056 , \11057 );
nand \U$10716 ( \11059 , \11058 , \2940 );
nand \U$10717 ( \11060 , \11052 , \11059 );
not \U$10718 ( \11061 , \10117 );
not \U$10719 ( \11062 , RIbb2e170_45);
not \U$10720 ( \11063 , \2946 );
or \U$10721 ( \11064 , \11062 , \11063 );
not \U$10722 ( \11065 , RIbb2e170_45);
nand \U$10723 ( \11066 , \893 , \11065 );
nand \U$10724 ( \11067 , \11064 , \11066 );
not \U$10725 ( \11068 , \11067 );
or \U$10726 ( \11069 , \11061 , \11068 );
nand \U$10727 ( \11070 , \10119 , \10606 );
nand \U$10728 ( \11071 , \11069 , \11070 );
xor \U$10729 ( \11072 , \11060 , \11071 );
not \U$10730 ( \11073 , \8995 );
not \U$10731 ( \11074 , \10716 );
or \U$10732 ( \11075 , \11073 , \11074 );
not \U$10733 ( \11076 , RIbb2e350_41);
not \U$10734 ( \11077 , \3981 );
or \U$10735 ( \11078 , \11076 , \11077 );
nand \U$10736 ( \11079 , \952 , \8357 );
nand \U$10737 ( \11080 , \11078 , \11079 );
nand \U$10738 ( \11081 , \11080 , \8362 );
nand \U$10739 ( \11082 , \11075 , \11081 );
and \U$10740 ( \11083 , \11072 , \11082 );
and \U$10741 ( \11084 , \11060 , \11071 );
or \U$10742 ( \11085 , \11083 , \11084 );
xor \U$10743 ( \11086 , \10912 , \10922 );
xor \U$10744 ( \11087 , \11086 , \10933 );
xor \U$10745 ( \11088 , \11085 , \11087 );
xor \U$10746 ( \11089 , \10561 , \10885 );
xor \U$10747 ( \11090 , \11089 , \10895 );
and \U$10748 ( \11091 , \11088 , \11090 );
and \U$10749 ( \11092 , \11085 , \11087 );
or \U$10750 ( \11093 , \11091 , \11092 );
not \U$10751 ( \11094 , \11093 );
xor \U$10752 ( \11095 , \10745 , \10788 );
xnor \U$10753 ( \11096 , \11095 , \10743 );
not \U$10754 ( \11097 , \11096 );
not \U$10755 ( \11098 , \11097 );
or \U$10756 ( \11099 , \11094 , \11098 );
not \U$10757 ( \11100 , \11096 );
not \U$10758 ( \11101 , \11093 );
not \U$10759 ( \11102 , \11101 );
or \U$10760 ( \11103 , \11100 , \11102 );
xor \U$10761 ( \11104 , \10765 , \10775 );
xor \U$10762 ( \11105 , \11104 , \10785 );
xor \U$10763 ( \11106 , \10728 , \10741 );
xor \U$10764 ( \11107 , \11106 , \10718 );
xor \U$10765 ( \11108 , \11105 , \11107 );
and \U$10766 ( \11109 , \10872 , \10844 );
not \U$10767 ( \11110 , \10872 );
and \U$10768 ( \11111 , \11110 , \10845 );
nor \U$10769 ( \11112 , \11109 , \11111 );
xor \U$10770 ( \11113 , \11112 , \10859 );
and \U$10771 ( \11114 , \11108 , \11113 );
and \U$10772 ( \11115 , \11105 , \11107 );
or \U$10773 ( \11116 , \11114 , \11115 );
nand \U$10774 ( \11117 , \11103 , \11116 );
nand \U$10775 ( \11118 , \11099 , \11117 );
nand \U$10776 ( \11119 , \11049 , \11118 );
nand \U$10777 ( \11120 , \11045 , \11119 );
xor \U$10778 ( \11121 , \10389 , \10379 );
xor \U$10779 ( \11122 , \11121 , \10402 );
not \U$10780 ( \11123 , \10477 );
not \U$10781 ( \11124 , \10463 );
or \U$10782 ( \11125 , \11123 , \11124 );
nand \U$10783 ( \11126 , \10476 , \10453 );
nand \U$10784 ( \11127 , \11125 , \11126 );
xor \U$10785 ( \11128 , \11127 , \10474 );
xor \U$10786 ( \11129 , \11122 , \11128 );
not \U$10787 ( \11130 , \10749 );
not \U$10788 ( \11131 , \11130 );
not \U$10789 ( \11132 , \5941 );
or \U$10790 ( \11133 , \11131 , \11132 );
not \U$10791 ( \11134 , \10755 );
nand \U$10792 ( \11135 , \11133 , \11134 );
nand \U$10793 ( \11136 , \10747 , \10758 );
not \U$10794 ( \11137 , \11136 );
and \U$10795 ( \11138 , \11135 , \11137 );
not \U$10796 ( \11139 , \11135 );
and \U$10797 ( \11140 , \11139 , \11136 );
nor \U$10798 ( \11141 , \11138 , \11140 );
buf \U$10799 ( \11142 , \11141 );
not \U$10800 ( \11143 , \11142 );
not \U$10801 ( \11144 , \11143 );
buf \U$10802 ( \11145 , \11144 );
and \U$10803 ( \11146 , \1394 , \11145 );
not \U$10804 ( \11147 , \1429 );
xor \U$10805 ( \11148 , \1313 , \10764 );
not \U$10806 ( \11149 , \11148 );
or \U$10807 ( \11150 , \11147 , \11149 );
nand \U$10808 ( \11151 , \10614 , \1376 );
nand \U$10809 ( \11152 , \11150 , \11151 );
xor \U$10810 ( \11153 , \11146 , \11152 );
not \U$10811 ( \11154 , \1265 );
not \U$10812 ( \11155 , \1290 );
not \U$10813 ( \11156 , \10306 );
or \U$10814 ( \11157 , \11155 , \11156 );
nand \U$10815 ( \11158 , \9841 , \1245 );
nand \U$10816 ( \11159 , \11157 , \11158 );
not \U$10817 ( \11160 , \11159 );
or \U$10818 ( \11161 , \11154 , \11160 );
nand \U$10819 ( \11162 , \10625 , \1294 );
nand \U$10820 ( \11163 , \11161 , \11162 );
and \U$10821 ( \11164 , \11153 , \11163 );
and \U$10822 ( \11165 , \11146 , \11152 );
or \U$10823 ( \11166 , \11164 , \11165 );
not \U$10824 ( \11167 , RIbb2e008_48);
and \U$10825 ( \11168 , \11167 , RIbb2e080_47);
and \U$10826 ( \11169 , \10113 , RIbb2e008_48);
nor \U$10827 ( \11170 , \11168 , \11169 );
and \U$10828 ( \11171 , RIbb2df90_49, \11167 );
not \U$10829 ( \11172 , RIbb2df90_49);
and \U$10830 ( \11173 , \11172 , RIbb2e008_48);
or \U$10831 ( \11174 , \11171 , \11173 );
nor \U$10832 ( \11175 , \11170 , \11174 );
buf \U$10833 ( \11176 , \11175 );
buf \U$10834 ( \11177 , \11174 );
or \U$10835 ( \11178 , \11176 , \11177 );
nand \U$10836 ( \11179 , \11178 , RIbb2e080_47);
not \U$10837 ( \11180 , \1011 );
and \U$10838 ( \11181 , RIbb2f160_11, \6231 );
not \U$10839 ( \11182 , RIbb2f160_11);
and \U$10840 ( \11183 , \11182 , \7111 );
or \U$10841 ( \11184 , \11181 , \11183 );
not \U$10842 ( \11185 , \11184 );
or \U$10843 ( \11186 , \11180 , \11185 );
nand \U$10844 ( \11187 , \10559 , \1077 );
nand \U$10845 ( \11188 , \11186 , \11187 );
xor \U$10846 ( \11189 , \11179 , \11188 );
not \U$10847 ( \11190 , \998 );
not \U$10848 ( \11191 , \10854 );
or \U$10849 ( \11192 , \11190 , \11191 );
not \U$10850 ( \11193 , RIbb2f070_13);
not \U$10851 ( \11194 , \4393 );
or \U$10852 ( \11195 , \11193 , \11194 );
nand \U$10853 ( \11196 , \6269 , \3421 );
nand \U$10854 ( \11197 , \11195 , \11196 );
nand \U$10855 ( \11198 , \11197 , \916 );
nand \U$10856 ( \11199 , \11192 , \11198 );
and \U$10857 ( \11200 , \11189 , \11199 );
and \U$10858 ( \11201 , \11179 , \11188 );
or \U$10859 ( \11202 , \11200 , \11201 );
xor \U$10860 ( \11203 , \11166 , \11202 );
not \U$10861 ( \11204 , \1147 );
not \U$10862 ( \11205 , \10590 );
or \U$10863 ( \11206 , \11204 , \11205 );
not \U$10864 ( \11207 , RIbb2f430_5);
not \U$10865 ( \11208 , \10175 );
or \U$10866 ( \11209 , \11207 , \11208 );
nand \U$10867 ( \11210 , \10178 , \1980 );
nand \U$10868 ( \11211 , \11209 , \11210 );
nand \U$10869 ( \11212 , \11211 , \1090 );
nand \U$10870 ( \11213 , \11206 , \11212 );
not \U$10871 ( \11214 , \1570 );
not \U$10872 ( \11215 , \10581 );
or \U$10873 ( \11216 , \11214 , \11215 );
not \U$10874 ( \11217 , RIbb2f250_9);
not \U$10875 ( \11218 , \10156 );
not \U$10876 ( \11219 , \11218 );
or \U$10877 ( \11220 , \11217 , \11219 );
nand \U$10878 ( \11221 , \10156 , \5064 );
nand \U$10879 ( \11222 , \11220 , \11221 );
nand \U$10880 ( \11223 , \11222 , \1533 );
nand \U$10881 ( \11224 , \11216 , \11223 );
xor \U$10882 ( \11225 , \11213 , \11224 );
not \U$10883 ( \11226 , \1737 );
not \U$10884 ( \11227 , \10568 );
or \U$10885 ( \11228 , \11226 , \11227 );
not \U$10886 ( \11229 , RIbb2f340_7);
not \U$10887 ( \11230 , \9071 );
or \U$10888 ( \11231 , \11229 , \11230 );
not \U$10889 ( \11232 , \7299 );
not \U$10890 ( \11233 , \11232 );
nand \U$10891 ( \11234 , \11233 , \2700 );
nand \U$10892 ( \11235 , \11231 , \11234 );
nand \U$10893 ( \11236 , \11235 , \1702 );
nand \U$10894 ( \11237 , \11228 , \11236 );
and \U$10895 ( \11238 , \11225 , \11237 );
and \U$10896 ( \11239 , \11213 , \11224 );
or \U$10897 ( \11240 , \11238 , \11239 );
and \U$10898 ( \11241 , \11203 , \11240 );
and \U$10899 ( \11242 , \11166 , \11202 );
or \U$10900 ( \11243 , \11241 , \11242 );
and \U$10901 ( \11244 , \11129 , \11243 );
and \U$10902 ( \11245 , \11122 , \11128 );
or \U$10903 ( \11246 , \11244 , \11245 );
xor \U$10904 ( \11247 , \10535 , \10544 );
xor \U$10905 ( \11248 , \11247 , \10633 );
xor \U$10906 ( \11249 , \11246 , \11248 );
xor \U$10907 ( \11250 , \10562 , \10597 );
xor \U$10908 ( \11251 , \11250 , \10630 );
xor \U$10909 ( \11252 , \10610 , \10616 );
xor \U$10910 ( \11253 , \11252 , \10627 );
not \U$10911 ( \11254 , \7103 );
and \U$10912 ( \11255 , RIbb2e440_39, \4595 );
not \U$10913 ( \11256 , RIbb2e440_39);
and \U$10914 ( \11257 , \11256 , \1038 );
or \U$10915 ( \11258 , \11255 , \11257 );
not \U$10916 ( \11259 , \11258 );
or \U$10917 ( \11260 , \11254 , \11259 );
nand \U$10918 ( \11261 , \10910 , \8450 );
nand \U$10919 ( \11262 , \11260 , \11261 );
not \U$10920 ( \11263 , \11262 );
not \U$10921 ( \11264 , \11263 );
not \U$10922 ( \11265 , \2925 );
not \U$10923 ( \11266 , \10841 );
or \U$10924 ( \11267 , \11265 , \11266 );
not \U$10925 ( \11268 , RIbb2e8f0_29);
not \U$10926 ( \11269 , \3822 );
or \U$10927 ( \11270 , \11268 , \11269 );
nand \U$10928 ( \11271 , \3821 , \2911 );
nand \U$10929 ( \11272 , \11270 , \11271 );
nand \U$10930 ( \11273 , \11272 , \2922 );
nand \U$10931 ( \11274 , \11267 , \11273 );
not \U$10932 ( \11275 , \11274 );
not \U$10933 ( \11276 , \11275 );
or \U$10934 ( \11277 , \11264 , \11276 );
not \U$10935 ( \11278 , \3465 );
not \U$10936 ( \11279 , \10931 );
or \U$10937 ( \11280 , \11278 , \11279 );
not \U$10938 ( \11281 , RIbb2e9e0_27);
not \U$10939 ( \11282 , \1853 );
or \U$10940 ( \11283 , \11281 , \11282 );
not \U$10941 ( \11284 , RIbb2e9e0_27);
nand \U$10942 ( \11285 , \4610 , \11284 );
nand \U$10943 ( \11286 , \11283 , \11285 );
nand \U$10944 ( \11287 , \11286 , \3445 );
nand \U$10945 ( \11288 , \11280 , \11287 );
nand \U$10946 ( \11289 , \11277 , \11288 );
nand \U$10947 ( \11290 , \11274 , \11262 );
nand \U$10948 ( \11291 , \11289 , \11290 );
xor \U$10949 ( \11292 , \11253 , \11291 );
not \U$10950 ( \11293 , \3887 );
not \U$10951 ( \11294 , RIbb2e710_33);
not \U$10952 ( \11295 , \1113 );
or \U$10953 ( \11296 , \11294 , \11295 );
nand \U$10954 ( \11297 , \4006 , \6058 );
nand \U$10955 ( \11298 , \11296 , \11297 );
not \U$10956 ( \11299 , \11298 );
or \U$10957 ( \11300 , \11293 , \11299 );
nand \U$10958 ( \11301 , \10675 , \4791 );
nand \U$10959 ( \11302 , \11300 , \11301 );
not \U$10960 ( \11303 , \836 );
not \U$10961 ( \11304 , \10881 );
or \U$10962 ( \11305 , \11303 , \11304 );
not \U$10963 ( \11306 , RIbb2ee90_17);
not \U$10964 ( \11307 , \4031 );
or \U$10965 ( \11308 , \11306 , \11307 );
nand \U$10966 ( \11309 , \4030 , \3699 );
nand \U$10967 ( \11310 , \11308 , \11309 );
nand \U$10968 ( \11311 , \11310 , \832 );
nand \U$10969 ( \11312 , \11305 , \11311 );
xor \U$10970 ( \11313 , \11302 , \11312 );
not \U$10971 ( \11314 , \3105 );
not \U$10972 ( \11315 , \10783 );
or \U$10973 ( \11316 , \11314 , \11315 );
and \U$10974 ( \11317 , RIbb2ef80_15, \4040 );
not \U$10975 ( \11318 , RIbb2ef80_15);
and \U$10976 ( \11319 , \11318 , \6013 );
or \U$10977 ( \11320 , \11317 , \11319 );
nand \U$10978 ( \11321 , \11320 , \1445 );
nand \U$10979 ( \11322 , \11316 , \11321 );
and \U$10980 ( \11323 , \11313 , \11322 );
and \U$10981 ( \11324 , \11302 , \11312 );
or \U$10982 ( \11325 , \11323 , \11324 );
and \U$10983 ( \11326 , \11292 , \11325 );
and \U$10984 ( \11327 , \11253 , \11291 );
or \U$10985 ( \11328 , \11326 , \11327 );
xor \U$10986 ( \11329 , \11251 , \11328 );
xor \U$10987 ( \11330 , \10572 , \10583 );
xor \U$10988 ( \11331 , \11330 , \10594 );
not \U$10989 ( \11332 , \5845 );
not \U$10990 ( \11333 , \10660 );
or \U$10991 ( \11334 , \11332 , \11333 );
not \U$10992 ( \11335 , RIbb2e620_35);
not \U$10993 ( \11336 , \3773 );
or \U$10994 ( \11337 , \11335 , \11336 );
not \U$10995 ( \11338 , RIbb2e620_35);
nand \U$10996 ( \11339 , \7033 , \11338 );
nand \U$10997 ( \11340 , \11337 , \11339 );
nand \U$10998 ( \11341 , \11340 , \4712 );
nand \U$10999 ( \11342 , \11334 , \11341 );
not \U$11000 ( \11343 , \11342 );
not \U$11001 ( \11344 , \3383 );
not \U$11002 ( \11345 , \10737 );
or \U$11003 ( \11346 , \11344 , \11345 );
not \U$11004 ( \11347 , RIbb2ebc0_23);
not \U$11005 ( \11348 , \4216 );
or \U$11006 ( \11349 , \11347 , \11348 );
nand \U$11007 ( \11350 , \3167 , \3396 );
nand \U$11008 ( \11351 , \11349 , \11350 );
nand \U$11009 ( \11352 , \11351 , \3406 );
nand \U$11010 ( \11353 , \11346 , \11352 );
not \U$11011 ( \11354 , \11353 );
or \U$11012 ( \11355 , \11343 , \11354 );
or \U$11013 ( \11356 , \11353 , \11342 );
not \U$11014 ( \11357 , \2078 );
not \U$11015 ( \11358 , \10686 );
or \U$11016 ( \11359 , \11357 , \11358 );
not \U$11017 ( \11360 , RIbb2ecb0_21);
not \U$11018 ( \11361 , \3203 );
or \U$11019 ( \11362 , \11360 , \11361 );
nand \U$11020 ( \11363 , \4640 , \849 );
nand \U$11021 ( \11364 , \11362 , \11363 );
nand \U$11022 ( \11365 , \11364 , \2077 );
nand \U$11023 ( \11366 , \11359 , \11365 );
nand \U$11024 ( \11367 , \11356 , \11366 );
nand \U$11025 ( \11368 , \11355 , \11367 );
xor \U$11026 ( \11369 , \11331 , \11368 );
not \U$11027 ( \11370 , \6251 );
and \U$11028 ( \11371 , \5130 , RIbb2e530_37);
not \U$11029 ( \11372 , \5130 );
and \U$11030 ( \11373 , \11372 , \8701 );
or \U$11031 ( \11374 , \11371 , \11373 );
not \U$11032 ( \11375 , \11374 );
or \U$11033 ( \11376 , \11370 , \11375 );
nand \U$11034 ( \11377 , \10920 , \6242 );
nand \U$11035 ( \11378 , \11376 , \11377 );
not \U$11036 ( \11379 , \10451 );
not \U$11037 ( \11380 , \10870 );
or \U$11038 ( \11381 , \11379 , \11380 );
not \U$11039 ( \11382 , RIbb2e260_43);
not \U$11040 ( \11383 , \7143 );
or \U$11041 ( \11384 , \11382 , \11383 );
nand \U$11042 ( \11385 , \3453 , \8347 );
nand \U$11043 ( \11386 , \11384 , \11385 );
nand \U$11044 ( \11387 , \11386 , \10449 );
nand \U$11045 ( \11388 , \11381 , \11387 );
xor \U$11046 ( \11389 , \11378 , \11388 );
not \U$11047 ( \11390 , \2963 );
not \U$11048 ( \11391 , \10724 );
or \U$11049 ( \11392 , \11390 , \11391 );
and \U$11050 ( \11393 , RIbb2ead0_25, \3319 );
not \U$11051 ( \11394 , RIbb2ead0_25);
and \U$11052 ( \11395 , \11394 , \3320 );
or \U$11053 ( \11396 , \11393 , \11395 );
nand \U$11054 ( \11397 , \11396 , \2980 );
nand \U$11055 ( \11398 , \11392 , \11397 );
and \U$11056 ( \11399 , \11389 , \11398 );
and \U$11057 ( \11400 , \11378 , \11388 );
or \U$11058 ( \11401 , \11399 , \11400 );
and \U$11059 ( \11402 , \11369 , \11401 );
and \U$11060 ( \11403 , \11331 , \11368 );
or \U$11061 ( \11404 , \11402 , \11403 );
and \U$11062 ( \11405 , \11329 , \11404 );
and \U$11063 ( \11406 , \11251 , \11328 );
or \U$11064 ( \11407 , \11405 , \11406 );
and \U$11065 ( \11408 , \11249 , \11407 );
and \U$11066 ( \11409 , \11246 , \11248 );
or \U$11067 ( \11410 , \11408 , \11409 );
or \U$11068 ( \11411 , \11120 , \11410 );
xor \U$11069 ( \11412 , \10817 , \10827 );
xor \U$11070 ( \11413 , \11412 , \10943 );
nand \U$11071 ( \11414 , \11411 , \11413 );
nand \U$11072 ( \11415 , \11120 , \11410 );
nand \U$11073 ( \11416 , \11414 , \11415 );
nand \U$11074 ( \11417 , \11020 , \11416 );
not \U$11075 ( \11418 , \10957 );
nand \U$11076 ( \11419 , \11418 , \11017 );
and \U$11077 ( \11420 , \11417 , \11419 );
xor \U$11078 ( \11421 , \10955 , \11420 );
xor \U$11079 ( \11422 , \10800 , \10802 );
xor \U$11080 ( \11423 , \11422 , \10805 );
and \U$11081 ( \11424 , \11421 , \11423 );
and \U$11082 ( \11425 , \10955 , \11420 );
or \U$11083 ( \11426 , \11424 , \11425 );
nand \U$11084 ( \11427 , \10809 , \11426 );
buf \U$11085 ( \11428 , \11427 );
xor \U$11086 ( \11429 , \10955 , \11420 );
xor \U$11087 ( \11430 , \11429 , \11423 );
buf \U$11088 ( \11431 , \11430 );
not \U$11089 ( \11432 , \11418 );
not \U$11090 ( \11433 , \11018 );
or \U$11091 ( \11434 , \11432 , \11433 );
nand \U$11092 ( \11435 , \11017 , \10957 );
nand \U$11093 ( \11436 , \11434 , \11435 );
xor \U$11094 ( \11437 , \11416 , \11436 );
xor \U$11095 ( \11438 , \10814 , \10951 );
xor \U$11096 ( \11439 , \11438 , \10946 );
or \U$11097 ( \11440 , \11437 , \11439 );
not \U$11098 ( \11441 , \11000 );
not \U$11099 ( \11442 , \10971 );
or \U$11100 ( \11443 , \11441 , \11442 );
or \U$11101 ( \11444 , \11000 , \10971 );
nand \U$11102 ( \11445 , \11443 , \11444 );
and \U$11103 ( \11446 , \11445 , \10983 );
not \U$11104 ( \11447 , \11445 );
not \U$11105 ( \11448 , \10983 );
and \U$11106 ( \11449 , \11447 , \11448 );
nor \U$11107 ( \11450 , \11446 , \11449 );
not \U$11108 ( \11451 , \11450 );
and \U$11109 ( \11452 , \10939 , \10834 );
not \U$11110 ( \11453 , \10939 );
and \U$11111 ( \11454 , \11453 , \10833 );
or \U$11112 ( \11455 , \11452 , \11454 );
and \U$11113 ( \11456 , \11455 , \10830 );
not \U$11114 ( \11457 , \11455 );
and \U$11115 ( \11458 , \11457 , \10941 );
nor \U$11116 ( \11459 , \11456 , \11458 );
nand \U$11117 ( \11460 , \11451 , \11459 );
not \U$11118 ( \11461 , \11460 );
xor \U$11119 ( \11462 , \11246 , \11248 );
xor \U$11120 ( \11463 , \11462 , \11407 );
not \U$11121 ( \11464 , \11463 );
or \U$11122 ( \11465 , \11461 , \11464 );
not \U$11123 ( \11466 , \11459 );
nand \U$11124 ( \11467 , \11466 , \11450 );
nand \U$11125 ( \11468 , \11465 , \11467 );
not \U$11126 ( \11469 , \11468 );
not \U$11127 ( \11470 , \11002 );
not \U$11128 ( \11471 , \11013 );
or \U$11129 ( \11472 , \11470 , \11471 );
or \U$11130 ( \11473 , \11013 , \11002 );
nand \U$11131 ( \11474 , \11472 , \11473 );
and \U$11132 ( \11475 , \11474 , \10960 );
not \U$11133 ( \11476 , \11474 );
not \U$11134 ( \11477 , \10960 );
and \U$11135 ( \11478 , \11476 , \11477 );
nor \U$11136 ( \11479 , \11475 , \11478 );
not \U$11137 ( \11480 , \11479 );
or \U$11138 ( \11481 , \11469 , \11480 );
xor \U$11139 ( \11482 , \11122 , \11128 );
xor \U$11140 ( \11483 , \11482 , \11243 );
not \U$11141 ( \11484 , \10690 );
not \U$11142 ( \11485 , \10678 );
or \U$11143 ( \11486 , \11484 , \11485 );
or \U$11144 ( \11487 , \10690 , \10678 );
nand \U$11145 ( \11488 , \11486 , \11487 );
xnor \U$11146 ( \11489 , \11488 , \10664 );
not \U$11147 ( \11490 , \11489 );
not \U$11148 ( \11491 , \11490 );
xor \U$11149 ( \11492 , \11166 , \11202 );
xor \U$11150 ( \11493 , \11492 , \11240 );
not \U$11151 ( \11494 , \11493 );
or \U$11152 ( \11495 , \11491 , \11494 );
not \U$11153 ( \11496 , \11489 );
not \U$11154 ( \11497 , \11493 );
not \U$11155 ( \11498 , \11497 );
or \U$11156 ( \11499 , \11496 , \11498 );
not \U$11157 ( \11500 , \998 );
not \U$11158 ( \11501 , \11197 );
or \U$11159 ( \11502 , \11500 , \11501 );
not \U$11160 ( \11503 , RIbb2f070_13);
not \U$11161 ( \11504 , \10552 );
or \U$11162 ( \11505 , \11503 , \11504 );
nand \U$11163 ( \11506 , \6202 , \1656 );
nand \U$11164 ( \11507 , \11505 , \11506 );
nand \U$11165 ( \11508 , \11507 , \916 );
nand \U$11166 ( \11509 , \11502 , \11508 );
not \U$11167 ( \11510 , \855 );
not \U$11168 ( \11511 , \10893 );
or \U$11169 ( \11512 , \11510 , \11511 );
not \U$11170 ( \11513 , RIbb2eda0_19);
not \U$11171 ( \11514 , \7018 );
or \U$11172 ( \11515 , \11513 , \11514 );
nand \U$11173 ( \11516 , \3654 , \5277 );
nand \U$11174 ( \11517 , \11515 , \11516 );
nand \U$11175 ( \11518 , \11517 , \853 );
nand \U$11176 ( \11519 , \11512 , \11518 );
xor \U$11177 ( \11520 , \11509 , \11519 );
not \U$11178 ( \11521 , \1737 );
not \U$11179 ( \11522 , \11235 );
or \U$11180 ( \11523 , \11521 , \11522 );
and \U$11181 ( \11524 , \9819 , \1734 );
not \U$11182 ( \11525 , \9819 );
and \U$11183 ( \11526 , \11525 , RIbb2f340_7);
or \U$11184 ( \11527 , \11524 , \11526 );
nand \U$11185 ( \11528 , \11527 , \1702 );
nand \U$11186 ( \11529 , \11523 , \11528 );
not \U$11187 ( \11530 , \11529 );
not \U$11188 ( \11531 , \1570 );
not \U$11189 ( \11532 , \11222 );
or \U$11190 ( \11533 , \11531 , \11532 );
buf \U$11191 ( \11534 , \6937 );
not \U$11192 ( \11535 , \11534 );
and \U$11193 ( \11536 , \11535 , RIbb2f250_9);
not \U$11194 ( \11537 , \11535 );
and \U$11195 ( \11538 , \11537 , \1554 );
or \U$11196 ( \11539 , \11536 , \11538 );
nand \U$11197 ( \11540 , \11539 , \1533 );
nand \U$11198 ( \11541 , \11533 , \11540 );
not \U$11199 ( \11542 , \11541 );
or \U$11200 ( \11543 , \11530 , \11542 );
not \U$11201 ( \11544 , \11541 );
not \U$11202 ( \11545 , \11544 );
not \U$11203 ( \11546 , \11529 );
not \U$11204 ( \11547 , \11546 );
or \U$11205 ( \11548 , \11545 , \11547 );
not \U$11206 ( \11549 , \1077 );
not \U$11207 ( \11550 , \11184 );
or \U$11208 ( \11551 , \11549 , \11550 );
not \U$11209 ( \11552 , RIbb2f160_11);
not \U$11210 ( \11553 , \5956 );
or \U$11211 ( \11554 , \11552 , \11553 );
nand \U$11212 ( \11555 , \5955 , \1043 );
nand \U$11213 ( \11556 , \11554 , \11555 );
nand \U$11214 ( \11557 , \11556 , \1011 );
nand \U$11215 ( \11558 , \11551 , \11557 );
nand \U$11216 ( \11559 , \11548 , \11558 );
nand \U$11217 ( \11560 , \11543 , \11559 );
and \U$11218 ( \11561 , \11520 , \11560 );
and \U$11219 ( \11562 , \11509 , \11519 );
or \U$11220 ( \11563 , \11561 , \11562 );
nand \U$11221 ( \11564 , \11499 , \11563 );
nand \U$11222 ( \11565 , \11495 , \11564 );
xor \U$11223 ( \11566 , \11483 , \11565 );
not \U$11224 ( \11567 , \596 );
not \U$11225 ( \11568 , \4361 );
or \U$11226 ( \11569 , \11567 , \11568 );
nand \U$11227 ( \11570 , RIbb2c208_112, RIbb32bf8_176);
nand \U$11228 ( \11571 , \11569 , \11570 );
nand \U$11229 ( \11572 , \595 , \540 );
not \U$11230 ( \11573 , \11572 );
and \U$11231 ( \11574 , \11571 , \11573 );
not \U$11232 ( \11575 , \11571 );
and \U$11233 ( \11576 , \11575 , \11572 );
nor \U$11234 ( \11577 , \11574 , \11576 );
buf \U$11235 ( \11578 , \11577 );
not \U$11236 ( \11579 , \11578 );
buf \U$11237 ( \11580 , \11579 );
not \U$11238 ( \11581 , \11580 );
and \U$11239 ( \11582 , \1313 , \11581 );
not \U$11240 ( \11583 , \1429 );
xor \U$11241 ( \11584 , \1394 , \11145 );
not \U$11242 ( \11585 , \11584 );
or \U$11243 ( \11586 , \11583 , \11585 );
nand \U$11244 ( \11587 , \11148 , \1376 );
nand \U$11245 ( \11588 , \11586 , \11587 );
or \U$11246 ( \11589 , \11582 , \11588 );
not \U$11247 ( \11590 , \4791 );
not \U$11248 ( \11591 , \11298 );
or \U$11249 ( \11592 , \11590 , \11591 );
not \U$11250 ( \11593 , RIbb2e710_33);
not \U$11251 ( \11594 , \3290 );
or \U$11252 ( \11595 , \11593 , \11594 );
nand \U$11253 ( \11596 , \1283 , \3877 );
nand \U$11254 ( \11597 , \11595 , \11596 );
nand \U$11255 ( \11598 , \11597 , \3887 );
nand \U$11256 ( \11599 , \11592 , \11598 );
nand \U$11257 ( \11600 , \11589 , \11599 );
nand \U$11258 ( \11601 , \11588 , \11582 );
nand \U$11259 ( \11602 , \11600 , \11601 );
not \U$11260 ( \11603 , \11602 );
not \U$11261 ( \11604 , \10119 );
not \U$11262 ( \11605 , \11067 );
or \U$11263 ( \11606 , \11604 , \11605 );
not \U$11264 ( \11607 , RIbb2e170_45);
not \U$11265 ( \11608 , \3262 );
or \U$11266 ( \11609 , \11607 , \11608 );
nand \U$11267 ( \11610 , \3261 , \9094 );
nand \U$11268 ( \11611 , \11609 , \11610 );
nand \U$11269 ( \11612 , \11611 , \10117 );
nand \U$11270 ( \11613 , \11606 , \11612 );
not \U$11271 ( \11614 , \1517 );
not \U$11272 ( \11615 , \11320 );
or \U$11273 ( \11616 , \11614 , \11615 );
and \U$11274 ( \11617 , RIbb2ef80_15, \4088 );
not \U$11275 ( \11618 , RIbb2ef80_15);
and \U$11276 ( \11619 , \11618 , \4324 );
or \U$11277 ( \11620 , \11617 , \11619 );
nand \U$11278 ( \11621 , \11620 , \1445 );
nand \U$11279 ( \11622 , \11616 , \11621 );
xor \U$11280 ( \11623 , \11613 , \11622 );
not \U$11281 ( \11624 , \836 );
not \U$11282 ( \11625 , \11310 );
or \U$11283 ( \11626 , \11624 , \11625 );
not \U$11284 ( \11627 , RIbb2ee90_17);
not \U$11285 ( \11628 , \3276 );
or \U$11286 ( \11629 , \11627 , \11628 );
nand \U$11287 ( \11630 , \3275 , \3699 );
nand \U$11288 ( \11631 , \11629 , \11630 );
nand \U$11289 ( \11632 , \11631 , \832 );
nand \U$11290 ( \11633 , \11626 , \11632 );
and \U$11291 ( \11634 , \11623 , \11633 );
and \U$11292 ( \11635 , \11613 , \11622 );
or \U$11293 ( \11636 , \11634 , \11635 );
not \U$11294 ( \11637 , \11636 );
or \U$11295 ( \11638 , \11603 , \11637 );
or \U$11296 ( \11639 , \11636 , \11602 );
xor \U$11297 ( \11640 , \11213 , \11224 );
xor \U$11298 ( \11641 , \11640 , \11237 );
nand \U$11299 ( \11642 , \11639 , \11641 );
nand \U$11300 ( \11643 , \11638 , \11642 );
xor \U$11301 ( \11644 , \11146 , \11152 );
xor \U$11302 ( \11645 , \11644 , \11163 );
xor \U$11303 ( \11646 , \11179 , \11188 );
xor \U$11304 ( \11647 , \11646 , \11199 );
xor \U$11305 ( \11648 , \11645 , \11647 );
not \U$11306 ( \11649 , \5845 );
not \U$11307 ( \11650 , \11340 );
or \U$11308 ( \11651 , \11649 , \11650 );
not \U$11309 ( \11652 , RIbb2e620_35);
not \U$11310 ( \11653 , \5988 );
or \U$11311 ( \11654 , \11652 , \11653 );
nand \U$11312 ( \11655 , \3053 , \6688 );
nand \U$11313 ( \11656 , \11654 , \11655 );
nand \U$11314 ( \11657 , \11656 , \4712 );
nand \U$11315 ( \11658 , \11651 , \11657 );
not \U$11316 ( \11659 , \2078 );
not \U$11317 ( \11660 , \11364 );
or \U$11318 ( \11661 , \11659 , \11660 );
not \U$11319 ( \11662 , RIbb2ecb0_21);
not \U$11320 ( \11663 , \3226 );
or \U$11321 ( \11664 , \11662 , \11663 );
nand \U$11322 ( \11665 , \3228 , \849 );
nand \U$11323 ( \11666 , \11664 , \11665 );
nand \U$11324 ( \11667 , \11666 , \2077 );
nand \U$11325 ( \11668 , \11661 , \11667 );
xor \U$11326 ( \11669 , \11658 , \11668 );
not \U$11327 ( \11670 , \853 );
not \U$11328 ( \11671 , RIbb2eda0_19);
not \U$11329 ( \11672 , \10096 );
or \U$11330 ( \11673 , \11671 , \11672 );
nand \U$11331 ( \11674 , \10095 , \1776 );
nand \U$11332 ( \11675 , \11673 , \11674 );
not \U$11333 ( \11676 , \11675 );
or \U$11334 ( \11677 , \11670 , \11676 );
nand \U$11335 ( \11678 , \11517 , \855 );
nand \U$11336 ( \11679 , \11677 , \11678 );
and \U$11337 ( \11680 , \11669 , \11679 );
and \U$11338 ( \11681 , \11658 , \11668 );
or \U$11339 ( \11682 , \11680 , \11681 );
and \U$11340 ( \11683 , \11648 , \11682 );
and \U$11341 ( \11684 , \11645 , \11647 );
or \U$11342 ( \11685 , \11683 , \11684 );
xor \U$11343 ( \11686 , \11643 , \11685 );
not \U$11344 ( \11687 , \11176 );
not \U$11345 ( \11688 , RIbb2e080_47);
not \U$11346 ( \11689 , \813 );
or \U$11347 ( \11690 , \11688 , \11689 );
nand \U$11348 ( \11691 , \10604 , \10113 );
nand \U$11349 ( \11692 , \11690 , \11691 );
not \U$11350 ( \11693 , \11692 );
or \U$11351 ( \11694 , \11687 , \11693 );
nand \U$11352 ( \11695 , \11177 , RIbb2e080_47);
nand \U$11353 ( \11696 , \11694 , \11695 );
not \U$11354 ( \11697 , \1147 );
not \U$11355 ( \11698 , \11211 );
or \U$11356 ( \11699 , \11697 , \11698 );
not \U$11357 ( \11700 , \9860 );
and \U$11358 ( \11701 , \11700 , RIbb2f430_5);
not \U$11359 ( \11702 , \11700 );
and \U$11360 ( \11703 , \11702 , \1647 );
or \U$11361 ( \11704 , \11701 , \11703 );
nand \U$11362 ( \11705 , \11704 , \1090 );
nand \U$11363 ( \11706 , \11699 , \11705 );
xor \U$11364 ( \11707 , \11696 , \11706 );
not \U$11365 ( \11708 , \1294 );
not \U$11366 ( \11709 , \11159 );
or \U$11367 ( \11710 , \11708 , \11709 );
and \U$11368 ( \11711 , \10301 , \1245 );
not \U$11369 ( \11712 , \10301 );
and \U$11370 ( \11713 , \11712 , \1246 );
or \U$11371 ( \11714 , \11711 , \11713 );
nand \U$11372 ( \11715 , \11714 , \1265 );
nand \U$11373 ( \11716 , \11710 , \11715 );
and \U$11374 ( \11717 , \11707 , \11716 );
and \U$11375 ( \11718 , \11696 , \11706 );
or \U$11376 ( \11719 , \11717 , \11718 );
not \U$11377 ( \11720 , \8450 );
not \U$11378 ( \11721 , \11258 );
or \U$11379 ( \11722 , \11720 , \11721 );
and \U$11380 ( \11723 , RIbb2e440_39, \1550 );
not \U$11381 ( \11724 , RIbb2e440_39);
and \U$11382 ( \11725 , \11724 , \1548 );
or \U$11383 ( \11726 , \11723 , \11725 );
nand \U$11384 ( \11727 , \11726 , \8445 );
nand \U$11385 ( \11728 , \11722 , \11727 );
not \U$11386 ( \11729 , \10451 );
not \U$11387 ( \11730 , \11386 );
or \U$11388 ( \11731 , \11729 , \11730 );
not \U$11389 ( \11732 , RIbb2e260_43);
not \U$11390 ( \11733 , \988 );
or \U$11391 ( \11734 , \11732 , \11733 );
nand \U$11392 ( \11735 , \987 , \10444 );
nand \U$11393 ( \11736 , \11734 , \11735 );
nand \U$11394 ( \11737 , \11736 , \10449 );
nand \U$11395 ( \11738 , \11731 , \11737 );
xor \U$11396 ( \11739 , \11728 , \11738 );
not \U$11397 ( \11740 , \3445 );
not \U$11398 ( \11741 , RIbb2e9e0_27);
not \U$11399 ( \11742 , \3310 );
or \U$11400 ( \11743 , \11741 , \11742 );
nand \U$11401 ( \11744 , \4450 , \3454 );
nand \U$11402 ( \11745 , \11743 , \11744 );
not \U$11403 ( \11746 , \11745 );
or \U$11404 ( \11747 , \11740 , \11746 );
nand \U$11405 ( \11748 , \11286 , \3465 );
nand \U$11406 ( \11749 , \11747 , \11748 );
and \U$11407 ( \11750 , \11739 , \11749 );
and \U$11408 ( \11751 , \11728 , \11738 );
or \U$11409 ( \11752 , \11750 , \11751 );
xor \U$11410 ( \11753 , \11719 , \11752 );
not \U$11411 ( \11754 , \2963 );
not \U$11412 ( \11755 , \11396 );
or \U$11413 ( \11756 , \11754 , \11755 );
and \U$11414 ( \11757 , RIbb2ead0_25, \3520 );
not \U$11415 ( \11758 , RIbb2ead0_25);
and \U$11416 ( \11759 , \11758 , \3343 );
or \U$11417 ( \11760 , \11757 , \11759 );
nand \U$11418 ( \11761 , \11760 , \2980 );
nand \U$11419 ( \11762 , \11756 , \11761 );
not \U$11420 ( \11763 , \6242 );
not \U$11421 ( \11764 , \11374 );
or \U$11422 ( \11765 , \11763 , \11764 );
not \U$11423 ( \11766 , RIbb2e530_37);
not \U$11424 ( \11767 , \1689 );
or \U$11425 ( \11768 , \11766 , \11767 );
nand \U$11426 ( \11769 , \3552 , \7243 );
nand \U$11427 ( \11770 , \11768 , \11769 );
nand \U$11428 ( \11771 , \11770 , \6251 );
nand \U$11429 ( \11772 , \11765 , \11771 );
xor \U$11430 ( \11773 , \11762 , \11772 );
not \U$11431 ( \11774 , \3383 );
not \U$11432 ( \11775 , \11351 );
or \U$11433 ( \11776 , \11774 , \11775 );
not \U$11434 ( \11777 , RIbb2ebc0_23);
not \U$11435 ( \11778 , \6301 );
or \U$11436 ( \11779 , \11777 , \11778 );
nand \U$11437 ( \11780 , \3620 , \3401 );
nand \U$11438 ( \11781 , \11779 , \11780 );
nand \U$11439 ( \11782 , \11781 , \3407 );
nand \U$11440 ( \11783 , \11776 , \11782 );
and \U$11441 ( \11784 , \11773 , \11783 );
and \U$11442 ( \11785 , \11762 , \11772 );
or \U$11443 ( \11786 , \11784 , \11785 );
and \U$11444 ( \11787 , \11753 , \11786 );
and \U$11445 ( \11788 , \11719 , \11752 );
or \U$11446 ( \11789 , \11787 , \11788 );
and \U$11447 ( \11790 , \11686 , \11789 );
and \U$11448 ( \11791 , \11643 , \11685 );
or \U$11449 ( \11792 , \11790 , \11791 );
and \U$11450 ( \11793 , \11566 , \11792 );
and \U$11451 ( \11794 , \11483 , \11565 );
or \U$11452 ( \11795 , \11793 , \11794 );
not \U$11453 ( \11796 , \11795 );
and \U$11454 ( \11797 , \11118 , \11042 );
not \U$11455 ( \11798 , \11118 );
and \U$11456 ( \11799 , \11798 , \11043 );
or \U$11457 ( \11800 , \11797 , \11799 );
xor \U$11458 ( \11801 , \11800 , \11039 );
not \U$11459 ( \11802 , \11801 );
or \U$11460 ( \11803 , \11796 , \11802 );
or \U$11461 ( \11804 , \11801 , \11795 );
xor \U$11462 ( \11805 , \11251 , \11328 );
xor \U$11463 ( \11806 , \11805 , \11404 );
not \U$11464 ( \11807 , \8995 );
not \U$11465 ( \11808 , \11080 );
or \U$11466 ( \11809 , \11807 , \11808 );
not \U$11467 ( \11810 , RIbb2e350_41);
not \U$11468 ( \11811 , \4284 );
or \U$11469 ( \11812 , \11810 , \11811 );
nand \U$11470 ( \11813 , \3099 , \7097 );
nand \U$11471 ( \11814 , \11812 , \11813 );
nand \U$11472 ( \11815 , \11814 , \8362 );
nand \U$11473 ( \11816 , \11809 , \11815 );
not \U$11474 ( \11817 , \2922 );
not \U$11475 ( \11818 , RIbb2e8f0_29);
not \U$11476 ( \11819 , \3575 );
or \U$11477 ( \11820 , \11818 , \11819 );
nand \U$11478 ( \11821 , \1339 , \3800 );
nand \U$11479 ( \11822 , \11820 , \11821 );
not \U$11480 ( \11823 , \11822 );
or \U$11481 ( \11824 , \11817 , \11823 );
nand \U$11482 ( \11825 , \11272 , \2925 );
nand \U$11483 ( \11826 , \11824 , \11825 );
xor \U$11484 ( \11827 , \11816 , \11826 );
not \U$11485 ( \11828 , \2941 );
not \U$11486 ( \11829 , \11058 );
or \U$11487 ( \11830 , \11828 , \11829 );
and \U$11488 ( \11831 , RIbb2e800_31, \1387 );
not \U$11489 ( \11832 , RIbb2e800_31);
and \U$11490 ( \11833 , \11832 , \4341 );
nor \U$11491 ( \11834 , \11831 , \11833 );
nand \U$11492 ( \11835 , \11834 , \2940 );
nand \U$11493 ( \11836 , \11830 , \11835 );
and \U$11494 ( \11837 , \11827 , \11836 );
and \U$11495 ( \11838 , \11816 , \11826 );
or \U$11496 ( \11839 , \11837 , \11838 );
xor \U$11497 ( \11840 , \11378 , \11388 );
xor \U$11498 ( \11841 , \11840 , \11398 );
xor \U$11499 ( \11842 , \11839 , \11841 );
xor \U$11500 ( \11843 , \11366 , \11353 );
xor \U$11501 ( \11844 , \11843 , \11342 );
and \U$11502 ( \11845 , \11842 , \11844 );
and \U$11503 ( \11846 , \11839 , \11841 );
or \U$11504 ( \11847 , \11845 , \11846 );
xor \U$11505 ( \11848 , \11253 , \11291 );
xor \U$11506 ( \11849 , \11848 , \11325 );
xor \U$11507 ( \11850 , \11847 , \11849 );
xor \U$11508 ( \11851 , \11288 , \11263 );
xnor \U$11509 ( \11852 , \11851 , \11275 );
not \U$11510 ( \11853 , \11852 );
xor \U$11511 ( \11854 , \11060 , \11071 );
xor \U$11512 ( \11855 , \11854 , \11082 );
buf \U$11513 ( \11856 , \11855 );
or \U$11514 ( \11857 , \11853 , \11856 );
xor \U$11515 ( \11858 , \11302 , \11312 );
xor \U$11516 ( \11859 , \11858 , \11322 );
nand \U$11517 ( \11860 , \11857 , \11859 );
nand \U$11518 ( \11861 , \11853 , \11856 );
nand \U$11519 ( \11862 , \11860 , \11861 );
and \U$11520 ( \11863 , \11850 , \11862 );
and \U$11521 ( \11864 , \11847 , \11849 );
or \U$11522 ( \11865 , \11863 , \11864 );
xor \U$11523 ( \11866 , \11806 , \11865 );
not \U$11524 ( \11867 , \11093 );
not \U$11525 ( \11868 , \11096 );
or \U$11526 ( \11869 , \11867 , \11868 );
or \U$11527 ( \11870 , \11096 , \11093 );
nand \U$11528 ( \11871 , \11869 , \11870 );
and \U$11529 ( \11872 , \11871 , \11116 );
not \U$11530 ( \11873 , \11871 );
not \U$11531 ( \11874 , \11116 );
and \U$11532 ( \11875 , \11873 , \11874 );
nor \U$11533 ( \11876 , \11872 , \11875 );
and \U$11534 ( \11877 , \11866 , \11876 );
and \U$11535 ( \11878 , \11806 , \11865 );
or \U$11536 ( \11879 , \11877 , \11878 );
nand \U$11537 ( \11880 , \11804 , \11879 );
nand \U$11538 ( \11881 , \11803 , \11880 );
not \U$11539 ( \11882 , \11479 );
not \U$11540 ( \11883 , \11468 );
nand \U$11541 ( \11884 , \11882 , \11883 );
nand \U$11542 ( \11885 , \11881 , \11884 );
nand \U$11543 ( \11886 , \11481 , \11885 );
nand \U$11544 ( \11887 , \11440 , \11886 );
nand \U$11545 ( \11888 , \11437 , \11439 );
nand \U$11546 ( \11889 , \11887 , \11888 );
not \U$11547 ( \11890 , \11889 );
nand \U$11548 ( \11891 , \11431 , \11890 );
and \U$11549 ( \11892 , \11428 , \11891 );
xor \U$11550 ( \11893 , \10010 , \10518 );
and \U$11551 ( \11894 , \11893 , \10808 );
and \U$11552 ( \11895 , \10010 , \10518 );
or \U$11553 ( \11896 , \11894 , \11895 );
not \U$11554 ( \11897 , \9776 );
not \U$11555 ( \11898 , \10009 );
or \U$11556 ( \11899 , \11897 , \11898 );
or \U$11557 ( \11900 , \9776 , \10009 );
nand \U$11558 ( \11901 , \11900 , \10006 );
nand \U$11559 ( \11902 , \11899 , \11901 );
not \U$11560 ( \11903 , \11902 );
xor \U$11561 ( \11904 , \9155 , \9224 );
xor \U$11562 ( \11905 , \11904 , \9488 );
not \U$11563 ( \11906 , \11905 );
not \U$11564 ( \11907 , \11906 );
or \U$11565 ( \11908 , \11903 , \11907 );
not \U$11566 ( \11909 , \11902 );
nand \U$11567 ( \11910 , \11905 , \11909 );
nand \U$11568 ( \11911 , \11908 , \11910 );
not \U$11569 ( \11912 , \10079 );
not \U$11570 ( \11913 , \10087 );
or \U$11571 ( \11914 , \11912 , \11913 );
not \U$11572 ( \11915 , \10080 );
not \U$11573 ( \11916 , \10086 );
or \U$11574 ( \11917 , \11915 , \11916 );
nand \U$11575 ( \11918 , \11917 , \10514 );
nand \U$11576 ( \11919 , \11914 , \11918 );
not \U$11577 ( \11920 , \11919 );
and \U$11578 ( \11921 , \11911 , \11920 );
not \U$11579 ( \11922 , \11911 );
and \U$11580 ( \11923 , \11922 , \11919 );
nor \U$11581 ( \11924 , \11921 , \11923 );
nand \U$11582 ( \11925 , \11896 , \11924 );
not \U$11583 ( \11926 , \11925 );
xor \U$11584 ( \11927 , \8796 , \9491 );
xor \U$11585 ( \11928 , \11927 , \9525 );
not \U$11586 ( \11929 , \11909 );
not \U$11587 ( \11930 , \11906 );
or \U$11588 ( \11931 , \11929 , \11930 );
nand \U$11589 ( \11932 , \11931 , \11919 );
nand \U$11590 ( \11933 , \11905 , \11902 );
nand \U$11591 ( \11934 , \11932 , \11933 );
nor \U$11592 ( \11935 , \11928 , \11934 );
nor \U$11593 ( \11936 , \11926 , \11935 );
not \U$11594 ( \11937 , \9647 );
not \U$11595 ( \11938 , \9659 );
or \U$11596 ( \11939 , \11937 , \11938 );
nand \U$11597 ( \11940 , \11939 , \9672 );
nand \U$11598 ( \11941 , \9660 , \9646 );
nand \U$11599 ( \11942 , \11940 , \11941 );
not \U$11600 ( \11943 , \11942 );
xor \U$11601 ( \11944 , \7526 , \7514 );
xnor \U$11602 ( \11945 , \11944 , \7529 );
nand \U$11603 ( \11946 , \11943 , \11945 );
and \U$11604 ( \11947 , \9675 , \11892 , \11936 , \11946 );
not \U$11605 ( \11948 , \11176 );
not \U$11606 ( \11949 , RIbb2e080_47);
not \U$11607 ( \11950 , \1475 );
or \U$11608 ( \11951 , \11949 , \11950 );
nand \U$11609 ( \11952 , \4558 , \10113 );
nand \U$11610 ( \11953 , \11951 , \11952 );
not \U$11611 ( \11954 , \11953 );
or \U$11612 ( \11955 , \11948 , \11954 );
not \U$11613 ( \11956 , RIbb2e080_47);
not \U$11614 ( \11957 , \3262 );
or \U$11615 ( \11958 , \11956 , \11957 );
not \U$11616 ( \11959 , RIbb2e080_47);
nand \U$11617 ( \11960 , \3261 , \11959 );
nand \U$11618 ( \11961 , \11958 , \11960 );
nand \U$11619 ( \11962 , \11961 , \11177 );
nand \U$11620 ( \11963 , \11955 , \11962 );
not \U$11621 ( \11964 , \2940 );
not \U$11622 ( \11965 , RIbb2e800_31);
not \U$11623 ( \11966 , \4609 );
or \U$11624 ( \11967 , \11965 , \11966 );
nand \U$11625 ( \11968 , \1852 , \8810 );
nand \U$11626 ( \11969 , \11967 , \11968 );
not \U$11627 ( \11970 , \11969 );
or \U$11628 ( \11971 , \11964 , \11970 );
not \U$11629 ( \11972 , RIbb2e800_31);
not \U$11630 ( \11973 , \6097 );
or \U$11631 ( \11974 , \11972 , \11973 );
not \U$11632 ( \11975 , RIbb2e800_31);
nand \U$11633 ( \11976 , \1339 , \11975 );
nand \U$11634 ( \11977 , \11974 , \11976 );
nand \U$11635 ( \11978 , \11977 , \3613 );
nand \U$11636 ( \11979 , \11971 , \11978 );
or \U$11637 ( \11980 , \11963 , \11979 );
not \U$11638 ( \11981 , \10449 );
not \U$11639 ( \11982 , RIbb2e260_43);
not \U$11640 ( \11983 , \4595 );
or \U$11641 ( \11984 , \11982 , \11983 );
nand \U$11642 ( \11985 , \1561 , \10444 );
nand \U$11643 ( \11986 , \11984 , \11985 );
not \U$11644 ( \11987 , \11986 );
or \U$11645 ( \11988 , \11981 , \11987 );
not \U$11646 ( \11989 , RIbb2e260_43);
not \U$11647 ( \11990 , \1070 );
or \U$11648 ( \11991 , \11989 , \11990 );
nand \U$11649 ( \11992 , \1071 , \8347 );
nand \U$11650 ( \11993 , \11991 , \11992 );
nand \U$11651 ( \11994 , \11993 , \10451 );
nand \U$11652 ( \11995 , \11988 , \11994 );
nand \U$11653 ( \11996 , \11980 , \11995 );
nand \U$11654 ( \11997 , \11979 , \11963 );
nand \U$11655 ( \11998 , \11996 , \11997 );
not \U$11656 ( \11999 , \10599 );
not \U$11657 ( \12000 , RIbb2e170_45);
not \U$11658 ( \12001 , \10421 );
or \U$11659 ( \12002 , \12000 , \12001 );
not \U$11660 ( \12003 , RIbb2e170_45);
nand \U$11661 ( \12004 , \952 , \12003 );
nand \U$11662 ( \12005 , \12002 , \12004 );
not \U$11663 ( \12006 , \12005 );
or \U$11664 ( \12007 , \11999 , \12006 );
not \U$11665 ( \12008 , RIbb2e170_45);
not \U$11666 ( \12009 , \992 );
or \U$11667 ( \12010 , \12008 , \12009 );
nand \U$11668 ( \12011 , \987 , \12003 );
nand \U$11669 ( \12012 , \12010 , \12011 );
nand \U$11670 ( \12013 , \12012 , \10119 );
nand \U$11671 ( \12014 , \12007 , \12013 );
not \U$11672 ( \12015 , \3887 );
not \U$11673 ( \12016 , RIbb2e710_33);
not \U$11674 ( \12017 , \1420 );
or \U$11675 ( \12018 , \12016 , \12017 );
not \U$11676 ( \12019 , RIbb2e710_33);
nand \U$11677 ( \12020 , \1421 , \12019 );
nand \U$11678 ( \12021 , \12018 , \12020 );
not \U$11679 ( \12022 , \12021 );
or \U$11680 ( \12023 , \12015 , \12022 );
buf \U$11681 ( \12024 , \1385 );
and \U$11682 ( \12025 , \12024 , RIbb2e710_33);
not \U$11683 ( \12026 , \12024 );
and \U$11684 ( \12027 , \12026 , \3877 );
or \U$11685 ( \12028 , \12025 , \12027 );
nand \U$11686 ( \12029 , \12028 , \4791 );
nand \U$11687 ( \12030 , \12023 , \12029 );
xor \U$11688 ( \12031 , \12014 , \12030 );
not \U$11689 ( \12032 , \5845 );
not \U$11690 ( \12033 , RIbb2e620_35);
not \U$11691 ( \12034 , \1284 );
or \U$11692 ( \12035 , \12033 , \12034 );
buf \U$11693 ( \12036 , \1280 );
not \U$11694 ( \12037 , \12036 );
not \U$11695 ( \12038 , \12037 );
nand \U$11696 ( \12039 , \12038 , \6002 );
nand \U$11697 ( \12040 , \12035 , \12039 );
not \U$11698 ( \12041 , \12040 );
or \U$11699 ( \12042 , \12032 , \12041 );
not \U$11700 ( \12043 , RIbb2e620_35);
not \U$11701 ( \12044 , \1170 );
or \U$11702 ( \12045 , \12043 , \12044 );
not \U$11703 ( \12046 , \3990 );
nand \U$11704 ( \12047 , \12046 , \11338 );
nand \U$11705 ( \12048 , \12045 , \12047 );
nand \U$11706 ( \12049 , \12048 , \4712 );
nand \U$11707 ( \12050 , \12042 , \12049 );
and \U$11708 ( \12051 , \12031 , \12050 );
and \U$11709 ( \12052 , \12014 , \12030 );
or \U$11710 ( \12053 , \12051 , \12052 );
or \U$11711 ( \12054 , \11998 , \12053 );
not \U$11712 ( \12055 , \2922 );
not \U$11713 ( \12056 , RIbb2e8f0_29);
not \U$11714 ( \12057 , \3319 );
or \U$11715 ( \12058 , \12056 , \12057 );
nand \U$11716 ( \12059 , \2225 , \4800 );
nand \U$11717 ( \12060 , \12058 , \12059 );
not \U$11718 ( \12061 , \12060 );
or \U$11719 ( \12062 , \12055 , \12061 );
not \U$11720 ( \12063 , RIbb2e8f0_29);
not \U$11721 ( \12064 , \4449 );
or \U$11722 ( \12065 , \12063 , \12064 );
nand \U$11723 ( \12066 , \4450 , \2949 );
nand \U$11724 ( \12067 , \12065 , \12066 );
nand \U$11725 ( \12068 , \12067 , \2925 );
nand \U$11726 ( \12069 , \12062 , \12068 );
not \U$11727 ( \12070 , \8362 );
not \U$11728 ( \12071 , RIbb2e350_41);
not \U$11729 ( \12072 , \5130 );
or \U$11730 ( \12073 , \12071 , \12072 );
nand \U$11731 ( \12074 , \3480 , \8357 );
nand \U$11732 ( \12075 , \12073 , \12074 );
not \U$11733 ( \12076 , \12075 );
or \U$11734 ( \12077 , \12070 , \12076 );
not \U$11735 ( \12078 , RIbb2e350_41);
not \U$11736 ( \12079 , \1549 );
or \U$11737 ( \12080 , \12078 , \12079 );
nand \U$11738 ( \12081 , \1548 , \7097 );
nand \U$11739 ( \12082 , \12080 , \12081 );
nand \U$11740 ( \12083 , \12082 , \8995 );
nand \U$11741 ( \12084 , \12077 , \12083 );
or \U$11742 ( \12085 , \12069 , \12084 );
not \U$11743 ( \12086 , \12085 );
not \U$11744 ( \12087 , \3445 );
not \U$11745 ( \12088 , RIbb2e9e0_27);
not \U$11746 ( \12089 , \4219 );
or \U$11747 ( \12090 , \12088 , \12089 );
nand \U$11748 ( \12091 , \3167 , \3454 );
nand \U$11749 ( \12092 , \12090 , \12091 );
not \U$11750 ( \12093 , \12092 );
or \U$11751 ( \12094 , \12087 , \12093 );
not \U$11752 ( \12095 , RIbb2e9e0_27);
buf \U$11753 ( \12096 , \3341 );
not \U$11754 ( \12097 , \12096 );
not \U$11755 ( \12098 , \12097 );
or \U$11756 ( \12099 , \12095 , \12098 );
nand \U$11757 ( \12100 , \3521 , \3454 );
nand \U$11758 ( \12101 , \12099 , \12100 );
nand \U$11759 ( \12102 , \12101 , \3465 );
nand \U$11760 ( \12103 , \12094 , \12102 );
not \U$11761 ( \12104 , \12103 );
or \U$11762 ( \12105 , \12086 , \12104 );
nand \U$11763 ( \12106 , \12069 , \12084 );
nand \U$11764 ( \12107 , \12105 , \12106 );
nand \U$11765 ( \12108 , \12054 , \12107 );
not \U$11766 ( \12109 , \11998 );
not \U$11767 ( \12110 , \12109 );
nand \U$11768 ( \12111 , \12110 , \12053 );
nand \U$11769 ( \12112 , \12108 , \12111 );
not \U$11770 ( \12113 , \998 );
not \U$11771 ( \12114 , RIbb2f070_13);
not \U$11772 ( \12115 , \6231 );
or \U$11773 ( \12116 , \12114 , \12115 );
nand \U$11774 ( \12117 , \6232 , \3421 );
nand \U$11775 ( \12118 , \12116 , \12117 );
not \U$11776 ( \12119 , \12118 );
or \U$11777 ( \12120 , \12113 , \12119 );
not \U$11778 ( \12121 , RIbb2f070_13);
not \U$11779 ( \12122 , \10577 );
or \U$11780 ( \12123 , \12121 , \12122 );
nand \U$11781 ( \12124 , \5957 , \906 );
nand \U$11782 ( \12125 , \12123 , \12124 );
nand \U$11783 ( \12126 , \12125 , \916 );
nand \U$11784 ( \12127 , \12120 , \12126 );
not \U$11785 ( \12128 , \12127 );
not \U$11786 ( \12129 , \1011 );
not \U$11787 ( \12130 , RIbb2f160_11);
not \U$11788 ( \12131 , \11535 );
or \U$11789 ( \12132 , \12130 , \12131 );
nand \U$11790 ( \12133 , \6939 , \1805 );
nand \U$11791 ( \12134 , \12132 , \12133 );
not \U$11792 ( \12135 , \12134 );
or \U$11793 ( \12136 , \12129 , \12135 );
not \U$11794 ( \12137 , RIbb2f160_11);
not \U$11795 ( \12138 , \11218 );
or \U$11796 ( \12139 , \12137 , \12138 );
nand \U$11797 ( \12140 , \8339 , \1805 );
nand \U$11798 ( \12141 , \12139 , \12140 );
nand \U$11799 ( \12142 , \12141 , \1077 );
nand \U$11800 ( \12143 , \12136 , \12142 );
not \U$11801 ( \12144 , \12143 );
or \U$11802 ( \12145 , \12128 , \12144 );
or \U$11803 ( \12146 , \12143 , \12127 );
not \U$11804 ( \12147 , \1445 );
and \U$11805 ( \12148 , RIbb2ef80_15, \10556 );
not \U$11806 ( \12149 , RIbb2ef80_15);
and \U$11807 ( \12150 , \12149 , \6202 );
or \U$11808 ( \12151 , \12148 , \12150 );
not \U$11809 ( \12152 , \12151 );
or \U$11810 ( \12153 , \12147 , \12152 );
not \U$11811 ( \12154 , \8375 );
and \U$11812 ( \12155 , RIbb2ef80_15, \12154 );
not \U$11813 ( \12156 , RIbb2ef80_15);
and \U$11814 ( \12157 , \12156 , \8375 );
or \U$11815 ( \12158 , \12155 , \12157 );
nand \U$11816 ( \12159 , \12158 , \1517 );
nand \U$11817 ( \12160 , \12153 , \12159 );
nand \U$11818 ( \12161 , \12146 , \12160 );
nand \U$11819 ( \12162 , \12145 , \12161 );
and \U$11820 ( \12163 , RIbb2df90_49, RIbb2df18_50);
xor \U$11821 ( \12164 , RIbb2dea0_51, RIbb2df18_50);
nor \U$11822 ( \12165 , RIbb2df90_49, RIbb2df18_50);
nor \U$11823 ( \12166 , \12163 , \12164 , \12165 );
buf \U$11824 ( \12167 , \12166 );
buf \U$11825 ( \12168 , \12164 );
buf \U$11826 ( \12169 , \12168 );
or \U$11827 ( \12170 , \12167 , \12169 );
nand \U$11828 ( \12171 , \12170 , RIbb2df90_49);
nand \U$11829 ( \12172 , \596 , \11570 );
xnor \U$11830 ( \12173 , \12172 , \4361 );
buf \U$11831 ( \12174 , \12173 );
buf \U$11832 ( \12175 , \12174 );
and \U$11833 ( \12176 , \1393 , \12175 );
xor \U$11834 ( \12177 , \12171 , \12176 );
not \U$11835 ( \12178 , \1517 );
not \U$11836 ( \12179 , \11620 );
or \U$11837 ( \12180 , \12178 , \12179 );
nand \U$11838 ( \12181 , \12158 , \1445 );
nand \U$11839 ( \12182 , \12180 , \12181 );
xor \U$11840 ( \12183 , \12177 , \12182 );
xor \U$11841 ( \12184 , \12162 , \12183 );
not \U$11842 ( \12185 , \1702 );
not \U$11843 ( \12186 , RIbb2f340_7);
not \U$11844 ( \12187 , \9279 );
or \U$11845 ( \12188 , \12186 , \12187 );
nand \U$11846 ( \12189 , \9860 , \1692 );
nand \U$11847 ( \12190 , \12188 , \12189 );
not \U$11848 ( \12191 , \12190 );
or \U$11849 ( \12192 , \12185 , \12191 );
not \U$11850 ( \12193 , RIbb2f340_7);
not \U$11851 ( \12194 , \8631 );
not \U$11852 ( \12195 , \12194 );
or \U$11853 ( \12196 , \12193 , \12195 );
nand \U$11854 ( \12197 , \8631 , \2700 );
nand \U$11855 ( \12198 , \12196 , \12197 );
nand \U$11856 ( \12199 , \12198 , \1737 );
nand \U$11857 ( \12200 , \12192 , \12199 );
not \U$11858 ( \12201 , \1570 );
not \U$11859 ( \12202 , RIbb2f250_9);
not \U$11860 ( \12203 , \9071 );
or \U$11861 ( \12204 , \12202 , \12203 );
nand \U$11862 ( \12205 , \9074 , \1566 );
nand \U$11863 ( \12206 , \12204 , \12205 );
not \U$11864 ( \12207 , \12206 );
or \U$11865 ( \12208 , \12201 , \12207 );
not \U$11866 ( \12209 , RIbb2f250_9);
not \U$11867 ( \12210 , \8318 );
buf \U$11868 ( \12211 , \12210 );
not \U$11869 ( \12212 , \12211 );
or \U$11870 ( \12213 , \12209 , \12212 );
not \U$11871 ( \12214 , \12211 );
nand \U$11872 ( \12215 , \12214 , \1566 );
nand \U$11873 ( \12216 , \12213 , \12215 );
nand \U$11874 ( \12217 , \12216 , \1533 );
nand \U$11875 ( \12218 , \12208 , \12217 );
xor \U$11876 ( \12219 , \12200 , \12218 );
not \U$11877 ( \12220 , \1147 );
not \U$11878 ( \12221 , RIbb2f430_5);
not \U$11879 ( \12222 , \9841 );
not \U$11880 ( \12223 , \12222 );
or \U$11881 ( \12224 , \12221 , \12223 );
nand \U$11882 ( \12225 , \9841 , \1085 );
nand \U$11883 ( \12226 , \12224 , \12225 );
not \U$11884 ( \12227 , \12226 );
or \U$11885 ( \12228 , \12220 , \12227 );
not \U$11886 ( \12229 , RIbb2f430_5);
not \U$11887 ( \12230 , \10301 );
not \U$11888 ( \12231 , \12230 );
or \U$11889 ( \12232 , \12229 , \12231 );
not \U$11890 ( \12233 , \10300 );
buf \U$11891 ( \12234 , \12233 );
not \U$11892 ( \12235 , \12234 );
nand \U$11893 ( \12236 , \12235 , \1647 );
nand \U$11894 ( \12237 , \12232 , \12236 );
nand \U$11895 ( \12238 , \12237 , \1090 );
nand \U$11896 ( \12239 , \12228 , \12238 );
and \U$11897 ( \12240 , \12219 , \12239 );
and \U$11898 ( \12241 , \12200 , \12218 );
or \U$11899 ( \12242 , \12240 , \12241 );
xor \U$11900 ( \12243 , \12184 , \12242 );
xor \U$11901 ( \12244 , \12112 , \12243 );
xor \U$11902 ( \12245 , \12160 , \12143 );
xor \U$11903 ( \12246 , \12245 , \12127 );
not \U$11904 ( \12247 , \1294 );
not \U$11905 ( \12248 , \1246 );
not \U$11906 ( \12249 , \10764 );
not \U$11907 ( \12250 , \12249 );
or \U$11908 ( \12251 , \12248 , \12250 );
nand \U$11909 ( \12252 , \10764 , \1245 );
nand \U$11910 ( \12253 , \12251 , \12252 );
not \U$11911 ( \12254 , \12253 );
or \U$11912 ( \12255 , \12247 , \12254 );
not \U$11913 ( \12256 , \1288 );
not \U$11914 ( \12257 , \11142 );
not \U$11915 ( \12258 , \12257 );
or \U$11916 ( \12259 , \12256 , \12258 );
not \U$11917 ( \12260 , \11142 );
not \U$11918 ( \12261 , \12260 );
nand \U$11919 ( \12262 , \12261 , \1244 );
nand \U$11920 ( \12263 , \12259 , \12262 );
nand \U$11921 ( \12264 , \12263 , \1265 );
nand \U$11922 ( \12265 , \12255 , \12264 );
not \U$11923 ( \12266 , \1376 );
xor \U$11924 ( \12267 , \1313 , \11581 );
not \U$11925 ( \12268 , \12267 );
or \U$11926 ( \12269 , \12266 , \12268 );
xor \U$11927 ( \12270 , \1393 , \12175 );
nand \U$11928 ( \12271 , \12270 , \1430 );
nand \U$11929 ( \12272 , \12269 , \12271 );
xor \U$11930 ( \12273 , \12265 , \12272 );
not \U$11931 ( \12274 , \12167 );
not \U$11932 ( \12275 , RIbb2df90_49);
not \U$11933 ( \12276 , \813 );
or \U$11934 ( \12277 , \12275 , \12276 );
not \U$11935 ( \12278 , RIbb2df90_49);
nand \U$11936 ( \12279 , \10604 , \12278 );
nand \U$11937 ( \12280 , \12277 , \12279 );
not \U$11938 ( \12281 , \12280 );
or \U$11939 ( \12282 , \12274 , \12281 );
not \U$11940 ( \12283 , \12168 );
not \U$11941 ( \12284 , \12283 );
buf \U$11942 ( \12285 , \12284 );
nand \U$11943 ( \12286 , \12285 , RIbb2df90_49);
nand \U$11944 ( \12287 , \12282 , \12286 );
xor \U$11945 ( \12288 , \12273 , \12287 );
xor \U$11946 ( \12289 , \12246 , \12288 );
not \U$11947 ( \12290 , \1376 );
not \U$11948 ( \12291 , \1313 );
buf \U$11949 ( \12292 , \448 );
not \U$11950 ( \12293 , \449 );
and \U$11951 ( \12294 , \12292 , \12293 );
not \U$11952 ( \12295 , \12294 );
buf \U$11953 ( \12296 , \591 );
not \U$11954 ( \12297 , \12296 );
nor \U$11955 ( \12298 , \12295 , \12297 );
not \U$11956 ( \12299 , \12298 );
not \U$11957 ( \12300 , \490 );
buf \U$11958 ( \12301 , \478 );
not \U$11959 ( \12302 , \12301 );
or \U$11960 ( \12303 , \12300 , \12302 );
not \U$11961 ( \12304 , \590 );
nand \U$11962 ( \12305 , \12303 , \12304 );
not \U$11963 ( \12306 , \12305 );
or \U$11964 ( \12307 , \12299 , \12306 );
buf \U$11965 ( \12308 , \443 );
and \U$11966 ( \12309 , \12308 , \12294 );
not \U$11967 ( \12310 , \12293 );
not \U$11968 ( \12311 , \560 );
or \U$11969 ( \12312 , \12310 , \12311 );
nand \U$11970 ( \12313 , \12312 , \565 );
nor \U$11971 ( \12314 , \12309 , \12313 );
nand \U$11972 ( \12315 , \12307 , \12314 );
nor \U$11973 ( \12316 , \563 , \568 );
and \U$11974 ( \12317 , \12315 , \12316 );
not \U$11975 ( \12318 , \12315 );
not \U$11976 ( \12319 , \12316 );
and \U$11977 ( \12320 , \12318 , \12319 );
nor \U$11978 ( \12321 , \12317 , \12320 );
not \U$11979 ( \12322 , \12321 );
buf \U$11980 ( \12323 , \12322 );
not \U$11981 ( \12324 , \12323 );
not \U$11982 ( \12325 , \12324 );
not \U$11983 ( \12326 , \12325 );
or \U$11984 ( \12327 , \12291 , \12326 );
nand \U$11985 ( \12328 , \12324 , \1392 );
nand \U$11986 ( \12329 , \12327 , \12328 );
not \U$11987 ( \12330 , \12329 );
or \U$11988 ( \12331 , \12290 , \12330 );
not \U$11989 ( \12332 , \12305 );
not \U$11990 ( \12333 , \12292 );
nor \U$11991 ( \12334 , \12333 , \12297 );
not \U$11992 ( \12335 , \12334 );
or \U$11993 ( \12336 , \12332 , \12335 );
nand \U$11994 ( \12337 , \12308 , \12292 );
not \U$11995 ( \12338 , \560 );
and \U$11996 ( \12339 , \12337 , \12338 );
nand \U$11997 ( \12340 , \12336 , \12339 );
nand \U$11998 ( \12341 , \12293 , \565 );
not \U$11999 ( \12342 , \12341 );
and \U$12000 ( \12343 , \12340 , \12342 );
not \U$12001 ( \12344 , \12340 );
and \U$12002 ( \12345 , \12344 , \12341 );
nor \U$12003 ( \12346 , \12343 , \12345 );
buf \U$12004 ( \12347 , \12346 );
not \U$12005 ( \12348 , \12347 );
not \U$12006 ( \12349 , \12348 );
xor \U$12007 ( \12350 , \1312 , \12349 );
nand \U$12008 ( \12351 , \12350 , \1429 );
nand \U$12009 ( \12352 , \12331 , \12351 );
not \U$12010 ( \12353 , \8450 );
and \U$12011 ( \12354 , RIbb2e440_39, \3370 );
not \U$12012 ( \12355 , RIbb2e440_39);
and \U$12013 ( \12356 , \12355 , \1687 );
or \U$12014 ( \12357 , \12354 , \12356 );
not \U$12015 ( \12358 , \12357 );
or \U$12016 ( \12359 , \12353 , \12358 );
and \U$12017 ( \12360 , RIbb2e440_39, \3773 );
not \U$12018 ( \12361 , RIbb2e440_39);
and \U$12019 ( \12362 , \12361 , \7033 );
or \U$12020 ( \12363 , \12360 , \12362 );
nand \U$12021 ( \12364 , \12363 , \8445 );
nand \U$12022 ( \12365 , \12359 , \12364 );
xor \U$12023 ( \12366 , \12352 , \12365 );
not \U$12024 ( \12367 , \2963 );
and \U$12025 ( \12368 , RIbb2ead0_25, \3143 );
not \U$12026 ( \12369 , RIbb2ead0_25);
and \U$12027 ( \12370 , \12369 , \3146 );
or \U$12028 ( \12371 , \12368 , \12370 );
not \U$12029 ( \12372 , \12371 );
or \U$12030 ( \12373 , \12367 , \12372 );
and \U$12031 ( \12374 , RIbb2ead0_25, \4639 );
not \U$12032 ( \12375 , RIbb2ead0_25);
and \U$12033 ( \12376 , \12375 , \4640 );
or \U$12034 ( \12377 , \12374 , \12376 );
nand \U$12035 ( \12378 , \12377 , \2980 );
nand \U$12036 ( \12379 , \12373 , \12378 );
and \U$12037 ( \12380 , \12366 , \12379 );
and \U$12038 ( \12381 , \12352 , \12365 );
or \U$12039 ( \12382 , \12380 , \12381 );
and \U$12040 ( \12383 , \12289 , \12382 );
and \U$12041 ( \12384 , \12246 , \12288 );
or \U$12042 ( \12385 , \12383 , \12384 );
and \U$12043 ( \12386 , \12244 , \12385 );
and \U$12044 ( \12387 , \12112 , \12243 );
or \U$12045 ( \12388 , \12386 , \12387 );
not \U$12046 ( \12389 , \11509 );
xor \U$12047 ( \12390 , \12171 , \12176 );
and \U$12048 ( \12391 , \12390 , \12182 );
and \U$12049 ( \12392 , \12171 , \12176 );
or \U$12050 ( \12393 , \12391 , \12392 );
xor \U$12051 ( \12394 , \12389 , \12393 );
not \U$12052 ( \12395 , \998 );
not \U$12053 ( \12396 , \11507 );
or \U$12054 ( \12397 , \12395 , \12396 );
nand \U$12055 ( \12398 , \12118 , \916 );
nand \U$12056 ( \12399 , \12397 , \12398 );
not \U$12057 ( \12400 , \1570 );
not \U$12058 ( \12401 , \11539 );
or \U$12059 ( \12402 , \12400 , \12401 );
nand \U$12060 ( \12403 , \12206 , \1533 );
nand \U$12061 ( \12404 , \12402 , \12403 );
nor \U$12062 ( \12405 , \12399 , \12404 );
and \U$12063 ( \12406 , \1077 , \11556 );
and \U$12064 ( \12407 , \12141 , \1011 );
nor \U$12065 ( \12408 , \12406 , \12407 );
or \U$12066 ( \12409 , \12405 , \12408 );
nand \U$12067 ( \12410 , \12399 , \12404 );
nand \U$12068 ( \12411 , \12409 , \12410 );
xor \U$12069 ( \12412 , \12394 , \12411 );
xor \U$12070 ( \12413 , \12162 , \12183 );
and \U$12071 ( \12414 , \12413 , \12242 );
and \U$12072 ( \12415 , \12162 , \12183 );
or \U$12073 ( \12416 , \12414 , \12415 );
xor \U$12074 ( \12417 , \12412 , \12416 );
xor \U$12075 ( \12418 , \12265 , \12272 );
and \U$12076 ( \12419 , \12418 , \12287 );
and \U$12077 ( \12420 , \12265 , \12272 );
or \U$12078 ( \12421 , \12419 , \12420 );
not \U$12079 ( \12422 , \1265 );
not \U$12080 ( \12423 , \12253 );
or \U$12081 ( \12424 , \12422 , \12423 );
nand \U$12082 ( \12425 , \11714 , \1294 );
nand \U$12083 ( \12426 , \12424 , \12425 );
not \U$12084 ( \12427 , \1090 );
not \U$12085 ( \12428 , \12226 );
or \U$12086 ( \12429 , \12427 , \12428 );
nand \U$12087 ( \12430 , \11704 , \1147 );
nand \U$12088 ( \12431 , \12429 , \12430 );
not \U$12089 ( \12432 , \12431 );
not \U$12090 ( \12433 , \1737 );
not \U$12091 ( \12434 , \11527 );
or \U$12092 ( \12435 , \12433 , \12434 );
nand \U$12093 ( \12436 , \12198 , \1702 );
nand \U$12094 ( \12437 , \12435 , \12436 );
not \U$12095 ( \12438 , \12437 );
and \U$12096 ( \12439 , \12432 , \12438 );
not \U$12097 ( \12440 , \12432 );
and \U$12098 ( \12441 , \12440 , \12437 );
nor \U$12099 ( \12442 , \12439 , \12441 );
xor \U$12100 ( \12443 , \12426 , \12442 );
xor \U$12101 ( \12444 , \12421 , \12443 );
not \U$12102 ( \12445 , \10117 );
not \U$12103 ( \12446 , \12012 );
or \U$12104 ( \12447 , \12445 , \12446 );
not \U$12105 ( \12448 , RIbb2e170_45);
not \U$12106 ( \12449 , \3451 );
or \U$12107 ( \12450 , \12448 , \12449 );
not \U$12108 ( \12451 , RIbb2e170_45);
nand \U$12109 ( \12452 , \1474 , \12451 );
nand \U$12110 ( \12453 , \12450 , \12452 );
nand \U$12111 ( \12454 , \12453 , \10119 );
nand \U$12112 ( \12455 , \12447 , \12454 );
not \U$12113 ( \12456 , \3465 );
not \U$12114 ( \12457 , RIbb2e9e0_27);
not \U$12115 ( \12458 , \3319 );
or \U$12116 ( \12459 , \12457 , \12458 );
nand \U$12117 ( \12460 , \2225 , \3454 );
nand \U$12118 ( \12461 , \12459 , \12460 );
not \U$12119 ( \12462 , \12461 );
or \U$12120 ( \12463 , \12456 , \12462 );
nand \U$12121 ( \12464 , \12101 , \3445 );
nand \U$12122 ( \12465 , \12463 , \12464 );
xor \U$12123 ( \12466 , \12455 , \12465 );
not \U$12124 ( \12467 , \2922 );
not \U$12125 ( \12468 , \12067 );
or \U$12126 ( \12469 , \12467 , \12468 );
not \U$12127 ( \12470 , RIbb2e8f0_29);
not \U$12128 ( \12471 , \1853 );
or \U$12129 ( \12472 , \12470 , \12471 );
nand \U$12130 ( \12473 , \1852 , \3265 );
nand \U$12131 ( \12474 , \12472 , \12473 );
nand \U$12132 ( \12475 , \12474 , \2925 );
nand \U$12133 ( \12476 , \12469 , \12475 );
and \U$12134 ( \12477 , \12466 , \12476 );
and \U$12135 ( \12478 , \12455 , \12465 );
or \U$12136 ( \12479 , \12477 , \12478 );
and \U$12137 ( \12480 , \12444 , \12479 );
and \U$12138 ( \12481 , \12421 , \12443 );
or \U$12139 ( \12482 , \12480 , \12481 );
xor \U$12140 ( \12483 , \12417 , \12482 );
xor \U$12141 ( \12484 , \12388 , \12483 );
not \U$12142 ( \12485 , \1702 );
not \U$12143 ( \12486 , RIbb2f340_7);
not \U$12144 ( \12487 , \10306 );
or \U$12145 ( \12488 , \12486 , \12487 );
nand \U$12146 ( \12489 , \9841 , \1692 );
nand \U$12147 ( \12490 , \12488 , \12489 );
not \U$12148 ( \12491 , \12490 );
or \U$12149 ( \12492 , \12485 , \12491 );
nand \U$12150 ( \12493 , \12190 , \1737 );
nand \U$12151 ( \12494 , \12492 , \12493 );
not \U$12152 ( \12495 , \1533 );
not \U$12153 ( \12496 , RIbb2f250_9);
not \U$12154 ( \12497 , \12194 );
or \U$12155 ( \12498 , \12496 , \12497 );
nand \U$12156 ( \12499 , \8631 , \1566 );
nand \U$12157 ( \12500 , \12498 , \12499 );
not \U$12158 ( \12501 , \12500 );
or \U$12159 ( \12502 , \12495 , \12501 );
nand \U$12160 ( \12503 , \12216 , \1570 );
nand \U$12161 ( \12504 , \12502 , \12503 );
xor \U$12162 ( \12505 , \12494 , \12504 );
not \U$12163 ( \12506 , \1077 );
not \U$12164 ( \12507 , \12134 );
or \U$12165 ( \12508 , \12506 , \12507 );
not \U$12166 ( \12509 , RIbb2f160_11);
not \U$12167 ( \12510 , \9071 );
or \U$12168 ( \12511 , \12509 , \12510 );
nand \U$12169 ( \12512 , \9074 , \1043 );
nand \U$12170 ( \12513 , \12511 , \12512 );
nand \U$12171 ( \12514 , \12513 , \1011 );
nand \U$12172 ( \12515 , \12508 , \12514 );
and \U$12173 ( \12516 , \12505 , \12515 );
and \U$12174 ( \12517 , \12494 , \12504 );
or \U$12175 ( \12518 , \12516 , \12517 );
not \U$12176 ( \12519 , \916 );
not \U$12177 ( \12520 , RIbb2f070_13);
not \U$12178 ( \12521 , \8338 );
or \U$12179 ( \12522 , \12520 , \12521 );
nand \U$12180 ( \12523 , \6604 , \1656 );
nand \U$12181 ( \12524 , \12522 , \12523 );
not \U$12182 ( \12525 , \12524 );
or \U$12183 ( \12526 , \12519 , \12525 );
nand \U$12184 ( \12527 , \12125 , \998 );
nand \U$12185 ( \12528 , \12526 , \12527 );
not \U$12186 ( \12529 , \1445 );
and \U$12187 ( \12530 , RIbb2ef80_15, \10126 );
not \U$12188 ( \12531 , RIbb2ef80_15);
and \U$12189 ( \12532 , \12531 , \6232 );
or \U$12190 ( \12533 , \12530 , \12532 );
not \U$12191 ( \12534 , \12533 );
or \U$12192 ( \12535 , \12529 , \12534 );
nand \U$12193 ( \12536 , \12151 , \1517 );
nand \U$12194 ( \12537 , \12535 , \12536 );
xor \U$12195 ( \12538 , \12528 , \12537 );
not \U$12196 ( \12539 , \836 );
not \U$12197 ( \12540 , RIbb2ee90_17);
not \U$12198 ( \12541 , \4325 );
or \U$12199 ( \12542 , \12540 , \12541 );
nand \U$12200 ( \12543 , \4089 , \3699 );
nand \U$12201 ( \12544 , \12542 , \12543 );
not \U$12202 ( \12545 , \12544 );
or \U$12203 ( \12546 , \12539 , \12545 );
not \U$12204 ( \12547 , RIbb2ee90_17);
not \U$12205 ( \12548 , \12154 );
or \U$12206 ( \12549 , \12547 , \12548 );
nand \U$12207 ( \12550 , \4394 , \816 );
nand \U$12208 ( \12551 , \12549 , \12550 );
nand \U$12209 ( \12552 , \12551 , \832 );
nand \U$12210 ( \12553 , \12546 , \12552 );
and \U$12211 ( \12554 , \12538 , \12553 );
and \U$12212 ( \12555 , \12528 , \12537 );
or \U$12213 ( \12556 , \12554 , \12555 );
xor \U$12214 ( \12557 , \12518 , \12556 );
not \U$12215 ( \12558 , \12167 );
not \U$12216 ( \12559 , RIbb2df90_49);
not \U$12217 ( \12560 , \1579 );
or \U$12218 ( \12561 , \12559 , \12560 );
nand \U$12219 ( \12562 , \892 , \12278 );
nand \U$12220 ( \12563 , \12561 , \12562 );
not \U$12221 ( \12564 , \12563 );
or \U$12222 ( \12565 , \12558 , \12564 );
nand \U$12223 ( \12566 , \12280 , \12285 );
nand \U$12224 ( \12567 , \12565 , \12566 );
not \U$12225 ( \12568 , \855 );
not \U$12226 ( \12569 , RIbb2eda0_19);
not \U$12227 ( \12570 , \4411 );
or \U$12228 ( \12571 , \12569 , \12570 );
nand \U$12229 ( \12572 , \3003 , \5277 );
nand \U$12230 ( \12573 , \12571 , \12572 );
not \U$12231 ( \12574 , \12573 );
or \U$12232 ( \12575 , \12568 , \12574 );
not \U$12233 ( \12576 , RIbb2eda0_19);
not \U$12234 ( \12577 , \10458 );
not \U$12235 ( \12578 , \12577 );
or \U$12236 ( \12579 , \12576 , \12578 );
nand \U$12237 ( \12580 , \10458 , \843 );
nand \U$12238 ( \12581 , \12579 , \12580 );
nand \U$12239 ( \12582 , \12581 , \853 );
nand \U$12240 ( \12583 , \12575 , \12582 );
xor \U$12241 ( \12584 , \12567 , \12583 );
not \U$12242 ( \12585 , \2078 );
not \U$12243 ( \12586 , RIbb2ecb0_21);
not \U$12244 ( \12587 , \5962 );
or \U$12245 ( \12588 , \12586 , \12587 );
nand \U$12246 ( \12589 , \10095 , \849 );
nand \U$12247 ( \12590 , \12588 , \12589 );
not \U$12248 ( \12591 , \12590 );
or \U$12249 ( \12592 , \12585 , \12591 );
not \U$12250 ( \12593 , RIbb2ecb0_21);
not \U$12251 ( \12594 , \8483 );
or \U$12252 ( \12595 , \12593 , \12594 );
not \U$12253 ( \12596 , \8483 );
nand \U$12254 ( \12597 , \12596 , \2254 );
nand \U$12255 ( \12598 , \12595 , \12597 );
nand \U$12256 ( \12599 , \12598 , \2077 );
nand \U$12257 ( \12600 , \12592 , \12599 );
and \U$12258 ( \12601 , \12584 , \12600 );
and \U$12259 ( \12602 , \12567 , \12583 );
or \U$12260 ( \12603 , \12601 , \12602 );
and \U$12261 ( \12604 , \12557 , \12603 );
and \U$12262 ( \12605 , \12518 , \12556 );
or \U$12263 ( \12606 , \12604 , \12605 );
xor \U$12264 ( \12607 , \12421 , \12443 );
xor \U$12265 ( \12608 , \12607 , \12479 );
xor \U$12266 ( \12609 , \12606 , \12608 );
not \U$12267 ( \12610 , \5845 );
and \U$12268 ( \12611 , \8501 , RIbb2e620_35);
not \U$12269 ( \12612 , \8501 );
and \U$12270 ( \12613 , \12612 , \3866 );
or \U$12271 ( \12614 , \12611 , \12613 );
not \U$12272 ( \12615 , \12614 );
or \U$12273 ( \12616 , \12610 , \12615 );
nand \U$12274 ( \12617 , \12040 , \4712 );
nand \U$12275 ( \12618 , \12616 , \12617 );
not \U$12276 ( \12619 , \836 );
not \U$12277 ( \12620 , RIbb2ee90_17);
not \U$12278 ( \12621 , \4040 );
or \U$12279 ( \12622 , \12620 , \12621 );
nand \U$12280 ( \12623 , \6013 , \2240 );
nand \U$12281 ( \12624 , \12622 , \12623 );
not \U$12282 ( \12625 , \12624 );
or \U$12283 ( \12626 , \12619 , \12625 );
nand \U$12284 ( \12627 , \12544 , \832 );
nand \U$12285 ( \12628 , \12626 , \12627 );
xor \U$12286 ( \12629 , \12618 , \12628 );
not \U$12287 ( \12630 , \855 );
not \U$12288 ( \12631 , RIbb2eda0_19);
not \U$12289 ( \12632 , \3045 );
or \U$12290 ( \12633 , \12631 , \12632 );
nand \U$12291 ( \12634 , \3046 , \1776 );
nand \U$12292 ( \12635 , \12633 , \12634 );
not \U$12293 ( \12636 , \12635 );
or \U$12294 ( \12637 , \12630 , \12636 );
nand \U$12295 ( \12638 , \12573 , \853 );
nand \U$12296 ( \12639 , \12637 , \12638 );
and \U$12297 ( \12640 , \12629 , \12639 );
and \U$12298 ( \12641 , \12618 , \12628 );
or \U$12299 ( \12642 , \12640 , \12641 );
not \U$12300 ( \12643 , \8445 );
not \U$12301 ( \12644 , \12357 );
or \U$12302 ( \12645 , \12643 , \12644 );
and \U$12303 ( \12646 , RIbb2e440_39, \3481 );
not \U$12304 ( \12647 , RIbb2e440_39);
and \U$12305 ( \12648 , \12647 , \3480 );
or \U$12306 ( \12649 , \12646 , \12648 );
nand \U$12307 ( \12650 , \12649 , \8450 );
nand \U$12308 ( \12651 , \12645 , \12650 );
not \U$12309 ( \12652 , \6251 );
not \U$12310 ( \12653 , RIbb2e530_37);
not \U$12311 ( \12654 , \3054 );
or \U$12312 ( \12655 , \12653 , \12654 );
nand \U$12313 ( \12656 , \1138 , \8701 );
nand \U$12314 ( \12657 , \12655 , \12656 );
not \U$12315 ( \12658 , \12657 );
or \U$12316 ( \12659 , \12652 , \12658 );
not \U$12317 ( \12660 , RIbb2e530_37);
not \U$12318 ( \12661 , \3239 );
or \U$12319 ( \12662 , \12660 , \12661 );
nand \U$12320 ( \12663 , \7033 , \6246 );
nand \U$12321 ( \12664 , \12662 , \12663 );
nand \U$12322 ( \12665 , \12664 , \6242 );
nand \U$12323 ( \12666 , \12659 , \12665 );
xor \U$12324 ( \12667 , \12651 , \12666 );
not \U$12325 ( \12668 , \2963 );
and \U$12326 ( \12669 , RIbb2ead0_25, \3168 );
not \U$12327 ( \12670 , RIbb2ead0_25);
and \U$12328 ( \12671 , \12670 , \4220 );
or \U$12329 ( \12672 , \12669 , \12671 );
not \U$12330 ( \12673 , \12672 );
or \U$12331 ( \12674 , \12668 , \12673 );
nand \U$12332 ( \12675 , \12371 , \2980 );
nand \U$12333 ( \12676 , \12674 , \12675 );
and \U$12334 ( \12677 , \12667 , \12676 );
and \U$12335 ( \12678 , \12651 , \12666 );
or \U$12336 ( \12679 , \12677 , \12678 );
xor \U$12337 ( \12680 , \12642 , \12679 );
not \U$12338 ( \12681 , RIbb2ddb0_53);
and \U$12339 ( \12682 , \12681 , RIbb2de28_52);
not \U$12340 ( \12683 , RIbb2de28_52);
and \U$12341 ( \12684 , \12683 , RIbb2ddb0_53);
nor \U$12342 ( \12685 , \12682 , \12684 );
and \U$12343 ( \12686 , RIbb2dea0_51, RIbb2de28_52);
not \U$12344 ( \12687 , RIbb2dea0_51);
and \U$12345 ( \12688 , \12687 , \12683 );
nor \U$12346 ( \12689 , \12686 , \12688 );
and \U$12347 ( \12690 , \12685 , \12689 );
not \U$12348 ( \12691 , \12685 );
buf \U$12349 ( \12692 , \12691 );
or \U$12350 ( \12693 , \12690 , \12692 );
nand \U$12351 ( \12694 , \12693 , RIbb2dea0_51);
and \U$12352 ( \12695 , \1312 , \12349 );
xor \U$12353 ( \12696 , \12694 , \12695 );
not \U$12354 ( \12697 , \1376 );
not \U$12355 ( \12698 , \12270 );
or \U$12356 ( \12699 , \12697 , \12698 );
nand \U$12357 ( \12700 , \12329 , \1429 );
nand \U$12358 ( \12701 , \12699 , \12700 );
and \U$12359 ( \12702 , \12696 , \12701 );
and \U$12360 ( \12703 , \12694 , \12695 );
or \U$12361 ( \12704 , \12702 , \12703 );
not \U$12362 ( \12705 , \2078 );
not \U$12363 ( \12706 , RIbb2ecb0_21);
not \U$12364 ( \12707 , \3762 );
not \U$12365 ( \12708 , \12707 );
or \U$12366 ( \12709 , \12706 , \12708 );
nand \U$12367 ( \12710 , \7021 , \849 );
nand \U$12368 ( \12711 , \12709 , \12710 );
not \U$12369 ( \12712 , \12711 );
or \U$12370 ( \12713 , \12705 , \12712 );
nand \U$12371 ( \12714 , \12590 , \2077 );
nand \U$12372 ( \12715 , \12713 , \12714 );
xor \U$12373 ( \12716 , \12704 , \12715 );
not \U$12374 ( \12717 , \3383 );
not \U$12375 ( \12718 , RIbb2ebc0_23);
not \U$12376 ( \12719 , \4639 );
or \U$12377 ( \12720 , \12718 , \12719 );
nand \U$12378 ( \12721 , \7009 , \2073 );
nand \U$12379 ( \12722 , \12720 , \12721 );
not \U$12380 ( \12723 , \12722 );
or \U$12381 ( \12724 , \12717 , \12723 );
not \U$12382 ( \12725 , RIbb2ebc0_23);
not \U$12383 ( \12726 , \3905 );
or \U$12384 ( \12727 , \12725 , \12726 );
nand \U$12385 ( \12728 , \3632 , \2073 );
nand \U$12386 ( \12729 , \12727 , \12728 );
nand \U$12387 ( \12730 , \12729 , \3407 );
nand \U$12388 ( \12731 , \12724 , \12730 );
and \U$12389 ( \12732 , \12716 , \12731 );
and \U$12390 ( \12733 , \12704 , \12715 );
or \U$12391 ( \12734 , \12732 , \12733 );
xor \U$12392 ( \12735 , \12680 , \12734 );
and \U$12393 ( \12736 , \12609 , \12735 );
and \U$12394 ( \12737 , \12606 , \12608 );
or \U$12395 ( \12738 , \12736 , \12737 );
xor \U$12396 ( \12739 , \12484 , \12738 );
not \U$12397 ( \12740 , \1737 );
not \U$12398 ( \12741 , \12490 );
or \U$12399 ( \12742 , \12740 , \12741 );
not \U$12400 ( \12743 , RIbb2f340_7);
not \U$12401 ( \12744 , \10300 );
not \U$12402 ( \12745 , \12744 );
or \U$12403 ( \12746 , \12743 , \12745 );
nand \U$12404 ( \12747 , \10301 , \1734 );
nand \U$12405 ( \12748 , \12746 , \12747 );
nand \U$12406 ( \12749 , \12748 , \1702 );
nand \U$12407 ( \12750 , \12742 , \12749 );
not \U$12408 ( \12751 , \12750 );
not \U$12409 ( \12752 , \1090 );
not \U$12410 ( \12753 , RIbb2f430_5);
not \U$12411 ( \12754 , \11142 );
not \U$12412 ( \12755 , \12754 );
not \U$12413 ( \12756 , \12755 );
not \U$12414 ( \12757 , \12756 );
or \U$12415 ( \12758 , \12753 , \12757 );
nand \U$12416 ( \12759 , \12261 , \1898 );
nand \U$12417 ( \12760 , \12758 , \12759 );
not \U$12418 ( \12761 , \12760 );
or \U$12419 ( \12762 , \12752 , \12761 );
not \U$12420 ( \12763 , RIbb2f430_5);
not \U$12421 ( \12764 , \10764 );
not \U$12422 ( \12765 , \12764 );
or \U$12423 ( \12766 , \12763 , \12765 );
nand \U$12424 ( \12767 , \10764 , \1980 );
nand \U$12425 ( \12768 , \12766 , \12767 );
nand \U$12426 ( \12769 , \12768 , \1147 );
nand \U$12427 ( \12770 , \12762 , \12769 );
not \U$12428 ( \12771 , \12770 );
or \U$12429 ( \12772 , \12751 , \12771 );
or \U$12430 ( \12773 , \12770 , \12750 );
buf \U$12431 ( \12774 , \12690 );
not \U$12432 ( \12775 , \12774 );
and \U$12433 ( \12776 , RIbb2dea0_51, \812 );
not \U$12434 ( \12777 , RIbb2dea0_51);
and \U$12435 ( \12778 , \12777 , \2251 );
or \U$12436 ( \12779 , \12776 , \12778 );
not \U$12437 ( \12780 , \12779 );
or \U$12438 ( \12781 , \12775 , \12780 );
nand \U$12439 ( \12782 , \12692 , RIbb2dea0_51);
nand \U$12440 ( \12783 , \12781 , \12782 );
nand \U$12441 ( \12784 , \12773 , \12783 );
nand \U$12442 ( \12785 , \12772 , \12784 );
not \U$12443 ( \12786 , \916 );
not \U$12444 ( \12787 , RIbb2f070_13);
not \U$12445 ( \12788 , \8639 );
or \U$12446 ( \12789 , \12787 , \12788 );
not \U$12447 ( \12790 , \8637 );
not \U$12448 ( \12791 , \12790 );
nand \U$12449 ( \12792 , \12791 , \906 );
nand \U$12450 ( \12793 , \12789 , \12792 );
not \U$12451 ( \12794 , \12793 );
or \U$12452 ( \12795 , \12786 , \12794 );
nand \U$12453 ( \12796 , \12524 , \998 );
nand \U$12454 ( \12797 , \12795 , \12796 );
not \U$12455 ( \12798 , \12797 );
not \U$12456 ( \12799 , \1011 );
not \U$12457 ( \12800 , RIbb2f160_11);
not \U$12458 ( \12801 , \9818 );
not \U$12459 ( \12802 , \12801 );
or \U$12460 ( \12803 , \12800 , \12802 );
nand \U$12461 ( \12804 , \9819 , \1805 );
nand \U$12462 ( \12805 , \12803 , \12804 );
not \U$12463 ( \12806 , \12805 );
or \U$12464 ( \12807 , \12799 , \12806 );
nand \U$12465 ( \12808 , \12513 , \1077 );
nand \U$12466 ( \12809 , \12807 , \12808 );
not \U$12467 ( \12810 , \12809 );
or \U$12468 ( \12811 , \12798 , \12810 );
or \U$12469 ( \12812 , \12809 , \12797 );
not \U$12470 ( \12813 , \1570 );
not \U$12471 ( \12814 , \12500 );
or \U$12472 ( \12815 , \12813 , \12814 );
not \U$12473 ( \12816 , RIbb2f250_9);
not \U$12474 ( \12817 , \9279 );
or \U$12475 ( \12818 , \12816 , \12817 );
not \U$12476 ( \12819 , \9277 );
buf \U$12477 ( \12820 , \12819 );
not \U$12478 ( \12821 , \12820 );
nand \U$12479 ( \12822 , \12821 , \1566 );
nand \U$12480 ( \12823 , \12818 , \12822 );
nand \U$12481 ( \12824 , \1533 , \12823 );
nand \U$12482 ( \12825 , \12815 , \12824 );
nand \U$12483 ( \12826 , \12812 , \12825 );
nand \U$12484 ( \12827 , \12811 , \12826 );
xor \U$12485 ( \12828 , \12785 , \12827 );
not \U$12486 ( \12829 , \1294 );
not \U$12487 ( \12830 , \1288 );
not \U$12488 ( \12831 , \11580 );
or \U$12489 ( \12832 , \12830 , \12831 );
nand \U$12490 ( \12833 , \11581 , \1244 );
nand \U$12491 ( \12834 , \12832 , \12833 );
not \U$12492 ( \12835 , \12834 );
or \U$12493 ( \12836 , \12829 , \12835 );
not \U$12494 ( \12837 , \1288 );
buf \U$12495 ( \12838 , \12174 );
not \U$12496 ( \12839 , \12838 );
not \U$12497 ( \12840 , \12839 );
or \U$12498 ( \12841 , \12837 , \12840 );
nand \U$12499 ( \12842 , \12838 , \1244 );
nand \U$12500 ( \12843 , \12841 , \12842 );
nand \U$12501 ( \12844 , \12843 , \1264 );
nand \U$12502 ( \12845 , \12836 , \12844 );
not \U$12503 ( \12846 , \6251 );
not \U$12504 ( \12847 , RIbb2e530_37);
not \U$12505 ( \12848 , \3290 );
or \U$12506 ( \12849 , \12847 , \12848 );
nand \U$12507 ( \12850 , \3291 , \8701 );
nand \U$12508 ( \12851 , \12849 , \12850 );
not \U$12509 ( \12852 , \12851 );
or \U$12510 ( \12853 , \12846 , \12852 );
not \U$12511 ( \12854 , RIbb2e530_37);
not \U$12512 ( \12855 , \8501 );
or \U$12513 ( \12856 , \12854 , \12855 );
nand \U$12514 ( \12857 , \4770 , \8701 );
nand \U$12515 ( \12858 , \12856 , \12857 );
nand \U$12516 ( \12859 , \12858 , \6242 );
nand \U$12517 ( \12860 , \12853 , \12859 );
xor \U$12518 ( \12861 , \12845 , \12860 );
not \U$12519 ( \12862 , \2077 );
not \U$12520 ( \12863 , RIbb2ecb0_21);
not \U$12521 ( \12864 , \3276 );
or \U$12522 ( \12865 , \12863 , \12864 );
nand \U$12523 ( \12866 , \3275 , \2254 );
nand \U$12524 ( \12867 , \12865 , \12866 );
not \U$12525 ( \12868 , \12867 );
or \U$12526 ( \12869 , \12862 , \12868 );
nand \U$12527 ( \12870 , \12598 , \2078 );
nand \U$12528 ( \12871 , \12869 , \12870 );
and \U$12529 ( \12872 , \12861 , \12871 );
and \U$12530 ( \12873 , \12845 , \12860 );
or \U$12531 ( \12874 , \12872 , \12873 );
and \U$12532 ( \12875 , \12828 , \12874 );
and \U$12533 ( \12876 , \12785 , \12827 );
or \U$12534 ( \12877 , \12875 , \12876 );
xor \U$12535 ( \12878 , \12494 , \12504 );
xor \U$12536 ( \12879 , \12878 , \12515 );
not \U$12537 ( \12880 , \12879 );
not \U$12538 ( \12881 , \1090 );
not \U$12539 ( \12882 , \12768 );
or \U$12540 ( \12883 , \12881 , \12882 );
nand \U$12541 ( \12884 , \12237 , \1147 );
nand \U$12542 ( \12885 , \12883 , \12884 );
not \U$12543 ( \12886 , \12885 );
not \U$12544 ( \12887 , \1264 );
not \U$12545 ( \12888 , \12834 );
or \U$12546 ( \12889 , \12887 , \12888 );
nand \U$12547 ( \12890 , \1294 , \12263 );
nand \U$12548 ( \12891 , \12889 , \12890 );
not \U$12549 ( \12892 , \12891 );
and \U$12550 ( \12893 , \12886 , \12892 );
not \U$12551 ( \12894 , \12886 );
and \U$12552 ( \12895 , \12894 , \12891 );
or \U$12553 ( \12896 , \12893 , \12895 );
not \U$12554 ( \12897 , \6251 );
not \U$12555 ( \12898 , \12858 );
or \U$12556 ( \12899 , \12897 , \12898 );
nand \U$12557 ( \12900 , \12657 , \6242 );
nand \U$12558 ( \12901 , \12899 , \12900 );
xor \U$12559 ( \12902 , \12896 , \12901 );
not \U$12560 ( \12903 , \12902 );
not \U$12561 ( \12904 , \12903 );
or \U$12562 ( \12905 , \12880 , \12904 );
xor \U$12563 ( \12906 , \12084 , \12103 );
xor \U$12564 ( \12907 , \12906 , \12069 );
not \U$12565 ( \12908 , \12879 );
nand \U$12566 ( \12909 , \12902 , \12908 );
nand \U$12567 ( \12910 , \12907 , \12909 );
nand \U$12568 ( \12911 , \12905 , \12910 );
xor \U$12569 ( \12912 , \12877 , \12911 );
not \U$12570 ( \12913 , \12892 );
not \U$12571 ( \12914 , \12886 );
or \U$12572 ( \12915 , \12913 , \12914 );
nand \U$12573 ( \12916 , \12915 , \12901 );
nand \U$12574 ( \12917 , \12885 , \12891 );
nand \U$12575 ( \12918 , \12916 , \12917 );
xor \U$12576 ( \12919 , \12200 , \12218 );
xor \U$12577 ( \12920 , \12919 , \12239 );
xor \U$12578 ( \12921 , \12918 , \12920 );
xor \U$12579 ( \12922 , \12651 , \12666 );
xor \U$12580 ( \12923 , \12922 , \12676 );
xor \U$12581 ( \12924 , \12921 , \12923 );
and \U$12582 ( \12925 , \12912 , \12924 );
and \U$12583 ( \12926 , \12877 , \12911 );
or \U$12584 ( \12927 , \12925 , \12926 );
xor \U$12585 ( \12928 , \12918 , \12920 );
and \U$12586 ( \12929 , \12928 , \12923 );
and \U$12587 ( \12930 , \12918 , \12920 );
or \U$12588 ( \12931 , \12929 , \12930 );
buf \U$12589 ( \12932 , \12321 );
buf \U$12590 ( \12933 , \12932 );
not \U$12591 ( \12934 , \12933 );
not \U$12592 ( \12935 , \12934 );
nand \U$12593 ( \12936 , \12935 , \1313 );
not \U$12594 ( \12937 , \8362 );
not \U$12595 ( \12938 , \12082 );
or \U$12596 ( \12939 , \12937 , \12938 );
not \U$12597 ( \12940 , RIbb2e350_41);
not \U$12598 ( \12941 , \1562 );
or \U$12599 ( \12942 , \12940 , \12941 );
nand \U$12600 ( \12943 , \1038 , \7097 );
nand \U$12601 ( \12944 , \12942 , \12943 );
nand \U$12602 ( \12945 , \12944 , \8995 );
nand \U$12603 ( \12946 , \12939 , \12945 );
xor \U$12604 ( \12947 , \12936 , \12946 );
not \U$12605 ( \12948 , \2940 );
not \U$12606 ( \12949 , \11977 );
or \U$12607 ( \12950 , \12948 , \12949 );
not \U$12608 ( \12951 , RIbb2e800_31);
not \U$12609 ( \12952 , \3822 );
or \U$12610 ( \12953 , \12951 , \12952 );
nand \U$12611 ( \12954 , \1421 , \9169 );
nand \U$12612 ( \12955 , \12953 , \12954 );
nand \U$12613 ( \12956 , \12955 , \2941 );
nand \U$12614 ( \12957 , \12950 , \12956 );
xor \U$12615 ( \12958 , \12947 , \12957 );
xor \U$12616 ( \12959 , \12455 , \12465 );
xor \U$12617 ( \12960 , \12959 , \12476 );
xor \U$12618 ( \12961 , \12958 , \12960 );
not \U$12619 ( \12962 , \11176 );
not \U$12620 ( \12963 , \11961 );
or \U$12621 ( \12964 , \12962 , \12963 );
buf \U$12622 ( \12965 , \11177 );
not \U$12623 ( \12966 , RIbb2e080_47);
not \U$12624 ( \12967 , \894 );
or \U$12625 ( \12968 , \12966 , \12967 );
not \U$12626 ( \12969 , \892 );
not \U$12627 ( \12970 , \12969 );
not \U$12628 ( \12971 , RIbb2e080_47);
nand \U$12629 ( \12972 , \12970 , \12971 );
nand \U$12630 ( \12973 , \12968 , \12972 );
nand \U$12631 ( \12974 , \12965 , \12973 );
nand \U$12632 ( \12975 , \12964 , \12974 );
not \U$12633 ( \12976 , \4791 );
not \U$12634 ( \12977 , RIbb2e710_33);
not \U$12635 ( \12978 , \11054 );
or \U$12636 ( \12979 , \12977 , \12978 );
nand \U$12637 ( \12980 , \3736 , \3877 );
nand \U$12638 ( \12981 , \12979 , \12980 );
not \U$12639 ( \12982 , \12981 );
or \U$12640 ( \12983 , \12976 , \12982 );
nand \U$12641 ( \12984 , \12028 , \3887 );
nand \U$12642 ( \12985 , \12983 , \12984 );
xor \U$12643 ( \12986 , \12975 , \12985 );
not \U$12644 ( \12987 , \10449 );
not \U$12645 ( \12988 , \11993 );
or \U$12646 ( \12989 , \12987 , \12988 );
not \U$12647 ( \12990 , RIbb2e260_43);
not \U$12648 ( \12991 , \2399 );
or \U$12649 ( \12992 , \12990 , \12991 );
not \U$12650 ( \12993 , \3981 );
nand \U$12651 ( \12994 , \12993 , \8347 );
nand \U$12652 ( \12995 , \12992 , \12994 );
nand \U$12653 ( \12996 , \12995 , \10451 );
nand \U$12654 ( \12997 , \12989 , \12996 );
xor \U$12655 ( \12998 , \12986 , \12997 );
and \U$12656 ( \12999 , \12961 , \12998 );
and \U$12657 ( \13000 , \12958 , \12960 );
or \U$12658 ( \13001 , \12999 , \13000 );
xor \U$12659 ( \13002 , \12931 , \13001 );
xor \U$12660 ( \13003 , \12936 , \12946 );
and \U$12661 ( \13004 , \13003 , \12957 );
and \U$12662 ( \13005 , \12936 , \12946 );
or \U$12663 ( \13006 , \13004 , \13005 );
not \U$12664 ( \13007 , \12404 );
not \U$12665 ( \13008 , \12408 );
or \U$12666 ( \13009 , \13007 , \13008 );
or \U$12667 ( \13010 , \12408 , \12404 );
nand \U$12668 ( \13011 , \13009 , \13010 );
xor \U$12669 ( \13012 , \12399 , \13011 );
xor \U$12670 ( \13013 , \13006 , \13012 );
xor \U$12671 ( \13014 , \12975 , \12985 );
and \U$12672 ( \13015 , \13014 , \12997 );
and \U$12673 ( \13016 , \12975 , \12985 );
or \U$12674 ( \13017 , \13015 , \13016 );
xor \U$12675 ( \13018 , \13013 , \13017 );
xor \U$12676 ( \13019 , \13002 , \13018 );
xor \U$12677 ( \13020 , \12927 , \13019 );
xor \U$12678 ( \13021 , \12606 , \12608 );
xor \U$12679 ( \13022 , \13021 , \12735 );
and \U$12680 ( \13023 , \13020 , \13022 );
and \U$12681 ( \13024 , \12927 , \13019 );
or \U$12682 ( \13025 , \13023 , \13024 );
xor \U$12683 ( \13026 , \12739 , \13025 );
or \U$12684 ( \13027 , \12679 , \12642 );
nand \U$12685 ( \13028 , \13027 , \12734 );
nand \U$12686 ( \13029 , \12679 , \12642 );
nand \U$12687 ( \13030 , \13028 , \13029 );
not \U$12688 ( \13031 , \1376 );
not \U$12689 ( \13032 , \11584 );
or \U$12690 ( \13033 , \13031 , \13032 );
nand \U$12691 ( \13034 , \12267 , \1429 );
nand \U$12692 ( \13035 , \13033 , \13034 );
not \U$12693 ( \13036 , \5845 );
not \U$12694 ( \13037 , \11656 );
or \U$12695 ( \13038 , \13036 , \13037 );
nand \U$12696 ( \13039 , \12614 , \4712 );
nand \U$12697 ( \13040 , \13038 , \13039 );
xor \U$12698 ( \13041 , \13035 , \13040 );
not \U$12699 ( \13042 , \853 );
not \U$12700 ( \13043 , \12635 );
or \U$12701 ( \13044 , \13042 , \13043 );
nand \U$12702 ( \13045 , \11675 , \855 );
nand \U$12703 ( \13046 , \13044 , \13045 );
xor \U$12704 ( \13047 , \13041 , \13046 );
not \U$12705 ( \13048 , \8995 );
not \U$12706 ( \13049 , \11814 );
or \U$12707 ( \13050 , \13048 , \13049 );
nand \U$12708 ( \13051 , \12944 , \8362 );
nand \U$12709 ( \13052 , \13050 , \13051 );
not \U$12710 ( \13053 , \10451 );
not \U$12711 ( \13054 , \11736 );
or \U$12712 ( \13055 , \13053 , \13054 );
nand \U$12713 ( \13056 , \12995 , \10449 );
nand \U$12714 ( \13057 , \13055 , \13056 );
xor \U$12715 ( \13058 , \13052 , \13057 );
not \U$12716 ( \13059 , \3613 );
not \U$12717 ( \13060 , \11834 );
or \U$12718 ( \13061 , \13059 , \13060 );
nand \U$12719 ( \13062 , \12955 , \2940 );
nand \U$12720 ( \13063 , \13061 , \13062 );
xor \U$12721 ( \13064 , \13058 , \13063 );
xor \U$12722 ( \13065 , \13047 , \13064 );
not \U$12723 ( \13066 , \6242 );
not \U$12724 ( \13067 , \11770 );
or \U$12725 ( \13068 , \13066 , \13067 );
nand \U$12726 ( \13069 , \12664 , \6251 );
nand \U$12727 ( \13070 , \13068 , \13069 );
not \U$12728 ( \13071 , \3383 );
not \U$12729 ( \13072 , \11781 );
or \U$12730 ( \13073 , \13071 , \13072 );
nand \U$12731 ( \13074 , \12722 , \3407 );
nand \U$12732 ( \13075 , \13073 , \13074 );
xor \U$12733 ( \13076 , \13070 , \13075 );
not \U$12734 ( \13077 , \2077 );
not \U$12735 ( \13078 , \12711 );
or \U$12736 ( \13079 , \13077 , \13078 );
nand \U$12737 ( \13080 , \11666 , \2078 );
nand \U$12738 ( \13081 , \13079 , \13080 );
xor \U$12739 ( \13082 , \13076 , \13081 );
and \U$12740 ( \13083 , \13065 , \13082 );
and \U$12741 ( \13084 , \13047 , \13064 );
or \U$12742 ( \13085 , \13083 , \13084 );
xor \U$12743 ( \13086 , \13030 , \13085 );
xor \U$12744 ( \13087 , \11696 , \11706 );
xor \U$12745 ( \13088 , \13087 , \11716 );
xor \U$12746 ( \13089 , \13070 , \13075 );
and \U$12747 ( \13090 , \13089 , \13081 );
and \U$12748 ( \13091 , \13070 , \13075 );
or \U$12749 ( \13092 , \13090 , \13091 );
xor \U$12750 ( \13093 , \13088 , \13092 );
xor \U$12751 ( \13094 , \13035 , \13040 );
and \U$12752 ( \13095 , \13094 , \13046 );
and \U$12753 ( \13096 , \13035 , \13040 );
or \U$12754 ( \13097 , \13095 , \13096 );
xor \U$12755 ( \13098 , \13093 , \13097 );
xor \U$12756 ( \13099 , \13086 , \13098 );
not \U$12757 ( \13100 , \13099 );
not \U$12758 ( \13101 , \12936 );
not \U$12759 ( \13102 , \8445 );
not \U$12760 ( \13103 , \12649 );
or \U$12761 ( \13104 , \13102 , \13103 );
nand \U$12762 ( \13105 , \11726 , \8450 );
nand \U$12763 ( \13106 , \13104 , \13105 );
xor \U$12764 ( \13107 , \13101 , \13106 );
not \U$12765 ( \13108 , \2963 );
not \U$12766 ( \13109 , \11760 );
or \U$12767 ( \13110 , \13108 , \13109 );
nand \U$12768 ( \13111 , \12672 , \2980 );
nand \U$12769 ( \13112 , \13110 , \13111 );
xor \U$12770 ( \13113 , \13107 , \13112 );
not \U$12771 ( \13114 , \13113 );
not \U$12772 ( \13115 , \10119 );
not \U$12773 ( \13116 , \11611 );
or \U$12774 ( \13117 , \13115 , \13116 );
nand \U$12775 ( \13118 , \12453 , \10599 );
nand \U$12776 ( \13119 , \13117 , \13118 );
not \U$12777 ( \13120 , \13119 );
not \U$12778 ( \13121 , \3465 );
not \U$12779 ( \13122 , \11745 );
or \U$12780 ( \13123 , \13121 , \13122 );
nand \U$12781 ( \13124 , \12461 , \3445 );
nand \U$12782 ( \13125 , \13123 , \13124 );
not \U$12783 ( \13126 , \13125 );
not \U$12784 ( \13127 , \13126 );
or \U$12785 ( \13128 , \13120 , \13127 );
or \U$12786 ( \13129 , \13126 , \13119 );
nand \U$12787 ( \13130 , \13128 , \13129 );
not \U$12788 ( \13131 , \2925 );
not \U$12789 ( \13132 , \11822 );
or \U$12790 ( \13133 , \13131 , \13132 );
nand \U$12791 ( \13134 , \12474 , \2922 );
nand \U$12792 ( \13135 , \13133 , \13134 );
not \U$12793 ( \13136 , \13135 );
and \U$12794 ( \13137 , \13130 , \13136 );
not \U$12795 ( \13138 , \13130 );
and \U$12796 ( \13139 , \13138 , \13135 );
nor \U$12797 ( \13140 , \13137 , \13139 );
not \U$12798 ( \13141 , \13140 );
or \U$12799 ( \13142 , \13114 , \13141 );
or \U$12800 ( \13143 , \13140 , \13113 );
nand \U$12801 ( \13144 , \13142 , \13143 );
not \U$12802 ( \13145 , \11176 );
not \U$12803 ( \13146 , \12973 );
or \U$12804 ( \13147 , \13145 , \13146 );
nand \U$12805 ( \13148 , \12965 , \11692 );
nand \U$12806 ( \13149 , \13147 , \13148 );
not \U$12807 ( \13150 , \4791 );
not \U$12808 ( \13151 , \11597 );
or \U$12809 ( \13152 , \13150 , \13151 );
nand \U$12810 ( \13153 , \12981 , \3887 );
nand \U$12811 ( \13154 , \13152 , \13153 );
xor \U$12812 ( \13155 , \13149 , \13154 );
not \U$12813 ( \13156 , \836 );
not \U$12814 ( \13157 , \11631 );
or \U$12815 ( \13158 , \13156 , \13157 );
nand \U$12816 ( \13159 , \12624 , \832 );
nand \U$12817 ( \13160 , \13158 , \13159 );
xor \U$12818 ( \13161 , \13155 , \13160 );
not \U$12819 ( \13162 , \13161 );
and \U$12820 ( \13163 , \13144 , \13162 );
not \U$12821 ( \13164 , \13144 );
and \U$12822 ( \13165 , \13164 , \13161 );
nor \U$12823 ( \13166 , \13163 , \13165 );
not \U$12824 ( \13167 , \13166 );
not \U$12825 ( \13168 , \13167 );
xor \U$12826 ( \13169 , \13047 , \13064 );
xor \U$12827 ( \13170 , \13169 , \13082 );
not \U$12828 ( \13171 , \13170 );
or \U$12829 ( \13172 , \13168 , \13171 );
or \U$12830 ( \13173 , \13170 , \13167 );
xor \U$12831 ( \13174 , \12704 , \12715 );
xor \U$12832 ( \13175 , \13174 , \12731 );
xor \U$12833 ( \13176 , \12694 , \12695 );
xor \U$12834 ( \13177 , \13176 , \12701 );
not \U$12835 ( \13178 , \3383 );
not \U$12836 ( \13179 , \12729 );
or \U$12837 ( \13180 , \13178 , \13179 );
not \U$12838 ( \13181 , RIbb2ebc0_23);
not \U$12839 ( \13182 , \3655 );
or \U$12840 ( \13183 , \13181 , \13182 );
nand \U$12841 ( \13184 , \3654 , \3388 );
nand \U$12842 ( \13185 , \13183 , \13184 );
nand \U$12843 ( \13186 , \13185 , \3406 );
nand \U$12844 ( \13187 , \13180 , \13186 );
xor \U$12845 ( \13188 , \13177 , \13187 );
nor \U$12846 ( \13189 , \12297 , \447 );
not \U$12847 ( \13190 , \13189 );
not \U$12848 ( \13191 , \490 );
not \U$12849 ( \13192 , \12301 );
or \U$12850 ( \13193 , \13191 , \13192 );
nand \U$12851 ( \13194 , \13193 , \12304 );
not \U$12852 ( \13195 , \13194 );
or \U$12853 ( \13196 , \13190 , \13195 );
not \U$12854 ( \13197 , \12308 );
not \U$12855 ( \13198 , \447 );
not \U$12856 ( \13199 , \13198 );
or \U$12857 ( \13200 , \13197 , \13199 );
nand \U$12858 ( \13201 , \13200 , \551 );
not \U$12859 ( \13202 , \13201 );
nand \U$12860 ( \13203 , \13196 , \13202 );
and \U$12861 ( \13204 , \556 , \559 );
and \U$12862 ( \13205 , \13203 , \13204 );
not \U$12863 ( \13206 , \13203 );
not \U$12864 ( \13207 , \13204 );
and \U$12865 ( \13208 , \13206 , \13207 );
nor \U$12866 ( \13209 , \13205 , \13208 );
buf \U$12867 ( \13210 , \13209 );
not \U$12868 ( \13211 , \13210 );
not \U$12869 ( \13212 , \13211 );
and \U$12870 ( \13213 , \13212 , \1394 );
not \U$12871 ( \13214 , \836 );
not \U$12872 ( \13215 , \12551 );
or \U$12873 ( \13216 , \13214 , \13215 );
not \U$12874 ( \13217 , RIbb2ee90_17);
not \U$12875 ( \13218 , \4698 );
or \U$12876 ( \13219 , \13217 , \13218 );
nand \U$12877 ( \13220 , \4697 , \822 );
nand \U$12878 ( \13221 , \13219 , \13220 );
nand \U$12879 ( \13222 , \13221 , \832 );
nand \U$12880 ( \13223 , \13216 , \13222 );
xor \U$12881 ( \13224 , \13213 , \13223 );
not \U$12882 ( \13225 , \1517 );
not \U$12883 ( \13226 , \12533 );
or \U$12884 ( \13227 , \13225 , \13226 );
and \U$12885 ( \13228 , RIbb2ef80_15, \5956 );
not \U$12886 ( \13229 , RIbb2ef80_15);
and \U$12887 ( \13230 , \13229 , \5955 );
or \U$12888 ( \13231 , \13228 , \13230 );
nand \U$12889 ( \13232 , \13231 , \1445 );
nand \U$12890 ( \13233 , \13227 , \13232 );
and \U$12891 ( \13234 , \13224 , \13233 );
and \U$12892 ( \13235 , \13213 , \13223 );
or \U$12893 ( \13236 , \13234 , \13235 );
and \U$12894 ( \13237 , \13188 , \13236 );
and \U$12895 ( \13238 , \13177 , \13187 );
or \U$12896 ( \13239 , \13237 , \13238 );
xor \U$12897 ( \13240 , \13175 , \13239 );
xor \U$12898 ( \13241 , \12618 , \12628 );
xor \U$12899 ( \13242 , \13241 , \12639 );
and \U$12900 ( \13243 , \13240 , \13242 );
and \U$12901 ( \13244 , \13175 , \13239 );
or \U$12902 ( \13245 , \13243 , \13244 );
nand \U$12903 ( \13246 , \13173 , \13245 );
nand \U$12904 ( \13247 , \13172 , \13246 );
xor \U$12905 ( \13248 , \12931 , \13001 );
and \U$12906 ( \13249 , \13248 , \13018 );
and \U$12907 ( \13250 , \12931 , \13001 );
or \U$12908 ( \13251 , \13249 , \13250 );
xnor \U$12909 ( \13252 , \13247 , \13251 );
not \U$12910 ( \13253 , \13252 );
or \U$12911 ( \13254 , \13100 , \13253 );
or \U$12912 ( \13255 , \13252 , \13099 );
nand \U$12913 ( \13256 , \13254 , \13255 );
xor \U$12914 ( \13257 , \13026 , \13256 );
xor \U$12915 ( \13258 , \12958 , \12960 );
xor \U$12916 ( \13259 , \13258 , \12998 );
xor \U$12917 ( \13260 , \13175 , \13239 );
xor \U$12918 ( \13261 , \13260 , \13242 );
xor \U$12919 ( \13262 , \13259 , \13261 );
xor \U$12920 ( \13263 , \13177 , \13187 );
xor \U$12921 ( \13264 , \13263 , \13236 );
xor \U$12922 ( \13265 , \12750 , \12770 );
xor \U$12923 ( \13266 , \13265 , \12783 );
xor \U$12924 ( \13267 , \13213 , \13223 );
xor \U$12925 ( \13268 , \13267 , \13233 );
xor \U$12926 ( \13269 , \13266 , \13268 );
xor \U$12927 ( \13270 , \12825 , \12797 );
xor \U$12928 ( \13271 , \13270 , \12809 );
and \U$12929 ( \13272 , \13269 , \13271 );
and \U$12930 ( \13273 , \13266 , \13268 );
or \U$12931 ( \13274 , \13272 , \13273 );
xor \U$12932 ( \13275 , \13264 , \13274 );
not \U$12933 ( \13276 , \2941 );
not \U$12934 ( \13277 , RIbb2e800_31);
not \U$12935 ( \13278 , \4449 );
or \U$12936 ( \13279 , \13277 , \13278 );
not \U$12937 ( \13280 , \2115 );
nand \U$12938 ( \13281 , \13280 , \9169 );
nand \U$12939 ( \13282 , \13279 , \13281 );
not \U$12940 ( \13283 , \13282 );
or \U$12941 ( \13284 , \13276 , \13283 );
not \U$12942 ( \13285 , RIbb2e800_31);
not \U$12943 ( \13286 , \2222 );
not \U$12944 ( \13287 , \13286 );
or \U$12945 ( \13288 , \13285 , \13287 );
not \U$12946 ( \13289 , \2222 );
not \U$12947 ( \13290 , \13289 );
nand \U$12948 ( \13291 , \13290 , \4096 );
nand \U$12949 ( \13292 , \13288 , \13291 );
nand \U$12950 ( \13293 , \13292 , \2940 );
nand \U$12951 ( \13294 , \13284 , \13293 );
buf \U$12952 ( \13295 , \12167 );
not \U$12953 ( \13296 , \13295 );
not \U$12954 ( \13297 , RIbb2df90_49);
not \U$12955 ( \13298 , \3451 );
or \U$12956 ( \13299 , \13297 , \13298 );
nand \U$12957 ( \13300 , \3450 , \12278 );
nand \U$12958 ( \13301 , \13299 , \13300 );
not \U$12959 ( \13302 , \13301 );
or \U$12960 ( \13303 , \13296 , \13302 );
not \U$12961 ( \13304 , RIbb2df90_49);
not \U$12962 ( \13305 , \8754 );
or \U$12963 ( \13306 , \13304 , \13305 );
not \U$12964 ( \13307 , \1508 );
not \U$12965 ( \13308 , \13307 );
nand \U$12966 ( \13309 , \13308 , \12278 );
nand \U$12967 ( \13310 , \13306 , \13309 );
nand \U$12968 ( \13311 , \13310 , \12285 );
nand \U$12969 ( \13312 , \13303 , \13311 );
xor \U$12970 ( \13313 , \13294 , \13312 );
not \U$12971 ( \13314 , \9099 );
not \U$12972 ( \13315 , RIbb2e260_43);
not \U$12973 ( \13316 , \5003 );
or \U$12974 ( \13317 , \13315 , \13316 );
nand \U$12975 ( \13318 , \1548 , \8347 );
nand \U$12976 ( \13319 , \13317 , \13318 );
not \U$12977 ( \13320 , \13319 );
or \U$12978 ( \13321 , \13314 , \13320 );
not \U$12979 ( \13322 , RIbb2e260_43);
not \U$12980 ( \13323 , \3479 );
or \U$12981 ( \13324 , \13322 , \13323 );
nand \U$12982 ( \13325 , \1730 , \8347 );
nand \U$12983 ( \13326 , \13324 , \13325 );
nand \U$12984 ( \13327 , \13326 , \9098 );
nand \U$12985 ( \13328 , \13321 , \13327 );
and \U$12986 ( \13329 , \13313 , \13328 );
and \U$12987 ( \13330 , \13294 , \13312 );
or \U$12988 ( \13331 , \13329 , \13330 );
not \U$12989 ( \13332 , \4712 );
not \U$12990 ( \13333 , RIbb2e620_35);
not \U$12991 ( \13334 , \3822 );
or \U$12992 ( \13335 , \13333 , \13334 );
nand \U$12993 ( \13336 , \1421 , \6002 );
nand \U$12994 ( \13337 , \13335 , \13336 );
not \U$12995 ( \13338 , \13337 );
or \U$12996 ( \13339 , \13332 , \13338 );
not \U$12997 ( \13340 , RIbb2e620_35);
not \U$12998 ( \13341 , \4339 );
or \U$12999 ( \13342 , \13340 , \13341 );
nand \U$13000 ( \13343 , \1386 , \3866 );
nand \U$13001 ( \13344 , \13342 , \13343 );
nand \U$13002 ( \13345 , \13344 , \5845 );
nand \U$13003 ( \13346 , \13339 , \13345 );
not \U$13004 ( \13347 , \13346 );
not \U$13005 ( \13348 , \3887 );
not \U$13006 ( \13349 , RIbb2e710_33);
not \U$13007 ( \13350 , \1853 );
or \U$13008 ( \13351 , \13349 , \13350 );
not \U$13009 ( \13352 , RIbb2e710_33);
nand \U$13010 ( \13353 , \4610 , \13352 );
nand \U$13011 ( \13354 , \13351 , \13353 );
not \U$13012 ( \13355 , \13354 );
or \U$13013 ( \13356 , \13348 , \13355 );
not \U$13014 ( \13357 , RIbb2e710_33);
not \U$13015 ( \13358 , \1338 );
not \U$13016 ( \13359 , \13358 );
or \U$13017 ( \13360 , \13357 , \13359 );
nand \U$13018 ( \13361 , \6096 , \3877 );
nand \U$13019 ( \13362 , \13360 , \13361 );
nand \U$13020 ( \13363 , \13362 , \4791 );
nand \U$13021 ( \13364 , \13356 , \13363 );
not \U$13022 ( \13365 , \13364 );
or \U$13023 ( \13366 , \13347 , \13365 );
or \U$13024 ( \13367 , \13364 , \13346 );
not \U$13025 ( \13368 , \10599 );
not \U$13026 ( \13369 , RIbb2e170_45);
not \U$13027 ( \13370 , \4595 );
or \U$13028 ( \13371 , \13369 , \13370 );
not \U$13029 ( \13372 , RIbb2e170_45);
nand \U$13030 ( \13373 , \1561 , \13372 );
nand \U$13031 ( \13374 , \13371 , \13373 );
not \U$13032 ( \13375 , \13374 );
or \U$13033 ( \13376 , \13368 , \13375 );
not \U$13034 ( \13377 , \13372 );
not \U$13035 ( \13378 , \3099 );
or \U$13036 ( \13379 , \13377 , \13378 );
not \U$13037 ( \13380 , \1886 );
nand \U$13038 ( \13381 , \13380 , RIbb2e170_45);
nand \U$13039 ( \13382 , \13379 , \13381 );
nand \U$13040 ( \13383 , \13382 , \10119 );
nand \U$13041 ( \13384 , \13376 , \13383 );
nand \U$13042 ( \13385 , \13367 , \13384 );
nand \U$13043 ( \13386 , \13366 , \13385 );
xor \U$13044 ( \13387 , \13331 , \13386 );
not \U$13045 ( \13388 , \8995 );
not \U$13046 ( \13389 , RIbb2e350_41);
not \U$13047 ( \13390 , \3368 );
or \U$13048 ( \13391 , \13389 , \13390 );
not \U$13049 ( \13392 , RIbb2e350_41);
nand \U$13050 ( \13393 , \1687 , \13392 );
nand \U$13051 ( \13394 , \13391 , \13393 );
not \U$13052 ( \13395 , \13394 );
or \U$13053 ( \13396 , \13388 , \13395 );
not \U$13054 ( \13397 , RIbb2e350_41);
not \U$13055 ( \13398 , \3238 );
or \U$13056 ( \13399 , \13397 , \13398 );
not \U$13057 ( \13400 , RIbb2e350_41);
nand \U$13058 ( \13401 , \3243 , \13400 );
nand \U$13059 ( \13402 , \13399 , \13401 );
nand \U$13060 ( \13403 , \13402 , \8362 );
nand \U$13061 ( \13404 , \13396 , \13403 );
not \U$13062 ( \13405 , \2925 );
not \U$13063 ( \13406 , RIbb2e8f0_29);
not \U$13064 ( \13407 , \3517 );
or \U$13065 ( \13408 , \13406 , \13407 );
nand \U$13066 ( \13409 , \12096 , \6970 );
nand \U$13067 ( \13410 , \13408 , \13409 );
not \U$13068 ( \13411 , \13410 );
or \U$13069 ( \13412 , \13405 , \13411 );
not \U$13070 ( \13413 , RIbb2e8f0_29);
not \U$13071 ( \13414 , \3166 );
not \U$13072 ( \13415 , \13414 );
or \U$13073 ( \13416 , \13413 , \13415 );
nand \U$13074 ( \13417 , \3951 , \3440 );
nand \U$13075 ( \13418 , \13416 , \13417 );
nand \U$13076 ( \13419 , \13418 , \2922 );
nand \U$13077 ( \13420 , \13412 , \13419 );
xor \U$13078 ( \13421 , \13404 , \13420 );
not \U$13079 ( \13422 , \3465 );
not \U$13080 ( \13423 , RIbb2e9e0_27);
not \U$13081 ( \13424 , \3143 );
or \U$13082 ( \13425 , \13423 , \13424 );
nand \U$13083 ( \13426 , \3146 , \6065 );
nand \U$13084 ( \13427 , \13425 , \13426 );
not \U$13085 ( \13428 , \13427 );
or \U$13086 ( \13429 , \13422 , \13428 );
not \U$13087 ( \13430 , RIbb2e9e0_27);
not \U$13088 ( \13431 , \4639 );
or \U$13089 ( \13432 , \13430 , \13431 );
nand \U$13090 ( \13433 , \3202 , \3454 );
nand \U$13091 ( \13434 , \13432 , \13433 );
nand \U$13092 ( \13435 , \13434 , \3445 );
nand \U$13093 ( \13436 , \13429 , \13435 );
and \U$13094 ( \13437 , \13421 , \13436 );
and \U$13095 ( \13438 , \13404 , \13420 );
or \U$13096 ( \13439 , \13437 , \13438 );
and \U$13097 ( \13440 , \13387 , \13439 );
and \U$13098 ( \13441 , \13331 , \13386 );
or \U$13099 ( \13442 , \13440 , \13441 );
and \U$13100 ( \13443 , \13275 , \13442 );
and \U$13101 ( \13444 , \13264 , \13274 );
or \U$13102 ( \13445 , \13443 , \13444 );
xnor \U$13103 ( \13446 , \13262 , \13445 );
not \U$13104 ( \13447 , \13446 );
not \U$13105 ( \13448 , \13447 );
xor \U$13106 ( \13449 , \12014 , \12030 );
xor \U$13107 ( \13450 , \13449 , \12050 );
xor \U$13108 ( \13451 , \12567 , \12583 );
xor \U$13109 ( \13452 , \13451 , \12600 );
xor \U$13110 ( \13453 , \13450 , \13452 );
xor \U$13111 ( \13454 , \11963 , \11995 );
xor \U$13112 ( \13455 , \13454 , \11979 );
xor \U$13113 ( \13456 , \13453 , \13455 );
xor \U$13114 ( \13457 , \12352 , \12365 );
xor \U$13115 ( \13458 , \13457 , \12379 );
xor \U$13116 ( \13459 , RIbb2dd38_54, RIbb2dcc0_55);
not \U$13117 ( \13460 , \13459 );
and \U$13118 ( \13461 , RIbb2dd38_54, RIbb2ddb0_53);
not \U$13119 ( \13462 , RIbb2dd38_54);
not \U$13120 ( \13463 , RIbb2ddb0_53);
and \U$13121 ( \13464 , \13462 , \13463 );
nor \U$13122 ( \13465 , \13461 , \13464 );
nand \U$13123 ( \13466 , \13460 , \13465 );
not \U$13124 ( \13467 , \13466 );
or \U$13125 ( \13468 , \13467 , \13459 );
nand \U$13126 ( \13469 , \13468 , RIbb2ddb0_53);
not \U$13127 ( \13470 , \1376 );
not \U$13128 ( \13471 , \12350 );
or \U$13129 ( \13472 , \13470 , \13471 );
not \U$13130 ( \13473 , \1393 );
buf \U$13131 ( \13474 , \13210 );
not \U$13132 ( \13475 , \13474 );
not \U$13133 ( \13476 , \13475 );
or \U$13134 ( \13477 , \13473 , \13476 );
nand \U$13135 ( \13478 , \13212 , \1392 );
nand \U$13136 ( \13479 , \13477 , \13478 );
nand \U$13137 ( \13480 , \13479 , \1429 );
nand \U$13138 ( \13481 , \13472 , \13480 );
xor \U$13139 ( \13482 , \13469 , \13481 );
not \U$13140 ( \13483 , \1294 );
not \U$13141 ( \13484 , \12843 );
or \U$13142 ( \13485 , \13483 , \13484 );
and \U$13143 ( \13486 , \1288 , \12934 );
not \U$13144 ( \13487 , \1288 );
and \U$13145 ( \13488 , \13487 , \12933 );
or \U$13146 ( \13489 , \13486 , \13488 );
nand \U$13147 ( \13490 , \13489 , \1264 );
nand \U$13148 ( \13491 , \13485 , \13490 );
and \U$13149 ( \13492 , \13482 , \13491 );
and \U$13150 ( \13493 , \13469 , \13481 );
or \U$13151 ( \13494 , \13492 , \13493 );
not \U$13152 ( \13495 , \1570 );
not \U$13153 ( \13496 , \12823 );
or \U$13154 ( \13497 , \13495 , \13496 );
not \U$13155 ( \13498 , \9840 );
and \U$13156 ( \13499 , \13498 , RIbb2f250_9);
not \U$13157 ( \13500 , \13498 );
and \U$13158 ( \13501 , \13500 , \1554 );
or \U$13159 ( \13502 , \13499 , \13501 );
nand \U$13160 ( \13503 , \13502 , \1533 );
nand \U$13161 ( \13504 , \13497 , \13503 );
not \U$13162 ( \13505 , \13504 );
not \U$13163 ( \13506 , \1147 );
not \U$13164 ( \13507 , \12760 );
or \U$13165 ( \13508 , \13506 , \13507 );
not \U$13166 ( \13509 , RIbb2f430_5);
not \U$13167 ( \13510 , \11579 );
or \U$13168 ( \13511 , \13509 , \13510 );
nand \U$13169 ( \13512 , \11578 , \1085 );
nand \U$13170 ( \13513 , \13511 , \13512 );
nand \U$13171 ( \13514 , \13513 , \1090 );
nand \U$13172 ( \13515 , \13508 , \13514 );
not \U$13173 ( \13516 , \13515 );
or \U$13174 ( \13517 , \13505 , \13516 );
or \U$13175 ( \13518 , \13515 , \13504 );
not \U$13176 ( \13519 , \1737 );
not \U$13177 ( \13520 , \12748 );
or \U$13178 ( \13521 , \13519 , \13520 );
not \U$13179 ( \13522 , RIbb2f340_7);
not \U$13180 ( \13523 , \12249 );
or \U$13181 ( \13524 , \13522 , \13523 );
buf \U$13182 ( \13525 , \10763 );
buf \U$13183 ( \13526 , \13525 );
nand \U$13184 ( \13527 , \13526 , \2700 );
nand \U$13185 ( \13528 , \13524 , \13527 );
nand \U$13186 ( \13529 , \13528 , \1702 );
nand \U$13187 ( \13530 , \13521 , \13529 );
nand \U$13188 ( \13531 , \13518 , \13530 );
nand \U$13189 ( \13532 , \13517 , \13531 );
xor \U$13190 ( \13533 , \13494 , \13532 );
not \U$13191 ( \13534 , \12296 );
not \U$13192 ( \13535 , \12305 );
or \U$13193 ( \13536 , \13534 , \13535 );
not \U$13194 ( \13537 , \12308 );
nand \U$13195 ( \13538 , \13536 , \13537 );
nand \U$13196 ( \13539 , \13198 , \551 );
not \U$13197 ( \13540 , \13539 );
and \U$13198 ( \13541 , \13538 , \13540 );
not \U$13199 ( \13542 , \13538 );
and \U$13200 ( \13543 , \13542 , \13539 );
nor \U$13201 ( \13544 , \13541 , \13543 );
buf \U$13202 ( \13545 , \13544 );
not \U$13203 ( \13546 , \13545 );
not \U$13204 ( \13547 , \13546 );
and \U$13205 ( \13548 , \13547 , \1394 );
not \U$13206 ( \13549 , \855 );
not \U$13207 ( \13550 , RIbb2eda0_19);
buf \U$13208 ( \13551 , \4085 );
not \U$13209 ( \13552 , \13551 );
not \U$13210 ( \13553 , \13552 );
or \U$13211 ( \13554 , \13550 , \13553 );
nand \U$13212 ( \13555 , \4086 , \843 );
nand \U$13213 ( \13556 , \13554 , \13555 );
not \U$13214 ( \13557 , \13556 );
or \U$13215 ( \13558 , \13549 , \13557 );
not \U$13216 ( \13559 , \4390 );
buf \U$13217 ( \13560 , \13559 );
and \U$13218 ( \13561 , \13560 , RIbb2eda0_19);
not \U$13219 ( \13562 , \13560 );
and \U$13220 ( \13563 , \13562 , \1776 );
or \U$13221 ( \13564 , \13561 , \13563 );
nand \U$13222 ( \13565 , \13564 , \853 );
nand \U$13223 ( \13566 , \13558 , \13565 );
xor \U$13224 ( \13567 , \13548 , \13566 );
not \U$13225 ( \13568 , \832 );
not \U$13226 ( \13569 , RIbb2ee90_17);
not \U$13227 ( \13570 , \10126 );
or \U$13228 ( \13571 , \13569 , \13570 );
nand \U$13229 ( \13572 , \7111 , \3057 );
nand \U$13230 ( \13573 , \13571 , \13572 );
not \U$13231 ( \13574 , \13573 );
or \U$13232 ( \13575 , \13568 , \13574 );
nand \U$13233 ( \13576 , \13221 , \836 );
nand \U$13234 ( \13577 , \13575 , \13576 );
and \U$13235 ( \13578 , \13567 , \13577 );
and \U$13236 ( \13579 , \13548 , \13566 );
or \U$13237 ( \13580 , \13578 , \13579 );
and \U$13238 ( \13581 , \13533 , \13580 );
and \U$13239 ( \13582 , \13494 , \13532 );
or \U$13240 ( \13583 , \13581 , \13582 );
xor \U$13241 ( \13584 , \13458 , \13583 );
xor \U$13242 ( \13585 , \12785 , \12827 );
xor \U$13243 ( \13586 , \13585 , \12874 );
xor \U$13244 ( \13587 , \13584 , \13586 );
xor \U$13245 ( \13588 , \13456 , \13587 );
not \U$13246 ( \13589 , \5845 );
not \U$13247 ( \13590 , \13337 );
or \U$13248 ( \13591 , \13589 , \13590 );
not \U$13249 ( \13592 , RIbb2e620_35);
not \U$13250 ( \13593 , \3494 );
or \U$13251 ( \13594 , \13592 , \13593 );
nand \U$13252 ( \13595 , \1337 , \6688 );
nand \U$13253 ( \13596 , \13594 , \13595 );
nand \U$13254 ( \13597 , \13596 , \4712 );
nand \U$13255 ( \13598 , \13591 , \13597 );
not \U$13256 ( \13599 , \12965 );
not \U$13257 ( \13600 , RIbb2e080_47);
not \U$13258 ( \13601 , \10421 );
or \U$13259 ( \13602 , \13600 , \13601 );
nand \U$13260 ( \13603 , \952 , \10113 );
nand \U$13261 ( \13604 , \13602 , \13603 );
not \U$13262 ( \13605 , \13604 );
or \U$13263 ( \13606 , \13599 , \13605 );
not \U$13264 ( \13607 , RIbb2e080_47);
not \U$13265 ( \13608 , \1069 );
or \U$13266 ( \13609 , \13607 , \13608 );
not \U$13267 ( \13610 , \1068 );
not \U$13268 ( \13611 , \13610 );
nand \U$13269 ( \13612 , \13611 , \10113 );
nand \U$13270 ( \13613 , \13609 , \13612 );
nand \U$13271 ( \13614 , \13613 , \11176 );
nand \U$13272 ( \13615 , \13606 , \13614 );
or \U$13273 ( \13616 , \13598 , \13615 );
not \U$13274 ( \13617 , \6251 );
not \U$13275 ( \13618 , RIbb2e530_37);
not \U$13276 ( \13619 , \1384 );
not \U$13277 ( \13620 , \13619 );
or \U$13278 ( \13621 , \13618 , \13620 );
nand \U$13279 ( \13622 , \1386 , \6246 );
nand \U$13280 ( \13623 , \13621 , \13622 );
not \U$13281 ( \13624 , \13623 );
or \U$13282 ( \13625 , \13617 , \13624 );
not \U$13283 ( \13626 , RIbb2e530_37);
not \U$13284 ( \13627 , \3990 );
or \U$13285 ( \13628 , \13626 , \13627 );
nand \U$13286 ( \13629 , \12046 , \7243 );
nand \U$13287 ( \13630 , \13628 , \13629 );
nand \U$13288 ( \13631 , \13630 , \6242 );
nand \U$13289 ( \13632 , \13625 , \13631 );
nand \U$13290 ( \13633 , \13616 , \13632 );
nand \U$13291 ( \13634 , \13598 , \13615 );
nand \U$13292 ( \13635 , \13633 , \13634 );
xor \U$13293 ( \13636 , \13504 , \13530 );
xor \U$13294 ( \13637 , \13636 , \13515 );
xor \U$13295 ( \13638 , \13635 , \13637 );
not \U$13296 ( \13639 , \4791 );
not \U$13297 ( \13640 , \13354 );
or \U$13298 ( \13641 , \13639 , \13640 );
not \U$13299 ( \13642 , RIbb2e710_33);
not \U$13300 ( \13643 , \9983 );
or \U$13301 ( \13644 , \13642 , \13643 );
nand \U$13302 ( \13645 , \3309 , \6844 );
nand \U$13303 ( \13646 , \13644 , \13645 );
nand \U$13304 ( \13647 , \13646 , \3887 );
nand \U$13305 ( \13648 , \13641 , \13647 );
not \U$13306 ( \13649 , \10119 );
not \U$13307 ( \13650 , \13374 );
or \U$13308 ( \13651 , \13649 , \13650 );
not \U$13309 ( \13652 , RIbb2e170_45);
not \U$13310 ( \13653 , \5003 );
or \U$13311 ( \13654 , \13652 , \13653 );
not \U$13312 ( \13655 , RIbb2e170_45);
nand \U$13313 ( \13656 , \13655 , \1547 );
nand \U$13314 ( \13657 , \13654 , \13656 );
nand \U$13315 ( \13658 , \13657 , \10599 );
nand \U$13316 ( \13659 , \13651 , \13658 );
xor \U$13317 ( \13660 , \13648 , \13659 );
not \U$13318 ( \13661 , \12285 );
not \U$13319 ( \13662 , \13301 );
or \U$13320 ( \13663 , \13661 , \13662 );
not \U$13321 ( \13664 , RIbb2df90_49);
not \U$13322 ( \13665 , \985 );
or \U$13323 ( \13666 , \13664 , \13665 );
nand \U$13324 ( \13667 , \984 , \12278 );
nand \U$13325 ( \13668 , \13666 , \13667 );
nand \U$13326 ( \13669 , \13668 , \12167 );
nand \U$13327 ( \13670 , \13663 , \13669 );
and \U$13328 ( \13671 , \13660 , \13670 );
and \U$13329 ( \13672 , \13648 , \13659 );
or \U$13330 ( \13673 , \13671 , \13672 );
and \U$13331 ( \13674 , \13638 , \13673 );
and \U$13332 ( \13675 , \13635 , \13637 );
or \U$13333 ( \13676 , \13674 , \13675 );
not \U$13334 ( \13677 , \1147 );
not \U$13335 ( \13678 , \13513 );
or \U$13336 ( \13679 , \13677 , \13678 );
not \U$13337 ( \13680 , \12174 );
and \U$13338 ( \13681 , RIbb2f430_5, \13680 );
not \U$13339 ( \13682 , RIbb2f430_5);
and \U$13340 ( \13683 , \13682 , \12175 );
or \U$13341 ( \13684 , \13681 , \13683 );
nand \U$13342 ( \13685 , \13684 , \1089 );
nand \U$13343 ( \13686 , \13679 , \13685 );
not \U$13344 ( \13687 , \1737 );
not \U$13345 ( \13688 , \13528 );
or \U$13346 ( \13689 , \13687 , \13688 );
and \U$13347 ( \13690 , RIbb2f340_7, \12257 );
not \U$13348 ( \13691 , RIbb2f340_7);
not \U$13349 ( \13692 , \12257 );
and \U$13350 ( \13693 , \13691 , \13692 );
or \U$13351 ( \13694 , \13690 , \13693 );
nand \U$13352 ( \13695 , \13694 , \1702 );
nand \U$13353 ( \13696 , \13689 , \13695 );
xor \U$13354 ( \13697 , \13686 , \13696 );
not \U$13355 ( \13698 , \8445 );
and \U$13356 ( \13699 , RIbb2e440_39, \1281 );
not \U$13357 ( \13700 , RIbb2e440_39);
and \U$13358 ( \13701 , \13700 , \1282 );
or \U$13359 ( \13702 , \13699 , \13701 );
not \U$13360 ( \13703 , \13702 );
or \U$13361 ( \13704 , \13698 , \13703 );
and \U$13362 ( \13705 , RIbb2e440_39, \1112 );
not \U$13363 ( \13706 , RIbb2e440_39);
not \U$13364 ( \13707 , \4765 );
not \U$13365 ( \13708 , \13707 );
and \U$13366 ( \13709 , \13706 , \13708 );
or \U$13367 ( \13710 , \13705 , \13709 );
nand \U$13368 ( \13711 , \13710 , \7104 );
nand \U$13369 ( \13712 , \13704 , \13711 );
and \U$13370 ( \13713 , \13697 , \13712 );
and \U$13371 ( \13714 , \13686 , \13696 );
or \U$13372 ( \13715 , \13713 , \13714 );
not \U$13373 ( \13716 , \12692 );
xor \U$13374 ( \13717 , RIbb2dea0_51, \892 );
not \U$13375 ( \13718 , \13717 );
or \U$13376 ( \13719 , \13716 , \13718 );
and \U$13377 ( \13720 , RIbb2dea0_51, \8754 );
not \U$13378 ( \13721 , RIbb2dea0_51);
and \U$13379 ( \13722 , \13721 , \1508 );
or \U$13380 ( \13723 , \13720 , \13722 );
nand \U$13381 ( \13724 , \13723 , \12774 );
nand \U$13382 ( \13725 , \13719 , \13724 );
not \U$13383 ( \13726 , \3406 );
not \U$13384 ( \13727 , RIbb2ebc0_23);
not \U$13385 ( \13728 , \3002 );
not \U$13386 ( \13729 , \13728 );
or \U$13387 ( \13730 , \13727 , \13729 );
not \U$13388 ( \13731 , \3000 );
not \U$13389 ( \13732 , \13731 );
nand \U$13390 ( \13733 , \13732 , \2073 );
nand \U$13391 ( \13734 , \13730 , \13733 );
not \U$13392 ( \13735 , \13734 );
or \U$13393 ( \13736 , \13726 , \13735 );
not \U$13394 ( \13737 , RIbb2ebc0_23);
not \U$13395 ( \13738 , \3044 );
not \U$13396 ( \13739 , \13738 );
or \U$13397 ( \13740 , \13737 , \13739 );
nand \U$13398 ( \13741 , \12596 , \2073 );
nand \U$13399 ( \13742 , \13740 , \13741 );
nand \U$13400 ( \13743 , \13742 , \3383 );
nand \U$13401 ( \13744 , \13736 , \13743 );
xor \U$13402 ( \13745 , \13725 , \13744 );
not \U$13403 ( \13746 , \2078 );
not \U$13404 ( \13747 , RIbb2ecb0_21);
not \U$13405 ( \13748 , \4752 );
or \U$13406 ( \13749 , \13747 , \13748 );
not \U$13407 ( \13750 , \4748 );
nand \U$13408 ( \13751 , \13750 , \849 );
nand \U$13409 ( \13752 , \13749 , \13751 );
not \U$13410 ( \13753 , \13752 );
or \U$13411 ( \13754 , \13746 , \13753 );
not \U$13412 ( \13755 , RIbb2ecb0_21);
not \U$13413 ( \13756 , \4324 );
not \U$13414 ( \13757 , \13756 );
or \U$13415 ( \13758 , \13755 , \13757 );
nand \U$13416 ( \13759 , \4086 , \2249 );
nand \U$13417 ( \13760 , \13758 , \13759 );
nand \U$13418 ( \13761 , \13760 , \2077 );
nand \U$13419 ( \13762 , \13754 , \13761 );
and \U$13420 ( \13763 , \13745 , \13762 );
and \U$13421 ( \13764 , \13725 , \13744 );
or \U$13422 ( \13765 , \13763 , \13764 );
xor \U$13423 ( \13766 , \13715 , \13765 );
not \U$13424 ( \13767 , \9099 );
not \U$13425 ( \13768 , \13326 );
or \U$13426 ( \13769 , \13767 , \13768 );
and \U$13427 ( \13770 , \1686 , RIbb2e260_43);
not \U$13428 ( \13771 , \1686 );
not \U$13429 ( \13772 , RIbb2e260_43);
and \U$13430 ( \13773 , \13771 , \13772 );
or \U$13431 ( \13774 , \13770 , \13773 );
nand \U$13432 ( \13775 , \13774 , \9098 );
nand \U$13433 ( \13776 , \13769 , \13775 );
not \U$13434 ( \13777 , \2941 );
not \U$13435 ( \13778 , \13292 );
or \U$13436 ( \13779 , \13777 , \13778 );
and \U$13437 ( \13780 , \3341 , \9169 );
not \U$13438 ( \13781 , \3341 );
and \U$13439 ( \13782 , \13781 , RIbb2e800_31);
or \U$13440 ( \13783 , \13780 , \13782 );
nand \U$13441 ( \13784 , \13783 , \2939 );
nand \U$13442 ( \13785 , \13779 , \13784 );
xor \U$13443 ( \13786 , \13776 , \13785 );
not \U$13444 ( \13787 , \2925 );
not \U$13445 ( \13788 , \13418 );
or \U$13446 ( \13789 , \13787 , \13788 );
not \U$13447 ( \13790 , RIbb2e8f0_29);
not \U$13448 ( \13791 , \3141 );
or \U$13449 ( \13792 , \13790 , \13791 );
nand \U$13450 ( \13793 , \3146 , \3440 );
nand \U$13451 ( \13794 , \13792 , \13793 );
nand \U$13452 ( \13795 , \13794 , \2922 );
nand \U$13453 ( \13796 , \13789 , \13795 );
and \U$13454 ( \13797 , \13786 , \13796 );
and \U$13455 ( \13798 , \13776 , \13785 );
or \U$13456 ( \13799 , \13797 , \13798 );
and \U$13457 ( \13800 , \13766 , \13799 );
and \U$13458 ( \13801 , \13715 , \13765 );
or \U$13459 ( \13802 , \13800 , \13801 );
or \U$13460 ( \13803 , \13676 , \13802 );
xor \U$13461 ( \13804 , \13548 , \13566 );
xor \U$13462 ( \13805 , \13804 , \13577 );
not \U$13463 ( \13806 , \1264 );
not \U$13464 ( \13807 , \1288 );
buf \U$13465 ( \13808 , \12346 );
not \U$13466 ( \13809 , \13808 );
not \U$13467 ( \13810 , \13809 );
or \U$13468 ( \13811 , \13807 , \13810 );
nand \U$13469 ( \13812 , \12347 , \1244 );
nand \U$13470 ( \13813 , \13811 , \13812 );
not \U$13471 ( \13814 , \13813 );
or \U$13472 ( \13815 , \13806 , \13814 );
nand \U$13473 ( \13816 , \13489 , \1294 );
nand \U$13474 ( \13817 , \13815 , \13816 );
not \U$13475 ( \13818 , \13817 );
not \U$13476 ( \13819 , \8995 );
not \U$13477 ( \13820 , \13402 );
or \U$13478 ( \13821 , \13819 , \13820 );
and \U$13479 ( \13822 , RIbb2e350_41, \8862 );
not \U$13480 ( \13823 , RIbb2e350_41);
and \U$13481 ( \13824 , \13823 , \3053 );
or \U$13482 ( \13825 , \13822 , \13824 );
nand \U$13483 ( \13826 , \13825 , \8362 );
nand \U$13484 ( \13827 , \13821 , \13826 );
xor \U$13485 ( \13828 , \13818 , \13827 );
not \U$13486 ( \13829 , \3465 );
not \U$13487 ( \13830 , \13434 );
or \U$13488 ( \13831 , \13829 , \13830 );
not \U$13489 ( \13832 , RIbb2e9e0_27);
not \U$13490 ( \13833 , \3905 );
or \U$13491 ( \13834 , \13832 , \13833 );
not \U$13492 ( \13835 , \3223 );
buf \U$13493 ( \13836 , \13835 );
not \U$13494 ( \13837 , \13836 );
nand \U$13495 ( \13838 , \13837 , \3454 );
nand \U$13496 ( \13839 , \13834 , \13838 );
nand \U$13497 ( \13840 , \13839 , \3445 );
nand \U$13498 ( \13841 , \13831 , \13840 );
and \U$13499 ( \13842 , \13828 , \13841 );
and \U$13500 ( \13843 , \13818 , \13827 );
or \U$13501 ( \13844 , \13842 , \13843 );
xor \U$13502 ( \13845 , \13805 , \13844 );
not \U$13503 ( \13846 , \998 );
not \U$13504 ( \13847 , \12793 );
or \U$13505 ( \13848 , \13846 , \13847 );
not \U$13506 ( \13849 , RIbb2f070_13);
not \U$13507 ( \13850 , \7296 );
not \U$13508 ( \13851 , \13850 );
or \U$13509 ( \13852 , \13849 , \13851 );
not \U$13510 ( \13853 , \7296 );
not \U$13511 ( \13854 , \13853 );
nand \U$13512 ( \13855 , \13854 , \3421 );
nand \U$13513 ( \13856 , \13852 , \13855 );
nand \U$13514 ( \13857 , \13856 , \916 );
nand \U$13515 ( \13858 , \13848 , \13857 );
not \U$13516 ( \13859 , \1077 );
not \U$13517 ( \13860 , \12805 );
or \U$13518 ( \13861 , \13859 , \13860 );
not \U$13519 ( \13862 , RIbb2f160_11);
not \U$13520 ( \13863 , \8630 );
not \U$13521 ( \13864 , \13863 );
or \U$13522 ( \13865 , \13862 , \13864 );
buf \U$13523 ( \13866 , \8630 );
nand \U$13524 ( \13867 , \13866 , \1048 );
nand \U$13525 ( \13868 , \13865 , \13867 );
nand \U$13526 ( \13869 , \13868 , \1011 );
nand \U$13527 ( \13870 , \13861 , \13869 );
xor \U$13528 ( \13871 , \13858 , \13870 );
not \U$13529 ( \13872 , \1517 );
not \U$13530 ( \13873 , \13231 );
or \U$13531 ( \13874 , \13872 , \13873 );
not \U$13532 ( \13875 , \6603 );
buf \U$13533 ( \13876 , \13875 );
and \U$13534 ( \13877 , RIbb2ef80_15, \13876 );
not \U$13535 ( \13878 , RIbb2ef80_15);
not \U$13536 ( \13879 , \8338 );
and \U$13537 ( \13880 , \13878 , \13879 );
or \U$13538 ( \13881 , \13877 , \13880 );
nand \U$13539 ( \13882 , \13881 , \1445 );
nand \U$13540 ( \13883 , \13874 , \13882 );
xor \U$13541 ( \13884 , \13871 , \13883 );
and \U$13542 ( \13885 , \13845 , \13884 );
and \U$13543 ( \13886 , \13805 , \13844 );
or \U$13544 ( \13887 , \13885 , \13886 );
nand \U$13545 ( \13888 , \13803 , \13887 );
nand \U$13546 ( \13889 , \13676 , \13802 );
nand \U$13547 ( \13890 , \13888 , \13889 );
and \U$13548 ( \13891 , \13588 , \13890 );
and \U$13549 ( \13892 , \13456 , \13587 );
or \U$13550 ( \13893 , \13891 , \13892 );
not \U$13551 ( \13894 , \13893 );
or \U$13552 ( \13895 , \13448 , \13894 );
not \U$13553 ( \13896 , \2980 );
and \U$13554 ( \13897 , RIbb2ead0_25, \12707 );
not \U$13555 ( \13898 , RIbb2ead0_25);
and \U$13556 ( \13899 , \13898 , \7021 );
or \U$13557 ( \13900 , \13897 , \13899 );
not \U$13558 ( \13901 , \13900 );
or \U$13559 ( \13902 , \13896 , \13901 );
not \U$13560 ( \13903 , \13835 );
not \U$13561 ( \13904 , \13903 );
and \U$13562 ( \13905 , RIbb2ead0_25, \13904 );
not \U$13563 ( \13906 , RIbb2ead0_25);
and \U$13564 ( \13907 , \13906 , \13837 );
or \U$13565 ( \13908 , \13905 , \13907 );
nand \U$13566 ( \13909 , \13908 , \2963 );
nand \U$13567 ( \13910 , \13902 , \13909 );
xor \U$13568 ( \13911 , \13817 , \13910 );
not \U$13569 ( \13912 , \1077 );
not \U$13570 ( \13913 , \13868 );
or \U$13571 ( \13914 , \13912 , \13913 );
not \U$13572 ( \13915 , RIbb2f160_11);
not \U$13573 ( \13916 , \9277 );
not \U$13574 ( \13917 , \13916 );
or \U$13575 ( \13918 , \13915 , \13917 );
not \U$13576 ( \13919 , \9277 );
not \U$13577 ( \13920 , \13919 );
nand \U$13578 ( \13921 , \13920 , \1048 );
nand \U$13579 ( \13922 , \13918 , \13921 );
nand \U$13580 ( \13923 , \13922 , \1011 );
nand \U$13581 ( \13924 , \13914 , \13923 );
not \U$13582 ( \13925 , \1570 );
not \U$13583 ( \13926 , \13502 );
or \U$13584 ( \13927 , \13925 , \13926 );
not \U$13585 ( \13928 , RIbb2f250_9);
not \U$13586 ( \13929 , \10300 );
not \U$13587 ( \13930 , \13929 );
or \U$13588 ( \13931 , \13928 , \13930 );
nand \U$13589 ( \13932 , \10300 , \1566 );
nand \U$13590 ( \13933 , \13931 , \13932 );
nand \U$13591 ( \13934 , \13933 , \1533 );
nand \U$13592 ( \13935 , \13927 , \13934 );
nor \U$13593 ( \13936 , \13924 , \13935 );
not \U$13594 ( \13937 , \13459 );
not \U$13595 ( \13938 , \13937 );
not \U$13596 ( \13939 , \12681 );
and \U$13597 ( \13940 , \13938 , \13939 );
not \U$13598 ( \13941 , RIbb2ddb0_53);
not \U$13599 ( \13942 , \13941 );
not \U$13600 ( \13943 , \811 );
or \U$13601 ( \13944 , \13942 , \13943 );
or \U$13602 ( \13945 , \811 , \13463 );
nand \U$13603 ( \13946 , \13944 , \13945 );
and \U$13604 ( \13947 , \13946 , \13467 );
nor \U$13605 ( \13948 , \13940 , \13947 );
or \U$13606 ( \13949 , \13936 , \13948 );
nand \U$13607 ( \13950 , \13924 , \13935 );
nand \U$13608 ( \13951 , \13949 , \13950 );
and \U$13609 ( \13952 , \13911 , \13951 );
and \U$13610 ( \13953 , \13817 , \13910 );
or \U$13611 ( \13954 , \13952 , \13953 );
xor \U$13612 ( \13955 , \13469 , \13481 );
xor \U$13613 ( \13956 , \13955 , \13491 );
not \U$13614 ( \13957 , \457 );
not \U$13615 ( \13958 , \419 );
nor \U$13616 ( \13959 , \13957 , \13958 );
not \U$13617 ( \13960 , \432 );
and \U$13618 ( \13961 , \13959 , \13960 );
not \U$13619 ( \13962 , \13961 );
not \U$13620 ( \13963 , \13194 );
or \U$13621 ( \13964 , \13962 , \13963 );
not \U$13622 ( \13965 , \13960 );
not \U$13623 ( \13966 , \423 );
or \U$13624 ( \13967 , \13965 , \13966 );
nand \U$13625 ( \13968 , \13967 , \437 );
not \U$13626 ( \13969 , \13968 );
nand \U$13627 ( \13970 , \13964 , \13969 );
nand \U$13628 ( \13971 , \436 , \440 );
not \U$13629 ( \13972 , \13971 );
and \U$13630 ( \13973 , \13970 , \13972 );
not \U$13631 ( \13974 , \13970 );
and \U$13632 ( \13975 , \13974 , \13971 );
nor \U$13633 ( \13976 , \13973 , \13975 );
buf \U$13634 ( \13977 , \13976 );
not \U$13635 ( \13978 , \13977 );
not \U$13636 ( \13979 , \13978 );
buf \U$13637 ( \13980 , \13979 );
and \U$13638 ( \13981 , \13980 , \1313 );
not \U$13639 ( \13982 , \1376 );
not \U$13640 ( \13983 , \13479 );
or \U$13641 ( \13984 , \13982 , \13983 );
not \U$13642 ( \13985 , \1312 );
not \U$13643 ( \13986 , \13545 );
not \U$13644 ( \13987 , \13986 );
or \U$13645 ( \13988 , \13985 , \13987 );
buf \U$13646 ( \13989 , \13545 );
not \U$13647 ( \13990 , \1312 );
nand \U$13648 ( \13991 , \13989 , \13990 );
nand \U$13649 ( \13992 , \13988 , \13991 );
nand \U$13650 ( \13993 , \13992 , \1429 );
nand \U$13651 ( \13994 , \13984 , \13993 );
xor \U$13652 ( \13995 , \13981 , \13994 );
not \U$13653 ( \13996 , \855 );
not \U$13654 ( \13997 , \13564 );
or \U$13655 ( \13998 , \13996 , \13997 );
not \U$13656 ( \13999 , RIbb2eda0_19);
not \U$13657 ( \14000 , \9020 );
not \U$13658 ( \14001 , \14000 );
or \U$13659 ( \14002 , \13999 , \14001 );
nand \U$13660 ( \14003 , \6198 , \3251 );
nand \U$13661 ( \14004 , \14002 , \14003 );
nand \U$13662 ( \14005 , \14004 , \853 );
nand \U$13663 ( \14006 , \13998 , \14005 );
and \U$13664 ( \14007 , \13995 , \14006 );
and \U$13665 ( \14008 , \13981 , \13994 );
or \U$13666 ( \14009 , \14007 , \14008 );
xor \U$13667 ( \14010 , \13956 , \14009 );
not \U$13668 ( \14011 , \1445 );
and \U$13669 ( \14012 , RIbb2ef80_15, \6938 );
not \U$13670 ( \14013 , RIbb2ef80_15);
and \U$13671 ( \14014 , \14013 , \6937 );
or \U$13672 ( \14015 , \14012 , \14014 );
not \U$13673 ( \14016 , \14015 );
or \U$13674 ( \14017 , \14011 , \14016 );
nand \U$13675 ( \14018 , \1517 , \13881 );
nand \U$13676 ( \14019 , \14017 , \14018 );
not \U$13677 ( \14020 , \14019 );
not \U$13678 ( \14021 , \14020 );
not \U$13679 ( \14022 , \916 );
not \U$13680 ( \14023 , RIbb2f070_13);
buf \U$13681 ( \14024 , \8318 );
not \U$13682 ( \14025 , \14024 );
not \U$13683 ( \14026 , \14025 );
or \U$13684 ( \14027 , \14023 , \14026 );
nand \U$13685 ( \14028 , \9818 , \3421 );
nand \U$13686 ( \14029 , \14027 , \14028 );
not \U$13687 ( \14030 , \14029 );
or \U$13688 ( \14031 , \14022 , \14030 );
nand \U$13689 ( \14032 , \13856 , \998 );
nand \U$13690 ( \14033 , \14031 , \14032 );
not \U$13691 ( \14034 , \14033 );
not \U$13692 ( \14035 , \14034 );
or \U$13693 ( \14036 , \14021 , \14035 );
not \U$13694 ( \14037 , \836 );
not \U$13695 ( \14038 , \13573 );
or \U$13696 ( \14039 , \14037 , \14038 );
not \U$13697 ( \14040 , RIbb2ee90_17);
not \U$13698 ( \14041 , \5954 );
not \U$13699 ( \14042 , \14041 );
or \U$13700 ( \14043 , \14040 , \14042 );
nand \U$13701 ( \14044 , \7308 , \2240 );
nand \U$13702 ( \14045 , \14043 , \14044 );
nand \U$13703 ( \14046 , \14045 , \832 );
nand \U$13704 ( \14047 , \14039 , \14046 );
nand \U$13705 ( \14048 , \14036 , \14047 );
nand \U$13706 ( \14049 , \14033 , \14019 );
nand \U$13707 ( \14050 , \14048 , \14049 );
and \U$13708 ( \14051 , \14010 , \14050 );
and \U$13709 ( \14052 , \13956 , \14009 );
or \U$13710 ( \14053 , \14051 , \14052 );
xor \U$13711 ( \14054 , \13954 , \14053 );
xor \U$13712 ( \14055 , \13494 , \13532 );
xor \U$13713 ( \14056 , \14055 , \13580 );
and \U$13714 ( \14057 , \14054 , \14056 );
and \U$13715 ( \14058 , \13954 , \14053 );
or \U$13716 ( \14059 , \14057 , \14058 );
xor \U$13717 ( \14060 , \13264 , \13274 );
xor \U$13718 ( \14061 , \14060 , \13442 );
xor \U$13719 ( \14062 , \14059 , \14061 );
xor \U$13720 ( \14063 , \13858 , \13870 );
and \U$13721 ( \14064 , \14063 , \13883 );
and \U$13722 ( \14065 , \13858 , \13870 );
or \U$13723 ( \14066 , \14064 , \14065 );
buf \U$13724 ( \14067 , \12774 );
not \U$13725 ( \14068 , \14067 );
not \U$13726 ( \14069 , \13717 );
or \U$13727 ( \14070 , \14068 , \14069 );
nand \U$13728 ( \14071 , \12779 , \12692 );
nand \U$13729 ( \14072 , \14070 , \14071 );
not \U$13730 ( \14073 , \12965 );
not \U$13731 ( \14074 , RIbb2e080_47);
not \U$13732 ( \14075 , \992 );
or \U$13733 ( \14076 , \14074 , \14075 );
nand \U$13734 ( \14077 , \987 , \10113 );
nand \U$13735 ( \14078 , \14076 , \14077 );
not \U$13736 ( \14079 , \14078 );
or \U$13737 ( \14080 , \14073 , \14079 );
nand \U$13738 ( \14081 , \13604 , \11176 );
nand \U$13739 ( \14082 , \14080 , \14081 );
xor \U$13740 ( \14083 , \14072 , \14082 );
not \U$13741 ( \14084 , \6242 );
not \U$13742 ( \14085 , \12851 );
or \U$13743 ( \14086 , \14084 , \14085 );
nand \U$13744 ( \14087 , \13630 , \6251 );
nand \U$13745 ( \14088 , \14086 , \14087 );
and \U$13746 ( \14089 , \14083 , \14088 );
and \U$13747 ( \14090 , \14072 , \14082 );
or \U$13748 ( \14091 , \14089 , \14090 );
xor \U$13749 ( \14092 , \14066 , \14091 );
not \U$13750 ( \14093 , \7104 );
and \U$13751 ( \14094 , RIbb2e440_39, \8862 );
not \U$13752 ( \14095 , RIbb2e440_39);
and \U$13753 ( \14096 , \14095 , \10673 );
or \U$13754 ( \14097 , \14094 , \14096 );
not \U$13755 ( \14098 , \14097 );
or \U$13756 ( \14099 , \14093 , \14098 );
nand \U$13757 ( \14100 , \13710 , \7103 );
nand \U$13758 ( \14101 , \14099 , \14100 );
not \U$13759 ( \14102 , \3383 );
not \U$13760 ( \14103 , RIbb2ebc0_23);
not \U$13761 ( \14104 , \5962 );
or \U$13762 ( \14105 , \14103 , \14104 );
nand \U$13763 ( \14106 , \10095 , \3396 );
nand \U$13764 ( \14107 , \14105 , \14106 );
not \U$13765 ( \14108 , \14107 );
or \U$13766 ( \14109 , \14102 , \14108 );
nand \U$13767 ( \14110 , \13742 , \3406 );
nand \U$13768 ( \14111 , \14109 , \14110 );
xor \U$13769 ( \14112 , \14101 , \14111 );
not \U$13770 ( \14113 , \2078 );
not \U$13771 ( \14114 , \12867 );
or \U$13772 ( \14115 , \14113 , \14114 );
nand \U$13773 ( \14116 , \13752 , \2077 );
nand \U$13774 ( \14117 , \14115 , \14116 );
and \U$13775 ( \14118 , \14112 , \14117 );
and \U$13776 ( \14119 , \14101 , \14111 );
or \U$13777 ( \14120 , \14118 , \14119 );
xor \U$13778 ( \14121 , \14092 , \14120 );
xor \U$13779 ( \14122 , \13266 , \13268 );
xor \U$13780 ( \14123 , \14122 , \13271 );
xor \U$13781 ( \14124 , \14121 , \14123 );
xor \U$13782 ( \14125 , \13294 , \13312 );
xor \U$13783 ( \14126 , \14125 , \13328 );
xor \U$13784 ( \14127 , \14101 , \14111 );
xor \U$13785 ( \14128 , \14127 , \14117 );
xor \U$13786 ( \14129 , \14126 , \14128 );
xor \U$13787 ( \14130 , \13384 , \13364 );
xor \U$13788 ( \14131 , \14130 , \13346 );
and \U$13789 ( \14132 , \14129 , \14131 );
and \U$13790 ( \14133 , \14126 , \14128 );
or \U$13791 ( \14134 , \14132 , \14133 );
and \U$13792 ( \14135 , \14124 , \14134 );
and \U$13793 ( \14136 , \14121 , \14123 );
or \U$13794 ( \14137 , \14135 , \14136 );
and \U$13795 ( \14138 , \14062 , \14137 );
and \U$13796 ( \14139 , \14059 , \14061 );
or \U$13797 ( \14140 , \14138 , \14139 );
not \U$13798 ( \14141 , \13893 );
nand \U$13799 ( \14142 , \14141 , \13446 );
nand \U$13800 ( \14143 , \14140 , \14142 );
nand \U$13801 ( \14144 , \13895 , \14143 );
not \U$13802 ( \14145 , \13445 );
or \U$13803 ( \14146 , \13261 , \13259 );
not \U$13804 ( \14147 , \14146 );
or \U$13805 ( \14148 , \14145 , \14147 );
nand \U$13806 ( \14149 , \13261 , \13259 );
nand \U$13807 ( \14150 , \14148 , \14149 );
xor \U$13808 ( \14151 , \13166 , \13170 );
xnor \U$13809 ( \14152 , \14151 , \13245 );
xor \U$13810 ( \14153 , \14150 , \14152 );
xor \U$13811 ( \14154 , \13458 , \13583 );
and \U$13812 ( \14155 , \14154 , \13586 );
and \U$13813 ( \14156 , \13458 , \13583 );
or \U$13814 ( \14157 , \14155 , \14156 );
not \U$13815 ( \14158 , \12167 );
not \U$13816 ( \14159 , \13310 );
or \U$13817 ( \14160 , \14158 , \14159 );
nand \U$13818 ( \14161 , \12563 , \12169 );
nand \U$13819 ( \14162 , \14160 , \14161 );
not \U$13820 ( \14163 , \855 );
not \U$13821 ( \14164 , \12581 );
or \U$13822 ( \14165 , \14163 , \14164 );
nand \U$13823 ( \14166 , \13556 , \853 );
nand \U$13824 ( \14167 , \14165 , \14166 );
xor \U$13825 ( \14168 , \14162 , \14167 );
not \U$13826 ( \14169 , \4712 );
not \U$13827 ( \14170 , \13344 );
or \U$13828 ( \14171 , \14169 , \14170 );
nand \U$13829 ( \14172 , \12048 , \5845 );
nand \U$13830 ( \14173 , \14171 , \14172 );
and \U$13831 ( \14174 , \14168 , \14173 );
and \U$13832 ( \14175 , \14162 , \14167 );
or \U$13833 ( \14176 , \14174 , \14175 );
not \U$13834 ( \14177 , \2940 );
not \U$13835 ( \14178 , \13282 );
or \U$13836 ( \14179 , \14177 , \14178 );
nand \U$13837 ( \14180 , \11969 , \3613 );
nand \U$13838 ( \14181 , \14179 , \14180 );
not \U$13839 ( \14182 , \11176 );
not \U$13840 ( \14183 , \14078 );
or \U$13841 ( \14184 , \14182 , \14183 );
nand \U$13842 ( \14185 , \11953 , \11177 );
nand \U$13843 ( \14186 , \14184 , \14185 );
xor \U$13844 ( \14187 , \14181 , \14186 );
not \U$13845 ( \14188 , \2922 );
not \U$13846 ( \14189 , \13410 );
or \U$13847 ( \14190 , \14188 , \14189 );
nand \U$13848 ( \14191 , \12060 , \2925 );
nand \U$13849 ( \14192 , \14190 , \14191 );
and \U$13850 ( \14193 , \14187 , \14192 );
and \U$13851 ( \14194 , \14181 , \14186 );
or \U$13852 ( \14195 , \14193 , \14194 );
xor \U$13853 ( \14196 , \14176 , \14195 );
not \U$13854 ( \14197 , \10449 );
not \U$13855 ( \14198 , \13319 );
or \U$13856 ( \14199 , \14197 , \14198 );
nand \U$13857 ( \14200 , \11986 , \10451 );
nand \U$13858 ( \14201 , \14199 , \14200 );
not \U$13859 ( \14202 , \10119 );
not \U$13860 ( \14203 , \12005 );
or \U$13861 ( \14204 , \14202 , \14203 );
nand \U$13862 ( \14205 , \13382 , \10117 );
nand \U$13863 ( \14206 , \14204 , \14205 );
xor \U$13864 ( \14207 , \14201 , \14206 );
not \U$13865 ( \14208 , \4791 );
not \U$13866 ( \14209 , \12021 );
or \U$13867 ( \14210 , \14208 , \14209 );
nand \U$13868 ( \14211 , \3887 , \13362 );
nand \U$13869 ( \14212 , \14210 , \14211 );
and \U$13870 ( \14213 , \14207 , \14212 );
and \U$13871 ( \14214 , \14201 , \14206 );
or \U$13872 ( \14215 , \14213 , \14214 );
xor \U$13873 ( \14216 , \14196 , \14215 );
not \U$13874 ( \14217 , \12908 );
not \U$13875 ( \14218 , \12903 );
or \U$13876 ( \14219 , \14217 , \14218 );
nand \U$13877 ( \14220 , \12902 , \12879 );
nand \U$13878 ( \14221 , \14219 , \14220 );
and \U$13879 ( \14222 , \14221 , \12907 );
not \U$13880 ( \14223 , \14221 );
not \U$13881 ( \14224 , \12907 );
and \U$13882 ( \14225 , \14223 , \14224 );
nor \U$13883 ( \14226 , \14222 , \14225 );
or \U$13884 ( \14227 , \14216 , \14226 );
not \U$13885 ( \14228 , \12352 );
not \U$13886 ( \14229 , \8361 );
not \U$13887 ( \14230 , \13394 );
or \U$13888 ( \14231 , \14229 , \14230 );
nand \U$13889 ( \14232 , \12075 , \8995 );
nand \U$13890 ( \14233 , \14231 , \14232 );
xor \U$13891 ( \14234 , \14228 , \14233 );
not \U$13892 ( \14235 , \3445 );
not \U$13893 ( \14236 , \13427 );
or \U$13894 ( \14237 , \14235 , \14236 );
nand \U$13895 ( \14238 , \12092 , \3465 );
nand \U$13896 ( \14239 , \14237 , \14238 );
and \U$13897 ( \14240 , \14234 , \14239 );
and \U$13898 ( \14241 , \14228 , \14233 );
or \U$13899 ( \14242 , \14240 , \14241 );
xor \U$13900 ( \14243 , \12528 , \12537 );
xor \U$13901 ( \14244 , \14243 , \12553 );
xor \U$13902 ( \14245 , \14242 , \14244 );
not \U$13903 ( \14246 , \2963 );
not \U$13904 ( \14247 , \12377 );
or \U$13905 ( \14248 , \14246 , \14247 );
nand \U$13906 ( \14249 , \13908 , \2980 );
nand \U$13907 ( \14250 , \14248 , \14249 );
not \U$13908 ( \14251 , \8445 );
not \U$13909 ( \14252 , \14097 );
or \U$13910 ( \14253 , \14251 , \14252 );
nand \U$13911 ( \14254 , \12363 , \8450 );
nand \U$13912 ( \14255 , \14253 , \14254 );
xor \U$13913 ( \14256 , \14250 , \14255 );
not \U$13914 ( \14257 , \3406 );
not \U$13915 ( \14258 , \14107 );
or \U$13916 ( \14259 , \14257 , \14258 );
nand \U$13917 ( \14260 , \13185 , \3383 );
nand \U$13918 ( \14261 , \14259 , \14260 );
and \U$13919 ( \14262 , \14256 , \14261 );
and \U$13920 ( \14263 , \14250 , \14255 );
or \U$13921 ( \14264 , \14262 , \14263 );
xor \U$13922 ( \14265 , \14245 , \14264 );
nand \U$13923 ( \14266 , \14227 , \14265 );
nand \U$13924 ( \14267 , \14216 , \14226 );
nand \U$13925 ( \14268 , \14266 , \14267 );
xor \U$13926 ( \14269 , \14157 , \14268 );
xor \U$13927 ( \14270 , \14066 , \14091 );
and \U$13928 ( \14271 , \14270 , \14120 );
and \U$13929 ( \14272 , \14066 , \14091 );
or \U$13930 ( \14273 , \14271 , \14272 );
xor \U$13931 ( \14274 , \14228 , \14233 );
xor \U$13932 ( \14275 , \14274 , \14239 );
xor \U$13933 ( \14276 , \14201 , \14206 );
xor \U$13934 ( \14277 , \14276 , \14212 );
xor \U$13935 ( \14278 , \14275 , \14277 );
xor \U$13936 ( \14279 , \14250 , \14255 );
xor \U$13937 ( \14280 , \14279 , \14261 );
and \U$13938 ( \14281 , \14278 , \14280 );
and \U$13939 ( \14282 , \14275 , \14277 );
or \U$13940 ( \14283 , \14281 , \14282 );
xor \U$13941 ( \14284 , \14273 , \14283 );
xor \U$13942 ( \14285 , \14162 , \14167 );
xor \U$13943 ( \14286 , \14285 , \14173 );
xor \U$13944 ( \14287 , \14181 , \14186 );
xor \U$13945 ( \14288 , \14287 , \14192 );
xor \U$13946 ( \14289 , \14286 , \14288 );
xor \U$13947 ( \14290 , \12845 , \12860 );
xor \U$13948 ( \14291 , \14290 , \12871 );
and \U$13949 ( \14292 , \14289 , \14291 );
and \U$13950 ( \14293 , \14286 , \14288 );
or \U$13951 ( \14294 , \14292 , \14293 );
and \U$13952 ( \14295 , \14284 , \14294 );
and \U$13953 ( \14296 , \14273 , \14283 );
or \U$13954 ( \14297 , \14295 , \14296 );
and \U$13955 ( \14298 , \14269 , \14297 );
and \U$13956 ( \14299 , \14157 , \14268 );
or \U$13957 ( \14300 , \14298 , \14299 );
xor \U$13958 ( \14301 , \14153 , \14300 );
xor \U$13959 ( \14302 , \14144 , \14301 );
xor \U$13960 ( \14303 , \12109 , \12107 );
xnor \U$13961 ( \14304 , \14303 , \12053 );
xor \U$13962 ( \14305 , \13450 , \13452 );
and \U$13963 ( \14306 , \14305 , \13455 );
and \U$13964 ( \14307 , \13450 , \13452 );
or \U$13965 ( \14308 , \14306 , \14307 );
xor \U$13966 ( \14309 , \14304 , \14308 );
xor \U$13967 ( \14310 , \12246 , \12288 );
xor \U$13968 ( \14311 , \14310 , \12382 );
xor \U$13969 ( \14312 , \14309 , \14311 );
not \U$13970 ( \14313 , \14312 );
not \U$13971 ( \14314 , \14244 );
not \U$13972 ( \14315 , \14264 );
or \U$13973 ( \14316 , \14314 , \14315 );
or \U$13974 ( \14317 , \14264 , \14244 );
nand \U$13975 ( \14318 , \14317 , \14242 );
nand \U$13976 ( \14319 , \14316 , \14318 );
xor \U$13977 ( \14320 , \12518 , \12556 );
xor \U$13978 ( \14321 , \14320 , \12603 );
xor \U$13979 ( \14322 , \14319 , \14321 );
xor \U$13980 ( \14323 , \14176 , \14195 );
and \U$13981 ( \14324 , \14323 , \14215 );
and \U$13982 ( \14325 , \14176 , \14195 );
or \U$13983 ( \14326 , \14324 , \14325 );
xor \U$13984 ( \14327 , \14322 , \14326 );
not \U$13985 ( \14328 , \14327 );
xor \U$13986 ( \14329 , \12877 , \12911 );
xor \U$13987 ( \14330 , \14329 , \12924 );
not \U$13988 ( \14331 , \14330 );
nand \U$13989 ( \14332 , \14328 , \14331 );
not \U$13990 ( \14333 , \14332 );
or \U$13991 ( \14334 , \14313 , \14333 );
nand \U$13992 ( \14335 , \14327 , \14330 );
nand \U$13993 ( \14336 , \14334 , \14335 );
xor \U$13994 ( \14337 , \14319 , \14321 );
and \U$13995 ( \14338 , \14337 , \14326 );
and \U$13996 ( \14339 , \14319 , \14321 );
or \U$13997 ( \14340 , \14338 , \14339 );
xor \U$13998 ( \14341 , \12112 , \12243 );
xor \U$13999 ( \14342 , \14341 , \12385 );
xor \U$14000 ( \14343 , \14340 , \14342 );
xor \U$14001 ( \14344 , \14304 , \14308 );
and \U$14002 ( \14345 , \14344 , \14311 );
and \U$14003 ( \14346 , \14304 , \14308 );
or \U$14004 ( \14347 , \14345 , \14346 );
xor \U$14005 ( \14348 , \14343 , \14347 );
xor \U$14006 ( \14349 , \14336 , \14348 );
xor \U$14007 ( \14350 , \12927 , \13019 );
xor \U$14008 ( \14351 , \14350 , \13022 );
xor \U$14009 ( \14352 , \14349 , \14351 );
and \U$14010 ( \14353 , \14302 , \14352 );
and \U$14011 ( \14354 , \14144 , \14301 );
or \U$14012 ( \14355 , \14353 , \14354 );
xor \U$14013 ( \14356 , \13257 , \14355 );
xor \U$14014 ( \14357 , \14150 , \14152 );
and \U$14015 ( \14358 , \14357 , \14300 );
and \U$14016 ( \14359 , \14150 , \14152 );
or \U$14017 ( \14360 , \14358 , \14359 );
xor \U$14018 ( \14361 , \13006 , \13012 );
and \U$14019 ( \14362 , \14361 , \13017 );
and \U$14020 ( \14363 , \13006 , \13012 );
or \U$14021 ( \14364 , \14362 , \14363 );
not \U$14022 ( \14365 , \12438 );
not \U$14023 ( \14366 , \12432 );
or \U$14024 ( \14367 , \14365 , \14366 );
nand \U$14025 ( \14368 , \14367 , \12426 );
nand \U$14026 ( \14369 , \12431 , \12437 );
nand \U$14027 ( \14370 , \14368 , \14369 );
xor \U$14028 ( \14371 , \13101 , \13106 );
and \U$14029 ( \14372 , \14371 , \13112 );
and \U$14030 ( \14373 , \13101 , \13106 );
or \U$14031 ( \14374 , \14372 , \14373 );
xor \U$14032 ( \14375 , \14370 , \14374 );
xor \U$14033 ( \14376 , \13052 , \13057 );
and \U$14034 ( \14377 , \14376 , \13063 );
and \U$14035 ( \14378 , \13052 , \13057 );
or \U$14036 ( \14379 , \14377 , \14378 );
xnor \U$14037 ( \14380 , \14375 , \14379 );
not \U$14038 ( \14381 , \14380 );
xor \U$14039 ( \14382 , \14364 , \14381 );
not \U$14040 ( \14383 , \13162 );
not \U$14041 ( \14384 , \13140 );
or \U$14042 ( \14385 , \14383 , \14384 );
nand \U$14043 ( \14386 , \14385 , \13113 );
not \U$14044 ( \14387 , \13140 );
nand \U$14045 ( \14388 , \14387 , \13161 );
nand \U$14046 ( \14389 , \14386 , \14388 );
xor \U$14047 ( \14390 , \14382 , \14389 );
xor \U$14048 ( \14391 , \13149 , \13154 );
and \U$14049 ( \14392 , \14391 , \13160 );
and \U$14050 ( \14393 , \13149 , \13154 );
or \U$14051 ( \14394 , \14392 , \14393 );
xor \U$14052 ( \14395 , \11728 , \11738 );
xor \U$14053 ( \14396 , \14395 , \11749 );
xor \U$14054 ( \14397 , \14394 , \14396 );
xor \U$14055 ( \14398 , \11762 , \11772 );
xor \U$14056 ( \14399 , \14398 , \11783 );
xnor \U$14057 ( \14400 , \14397 , \14399 );
xor \U$14058 ( \14401 , \11658 , \11668 );
xor \U$14059 ( \14402 , \14401 , \11679 );
xor \U$14060 ( \14403 , \11816 , \11826 );
xor \U$14061 ( \14404 , \14403 , \11836 );
not \U$14062 ( \14405 , \14404 );
and \U$14063 ( \14406 , \14402 , \14405 );
not \U$14064 ( \14407 , \14402 );
and \U$14065 ( \14408 , \14407 , \14404 );
or \U$14066 ( \14409 , \14406 , \14408 );
xor \U$14067 ( \14410 , \11613 , \11622 );
xor \U$14068 ( \14411 , \14410 , \11633 );
and \U$14069 ( \14412 , \14409 , \14411 );
not \U$14070 ( \14413 , \14409 );
not \U$14071 ( \14414 , \14411 );
and \U$14072 ( \14415 , \14413 , \14414 );
nor \U$14073 ( \14416 , \14412 , \14415 );
xnor \U$14074 ( \14417 , \14400 , \14416 );
not \U$14075 ( \14418 , \13136 );
not \U$14076 ( \14419 , \13126 );
or \U$14077 ( \14420 , \14418 , \14419 );
nand \U$14078 ( \14421 , \14420 , \13119 );
nand \U$14079 ( \14422 , \13125 , \13135 );
nand \U$14080 ( \14423 , \14421 , \14422 );
not \U$14081 ( \14424 , \11541 );
not \U$14082 ( \14425 , \11546 );
or \U$14083 ( \14426 , \14424 , \14425 );
nand \U$14084 ( \14427 , \11544 , \11529 );
nand \U$14085 ( \14428 , \14426 , \14427 );
not \U$14086 ( \14429 , \11558 );
and \U$14087 ( \14430 , \14428 , \14429 );
not \U$14088 ( \14431 , \14428 );
and \U$14089 ( \14432 , \14431 , \11558 );
nor \U$14090 ( \14433 , \14430 , \14432 );
and \U$14091 ( \14434 , \14423 , \14433 );
not \U$14092 ( \14435 , \14423 );
not \U$14093 ( \14436 , \14433 );
and \U$14094 ( \14437 , \14435 , \14436 );
or \U$14095 ( \14438 , \14434 , \14437 );
xor \U$14096 ( \14439 , \11582 , \11588 );
xnor \U$14097 ( \14440 , \14439 , \11599 );
and \U$14098 ( \14441 , \14438 , \14440 );
not \U$14099 ( \14442 , \14438 );
not \U$14100 ( \14443 , \14440 );
and \U$14101 ( \14444 , \14442 , \14443 );
nor \U$14102 ( \14445 , \14441 , \14444 );
not \U$14103 ( \14446 , \14445 );
and \U$14104 ( \14447 , \14417 , \14446 );
not \U$14105 ( \14448 , \14417 );
and \U$14106 ( \14449 , \14448 , \14445 );
nor \U$14107 ( \14450 , \14447 , \14449 );
xor \U$14108 ( \14451 , \14390 , \14450 );
xor \U$14109 ( \14452 , \14340 , \14342 );
and \U$14110 ( \14453 , \14452 , \14347 );
and \U$14111 ( \14454 , \14340 , \14342 );
or \U$14112 ( \14455 , \14453 , \14454 );
xor \U$14113 ( \14456 , \14451 , \14455 );
xor \U$14114 ( \14457 , \14360 , \14456 );
xor \U$14115 ( \14458 , \14336 , \14348 );
and \U$14116 ( \14459 , \14458 , \14351 );
and \U$14117 ( \14460 , \14336 , \14348 );
or \U$14118 ( \14461 , \14459 , \14460 );
xor \U$14119 ( \14462 , \14457 , \14461 );
xor \U$14120 ( \14463 , \14356 , \14462 );
and \U$14121 ( \14464 , \14327 , \14330 );
not \U$14122 ( \14465 , \14327 );
and \U$14123 ( \14466 , \14465 , \14331 );
nor \U$14124 ( \14467 , \14464 , \14466 );
and \U$14125 ( \14468 , \14467 , \14312 );
not \U$14126 ( \14469 , \14467 );
not \U$14127 ( \14470 , \14312 );
and \U$14128 ( \14471 , \14469 , \14470 );
nor \U$14129 ( \14472 , \14468 , \14471 );
xor \U$14130 ( \14473 , \14157 , \14268 );
xor \U$14131 ( \14474 , \14473 , \14297 );
xor \U$14132 ( \14475 , \14472 , \14474 );
xor \U$14133 ( \14476 , \13331 , \13386 );
xor \U$14134 ( \14477 , \14476 , \13439 );
xor \U$14135 ( \14478 , \14286 , \14288 );
xor \U$14136 ( \14479 , \14478 , \14291 );
xor \U$14137 ( \14480 , \14477 , \14479 );
xor \U$14138 ( \14481 , \14275 , \14277 );
xor \U$14139 ( \14482 , \14481 , \14280 );
and \U$14140 ( \14483 , \14480 , \14482 );
and \U$14141 ( \14484 , \14477 , \14479 );
or \U$14142 ( \14485 , \14483 , \14484 );
xor \U$14143 ( \14486 , \14273 , \14283 );
xor \U$14144 ( \14487 , \14486 , \14294 );
xor \U$14145 ( \14488 , \14485 , \14487 );
xor \U$14146 ( \14489 , \14216 , \14226 );
xor \U$14147 ( \14490 , \14489 , \14265 );
and \U$14148 ( \14491 , \14488 , \14490 );
and \U$14149 ( \14492 , \14485 , \14487 );
or \U$14150 ( \14493 , \14491 , \14492 );
and \U$14151 ( \14494 , \14475 , \14493 );
and \U$14152 ( \14495 , \14472 , \14474 );
or \U$14153 ( \14496 , \14494 , \14495 );
xor \U$14154 ( \14497 , \14072 , \14082 );
xor \U$14155 ( \14498 , \14497 , \14088 );
xor \U$14156 ( \14499 , \13404 , \13420 );
xor \U$14157 ( \14500 , \14499 , \13436 );
xor \U$14158 ( \14501 , \14498 , \14500 );
not \U$14159 ( \14502 , \1393 );
not \U$14160 ( \14503 , \13977 );
not \U$14161 ( \14504 , \14503 );
or \U$14162 ( \14505 , \14502 , \14504 );
buf \U$14163 ( \14506 , \13977 );
nand \U$14164 ( \14507 , \14506 , \13990 );
nand \U$14165 ( \14508 , \14505 , \14507 );
not \U$14166 ( \14509 , \14508 );
not \U$14167 ( \14510 , \1428 );
or \U$14168 ( \14511 , \14509 , \14510 );
nand \U$14169 ( \14512 , \13992 , \1376 );
nand \U$14170 ( \14513 , \14511 , \14512 );
not \U$14171 ( \14514 , \14513 );
not \U$14172 ( \14515 , \13959 );
not \U$14173 ( \14516 , \13194 );
or \U$14174 ( \14517 , \14515 , \14516 );
not \U$14175 ( \14518 , \423 );
nand \U$14176 ( \14519 , \14517 , \14518 );
nand \U$14177 ( \14520 , \13960 , \437 );
not \U$14178 ( \14521 , \14520 );
and \U$14179 ( \14522 , \14519 , \14521 );
not \U$14180 ( \14523 , \14519 );
and \U$14181 ( \14524 , \14523 , \14520 );
nor \U$14182 ( \14525 , \14522 , \14524 );
buf \U$14183 ( \14526 , \14525 );
buf \U$14184 ( \14527 , \14526 );
not \U$14185 ( \14528 , \14527 );
not \U$14186 ( \14529 , \14528 );
nand \U$14187 ( \14530 , \14529 , \1394 );
nand \U$14188 ( \14531 , \14514 , \14530 );
not \U$14189 ( \14532 , \14531 );
not \U$14190 ( \14533 , \2078 );
not \U$14191 ( \14534 , \13760 );
or \U$14192 ( \14535 , \14533 , \14534 );
not \U$14193 ( \14536 , \4390 );
and \U$14194 ( \14537 , \14536 , RIbb2ecb0_21);
not \U$14195 ( \14538 , \14536 );
and \U$14196 ( \14539 , \14538 , \849 );
or \U$14197 ( \14540 , \14537 , \14539 );
nand \U$14198 ( \14541 , \14540 , \2077 );
nand \U$14199 ( \14542 , \14535 , \14541 );
not \U$14200 ( \14543 , \14542 );
or \U$14201 ( \14544 , \14532 , \14543 );
not \U$14202 ( \14545 , \14530 );
nand \U$14203 ( \14546 , \14545 , \14513 );
nand \U$14204 ( \14547 , \14544 , \14546 );
not \U$14205 ( \14548 , \1011 );
not \U$14206 ( \14549 , RIbb2f160_11);
buf \U$14207 ( \14550 , \13498 );
not \U$14208 ( \14551 , \14550 );
or \U$14209 ( \14552 , \14549 , \14551 );
not \U$14210 ( \14553 , \14550 );
nand \U$14211 ( \14554 , \14553 , \1048 );
nand \U$14212 ( \14555 , \14552 , \14554 );
not \U$14213 ( \14556 , \14555 );
or \U$14214 ( \14557 , \14548 , \14556 );
nand \U$14215 ( \14558 , \13922 , \1077 );
nand \U$14216 ( \14559 , \14557 , \14558 );
not \U$14217 ( \14560 , \14559 );
not \U$14218 ( \14561 , \1533 );
not \U$14219 ( \14562 , RIbb2f250_9);
not \U$14220 ( \14563 , \10764 );
not \U$14221 ( \14564 , \14563 );
or \U$14222 ( \14565 , \14562 , \14564 );
nand \U$14223 ( \14566 , \10764 , \1554 );
nand \U$14224 ( \14567 , \14565 , \14566 );
not \U$14225 ( \14568 , \14567 );
or \U$14226 ( \14569 , \14561 , \14568 );
nand \U$14227 ( \14570 , \13933 , \1570 );
nand \U$14228 ( \14571 , \14569 , \14570 );
not \U$14229 ( \14572 , \14571 );
or \U$14230 ( \14573 , \14560 , \14572 );
not \U$14231 ( \14574 , \14559 );
not \U$14232 ( \14575 , \14574 );
not \U$14233 ( \14576 , \14571 );
not \U$14234 ( \14577 , \14576 );
or \U$14235 ( \14578 , \14575 , \14577 );
not \U$14236 ( \14579 , \998 );
not \U$14237 ( \14580 , \14029 );
or \U$14238 ( \14581 , \14579 , \14580 );
not \U$14239 ( \14582 , RIbb2f070_13);
not \U$14240 ( \14583 , \10175 );
or \U$14241 ( \14584 , \14582 , \14583 );
nand \U$14242 ( \14585 , \13866 , \3421 );
nand \U$14243 ( \14586 , \14584 , \14585 );
nand \U$14244 ( \14587 , \14586 , \916 );
nand \U$14245 ( \14588 , \14581 , \14587 );
nand \U$14246 ( \14589 , \14578 , \14588 );
nand \U$14247 ( \14590 , \14573 , \14589 );
xor \U$14248 ( \14591 , \14547 , \14590 );
xor \U$14249 ( \14592 , \13981 , \13994 );
xor \U$14250 ( \14593 , \14592 , \14006 );
and \U$14251 ( \14594 , \14591 , \14593 );
and \U$14252 ( \14595 , \14547 , \14590 );
or \U$14253 ( \14596 , \14594 , \14595 );
and \U$14254 ( \14597 , \14501 , \14596 );
and \U$14255 ( \14598 , \14498 , \14500 );
or \U$14256 ( \14599 , \14597 , \14598 );
xor \U$14257 ( \14600 , \13817 , \13910 );
xor \U$14258 ( \14601 , \14600 , \13951 );
not \U$14259 ( \14602 , RIbb2dbd0_57);
and \U$14260 ( \14603 , \14602 , RIbb2dc48_56);
not \U$14261 ( \14604 , RIbb2dc48_56);
and \U$14262 ( \14605 , \14604 , RIbb2dbd0_57);
nor \U$14263 ( \14606 , \14603 , \14605 );
not \U$14264 ( \14607 , \14606 );
and \U$14265 ( \14608 , RIbb2dcc0_55, RIbb2dc48_56);
not \U$14266 ( \14609 , RIbb2dcc0_55);
and \U$14267 ( \14610 , \14609 , \14604 );
nor \U$14268 ( \14611 , \14608 , \14610 );
and \U$14269 ( \14612 , \14606 , \14611 );
buf \U$14270 ( \14613 , \14612 );
not \U$14271 ( \14614 , \14613 );
not \U$14272 ( \14615 , \14614 );
or \U$14273 ( \14616 , \14607 , \14615 );
nand \U$14274 ( \14617 , \14616 , RIbb2dcc0_55);
not \U$14275 ( \14618 , \1294 );
not \U$14276 ( \14619 , \13813 );
or \U$14277 ( \14620 , \14618 , \14619 );
not \U$14278 ( \14621 , \1288 );
not \U$14279 ( \14622 , \13475 );
or \U$14280 ( \14623 , \14621 , \14622 );
not \U$14281 ( \14624 , \13210 );
not \U$14282 ( \14625 , \14624 );
nand \U$14283 ( \14626 , \14625 , \1244 );
nand \U$14284 ( \14627 , \14623 , \14626 );
nand \U$14285 ( \14628 , \14627 , \1264 );
nand \U$14286 ( \14629 , \14620 , \14628 );
xor \U$14287 ( \14630 , \14617 , \14629 );
not \U$14288 ( \14631 , \1147 );
not \U$14289 ( \14632 , \13684 );
or \U$14290 ( \14633 , \14631 , \14632 );
not \U$14291 ( \14634 , RIbb2f430_5);
not \U$14292 ( \14635 , \12322 );
not \U$14293 ( \14636 , \14635 );
not \U$14294 ( \14637 , \14636 );
or \U$14295 ( \14638 , \14634 , \14637 );
nand \U$14296 ( \14639 , \14635 , \1898 );
nand \U$14297 ( \14640 , \14638 , \14639 );
nand \U$14298 ( \14641 , \14640 , \1089 );
nand \U$14299 ( \14642 , \14633 , \14641 );
and \U$14300 ( \14643 , \14630 , \14642 );
and \U$14301 ( \14644 , \14617 , \14629 );
or \U$14302 ( \14645 , \14643 , \14644 );
not \U$14303 ( \14646 , \2963 );
not \U$14304 ( \14647 , \13900 );
or \U$14305 ( \14648 , \14646 , \14647 );
and \U$14306 ( \14649 , RIbb2ead0_25, \5962 );
not \U$14307 ( \14650 , RIbb2ead0_25);
and \U$14308 ( \14651 , \14650 , \10095 );
or \U$14309 ( \14652 , \14649 , \14651 );
nand \U$14310 ( \14653 , \14652 , \2980 );
nand \U$14311 ( \14654 , \14648 , \14653 );
xor \U$14312 ( \14655 , \14645 , \14654 );
not \U$14313 ( \14656 , \855 );
not \U$14314 ( \14657 , \14004 );
or \U$14315 ( \14658 , \14656 , \14657 );
not \U$14316 ( \14659 , RIbb2eda0_19);
not \U$14317 ( \14660 , \6231 );
or \U$14318 ( \14661 , \14659 , \14660 );
nand \U$14319 ( \14662 , \8387 , \1776 );
nand \U$14320 ( \14663 , \14661 , \14662 );
nand \U$14321 ( \14664 , \14663 , \853 );
nand \U$14322 ( \14665 , \14658 , \14664 );
not \U$14323 ( \14666 , \1517 );
not \U$14324 ( \14667 , \14015 );
or \U$14325 ( \14668 , \14666 , \14667 );
not \U$14326 ( \14669 , RIbb2ef80_15);
not \U$14327 ( \14670 , \9070 );
or \U$14328 ( \14671 , \14669 , \14670 );
not \U$14329 ( \14672 , \7296 );
not \U$14330 ( \14673 , \14672 );
nand \U$14331 ( \14674 , \14673 , \2356 );
nand \U$14332 ( \14675 , \14671 , \14674 );
nand \U$14333 ( \14676 , \14675 , \1445 );
nand \U$14334 ( \14677 , \14668 , \14676 );
nor \U$14335 ( \14678 , \14665 , \14677 );
not \U$14336 ( \14679 , \832 );
not \U$14337 ( \14680 , RIbb2ee90_17);
not \U$14338 ( \14681 , \8338 );
or \U$14339 ( \14682 , \14680 , \14681 );
nand \U$14340 ( \14683 , \6604 , \822 );
nand \U$14341 ( \14684 , \14682 , \14683 );
not \U$14342 ( \14685 , \14684 );
or \U$14343 ( \14686 , \14679 , \14685 );
nand \U$14344 ( \14687 , \14045 , \836 );
nand \U$14345 ( \14688 , \14686 , \14687 );
not \U$14346 ( \14689 , \14688 );
or \U$14347 ( \14690 , \14678 , \14689 );
nand \U$14348 ( \14691 , \14665 , \14677 );
nand \U$14349 ( \14692 , \14690 , \14691 );
and \U$14350 ( \14693 , \14655 , \14692 );
and \U$14351 ( \14694 , \14645 , \14654 );
or \U$14352 ( \14695 , \14693 , \14694 );
xor \U$14353 ( \14696 , \14601 , \14695 );
xor \U$14354 ( \14697 , \13956 , \14009 );
xor \U$14355 ( \14698 , \14697 , \14050 );
and \U$14356 ( \14699 , \14696 , \14698 );
and \U$14357 ( \14700 , \14601 , \14695 );
or \U$14358 ( \14701 , \14699 , \14700 );
xor \U$14359 ( \14702 , \14599 , \14701 );
xor \U$14360 ( \14703 , \13954 , \14053 );
xor \U$14361 ( \14704 , \14703 , \14056 );
and \U$14362 ( \14705 , \14702 , \14704 );
and \U$14363 ( \14706 , \14599 , \14701 );
or \U$14364 ( \14707 , \14705 , \14706 );
xor \U$14365 ( \14708 , \13456 , \13587 );
xor \U$14366 ( \14709 , \14708 , \13890 );
xor \U$14367 ( \14710 , \14707 , \14709 );
not \U$14368 ( \14711 , \3886 );
not \U$14369 ( \14712 , RIbb2e710_33);
not \U$14370 ( \14713 , \13286 );
or \U$14371 ( \14714 , \14712 , \14713 );
nand \U$14372 ( \14715 , \2222 , \12019 );
nand \U$14373 ( \14716 , \14714 , \14715 );
not \U$14374 ( \14717 , \14716 );
or \U$14375 ( \14718 , \14711 , \14717 );
nand \U$14376 ( \14719 , \13646 , \4790 );
nand \U$14377 ( \14720 , \14718 , \14719 );
not \U$14378 ( \14721 , \5845 );
not \U$14379 ( \14722 , \13596 );
or \U$14380 ( \14723 , \14721 , \14722 );
not \U$14381 ( \14724 , RIbb2e620_35);
not \U$14382 ( \14725 , \1851 );
not \U$14383 ( \14726 , \14725 );
or \U$14384 ( \14727 , \14724 , \14726 );
nand \U$14385 ( \14728 , \1851 , \3866 );
nand \U$14386 ( \14729 , \14727 , \14728 );
nand \U$14387 ( \14730 , \14729 , \4712 );
nand \U$14388 ( \14731 , \14723 , \14730 );
xor \U$14389 ( \14732 , \14720 , \14731 );
not \U$14390 ( \14733 , \14067 );
not \U$14391 ( \14734 , \3450 );
and \U$14392 ( \14735 , RIbb2dea0_51, \14734 );
not \U$14393 ( \14736 , RIbb2dea0_51);
and \U$14394 ( \14737 , \14736 , \3450 );
or \U$14395 ( \14738 , \14735 , \14737 );
not \U$14396 ( \14739 , \14738 );
or \U$14397 ( \14740 , \14733 , \14739 );
nand \U$14398 ( \14741 , \13723 , \12692 );
nand \U$14399 ( \14742 , \14740 , \14741 );
and \U$14400 ( \14743 , \14732 , \14742 );
and \U$14401 ( \14744 , \14720 , \14731 );
or \U$14402 ( \14745 , \14743 , \14744 );
buf \U$14403 ( \14746 , \14745 );
not \U$14404 ( \14747 , \14746 );
not \U$14405 ( \14748 , \12167 );
xor \U$14406 ( \14749 , RIbb2df90_49, \950 );
not \U$14407 ( \14750 , \14749 );
or \U$14408 ( \14751 , \14748 , \14750 );
not \U$14409 ( \14752 , \12283 );
nand \U$14410 ( \14753 , \13668 , \14752 );
nand \U$14411 ( \14754 , \14751 , \14753 );
not \U$14412 ( \14755 , \14754 );
not \U$14413 ( \14756 , \11176 );
and \U$14414 ( \14757 , RIbb2e080_47, \1559 );
not \U$14415 ( \14758 , RIbb2e080_47);
and \U$14416 ( \14759 , \14758 , \1560 );
or \U$14417 ( \14760 , \14757 , \14759 );
not \U$14418 ( \14761 , \14760 );
or \U$14419 ( \14762 , \14756 , \14761 );
nand \U$14420 ( \14763 , \13613 , \11177 );
nand \U$14421 ( \14764 , \14762 , \14763 );
not \U$14422 ( \14765 , \14764 );
or \U$14423 ( \14766 , \14755 , \14765 );
not \U$14424 ( \14767 , \14754 );
not \U$14425 ( \14768 , \14767 );
not \U$14426 ( \14769 , \14764 );
not \U$14427 ( \14770 , \14769 );
or \U$14428 ( \14771 , \14768 , \14770 );
not \U$14429 ( \14772 , \6242 );
not \U$14430 ( \14773 , \13623 );
or \U$14431 ( \14774 , \14772 , \14773 );
not \U$14432 ( \14775 , RIbb2e530_37);
not \U$14433 ( \14776 , \1420 );
or \U$14434 ( \14777 , \14775 , \14776 );
nand \U$14435 ( \14778 , \1421 , \8701 );
nand \U$14436 ( \14779 , \14777 , \14778 );
nand \U$14437 ( \14780 , \14779 , \6251 );
nand \U$14438 ( \14781 , \14774 , \14780 );
nand \U$14439 ( \14782 , \14771 , \14781 );
nand \U$14440 ( \14783 , \14766 , \14782 );
not \U$14441 ( \14784 , \14783 );
or \U$14442 ( \14785 , \14747 , \14784 );
or \U$14443 ( \14786 , \14746 , \14783 );
not \U$14444 ( \14787 , \2922 );
not \U$14445 ( \14788 , RIbb2e8f0_29);
not \U$14446 ( \14789 , \4638 );
or \U$14447 ( \14790 , \14788 , \14789 );
not \U$14448 ( \14791 , \4637 );
not \U$14449 ( \14792 , \14791 );
nand \U$14450 ( \14793 , \14792 , \3440 );
nand \U$14451 ( \14794 , \14790 , \14793 );
not \U$14452 ( \14795 , \14794 );
or \U$14453 ( \14796 , \14787 , \14795 );
nand \U$14454 ( \14797 , \13794 , \2925 );
nand \U$14455 ( \14798 , \14796 , \14797 );
not \U$14456 ( \14799 , \14798 );
not \U$14457 ( \14800 , \2939 );
not \U$14458 ( \14801 , RIbb2e800_31);
not \U$14459 ( \14802 , \4219 );
or \U$14460 ( \14803 , \14801 , \14802 );
nand \U$14461 ( \14804 , \3166 , \2917 );
nand \U$14462 ( \14805 , \14803 , \14804 );
not \U$14463 ( \14806 , \14805 );
or \U$14464 ( \14807 , \14800 , \14806 );
nand \U$14465 ( \14808 , \13783 , \2941 );
nand \U$14466 ( \14809 , \14807 , \14808 );
buf \U$14467 ( \14810 , \14809 );
not \U$14468 ( \14811 , \14810 );
or \U$14469 ( \14812 , \14799 , \14811 );
or \U$14470 ( \14813 , \14810 , \14798 );
not \U$14471 ( \14814 , \10119 );
not \U$14472 ( \14815 , \13657 );
or \U$14473 ( \14816 , \14814 , \14815 );
not \U$14474 ( \14817 , RIbb2e170_45);
not \U$14475 ( \14818 , \1729 );
not \U$14476 ( \14819 , \14818 );
not \U$14477 ( \14820 , \14819 );
or \U$14478 ( \14821 , \14817 , \14820 );
nand \U$14479 ( \14822 , \14818 , \11065 );
nand \U$14480 ( \14823 , \14821 , \14822 );
nand \U$14481 ( \14824 , \14823 , \10599 );
nand \U$14482 ( \14825 , \14816 , \14824 );
nand \U$14483 ( \14826 , \14813 , \14825 );
nand \U$14484 ( \14827 , \14812 , \14826 );
nand \U$14485 ( \14828 , \14786 , \14827 );
nand \U$14486 ( \14829 , \14785 , \14828 );
xor \U$14487 ( \14830 , \13948 , \13935 );
xor \U$14488 ( \14831 , \14830 , \13924 );
not \U$14489 ( \14832 , \14831 );
not \U$14490 ( \14833 , \14832 );
not \U$14491 ( \14834 , \1147 );
not \U$14492 ( \14835 , \14640 );
or \U$14493 ( \14836 , \14834 , \14835 );
not \U$14494 ( \14837 , RIbb2f430_5);
not \U$14495 ( \14838 , \13808 );
not \U$14496 ( \14839 , \14838 );
not \U$14497 ( \14840 , \14839 );
not \U$14498 ( \14841 , \14840 );
or \U$14499 ( \14842 , \14837 , \14841 );
buf \U$14500 ( \14843 , \13808 );
buf \U$14501 ( \14844 , \14843 );
nand \U$14502 ( \14845 , \14844 , \1980 );
nand \U$14503 ( \14846 , \14842 , \14845 );
nand \U$14504 ( \14847 , \14846 , \1089 );
nand \U$14505 ( \14848 , \14836 , \14847 );
not \U$14506 ( \14849 , \14848 );
not \U$14507 ( \14850 , \9098 );
not \U$14508 ( \14851 , RIbb2e260_43);
not \U$14509 ( \14852 , \1641 );
or \U$14510 ( \14853 , \14851 , \14852 );
nand \U$14511 ( \14854 , \8856 , \9847 );
nand \U$14512 ( \14855 , \14853 , \14854 );
not \U$14513 ( \14856 , \14855 );
or \U$14514 ( \14857 , \14850 , \14856 );
nand \U$14515 ( \14858 , \13774 , \9099 );
nand \U$14516 ( \14859 , \14857 , \14858 );
not \U$14517 ( \14860 , \14859 );
or \U$14518 ( \14861 , \14849 , \14860 );
or \U$14519 ( \14862 , \14859 , \14848 );
not \U$14520 ( \14863 , \3465 );
not \U$14521 ( \14864 , \13839 );
or \U$14522 ( \14865 , \14863 , \14864 );
not \U$14523 ( \14866 , RIbb2e9e0_27);
not \U$14524 ( \14867 , \12707 );
or \U$14525 ( \14868 , \14866 , \14867 );
nand \U$14526 ( \14869 , \7021 , \6065 );
nand \U$14527 ( \14870 , \14868 , \14869 );
nand \U$14528 ( \14871 , \14870 , \3445 );
nand \U$14529 ( \14872 , \14865 , \14871 );
nand \U$14530 ( \14873 , \14862 , \14872 );
nand \U$14531 ( \14874 , \14861 , \14873 );
not \U$14532 ( \14875 , \14874 );
or \U$14533 ( \14876 , \14833 , \14875 );
or \U$14534 ( \14877 , \14874 , \14832 );
xor \U$14535 ( \14878 , \13686 , \13696 );
xor \U$14536 ( \14879 , \14878 , \13712 );
nand \U$14537 ( \14880 , \14877 , \14879 );
nand \U$14538 ( \14881 , \14876 , \14880 );
xor \U$14539 ( \14882 , \14829 , \14881 );
not \U$14540 ( \14883 , \1702 );
not \U$14541 ( \14884 , RIbb2f340_7);
buf \U$14542 ( \14885 , \11578 );
not \U$14543 ( \14886 , \14885 );
not \U$14544 ( \14887 , \14886 );
or \U$14545 ( \14888 , \14884 , \14887 );
nand \U$14546 ( \14889 , \14885 , \1734 );
nand \U$14547 ( \14890 , \14888 , \14889 );
not \U$14548 ( \14891 , \14890 );
or \U$14549 ( \14892 , \14883 , \14891 );
nand \U$14550 ( \14893 , \13694 , \1737 );
nand \U$14551 ( \14894 , \14892 , \14893 );
not \U$14552 ( \14895 , \8362 );
not \U$14553 ( \14896 , RIbb2e350_41);
not \U$14554 ( \14897 , \4766 );
or \U$14555 ( \14898 , \14896 , \14897 );
not \U$14556 ( \14899 , RIbb2e350_41);
nand \U$14557 ( \14900 , \14899 , \13708 );
nand \U$14558 ( \14901 , \14898 , \14900 );
not \U$14559 ( \14902 , \14901 );
or \U$14560 ( \14903 , \14895 , \14902 );
nand \U$14561 ( \14904 , \13825 , \8354 );
nand \U$14562 ( \14905 , \14903 , \14904 );
xor \U$14563 ( \14906 , \14894 , \14905 );
not \U$14564 ( \14907 , \2963 );
not \U$14565 ( \14908 , \14652 );
or \U$14566 ( \14909 , \14907 , \14908 );
and \U$14567 ( \14910 , RIbb2ead0_25, \8483 );
not \U$14568 ( \14911 , RIbb2ead0_25);
not \U$14569 ( \14912 , \13738 );
and \U$14570 ( \14913 , \14911 , \14912 );
or \U$14571 ( \14914 , \14910 , \14913 );
nand \U$14572 ( \14915 , \14914 , \2980 );
nand \U$14573 ( \14916 , \14909 , \14915 );
and \U$14574 ( \14917 , \14906 , \14916 );
and \U$14575 ( \14918 , \14894 , \14905 );
or \U$14576 ( \14919 , \14917 , \14918 );
buf \U$14577 ( \14920 , \13467 );
not \U$14578 ( \14921 , \14920 );
not \U$14579 ( \14922 , RIbb2ddb0_53);
not \U$14580 ( \14923 , \12969 );
or \U$14581 ( \14924 , \14922 , \14923 );
nand \U$14582 ( \14925 , \892 , \12681 );
nand \U$14583 ( \14926 , \14924 , \14925 );
not \U$14584 ( \14927 , \14926 );
or \U$14585 ( \14928 , \14921 , \14927 );
buf \U$14586 ( \14929 , \13459 );
buf \U$14587 ( \14930 , \14929 );
nand \U$14588 ( \14931 , \13946 , \14930 );
nand \U$14589 ( \14932 , \14928 , \14931 );
not \U$14590 ( \14933 , \8450 );
not \U$14591 ( \14934 , \13702 );
or \U$14592 ( \14935 , \14933 , \14934 );
and \U$14593 ( \14936 , RIbb2e440_39, \3990 );
not \U$14594 ( \14937 , RIbb2e440_39);
and \U$14595 ( \14938 , \14937 , \1169 );
or \U$14596 ( \14939 , \14936 , \14938 );
nand \U$14597 ( \14940 , \14939 , \7103 );
nand \U$14598 ( \14941 , \14935 , \14940 );
xor \U$14599 ( \14942 , \14932 , \14941 );
not \U$14600 ( \14943 , \3406 );
not \U$14601 ( \14944 , RIbb2ebc0_23);
not \U$14602 ( \14945 , \12577 );
or \U$14603 ( \14946 , \14944 , \14945 );
nand \U$14604 ( \14947 , \3091 , \3401 );
nand \U$14605 ( \14948 , \14946 , \14947 );
not \U$14606 ( \14949 , \14948 );
or \U$14607 ( \14950 , \14943 , \14949 );
nand \U$14608 ( \14951 , \13734 , \3383 );
nand \U$14609 ( \14952 , \14950 , \14951 );
and \U$14610 ( \14953 , \14942 , \14952 );
and \U$14611 ( \14954 , \14932 , \14941 );
or \U$14612 ( \14955 , \14953 , \14954 );
xor \U$14613 ( \14956 , \14919 , \14955 );
and \U$14614 ( \14957 , \14034 , \14020 );
not \U$14615 ( \14958 , \14034 );
and \U$14616 ( \14959 , \14958 , \14019 );
nor \U$14617 ( \14960 , \14957 , \14959 );
xor \U$14618 ( \14961 , \14960 , \14047 );
and \U$14619 ( \14962 , \14956 , \14961 );
and \U$14620 ( \14963 , \14919 , \14955 );
or \U$14621 ( \14964 , \14962 , \14963 );
and \U$14622 ( \14965 , \14882 , \14964 );
and \U$14623 ( \14966 , \14829 , \14881 );
or \U$14624 ( \14967 , \14965 , \14966 );
xor \U$14625 ( \14968 , \13715 , \13765 );
xor \U$14626 ( \14969 , \14968 , \13799 );
xor \U$14627 ( \14970 , \13805 , \13844 );
xor \U$14628 ( \14971 , \14970 , \13884 );
xor \U$14629 ( \14972 , \14969 , \14971 );
xor \U$14630 ( \14973 , \13648 , \13659 );
xor \U$14631 ( \14974 , \14973 , \13670 );
xor \U$14632 ( \14975 , \13725 , \13744 );
xor \U$14633 ( \14976 , \14975 , \13762 );
or \U$14634 ( \14977 , \14974 , \14976 );
xor \U$14635 ( \14978 , \13776 , \13785 );
xor \U$14636 ( \14979 , \14978 , \13796 );
nand \U$14637 ( \14980 , \14977 , \14979 );
nand \U$14638 ( \14981 , \14974 , \14976 );
nand \U$14639 ( \14982 , \14980 , \14981 );
and \U$14640 ( \14983 , \14972 , \14982 );
and \U$14641 ( \14984 , \14969 , \14971 );
or \U$14642 ( \14985 , \14983 , \14984 );
xor \U$14643 ( \14986 , \14967 , \14985 );
xor \U$14644 ( \14987 , \13887 , \13802 );
xor \U$14645 ( \14988 , \14987 , \13676 );
and \U$14646 ( \14989 , \14986 , \14988 );
and \U$14647 ( \14990 , \14967 , \14985 );
or \U$14648 ( \14991 , \14989 , \14990 );
and \U$14649 ( \14992 , \14710 , \14991 );
and \U$14650 ( \14993 , \14707 , \14709 );
or \U$14651 ( \14994 , \14992 , \14993 );
not \U$14652 ( \14995 , \14140 );
not \U$14653 ( \14996 , \14995 );
not \U$14654 ( \14997 , \13893 );
not \U$14655 ( \14998 , \13446 );
or \U$14656 ( \14999 , \14997 , \14998 );
or \U$14657 ( \15000 , \13893 , \13446 );
nand \U$14658 ( \15001 , \14999 , \15000 );
not \U$14659 ( \15002 , \15001 );
or \U$14660 ( \15003 , \14996 , \15002 );
or \U$14661 ( \15004 , \15001 , \14995 );
nand \U$14662 ( \15005 , \15003 , \15004 );
xor \U$14663 ( \15006 , \14994 , \15005 );
xor \U$14664 ( \15007 , \14485 , \14487 );
xor \U$14665 ( \15008 , \15007 , \14490 );
xor \U$14666 ( \15009 , \14121 , \14123 );
xor \U$14667 ( \15010 , \15009 , \14134 );
xor \U$14668 ( \15011 , \13635 , \13637 );
xor \U$14669 ( \15012 , \15011 , \13673 );
xor \U$14670 ( \15013 , \13818 , \13827 );
xor \U$14671 ( \15014 , \15013 , \13841 );
xor \U$14672 ( \15015 , \13615 , \13632 );
xor \U$14673 ( \15016 , \15015 , \13598 );
xor \U$14674 ( \15017 , \15014 , \15016 );
not \U$14675 ( \15018 , \13958 );
nand \U$14676 ( \15019 , \15018 , \422 );
not \U$14677 ( \15020 , \15019 );
not \U$14678 ( \15021 , \457 );
not \U$14679 ( \15022 , \12305 );
or \U$14680 ( \15023 , \15021 , \15022 );
nand \U$14681 ( \15024 , RIbb2be48_120, RIbb32fb8_184);
nand \U$14682 ( \15025 , \15023 , \15024 );
not \U$14683 ( \15026 , \15025 );
or \U$14684 ( \15027 , \15020 , \15026 );
or \U$14685 ( \15028 , \15025 , \15019 );
nand \U$14686 ( \15029 , \15027 , \15028 );
buf \U$14687 ( \15030 , \15029 );
not \U$14688 ( \15031 , \15030 );
not \U$14689 ( \15032 , \15031 );
and \U$14690 ( \15033 , \15032 , \1312 );
not \U$14691 ( \15034 , \1429 );
not \U$14692 ( \15035 , \1393 );
buf \U$14693 ( \15036 , \14526 );
not \U$14694 ( \15037 , \15036 );
not \U$14695 ( \15038 , \15037 );
or \U$14696 ( \15039 , \15035 , \15038 );
nand \U$14697 ( \15040 , \15036 , \1392 );
nand \U$14698 ( \15041 , \15039 , \15040 );
not \U$14699 ( \15042 , \15041 );
or \U$14700 ( \15043 , \15034 , \15042 );
nand \U$14701 ( \15044 , \14508 , \1376 );
nand \U$14702 ( \15045 , \15043 , \15044 );
xor \U$14703 ( \15046 , \15033 , \15045 );
not \U$14704 ( \15047 , \1294 );
not \U$14705 ( \15048 , \14627 );
or \U$14706 ( \15049 , \15047 , \15048 );
not \U$14707 ( \15050 , \1288 );
not \U$14708 ( \15051 , \13989 );
not \U$14709 ( \15052 , \15051 );
or \U$14710 ( \15053 , \15050 , \15052 );
not \U$14711 ( \15054 , \13545 );
not \U$14712 ( \15055 , \15054 );
nand \U$14713 ( \15056 , \15055 , \1244 );
nand \U$14714 ( \15057 , \15053 , \15056 );
nand \U$14715 ( \15058 , \15057 , \1264 );
nand \U$14716 ( \15059 , \15049 , \15058 );
and \U$14717 ( \15060 , \15046 , \15059 );
and \U$14718 ( \15061 , \15033 , \15045 );
or \U$14719 ( \15062 , \15060 , \15061 );
not \U$14720 ( \15063 , \836 );
not \U$14721 ( \15064 , \14684 );
or \U$14722 ( \15065 , \15063 , \15064 );
not \U$14723 ( \15066 , \6937 );
and \U$14724 ( \15067 , RIbb2ee90_17, \15066 );
not \U$14725 ( \15068 , RIbb2ee90_17);
and \U$14726 ( \15069 , \15068 , \12791 );
or \U$14727 ( \15070 , \15067 , \15069 );
nand \U$14728 ( \15071 , \15070 , \832 );
nand \U$14729 ( \15072 , \15065 , \15071 );
not \U$14730 ( \15073 , \15072 );
not \U$14731 ( \15074 , \2077 );
not \U$14732 ( \15075 , RIbb2ecb0_21);
not \U$14733 ( \15076 , \9023 );
or \U$14734 ( \15077 , \15075 , \15076 );
not \U$14735 ( \15078 , \14000 );
nand \U$14736 ( \15079 , \15078 , \2067 );
nand \U$14737 ( \15080 , \15077 , \15079 );
not \U$14738 ( \15081 , \15080 );
or \U$14739 ( \15082 , \15074 , \15081 );
nand \U$14740 ( \15083 , \14540 , \2078 );
nand \U$14741 ( \15084 , \15082 , \15083 );
not \U$14742 ( \15085 , \15084 );
or \U$14743 ( \15086 , \15073 , \15085 );
or \U$14744 ( \15087 , \15084 , \15072 );
not \U$14745 ( \15088 , \855 );
not \U$14746 ( \15089 , \14663 );
or \U$14747 ( \15090 , \15088 , \15089 );
not \U$14748 ( \15091 , RIbb2eda0_19);
not \U$14749 ( \15092 , \14041 );
or \U$14750 ( \15093 , \15091 , \15092 );
nand \U$14751 ( \15094 , \7308 , \1776 );
nand \U$14752 ( \15095 , \15093 , \15094 );
nand \U$14753 ( \15096 , \15095 , \853 );
nand \U$14754 ( \15097 , \15090 , \15096 );
nand \U$14755 ( \15098 , \15087 , \15097 );
nand \U$14756 ( \15099 , \15086 , \15098 );
xor \U$14757 ( \15100 , \15062 , \15099 );
not \U$14758 ( \15101 , \1011 );
not \U$14759 ( \15102 , RIbb2f160_11);
not \U$14760 ( \15103 , \13929 );
or \U$14761 ( \15104 , \15102 , \15103 );
not \U$14762 ( \15105 , \10300 );
buf \U$14763 ( \15106 , \15105 );
not \U$14764 ( \15107 , \15106 );
nand \U$14765 ( \15108 , \15107 , \1043 );
nand \U$14766 ( \15109 , \15104 , \15108 );
not \U$14767 ( \15110 , \15109 );
or \U$14768 ( \15111 , \15101 , \15110 );
nand \U$14769 ( \15112 , \14555 , \1077 );
nand \U$14770 ( \15113 , \15111 , \15112 );
not \U$14771 ( \15114 , \1517 );
not \U$14772 ( \15115 , \14675 );
or \U$14773 ( \15116 , \15114 , \15115 );
and \U$14774 ( \15117 , RIbb2ef80_15, \12210 );
not \U$14775 ( \15118 , RIbb2ef80_15);
and \U$14776 ( \15119 , \15118 , \9818 );
or \U$14777 ( \15120 , \15117 , \15119 );
nand \U$14778 ( \15121 , \15120 , \1445 );
nand \U$14779 ( \15122 , \15116 , \15121 );
xor \U$14780 ( \15123 , \15113 , \15122 );
not \U$14781 ( \15124 , \916 );
not \U$14782 ( \15125 , RIbb2f070_13);
not \U$14783 ( \15126 , \12820 );
or \U$14784 ( \15127 , \15125 , \15126 );
not \U$14785 ( \15128 , \9857 );
nand \U$14786 ( \15129 , \15128 , \1656 );
nand \U$14787 ( \15130 , \15127 , \15129 );
not \U$14788 ( \15131 , \15130 );
or \U$14789 ( \15132 , \15124 , \15131 );
nand \U$14790 ( \15133 , \14586 , \998 );
nand \U$14791 ( \15134 , \15132 , \15133 );
and \U$14792 ( \15135 , \15123 , \15134 );
and \U$14793 ( \15136 , \15113 , \15122 );
or \U$14794 ( \15137 , \15135 , \15136 );
and \U$14795 ( \15138 , \15100 , \15137 );
and \U$14796 ( \15139 , \15062 , \15099 );
or \U$14797 ( \15140 , \15138 , \15139 );
and \U$14798 ( \15141 , \15017 , \15140 );
and \U$14799 ( \15142 , \15014 , \15016 );
or \U$14800 ( \15143 , \15141 , \15142 );
xor \U$14801 ( \15144 , \15012 , \15143 );
xor \U$14802 ( \15145 , \14498 , \14500 );
xor \U$14803 ( \15146 , \15145 , \14596 );
and \U$14804 ( \15147 , \15144 , \15146 );
and \U$14805 ( \15148 , \15012 , \15143 );
or \U$14806 ( \15149 , \15147 , \15148 );
xor \U$14807 ( \15150 , \15010 , \15149 );
xor \U$14808 ( \15151 , \14126 , \14128 );
xor \U$14809 ( \15152 , \15151 , \14131 );
xor \U$14810 ( \15153 , \14601 , \14695 );
xor \U$14811 ( \15154 , \15153 , \14698 );
xor \U$14812 ( \15155 , \15152 , \15154 );
xor \U$14813 ( \15156 , \14645 , \14654 );
xor \U$14814 ( \15157 , \15156 , \14692 );
xor \U$14815 ( \15158 , \14617 , \14629 );
xor \U$14816 ( \15159 , \15158 , \14642 );
xor \U$14817 ( \15160 , \14513 , \14530 );
not \U$14818 ( \15161 , \14542 );
xor \U$14819 ( \15162 , \15160 , \15161 );
xor \U$14820 ( \15163 , \15159 , \15162 );
not \U$14821 ( \15164 , \1737 );
not \U$14822 ( \15165 , \14890 );
or \U$14823 ( \15166 , \15164 , \15165 );
not \U$14824 ( \15167 , RIbb2f340_7);
not \U$14825 ( \15168 , \12839 );
or \U$14826 ( \15169 , \15167 , \15168 );
nand \U$14827 ( \15170 , \12175 , \1734 );
nand \U$14828 ( \15171 , \15169 , \15170 );
nand \U$14829 ( \15172 , \15171 , \1702 );
nand \U$14830 ( \15173 , \15166 , \15172 );
not \U$14831 ( \15174 , \14613 );
and \U$14832 ( \15175 , RIbb2dcc0_55, \812 );
not \U$14833 ( \15176 , RIbb2dcc0_55);
and \U$14834 ( \15177 , \15176 , \811 );
or \U$14835 ( \15178 , \15175 , \15177 );
not \U$14836 ( \15179 , \15178 );
or \U$14837 ( \15180 , \15174 , \15179 );
not \U$14838 ( \15181 , \14606 );
buf \U$14839 ( \15182 , \15181 );
nand \U$14840 ( \15183 , \15182 , RIbb2dcc0_55);
nand \U$14841 ( \15184 , \15180 , \15183 );
xor \U$14842 ( \15185 , \15173 , \15184 );
not \U$14843 ( \15186 , \1533 );
not \U$14844 ( \15187 , RIbb2f250_9);
buf \U$14845 ( \15188 , \12754 );
not \U$14846 ( \15189 , \15188 );
or \U$14847 ( \15190 , \15187 , \15189 );
nand \U$14848 ( \15191 , \11144 , \1566 );
nand \U$14849 ( \15192 , \15190 , \15191 );
not \U$14850 ( \15193 , \15192 );
or \U$14851 ( \15194 , \15186 , \15193 );
nand \U$14852 ( \15195 , \1570 , \14567 );
nand \U$14853 ( \15196 , \15194 , \15195 );
and \U$14854 ( \15197 , \15185 , \15196 );
and \U$14855 ( \15198 , \15173 , \15184 );
or \U$14856 ( \15199 , \15197 , \15198 );
and \U$14857 ( \15200 , \15163 , \15199 );
and \U$14858 ( \15201 , \15159 , \15162 );
or \U$14859 ( \15202 , \15200 , \15201 );
xor \U$14860 ( \15203 , \15157 , \15202 );
xor \U$14861 ( \15204 , \14547 , \14590 );
xor \U$14862 ( \15205 , \15204 , \14593 );
and \U$14863 ( \15206 , \15203 , \15205 );
and \U$14864 ( \15207 , \15157 , \15202 );
or \U$14865 ( \15208 , \15206 , \15207 );
and \U$14866 ( \15209 , \15155 , \15208 );
and \U$14867 ( \15210 , \15152 , \15154 );
or \U$14868 ( \15211 , \15209 , \15210 );
and \U$14869 ( \15212 , \15150 , \15211 );
and \U$14870 ( \15213 , \15010 , \15149 );
or \U$14871 ( \15214 , \15212 , \15213 );
or \U$14872 ( \15215 , \15008 , \15214 );
xor \U$14873 ( \15216 , \14059 , \14061 );
xor \U$14874 ( \15217 , \15216 , \14137 );
nand \U$14875 ( \15218 , \15215 , \15217 );
nand \U$14876 ( \15219 , \15008 , \15214 );
nand \U$14877 ( \15220 , \15218 , \15219 );
and \U$14878 ( \15221 , \15006 , \15220 );
and \U$14879 ( \15222 , \14994 , \15005 );
or \U$14880 ( \15223 , \15221 , \15222 );
xor \U$14881 ( \15224 , \14496 , \15223 );
xor \U$14882 ( \15225 , \14144 , \14301 );
xor \U$14883 ( \15226 , \15225 , \14352 );
and \U$14884 ( \15227 , \15224 , \15226 );
and \U$14885 ( \15228 , \14496 , \15223 );
or \U$14886 ( \15229 , \15227 , \15228 );
or \U$14887 ( \15230 , \14463 , \15229 );
xor \U$14888 ( \15231 , \12739 , \13025 );
and \U$14889 ( \15232 , \15231 , \13256 );
and \U$14890 ( \15233 , \12739 , \13025 );
or \U$14891 ( \15234 , \15232 , \15233 );
xor \U$14892 ( \15235 , \14390 , \14450 );
and \U$14893 ( \15236 , \15235 , \14455 );
and \U$14894 ( \15237 , \14390 , \14450 );
or \U$14895 ( \15238 , \15236 , \15237 );
not \U$14896 ( \15239 , \14445 );
not \U$14897 ( \15240 , \14400 );
or \U$14898 ( \15241 , \15239 , \15240 );
nand \U$14899 ( \15242 , \15241 , \14416 );
not \U$14900 ( \15243 , \14400 );
nand \U$14901 ( \15244 , \15243 , \14446 );
nand \U$14902 ( \15245 , \15242 , \15244 );
xor \U$14903 ( \15246 , \11645 , \11647 );
xor \U$14904 ( \15247 , \15246 , \11682 );
xor \U$14905 ( \15248 , \11839 , \11841 );
xor \U$14906 ( \15249 , \15248 , \11844 );
xor \U$14907 ( \15250 , \15247 , \15249 );
xor \U$14908 ( \15251 , \11855 , \11852 );
xor \U$14909 ( \15252 , \15251 , \11859 );
xnor \U$14910 ( \15253 , \15250 , \15252 );
xor \U$14911 ( \15254 , \15245 , \15253 );
xor \U$14912 ( \15255 , \12389 , \12393 );
and \U$14913 ( \15256 , \15255 , \12411 );
and \U$14914 ( \15257 , \12389 , \12393 );
or \U$14915 ( \15258 , \15256 , \15257 );
xor \U$14916 ( \15259 , \11509 , \11519 );
xor \U$14917 ( \15260 , \15259 , \11560 );
xor \U$14918 ( \15261 , \15258 , \15260 );
buf \U$14919 ( \15262 , \14370 );
or \U$14920 ( \15263 , \15262 , \14374 );
nand \U$14921 ( \15264 , \15263 , \14379 );
nand \U$14922 ( \15265 , \14374 , \15262 );
nand \U$14923 ( \15266 , \15264 , \15265 );
xor \U$14924 ( \15267 , \15261 , \15266 );
xor \U$14925 ( \15268 , \12412 , \12416 );
and \U$14926 ( \15269 , \15268 , \12482 );
and \U$14927 ( \15270 , \12412 , \12416 );
or \U$14928 ( \15271 , \15269 , \15270 );
xor \U$14929 ( \15272 , \15267 , \15271 );
xor \U$14930 ( \15273 , \13030 , \13085 );
and \U$14931 ( \15274 , \15273 , \13098 );
and \U$14932 ( \15275 , \13030 , \13085 );
or \U$14933 ( \15276 , \15274 , \15275 );
xor \U$14934 ( \15277 , \15272 , \15276 );
xor \U$14935 ( \15278 , \15254 , \15277 );
xor \U$14936 ( \15279 , \15238 , \15278 );
xor \U$14937 ( \15280 , \12388 , \12483 );
and \U$14938 ( \15281 , \15280 , \12738 );
and \U$14939 ( \15282 , \12388 , \12483 );
or \U$14940 ( \15283 , \15281 , \15282 );
not \U$14941 ( \15284 , \13251 );
not \U$14942 ( \15285 , \13099 );
or \U$14943 ( \15286 , \15284 , \15285 );
or \U$14944 ( \15287 , \13099 , \13251 );
nand \U$14945 ( \15288 , \15287 , \13247 );
nand \U$14946 ( \15289 , \15286 , \15288 );
xor \U$14947 ( \15290 , \15283 , \15289 );
not \U$14948 ( \15291 , \14436 );
not \U$14949 ( \15292 , \14443 );
or \U$14950 ( \15293 , \15291 , \15292 );
not \U$14951 ( \15294 , \14440 );
not \U$14952 ( \15295 , \14433 );
or \U$14953 ( \15296 , \15294 , \15295 );
nand \U$14954 ( \15297 , \15296 , \14423 );
nand \U$14955 ( \15298 , \15293 , \15297 );
or \U$14956 ( \15299 , \13088 , \13097 );
nand \U$14957 ( \15300 , \15299 , \13092 );
nand \U$14958 ( \15301 , \13097 , \13088 );
nand \U$14959 ( \15302 , \15300 , \15301 );
xor \U$14960 ( \15303 , \15298 , \15302 );
xor \U$14961 ( \15304 , \11719 , \11752 );
xor \U$14962 ( \15305 , \15304 , \11786 );
xor \U$14963 ( \15306 , \15303 , \15305 );
not \U$14964 ( \15307 , \14364 );
not \U$14965 ( \15308 , \14381 );
or \U$14966 ( \15309 , \15307 , \15308 );
not \U$14967 ( \15310 , \14364 );
not \U$14968 ( \15311 , \15310 );
not \U$14969 ( \15312 , \14380 );
or \U$14970 ( \15313 , \15311 , \15312 );
nand \U$14971 ( \15314 , \15313 , \14389 );
nand \U$14972 ( \15315 , \15309 , \15314 );
and \U$14973 ( \15316 , \15306 , \15315 );
not \U$14974 ( \15317 , \15306 );
not \U$14975 ( \15318 , \15315 );
and \U$14976 ( \15319 , \15317 , \15318 );
nor \U$14977 ( \15320 , \15316 , \15319 );
not \U$14978 ( \15321 , \14396 );
not \U$14979 ( \15322 , \14399 );
or \U$14980 ( \15323 , \15321 , \15322 );
or \U$14981 ( \15324 , \14399 , \14396 );
nand \U$14982 ( \15325 , \15324 , \14394 );
nand \U$14983 ( \15326 , \15323 , \15325 );
or \U$14984 ( \15327 , \14404 , \14411 );
nand \U$14985 ( \15328 , \15327 , \14402 );
nand \U$14986 ( \15329 , \14404 , \14411 );
nand \U$14987 ( \15330 , \15328 , \15329 );
xor \U$14988 ( \15331 , \15326 , \15330 );
not \U$14989 ( \15332 , \11636 );
xnor \U$14990 ( \15333 , \11602 , \11641 );
not \U$14991 ( \15334 , \15333 );
or \U$14992 ( \15335 , \15332 , \15334 );
or \U$14993 ( \15336 , \15333 , \11636 );
nand \U$14994 ( \15337 , \15335 , \15336 );
xnor \U$14995 ( \15338 , \15331 , \15337 );
not \U$14996 ( \15339 , \15338 );
and \U$14997 ( \15340 , \15320 , \15339 );
not \U$14998 ( \15341 , \15320 );
and \U$14999 ( \15342 , \15341 , \15338 );
nor \U$15000 ( \15343 , \15340 , \15342 );
xor \U$15001 ( \15344 , \15290 , \15343 );
xor \U$15002 ( \15345 , \15279 , \15344 );
xor \U$15003 ( \15346 , \15234 , \15345 );
xor \U$15004 ( \15347 , \14360 , \14456 );
and \U$15005 ( \15348 , \15347 , \14461 );
and \U$15006 ( \15349 , \14360 , \14456 );
or \U$15007 ( \15350 , \15348 , \15349 );
xor \U$15008 ( \15351 , \15346 , \15350 );
xor \U$15009 ( \15352 , \13257 , \14355 );
and \U$15010 ( \15353 , \15352 , \14462 );
and \U$15011 ( \15354 , \13257 , \14355 );
or \U$15012 ( \15355 , \15353 , \15354 );
nor \U$15013 ( \15356 , \15351 , \15355 );
not \U$15014 ( \15357 , \15356 );
xor \U$15015 ( \15358 , \14496 , \15223 );
xor \U$15016 ( \15359 , \15358 , \15226 );
xor \U$15017 ( \15360 , \14707 , \14709 );
xor \U$15018 ( \15361 , \15360 , \14991 );
not \U$15019 ( \15362 , \15361 );
xor \U$15020 ( \15363 , \14477 , \14479 );
xor \U$15021 ( \15364 , \15363 , \14482 );
xor \U$15022 ( \15365 , \14599 , \14701 );
xor \U$15023 ( \15366 , \15365 , \14704 );
xor \U$15024 ( \15367 , \15364 , \15366 );
xor \U$15025 ( \15368 , \14831 , \14879 );
xor \U$15026 ( \15369 , \15368 , \14874 );
not \U$15027 ( \15370 , \15369 );
not \U$15028 ( \15371 , \15370 );
xor \U$15029 ( \15372 , \14720 , \14731 );
xor \U$15030 ( \15373 , \15372 , \14742 );
not \U$15031 ( \15374 , \15373 );
xor \U$15032 ( \15375 , \14809 , \14825 );
xnor \U$15033 ( \15376 , \15375 , \14798 );
not \U$15034 ( \15377 , \15376 );
not \U$15035 ( \15378 , \15377 );
or \U$15036 ( \15379 , \15374 , \15378 );
not \U$15037 ( \15380 , \15376 );
or \U$15038 ( \15381 , \15373 , \15380 );
xor \U$15039 ( \15382 , \14932 , \14941 );
xor \U$15040 ( \15383 , \15382 , \14952 );
nand \U$15041 ( \15384 , \15381 , \15383 );
nand \U$15042 ( \15385 , \15379 , \15384 );
not \U$15043 ( \15386 , \15385 );
or \U$15044 ( \15387 , \15371 , \15386 );
or \U$15045 ( \15388 , \15370 , \15385 );
xor \U$15046 ( \15389 , \14848 , \14859 );
xnor \U$15047 ( \15390 , \15389 , \14872 );
not \U$15048 ( \15391 , \15390 );
not \U$15049 ( \15392 , \15391 );
not \U$15050 ( \15393 , \14848 );
not \U$15051 ( \15394 , \15393 );
not \U$15052 ( \15395 , \2940 );
not \U$15053 ( \15396 , RIbb2e800_31);
not \U$15054 ( \15397 , \3140 );
not \U$15055 ( \15398 , \15397 );
not \U$15056 ( \15399 , \15398 );
or \U$15057 ( \15400 , \15396 , \15399 );
nand \U$15058 ( \15401 , \3139 , \9169 );
nand \U$15059 ( \15402 , \15400 , \15401 );
not \U$15060 ( \15403 , \15402 );
or \U$15061 ( \15404 , \15395 , \15403 );
nand \U$15062 ( \15405 , \14805 , \3613 );
nand \U$15063 ( \15406 , \15404 , \15405 );
not \U$15064 ( \15407 , \15406 );
or \U$15065 ( \15408 , \15394 , \15407 );
not \U$15066 ( \15409 , \14848 );
not \U$15067 ( \15410 , \15406 );
not \U$15068 ( \15411 , \15410 );
or \U$15069 ( \15412 , \15409 , \15411 );
not \U$15070 ( \15413 , \2922 );
not \U$15071 ( \15414 , RIbb2e8f0_29);
not \U$15072 ( \15415 , \6173 );
or \U$15073 ( \15416 , \15414 , \15415 );
nand \U$15074 ( \15417 , \13903 , \2911 );
nand \U$15075 ( \15418 , \15416 , \15417 );
not \U$15076 ( \15419 , \15418 );
or \U$15077 ( \15420 , \15413 , \15419 );
nand \U$15078 ( \15421 , \14794 , \2925 );
nand \U$15079 ( \15422 , \15420 , \15421 );
nand \U$15080 ( \15423 , \15412 , \15422 );
nand \U$15081 ( \15424 , \15408 , \15423 );
not \U$15082 ( \15425 , \15424 );
or \U$15083 ( \15426 , \15392 , \15425 );
or \U$15084 ( \15427 , \15424 , \15391 );
not \U$15085 ( \15428 , \10449 );
not \U$15086 ( \15429 , RIbb2e260_43);
not \U$15087 ( \15430 , \8862 );
or \U$15088 ( \15431 , \15429 , \15430 );
nand \U$15089 ( \15432 , \1137 , \8347 );
nand \U$15090 ( \15433 , \15431 , \15432 );
not \U$15091 ( \15434 , \15433 );
or \U$15092 ( \15435 , \15428 , \15434 );
nand \U$15093 ( \15436 , \14855 , \9099 );
nand \U$15094 ( \15437 , \15435 , \15436 );
not \U$15095 ( \15438 , \15437 );
not \U$15096 ( \15439 , \3445 );
not \U$15097 ( \15440 , RIbb2e9e0_27);
not \U$15098 ( \15441 , \4021 );
or \U$15099 ( \15442 , \15440 , \15441 );
not \U$15100 ( \15443 , \4020 );
not \U$15101 ( \15444 , \15443 );
nand \U$15102 ( \15445 , \15444 , \4598 );
nand \U$15103 ( \15446 , \15442 , \15445 );
not \U$15104 ( \15447 , \15446 );
or \U$15105 ( \15448 , \15439 , \15447 );
nand \U$15106 ( \15449 , \14870 , \3465 );
nand \U$15107 ( \15450 , \15448 , \15449 );
not \U$15108 ( \15451 , \15450 );
or \U$15109 ( \15452 , \15438 , \15451 );
or \U$15110 ( \15453 , \15450 , \15437 );
not \U$15111 ( \15454 , \1264 );
not \U$15112 ( \15455 , \1288 );
buf \U$15113 ( \15456 , \13978 );
not \U$15114 ( \15457 , \15456 );
or \U$15115 ( \15458 , \15455 , \15457 );
nand \U$15116 ( \15459 , \13977 , \1244 );
nand \U$15117 ( \15460 , \15458 , \15459 );
not \U$15118 ( \15461 , \15460 );
or \U$15119 ( \15462 , \15454 , \15461 );
nand \U$15120 ( \15463 , \15057 , \1294 );
nand \U$15121 ( \15464 , \15462 , \15463 );
not \U$15122 ( \15465 , \1376 );
not \U$15123 ( \15466 , \15041 );
or \U$15124 ( \15467 , \15465 , \15466 );
not \U$15125 ( \15468 , \1393 );
not \U$15126 ( \15469 , \15029 );
not \U$15127 ( \15470 , \15469 );
not \U$15128 ( \15471 , \15470 );
not \U$15129 ( \15472 , \15471 );
or \U$15130 ( \15473 , \15468 , \15472 );
buf \U$15131 ( \15474 , \15470 );
nand \U$15132 ( \15475 , \15474 , \13990 );
nand \U$15133 ( \15476 , \15473 , \15475 );
nand \U$15134 ( \15477 , \15476 , \1429 );
nand \U$15135 ( \15478 , \15467 , \15477 );
xor \U$15136 ( \15479 , \15464 , \15478 );
not \U$15137 ( \15480 , \1737 );
not \U$15138 ( \15481 , \15171 );
or \U$15139 ( \15482 , \15480 , \15481 );
not \U$15140 ( \15483 , RIbb2f340_7);
buf \U$15141 ( \15484 , \12323 );
not \U$15142 ( \15485 , \15484 );
or \U$15143 ( \15486 , \15483 , \15485 );
nand \U$15144 ( \15487 , \12933 , \2700 );
nand \U$15145 ( \15488 , \15486 , \15487 );
nand \U$15146 ( \15489 , \15488 , \1702 );
nand \U$15147 ( \15490 , \15482 , \15489 );
and \U$15148 ( \15491 , \15479 , \15490 );
and \U$15149 ( \15492 , \15464 , \15478 );
or \U$15150 ( \15493 , \15491 , \15492 );
nand \U$15151 ( \15494 , \15453 , \15493 );
nand \U$15152 ( \15495 , \15452 , \15494 );
nand \U$15153 ( \15496 , \15427 , \15495 );
nand \U$15154 ( \15497 , \15426 , \15496 );
nand \U$15155 ( \15498 , \15388 , \15497 );
nand \U$15156 ( \15499 , \15387 , \15498 );
not \U$15157 ( \15500 , \15499 );
xor \U$15158 ( \15501 , \14829 , \14881 );
xor \U$15159 ( \15502 , \15501 , \14964 );
not \U$15160 ( \15503 , \15502 );
or \U$15161 ( \15504 , \15500 , \15503 );
or \U$15162 ( \15505 , \15502 , \15499 );
not \U$15163 ( \15506 , \14688 );
not \U$15164 ( \15507 , \14677 );
not \U$15165 ( \15508 , \15507 );
or \U$15166 ( \15509 , \15506 , \15508 );
or \U$15167 ( \15510 , \15507 , \14688 );
nand \U$15168 ( \15511 , \15509 , \15510 );
not \U$15169 ( \15512 , \14665 );
and \U$15170 ( \15513 , \15511 , \15512 );
not \U$15171 ( \15514 , \15511 );
and \U$15172 ( \15515 , \15514 , \14665 );
nor \U$15173 ( \15516 , \15513 , \15515 );
not \U$15174 ( \15517 , \15516 );
not \U$15175 ( \15518 , \15517 );
not \U$15176 ( \15519 , \14588 );
not \U$15177 ( \15520 , \14574 );
or \U$15178 ( \15521 , \15519 , \15520 );
or \U$15179 ( \15522 , \14588 , \14574 );
nand \U$15180 ( \15523 , \15521 , \15522 );
and \U$15181 ( \15524 , \15523 , \14576 );
not \U$15182 ( \15525 , \15523 );
and \U$15183 ( \15526 , \15525 , \14571 );
nor \U$15184 ( \15527 , \15524 , \15526 );
not \U$15185 ( \15528 , \15527 );
not \U$15186 ( \15529 , \15528 );
or \U$15187 ( \15530 , \15518 , \15529 );
not \U$15188 ( \15531 , \15527 );
not \U$15189 ( \15532 , \15516 );
or \U$15190 ( \15533 , \15531 , \15532 );
not \U$15191 ( \15534 , \10599 );
not \U$15192 ( \15535 , RIbb2e170_45);
not \U$15193 ( \15536 , \3370 );
or \U$15194 ( \15537 , \15535 , \15536 );
nand \U$15195 ( \15538 , \1687 , \9094 );
nand \U$15196 ( \15539 , \15537 , \15538 );
not \U$15197 ( \15540 , \15539 );
or \U$15198 ( \15541 , \15534 , \15540 );
nand \U$15199 ( \15542 , \14823 , \10119 );
nand \U$15200 ( \15543 , \15541 , \15542 );
not \U$15201 ( \15544 , \3887 );
not \U$15202 ( \15545 , RIbb2e710_33);
not \U$15203 ( \15546 , \3517 );
or \U$15204 ( \15547 , \15545 , \15546 );
nand \U$15205 ( \15548 , \12096 , \4785 );
nand \U$15206 ( \15549 , \15547 , \15548 );
not \U$15207 ( \15550 , \15549 );
or \U$15208 ( \15551 , \15544 , \15550 );
nand \U$15209 ( \15552 , \14716 , \4075 );
nand \U$15210 ( \15553 , \15551 , \15552 );
xor \U$15211 ( \15554 , \15543 , \15553 );
not \U$15212 ( \15555 , \12774 );
not \U$15213 ( \15556 , \984 );
and \U$15214 ( \15557 , RIbb2dea0_51, \15556 );
not \U$15215 ( \15558 , RIbb2dea0_51);
and \U$15216 ( \15559 , \15558 , \986 );
or \U$15217 ( \15560 , \15557 , \15559 );
not \U$15218 ( \15561 , \15560 );
or \U$15219 ( \15562 , \15555 , \15561 );
buf \U$15220 ( \15563 , \14738 );
nand \U$15221 ( \15564 , \15563 , \12692 );
nand \U$15222 ( \15565 , \15562 , \15564 );
and \U$15223 ( \15566 , \15554 , \15565 );
and \U$15224 ( \15567 , \15543 , \15553 );
or \U$15225 ( \15568 , \15566 , \15567 );
nand \U$15226 ( \15569 , \15533 , \15568 );
nand \U$15227 ( \15570 , \15530 , \15569 );
buf \U$15228 ( \15571 , \15570 );
not \U$15229 ( \15572 , \15571 );
xor \U$15230 ( \15573 , \14919 , \14955 );
xor \U$15231 ( \15574 , \15573 , \14961 );
not \U$15232 ( \15575 , \15574 );
or \U$15233 ( \15576 , \15572 , \15575 );
or \U$15234 ( \15577 , \15574 , \15571 );
not \U$15235 ( \15578 , \8362 );
not \U$15236 ( \15579 , RIbb2e350_41);
not \U$15237 ( \15580 , \3290 );
or \U$15238 ( \15581 , \15579 , \15580 );
not \U$15239 ( \15582 , \1280 );
not \U$15240 ( \15583 , \15582 );
nand \U$15241 ( \15584 , \15583 , \8357 );
nand \U$15242 ( \15585 , \15581 , \15584 );
not \U$15243 ( \15586 , \15585 );
or \U$15244 ( \15587 , \15578 , \15586 );
nand \U$15245 ( \15588 , \14901 , \8354 );
nand \U$15246 ( \15589 , \15587 , \15588 );
not \U$15247 ( \15590 , \15589 );
not \U$15248 ( \15591 , \3383 );
not \U$15249 ( \15592 , \14948 );
or \U$15250 ( \15593 , \15591 , \15592 );
not \U$15251 ( \15594 , RIbb2ebc0_23);
not \U$15252 ( \15595 , \4325 );
or \U$15253 ( \15596 , \15594 , \15595 );
nand \U$15254 ( \15597 , \4085 , \3388 );
nand \U$15255 ( \15598 , \15596 , \15597 );
nand \U$15256 ( \15599 , \15598 , \3406 );
nand \U$15257 ( \15600 , \15593 , \15599 );
not \U$15258 ( \15601 , \15600 );
or \U$15259 ( \15602 , \15590 , \15601 );
or \U$15260 ( \15603 , \15600 , \15589 );
not \U$15261 ( \15604 , \2980 );
not \U$15262 ( \15605 , \3274 );
and \U$15263 ( \15606 , RIbb2ead0_25, \15605 );
not \U$15264 ( \15607 , RIbb2ead0_25);
and \U$15265 ( \15608 , \15607 , \3274 );
or \U$15266 ( \15609 , \15606 , \15608 );
not \U$15267 ( \15610 , \15609 );
or \U$15268 ( \15611 , \15604 , \15610 );
nand \U$15269 ( \15612 , \14914 , \2963 );
nand \U$15270 ( \15613 , \15611 , \15612 );
nand \U$15271 ( \15614 , \15603 , \15613 );
nand \U$15272 ( \15615 , \15602 , \15614 );
not \U$15273 ( \15616 , \15615 );
not \U$15274 ( \15617 , \4712 );
not \U$15275 ( \15618 , RIbb2e620_35);
not \U$15276 ( \15619 , \3563 );
or \U$15277 ( \15620 , \15618 , \15619 );
nand \U$15278 ( \15621 , \2114 , \6002 );
nand \U$15279 ( \15622 , \15620 , \15621 );
not \U$15280 ( \15623 , \15622 );
or \U$15281 ( \15624 , \15617 , \15623 );
nand \U$15282 ( \15625 , \14729 , \5845 );
nand \U$15283 ( \15626 , \15624 , \15625 );
not \U$15284 ( \15627 , \11176 );
not \U$15285 ( \15628 , RIbb2e080_47);
not \U$15286 ( \15629 , \1548 );
not \U$15287 ( \15630 , \15629 );
or \U$15288 ( \15631 , \15628 , \15630 );
not \U$15289 ( \15632 , RIbb2e080_47);
nand \U$15290 ( \15633 , \1548 , \15632 );
nand \U$15291 ( \15634 , \15631 , \15633 );
not \U$15292 ( \15635 , \15634 );
or \U$15293 ( \15636 , \15627 , \15635 );
nand \U$15294 ( \15637 , \14760 , \12965 );
nand \U$15295 ( \15638 , \15636 , \15637 );
or \U$15296 ( \15639 , \15626 , \15638 );
not \U$15297 ( \15640 , \6242 );
not \U$15298 ( \15641 , \14779 );
or \U$15299 ( \15642 , \15640 , \15641 );
not \U$15300 ( \15643 , RIbb2e530_37);
not \U$15301 ( \15644 , \6095 );
or \U$15302 ( \15645 , \15643 , \15644 );
nand \U$15303 ( \15646 , \3495 , \6246 );
nand \U$15304 ( \15647 , \15645 , \15646 );
nand \U$15305 ( \15648 , \15647 , \6251 );
nand \U$15306 ( \15649 , \15642 , \15648 );
nand \U$15307 ( \15650 , \15639 , \15649 );
nand \U$15308 ( \15651 , \15626 , \15638 );
nand \U$15309 ( \15652 , \15650 , \15651 );
not \U$15310 ( \15653 , \15652 );
or \U$15311 ( \15654 , \15616 , \15653 );
not \U$15312 ( \15655 , \15615 );
not \U$15313 ( \15656 , \15655 );
not \U$15314 ( \15657 , \15652 );
not \U$15315 ( \15658 , \15657 );
or \U$15316 ( \15659 , \15656 , \15658 );
not \U$15317 ( \15660 , \12167 );
not \U$15318 ( \15661 , RIbb2df90_49);
not \U$15319 ( \15662 , \1069 );
or \U$15320 ( \15663 , \15661 , \15662 );
nand \U$15321 ( \15664 , \13611 , \12278 );
nand \U$15322 ( \15665 , \15663 , \15664 );
not \U$15323 ( \15666 , \15665 );
or \U$15324 ( \15667 , \15660 , \15666 );
nand \U$15325 ( \15668 , \14749 , \12284 );
nand \U$15326 ( \15669 , \15667 , \15668 );
not \U$15327 ( \15670 , \7103 );
and \U$15328 ( \15671 , RIbb2e440_39, \4339 );
not \U$15329 ( \15672 , RIbb2e440_39);
and \U$15330 ( \15673 , \15672 , \1386 );
or \U$15331 ( \15674 , \15671 , \15673 );
not \U$15332 ( \15675 , \15674 );
or \U$15333 ( \15676 , \15670 , \15675 );
nand \U$15334 ( \15677 , \14939 , \8450 );
nand \U$15335 ( \15678 , \15676 , \15677 );
nor \U$15336 ( \15679 , \15669 , \15678 );
not \U$15337 ( \15680 , \14920 );
not \U$15338 ( \15681 , RIbb2ddb0_53);
not \U$15339 ( \15682 , \13307 );
or \U$15340 ( \15683 , \15681 , \15682 );
nand \U$15341 ( \15684 , \8755 , \13463 );
nand \U$15342 ( \15685 , \15683 , \15684 );
not \U$15343 ( \15686 , \15685 );
or \U$15344 ( \15687 , \15680 , \15686 );
not \U$15345 ( \15688 , \13937 );
nand \U$15346 ( \15689 , \14926 , \15688 );
nand \U$15347 ( \15690 , \15687 , \15689 );
not \U$15348 ( \15691 , \15690 );
or \U$15349 ( \15692 , \15679 , \15691 );
nand \U$15350 ( \15693 , \15669 , \15678 );
nand \U$15351 ( \15694 , \15692 , \15693 );
nand \U$15352 ( \15695 , \15659 , \15694 );
nand \U$15353 ( \15696 , \15654 , \15695 );
nand \U$15354 ( \15697 , \15577 , \15696 );
nand \U$15355 ( \15698 , \15576 , \15697 );
nand \U$15356 ( \15699 , \15505 , \15698 );
nand \U$15357 ( \15700 , \15504 , \15699 );
and \U$15358 ( \15701 , \15367 , \15700 );
and \U$15359 ( \15702 , \15364 , \15366 );
or \U$15360 ( \15703 , \15701 , \15702 );
not \U$15361 ( \15704 , \15703 );
nand \U$15362 ( \15705 , \15362 , \15704 );
not \U$15363 ( \15706 , \15705 );
xor \U$15364 ( \15707 , \14967 , \14985 );
xor \U$15365 ( \15708 , \15707 , \14988 );
xor \U$15366 ( \15709 , \14969 , \14971 );
xor \U$15367 ( \15710 , \15709 , \14982 );
xor \U$15368 ( \15711 , \14745 , \14827 );
xnor \U$15369 ( \15712 , \15711 , \14783 );
not \U$15370 ( \15713 , \15712 );
xor \U$15371 ( \15714 , \14976 , \14979 );
not \U$15372 ( \15715 , \14974 );
and \U$15373 ( \15716 , \15714 , \15715 );
not \U$15374 ( \15717 , \15714 );
and \U$15375 ( \15718 , \15717 , \14974 );
nor \U$15376 ( \15719 , \15716 , \15718 );
not \U$15377 ( \15720 , \15719 );
or \U$15378 ( \15721 , \15713 , \15720 );
xor \U$15379 ( \15722 , \14894 , \14905 );
xor \U$15380 ( \15723 , \15722 , \14916 );
not \U$15381 ( \15724 , \15723 );
not \U$15382 ( \15725 , \15724 );
not \U$15383 ( \15726 , \15725 );
not \U$15384 ( \15727 , \14764 );
not \U$15385 ( \15728 , \14767 );
or \U$15386 ( \15729 , \15727 , \15728 );
or \U$15387 ( \15730 , \14764 , \14767 );
nand \U$15388 ( \15731 , \15729 , \15730 );
xnor \U$15389 ( \15732 , \15731 , \14781 );
not \U$15390 ( \15733 , \15732 );
not \U$15391 ( \15734 , \15733 );
or \U$15392 ( \15735 , \15726 , \15734 );
or \U$15393 ( \15736 , \15733 , \15725 );
xor \U$15394 ( \15737 , RIbb2db58_58, RIbb2dae0_59);
buf \U$15395 ( \15738 , \15737 );
not \U$15396 ( \15739 , \15738 );
not \U$15397 ( \15740 , \15739 );
not \U$15398 ( \15741 , RIbb2dbd0_57);
and \U$15399 ( \15742 , RIbb2db58_58, \15741 );
not \U$15400 ( \15743 , RIbb2db58_58);
and \U$15401 ( \15744 , \15743 , RIbb2dbd0_57);
nor \U$15402 ( \15745 , \15742 , \15744 );
nor \U$15403 ( \15746 , \15745 , \15737 );
not \U$15404 ( \15747 , \15746 );
not \U$15405 ( \15748 , \15747 );
or \U$15406 ( \15749 , \15740 , \15748 );
nand \U$15407 ( \15750 , \15749 , RIbb2dbd0_57);
and \U$15408 ( \15751 , \457 , \15024 );
xor \U$15409 ( \15752 , \13194 , \15751 );
buf \U$15410 ( \15753 , \15752 );
not \U$15411 ( \15754 , \15753 );
buf \U$15412 ( \15755 , \15754 );
not \U$15413 ( \15756 , \15755 );
and \U$15414 ( \15757 , \15756 , \1393 );
xor \U$15415 ( \15758 , \15750 , \15757 );
not \U$15416 ( \15759 , \1089 );
not \U$15417 ( \15760 , RIbb2f430_5);
not \U$15418 ( \15761 , \13474 );
not \U$15419 ( \15762 , \15761 );
or \U$15420 ( \15763 , \15760 , \15762 );
nand \U$15421 ( \15764 , \14625 , \1980 );
nand \U$15422 ( \15765 , \15763 , \15764 );
not \U$15423 ( \15766 , \15765 );
or \U$15424 ( \15767 , \15759 , \15766 );
nand \U$15425 ( \15768 , \14846 , \1147 );
nand \U$15426 ( \15769 , \15767 , \15768 );
and \U$15427 ( \15770 , \15758 , \15769 );
and \U$15428 ( \15771 , \15750 , \15757 );
or \U$15429 ( \15772 , \15770 , \15771 );
not \U$15430 ( \15773 , \832 );
not \U$15431 ( \15774 , RIbb2ee90_17);
not \U$15432 ( \15775 , \13853 );
or \U$15433 ( \15776 , \15774 , \15775 );
nand \U$15434 ( \15777 , \14673 , \859 );
nand \U$15435 ( \15778 , \15776 , \15777 );
not \U$15436 ( \15779 , \15778 );
or \U$15437 ( \15780 , \15773 , \15779 );
nand \U$15438 ( \15781 , \15070 , \836 );
nand \U$15439 ( \15782 , \15780 , \15781 );
not \U$15440 ( \15783 , \1517 );
not \U$15441 ( \15784 , \15120 );
or \U$15442 ( \15785 , \15783 , \15784 );
not \U$15443 ( \15786 , \8630 );
and \U$15444 ( \15787 , RIbb2ef80_15, \15786 );
not \U$15445 ( \15788 , RIbb2ef80_15);
and \U$15446 ( \15789 , \15788 , \13866 );
or \U$15447 ( \15790 , \15787 , \15789 );
nand \U$15448 ( \15791 , \15790 , \1445 );
nand \U$15449 ( \15792 , \15785 , \15791 );
or \U$15450 ( \15793 , \15782 , \15792 );
not \U$15451 ( \15794 , \853 );
not \U$15452 ( \15795 , RIbb2eda0_19);
not \U$15453 ( \15796 , \8337 );
not \U$15454 ( \15797 , \15796 );
not \U$15455 ( \15798 , \15797 );
or \U$15456 ( \15799 , \15795 , \15798 );
nand \U$15457 ( \15800 , \13879 , \1776 );
nand \U$15458 ( \15801 , \15799 , \15800 );
not \U$15459 ( \15802 , \15801 );
or \U$15460 ( \15803 , \15794 , \15802 );
nand \U$15461 ( \15804 , \15095 , \855 );
nand \U$15462 ( \15805 , \15803 , \15804 );
nand \U$15463 ( \15806 , \15793 , \15805 );
nand \U$15464 ( \15807 , \15782 , \15792 );
nand \U$15465 ( \15808 , \15806 , \15807 );
xor \U$15466 ( \15809 , \15772 , \15808 );
and \U$15467 ( \15810 , \483 , \489 );
not \U$15468 ( \15811 , \15810 );
not \U$15469 ( \15812 , \12301 );
or \U$15470 ( \15813 , \15811 , \15812 );
and \U$15471 ( \15814 , \581 , \489 );
nor \U$15472 ( \15815 , \15814 , \585 );
nand \U$15473 ( \15816 , \15813 , \15815 );
nand \U$15474 ( \15817 , \486 , \587 );
not \U$15475 ( \15818 , \15817 );
and \U$15476 ( \15819 , \15816 , \15818 );
not \U$15477 ( \15820 , \15816 );
and \U$15478 ( \15821 , \15820 , \15817 );
nor \U$15479 ( \15822 , \15819 , \15821 );
not \U$15480 ( \15823 , \15822 );
buf \U$15481 ( \15824 , \15823 );
not \U$15482 ( \15825 , \15824 );
and \U$15483 ( \15826 , \15825 , \1393 );
not \U$15484 ( \15827 , \3383 );
not \U$15485 ( \15828 , \15598 );
or \U$15486 ( \15829 , \15827 , \15828 );
not \U$15487 ( \15830 , RIbb2ebc0_23);
not \U$15488 ( \15831 , \13560 );
or \U$15489 ( \15832 , \15830 , \15831 );
nand \U$15490 ( \15833 , \8375 , \3388 );
nand \U$15491 ( \15834 , \15832 , \15833 );
nand \U$15492 ( \15835 , \15834 , \3406 );
nand \U$15493 ( \15836 , \15829 , \15835 );
xor \U$15494 ( \15837 , \15826 , \15836 );
not \U$15495 ( \15838 , \2077 );
not \U$15496 ( \15839 , RIbb2ecb0_21);
not \U$15497 ( \15840 , \9109 );
or \U$15498 ( \15841 , \15839 , \15840 );
nand \U$15499 ( \15842 , \7111 , \849 );
nand \U$15500 ( \15843 , \15841 , \15842 );
not \U$15501 ( \15844 , \15843 );
or \U$15502 ( \15845 , \15838 , \15844 );
nand \U$15503 ( \15846 , \15080 , \2078 );
nand \U$15504 ( \15847 , \15845 , \15846 );
and \U$15505 ( \15848 , \15837 , \15847 );
and \U$15506 ( \15849 , \15826 , \15836 );
or \U$15507 ( \15850 , \15848 , \15849 );
and \U$15508 ( \15851 , \15809 , \15850 );
and \U$15509 ( \15852 , \15772 , \15808 );
or \U$15510 ( \15853 , \15851 , \15852 );
nand \U$15511 ( \15854 , \15736 , \15853 );
nand \U$15512 ( \15855 , \15735 , \15854 );
nand \U$15513 ( \15856 , \15721 , \15855 );
not \U$15514 ( \15857 , \15712 );
not \U$15515 ( \15858 , \15719 );
nand \U$15516 ( \15859 , \15857 , \15858 );
nand \U$15517 ( \15860 , \15856 , \15859 );
xor \U$15518 ( \15861 , \15710 , \15860 );
xor \U$15519 ( \15862 , \15012 , \15143 );
xor \U$15520 ( \15863 , \15862 , \15146 );
and \U$15521 ( \15864 , \15861 , \15863 );
and \U$15522 ( \15865 , \15710 , \15860 );
or \U$15523 ( \15866 , \15864 , \15865 );
xor \U$15524 ( \15867 , \15708 , \15866 );
xor \U$15525 ( \15868 , \15010 , \15149 );
xor \U$15526 ( \15869 , \15868 , \15211 );
and \U$15527 ( \15870 , \15867 , \15869 );
and \U$15528 ( \15871 , \15708 , \15866 );
or \U$15529 ( \15872 , \15870 , \15871 );
not \U$15530 ( \15873 , \15872 );
or \U$15531 ( \15874 , \15706 , \15873 );
not \U$15532 ( \15875 , \15362 );
nand \U$15533 ( \15876 , \15875 , \15703 );
nand \U$15534 ( \15877 , \15874 , \15876 );
xor \U$15535 ( \15878 , \14472 , \14474 );
xor \U$15536 ( \15879 , \15878 , \14493 );
buf \U$15537 ( \15880 , \15879 );
or \U$15538 ( \15881 , \15877 , \15880 );
xor \U$15539 ( \15882 , \14994 , \15005 );
xor \U$15540 ( \15883 , \15882 , \15220 );
nand \U$15541 ( \15884 , \15881 , \15883 );
nand \U$15542 ( \15885 , \15877 , \15880 );
nand \U$15543 ( \15886 , \15884 , \15885 );
or \U$15544 ( \15887 , \15359 , \15886 );
and \U$15545 ( \15888 , \15230 , \15357 , \15887 );
not \U$15546 ( \15889 , \15247 );
not \U$15547 ( \15890 , \15252 );
not \U$15548 ( \15891 , \15890 );
or \U$15549 ( \15892 , \15889 , \15891 );
or \U$15550 ( \15893 , \15890 , \15247 );
nand \U$15551 ( \15894 , \15893 , \15249 );
nand \U$15552 ( \15895 , \15892 , \15894 );
xor \U$15553 ( \15896 , \11331 , \11368 );
xor \U$15554 ( \15897 , \15896 , \11401 );
xor \U$15555 ( \15898 , \11085 , \11087 );
xor \U$15556 ( \15899 , \15898 , \11090 );
xor \U$15557 ( \15900 , \15897 , \15899 );
xor \U$15558 ( \15901 , \11105 , \11107 );
xor \U$15559 ( \15902 , \15901 , \11113 );
xor \U$15560 ( \15903 , \15900 , \15902 );
xor \U$15561 ( \15904 , \15895 , \15903 );
xor \U$15562 ( \15905 , \15267 , \15271 );
and \U$15563 ( \15906 , \15905 , \15276 );
and \U$15564 ( \15907 , \15267 , \15271 );
or \U$15565 ( \15908 , \15906 , \15907 );
xnor \U$15566 ( \15909 , \15904 , \15908 );
not \U$15567 ( \15910 , \15909 );
xor \U$15568 ( \15911 , \15245 , \15253 );
and \U$15569 ( \15912 , \15911 , \15277 );
and \U$15570 ( \15913 , \15245 , \15253 );
or \U$15571 ( \15914 , \15912 , \15913 );
not \U$15572 ( \15915 , \15914 );
or \U$15573 ( \15916 , \15910 , \15915 );
or \U$15574 ( \15917 , \15914 , \15909 );
nand \U$15575 ( \15918 , \15916 , \15917 );
xor \U$15576 ( \15919 , \15283 , \15289 );
and \U$15577 ( \15920 , \15919 , \15343 );
and \U$15578 ( \15921 , \15283 , \15289 );
or \U$15579 ( \15922 , \15920 , \15921 );
not \U$15580 ( \15923 , \15922 );
and \U$15581 ( \15924 , \15918 , \15923 );
not \U$15582 ( \15925 , \15918 );
and \U$15583 ( \15926 , \15925 , \15922 );
or \U$15584 ( \15927 , \15924 , \15926 );
not \U$15585 ( \15928 , \15927 );
not \U$15586 ( \15929 , \15339 );
not \U$15587 ( \15930 , \15315 );
or \U$15588 ( \15931 , \15929 , \15930 );
not \U$15589 ( \15932 , \15318 );
not \U$15590 ( \15933 , \15338 );
or \U$15591 ( \15934 , \15932 , \15933 );
nand \U$15592 ( \15935 , \15934 , \15306 );
nand \U$15593 ( \15936 , \15931 , \15935 );
xor \U$15594 ( \15937 , \15298 , \15302 );
and \U$15595 ( \15938 , \15937 , \15305 );
and \U$15596 ( \15939 , \15298 , \15302 );
or \U$15597 ( \15940 , \15938 , \15939 );
not \U$15598 ( \15941 , \15940 );
not \U$15599 ( \15942 , \15941 );
not \U$15600 ( \15943 , \11497 );
not \U$15601 ( \15944 , \11563 );
not \U$15602 ( \15945 , \11489 );
or \U$15603 ( \15946 , \15944 , \15945 );
or \U$15604 ( \15947 , \11563 , \11489 );
nand \U$15605 ( \15948 , \15946 , \15947 );
not \U$15606 ( \15949 , \15948 );
and \U$15607 ( \15950 , \15943 , \15949 );
and \U$15608 ( \15951 , \15948 , \11497 );
nor \U$15609 ( \15952 , \15950 , \15951 );
not \U$15610 ( \15953 , \15952 );
not \U$15611 ( \15954 , \15953 );
xor \U$15612 ( \15955 , \15258 , \15260 );
and \U$15613 ( \15956 , \15955 , \15266 );
and \U$15614 ( \15957 , \15258 , \15260 );
or \U$15615 ( \15958 , \15956 , \15957 );
not \U$15616 ( \15959 , \15958 );
not \U$15617 ( \15960 , \15959 );
or \U$15618 ( \15961 , \15954 , \15960 );
nand \U$15619 ( \15962 , \15958 , \15952 );
nand \U$15620 ( \15963 , \15961 , \15962 );
not \U$15621 ( \15964 , \15963 );
or \U$15622 ( \15965 , \15942 , \15964 );
or \U$15623 ( \15966 , \15963 , \15941 );
nand \U$15624 ( \15967 , \15965 , \15966 );
xor \U$15625 ( \15968 , \15936 , \15967 );
xor \U$15626 ( \15969 , \11643 , \11685 );
xor \U$15627 ( \15970 , \15969 , \11789 );
not \U$15628 ( \15971 , \15337 );
not \U$15629 ( \15972 , \15326 );
or \U$15630 ( \15973 , \15971 , \15972 );
or \U$15631 ( \15974 , \15326 , \15337 );
nand \U$15632 ( \15975 , \15974 , \15330 );
nand \U$15633 ( \15976 , \15973 , \15975 );
xor \U$15634 ( \15977 , \15970 , \15976 );
xor \U$15635 ( \15978 , \11847 , \11849 );
xor \U$15636 ( \15979 , \15978 , \11862 );
xor \U$15637 ( \15980 , \15977 , \15979 );
xnor \U$15638 ( \15981 , \15968 , \15980 );
not \U$15639 ( \15982 , \15981 );
not \U$15640 ( \15983 , \15982 );
or \U$15641 ( \15984 , \15928 , \15983 );
not \U$15642 ( \15985 , \15981 );
and \U$15643 ( \15986 , \15918 , \15923 );
not \U$15644 ( \15987 , \15918 );
and \U$15645 ( \15988 , \15987 , \15922 );
nor \U$15646 ( \15989 , \15986 , \15988 );
not \U$15647 ( \15990 , \15989 );
or \U$15648 ( \15991 , \15985 , \15990 );
xor \U$15649 ( \15992 , \15238 , \15278 );
and \U$15650 ( \15993 , \15992 , \15344 );
and \U$15651 ( \15994 , \15238 , \15278 );
or \U$15652 ( \15995 , \15993 , \15994 );
nand \U$15653 ( \15996 , \15991 , \15995 );
nand \U$15654 ( \15997 , \15984 , \15996 );
xor \U$15655 ( \15998 , \11483 , \11565 );
xor \U$15656 ( \15999 , \15998 , \11792 );
xor \U$15657 ( \16000 , \15970 , \15976 );
and \U$15658 ( \16001 , \16000 , \15979 );
and \U$15659 ( \16002 , \15970 , \15976 );
or \U$15660 ( \16003 , \16001 , \16002 );
xor \U$15661 ( \16004 , \15999 , \16003 );
xor \U$15662 ( \16005 , \11806 , \11865 );
xor \U$15663 ( \16006 , \16005 , \11876 );
xor \U$15664 ( \16007 , \16004 , \16006 );
not \U$15665 ( \16008 , \15895 );
not \U$15666 ( \16009 , \16008 );
not \U$15667 ( \16010 , \15903 );
not \U$15668 ( \16011 , \16010 );
or \U$15669 ( \16012 , \16009 , \16011 );
nand \U$15670 ( \16013 , \16012 , \15908 );
not \U$15671 ( \16014 , \16008 );
nand \U$15672 ( \16015 , \16014 , \15903 );
nand \U$15673 ( \16016 , \16013 , \16015 );
xor \U$15674 ( \16017 , \15897 , \15899 );
and \U$15675 ( \16018 , \16017 , \15902 );
and \U$15676 ( \16019 , \15897 , \15899 );
or \U$15677 ( \16020 , \16018 , \16019 );
not \U$15678 ( \16021 , \15953 );
not \U$15679 ( \16022 , \15958 );
or \U$15680 ( \16023 , \16021 , \16022 );
not \U$15681 ( \16024 , \15952 );
not \U$15682 ( \16025 , \15959 );
or \U$15683 ( \16026 , \16024 , \16025 );
nand \U$15684 ( \16027 , \16026 , \15940 );
nand \U$15685 ( \16028 , \16023 , \16027 );
xor \U$15686 ( \16029 , \16020 , \16028 );
not \U$15687 ( \16030 , \11033 );
not \U$15688 ( \16031 , \16030 );
not \U$15689 ( \16032 , \11028 );
or \U$15690 ( \16033 , \16031 , \16032 );
not \U$15691 ( \16034 , \11028 );
nand \U$15692 ( \16035 , \16034 , \11033 );
nand \U$15693 ( \16036 , \16033 , \16035 );
and \U$15694 ( \16037 , \16036 , \11036 );
not \U$15695 ( \16038 , \16036 );
not \U$15696 ( \16039 , \11036 );
and \U$15697 ( \16040 , \16038 , \16039 );
nor \U$15698 ( \16041 , \16037 , \16040 );
xor \U$15699 ( \16042 , \16029 , \16041 );
xor \U$15700 ( \16043 , \16016 , \16042 );
or \U$15701 ( \16044 , \15936 , \15967 );
nand \U$15702 ( \16045 , \16044 , \15980 );
nand \U$15703 ( \16046 , \15936 , \15967 );
nand \U$15704 ( \16047 , \16045 , \16046 );
xor \U$15705 ( \16048 , \16043 , \16047 );
xor \U$15706 ( \16049 , \16007 , \16048 );
not \U$15707 ( \16050 , \15914 );
not \U$15708 ( \16051 , \15909 );
not \U$15709 ( \16052 , \16051 );
or \U$15710 ( \16053 , \16050 , \16052 );
not \U$15711 ( \16054 , \15909 );
not \U$15712 ( \16055 , \15914 );
not \U$15713 ( \16056 , \16055 );
or \U$15714 ( \16057 , \16054 , \16056 );
nand \U$15715 ( \16058 , \16057 , \15922 );
nand \U$15716 ( \16059 , \16053 , \16058 );
xor \U$15717 ( \16060 , \16049 , \16059 );
or \U$15718 ( \16061 , \15997 , \16060 );
xor \U$15719 ( \16062 , \11795 , \11879 );
xnor \U$15720 ( \16063 , \16062 , \11801 );
xor \U$15721 ( \16064 , \16016 , \16042 );
and \U$15722 ( \16065 , \16064 , \16047 );
and \U$15723 ( \16066 , \16016 , \16042 );
or \U$15724 ( \16067 , \16065 , \16066 );
not \U$15725 ( \16068 , \16067 );
xor \U$15726 ( \16069 , \16063 , \16068 );
not \U$15727 ( \16070 , \11450 );
not \U$15728 ( \16071 , \11459 );
or \U$15729 ( \16072 , \16070 , \16071 );
or \U$15730 ( \16073 , \11459 , \11450 );
nand \U$15731 ( \16074 , \16072 , \16073 );
not \U$15732 ( \16075 , \11463 );
and \U$15733 ( \16076 , \16074 , \16075 );
not \U$15734 ( \16077 , \16074 );
and \U$15735 ( \16078 , \16077 , \11463 );
nor \U$15736 ( \16079 , \16076 , \16078 );
xor \U$15737 ( \16080 , \16020 , \16028 );
and \U$15738 ( \16081 , \16080 , \16041 );
and \U$15739 ( \16082 , \16020 , \16028 );
or \U$15740 ( \16083 , \16081 , \16082 );
xor \U$15741 ( \16084 , \16079 , \16083 );
xor \U$15742 ( \16085 , \15999 , \16003 );
and \U$15743 ( \16086 , \16085 , \16006 );
and \U$15744 ( \16087 , \15999 , \16003 );
or \U$15745 ( \16088 , \16086 , \16087 );
xor \U$15746 ( \16089 , \16084 , \16088 );
xor \U$15747 ( \16090 , \16069 , \16089 );
xor \U$15748 ( \16091 , \16007 , \16048 );
and \U$15749 ( \16092 , \16091 , \16059 );
and \U$15750 ( \16093 , \16007 , \16048 );
or \U$15751 ( \16094 , \16092 , \16093 );
not \U$15752 ( \16095 , \16094 );
nand \U$15753 ( \16096 , \16090 , \16095 );
xor \U$15754 ( \16097 , \11120 , \11410 );
xor \U$15755 ( \16098 , \16097 , \11413 );
xor \U$15756 ( \16099 , \11883 , \11479 );
xor \U$15757 ( \16100 , \16099 , \11881 );
xor \U$15758 ( \16101 , \16098 , \16100 );
not \U$15759 ( \16102 , \16079 );
not \U$15760 ( \16103 , \16102 );
not \U$15761 ( \16104 , \16088 );
or \U$15762 ( \16105 , \16103 , \16104 );
or \U$15763 ( \16106 , \16088 , \16102 );
nand \U$15764 ( \16107 , \16106 , \16083 );
nand \U$15765 ( \16108 , \16105 , \16107 );
xor \U$15766 ( \16109 , \16101 , \16108 );
xor \U$15767 ( \16110 , \16063 , \16068 );
and \U$15768 ( \16111 , \16110 , \16089 );
and \U$15769 ( \16112 , \16063 , \16068 );
or \U$15770 ( \16113 , \16111 , \16112 );
nand \U$15771 ( \16114 , \16109 , \16113 );
not \U$15772 ( \16115 , \16098 );
not \U$15773 ( \16116 , \16100 );
not \U$15774 ( \16117 , \16116 );
or \U$15775 ( \16118 , \16115 , \16117 );
not \U$15776 ( \16119 , \16098 );
nand \U$15777 ( \16120 , \16119 , \16100 );
nand \U$15778 ( \16121 , \16108 , \16120 );
nand \U$15779 ( \16122 , \16118 , \16121 );
not \U$15780 ( \16123 , \16122 );
xor \U$15781 ( \16124 , \11439 , \11886 );
xnor \U$15782 ( \16125 , \16124 , \11437 );
nand \U$15783 ( \16126 , \16123 , \16125 );
and \U$15784 ( \16127 , \16061 , \16096 , \16114 , \16126 );
xor \U$15785 ( \16128 , \15234 , \15345 );
and \U$15786 ( \16129 , \16128 , \15350 );
and \U$15787 ( \16130 , \15234 , \15345 );
or \U$15788 ( \16131 , \16129 , \16130 );
not \U$15789 ( \16132 , \16131 );
not \U$15790 ( \16133 , \15927 );
not \U$15791 ( \16134 , \15981 );
or \U$15792 ( \16135 , \16133 , \16134 );
nand \U$15793 ( \16136 , \15989 , \15982 );
nand \U$15794 ( \16137 , \16135 , \16136 );
xnor \U$15795 ( \16138 , \16137 , \15995 );
nand \U$15796 ( \16139 , \16132 , \16138 );
and \U$15797 ( \16140 , \11947 , \15888 , \16127 , \16139 );
not \U$15798 ( \16141 , \16140 );
not \U$15799 ( \16142 , \2925 );
not \U$15800 ( \16143 , RIbb2e8f0_29);
not \U$15801 ( \16144 , \4752 );
or \U$15802 ( \16145 , \16143 , \16144 );
nand \U$15803 ( \16146 , \10458 , \3440 );
nand \U$15804 ( \16147 , \16145 , \16146 );
not \U$15805 ( \16148 , \16147 );
or \U$15806 ( \16149 , \16142 , \16148 );
not \U$15807 ( \16150 , RIbb2e8f0_29);
not \U$15808 ( \16151 , \13756 );
or \U$15809 ( \16152 , \16150 , \16151 );
buf \U$15810 ( \16153 , \13551 );
nand \U$15811 ( \16154 , \16153 , \2911 );
nand \U$15812 ( \16155 , \16152 , \16154 );
nand \U$15813 ( \16156 , \16155 , \2922 );
nand \U$15814 ( \16157 , \16149 , \16156 );
not \U$15815 ( \16158 , \16157 );
not \U$15816 ( \16159 , \11176 );
not \U$15817 ( \16160 , RIbb2e080_47);
not \U$15818 ( \16161 , \3290 );
or \U$15819 ( \16162 , \16160 , \16161 );
not \U$15820 ( \16163 , RIbb2e080_47);
nand \U$15821 ( \16164 , \1282 , \16163 );
nand \U$15822 ( \16165 , \16162 , \16164 );
not \U$15823 ( \16166 , \16165 );
or \U$15824 ( \16167 , \16159 , \16166 );
not \U$15825 ( \16168 , RIbb2e080_47);
not \U$15826 ( \16169 , \3066 );
or \U$15827 ( \16170 , \16168 , \16169 );
not \U$15828 ( \16171 , RIbb2e080_47);
nand \U$15829 ( \16172 , \4006 , \16171 );
nand \U$15830 ( \16173 , \16170 , \16172 );
nand \U$15831 ( \16174 , \16173 , \11177 );
nand \U$15832 ( \16175 , \16167 , \16174 );
not \U$15833 ( \16176 , \16175 );
or \U$15834 ( \16177 , \16158 , \16176 );
or \U$15835 ( \16178 , \16175 , \16157 );
not \U$15836 ( \16179 , \3613 );
not \U$15837 ( \16180 , \4028 );
not \U$15838 ( \16181 , \16180 );
not \U$15839 ( \16182 , \2917 );
and \U$15840 ( \16183 , \16181 , \16182 );
not \U$15841 ( \16184 , \3044 );
not \U$15842 ( \16185 , \16184 );
and \U$15843 ( \16186 , \16185 , \8810 );
nor \U$15844 ( \16187 , \16183 , \16186 );
nor \U$15845 ( \16188 , \16179 , \16187 );
not \U$15846 ( \16189 , \2940 );
nand \U$15847 ( \16190 , \15605 , RIbb2e800_31);
nand \U$15848 ( \16191 , \13732 , \9169 );
and \U$15849 ( \16192 , \16190 , \16191 );
nor \U$15850 ( \16193 , \16189 , \16192 );
nor \U$15851 ( \16194 , \16188 , \16193 );
not \U$15852 ( \16195 , \16194 );
nand \U$15853 ( \16196 , \16178 , \16195 );
nand \U$15854 ( \16197 , \16177 , \16196 );
not \U$15855 ( \16198 , \14920 );
not \U$15856 ( \16199 , RIbb2ddb0_53);
not \U$15857 ( \16200 , \5003 );
or \U$15858 ( \16201 , \16199 , \16200 );
nand \U$15859 ( \16202 , \1548 , \12681 );
nand \U$15860 ( \16203 , \16201 , \16202 );
not \U$15861 ( \16204 , \16203 );
or \U$15862 ( \16205 , \16198 , \16204 );
not \U$15863 ( \16206 , RIbb2ddb0_53);
not \U$15864 ( \16207 , \1036 );
not \U$15865 ( \16208 , \16207 );
or \U$15866 ( \16209 , \16206 , \16208 );
not \U$15867 ( \16210 , RIbb2ddb0_53);
nand \U$15868 ( \16211 , \1560 , \16210 );
nand \U$15869 ( \16212 , \16209 , \16211 );
nand \U$15870 ( \16213 , \16212 , \14930 );
nand \U$15871 ( \16214 , \16205 , \16213 );
not \U$15872 ( \16215 , \10451 );
not \U$15873 ( \16216 , RIbb2e260_43);
not \U$15874 ( \16217 , \3822 );
or \U$15875 ( \16218 , \16216 , \16217 );
nand \U$15876 ( \16219 , \3821 , \8347 );
nand \U$15877 ( \16220 , \16218 , \16219 );
not \U$15878 ( \16221 , \16220 );
or \U$15879 ( \16222 , \16215 , \16221 );
not \U$15880 ( \16223 , RIbb2e260_43);
not \U$15881 ( \16224 , \6095 );
or \U$15882 ( \16225 , \16223 , \16224 );
nand \U$15883 ( \16226 , \1338 , \8347 );
nand \U$15884 ( \16227 , \16225 , \16226 );
nand \U$15885 ( \16228 , \16227 , \9098 );
nand \U$15886 ( \16229 , \16222 , \16228 );
xor \U$15887 ( \16230 , \16214 , \16229 );
not \U$15888 ( \16231 , \8362 );
not \U$15889 ( \16232 , RIbb2e350_41);
not \U$15890 ( \16233 , \4449 );
or \U$15891 ( \16234 , \16232 , \16233 );
not \U$15892 ( \16235 , \3563 );
nand \U$15893 ( \16236 , \16235 , \9402 );
nand \U$15894 ( \16237 , \16234 , \16236 );
not \U$15895 ( \16238 , \16237 );
or \U$15896 ( \16239 , \16231 , \16238 );
not \U$15897 ( \16240 , RIbb2e350_41);
not \U$15898 ( \16241 , \4609 );
or \U$15899 ( \16242 , \16240 , \16241 );
nand \U$15900 ( \16243 , \4610 , \7097 );
nand \U$15901 ( \16244 , \16242 , \16243 );
nand \U$15902 ( \16245 , \16244 , \8995 );
nand \U$15903 ( \16246 , \16239 , \16245 );
and \U$15904 ( \16247 , \16230 , \16246 );
and \U$15905 ( \16248 , \16214 , \16229 );
or \U$15906 ( \16249 , \16247 , \16248 );
not \U$15907 ( \16250 , \16249 );
xor \U$15908 ( \16251 , \16197 , \16250 );
and \U$15909 ( \16252 , RIbb2da68_60, RIbb2d9f0_61);
not \U$15910 ( \16253 , RIbb2da68_60);
not \U$15911 ( \16254 , RIbb2d9f0_61);
and \U$15912 ( \16255 , \16253 , \16254 );
nor \U$15913 ( \16256 , \16252 , \16255 );
buf \U$15914 ( \16257 , \16256 );
not \U$15915 ( \16258 , \16257 );
and \U$15916 ( \16259 , RIbb2dae0_59, \1579 );
not \U$15917 ( \16260 , RIbb2dae0_59);
and \U$15918 ( \16261 , \16260 , \893 );
or \U$15919 ( \16262 , \16259 , \16261 );
not \U$15920 ( \16263 , \16262 );
or \U$15921 ( \16264 , \16258 , \16263 );
and \U$15922 ( \16265 , RIbb2dae0_59, \13307 );
not \U$15923 ( \16266 , RIbb2dae0_59);
and \U$15924 ( \16267 , \16266 , \1508 );
or \U$15925 ( \16268 , \16265 , \16267 );
xnor \U$15926 ( \16269 , RIbb2da68_60, RIbb2dae0_59);
nor \U$15927 ( \16270 , \16269 , \16256 );
buf \U$15928 ( \16271 , \16270 );
nand \U$15929 ( \16272 , \16268 , \16271 );
nand \U$15930 ( \16273 , \16264 , \16272 );
not \U$15931 ( \16274 , \14613 );
and \U$15932 ( \16275 , RIbb2dcc0_55, \1069 );
not \U$15933 ( \16276 , RIbb2dcc0_55);
not \U$15934 ( \16277 , \1069 );
and \U$15935 ( \16278 , \16276 , \16277 );
or \U$15936 ( \16279 , \16275 , \16278 );
not \U$15937 ( \16280 , \16279 );
or \U$15938 ( \16281 , \16274 , \16280 );
and \U$15939 ( \16282 , RIbb2dcc0_55, \10421 );
not \U$15940 ( \16283 , RIbb2dcc0_55);
and \U$15941 ( \16284 , \16283 , \956 );
or \U$15942 ( \16285 , \16282 , \16284 );
nand \U$15943 ( \16286 , \16285 , \15181 );
nand \U$15944 ( \16287 , \16281 , \16286 );
xor \U$15945 ( \16288 , \16273 , \16287 );
not \U$15946 ( \16289 , \10599 );
not \U$15947 ( \16290 , RIbb2e170_45);
not \U$15948 ( \16291 , \13619 );
or \U$15949 ( \16292 , \16290 , \16291 );
nand \U$15950 ( \16293 , \1386 , \12003 );
nand \U$15951 ( \16294 , \16292 , \16293 );
not \U$15952 ( \16295 , \16294 );
or \U$15953 ( \16296 , \16289 , \16295 );
not \U$15954 ( \16297 , RIbb2e170_45);
not \U$15955 ( \16298 , \1170 );
or \U$15956 ( \16299 , \16297 , \16298 );
nand \U$15957 ( \16300 , \12046 , \12451 );
nand \U$15958 ( \16301 , \16299 , \16300 );
nand \U$15959 ( \16302 , \16301 , \10119 );
nand \U$15960 ( \16303 , \16296 , \16302 );
and \U$15961 ( \16304 , \16288 , \16303 );
and \U$15962 ( \16305 , \16273 , \16287 );
or \U$15963 ( \16306 , \16304 , \16305 );
xnor \U$15964 ( \16307 , \16251 , \16306 );
not \U$15965 ( \16308 , \1702 );
not \U$15966 ( \16309 , \14526 );
and \U$15967 ( \16310 , \16309 , RIbb2f340_7);
not \U$15968 ( \16311 , \16309 );
and \U$15969 ( \16312 , \16311 , \1734 );
or \U$15970 ( \16313 , \16310 , \16312 );
not \U$15971 ( \16314 , \16313 );
or \U$15972 ( \16315 , \16308 , \16314 );
not \U$15973 ( \16316 , RIbb2f340_7);
not \U$15974 ( \16317 , \13976 );
not \U$15975 ( \16318 , \16317 );
or \U$15976 ( \16319 , \16316 , \16318 );
not \U$15977 ( \16320 , \16317 );
nand \U$15978 ( \16321 , \16320 , \1692 );
nand \U$15979 ( \16322 , \16319 , \16321 );
nand \U$15980 ( \16323 , \16322 , \1737 );
nand \U$15981 ( \16324 , \16315 , \16323 );
not \U$15982 ( \16325 , \3465 );
not \U$15983 ( \16326 , RIbb2e9e0_27);
not \U$15984 ( \16327 , \13560 );
or \U$15985 ( \16328 , \16326 , \16327 );
nand \U$15986 ( \16329 , \8375 , \3454 );
nand \U$15987 ( \16330 , \16328 , \16329 );
not \U$15988 ( \16331 , \16330 );
or \U$15989 ( \16332 , \16325 , \16331 );
not \U$15990 ( \16333 , \4598 );
not \U$15991 ( \16334 , \4697 );
or \U$15992 ( \16335 , \16333 , \16334 );
not \U$15993 ( \16336 , \6198 );
nand \U$15994 ( \16337 , \16336 , RIbb2e9e0_27);
nand \U$15995 ( \16338 , \16335 , \16337 );
nand \U$15996 ( \16339 , \16338 , \3445 );
nand \U$15997 ( \16340 , \16332 , \16339 );
xor \U$15998 ( \16341 , \16324 , \16340 );
and \U$15999 ( \16342 , RIbb2ead0_25, \14041 );
not \U$16000 ( \16343 , RIbb2ead0_25);
and \U$16001 ( \16344 , \16343 , \7308 );
or \U$16002 ( \16345 , \16342 , \16344 );
not \U$16003 ( \16346 , \16345 );
or \U$16004 ( \16347 , \16346 , \6131 );
and \U$16005 ( \16348 , RIbb2ead0_25, \10126 );
not \U$16006 ( \16349 , RIbb2ead0_25);
and \U$16007 ( \16350 , \16349 , \8387 );
or \U$16008 ( \16351 , \16348 , \16350 );
not \U$16009 ( \16352 , \16351 );
not \U$16010 ( \16353 , \2963 );
or \U$16011 ( \16354 , \16352 , \16353 );
nand \U$16012 ( \16355 , \16347 , \16354 );
xor \U$16013 ( \16356 , \16341 , \16355 );
not \U$16014 ( \16357 , \14613 );
and \U$16015 ( \16358 , RIbb2dcc0_55, \1559 );
not \U$16016 ( \16359 , RIbb2dcc0_55);
and \U$16017 ( \16360 , \16359 , \1037 );
or \U$16018 ( \16361 , \16358 , \16360 );
not \U$16019 ( \16362 , \16361 );
or \U$16020 ( \16363 , \16357 , \16362 );
nand \U$16021 ( \16364 , \16279 , \15181 );
nand \U$16022 ( \16365 , \16363 , \16364 );
not \U$16023 ( \16366 , \16365 );
not \U$16024 ( \16367 , \16366 );
not \U$16025 ( \16368 , \9098 );
not \U$16026 ( \16369 , RIbb2e260_43);
not \U$16027 ( \16370 , \4609 );
or \U$16028 ( \16371 , \16369 , \16370 );
nand \U$16029 ( \16372 , \1852 , \10444 );
nand \U$16030 ( \16373 , \16371 , \16372 );
not \U$16031 ( \16374 , \16373 );
or \U$16032 ( \16375 , \16368 , \16374 );
nand \U$16033 ( \16376 , \16227 , \9099 );
nand \U$16034 ( \16377 , \16375 , \16376 );
not \U$16035 ( \16378 , \16377 );
not \U$16036 ( \16379 , \16378 );
or \U$16037 ( \16380 , \16367 , \16379 );
not \U$16038 ( \16381 , \10119 );
not \U$16039 ( \16382 , \16294 );
or \U$16040 ( \16383 , \16381 , \16382 );
not \U$16041 ( \16384 , RIbb2e170_45);
not \U$16042 ( \16385 , \3822 );
or \U$16043 ( \16386 , \16384 , \16385 );
nand \U$16044 ( \16387 , \3821 , \12003 );
nand \U$16045 ( \16388 , \16386 , \16387 );
nand \U$16046 ( \16389 , \16388 , \10117 );
nand \U$16047 ( \16390 , \16383 , \16389 );
nand \U$16048 ( \16391 , \16380 , \16390 );
nand \U$16049 ( \16392 , \16377 , \16365 );
nand \U$16050 ( \16393 , \16391 , \16392 );
xor \U$16051 ( \16394 , \16356 , \16393 );
not \U$16052 ( \16395 , \5845 );
not \U$16053 ( \16396 , \3201 );
not \U$16054 ( \16397 , \6002 );
and \U$16055 ( \16398 , \16396 , \16397 );
not \U$16056 ( \16399 , \4637 );
not \U$16057 ( \16400 , \16399 );
and \U$16058 ( \16401 , \16400 , \6002 );
nor \U$16059 ( \16402 , \16398 , \16401 );
nor \U$16060 ( \16403 , \16395 , \16402 );
not \U$16061 ( \16404 , RIbb2e620_35);
not \U$16062 ( \16405 , \13836 );
or \U$16063 ( \16406 , \16404 , \16405 );
nand \U$16064 ( \16407 , \13903 , \6002 );
nand \U$16065 ( \16408 , \16406 , \16407 );
not \U$16066 ( \16409 , \16408 );
nor \U$16067 ( \16410 , \16409 , \4713 );
nor \U$16068 ( \16411 , \16403 , \16410 );
not \U$16069 ( \16412 , \16411 );
not \U$16070 ( \16413 , \13295 );
not \U$16071 ( \16414 , RIbb2df90_49);
not \U$16072 ( \16415 , \7424 );
or \U$16073 ( \16416 , \16414 , \16415 );
nand \U$16074 ( \16417 , \10673 , \12278 );
nand \U$16075 ( \16418 , \16416 , \16417 );
not \U$16076 ( \16419 , \16418 );
or \U$16077 ( \16420 , \16413 , \16419 );
not \U$16078 ( \16421 , \12278 );
not \U$16079 ( \16422 , \3243 );
or \U$16080 ( \16423 , \16421 , \16422 );
not \U$16081 ( \16424 , \1642 );
nand \U$16082 ( \16425 , \16424 , RIbb2df90_49);
nand \U$16083 ( \16426 , \16423 , \16425 );
buf \U$16084 ( \16427 , \12168 );
nand \U$16085 ( \16428 , \16426 , \16427 );
nand \U$16086 ( \16429 , \16420 , \16428 );
not \U$16087 ( \16430 , \16429 );
not \U$16088 ( \16431 , \6242 );
not \U$16089 ( \16432 , RIbb2e530_37);
not \U$16090 ( \16433 , \3952 );
or \U$16091 ( \16434 , \16432 , \16433 );
nand \U$16092 ( \16435 , \3951 , \4708 );
nand \U$16093 ( \16436 , \16434 , \16435 );
not \U$16094 ( \16437 , \16436 );
or \U$16095 ( \16438 , \16431 , \16437 );
not \U$16096 ( \16439 , RIbb2e530_37);
not \U$16097 ( \16440 , \6301 );
or \U$16098 ( \16441 , \16439 , \16440 );
nand \U$16099 ( \16442 , \15397 , \6246 );
nand \U$16100 ( \16443 , \16441 , \16442 );
nand \U$16101 ( \16444 , \16443 , \6251 );
nand \U$16102 ( \16445 , \16438 , \16444 );
not \U$16103 ( \16446 , \16445 );
not \U$16104 ( \16447 , \16446 );
or \U$16105 ( \16448 , \16430 , \16447 );
or \U$16106 ( \16449 , \16446 , \16429 );
nand \U$16107 ( \16450 , \16448 , \16449 );
xor \U$16108 ( \16451 , \16412 , \16450 );
and \U$16109 ( \16452 , \16394 , \16451 );
and \U$16110 ( \16453 , \16356 , \16393 );
or \U$16111 ( \16454 , \16452 , \16453 );
or \U$16112 ( \16455 , \16307 , \16454 );
not \U$16113 ( \16456 , \2078 );
not \U$16114 ( \16457 , RIbb2ecb0_21);
not \U$16115 ( \16458 , \9791 );
or \U$16116 ( \16459 , \16457 , \16458 );
nand \U$16117 ( \16460 , \11534 , \2067 );
nand \U$16118 ( \16461 , \16459 , \16460 );
not \U$16119 ( \16462 , \16461 );
or \U$16120 ( \16463 , \16456 , \16462 );
not \U$16121 ( \16464 , RIbb2ecb0_21);
not \U$16122 ( \16465 , \13853 );
or \U$16123 ( \16466 , \16464 , \16465 );
nand \U$16124 ( \16467 , \13854 , \2249 );
nand \U$16125 ( \16468 , \16466 , \16467 );
nand \U$16126 ( \16469 , \16468 , \2077 );
nand \U$16127 ( \16470 , \16463 , \16469 );
not \U$16128 ( \16471 , \836 );
not \U$16129 ( \16472 , RIbb2ee90_17);
not \U$16130 ( \16473 , \9279 );
or \U$16131 ( \16474 , \16472 , \16473 );
not \U$16132 ( \16475 , \13916 );
nand \U$16133 ( \16476 , \16475 , \859 );
nand \U$16134 ( \16477 , \16474 , \16476 );
not \U$16135 ( \16478 , \16477 );
or \U$16136 ( \16479 , \16471 , \16478 );
not \U$16137 ( \16480 , RIbb2ee90_17);
not \U$16138 ( \16481 , \12222 );
or \U$16139 ( \16482 , \16480 , \16481 );
nand \U$16140 ( \16483 , \9841 , \859 );
nand \U$16141 ( \16484 , \16482 , \16483 );
nand \U$16142 ( \16485 , \16484 , \832 );
nand \U$16143 ( \16486 , \16479 , \16485 );
and \U$16144 ( \16487 , \16470 , \16486 );
not \U$16145 ( \16488 , \16470 );
not \U$16146 ( \16489 , \16486 );
and \U$16147 ( \16490 , \16488 , \16489 );
nor \U$16148 ( \16491 , \16487 , \16490 );
not \U$16149 ( \16492 , \855 );
not \U$16150 ( \16493 , RIbb2eda0_19);
not \U$16151 ( \16494 , \8320 );
or \U$16152 ( \16495 , \16493 , \16494 );
nand \U$16153 ( \16496 , \9819 , \1776 );
nand \U$16154 ( \16497 , \16495 , \16496 );
not \U$16155 ( \16498 , \16497 );
or \U$16156 ( \16499 , \16492 , \16498 );
not \U$16157 ( \16500 , \1779 );
not \U$16158 ( \16501 , RIbb2eda0_19);
not \U$16159 ( \16502 , \13863 );
or \U$16160 ( \16503 , \16501 , \16502 );
nand \U$16161 ( \16504 , \13866 , \3251 );
nand \U$16162 ( \16505 , \16503 , \16504 );
nand \U$16163 ( \16506 , \16500 , \16505 );
nand \U$16164 ( \16507 , \16499 , \16506 );
not \U$16165 ( \16508 , \16507 );
and \U$16166 ( \16509 , \16491 , \16508 );
not \U$16167 ( \16510 , \16491 );
and \U$16168 ( \16511 , \16510 , \16507 );
nor \U$16169 ( \16512 , \16509 , \16511 );
not \U$16170 ( \16513 , \16512 );
not \U$16171 ( \16514 , \16513 );
not \U$16172 ( \16515 , \16445 );
not \U$16173 ( \16516 , \16412 );
or \U$16174 ( \16517 , \16515 , \16516 );
not \U$16175 ( \16518 , \16411 );
not \U$16176 ( \16519 , \16446 );
or \U$16177 ( \16520 , \16518 , \16519 );
nand \U$16178 ( \16521 , \16520 , \16429 );
nand \U$16179 ( \16522 , \16517 , \16521 );
not \U$16180 ( \16523 , \16522 );
not \U$16181 ( \16524 , \16523 );
or \U$16182 ( \16525 , \16514 , \16524 );
nand \U$16183 ( \16526 , \16522 , \16512 );
nand \U$16184 ( \16527 , \16525 , \16526 );
and \U$16185 ( \16528 , RIbb2d900_63, RIbb2d978_62);
not \U$16186 ( \16529 , RIbb2d900_63);
not \U$16187 ( \16530 , RIbb2d978_62);
and \U$16188 ( \16531 , \16529 , \16530 );
nor \U$16189 ( \16532 , \16528 , \16531 );
buf \U$16190 ( \16533 , \16532 );
not \U$16191 ( \16534 , \16533 );
not \U$16192 ( \16535 , \16534 );
and \U$16193 ( \16536 , \16530 , RIbb2d9f0_61);
not \U$16194 ( \16537 , RIbb2d9f0_61);
and \U$16195 ( \16538 , \16537 , RIbb2d978_62);
nor \U$16196 ( \16539 , \16536 , \16538 );
nor \U$16197 ( \16540 , \16539 , \16532 );
buf \U$16198 ( \16541 , \16540 );
not \U$16199 ( \16542 , \16541 );
not \U$16200 ( \16543 , \16542 );
or \U$16201 ( \16544 , \16535 , \16543 );
nand \U$16202 ( \16545 , \16544 , RIbb2d9f0_61);
not \U$16203 ( \16546 , \482 );
nand \U$16204 ( \16547 , \16546 , \577 );
not \U$16205 ( \16548 , \16547 );
not \U$16206 ( \16549 , \12301 );
or \U$16207 ( \16550 , \16548 , \16549 );
or \U$16208 ( \16551 , \16547 , \12301 );
nand \U$16209 ( \16552 , \16550 , \16551 );
buf \U$16210 ( \16553 , \16552 );
not \U$16211 ( \16554 , \16553 );
buf \U$16212 ( \16555 , \16554 );
not \U$16213 ( \16556 , \16555 );
and \U$16214 ( \16557 , \1312 , \16556 );
xor \U$16215 ( \16558 , \16545 , \16557 );
not \U$16216 ( \16559 , \1261 );
not \U$16217 ( \16560 , \1288 );
not \U$16218 ( \16561 , \15752 );
not \U$16219 ( \16562 , \16561 );
not \U$16220 ( \16563 , \16562 );
not \U$16221 ( \16564 , \16563 );
or \U$16222 ( \16565 , \16560 , \16564 );
buf \U$16223 ( \16566 , \15752 );
not \U$16224 ( \16567 , \16566 );
not \U$16225 ( \16568 , \16567 );
not \U$16226 ( \16569 , \1253 );
nand \U$16227 ( \16570 , \16568 , \16569 );
nand \U$16228 ( \16571 , \16565 , \16570 );
not \U$16229 ( \16572 , \16571 );
or \U$16230 ( \16573 , \16559 , \16572 );
not \U$16231 ( \16574 , \1288 );
buf \U$16232 ( \16575 , \15822 );
buf \U$16233 ( \16576 , \16575 );
not \U$16234 ( \16577 , \16576 );
not \U$16235 ( \16578 , \16577 );
or \U$16236 ( \16579 , \16574 , \16578 );
nand \U$16237 ( \16580 , \16576 , \16569 );
nand \U$16238 ( \16581 , \16579 , \16580 );
nand \U$16239 ( \16582 , \16581 , \1264 );
nand \U$16240 ( \16583 , \16573 , \16582 );
xor \U$16241 ( \16584 , \16558 , \16583 );
not \U$16242 ( \16585 , \1517 );
and \U$16243 ( \16586 , RIbb2ef80_15, \12230 );
not \U$16244 ( \16587 , RIbb2ef80_15);
and \U$16245 ( \16588 , \16587 , \10301 );
or \U$16246 ( \16589 , \16586 , \16588 );
not \U$16247 ( \16590 , \16589 );
or \U$16248 ( \16591 , \16585 , \16590 );
and \U$16249 ( \16592 , RIbb2ef80_15, \14563 );
not \U$16250 ( \16593 , RIbb2ef80_15);
and \U$16251 ( \16594 , \16593 , \10764 );
or \U$16252 ( \16595 , \16592 , \16594 );
nand \U$16253 ( \16596 , \16595 , \1445 );
nand \U$16254 ( \16597 , \16591 , \16596 );
xor \U$16255 ( \16598 , \16584 , \16597 );
not \U$16256 ( \16599 , \998 );
not \U$16257 ( \16600 , RIbb2f070_13);
not \U$16258 ( \16601 , \11144 );
not \U$16259 ( \16602 , \16601 );
or \U$16260 ( \16603 , \16600 , \16602 );
not \U$16261 ( \16604 , \15188 );
nand \U$16262 ( \16605 , \16604 , \3421 );
nand \U$16263 ( \16606 , \16603 , \16605 );
not \U$16264 ( \16607 , \16606 );
or \U$16265 ( \16608 , \16599 , \16607 );
not \U$16266 ( \16609 , RIbb2f070_13);
not \U$16267 ( \16610 , \11580 );
or \U$16268 ( \16611 , \16609 , \16610 );
nand \U$16269 ( \16612 , \14885 , \906 );
nand \U$16270 ( \16613 , \16611 , \16612 );
nand \U$16271 ( \16614 , \16613 , \916 );
nand \U$16272 ( \16615 , \16608 , \16614 );
xor \U$16273 ( \16616 , \16598 , \16615 );
not \U$16274 ( \16617 , \16616 );
and \U$16275 ( \16618 , \16527 , \16617 );
not \U$16276 ( \16619 , \16527 );
and \U$16277 ( \16620 , \16619 , \16616 );
nor \U$16278 ( \16621 , \16618 , \16620 );
not \U$16279 ( \16622 , \16621 );
nand \U$16280 ( \16623 , \16455 , \16622 );
nand \U$16281 ( \16624 , \16307 , \16454 );
nand \U$16282 ( \16625 , \16623 , \16624 );
not \U$16283 ( \16626 , \12692 );
and \U$16284 ( \16627 , RIbb2dea0_51, \3479 );
not \U$16285 ( \16628 , RIbb2dea0_51);
and \U$16286 ( \16629 , \16628 , \1730 );
or \U$16287 ( \16630 , \16627 , \16629 );
not \U$16288 ( \16631 , \16630 );
or \U$16289 ( \16632 , \16626 , \16631 );
not \U$16290 ( \16633 , \3363 );
and \U$16291 ( \16634 , RIbb2dea0_51, \16633 );
not \U$16292 ( \16635 , RIbb2dea0_51);
and \U$16293 ( \16636 , \16635 , \3369 );
or \U$16294 ( \16637 , \16634 , \16636 );
nand \U$16295 ( \16638 , \16637 , \12774 );
nand \U$16296 ( \16639 , \16632 , \16638 );
not \U$16297 ( \16640 , \16639 );
not \U$16298 ( \16641 , \8450 );
and \U$16299 ( \16642 , RIbb2e440_39, \13289 );
not \U$16300 ( \16643 , RIbb2e440_39);
and \U$16301 ( \16644 , \16643 , \13290 );
or \U$16302 ( \16645 , \16642 , \16644 );
not \U$16303 ( \16646 , \16645 );
or \U$16304 ( \16647 , \16641 , \16646 );
and \U$16305 ( \16648 , RIbb2e440_39, \12097 );
not \U$16306 ( \16649 , RIbb2e440_39);
and \U$16307 ( \16650 , \16649 , \12096 );
or \U$16308 ( \16651 , \16648 , \16650 );
nand \U$16309 ( \16652 , \16651 , \7103 );
nand \U$16310 ( \16653 , \16647 , \16652 );
not \U$16311 ( \16654 , \16653 );
not \U$16312 ( \16655 , \16654 );
or \U$16313 ( \16656 , \16640 , \16655 );
not \U$16314 ( \16657 , \16639 );
nand \U$16315 ( \16658 , \16657 , \16653 );
nand \U$16316 ( \16659 , \16656 , \16658 );
not \U$16317 ( \16660 , \15738 );
not \U$16318 ( \16661 , RIbb2dbd0_57);
not \U$16319 ( \16662 , \3451 );
or \U$16320 ( \16663 , \16661 , \16662 );
nand \U$16321 ( \16664 , \3450 , \14602 );
nand \U$16322 ( \16665 , \16663 , \16664 );
not \U$16323 ( \16666 , \16665 );
or \U$16324 ( \16667 , \16660 , \16666 );
not \U$16325 ( \16668 , RIbb2dbd0_57);
not \U$16326 ( \16669 , \988 );
or \U$16327 ( \16670 , \16668 , \16669 );
not \U$16328 ( \16671 , RIbb2dbd0_57);
nand \U$16329 ( \16672 , \987 , \16671 );
nand \U$16330 ( \16673 , \16670 , \16672 );
not \U$16331 ( \16674 , \15747 );
buf \U$16332 ( \16675 , \16674 );
nand \U$16333 ( \16676 , \16673 , \16675 );
nand \U$16334 ( \16677 , \16667 , \16676 );
not \U$16335 ( \16678 , \16677 );
and \U$16336 ( \16679 , \16659 , \16678 );
not \U$16337 ( \16680 , \16659 );
and \U$16338 ( \16681 , \16680 , \16677 );
nor \U$16339 ( \16682 , \16679 , \16681 );
not \U$16340 ( \16683 , \16682 );
xor \U$16341 ( \16684 , \16214 , \16229 );
xor \U$16342 ( \16685 , \16684 , \16246 );
not \U$16343 ( \16686 , \16685 );
not \U$16344 ( \16687 , \16686 );
or \U$16345 ( \16688 , \16683 , \16687 );
not \U$16346 ( \16689 , \461 );
not \U$16347 ( \16690 , \16689 );
buf \U$16348 ( \16691 , \468 );
not \U$16349 ( \16692 , \16691 );
or \U$16350 ( \16693 , \16690 , \16692 );
buf \U$16351 ( \16694 , \472 );
nand \U$16352 ( \16695 , \16693 , \16694 );
not \U$16353 ( \16696 , \460 );
and \U$16354 ( \16697 , \16696 , \475 );
and \U$16355 ( \16698 , \16695 , \16697 );
not \U$16356 ( \16699 , \16695 );
not \U$16357 ( \16700 , \16697 );
and \U$16358 ( \16701 , \16699 , \16700 );
nor \U$16359 ( \16702 , \16698 , \16701 );
buf \U$16360 ( \16703 , \16702 );
buf \U$16361 ( \16704 , \16703 );
and \U$16362 ( \16705 , \1393 , \16704 );
buf \U$16363 ( \16706 , \16553 );
not \U$16364 ( \16707 , \16706 );
not \U$16365 ( \16708 , \13990 );
or \U$16366 ( \16709 , \16707 , \16708 );
not \U$16367 ( \16710 , \16553 );
nand \U$16368 ( \16711 , \1312 , \16710 );
nand \U$16369 ( \16712 , \16709 , \16711 );
not \U$16370 ( \16713 , \16712 );
not \U$16371 ( \16714 , \1428 );
or \U$16372 ( \16715 , \16713 , \16714 );
not \U$16373 ( \16716 , \16546 );
not \U$16374 ( \16717 , \12301 );
or \U$16375 ( \16718 , \16716 , \16717 );
nand \U$16376 ( \16719 , \16718 , \577 );
not \U$16377 ( \16720 , \580 );
nor \U$16378 ( \16721 , \16720 , \578 );
and \U$16379 ( \16722 , \16719 , \16721 );
not \U$16380 ( \16723 , \16719 );
not \U$16381 ( \16724 , \16721 );
and \U$16382 ( \16725 , \16723 , \16724 );
nor \U$16383 ( \16726 , \16722 , \16725 );
not \U$16384 ( \16727 , \16726 );
buf \U$16385 ( \16728 , \16727 );
not \U$16386 ( \16729 , \16728 );
xor \U$16387 ( \16730 , \1312 , \16729 );
nand \U$16388 ( \16731 , \16730 , \1375 );
nand \U$16389 ( \16732 , \16715 , \16731 );
xor \U$16390 ( \16733 , \16705 , \16732 );
not \U$16391 ( \16734 , \1288 );
not \U$16392 ( \16735 , \483 );
not \U$16393 ( \16736 , \12301 );
or \U$16394 ( \16737 , \16735 , \16736 );
not \U$16395 ( \16738 , \581 );
nand \U$16396 ( \16739 , \16737 , \16738 );
nand \U$16397 ( \16740 , \489 , \584 );
not \U$16398 ( \16741 , \16740 );
and \U$16399 ( \16742 , \16739 , \16741 );
not \U$16400 ( \16743 , \16739 );
and \U$16401 ( \16744 , \16743 , \16740 );
nor \U$16402 ( \16745 , \16742 , \16744 );
not \U$16403 ( \16746 , \16745 );
buf \U$16404 ( \16747 , \16746 );
buf \U$16405 ( \16748 , \16747 );
not \U$16406 ( \16749 , \16748 );
or \U$16407 ( \16750 , \16734 , \16749 );
not \U$16408 ( \16751 , \16747 );
nand \U$16409 ( \16752 , \16751 , \16569 );
nand \U$16410 ( \16753 , \16750 , \16752 );
not \U$16411 ( \16754 , \16753 );
not \U$16412 ( \16755 , \1264 );
or \U$16413 ( \16756 , \16754 , \16755 );
nand \U$16414 ( \16757 , \16581 , \1261 );
nand \U$16415 ( \16758 , \16756 , \16757 );
not \U$16416 ( \16759 , \16758 );
xor \U$16417 ( \16760 , \16733 , \16759 );
not \U$16418 ( \16761 , \1077 );
not \U$16419 ( \16762 , \14843 );
not \U$16420 ( \16763 , \1043 );
and \U$16421 ( \16764 , \16762 , \16763 );
not \U$16422 ( \16765 , \14838 );
and \U$16423 ( \16766 , \16765 , \1805 );
nor \U$16424 ( \16767 , \16764 , \16766 );
not \U$16425 ( \16768 , \16767 );
not \U$16426 ( \16769 , \16768 );
or \U$16427 ( \16770 , \16761 , \16769 );
not \U$16428 ( \16771 , RIbb2f160_11);
not \U$16429 ( \16772 , \13475 );
or \U$16430 ( \16773 , \16771 , \16772 );
nand \U$16431 ( \16774 , \13474 , \1048 );
nand \U$16432 ( \16775 , \16773 , \16774 );
nand \U$16433 ( \16776 , \16775 , \1011 );
nand \U$16434 ( \16777 , \16770 , \16776 );
not \U$16435 ( \16778 , \1737 );
not \U$16436 ( \16779 , \16313 );
or \U$16437 ( \16780 , \16778 , \16779 );
not \U$16438 ( \16781 , RIbb2f340_7);
not \U$16439 ( \16782 , \15469 );
not \U$16440 ( \16783 , \16782 );
not \U$16441 ( \16784 , \16783 );
or \U$16442 ( \16785 , \16781 , \16784 );
nand \U$16443 ( \16786 , \15474 , \1734 );
nand \U$16444 ( \16787 , \16785 , \16786 );
nand \U$16445 ( \16788 , \16787 , \1702 );
nand \U$16446 ( \16789 , \16780 , \16788 );
and \U$16447 ( \16790 , \16777 , \16789 );
xor \U$16448 ( \16791 , \16760 , \16790 );
not \U$16449 ( \16792 , \4791 );
not \U$16450 ( \16793 , RIbb2e710_33);
not \U$16451 ( \16794 , \12707 );
or \U$16452 ( \16795 , \16793 , \16794 );
nand \U$16453 ( \16796 , \3654 , \2935 );
nand \U$16454 ( \16797 , \16795 , \16796 );
not \U$16455 ( \16798 , \16797 );
or \U$16456 ( \16799 , \16792 , \16798 );
not \U$16457 ( \16800 , RIbb2e710_33);
not \U$16458 ( \16801 , \4015 );
or \U$16459 ( \16802 , \16800 , \16801 );
not \U$16460 ( \16803 , RIbb2e710_33);
nand \U$16461 ( \16804 , \3022 , \16803 );
nand \U$16462 ( \16805 , \16802 , \16804 );
nand \U$16463 ( \16806 , \16805 , \3887 );
nand \U$16464 ( \16807 , \16799 , \16806 );
xor \U$16465 ( \16808 , \16791 , \16807 );
nand \U$16466 ( \16809 , \16688 , \16808 );
nand \U$16467 ( \16810 , \16683 , \16687 );
nand \U$16468 ( \16811 , \16809 , \16810 );
nand \U$16469 ( \16812 , \16689 , \16694 );
not \U$16470 ( \16813 , \16812 );
and \U$16471 ( \16814 , \16691 , \16813 );
not \U$16472 ( \16815 , \16691 );
and \U$16473 ( \16816 , \16815 , \16812 );
nor \U$16474 ( \16817 , \16814 , \16816 );
buf \U$16475 ( \16818 , \16817 );
not \U$16476 ( \16819 , \16818 );
buf \U$16477 ( \16820 , \16819 );
not \U$16478 ( \16821 , \16820 );
and \U$16479 ( \16822 , \1393 , \16821 );
not \U$16480 ( \16823 , \1261 );
not \U$16481 ( \16824 , \16753 );
or \U$16482 ( \16825 , \16823 , \16824 );
not \U$16483 ( \16826 , \1288 );
not \U$16484 ( \16827 , \16727 );
or \U$16485 ( \16828 , \16826 , \16827 );
not \U$16486 ( \16829 , \16727 );
nand \U$16487 ( \16830 , \16829 , \1244 );
nand \U$16488 ( \16831 , \16828 , \16830 );
nand \U$16489 ( \16832 , \16831 , \1264 );
nand \U$16490 ( \16833 , \16825 , \16832 );
xor \U$16491 ( \16834 , \16822 , \16833 );
not \U$16492 ( \16835 , \1147 );
not \U$16493 ( \16836 , RIbb2f430_5);
not \U$16494 ( \16837 , \16567 );
or \U$16495 ( \16838 , \16836 , \16837 );
nand \U$16496 ( \16839 , \16568 , \1980 );
nand \U$16497 ( \16840 , \16838 , \16839 );
not \U$16498 ( \16841 , \16840 );
or \U$16499 ( \16842 , \16835 , \16841 );
not \U$16500 ( \16843 , RIbb2f430_5);
not \U$16501 ( \16844 , \16575 );
not \U$16502 ( \16845 , \16844 );
or \U$16503 ( \16846 , \16843 , \16845 );
nand \U$16504 ( \16847 , \16575 , \1898 );
nand \U$16505 ( \16848 , \16846 , \16847 );
nand \U$16506 ( \16849 , \16848 , \1089 );
nand \U$16507 ( \16850 , \16842 , \16849 );
xor \U$16508 ( \16851 , \16834 , \16850 );
not \U$16509 ( \16852 , \1089 );
not \U$16510 ( \16853 , RIbb2f430_5);
not \U$16511 ( \16854 , \16747 );
or \U$16512 ( \16855 , \16853 , \16854 );
not \U$16513 ( \16856 , \16747 );
nand \U$16514 ( \16857 , \16856 , \1980 );
nand \U$16515 ( \16858 , \16855 , \16857 );
not \U$16516 ( \16859 , \16858 );
or \U$16517 ( \16860 , \16852 , \16859 );
nand \U$16518 ( \16861 , \16848 , \1147 );
nand \U$16519 ( \16862 , \16860 , \16861 );
not \U$16520 ( \16863 , \998 );
not \U$16521 ( \16864 , RIbb2f070_13);
not \U$16522 ( \16865 , \12932 );
not \U$16523 ( \16866 , \16865 );
or \U$16524 ( \16867 , \16864 , \16866 );
nand \U$16525 ( \16868 , \14635 , \1656 );
nand \U$16526 ( \16869 , \16867 , \16868 );
not \U$16527 ( \16870 , \16869 );
or \U$16528 ( \16871 , \16863 , \16870 );
not \U$16529 ( \16872 , RIbb2f070_13);
not \U$16530 ( \16873 , \13809 );
or \U$16531 ( \16874 , \16872 , \16873 );
nand \U$16532 ( \16875 , \14839 , \1656 );
nand \U$16533 ( \16876 , \16874 , \16875 );
nand \U$16534 ( \16877 , \16876 , \916 );
nand \U$16535 ( \16878 , \16871 , \16877 );
xor \U$16536 ( \16879 , \16862 , \16878 );
not \U$16537 ( \16880 , \1737 );
not \U$16538 ( \16881 , \16787 );
or \U$16539 ( \16882 , \16880 , \16881 );
not \U$16540 ( \16883 , RIbb2f340_7);
not \U$16541 ( \16884 , \16563 );
or \U$16542 ( \16885 , \16883 , \16884 );
nand \U$16543 ( \16886 , \15753 , \1734 );
nand \U$16544 ( \16887 , \16885 , \16886 );
nand \U$16545 ( \16888 , \16887 , \1702 );
nand \U$16546 ( \16889 , \16882 , \16888 );
and \U$16547 ( \16890 , \16879 , \16889 );
and \U$16548 ( \16891 , \16862 , \16878 );
or \U$16549 ( \16892 , \16890 , \16891 );
xor \U$16550 ( \16893 , \16851 , \16892 );
not \U$16551 ( \16894 , \5845 );
not \U$16552 ( \16895 , \16408 );
or \U$16553 ( \16896 , \16894 , \16895 );
not \U$16554 ( \16897 , RIbb2e620_35);
not \U$16555 ( \16898 , \3653 );
not \U$16556 ( \16899 , \16898 );
or \U$16557 ( \16900 , \16897 , \16899 );
nand \U$16558 ( \16901 , \3654 , \6002 );
nand \U$16559 ( \16902 , \16900 , \16901 );
nand \U$16560 ( \16903 , \16902 , \4712 );
nand \U$16561 ( \16904 , \16896 , \16903 );
and \U$16562 ( \16905 , \16893 , \16904 );
and \U$16563 ( \16906 , \16851 , \16892 );
or \U$16564 ( \16907 , \16905 , \16906 );
xor \U$16565 ( \16908 , \16273 , \16287 );
xor \U$16566 ( \16909 , \16908 , \16303 );
xor \U$16567 ( \16910 , \16907 , \16909 );
xor \U$16568 ( \16911 , \16194 , \16175 );
xnor \U$16569 ( \16912 , \16911 , \16157 );
and \U$16570 ( \16913 , \16910 , \16912 );
and \U$16571 ( \16914 , \16907 , \16909 );
or \U$16572 ( \16915 , \16913 , \16914 );
xor \U$16573 ( \16916 , \16811 , \16915 );
not \U$16574 ( \16917 , \3465 );
not \U$16575 ( \16918 , RIbb2e9e0_27);
not \U$16576 ( \16919 , \4087 );
or \U$16577 ( \16920 , \16918 , \16919 );
nand \U$16578 ( \16921 , \16153 , \3454 );
nand \U$16579 ( \16922 , \16920 , \16921 );
not \U$16580 ( \16923 , \16922 );
or \U$16581 ( \16924 , \16917 , \16923 );
nand \U$16582 ( \16925 , \16330 , \3445 );
nand \U$16583 ( \16926 , \16924 , \16925 );
not \U$16584 ( \16927 , \2963 );
not \U$16585 ( \16928 , RIbb2ead0_25);
not \U$16586 ( \16929 , \9023 );
or \U$16587 ( \16930 , \16928 , \16929 );
not \U$16588 ( \16931 , RIbb2ead0_25);
nand \U$16589 ( \16932 , \16931 , \6198 );
nand \U$16590 ( \16933 , \16930 , \16932 );
not \U$16591 ( \16934 , \16933 );
or \U$16592 ( \16935 , \16927 , \16934 );
nand \U$16593 ( \16936 , \16351 , \2980 );
nand \U$16594 ( \16937 , \16935 , \16936 );
not \U$16595 ( \16938 , \16937 );
xor \U$16596 ( \16939 , \16926 , \16938 );
not \U$16597 ( \16940 , RIbb2ebc0_23);
not \U$16598 ( \16941 , \8338 );
or \U$16599 ( \16942 , \16940 , \16941 );
not \U$16600 ( \16943 , \8338 );
nand \U$16601 ( \16944 , \16943 , \2073 );
nand \U$16602 ( \16945 , \16942 , \16944 );
not \U$16603 ( \16946 , \16945 );
not \U$16604 ( \16947 , \3406 );
nor \U$16605 ( \16948 , \16946 , \16947 );
not \U$16606 ( \16949 , RIbb2ebc0_23);
not \U$16607 ( \16950 , \9010 );
or \U$16608 ( \16951 , \16949 , \16950 );
not \U$16609 ( \16952 , \14041 );
nand \U$16610 ( \16953 , \16952 , \3388 );
nand \U$16611 ( \16954 , \16951 , \16953 );
and \U$16612 ( \16955 , \16954 , \3383 );
nor \U$16613 ( \16956 , \16948 , \16955 );
xnor \U$16614 ( \16957 , \16939 , \16956 );
not \U$16615 ( \16958 , \16957 );
not \U$16616 ( \16959 , \16958 );
not \U$16617 ( \16960 , \16678 );
not \U$16618 ( \16961 , \16654 );
or \U$16619 ( \16962 , \16960 , \16961 );
nand \U$16620 ( \16963 , \16962 , \16639 );
nand \U$16621 ( \16964 , \16653 , \16677 );
nand \U$16622 ( \16965 , \16963 , \16964 );
not \U$16623 ( \16966 , \16965 );
not \U$16624 ( \16967 , \16966 );
or \U$16625 ( \16968 , \16959 , \16967 );
nand \U$16626 ( \16969 , \16965 , \16957 );
nand \U$16627 ( \16970 , \16968 , \16969 );
not \U$16628 ( \16971 , RIbb2e620_35);
not \U$16629 ( \16972 , \6301 );
or \U$16630 ( \16973 , \16971 , \16972 );
nand \U$16631 ( \16974 , \9707 , \6002 );
nand \U$16632 ( \16975 , \16973 , \16974 );
not \U$16633 ( \16976 , \16975 );
not \U$16634 ( \16977 , \5845 );
or \U$16635 ( \16978 , \16976 , \16977 );
not \U$16636 ( \16979 , \16402 );
nand \U$16637 ( \16980 , \16979 , \4712 );
nand \U$16638 ( \16981 , \16978 , \16980 );
not \U$16639 ( \16982 , \12285 );
not \U$16640 ( \16983 , RIbb2df90_49);
not \U$16641 ( \16984 , \3370 );
or \U$16642 ( \16985 , \16983 , \16984 );
nand \U$16643 ( \16986 , \1687 , \12278 );
nand \U$16644 ( \16987 , \16985 , \16986 );
not \U$16645 ( \16988 , \16987 );
or \U$16646 ( \16989 , \16982 , \16988 );
nand \U$16647 ( \16990 , \16426 , \12167 );
nand \U$16648 ( \16991 , \16989 , \16990 );
xor \U$16649 ( \16992 , \16981 , \16991 );
not \U$16650 ( \16993 , \6251 );
not \U$16651 ( \16994 , \16436 );
or \U$16652 ( \16995 , \16993 , \16994 );
not \U$16653 ( \16996 , RIbb2e530_37);
not \U$16654 ( \16997 , \3516 );
or \U$16655 ( \16998 , \16996 , \16997 );
nand \U$16656 ( \16999 , \12096 , \8701 );
nand \U$16657 ( \17000 , \16998 , \16999 );
nand \U$16658 ( \17001 , \17000 , \6242 );
nand \U$16659 ( \17002 , \16995 , \17001 );
xor \U$16660 ( \17003 , \16992 , \17002 );
and \U$16661 ( \17004 , \16970 , \17003 );
not \U$16662 ( \17005 , \16970 );
not \U$16663 ( \17006 , \17003 );
and \U$16664 ( \17007 , \17005 , \17006 );
nor \U$16665 ( \17008 , \17004 , \17007 );
and \U$16666 ( \17009 , \16916 , \17008 );
and \U$16667 ( \17010 , \16811 , \16915 );
or \U$16668 ( \17011 , \17009 , \17010 );
xor \U$16669 ( \17012 , \16625 , \17011 );
not \U$16670 ( \17013 , \16958 );
not \U$16671 ( \17014 , \16965 );
or \U$16672 ( \17015 , \17013 , \17014 );
not \U$16673 ( \17016 , \16957 );
not \U$16674 ( \17017 , \16966 );
or \U$16675 ( \17018 , \17016 , \17017 );
nand \U$16676 ( \17019 , \17018 , \17003 );
nand \U$16677 ( \17020 , \17015 , \17019 );
not \U$16678 ( \17021 , \17020 );
not \U$16679 ( \17022 , \17021 );
not \U$16680 ( \17023 , \16271 );
not \U$16681 ( \17024 , RIbb2dae0_59);
and \U$16682 ( \17025 , \811 , \17024 );
not \U$16683 ( \17026 , \811 );
and \U$16684 ( \17027 , \17026 , RIbb2dae0_59);
or \U$16685 ( \17028 , \17025 , \17027 );
not \U$16686 ( \17029 , \17028 );
or \U$16687 ( \17030 , \17023 , \17029 );
nand \U$16688 ( \17031 , \16257 , RIbb2dae0_59);
nand \U$16689 ( \17032 , \17030 , \17031 );
not \U$16690 ( \17033 , \1517 );
and \U$16691 ( \17034 , RIbb2ef80_15, \10306 );
not \U$16692 ( \17035 , RIbb2ef80_15);
and \U$16693 ( \17036 , \17035 , \9841 );
or \U$16694 ( \17037 , \17034 , \17036 );
not \U$16695 ( \17038 , \17037 );
or \U$16696 ( \17039 , \17033 , \17038 );
not \U$16697 ( \17040 , \12230 );
xor \U$16698 ( \17041 , RIbb2ef80_15, \17040 );
nand \U$16699 ( \17042 , \17041 , \1445 );
nand \U$16700 ( \17043 , \17039 , \17042 );
xor \U$16701 ( \17044 , \17032 , \17043 );
not \U$16702 ( \17045 , \916 );
not \U$16703 ( \17046 , \16606 );
or \U$16704 ( \17047 , \17045 , \17046 );
not \U$16705 ( \17048 , RIbb2f070_13);
not \U$16706 ( \17049 , \14563 );
or \U$16707 ( \17050 , \17048 , \17049 );
nand \U$16708 ( \17051 , \10764 , \906 );
nand \U$16709 ( \17052 , \17050 , \17051 );
nand \U$16710 ( \17053 , \17052 , \998 );
nand \U$16711 ( \17054 , \17047 , \17053 );
not \U$16712 ( \17055 , \17054 );
xor \U$16713 ( \17056 , \17044 , \17055 );
not \U$16714 ( \17057 , \2077 );
not \U$16715 ( \17058 , \16461 );
or \U$16716 ( \17059 , \17057 , \17058 );
not \U$16717 ( \17060 , RIbb2ecb0_21);
not \U$16718 ( \17061 , \8338 );
or \U$16719 ( \17062 , \17060 , \17061 );
nand \U$16720 ( \17063 , \8339 , \2067 );
nand \U$16721 ( \17064 , \17062 , \17063 );
nand \U$16722 ( \17065 , \17064 , \2078 );
nand \U$16723 ( \17066 , \17059 , \17065 );
not \U$16724 ( \17067 , \854 );
not \U$16725 ( \17068 , RIbb2eda0_19);
not \U$16726 ( \17069 , \13850 );
or \U$16727 ( \17070 , \17068 , \17069 );
nand \U$16728 ( \17071 , \13854 , \1776 );
nand \U$16729 ( \17072 , \17070 , \17071 );
not \U$16730 ( \17073 , \17072 );
or \U$16731 ( \17074 , \17067 , \17073 );
nand \U$16732 ( \17075 , \16497 , \853 );
nand \U$16733 ( \17076 , \17074 , \17075 );
xor \U$16734 ( \17077 , \17066 , \17076 );
not \U$16735 ( \17078 , \836 );
not \U$16736 ( \17079 , \822 );
not \U$16737 ( \17080 , \10178 );
or \U$16738 ( \17081 , \17079 , \17080 );
not \U$16739 ( \17082 , \13866 );
nand \U$16740 ( \17083 , \17082 , RIbb2ee90_17);
nand \U$16741 ( \17084 , \17081 , \17083 );
not \U$16742 ( \17085 , \17084 );
or \U$16743 ( \17086 , \17078 , \17085 );
nand \U$16744 ( \17087 , \16477 , \832 );
nand \U$16745 ( \17088 , \17086 , \17087 );
xor \U$16746 ( \17089 , \17077 , \17088 );
xor \U$16747 ( \17090 , \17056 , \17089 );
not \U$16748 ( \17091 , \16674 );
not \U$16749 ( \17092 , \16665 );
or \U$16750 ( \17093 , \17091 , \17092 );
not \U$16751 ( \17094 , RIbb2dbd0_57);
not \U$16752 ( \17095 , \8754 );
or \U$16753 ( \17096 , \17094 , \17095 );
not \U$16754 ( \17097 , RIbb2dbd0_57);
nand \U$16755 ( \17098 , \13308 , \17097 );
nand \U$16756 ( \17099 , \17096 , \17098 );
buf \U$16757 ( \17100 , \15738 );
nand \U$16758 ( \17101 , \17099 , \17100 );
nand \U$16759 ( \17102 , \17093 , \17101 );
not \U$16760 ( \17103 , \14067 );
not \U$16761 ( \17104 , \16630 );
or \U$16762 ( \17105 , \17103 , \17104 );
and \U$16763 ( \17106 , RIbb2dea0_51, \5003 );
not \U$16764 ( \17107 , RIbb2dea0_51);
and \U$16765 ( \17108 , \17107 , \1548 );
or \U$16766 ( \17109 , \17106 , \17108 );
nand \U$16767 ( \17110 , \17109 , \12692 );
nand \U$16768 ( \17111 , \17105 , \17110 );
xor \U$16769 ( \17112 , \17102 , \17111 );
not \U$16770 ( \17113 , \7104 );
not \U$16771 ( \17114 , \16235 );
not \U$16772 ( \17115 , \10908 );
and \U$16773 ( \17116 , \17114 , \17115 );
and \U$16774 ( \17117 , \13280 , \10908 );
nor \U$16775 ( \17118 , \17116 , \17117 );
not \U$16776 ( \17119 , \17118 );
not \U$16777 ( \17120 , \17119 );
or \U$16778 ( \17121 , \17113 , \17120 );
nand \U$16779 ( \17122 , \16645 , \8445 );
nand \U$16780 ( \17123 , \17121 , \17122 );
and \U$16781 ( \17124 , \17112 , \17123 );
and \U$16782 ( \17125 , \17102 , \17111 );
or \U$16783 ( \17126 , \17124 , \17125 );
xor \U$16784 ( \17127 , \17090 , \17126 );
not \U$16785 ( \17128 , \17127 );
not \U$16786 ( \17129 , \17128 );
or \U$16787 ( \17130 , \17022 , \17129 );
nand \U$16788 ( \17131 , \17127 , \17020 );
nand \U$16789 ( \17132 , \17130 , \17131 );
not \U$16790 ( \17133 , \14613 );
not \U$16791 ( \17134 , \16285 );
or \U$16792 ( \17135 , \17133 , \17134 );
and \U$16793 ( \17136 , RIbb2dcc0_55, \15556 );
not \U$16794 ( \17137 , RIbb2dcc0_55);
and \U$16795 ( \17138 , \17137 , \986 );
or \U$16796 ( \17139 , \17136 , \17138 );
nand \U$16797 ( \17140 , \17139 , \15182 );
nand \U$16798 ( \17141 , \17135 , \17140 );
not \U$16799 ( \17142 , \17141 );
not \U$16800 ( \17143 , \16271 );
not \U$16801 ( \17144 , \16262 );
or \U$16802 ( \17145 , \17143 , \17144 );
nand \U$16803 ( \17146 , \16257 , \17028 );
nand \U$16804 ( \17147 , \17145 , \17146 );
not \U$16805 ( \17148 , \17147 );
or \U$16806 ( \17149 , \17142 , \17148 );
not \U$16807 ( \17150 , \17147 );
not \U$16808 ( \17151 , \17150 );
not \U$16809 ( \17152 , \17141 );
not \U$16810 ( \17153 , \17152 );
or \U$16811 ( \17154 , \17151 , \17153 );
not \U$16812 ( \17155 , \10119 );
not \U$16813 ( \17156 , RIbb2e170_45);
not \U$16814 ( \17157 , \3290 );
or \U$16815 ( \17158 , \17156 , \17157 );
nand \U$16816 ( \17159 , \1283 , \9094 );
nand \U$16817 ( \17160 , \17158 , \17159 );
not \U$16818 ( \17161 , \17160 );
or \U$16819 ( \17162 , \17155 , \17161 );
nand \U$16820 ( \17163 , \16301 , \10117 );
nand \U$16821 ( \17164 , \17162 , \17163 );
nand \U$16822 ( \17165 , \17154 , \17164 );
nand \U$16823 ( \17166 , \17149 , \17165 );
not \U$16824 ( \17167 , \11176 );
not \U$16825 ( \17168 , \16173 );
or \U$16826 ( \17169 , \17167 , \17168 );
and \U$16827 ( \17170 , RIbb2e080_47, \3054 );
not \U$16828 ( \17171 , RIbb2e080_47);
and \U$16829 ( \17172 , \17171 , \10673 );
or \U$16830 ( \17173 , \17170 , \17172 );
nand \U$16831 ( \17174 , \17173 , \12965 );
nand \U$16832 ( \17175 , \17169 , \17174 );
buf \U$16833 ( \17176 , \17175 );
not \U$16834 ( \17177 , \17176 );
not \U$16835 ( \17178 , \2925 );
not \U$16836 ( \17179 , RIbb2e8f0_29);
not \U$16837 ( \17180 , \3276 );
or \U$16838 ( \17181 , \17179 , \17180 );
nand \U$16839 ( \17182 , \3003 , \3800 );
nand \U$16840 ( \17183 , \17181 , \17182 );
not \U$16841 ( \17184 , \17183 );
or \U$16842 ( \17185 , \17178 , \17184 );
nand \U$16843 ( \17186 , \16147 , \2922 );
nand \U$16844 ( \17187 , \17185 , \17186 );
not \U$16845 ( \17188 , \17187 );
or \U$16846 ( \17189 , \17177 , \17188 );
or \U$16847 ( \17190 , \17176 , \17187 );
not \U$16848 ( \17191 , \2940 );
not \U$16849 ( \17192 , \16187 );
not \U$16850 ( \17193 , \17192 );
or \U$16851 ( \17194 , \17191 , \17193 );
not \U$16852 ( \17195 , RIbb2e800_31);
not \U$16853 ( \17196 , \15443 );
or \U$16854 ( \17197 , \17195 , \17196 );
nand \U$16855 ( \17198 , \3022 , \9169 );
nand \U$16856 ( \17199 , \17197 , \17198 );
nand \U$16857 ( \17200 , \17199 , \2941 );
nand \U$16858 ( \17201 , \17194 , \17200 );
nand \U$16859 ( \17202 , \17190 , \17201 );
nand \U$16860 ( \17203 , \17189 , \17202 );
xor \U$16861 ( \17204 , \17166 , \17203 );
not \U$16862 ( \17205 , \8995 );
not \U$16863 ( \17206 , RIbb2e350_41);
not \U$16864 ( \17207 , \1337 );
not \U$16865 ( \17208 , \17207 );
or \U$16866 ( \17209 , \17206 , \17208 );
nand \U$16867 ( \17210 , \3495 , \9402 );
nand \U$16868 ( \17211 , \17209 , \17210 );
not \U$16869 ( \17212 , \17211 );
or \U$16870 ( \17213 , \17205 , \17212 );
nand \U$16871 ( \17214 , \8362 , \16244 );
nand \U$16872 ( \17215 , \17213 , \17214 );
not \U$16873 ( \17216 , \14930 );
not \U$16874 ( \17217 , RIbb2ddb0_53);
not \U$16875 ( \17218 , \1070 );
or \U$16876 ( \17219 , \17217 , \17218 );
nand \U$16877 ( \17220 , \1886 , \13463 );
nand \U$16878 ( \17221 , \17219 , \17220 );
not \U$16879 ( \17222 , \17221 );
or \U$16880 ( \17223 , \17216 , \17222 );
nand \U$16881 ( \17224 , \16212 , \13467 );
nand \U$16882 ( \17225 , \17223 , \17224 );
or \U$16883 ( \17226 , \17215 , \17225 );
not \U$16884 ( \17227 , \10451 );
not \U$16885 ( \17228 , RIbb2e260_43);
not \U$16886 ( \17229 , \12024 );
or \U$16887 ( \17230 , \17228 , \17229 );
not \U$16888 ( \17231 , RIbb2e260_43);
nand \U$16889 ( \17232 , \4340 , \17231 );
nand \U$16890 ( \17233 , \17230 , \17232 );
not \U$16891 ( \17234 , \17233 );
or \U$16892 ( \17235 , \17227 , \17234 );
nand \U$16893 ( \17236 , \16220 , \10449 );
nand \U$16894 ( \17237 , \17235 , \17236 );
nand \U$16895 ( \17238 , \17226 , \17237 );
nand \U$16896 ( \17239 , \17215 , \17225 );
nand \U$16897 ( \17240 , \17238 , \17239 );
xor \U$16898 ( \17241 , \17204 , \17240 );
and \U$16899 ( \17242 , \17132 , \17241 );
not \U$16900 ( \17243 , \17132 );
not \U$16901 ( \17244 , \17241 );
and \U$16902 ( \17245 , \17243 , \17244 );
nor \U$16903 ( \17246 , \17242 , \17245 );
xor \U$16904 ( \17247 , \17012 , \17246 );
xor \U$16905 ( \17248 , \16811 , \16915 );
xor \U$16906 ( \17249 , \17248 , \17008 );
xor \U$16907 ( \17250 , \16907 , \16909 );
xor \U$16908 ( \17251 , \17250 , \16912 );
not \U$16909 ( \17252 , \17251 );
and \U$16910 ( \17253 , \16682 , \16685 );
not \U$16911 ( \17254 , \16682 );
and \U$16912 ( \17255 , \17254 , \16686 );
nor \U$16913 ( \17256 , \17253 , \17255 );
xor \U$16914 ( \17257 , \17256 , \16808 );
buf \U$16915 ( \17258 , \17257 );
nand \U$16916 ( \17259 , \17252 , \17258 );
not \U$16917 ( \17260 , \17259 );
xor \U$16918 ( \17261 , \16777 , \16789 );
not \U$16919 ( \17262 , RIbb2d900_63);
not \U$16920 ( \17263 , \17262 );
not \U$16921 ( \17264 , RIbb2d888_64);
not \U$16922 ( \17265 , \17264 );
and \U$16923 ( \17266 , \17263 , \17265 );
not \U$16924 ( \17267 , RIbb2d900_63);
not \U$16925 ( \17268 , \812 );
or \U$16926 ( \17269 , \17267 , \17268 );
not \U$16927 ( \17270 , RIbb2d900_63);
nand \U$16928 ( \17271 , \811 , \17270 );
nand \U$16929 ( \17272 , \17269 , \17271 );
and \U$16930 ( \17273 , \17264 , RIbb2d900_63);
buf \U$16931 ( \17274 , \17273 );
buf \U$16932 ( \17275 , \17274 );
and \U$16933 ( \17276 , \17272 , \17275 );
nor \U$16934 ( \17277 , \17266 , \17276 );
not \U$16935 ( \17278 , \17277 );
not \U$16936 ( \17279 , \1517 );
and \U$16937 ( \17280 , RIbb2ef80_15, \14885 );
not \U$16938 ( \17281 , RIbb2ef80_15);
and \U$16939 ( \17282 , \17281 , \11580 );
nor \U$16940 ( \17283 , \17280 , \17282 );
not \U$16941 ( \17284 , \17283 );
or \U$16942 ( \17285 , \17279 , \17284 );
not \U$16943 ( \17286 , \1575 );
not \U$16944 ( \17287 , \13680 );
xor \U$16945 ( \17288 , RIbb2ef80_15, \17287 );
nand \U$16946 ( \17289 , \17286 , \17288 );
nand \U$16947 ( \17290 , \17285 , \17289 );
or \U$16948 ( \17291 , \17278 , \17290 );
not \U$16949 ( \17292 , \832 );
not \U$16950 ( \17293 , RIbb2ee90_17);
not \U$16951 ( \17294 , \11142 );
not \U$16952 ( \17295 , \17294 );
or \U$16953 ( \17296 , \17293 , \17295 );
not \U$16954 ( \17297 , \12260 );
nand \U$16955 ( \17298 , \17297 , \3057 );
nand \U$16956 ( \17299 , \17296 , \17298 );
not \U$16957 ( \17300 , \17299 );
or \U$16958 ( \17301 , \17292 , \17300 );
not \U$16959 ( \17302 , RIbb2ee90_17);
not \U$16960 ( \17303 , \12764 );
or \U$16961 ( \17304 , \17302 , \17303 );
nand \U$16962 ( \17305 , \13525 , \3057 );
nand \U$16963 ( \17306 , \17304 , \17305 );
nand \U$16964 ( \17307 , \17306 , \836 );
nand \U$16965 ( \17308 , \17301 , \17307 );
nand \U$16966 ( \17309 , \17291 , \17308 );
nand \U$16967 ( \17310 , \17290 , \17278 );
nand \U$16968 ( \17311 , \17309 , \17310 );
xor \U$16969 ( \17312 , \17261 , \17311 );
not \U$16970 ( \17313 , \1570 );
not \U$16971 ( \17314 , RIbb2f250_9);
buf \U$16972 ( \17315 , \13546 );
not \U$16973 ( \17316 , \17315 );
or \U$16974 ( \17317 , \17314 , \17316 );
nand \U$16975 ( \17318 , \13547 , \5064 );
nand \U$16976 ( \17319 , \17317 , \17318 );
not \U$16977 ( \17320 , \17319 );
or \U$16978 ( \17321 , \17313 , \17320 );
not \U$16979 ( \17322 , RIbb2f250_9);
not \U$16980 ( \17323 , \14503 );
or \U$16981 ( \17324 , \17322 , \17323 );
nand \U$16982 ( \17325 , \16320 , \1554 );
nand \U$16983 ( \17326 , \17324 , \17325 );
nand \U$16984 ( \17327 , \17326 , \1533 );
nand \U$16985 ( \17328 , \17321 , \17327 );
not \U$16986 ( \17329 , \998 );
not \U$16987 ( \17330 , RIbb2f070_13);
not \U$16988 ( \17331 , \13680 );
or \U$16989 ( \17332 , \17330 , \17331 );
nand \U$16990 ( \17333 , \12175 , \906 );
nand \U$16991 ( \17334 , \17332 , \17333 );
not \U$16992 ( \17335 , \17334 );
or \U$16993 ( \17336 , \17329 , \17335 );
nand \U$16994 ( \17337 , \16869 , \916 );
nand \U$16995 ( \17338 , \17336 , \17337 );
xor \U$16996 ( \17339 , \17328 , \17338 );
not \U$16997 ( \17340 , \3445 );
not \U$16998 ( \17341 , \8387 );
and \U$16999 ( \17342 , RIbb2e9e0_27, \17341 );
not \U$17000 ( \17343 , RIbb2e9e0_27);
and \U$17001 ( \17344 , \17343 , \7111 );
or \U$17002 ( \17345 , \17342 , \17344 );
not \U$17003 ( \17346 , \17345 );
or \U$17004 ( \17347 , \17340 , \17346 );
nand \U$17005 ( \17348 , \16338 , \3465 );
nand \U$17006 ( \17349 , \17347 , \17348 );
xor \U$17007 ( \17350 , \17339 , \17349 );
xor \U$17008 ( \17351 , \17312 , \17350 );
not \U$17009 ( \17352 , \17275 );
xor \U$17010 ( \17353 , RIbb2d900_63, \892 );
not \U$17011 ( \17354 , \17353 );
or \U$17012 ( \17355 , \17352 , \17354 );
nand \U$17013 ( \17356 , \17272 , RIbb2d888_64);
nand \U$17014 ( \17357 , \17355 , \17356 );
not \U$17015 ( \17358 , \12284 );
not \U$17016 ( \17359 , RIbb2df90_49);
not \U$17017 ( \17360 , \12037 );
or \U$17018 ( \17361 , \17359 , \17360 );
not \U$17019 ( \17362 , RIbb2df90_49);
nand \U$17020 ( \17363 , \17362 , \12036 );
nand \U$17021 ( \17364 , \17361 , \17363 );
not \U$17022 ( \17365 , \17364 );
or \U$17023 ( \17366 , \17358 , \17365 );
and \U$17024 ( \17367 , \12278 , \1170 );
not \U$17025 ( \17368 , \12278 );
not \U$17026 ( \17369 , \1169 );
not \U$17027 ( \17370 , \17369 );
and \U$17028 ( \17371 , \17368 , \17370 );
nor \U$17029 ( \17372 , \17367 , \17371 );
nand \U$17030 ( \17373 , \17372 , \12167 );
nand \U$17031 ( \17374 , \17366 , \17373 );
xor \U$17032 ( \17375 , \17357 , \17374 );
not \U$17033 ( \17376 , \11177 );
not \U$17034 ( \17377 , RIbb2e080_47);
not \U$17035 ( \17378 , \12024 );
or \U$17036 ( \17379 , \17377 , \17378 );
not \U$17037 ( \17380 , \13619 );
nand \U$17038 ( \17381 , \17380 , \11959 );
nand \U$17039 ( \17382 , \17379 , \17381 );
not \U$17040 ( \17383 , \17382 );
or \U$17041 ( \17384 , \17376 , \17383 );
not \U$17042 ( \17385 , RIbb2e080_47);
not \U$17043 ( \17386 , \1419 );
not \U$17044 ( \17387 , \17386 );
or \U$17045 ( \17388 , \17385 , \17387 );
nand \U$17046 ( \17389 , \3821 , \10113 );
nand \U$17047 ( \17390 , \17388 , \17389 );
nand \U$17048 ( \17391 , \17390 , \11176 );
nand \U$17049 ( \17392 , \17384 , \17391 );
and \U$17050 ( \17393 , \17375 , \17392 );
and \U$17051 ( \17394 , \17357 , \17374 );
or \U$17052 ( \17395 , \17393 , \17394 );
not \U$17053 ( \17396 , \17395 );
buf \U$17054 ( \17397 , \15738 );
not \U$17055 ( \17398 , \17397 );
not \U$17056 ( \17399 , RIbb2dbd0_57);
not \U$17057 ( \17400 , \4284 );
or \U$17058 ( \17401 , \17399 , \17400 );
nand \U$17059 ( \17402 , \1886 , \14602 );
nand \U$17060 ( \17403 , \17401 , \17402 );
not \U$17061 ( \17404 , \17403 );
or \U$17062 ( \17405 , \17398 , \17404 );
not \U$17063 ( \17406 , RIbb2dbd0_57);
not \U$17064 ( \17407 , \1560 );
not \U$17065 ( \17408 , \17407 );
or \U$17066 ( \17409 , \17406 , \17408 );
not \U$17067 ( \17410 , \16207 );
not \U$17068 ( \17411 , RIbb2dbd0_57);
nand \U$17069 ( \17412 , \17410 , \17411 );
nand \U$17070 ( \17413 , \17409 , \17412 );
nand \U$17071 ( \17414 , \17413 , \16675 );
nand \U$17072 ( \17415 , \17405 , \17414 );
not \U$17073 ( \17416 , \17415 );
not \U$17074 ( \17417 , \17416 );
not \U$17075 ( \17418 , \3887 );
not \U$17076 ( \17419 , RIbb2e710_33);
not \U$17077 ( \17420 , \3090 );
or \U$17078 ( \17421 , \17419 , \17420 );
nand \U$17079 ( \17422 , \3091 , \13352 );
nand \U$17080 ( \17423 , \17421 , \17422 );
not \U$17081 ( \17424 , \17423 );
or \U$17082 ( \17425 , \17418 , \17424 );
not \U$17083 ( \17426 , RIbb2e710_33);
not \U$17084 ( \17427 , \13731 );
or \U$17085 ( \17428 , \17426 , \17427 );
nand \U$17086 ( \17429 , \13732 , \3864 );
nand \U$17087 ( \17430 , \17428 , \17429 );
nand \U$17088 ( \17431 , \17430 , \4791 );
nand \U$17089 ( \17432 , \17425 , \17431 );
not \U$17090 ( \17433 , \17432 );
not \U$17091 ( \17434 , \17433 );
or \U$17092 ( \17435 , \17417 , \17434 );
not \U$17093 ( \17436 , \836 );
not \U$17094 ( \17437 , \17299 );
or \U$17095 ( \17438 , \17436 , \17437 );
not \U$17096 ( \17439 , RIbb2ee90_17);
not \U$17097 ( \17440 , \11578 );
not \U$17098 ( \17441 , \17440 );
or \U$17099 ( \17442 , \17439 , \17441 );
nand \U$17100 ( \17443 , \11578 , \3057 );
nand \U$17101 ( \17444 , \17442 , \17443 );
nand \U$17102 ( \17445 , \17444 , \832 );
nand \U$17103 ( \17446 , \17438 , \17445 );
nand \U$17104 ( \17447 , \17435 , \17446 );
not \U$17105 ( \17448 , \17416 );
nand \U$17106 ( \17449 , \17448 , \17432 );
nand \U$17107 ( \17450 , \17447 , \17449 );
not \U$17108 ( \17451 , \17450 );
or \U$17109 ( \17452 , \17396 , \17451 );
or \U$17110 ( \17453 , \17450 , \17395 );
not \U$17111 ( \17454 , \8362 );
not \U$17112 ( \17455 , RIbb2e350_41);
not \U$17113 ( \17456 , \4219 );
or \U$17114 ( \17457 , \17455 , \17456 );
nand \U$17115 ( \17458 , \3166 , \13392 );
nand \U$17116 ( \17459 , \17457 , \17458 );
not \U$17117 ( \17460 , \17459 );
or \U$17118 ( \17461 , \17454 , \17460 );
not \U$17119 ( \17462 , RIbb2e350_41);
not \U$17120 ( \17463 , \3516 );
or \U$17121 ( \17464 , \17462 , \17463 );
nand \U$17122 ( \17465 , \3341 , \7097 );
nand \U$17123 ( \17466 , \17464 , \17465 );
nand \U$17124 ( \17467 , \17466 , \8353 );
nand \U$17125 ( \17468 , \17461 , \17467 );
not \U$17126 ( \17469 , \17468 );
buf \U$17127 ( \17470 , \16257 );
not \U$17128 ( \17471 , \17470 );
and \U$17129 ( \17472 , RIbb2dae0_59, \15556 );
not \U$17130 ( \17473 , RIbb2dae0_59);
not \U$17131 ( \17474 , \15556 );
and \U$17132 ( \17475 , \17473 , \17474 );
or \U$17133 ( \17476 , \17472 , \17475 );
not \U$17134 ( \17477 , \17476 );
or \U$17135 ( \17478 , \17471 , \17477 );
xor \U$17136 ( \17479 , RIbb2dae0_59, \950 );
nand \U$17137 ( \17480 , \17479 , \16271 );
nand \U$17138 ( \17481 , \17478 , \17480 );
not \U$17139 ( \17482 , \17481 );
or \U$17140 ( \17483 , \17469 , \17482 );
or \U$17141 ( \17484 , \17481 , \17468 );
not \U$17142 ( \17485 , \9099 );
not \U$17143 ( \17486 , RIbb2e260_43);
not \U$17144 ( \17487 , \9983 );
or \U$17145 ( \17488 , \17486 , \17487 );
nand \U$17146 ( \17489 , \16235 , \13772 );
nand \U$17147 ( \17490 , \17488 , \17489 );
not \U$17148 ( \17491 , \17490 );
or \U$17149 ( \17492 , \17485 , \17491 );
not \U$17150 ( \17493 , RIbb2e260_43);
not \U$17151 ( \17494 , \13289 );
or \U$17152 ( \17495 , \17493 , \17494 );
nand \U$17153 ( \17496 , \2222 , \8347 );
nand \U$17154 ( \17497 , \17495 , \17496 );
nand \U$17155 ( \17498 , \17497 , \9098 );
nand \U$17156 ( \17499 , \17492 , \17498 );
nand \U$17157 ( \17500 , \17484 , \17499 );
nand \U$17158 ( \17501 , \17483 , \17500 );
nand \U$17159 ( \17502 , \17453 , \17501 );
nand \U$17160 ( \17503 , \17452 , \17502 );
xor \U$17161 ( \17504 , \17351 , \17503 );
xor \U$17162 ( \17505 , RIbb33378_192, RIbb31578_128);
buf \U$17163 ( \17506 , \17505 );
and \U$17164 ( \17507 , \1312 , \17506 );
not \U$17165 ( \17508 , \467 );
buf \U$17166 ( \17509 , \465 );
nor \U$17167 ( \17510 , \17508 , \17509 );
buf \U$17168 ( \17511 , \464 );
not \U$17169 ( \17512 , \17511 );
and \U$17170 ( \17513 , \17510 , \17512 );
not \U$17171 ( \17514 , \17510 );
and \U$17172 ( \17515 , \17514 , \17511 );
nor \U$17173 ( \17516 , \17513 , \17515 );
buf \U$17174 ( \17517 , \17516 );
buf \U$17175 ( \17518 , \17517 );
not \U$17176 ( \17519 , \17518 );
buf \U$17177 ( \17520 , \17519 );
and \U$17178 ( \17521 , \17520 , \13990 );
not \U$17179 ( \17522 , \17520 );
not \U$17180 ( \17523 , \1391 );
and \U$17181 ( \17524 , \17522 , \17523 );
nor \U$17182 ( \17525 , \17521 , \17524 );
not \U$17183 ( \17526 , \17525 );
not \U$17184 ( \17527 , \1428 );
or \U$17185 ( \17528 , \17526 , \17527 );
buf \U$17186 ( \17529 , \16817 );
not \U$17187 ( \17530 , \17529 );
not \U$17188 ( \17531 , \1392 );
or \U$17189 ( \17532 , \17530 , \17531 );
nand \U$17190 ( \17533 , \17523 , \16820 );
nand \U$17191 ( \17534 , \17532 , \17533 );
nand \U$17192 ( \17535 , \1375 , \17534 );
nand \U$17193 ( \17536 , \17528 , \17535 );
xor \U$17194 ( \17537 , \17507 , \17536 );
not \U$17195 ( \17538 , \1737 );
not \U$17196 ( \17539 , \16887 );
or \U$17197 ( \17540 , \17538 , \17539 );
not \U$17198 ( \17541 , RIbb2f340_7);
not \U$17199 ( \17542 , \15824 );
or \U$17200 ( \17543 , \17541 , \17542 );
nand \U$17201 ( \17544 , \16576 , \1734 );
nand \U$17202 ( \17545 , \17543 , \17544 );
nand \U$17203 ( \17546 , \17545 , \1702 );
nand \U$17204 ( \17547 , \17540 , \17546 );
xor \U$17205 ( \17548 , \17537 , \17547 );
not \U$17206 ( \17549 , \14930 );
not \U$17207 ( \17550 , RIbb2ddb0_53);
not \U$17208 ( \17551 , \16633 );
or \U$17209 ( \17552 , \17550 , \17551 );
nand \U$17210 ( \17553 , \3369 , \13941 );
nand \U$17211 ( \17554 , \17552 , \17553 );
not \U$17212 ( \17555 , \17554 );
or \U$17213 ( \17556 , \17549 , \17555 );
not \U$17214 ( \17557 , RIbb2ddb0_53);
not \U$17215 ( \17558 , \1641 );
or \U$17216 ( \17559 , \17557 , \17558 );
nand \U$17217 ( \17560 , \8856 , \12681 );
nand \U$17218 ( \17561 , \17559 , \17560 );
not \U$17219 ( \17562 , \13466 );
buf \U$17220 ( \17563 , \17562 );
nand \U$17221 ( \17564 , \17561 , \17563 );
nand \U$17222 ( \17565 , \17556 , \17564 );
xor \U$17223 ( \17566 , \17548 , \17565 );
not \U$17224 ( \17567 , \7104 );
not \U$17225 ( \17568 , \3139 );
and \U$17226 ( \17569 , RIbb2e440_39, \17568 );
not \U$17227 ( \17570 , RIbb2e440_39);
and \U$17228 ( \17571 , \17570 , \3139 );
or \U$17229 ( \17572 , \17569 , \17571 );
not \U$17230 ( \17573 , \17572 );
or \U$17231 ( \17574 , \17567 , \17573 );
and \U$17232 ( \17575 , RIbb2e440_39, \16399 );
not \U$17233 ( \17576 , RIbb2e440_39);
and \U$17234 ( \17577 , \17576 , \4637 );
or \U$17235 ( \17578 , \17575 , \17577 );
nand \U$17236 ( \17579 , \17578 , \7103 );
nand \U$17237 ( \17580 , \17574 , \17579 );
and \U$17238 ( \17581 , \17566 , \17580 );
and \U$17239 ( \17582 , \17548 , \17565 );
or \U$17240 ( \17583 , \17581 , \17582 );
not \U$17241 ( \17584 , \6242 );
not \U$17242 ( \17585 , RIbb2e530_37);
not \U$17243 ( \17586 , \6172 );
or \U$17244 ( \17587 , \17585 , \17586 );
nand \U$17245 ( \17588 , \13903 , \6246 );
nand \U$17246 ( \17589 , \17587 , \17588 );
not \U$17247 ( \17590 , \17589 );
or \U$17248 ( \17591 , \17584 , \17590 );
not \U$17249 ( \17592 , RIbb2e530_37);
not \U$17250 ( \17593 , \16898 );
or \U$17251 ( \17594 , \17592 , \17593 );
nand \U$17252 ( \17595 , \3653 , \6246 );
nand \U$17253 ( \17596 , \17594 , \17595 );
nand \U$17254 ( \17597 , \6251 , \17596 );
nand \U$17255 ( \17598 , \17591 , \17597 );
not \U$17256 ( \17599 , \12692 );
and \U$17257 ( \17600 , RIbb2dea0_51, \8862 );
not \U$17258 ( \17601 , RIbb2dea0_51);
and \U$17259 ( \17602 , \17601 , \1137 );
or \U$17260 ( \17603 , \17600 , \17602 );
not \U$17261 ( \17604 , \17603 );
or \U$17262 ( \17605 , \17599 , \17604 );
not \U$17263 ( \17606 , RIbb2dea0_51);
not \U$17264 ( \17607 , \1112 );
or \U$17265 ( \17608 , \17606 , \17607 );
not \U$17266 ( \17609 , RIbb2dea0_51);
nand \U$17267 ( \17610 , \17609 , \4769 );
nand \U$17268 ( \17611 , \17608 , \17610 );
nand \U$17269 ( \17612 , \17611 , \14067 );
nand \U$17270 ( \17613 , \17605 , \17612 );
xor \U$17271 ( \17614 , \17598 , \17613 );
not \U$17272 ( \17615 , \4712 );
not \U$17273 ( \17616 , RIbb2e620_35);
not \U$17274 ( \17617 , \3045 );
or \U$17275 ( \17618 , \17616 , \17617 );
nand \U$17276 ( \17619 , \12596 , \3866 );
nand \U$17277 ( \17620 , \17618 , \17619 );
not \U$17278 ( \17621 , \17620 );
or \U$17279 ( \17622 , \17615 , \17621 );
not \U$17280 ( \17623 , RIbb2e620_35);
not \U$17281 ( \17624 , \3023 );
or \U$17282 ( \17625 , \17623 , \17624 );
nand \U$17283 ( \17626 , \3022 , \3866 );
nand \U$17284 ( \17627 , \17625 , \17626 );
nand \U$17285 ( \17628 , \17627 , \5845 );
nand \U$17286 ( \17629 , \17622 , \17628 );
and \U$17287 ( \17630 , \17614 , \17629 );
and \U$17288 ( \17631 , \17598 , \17613 );
or \U$17289 ( \17632 , \17630 , \17631 );
xor \U$17290 ( \17633 , \17583 , \17632 );
xor \U$17291 ( \17634 , \17277 , \17290 );
xnor \U$17292 ( \17635 , \17634 , \17308 );
and \U$17293 ( \17636 , \17633 , \17635 );
and \U$17294 ( \17637 , \17583 , \17632 );
or \U$17295 ( \17638 , \17636 , \17637 );
and \U$17296 ( \17639 , \17504 , \17638 );
and \U$17297 ( \17640 , \17351 , \17503 );
or \U$17298 ( \17641 , \17639 , \17640 );
not \U$17299 ( \17642 , \17641 );
or \U$17300 ( \17643 , \17260 , \17642 );
not \U$17301 ( \17644 , \17258 );
nand \U$17302 ( \17645 , \17644 , \17251 );
nand \U$17303 ( \17646 , \17643 , \17645 );
xor \U$17304 ( \17647 , \17249 , \17646 );
xor \U$17305 ( \17648 , \17102 , \17111 );
xor \U$17306 ( \17649 , \17648 , \17123 );
not \U$17307 ( \17650 , \17649 );
not \U$17308 ( \17651 , \17650 );
xor \U$17309 ( \17652 , \17175 , \17201 );
xnor \U$17310 ( \17653 , \17652 , \17187 );
not \U$17311 ( \17654 , \17653 );
not \U$17312 ( \17655 , \17654 );
or \U$17313 ( \17656 , \17651 , \17655 );
nand \U$17314 ( \17657 , \17653 , \17649 );
nand \U$17315 ( \17658 , \17656 , \17657 );
xor \U$17316 ( \17659 , \16705 , \16732 );
and \U$17317 ( \17660 , \17659 , \16759 );
and \U$17318 ( \17661 , \16705 , \16732 );
or \U$17319 ( \17662 , \17660 , \17661 );
not \U$17320 ( \17663 , \12321 );
not \U$17321 ( \17664 , \17663 );
not \U$17322 ( \17665 , \17664 );
not \U$17323 ( \17666 , \1805 );
and \U$17324 ( \17667 , \17665 , \17666 );
and \U$17325 ( \17668 , \14635 , \1048 );
nor \U$17326 ( \17669 , \17667 , \17668 );
not \U$17327 ( \17670 , \17669 );
not \U$17328 ( \17671 , \1943 );
and \U$17329 ( \17672 , \17670 , \17671 );
nor \U$17330 ( \17673 , \16767 , \2122 );
nor \U$17331 ( \17674 , \17672 , \17673 );
not \U$17332 ( \17675 , \17674 );
not \U$17333 ( \17676 , \17675 );
not \U$17334 ( \17677 , \1147 );
not \U$17335 ( \17678 , RIbb2f430_5);
not \U$17336 ( \17679 , \15471 );
or \U$17337 ( \17680 , \17678 , \17679 );
buf \U$17338 ( \17681 , \15469 );
not \U$17339 ( \17682 , \17681 );
nand \U$17340 ( \17683 , \17682 , \1085 );
nand \U$17341 ( \17684 , \17680 , \17683 );
not \U$17342 ( \17685 , \17684 );
or \U$17343 ( \17686 , \17677 , \17685 );
nand \U$17344 ( \17687 , \16840 , \1089 );
nand \U$17345 ( \17688 , \17686 , \17687 );
not \U$17346 ( \17689 , \17688 );
or \U$17347 ( \17690 , \17676 , \17689 );
not \U$17348 ( \17691 , \17688 );
not \U$17349 ( \17692 , \17691 );
not \U$17350 ( \17693 , \17674 );
or \U$17351 ( \17694 , \17692 , \17693 );
not \U$17352 ( \17695 , \1570 );
not \U$17353 ( \17696 , RIbb2f250_9);
not \U$17354 ( \17697 , \13475 );
or \U$17355 ( \17698 , \17696 , \17697 );
nand \U$17356 ( \17699 , \13212 , \1566 );
nand \U$17357 ( \17700 , \17698 , \17699 );
not \U$17358 ( \17701 , \17700 );
or \U$17359 ( \17702 , \17695 , \17701 );
nand \U$17360 ( \17703 , \17319 , \1533 );
nand \U$17361 ( \17704 , \17702 , \17703 );
nand \U$17362 ( \17705 , \17694 , \17704 );
nand \U$17363 ( \17706 , \17690 , \17705 );
xor \U$17364 ( \17707 , \17662 , \17706 );
not \U$17365 ( \17708 , \3887 );
not \U$17366 ( \17709 , \16797 );
or \U$17367 ( \17710 , \17708 , \17709 );
not \U$17368 ( \17711 , RIbb2e710_33);
not \U$17369 ( \17712 , \13904 );
or \U$17370 ( \17713 , \17711 , \17712 );
nand \U$17371 ( \17714 , \3228 , \2935 );
nand \U$17372 ( \17715 , \17713 , \17714 );
nand \U$17373 ( \17716 , \17715 , \4791 );
nand \U$17374 ( \17717 , \17710 , \17716 );
xor \U$17375 ( \17718 , \17707 , \17717 );
and \U$17376 ( \17719 , \17658 , \17718 );
not \U$17377 ( \17720 , \17658 );
not \U$17378 ( \17721 , \17718 );
and \U$17379 ( \17722 , \17720 , \17721 );
nor \U$17380 ( \17723 , \17719 , \17722 );
xor \U$17381 ( \17724 , \16760 , \16790 );
and \U$17382 ( \17725 , \17724 , \16807 );
and \U$17383 ( \17726 , \16760 , \16790 );
or \U$17384 ( \17727 , \17725 , \17726 );
not \U$17385 ( \17728 , \17147 );
not \U$17386 ( \17729 , \17152 );
or \U$17387 ( \17730 , \17728 , \17729 );
nand \U$17388 ( \17731 , \17141 , \17150 );
nand \U$17389 ( \17732 , \17730 , \17731 );
xor \U$17390 ( \17733 , \17164 , \17732 );
xor \U$17391 ( \17734 , \17727 , \17733 );
xor \U$17392 ( \17735 , \17225 , \17215 );
xor \U$17393 ( \17736 , \17735 , \17237 );
xor \U$17394 ( \17737 , \17734 , \17736 );
xor \U$17395 ( \17738 , \17723 , \17737 );
xor \U$17396 ( \17739 , \17328 , \17338 );
and \U$17397 ( \17740 , \17739 , \17349 );
and \U$17398 ( \17741 , \17328 , \17338 );
or \U$17399 ( \17742 , \17740 , \17741 );
not \U$17400 ( \17743 , \1312 );
not \U$17401 ( \17744 , \17516 );
buf \U$17402 ( \17745 , \17744 );
nor \U$17403 ( \17746 , \17743 , \17745 );
not \U$17404 ( \17747 , \17534 );
not \U$17405 ( \17748 , \1428 );
or \U$17406 ( \17749 , \17747 , \17748 );
not \U$17407 ( \17750 , \16703 );
not \U$17408 ( \17751 , \17750 );
not \U$17409 ( \17752 , \17751 );
not \U$17410 ( \17753 , \13990 );
or \U$17411 ( \17754 , \17752 , \17753 );
not \U$17412 ( \17755 , \16703 );
buf \U$17413 ( \17756 , \17755 );
nand \U$17414 ( \17757 , \17523 , \17756 );
nand \U$17415 ( \17758 , \17754 , \17757 );
nand \U$17416 ( \17759 , \1375 , \17758 );
nand \U$17417 ( \17760 , \17749 , \17759 );
xor \U$17418 ( \17761 , \17746 , \17760 );
not \U$17419 ( \17762 , \1261 );
not \U$17420 ( \17763 , \16831 );
or \U$17421 ( \17764 , \17762 , \17763 );
not \U$17422 ( \17765 , \16556 );
not \U$17423 ( \17766 , \1243 );
or \U$17424 ( \17767 , \17765 , \17766 );
not \U$17425 ( \17768 , \16706 );
nand \U$17426 ( \17769 , \1288 , \17768 );
nand \U$17427 ( \17770 , \17767 , \17769 );
nand \U$17428 ( \17771 , \1264 , \17770 );
nand \U$17429 ( \17772 , \17764 , \17771 );
and \U$17430 ( \17773 , \17761 , \17772 );
and \U$17431 ( \17774 , \17746 , \17760 );
or \U$17432 ( \17775 , \17773 , \17774 );
not \U$17433 ( \17776 , \17758 );
not \U$17434 ( \17777 , \1428 );
or \U$17435 ( \17778 , \17776 , \17777 );
nand \U$17436 ( \17779 , \1375 , \16712 );
nand \U$17437 ( \17780 , \17778 , \17779 );
nor \U$17438 ( \17781 , \17780 , \17262 );
not \U$17439 ( \17782 , \17781 );
nand \U$17440 ( \17783 , \17780 , \17262 );
nand \U$17441 ( \17784 , \17782 , \17783 );
xor \U$17442 ( \17785 , \17775 , \17784 );
not \U$17443 ( \17786 , \2925 );
not \U$17444 ( \17787 , \16155 );
or \U$17445 ( \17788 , \17786 , \17787 );
not \U$17446 ( \17789 , RIbb2e8f0_29);
not \U$17447 ( \17790 , \4392 );
or \U$17448 ( \17791 , \17789 , \17790 );
nand \U$17449 ( \17792 , \8375 , \2949 );
nand \U$17450 ( \17793 , \17791 , \17792 );
nand \U$17451 ( \17794 , \17793 , \2922 );
nand \U$17452 ( \17795 , \17788 , \17794 );
and \U$17453 ( \17796 , \17785 , \17795 );
and \U$17454 ( \17797 , \17775 , \17784 );
or \U$17455 ( \17798 , \17796 , \17797 );
xor \U$17456 ( \17799 , \17742 , \17798 );
not \U$17457 ( \17800 , \3383 );
not \U$17458 ( \17801 , RIbb2ebc0_23);
not \U$17459 ( \17802 , \6938 );
or \U$17460 ( \17803 , \17801 , \17802 );
nand \U$17461 ( \17804 , \11534 , \2073 );
nand \U$17462 ( \17805 , \17803 , \17804 );
not \U$17463 ( \17806 , \17805 );
or \U$17464 ( \17807 , \17800 , \17806 );
not \U$17465 ( \17808 , RIbb2ebc0_23);
not \U$17466 ( \17809 , \13853 );
or \U$17467 ( \17810 , \17808 , \17809 );
not \U$17468 ( \17811 , \7296 );
not \U$17469 ( \17812 , \17811 );
nand \U$17470 ( \17813 , \17812 , \3388 );
nand \U$17471 ( \17814 , \17810 , \17813 );
nand \U$17472 ( \17815 , \17814 , \3406 );
nand \U$17473 ( \17816 , \17807 , \17815 );
not \U$17474 ( \17817 , \17816 );
not \U$17475 ( \17818 , \2078 );
not \U$17476 ( \17819 , RIbb2ecb0_21);
not \U$17477 ( \17820 , \12210 );
or \U$17478 ( \17821 , \17819 , \17820 );
nand \U$17479 ( \17822 , \9818 , \849 );
nand \U$17480 ( \17823 , \17821 , \17822 );
not \U$17481 ( \17824 , \17823 );
or \U$17482 ( \17825 , \17818 , \17824 );
not \U$17483 ( \17826 , RIbb2ecb0_21);
not \U$17484 ( \17827 , \15786 );
or \U$17485 ( \17828 , \17826 , \17827 );
nand \U$17486 ( \17829 , \8630 , \2249 );
nand \U$17487 ( \17830 , \17828 , \17829 );
nand \U$17488 ( \17831 , \17830 , \2077 );
nand \U$17489 ( \17832 , \17825 , \17831 );
not \U$17490 ( \17833 , \17832 );
or \U$17491 ( \17834 , \17817 , \17833 );
not \U$17492 ( \17835 , \17832 );
not \U$17493 ( \17836 , \17835 );
not \U$17494 ( \17837 , \17816 );
not \U$17495 ( \17838 , \17837 );
or \U$17496 ( \17839 , \17836 , \17838 );
not \U$17497 ( \17840 , \16345 );
not \U$17498 ( \17841 , \2963 );
or \U$17499 ( \17842 , \17840 , \17841 );
and \U$17500 ( \17843 , RIbb2ead0_25, \15797 );
not \U$17501 ( \17844 , RIbb2ead0_25);
and \U$17502 ( \17845 , \17844 , \6604 );
or \U$17503 ( \17846 , \17843 , \17845 );
nand \U$17504 ( \17847 , \17846 , \2980 );
nand \U$17505 ( \17848 , \17842 , \17847 );
nand \U$17506 ( \17849 , \17839 , \17848 );
nand \U$17507 ( \17850 , \17834 , \17849 );
xor \U$17508 ( \17851 , \17799 , \17850 );
not \U$17509 ( \17852 , \17688 );
not \U$17510 ( \17853 , \17674 );
or \U$17511 ( \17854 , \17852 , \17853 );
nand \U$17512 ( \17855 , \17675 , \17691 );
nand \U$17513 ( \17856 , \17854 , \17855 );
xor \U$17514 ( \17857 , \17856 , \17704 );
not \U$17515 ( \17858 , \1445 );
and \U$17516 ( \17859 , RIbb2ef80_15, \14886 );
not \U$17517 ( \17860 , RIbb2ef80_15);
and \U$17518 ( \17861 , \17860 , \11581 );
or \U$17519 ( \17862 , \17859 , \17861 );
not \U$17520 ( \17863 , \17862 );
or \U$17521 ( \17864 , \17858 , \17863 );
and \U$17522 ( \17865 , RIbb2ef80_15, \15188 );
not \U$17523 ( \17866 , RIbb2ef80_15);
and \U$17524 ( \17867 , \17866 , \11144 );
or \U$17525 ( \17868 , \17865 , \17867 );
nand \U$17526 ( \17869 , \17868 , \1517 );
nand \U$17527 ( \17870 , \17864 , \17869 );
not \U$17528 ( \17871 , \17870 );
not \U$17529 ( \17872 , \853 );
not \U$17530 ( \17873 , RIbb2eda0_19);
not \U$17531 ( \17874 , \10306 );
or \U$17532 ( \17875 , \17873 , \17874 );
nand \U$17533 ( \17876 , \9841 , \1776 );
nand \U$17534 ( \17877 , \17875 , \17876 );
not \U$17535 ( \17878 , \17877 );
or \U$17536 ( \17879 , \17872 , \17878 );
not \U$17537 ( \17880 , RIbb2eda0_19);
not \U$17538 ( \17881 , \13916 );
or \U$17539 ( \17882 , \17880 , \17881 );
nand \U$17540 ( \17883 , \16475 , \3251 );
nand \U$17541 ( \17884 , \17882 , \17883 );
nand \U$17542 ( \17885 , \17884 , \855 );
nand \U$17543 ( \17886 , \17879 , \17885 );
not \U$17544 ( \17887 , \17886 );
nand \U$17545 ( \17888 , \17871 , \17887 );
not \U$17546 ( \17889 , \17888 );
not \U$17547 ( \17890 , \832 );
not \U$17548 ( \17891 , \17306 );
or \U$17549 ( \17892 , \17890 , \17891 );
not \U$17550 ( \17893 , RIbb2ee90_17);
not \U$17551 ( \17894 , \12230 );
or \U$17552 ( \17895 , \17893 , \17894 );
not \U$17553 ( \17896 , \15105 );
nand \U$17554 ( \17897 , \17896 , \816 );
nand \U$17555 ( \17898 , \17895 , \17897 );
nand \U$17556 ( \17899 , \17898 , \836 );
nand \U$17557 ( \17900 , \17892 , \17899 );
not \U$17558 ( \17901 , \17900 );
or \U$17559 ( \17902 , \17889 , \17901 );
nand \U$17560 ( \17903 , \17886 , \17870 );
nand \U$17561 ( \17904 , \17902 , \17903 );
xor \U$17562 ( \17905 , \17857 , \17904 );
not \U$17563 ( \17906 , \3887 );
not \U$17564 ( \17907 , RIbb2e710_33);
not \U$17565 ( \17908 , \3045 );
or \U$17566 ( \17909 , \17907 , \17908 );
not \U$17567 ( \17910 , \3044 );
not \U$17568 ( \17911 , \17910 );
nand \U$17569 ( \17912 , \17911 , \13352 );
nand \U$17570 ( \17913 , \17909 , \17912 );
not \U$17571 ( \17914 , \17913 );
or \U$17572 ( \17915 , \17906 , \17914 );
not \U$17573 ( \17916 , \3871 );
nand \U$17574 ( \17917 , \17916 , \16805 );
nand \U$17575 ( \17918 , \17915 , \17917 );
not \U$17576 ( \17919 , \17918 );
not \U$17577 ( \17920 , \17919 );
not \U$17578 ( \17921 , \2940 );
not \U$17579 ( \17922 , RIbb2e800_31);
not \U$17580 ( \17923 , \4752 );
or \U$17581 ( \17924 , \17922 , \17923 );
nand \U$17582 ( \17925 , \3089 , \9169 );
nand \U$17583 ( \17926 , \17924 , \17925 );
not \U$17584 ( \17927 , \17926 );
or \U$17585 ( \17928 , \17921 , \17927 );
not \U$17586 ( \17929 , RIbb2e800_31);
not \U$17587 ( \17930 , \13731 );
or \U$17588 ( \17931 , \17929 , \17930 );
nand \U$17589 ( \17932 , \17931 , \16191 );
nand \U$17590 ( \17933 , \17932 , \3613 );
nand \U$17591 ( \17934 , \17928 , \17933 );
not \U$17592 ( \17935 , \17934 );
not \U$17593 ( \17936 , \17935 );
or \U$17594 ( \17937 , \17920 , \17936 );
not \U$17595 ( \17938 , \12167 );
not \U$17596 ( \17939 , RIbb2df90_49);
not \U$17597 ( \17940 , \3066 );
or \U$17598 ( \17941 , \17939 , \17940 );
nand \U$17599 ( \17942 , \3067 , \12278 );
nand \U$17600 ( \17943 , \17941 , \17942 );
not \U$17601 ( \17944 , \17943 );
or \U$17602 ( \17945 , \17938 , \17944 );
nand \U$17603 ( \17946 , \16418 , \16427 );
nand \U$17604 ( \17947 , \17945 , \17946 );
nand \U$17605 ( \17948 , \17937 , \17947 );
nand \U$17606 ( \17949 , \17934 , \17918 );
nand \U$17607 ( \17950 , \17948 , \17949 );
xor \U$17608 ( \17951 , \17905 , \17950 );
xor \U$17609 ( \17952 , \17851 , \17951 );
not \U$17610 ( \17953 , \15181 );
not \U$17611 ( \17954 , \16361 );
or \U$17612 ( \17955 , \17953 , \17954 );
not \U$17613 ( \17956 , RIbb2dcc0_55);
not \U$17614 ( \17957 , \5003 );
or \U$17615 ( \17958 , \17956 , \17957 );
not \U$17616 ( \17959 , RIbb2dcc0_55);
nand \U$17617 ( \17960 , \1548 , \17959 );
nand \U$17618 ( \17961 , \17958 , \17960 );
nand \U$17619 ( \17962 , \17961 , \14613 );
nand \U$17620 ( \17963 , \17955 , \17962 );
not \U$17621 ( \17964 , \10119 );
not \U$17622 ( \17965 , \16388 );
or \U$17623 ( \17966 , \17964 , \17965 );
not \U$17624 ( \17967 , RIbb2e170_45);
not \U$17625 ( \17968 , \13358 );
or \U$17626 ( \17969 , \17967 , \17968 );
not \U$17627 ( \17970 , RIbb2e170_45);
nand \U$17628 ( \17971 , \6096 , \17970 );
nand \U$17629 ( \17972 , \17969 , \17971 );
nand \U$17630 ( \17973 , \17972 , \10117 );
nand \U$17631 ( \17974 , \17966 , \17973 );
xor \U$17632 ( \17975 , \17963 , \17974 );
not \U$17633 ( \17976 , \10451 );
not \U$17634 ( \17977 , \16373 );
or \U$17635 ( \17978 , \17976 , \17977 );
nand \U$17636 ( \17979 , \17490 , \9098 );
nand \U$17637 ( \17980 , \17978 , \17979 );
and \U$17638 ( \17981 , \17975 , \17980 );
and \U$17639 ( \17982 , \17963 , \17974 );
or \U$17640 ( \17983 , \17981 , \17982 );
not \U$17641 ( \17984 , \3613 );
not \U$17642 ( \17985 , \17926 );
or \U$17643 ( \17986 , \17984 , \17985 );
not \U$17644 ( \17987 , RIbb2e800_31);
not \U$17645 ( \17988 , \13552 );
or \U$17646 ( \17989 , \17987 , \17988 );
nand \U$17647 ( \17990 , \13551 , \9169 );
nand \U$17648 ( \17991 , \17989 , \17990 );
nand \U$17649 ( \17992 , \17991 , \2939 );
nand \U$17650 ( \17993 , \17986 , \17992 );
not \U$17651 ( \17994 , \4075 );
not \U$17652 ( \17995 , \17913 );
or \U$17653 ( \17996 , \17994 , \17995 );
nand \U$17654 ( \17997 , \3887 , \17430 );
nand \U$17655 ( \17998 , \17996 , \17997 );
xor \U$17656 ( \17999 , \17993 , \17998 );
not \U$17657 ( \18000 , \12285 );
not \U$17658 ( \18001 , \17943 );
or \U$17659 ( \18002 , \18000 , \18001 );
nand \U$17660 ( \18003 , \17364 , \12167 );
nand \U$17661 ( \18004 , \18002 , \18003 );
and \U$17662 ( \18005 , \17999 , \18004 );
and \U$17663 ( \18006 , \17993 , \17998 );
or \U$17664 ( \18007 , \18005 , \18006 );
nor \U$17665 ( \18008 , \17983 , \18007 );
not \U$17666 ( \18009 , \8354 );
not \U$17667 ( \18010 , RIbb2e350_41);
not \U$17668 ( \18011 , \13286 );
or \U$17669 ( \18012 , \18010 , \18011 );
nand \U$17670 ( \18013 , \2222 , \9402 );
nand \U$17671 ( \18014 , \18012 , \18013 );
not \U$17672 ( \18015 , \18014 );
or \U$17673 ( \18016 , \18009 , \18015 );
nand \U$17674 ( \18017 , \17466 , \8361 );
nand \U$17675 ( \18018 , \18016 , \18017 );
not \U$17676 ( \18019 , \16271 );
not \U$17677 ( \18020 , \17476 );
or \U$17678 ( \18021 , \18019 , \18020 );
and \U$17679 ( \18022 , RIbb2dae0_59, \14734 );
not \U$17680 ( \18023 , RIbb2dae0_59);
and \U$17681 ( \18024 , \18023 , \3450 );
or \U$17682 ( \18025 , \18022 , \18024 );
nand \U$17683 ( \18026 , \18025 , \16257 );
nand \U$17684 ( \18027 , \18021 , \18026 );
or \U$17685 ( \18028 , \18018 , \18027 );
not \U$17686 ( \18029 , \14920 );
not \U$17687 ( \18030 , \17554 );
or \U$17688 ( \18031 , \18029 , \18030 );
not \U$17689 ( \18032 , RIbb2ddb0_53);
not \U$17690 ( \18033 , \14819 );
or \U$17691 ( \18034 , \18032 , \18033 );
nand \U$17692 ( \18035 , \3484 , \13463 );
nand \U$17693 ( \18036 , \18034 , \18035 );
nand \U$17694 ( \18037 , \18036 , \14929 );
nand \U$17695 ( \18038 , \18031 , \18037 );
nand \U$17696 ( \18039 , \18028 , \18038 );
nand \U$17697 ( \18040 , \18018 , \18027 );
and \U$17698 ( \18041 , \18039 , \18040 );
or \U$17699 ( \18042 , \18008 , \18041 );
nand \U$17700 ( \18043 , \17983 , \18007 );
nand \U$17701 ( \18044 , \18042 , \18043 );
and \U$17702 ( \18045 , \17952 , \18044 );
and \U$17703 ( \18046 , \17851 , \17951 );
or \U$17704 ( \18047 , \18045 , \18046 );
xor \U$17705 ( \18048 , \17738 , \18047 );
and \U$17706 ( \18049 , \17647 , \18048 );
and \U$17707 ( \18050 , \17249 , \17646 );
or \U$17708 ( \18051 , \18049 , \18050 );
xor \U$17709 ( \18052 , \17247 , \18051 );
xor \U$17710 ( \18053 , \16545 , \16557 );
and \U$17711 ( \18054 , \18053 , \16583 );
and \U$17712 ( \18055 , \16545 , \16557 );
or \U$17713 ( \18056 , \18054 , \18055 );
not \U$17714 ( \18057 , \3383 );
not \U$17715 ( \18058 , RIbb2ebc0_23);
not \U$17716 ( \18059 , \10126 );
or \U$17717 ( \18060 , \18058 , \18059 );
nand \U$17718 ( \18061 , \8387 , \3396 );
nand \U$17719 ( \18062 , \18060 , \18061 );
not \U$17720 ( \18063 , \18062 );
or \U$17721 ( \18064 , \18057 , \18063 );
nand \U$17722 ( \18065 , \16954 , \3406 );
nand \U$17723 ( \18066 , \18064 , \18065 );
xor \U$17724 ( \18067 , \18056 , \18066 );
not \U$17725 ( \18068 , \2963 );
not \U$17726 ( \18069 , RIbb2ead0_25);
not \U$17727 ( \18070 , \4393 );
or \U$17728 ( \18071 , \18069 , \18070 );
not \U$17729 ( \18072 , RIbb2ead0_25);
nand \U$17730 ( \18073 , \18072 , \6269 );
nand \U$17731 ( \18074 , \18071 , \18073 );
not \U$17732 ( \18075 , \18074 );
or \U$17733 ( \18076 , \18068 , \18075 );
nand \U$17734 ( \18077 , \16933 , \2980 );
nand \U$17735 ( \18078 , \18076 , \18077 );
xor \U$17736 ( \18079 , \18067 , \18078 );
not \U$17737 ( \18080 , \17002 );
not \U$17738 ( \18081 , \16981 );
or \U$17739 ( \18082 , \18080 , \18081 );
or \U$17740 ( \18083 , \16981 , \17002 );
nand \U$17741 ( \18084 , \18083 , \16991 );
nand \U$17742 ( \18085 , \18082 , \18084 );
xor \U$17743 ( \18086 , \18079 , \18085 );
not \U$17744 ( \18087 , \16730 );
not \U$17745 ( \18088 , \1428 );
or \U$17746 ( \18089 , \18087 , \18088 );
not \U$17747 ( \18090 , \1312 );
not \U$17748 ( \18091 , \16747 );
or \U$17749 ( \18092 , \18090 , \18091 );
not \U$17750 ( \18093 , \16748 );
nand \U$17751 ( \18094 , \18093 , \13990 );
nand \U$17752 ( \18095 , \18092 , \18094 );
nand \U$17753 ( \18096 , \18095 , \1375 );
nand \U$17754 ( \18097 , \18089 , \18096 );
xor \U$17755 ( \18098 , \18097 , \16758 );
not \U$17756 ( \18099 , \1570 );
not \U$17757 ( \18100 , RIbb2f250_9);
not \U$17758 ( \18101 , \12348 );
or \U$17759 ( \18102 , \18100 , \18101 );
nand \U$17760 ( \18103 , \14839 , \1566 );
nand \U$17761 ( \18104 , \18102 , \18103 );
not \U$17762 ( \18105 , \18104 );
or \U$17763 ( \18106 , \18099 , \18105 );
nand \U$17764 ( \18107 , \17700 , \1533 );
nand \U$17765 ( \18108 , \18106 , \18107 );
and \U$17766 ( \18109 , \18098 , \18108 );
and \U$17767 ( \18110 , \18097 , \16758 );
or \U$17768 ( \18111 , \18109 , \18110 );
not \U$17769 ( \18112 , \12965 );
not \U$17770 ( \18113 , RIbb2e080_47);
not \U$17771 ( \18114 , \3238 );
or \U$17772 ( \18115 , \18113 , \18114 );
nand \U$17773 ( \18116 , \3243 , \16171 );
nand \U$17774 ( \18117 , \18115 , \18116 );
not \U$17775 ( \18118 , \18117 );
or \U$17776 ( \18119 , \18112 , \18118 );
nand \U$17777 ( \18120 , \17173 , \11176 );
nand \U$17778 ( \18121 , \18119 , \18120 );
xor \U$17779 ( \18122 , \18111 , \18121 );
not \U$17780 ( \18123 , \2940 );
not \U$17781 ( \18124 , \17199 );
or \U$17782 ( \18125 , \18123 , \18124 );
not \U$17783 ( \18126 , RIbb2e800_31);
not \U$17784 ( \18127 , \3655 );
or \U$17785 ( \18128 , \18126 , \18127 );
nand \U$17786 ( \18129 , \3762 , \11975 );
nand \U$17787 ( \18130 , \18128 , \18129 );
nand \U$17788 ( \18131 , \18130 , \2941 );
nand \U$17789 ( \18132 , \18125 , \18131 );
xor \U$17790 ( \18133 , \18122 , \18132 );
xnor \U$17791 ( \18134 , \18086 , \18133 );
not \U$17792 ( \18135 , \18134 );
not \U$17793 ( \18136 , \17649 );
not \U$17794 ( \18137 , \17654 );
or \U$17795 ( \18138 , \18136 , \18137 );
or \U$17796 ( \18139 , \17654 , \17649 );
nand \U$17797 ( \18140 , \18139 , \17718 );
nand \U$17798 ( \18141 , \18138 , \18140 );
not \U$17799 ( \18142 , \18141 );
or \U$17800 ( \18143 , \18135 , \18142 );
or \U$17801 ( \18144 , \18134 , \18141 );
nand \U$17802 ( \18145 , \18143 , \18144 );
xor \U$17803 ( \18146 , \17727 , \17733 );
and \U$17804 ( \18147 , \18146 , \17736 );
and \U$17805 ( \18148 , \17727 , \17733 );
or \U$17806 ( \18149 , \18147 , \18148 );
and \U$17807 ( \18150 , \18145 , \18149 );
not \U$17808 ( \18151 , \18145 );
not \U$17809 ( \18152 , \18149 );
and \U$17810 ( \18153 , \18151 , \18152 );
nor \U$17811 ( \18154 , \18150 , \18153 );
xor \U$17812 ( \18155 , \17662 , \17706 );
and \U$17813 ( \18156 , \18155 , \17717 );
and \U$17814 ( \18157 , \17662 , \17706 );
or \U$17815 ( \18158 , \18156 , \18157 );
not \U$17816 ( \18159 , \7104 );
not \U$17817 ( \18160 , \4610 );
not \U$17818 ( \18161 , \10908 );
and \U$17819 ( \18162 , \18160 , \18161 );
and \U$17820 ( \18163 , \3810 , \10908 );
nor \U$17821 ( \18164 , \18162 , \18163 );
nor \U$17822 ( \18165 , \18159 , \18164 );
not \U$17823 ( \18166 , \7103 );
nor \U$17824 ( \18167 , \18166 , \17118 );
nor \U$17825 ( \18168 , \18165 , \18167 );
not \U$17826 ( \18169 , \18168 );
not \U$17827 ( \18170 , \15181 );
not \U$17828 ( \18171 , RIbb2dcc0_55);
not \U$17829 ( \18172 , \14734 );
or \U$17830 ( \18173 , \18171 , \18172 );
not \U$17831 ( \18174 , RIbb2dcc0_55);
nand \U$17832 ( \18175 , \3450 , \18174 );
nand \U$17833 ( \18176 , \18173 , \18175 );
not \U$17834 ( \18177 , \18176 );
or \U$17835 ( \18178 , \18170 , \18177 );
nand \U$17836 ( \18179 , \17139 , \14613 );
nand \U$17837 ( \18180 , \18178 , \18179 );
not \U$17838 ( \18181 , \6241 );
and \U$17839 ( \18182 , \13286 , RIbb2e530_37);
not \U$17840 ( \18183 , \13286 );
and \U$17841 ( \18184 , \18183 , \4708 );
or \U$17842 ( \18185 , \18182 , \18184 );
not \U$17843 ( \18186 , \18185 );
or \U$17844 ( \18187 , \18181 , \18186 );
not \U$17845 ( \18188 , \6252 );
nand \U$17846 ( \18189 , \18188 , \17000 );
nand \U$17847 ( \18190 , \18187 , \18189 );
and \U$17848 ( \18191 , \18180 , \18190 );
not \U$17849 ( \18192 , \18180 );
not \U$17850 ( \18193 , \18190 );
and \U$17851 ( \18194 , \18192 , \18193 );
nor \U$17852 ( \18195 , \18191 , \18194 );
not \U$17853 ( \18196 , \18195 );
or \U$17854 ( \18197 , \18169 , \18196 );
or \U$17855 ( \18198 , \18168 , \18195 );
nand \U$17856 ( \18199 , \18197 , \18198 );
xor \U$17857 ( \18200 , \18158 , \18199 );
not \U$17858 ( \18201 , \14067 );
not \U$17859 ( \18202 , \17109 );
or \U$17860 ( \18203 , \18201 , \18202 );
not \U$17861 ( \18204 , \1037 );
and \U$17862 ( \18205 , RIbb2dea0_51, \18204 );
not \U$17863 ( \18206 , RIbb2dea0_51);
and \U$17864 ( \18207 , \18206 , \1037 );
or \U$17865 ( \18208 , \18205 , \18207 );
nand \U$17866 ( \18209 , \18208 , \12692 );
nand \U$17867 ( \18210 , \18203 , \18209 );
not \U$17868 ( \18211 , \14930 );
not \U$17869 ( \18212 , RIbb2ddb0_53);
not \U$17870 ( \18213 , \951 );
or \U$17871 ( \18214 , \18212 , \18213 );
nand \U$17872 ( \18215 , \956 , \13941 );
nand \U$17873 ( \18216 , \18214 , \18215 );
not \U$17874 ( \18217 , \18216 );
or \U$17875 ( \18218 , \18211 , \18217 );
nand \U$17876 ( \18219 , \17221 , \17562 );
nand \U$17877 ( \18220 , \18218 , \18219 );
xor \U$17878 ( \18221 , \18210 , \18220 );
not \U$17879 ( \18222 , \8354 );
and \U$17880 ( \18223 , \17386 , RIbb2e350_41);
not \U$17881 ( \18224 , \17386 );
and \U$17882 ( \18225 , \18224 , \7097 );
or \U$17883 ( \18226 , \18223 , \18225 );
not \U$17884 ( \18227 , \18226 );
or \U$17885 ( \18228 , \18222 , \18227 );
nand \U$17886 ( \18229 , \17211 , \8362 );
nand \U$17887 ( \18230 , \18228 , \18229 );
xor \U$17888 ( \18231 , \18221 , \18230 );
xor \U$17889 ( \18232 , \18200 , \18231 );
not \U$17890 ( \18233 , \1077 );
not \U$17891 ( \18234 , RIbb2f160_11);
not \U$17892 ( \18235 , \11580 );
or \U$17893 ( \18236 , \18234 , \18235 );
nand \U$17894 ( \18237 , \14885 , \1048 );
nand \U$17895 ( \18238 , \18236 , \18237 );
not \U$17896 ( \18239 , \18238 );
or \U$17897 ( \18240 , \18233 , \18239 );
not \U$17898 ( \18241 , RIbb2f160_11);
not \U$17899 ( \18242 , \12839 );
or \U$17900 ( \18243 , \18241 , \18242 );
nand \U$17901 ( \18244 , \12175 , \1805 );
nand \U$17902 ( \18245 , \18243 , \18244 );
nand \U$17903 ( \18246 , \18245 , \1011 );
nand \U$17904 ( \18247 , \18240 , \18246 );
not \U$17905 ( \18248 , \2922 );
not \U$17906 ( \18249 , \17183 );
or \U$17907 ( \18250 , \18248 , \18249 );
not \U$17908 ( \18251 , RIbb2e8f0_29);
not \U$17909 ( \18252 , \3045 );
or \U$17910 ( \18253 , \18251 , \18252 );
nand \U$17911 ( \18254 , \16185 , \3440 );
nand \U$17912 ( \18255 , \18253 , \18254 );
nand \U$17913 ( \18256 , \18255 , \2925 );
nand \U$17914 ( \18257 , \18250 , \18256 );
xor \U$17915 ( \18258 , \18247 , \18257 );
not \U$17916 ( \18259 , \10599 );
not \U$17917 ( \18260 , \17160 );
or \U$17918 ( \18261 , \18259 , \18260 );
not \U$17919 ( \18262 , RIbb2e170_45);
not \U$17920 ( \18263 , \3066 );
or \U$17921 ( \18264 , \18262 , \18263 );
nand \U$17922 ( \18265 , \4006 , \9094 );
nand \U$17923 ( \18266 , \18264 , \18265 );
nand \U$17924 ( \18267 , \18266 , \10119 );
nand \U$17925 ( \18268 , \18261 , \18267 );
xor \U$17926 ( \18269 , \18258 , \18268 );
not \U$17927 ( \18270 , \5845 );
not \U$17928 ( \18271 , RIbb2e620_35);
not \U$17929 ( \18272 , \3952 );
or \U$17930 ( \18273 , \18271 , \18272 );
nand \U$17931 ( \18274 , \3951 , \6002 );
nand \U$17932 ( \18275 , \18273 , \18274 );
not \U$17933 ( \18276 , \18275 );
or \U$17934 ( \18277 , \18270 , \18276 );
nand \U$17935 ( \18278 , \16975 , \4712 );
nand \U$17936 ( \18279 , \18277 , \18278 );
not \U$17937 ( \18280 , \13295 );
not \U$17938 ( \18281 , \16987 );
or \U$17939 ( \18282 , \18280 , \18281 );
not \U$17940 ( \18283 , RIbb2df90_49);
not \U$17941 ( \18284 , \3479 );
or \U$17942 ( \18285 , \18283 , \18284 );
nand \U$17943 ( \18286 , \3480 , \12278 );
nand \U$17944 ( \18287 , \18285 , \18286 );
nand \U$17945 ( \18288 , \18287 , \12285 );
nand \U$17946 ( \18289 , \18282 , \18288 );
xor \U$17947 ( \18290 , \18279 , \18289 );
not \U$17948 ( \18291 , \4791 );
not \U$17949 ( \18292 , \16400 );
not \U$17950 ( \18293 , \3877 );
and \U$17951 ( \18294 , \18292 , \18293 );
not \U$17952 ( \18295 , RIbb2e710_33);
and \U$17953 ( \18296 , \3202 , \18295 );
nor \U$17954 ( \18297 , \18294 , \18296 );
not \U$17955 ( \18298 , \18297 );
not \U$17956 ( \18299 , \18298 );
or \U$17957 ( \18300 , \18291 , \18299 );
nand \U$17958 ( \18301 , \17715 , \3887 );
nand \U$17959 ( \18302 , \18300 , \18301 );
xor \U$17960 ( \18303 , \18290 , \18302 );
xor \U$17961 ( \18304 , \18269 , \18303 );
not \U$17962 ( \18305 , \10449 );
not \U$17963 ( \18306 , \17233 );
or \U$17964 ( \18307 , \18305 , \18306 );
not \U$17965 ( \18308 , RIbb2e260_43);
not \U$17966 ( \18309 , \11054 );
or \U$17967 ( \18310 , \18308 , \18309 );
nand \U$17968 ( \18311 , \3109 , \17231 );
nand \U$17969 ( \18312 , \18310 , \18311 );
nand \U$17970 ( \18313 , \18312 , \9099 );
nand \U$17971 ( \18314 , \18307 , \18313 );
not \U$17972 ( \18315 , \17100 );
not \U$17973 ( \18316 , RIbb2dbd0_57);
not \U$17974 ( \18317 , \12969 );
or \U$17975 ( \18318 , \18316 , \18317 );
nand \U$17976 ( \18319 , \12970 , \15741 );
nand \U$17977 ( \18320 , \18318 , \18319 );
not \U$17978 ( \18321 , \18320 );
or \U$17979 ( \18322 , \18315 , \18321 );
nand \U$17980 ( \18323 , \17099 , \16675 );
nand \U$17981 ( \18324 , \18322 , \18323 );
not \U$17982 ( \18325 , \18324 );
and \U$17983 ( \18326 , \18314 , \18325 );
not \U$17984 ( \18327 , \18314 );
and \U$17985 ( \18328 , \18327 , \18324 );
or \U$17986 ( \18329 , \18326 , \18328 );
not \U$17987 ( \18330 , \3465 );
not \U$17988 ( \18331 , RIbb2e9e0_27);
not \U$17989 ( \18332 , \4748 );
or \U$17990 ( \18333 , \18331 , \18332 );
nand \U$17991 ( \18334 , \10458 , \3454 );
nand \U$17992 ( \18335 , \18333 , \18334 );
not \U$17993 ( \18336 , \18335 );
or \U$17994 ( \18337 , \18330 , \18336 );
nand \U$17995 ( \18338 , \16922 , \3445 );
nand \U$17996 ( \18339 , \18337 , \18338 );
and \U$17997 ( \18340 , \18329 , \18339 );
not \U$17998 ( \18341 , \18329 );
not \U$17999 ( \18342 , \18339 );
and \U$18000 ( \18343 , \18341 , \18342 );
nor \U$18001 ( \18344 , \18340 , \18343 );
xor \U$18002 ( \18345 , \18304 , \18344 );
xor \U$18003 ( \18346 , \18232 , \18345 );
xor \U$18004 ( \18347 , \18097 , \16758 );
xor \U$18005 ( \18348 , \18347 , \18108 );
not \U$18006 ( \18349 , \1089 );
not \U$18007 ( \18350 , \17684 );
or \U$18008 ( \18351 , \18349 , \18350 );
not \U$18009 ( \18352 , RIbb2f430_5);
not \U$18010 ( \18353 , \14526 );
not \U$18011 ( \18354 , \18353 );
or \U$18012 ( \18355 , \18352 , \18354 );
nand \U$18013 ( \18356 , \14527 , \1085 );
nand \U$18014 ( \18357 , \18355 , \18356 );
nand \U$18015 ( \18358 , \18357 , \1147 );
nand \U$18016 ( \18359 , \18351 , \18358 );
not \U$18017 ( \18360 , \1737 );
not \U$18018 ( \18361 , RIbb2f340_7);
not \U$18019 ( \18362 , \15054 );
or \U$18020 ( \18363 , \18361 , \18362 );
nand \U$18021 ( \18364 , \15055 , \2700 );
nand \U$18022 ( \18365 , \18363 , \18364 );
not \U$18023 ( \18366 , \18365 );
or \U$18024 ( \18367 , \18360 , \18366 );
nand \U$18025 ( \18368 , \16322 , \1702 );
nand \U$18026 ( \18369 , \18367 , \18368 );
xor \U$18027 ( \18370 , \18359 , \18369 );
not \U$18028 ( \18371 , \1077 );
not \U$18029 ( \18372 , \18245 );
or \U$18030 ( \18373 , \18371 , \18372 );
not \U$18031 ( \18374 , \17669 );
nand \U$18032 ( \18375 , \18374 , \1011 );
nand \U$18033 ( \18376 , \18373 , \18375 );
xor \U$18034 ( \18377 , \18370 , \18376 );
xor \U$18035 ( \18378 , \18348 , \18377 );
not \U$18036 ( \18379 , \998 );
not \U$18037 ( \18380 , \16613 );
or \U$18038 ( \18381 , \18379 , \18380 );
nand \U$18039 ( \18382 , \17334 , \916 );
nand \U$18040 ( \18383 , \18381 , \18382 );
not \U$18041 ( \18384 , \16541 );
not \U$18042 ( \18385 , RIbb2d9f0_61);
not \U$18043 ( \18386 , \813 );
or \U$18044 ( \18387 , \18385 , \18386 );
not \U$18045 ( \18388 , \812 );
nand \U$18046 ( \18389 , \18388 , \16537 );
nand \U$18047 ( \18390 , \18387 , \18389 );
not \U$18048 ( \18391 , \18390 );
or \U$18049 ( \18392 , \18384 , \18391 );
nand \U$18050 ( \18393 , \16533 , RIbb2d9f0_61);
nand \U$18051 ( \18394 , \18392 , \18393 );
xor \U$18052 ( \18395 , \18383 , \18394 );
not \U$18053 ( \18396 , \1445 );
not \U$18054 ( \18397 , \17868 );
or \U$18055 ( \18398 , \18396 , \18397 );
nand \U$18056 ( \18399 , \16595 , \1517 );
nand \U$18057 ( \18400 , \18398 , \18399 );
and \U$18058 ( \18401 , \18395 , \18400 );
and \U$18059 ( \18402 , \18383 , \18394 );
or \U$18060 ( \18403 , \18401 , \18402 );
and \U$18061 ( \18404 , \18378 , \18403 );
and \U$18062 ( \18405 , \18348 , \18377 );
or \U$18063 ( \18406 , \18404 , \18405 );
xor \U$18064 ( \18407 , \16324 , \16340 );
and \U$18065 ( \18408 , \18407 , \16355 );
and \U$18066 ( \18409 , \16324 , \16340 );
or \U$18067 ( \18410 , \18408 , \18409 );
not \U$18068 ( \18411 , \18410 );
not \U$18069 ( \18412 , \854 );
not \U$18070 ( \18413 , \16505 );
or \U$18071 ( \18414 , \18412 , \18413 );
nand \U$18072 ( \18415 , \17884 , \853 );
nand \U$18073 ( \18416 , \18414 , \18415 );
not \U$18074 ( \18417 , \18416 );
not \U$18075 ( \18418 , \2077 );
not \U$18076 ( \18419 , \17823 );
or \U$18077 ( \18420 , \18418 , \18419 );
nand \U$18078 ( \18421 , \16468 , \2078 );
nand \U$18079 ( \18422 , \18420 , \18421 );
not \U$18080 ( \18423 , \18422 );
or \U$18081 ( \18424 , \18417 , \18423 );
not \U$18082 ( \18425 , \18416 );
not \U$18083 ( \18426 , \18425 );
not \U$18084 ( \18427 , \18422 );
not \U$18085 ( \18428 , \18427 );
or \U$18086 ( \18429 , \18426 , \18428 );
not \U$18087 ( \18430 , \836 );
not \U$18088 ( \18431 , \16484 );
or \U$18089 ( \18432 , \18430 , \18431 );
nand \U$18090 ( \18433 , \17898 , \832 );
nand \U$18091 ( \18434 , \18432 , \18433 );
nand \U$18092 ( \18435 , \18429 , \18434 );
nand \U$18093 ( \18436 , \18424 , \18435 );
not \U$18094 ( \18437 , \18436 );
or \U$18095 ( \18438 , \18411 , \18437 );
or \U$18096 ( \18439 , \18436 , \18410 );
not \U$18097 ( \18440 , \17781 );
not \U$18098 ( \18441 , \18440 );
not \U$18099 ( \18442 , \3406 );
not \U$18100 ( \18443 , \17805 );
or \U$18101 ( \18444 , \18442 , \18443 );
nand \U$18102 ( \18445 , \16945 , \3383 );
nand \U$18103 ( \18446 , \18444 , \18445 );
not \U$18104 ( \18447 , \18446 );
or \U$18105 ( \18448 , \18441 , \18447 );
or \U$18106 ( \18449 , \18446 , \18440 );
xor \U$18107 ( \18450 , \16822 , \16833 );
and \U$18108 ( \18451 , \18450 , \16850 );
and \U$18109 ( \18452 , \16822 , \16833 );
or \U$18110 ( \18453 , \18451 , \18452 );
nand \U$18111 ( \18454 , \18449 , \18453 );
nand \U$18112 ( \18455 , \18448 , \18454 );
nand \U$18113 ( \18456 , \18439 , \18455 );
nand \U$18114 ( \18457 , \18438 , \18456 );
xor \U$18115 ( \18458 , \18406 , \18457 );
nor \U$18116 ( \18459 , \16249 , \16197 );
not \U$18117 ( \18460 , \16306 );
or \U$18118 ( \18461 , \18459 , \18460 );
nand \U$18119 ( \18462 , \16249 , \16197 );
nand \U$18120 ( \18463 , \18461 , \18462 );
xor \U$18121 ( \18464 , \18458 , \18463 );
xor \U$18122 ( \18465 , \18346 , \18464 );
not \U$18123 ( \18466 , \18465 );
and \U$18124 ( \18467 , \18154 , \18466 );
not \U$18125 ( \18468 , \18154 );
and \U$18126 ( \18469 , \18468 , \18465 );
nor \U$18127 ( \18470 , \18467 , \18469 );
not \U$18128 ( \18471 , \18470 );
xor \U$18129 ( \18472 , \17723 , \17737 );
and \U$18130 ( \18473 , \18472 , \18047 );
and \U$18131 ( \18474 , \17723 , \17737 );
or \U$18132 ( \18475 , \18473 , \18474 );
not \U$18133 ( \18476 , \18475 );
and \U$18134 ( \18477 , \18471 , \18476 );
and \U$18135 ( \18478 , \18470 , \18475 );
nor \U$18136 ( \18479 , \18477 , \18478 );
not \U$18137 ( \18480 , \18479 );
xor \U$18138 ( \18481 , \18052 , \18480 );
xor \U$18139 ( \18482 , \17261 , \17311 );
and \U$18140 ( \18483 , \18482 , \17350 );
and \U$18141 ( \18484 , \17261 , \17311 );
or \U$18142 ( \18485 , \18483 , \18484 );
not \U$18143 ( \18486 , \18485 );
and \U$18144 ( \18487 , \17848 , \17816 );
not \U$18145 ( \18488 , \17848 );
and \U$18146 ( \18489 , \18488 , \17837 );
nor \U$18147 ( \18490 , \18487 , \18489 );
and \U$18148 ( \18491 , \18490 , \17835 );
not \U$18149 ( \18492 , \18490 );
and \U$18150 ( \18493 , \18492 , \17832 );
nor \U$18151 ( \18494 , \18491 , \18493 );
not \U$18152 ( \18495 , \18494 );
xor \U$18153 ( \18496 , \17900 , \17887 );
xor \U$18154 ( \18497 , \18496 , \17870 );
not \U$18155 ( \18498 , \18497 );
or \U$18156 ( \18499 , \18495 , \18498 );
not \U$18157 ( \18500 , \8445 );
not \U$18158 ( \18501 , \17572 );
or \U$18159 ( \18502 , \18500 , \18501 );
and \U$18160 ( \18503 , RIbb2e440_39, \13414 );
not \U$18161 ( \18504 , RIbb2e440_39);
and \U$18162 ( \18505 , \18504 , \3951 );
or \U$18163 ( \18506 , \18503 , \18505 );
nand \U$18164 ( \18507 , \18506 , \8450 );
nand \U$18165 ( \18508 , \18502 , \18507 );
not \U$18166 ( \18509 , \14067 );
not \U$18167 ( \18510 , \17603 );
or \U$18168 ( \18511 , \18509 , \18510 );
and \U$18169 ( \18512 , RIbb2dea0_51, \3242 );
not \U$18170 ( \18513 , RIbb2dea0_51);
and \U$18171 ( \18514 , \18513 , \8856 );
or \U$18172 ( \18515 , \18512 , \18514 );
nand \U$18173 ( \18516 , \18515 , \12692 );
nand \U$18174 ( \18517 , \18511 , \18516 );
nor \U$18175 ( \18518 , \18508 , \18517 );
not \U$18176 ( \18519 , RIbb2e530_37);
not \U$18177 ( \18520 , \4638 );
or \U$18178 ( \18521 , \18519 , \18520 );
nand \U$18179 ( \18522 , \3202 , \4708 );
nand \U$18180 ( \18523 , \18521 , \18522 );
and \U$18181 ( \18524 , \6242 , \18523 );
and \U$18182 ( \18525 , \17589 , \6251 );
nor \U$18183 ( \18526 , \18524 , \18525 );
or \U$18184 ( \18527 , \18518 , \18526 );
nand \U$18185 ( \18528 , \18508 , \18517 );
nand \U$18186 ( \18529 , \18527 , \18528 );
nand \U$18187 ( \18530 , \18499 , \18529 );
not \U$18188 ( \18531 , \18497 );
not \U$18189 ( \18532 , \18494 );
nand \U$18190 ( \18533 , \18531 , \18532 );
nand \U$18191 ( \18534 , \18530 , \18533 );
not \U$18192 ( \18535 , \18534 );
or \U$18193 ( \18536 , \18486 , \18535 );
or \U$18194 ( \18537 , \18534 , \18485 );
not \U$18195 ( \18538 , \1570 );
not \U$18196 ( \18539 , \17326 );
or \U$18197 ( \18540 , \18538 , \18539 );
not \U$18198 ( \18541 , RIbb2f250_9);
not \U$18199 ( \18542 , \16309 );
or \U$18200 ( \18543 , \18541 , \18542 );
nand \U$18201 ( \18544 , \14526 , \1554 );
nand \U$18202 ( \18545 , \18543 , \18544 );
nand \U$18203 ( \18546 , \18545 , \1533 );
nand \U$18204 ( \18547 , \18540 , \18546 );
not \U$18205 ( \18548 , \1077 );
not \U$18206 ( \18549 , \16775 );
or \U$18207 ( \18550 , \18548 , \18549 );
not \U$18208 ( \18551 , RIbb2f160_11);
not \U$18209 ( \18552 , \13545 );
not \U$18210 ( \18553 , \18552 );
or \U$18211 ( \18554 , \18551 , \18553 );
nand \U$18212 ( \18555 , \13545 , \1805 );
nand \U$18213 ( \18556 , \18554 , \18555 );
nand \U$18214 ( \18557 , \18556 , \1011 );
nand \U$18215 ( \18558 , \18550 , \18557 );
xor \U$18216 ( \18559 , \18547 , \18558 );
not \U$18217 ( \18560 , \3445 );
not \U$18218 ( \18561 , RIbb2e9e0_27);
not \U$18219 ( \18562 , \9010 );
or \U$18220 ( \18563 , \18561 , \18562 );
not \U$18221 ( \18564 , \5954 );
not \U$18222 ( \18565 , \18564 );
nand \U$18223 ( \18566 , \18565 , \4598 );
nand \U$18224 ( \18567 , \18563 , \18566 );
not \U$18225 ( \18568 , \18567 );
or \U$18226 ( \18569 , \18560 , \18568 );
nand \U$18227 ( \18570 , \17345 , \3465 );
nand \U$18228 ( \18571 , \18569 , \18570 );
and \U$18229 ( \18572 , \18559 , \18571 );
and \U$18230 ( \18573 , \18547 , \18558 );
or \U$18231 ( \18574 , \18572 , \18573 );
not \U$18232 ( \18575 , \18574 );
not \U$18233 ( \18576 , \2077 );
not \U$18234 ( \18577 , RIbb2ecb0_21);
not \U$18235 ( \18578 , \9277 );
not \U$18236 ( \18579 , \18578 );
or \U$18237 ( \18580 , \18577 , \18579 );
not \U$18238 ( \18581 , RIbb2ecb0_21);
nand \U$18239 ( \18582 , \18581 , \9278 );
nand \U$18240 ( \18583 , \18580 , \18582 );
not \U$18241 ( \18584 , \18583 );
or \U$18242 ( \18585 , \18576 , \18584 );
nand \U$18243 ( \18586 , \17830 , \2078 );
nand \U$18244 ( \18587 , \18585 , \18586 );
not \U$18245 ( \18588 , \3383 );
not \U$18246 ( \18589 , \17814 );
or \U$18247 ( \18590 , \18588 , \18589 );
not \U$18248 ( \18591 , RIbb2ebc0_23);
not \U$18249 ( \18592 , \14025 );
or \U$18250 ( \18593 , \18591 , \18592 );
nand \U$18251 ( \18594 , \9818 , \2073 );
nand \U$18252 ( \18595 , \18593 , \18594 );
nand \U$18253 ( \18596 , \18595 , \3406 );
nand \U$18254 ( \18597 , \18590 , \18596 );
or \U$18255 ( \18598 , \18587 , \18597 );
not \U$18256 ( \18599 , \854 );
not \U$18257 ( \18600 , \17877 );
or \U$18258 ( \18601 , \18599 , \18600 );
not \U$18259 ( \18602 , RIbb2eda0_19);
not \U$18260 ( \18603 , \13929 );
or \U$18261 ( \18604 , \18602 , \18603 );
nand \U$18262 ( \18605 , \10301 , \843 );
nand \U$18263 ( \18606 , \18604 , \18605 );
nand \U$18264 ( \18607 , \18606 , \853 );
nand \U$18265 ( \18608 , \18601 , \18607 );
nand \U$18266 ( \18609 , \18598 , \18608 );
nand \U$18267 ( \18610 , \18597 , \18587 );
nand \U$18268 ( \18611 , \18609 , \18610 );
not \U$18269 ( \18612 , \18611 );
or \U$18270 ( \18613 , \18575 , \18612 );
or \U$18271 ( \18614 , \18611 , \18574 );
xor \U$18272 ( \18615 , \17507 , \17536 );
and \U$18273 ( \18616 , \18615 , \17547 );
and \U$18274 ( \18617 , \17507 , \17536 );
or \U$18275 ( \18618 , \18616 , \18617 );
not \U$18276 ( \18619 , \2925 );
not \U$18277 ( \18620 , \17793 );
or \U$18278 ( \18621 , \18619 , \18620 );
not \U$18279 ( \18622 , RIbb2e8f0_29);
not \U$18280 ( \18623 , \4696 );
not \U$18281 ( \18624 , \18623 );
not \U$18282 ( \18625 , \18624 );
or \U$18283 ( \18626 , \18622 , \18625 );
nand \U$18284 ( \18627 , \9022 , \2949 );
nand \U$18285 ( \18628 , \18626 , \18627 );
nand \U$18286 ( \18629 , \18628 , \2922 );
nand \U$18287 ( \18630 , \18621 , \18629 );
xor \U$18288 ( \18631 , \18618 , \18630 );
not \U$18289 ( \18632 , \2980 );
not \U$18290 ( \18633 , RIbb2ead0_25);
not \U$18291 ( \18634 , \8639 );
or \U$18292 ( \18635 , \18633 , \18634 );
not \U$18293 ( \18636 , RIbb2ead0_25);
nand \U$18294 ( \18637 , \8638 , \18636 );
nand \U$18295 ( \18638 , \18635 , \18637 );
not \U$18296 ( \18639 , \18638 );
or \U$18297 ( \18640 , \18632 , \18639 );
nand \U$18298 ( \18641 , \17846 , \2963 );
nand \U$18299 ( \18642 , \18640 , \18641 );
and \U$18300 ( \18643 , \18631 , \18642 );
and \U$18301 ( \18644 , \18618 , \18630 );
or \U$18302 ( \18645 , \18643 , \18644 );
nand \U$18303 ( \18646 , \18614 , \18645 );
nand \U$18304 ( \18647 , \18613 , \18646 );
nand \U$18305 ( \18648 , \18537 , \18647 );
nand \U$18306 ( \18649 , \18536 , \18648 );
xor \U$18307 ( \18650 , \18348 , \18377 );
xor \U$18308 ( \18651 , \18650 , \18403 );
xor \U$18309 ( \18652 , \17781 , \18453 );
xnor \U$18310 ( \18653 , \18652 , \18446 );
xor \U$18311 ( \18654 , \18383 , \18394 );
xor \U$18312 ( \18655 , \18654 , \18400 );
xor \U$18313 ( \18656 , \18653 , \18655 );
xor \U$18314 ( \18657 , \18416 , \18427 );
xnor \U$18315 ( \18658 , \18657 , \18434 );
and \U$18316 ( \18659 , \18656 , \18658 );
and \U$18317 ( \18660 , \18653 , \18655 );
or \U$18318 ( \18661 , \18659 , \18660 );
xor \U$18319 ( \18662 , \18651 , \18661 );
xor \U$18320 ( \18663 , \18455 , \18436 );
xor \U$18321 ( \18664 , \18663 , \18410 );
xor \U$18322 ( \18665 , \18662 , \18664 );
xor \U$18323 ( \18666 , \18649 , \18665 );
xor \U$18324 ( \18667 , \17742 , \17798 );
and \U$18325 ( \18668 , \18667 , \17850 );
and \U$18326 ( \18669 , \17742 , \17798 );
or \U$18327 ( \18670 , \18668 , \18669 );
xor \U$18328 ( \18671 , \17857 , \17904 );
and \U$18329 ( \18672 , \18671 , \17950 );
and \U$18330 ( \18673 , \17857 , \17904 );
or \U$18331 ( \18674 , \18672 , \18673 );
xor \U$18332 ( \18675 , \18670 , \18674 );
not \U$18333 ( \18676 , \14067 );
not \U$18334 ( \18677 , \18515 );
or \U$18335 ( \18678 , \18676 , \18677 );
nand \U$18336 ( \18679 , \16637 , \12692 );
nand \U$18337 ( \18680 , \18678 , \18679 );
not \U$18338 ( \18681 , \8450 );
not \U$18339 ( \18682 , \16651 );
or \U$18340 ( \18683 , \18681 , \18682 );
nand \U$18341 ( \18684 , \18506 , \8445 );
nand \U$18342 ( \18685 , \18683 , \18684 );
xor \U$18343 ( \18686 , \18680 , \18685 );
not \U$18344 ( \18687 , \6251 );
not \U$18345 ( \18688 , \18523 );
or \U$18346 ( \18689 , \18687 , \18688 );
nand \U$18347 ( \18690 , \16443 , \6242 );
nand \U$18348 ( \18691 , \18689 , \18690 );
and \U$18349 ( \18692 , \18686 , \18691 );
and \U$18350 ( \18693 , \18680 , \18685 );
or \U$18351 ( \18694 , \18692 , \18693 );
not \U$18352 ( \18695 , \8361 );
not \U$18353 ( \18696 , \18014 );
or \U$18354 ( \18697 , \18695 , \18696 );
nand \U$18355 ( \18698 , \16237 , \8995 );
nand \U$18356 ( \18699 , \18697 , \18698 );
not \U$18357 ( \18700 , \18699 );
not \U$18358 ( \18701 , \16271 );
not \U$18359 ( \18702 , \18025 );
or \U$18360 ( \18703 , \18701 , \18702 );
nand \U$18361 ( \18704 , \16268 , \17470 );
nand \U$18362 ( \18705 , \18703 , \18704 );
not \U$18363 ( \18706 , \18705 );
or \U$18364 ( \18707 , \18700 , \18706 );
or \U$18365 ( \18708 , \18699 , \18705 );
not \U$18366 ( \18709 , \13467 );
not \U$18367 ( \18710 , \18036 );
or \U$18368 ( \18711 , \18709 , \18710 );
nand \U$18369 ( \18712 , \16203 , \14930 );
nand \U$18370 ( \18713 , \18711 , \18712 );
nand \U$18371 ( \18714 , \18708 , \18713 );
nand \U$18372 ( \18715 , \18707 , \18714 );
xor \U$18373 ( \18716 , \18694 , \18715 );
buf \U$18374 ( \18717 , \16541 );
not \U$18375 ( \18718 , \18717 );
not \U$18376 ( \18719 , RIbb2d9f0_61);
not \U$18377 ( \18720 , \1579 );
or \U$18378 ( \18721 , \18719 , \18720 );
not \U$18379 ( \18722 , \1579 );
nand \U$18380 ( \18723 , \18722 , \16254 );
nand \U$18381 ( \18724 , \18721 , \18723 );
not \U$18382 ( \18725 , \18724 );
or \U$18383 ( \18726 , \18718 , \18725 );
nand \U$18384 ( \18727 , \18390 , \16533 );
nand \U$18385 ( \18728 , \18726 , \18727 );
not \U$18386 ( \18729 , \11177 );
not \U$18387 ( \18730 , \16165 );
or \U$18388 ( \18731 , \18729 , \18730 );
not \U$18389 ( \18732 , RIbb2e080_47);
not \U$18390 ( \18733 , \3990 );
or \U$18391 ( \18734 , \18732 , \18733 );
nand \U$18392 ( \18735 , \3109 , \10113 );
nand \U$18393 ( \18736 , \18734 , \18735 );
nand \U$18394 ( \18737 , \18736 , \11176 );
nand \U$18395 ( \18738 , \18731 , \18737 );
xor \U$18396 ( \18739 , \18728 , \18738 );
not \U$18397 ( \18740 , \16675 );
not \U$18398 ( \18741 , RIbb2dbd0_57);
not \U$18399 ( \18742 , \10421 );
or \U$18400 ( \18743 , \18741 , \18742 );
nand \U$18401 ( \18744 , \956 , \14602 );
nand \U$18402 ( \18745 , \18743 , \18744 );
not \U$18403 ( \18746 , \18745 );
or \U$18404 ( \18747 , \18740 , \18746 );
nand \U$18405 ( \18748 , \16673 , \17100 );
nand \U$18406 ( \18749 , \18747 , \18748 );
and \U$18407 ( \18750 , \18739 , \18749 );
and \U$18408 ( \18751 , \18728 , \18738 );
or \U$18409 ( \18752 , \18750 , \18751 );
and \U$18410 ( \18753 , \18716 , \18752 );
and \U$18411 ( \18754 , \18694 , \18715 );
or \U$18412 ( \18755 , \18753 , \18754 );
xor \U$18413 ( \18756 , \18675 , \18755 );
xor \U$18414 ( \18757 , \18666 , \18756 );
not \U$18415 ( \18758 , \18757 );
not \U$18416 ( \18759 , \18758 );
not \U$18417 ( \18760 , \18759 );
xor \U$18418 ( \18761 , \18647 , \18485 );
xnor \U$18419 ( \18762 , \18761 , \18534 );
not \U$18420 ( \18763 , \18762 );
not \U$18421 ( \18764 , \18763 );
xor \U$18422 ( \18765 , \16862 , \16878 );
xor \U$18423 ( \18766 , \18765 , \16889 );
xor \U$18424 ( \18767 , \18547 , \18558 );
xor \U$18425 ( \18768 , \18767 , \18571 );
xor \U$18426 ( \18769 , \18766 , \18768 );
not \U$18427 ( \18770 , \2077 );
not \U$18428 ( \18771 , RIbb2ecb0_21);
not \U$18429 ( \18772 , \14550 );
or \U$18430 ( \18773 , \18771 , \18772 );
nand \U$18431 ( \18774 , \9841 , \2067 );
nand \U$18432 ( \18775 , \18773 , \18774 );
not \U$18433 ( \18776 , \18775 );
or \U$18434 ( \18777 , \18770 , \18776 );
nand \U$18435 ( \18778 , \2078 , \18583 );
nand \U$18436 ( \18779 , \18777 , \18778 );
not \U$18437 ( \18780 , \18779 );
not \U$18438 ( \18781 , \3613 );
not \U$18439 ( \18782 , \17991 );
or \U$18440 ( \18783 , \18781 , \18782 );
not \U$18441 ( \18784 , RIbb2e800_31);
not \U$18442 ( \18785 , \4392 );
or \U$18443 ( \18786 , \18784 , \18785 );
nand \U$18444 ( \18787 , \8375 , \2917 );
nand \U$18445 ( \18788 , \18786 , \18787 );
nand \U$18446 ( \18789 , \18788 , \2940 );
nand \U$18447 ( \18790 , \18783 , \18789 );
not \U$18448 ( \18791 , \18790 );
or \U$18449 ( \18792 , \18780 , \18791 );
not \U$18450 ( \18793 , \18790 );
not \U$18451 ( \18794 , \18793 );
not \U$18452 ( \18795 , \18779 );
not \U$18453 ( \18796 , \18795 );
or \U$18454 ( \18797 , \18794 , \18796 );
not \U$18455 ( \18798 , \854 );
not \U$18456 ( \18799 , \18606 );
or \U$18457 ( \18800 , \18798 , \18799 );
not \U$18458 ( \18801 , RIbb2eda0_19);
not \U$18459 ( \18802 , \13525 );
not \U$18460 ( \18803 , \18802 );
or \U$18461 ( \18804 , \18801 , \18803 );
nand \U$18462 ( \18805 , \10764 , \1776 );
nand \U$18463 ( \18806 , \18804 , \18805 );
nand \U$18464 ( \18807 , \18806 , \853 );
nand \U$18465 ( \18808 , \18800 , \18807 );
nand \U$18466 ( \18809 , \18797 , \18808 );
nand \U$18467 ( \18810 , \18792 , \18809 );
and \U$18468 ( \18811 , \18769 , \18810 );
and \U$18469 ( \18812 , \18766 , \18768 );
or \U$18470 ( \18813 , \18811 , \18812 );
not \U$18471 ( \18814 , \1570 );
not \U$18472 ( \18815 , \18545 );
or \U$18473 ( \18816 , \18814 , \18815 );
not \U$18474 ( \18817 , RIbb2f250_9);
not \U$18475 ( \18818 , \15031 );
or \U$18476 ( \18819 , \18817 , \18818 );
nand \U$18477 ( \18820 , \15030 , \1554 );
nand \U$18478 ( \18821 , \18819 , \18820 );
nand \U$18479 ( \18822 , \18821 , \1533 );
nand \U$18480 ( \18823 , \18816 , \18822 );
not \U$18481 ( \18824 , \18823 );
not \U$18482 ( \18825 , \1077 );
not \U$18483 ( \18826 , \18556 );
or \U$18484 ( \18827 , \18825 , \18826 );
not \U$18485 ( \18828 , RIbb2f160_11);
not \U$18486 ( \18829 , \13977 );
not \U$18487 ( \18830 , \18829 );
or \U$18488 ( \18831 , \18828 , \18830 );
nand \U$18489 ( \18832 , \13977 , \1048 );
nand \U$18490 ( \18833 , \18831 , \18832 );
nand \U$18491 ( \18834 , \18833 , \1011 );
nand \U$18492 ( \18835 , \18827 , \18834 );
not \U$18493 ( \18836 , \18835 );
nand \U$18494 ( \18837 , \18824 , \18836 );
not \U$18495 ( \18838 , \18837 );
not \U$18496 ( \18839 , \1517 );
not \U$18497 ( \18840 , \17288 );
or \U$18498 ( \18841 , \18839 , \18840 );
not \U$18499 ( \18842 , \12932 );
and \U$18500 ( \18843 , RIbb2ef80_15, \18842 );
not \U$18501 ( \18844 , RIbb2ef80_15);
and \U$18502 ( \18845 , \18844 , \14635 );
or \U$18503 ( \18846 , \18843 , \18845 );
nand \U$18504 ( \18847 , \18846 , \1445 );
nand \U$18505 ( \18848 , \18841 , \18847 );
not \U$18506 ( \18849 , \18848 );
or \U$18507 ( \18850 , \18838 , \18849 );
nand \U$18508 ( \18851 , \18835 , \18823 );
nand \U$18509 ( \18852 , \18850 , \18851 );
not \U$18510 ( \18853 , \998 );
not \U$18511 ( \18854 , \16876 );
or \U$18512 ( \18855 , \18853 , \18854 );
not \U$18513 ( \18856 , RIbb2f070_13);
not \U$18514 ( \18857 , \13210 );
not \U$18515 ( \18858 , \18857 );
or \U$18516 ( \18859 , \18856 , \18858 );
nand \U$18517 ( \18860 , \13210 , \906 );
nand \U$18518 ( \18861 , \18859 , \18860 );
nand \U$18519 ( \18862 , \18861 , \916 );
nand \U$18520 ( \18863 , \18855 , \18862 );
not \U$18521 ( \18864 , \2925 );
not \U$18522 ( \18865 , \18628 );
or \U$18523 ( \18866 , \18864 , \18865 );
and \U$18524 ( \18867 , \9108 , RIbb2e8f0_29);
not \U$18525 ( \18868 , \9108 );
and \U$18526 ( \18869 , \18868 , \2949 );
or \U$18527 ( \18870 , \18867 , \18869 );
nand \U$18528 ( \18871 , \18870 , \2922 );
nand \U$18529 ( \18872 , \18866 , \18871 );
xor \U$18530 ( \18873 , \18863 , \18872 );
not \U$18531 ( \18874 , \3445 );
not \U$18532 ( \18875 , RIbb2e9e0_27);
not \U$18533 ( \18876 , \6943 );
or \U$18534 ( \18877 , \18875 , \18876 );
nand \U$18535 ( \18878 , \16943 , \3454 );
nand \U$18536 ( \18879 , \18877 , \18878 );
not \U$18537 ( \18880 , \18879 );
or \U$18538 ( \18881 , \18874 , \18880 );
nand \U$18539 ( \18882 , \18567 , \3465 );
nand \U$18540 ( \18883 , \18881 , \18882 );
and \U$18541 ( \18884 , \18873 , \18883 );
and \U$18542 ( \18885 , \18863 , \18872 );
or \U$18543 ( \18886 , \18884 , \18885 );
xor \U$18544 ( \18887 , \18852 , \18886 );
not \U$18545 ( \18888 , \2963 );
not \U$18546 ( \18889 , \18638 );
or \U$18547 ( \18890 , \18888 , \18889 );
and \U$18548 ( \18891 , RIbb2ead0_25, \13850 );
not \U$18549 ( \18892 , RIbb2ead0_25);
and \U$18550 ( \18893 , \18892 , \7296 );
or \U$18551 ( \18894 , \18891 , \18893 );
nand \U$18552 ( \18895 , \18894 , \2980 );
nand \U$18553 ( \18896 , \18890 , \18895 );
not \U$18554 ( \18897 , \3383 );
not \U$18555 ( \18898 , \18595 );
or \U$18556 ( \18899 , \18897 , \18898 );
not \U$18557 ( \18900 , RIbb2ebc0_23);
not \U$18558 ( \18901 , \13863 );
or \U$18559 ( \18902 , \18900 , \18901 );
nand \U$18560 ( \18903 , \8630 , \3401 );
nand \U$18561 ( \18904 , \18902 , \18903 );
nand \U$18562 ( \18905 , \18904 , \3406 );
nand \U$18563 ( \18906 , \18899 , \18905 );
nor \U$18564 ( \18907 , \18896 , \18906 );
not \U$18565 ( \18908 , \16817 );
not \U$18566 ( \18909 , \18908 );
not \U$18567 ( \18910 , \18909 );
not \U$18568 ( \18911 , \1243 );
or \U$18569 ( \18912 , \18910 , \18911 );
not \U$18570 ( \18913 , \1243 );
nand \U$18571 ( \18914 , \18913 , \16820 );
nand \U$18572 ( \18915 , \18912 , \18914 );
not \U$18573 ( \18916 , \18915 );
not \U$18574 ( \18917 , \1264 );
or \U$18575 ( \18918 , \18916 , \18917 );
not \U$18576 ( \18919 , \1243 );
not \U$18577 ( \18920 , \17750 );
not \U$18578 ( \18921 , \18920 );
or \U$18579 ( \18922 , \18919 , \18921 );
buf \U$18580 ( \18923 , \16703 );
not \U$18581 ( \18924 , \18923 );
nand \U$18582 ( \18925 , \18913 , \18924 );
nand \U$18583 ( \18926 , \18922 , \18925 );
nand \U$18584 ( \18927 , \18926 , \1261 );
nand \U$18585 ( \18928 , \18918 , \18927 );
not \U$18586 ( \18929 , \17506 );
and \U$18587 ( \18930 , \18929 , \1392 );
not \U$18588 ( \18931 , \18929 );
and \U$18589 ( \18932 , \18931 , \17523 );
nor \U$18590 ( \18933 , \18930 , \18932 );
not \U$18591 ( \18934 , \18933 );
not \U$18592 ( \18935 , \1428 );
or \U$18593 ( \18936 , \18934 , \18935 );
nand \U$18594 ( \18937 , \1375 , \17525 );
nand \U$18595 ( \18938 , \18936 , \18937 );
xor \U$18596 ( \18939 , \18928 , \18938 );
not \U$18597 ( \18940 , \1147 );
not \U$18598 ( \18941 , RIbb2f430_5);
not \U$18599 ( \18942 , \16728 );
or \U$18600 ( \18943 , \18941 , \18942 );
nand \U$18601 ( \18944 , \16829 , \1980 );
nand \U$18602 ( \18945 , \18943 , \18944 );
not \U$18603 ( \18946 , \18945 );
or \U$18604 ( \18947 , \18940 , \18946 );
not \U$18605 ( \18948 , RIbb2f430_5);
not \U$18606 ( \18949 , \16710 );
or \U$18607 ( \18950 , \18948 , \18949 );
nand \U$18608 ( \18951 , \16706 , \1980 );
nand \U$18609 ( \18952 , \18950 , \18951 );
nand \U$18610 ( \18953 , \18952 , \1089 );
nand \U$18611 ( \18954 , \18947 , \18953 );
and \U$18612 ( \18955 , \18939 , \18954 );
and \U$18613 ( \18956 , \18928 , \18938 );
or \U$18614 ( \18957 , \18955 , \18956 );
not \U$18615 ( \18958 , \18957 );
or \U$18616 ( \18959 , \18907 , \18958 );
nand \U$18617 ( \18960 , \18896 , \18906 );
nand \U$18618 ( \18961 , \18959 , \18960 );
and \U$18619 ( \18962 , \18887 , \18961 );
and \U$18620 ( \18963 , \18852 , \18886 );
or \U$18621 ( \18964 , \18962 , \18963 );
xor \U$18622 ( \18965 , \18813 , \18964 );
xor \U$18623 ( \18966 , \18587 , \18597 );
xnor \U$18624 ( \18967 , \18966 , \18608 );
not \U$18625 ( \18968 , \18967 );
not \U$18626 ( \18969 , \10119 );
not \U$18627 ( \18970 , \17972 );
or \U$18628 ( \18971 , \18969 , \18970 );
not \U$18629 ( \18972 , RIbb2e170_45);
not \U$18630 ( \18973 , \1853 );
or \U$18631 ( \18974 , \18972 , \18973 );
nand \U$18632 ( \18975 , \4610 , \12003 );
nand \U$18633 ( \18976 , \18974 , \18975 );
nand \U$18634 ( \18977 , \18976 , \10599 );
nand \U$18635 ( \18978 , \18971 , \18977 );
not \U$18636 ( \18979 , \16541 );
not \U$18637 ( \18980 , RIbb2d9f0_61);
not \U$18638 ( \18981 , \14734 );
or \U$18639 ( \18982 , \18980 , \18981 );
nand \U$18640 ( \18983 , \3450 , \16537 );
nand \U$18641 ( \18984 , \18982 , \18983 );
not \U$18642 ( \18985 , \18984 );
or \U$18643 ( \18986 , \18979 , \18985 );
not \U$18644 ( \18987 , RIbb2d9f0_61);
not \U$18645 ( \18988 , \1509 );
or \U$18646 ( \18989 , \18987 , \18988 );
nand \U$18647 ( \18990 , \13308 , \16254 );
nand \U$18648 ( \18991 , \18989 , \18990 );
nand \U$18649 ( \18992 , \18991 , \16533 );
nand \U$18650 ( \18993 , \18986 , \18992 );
xor \U$18651 ( \18994 , \18978 , \18993 );
not \U$18652 ( \18995 , \14613 );
xnor \U$18653 ( \18996 , RIbb2dcc0_55, \3479 );
not \U$18654 ( \18997 , \18996 );
or \U$18655 ( \18998 , \18995 , \18997 );
nand \U$18656 ( \18999 , \17961 , \15181 );
nand \U$18657 ( \19000 , \18998 , \18999 );
and \U$18658 ( \19001 , \18994 , \19000 );
and \U$18659 ( \19002 , \18978 , \18993 );
or \U$18660 ( \19003 , \19001 , \19002 );
or \U$18661 ( \19004 , \18968 , \19003 );
xor \U$18662 ( \19005 , \18618 , \18630 );
xor \U$18663 ( \19006 , \19005 , \18642 );
nand \U$18664 ( \19007 , \19004 , \19006 );
nand \U$18665 ( \19008 , \18968 , \19003 );
nand \U$18666 ( \19009 , \19007 , \19008 );
and \U$18667 ( \19010 , \18965 , \19009 );
and \U$18668 ( \19011 , \18813 , \18964 );
or \U$18669 ( \19012 , \19010 , \19011 );
not \U$18670 ( \19013 , \19012 );
or \U$18671 ( \19014 , \18764 , \19013 );
not \U$18672 ( \19015 , \18762 );
not \U$18673 ( \19016 , \19012 );
not \U$18674 ( \19017 , \19016 );
or \U$18675 ( \19018 , \19015 , \19017 );
xor \U$18676 ( \19019 , \18611 , \18645 );
xor \U$18677 ( \19020 , \19019 , \18574 );
not \U$18678 ( \19021 , \18494 );
not \U$18679 ( \19022 , \18497 );
not \U$18680 ( \19023 , \19022 );
or \U$18681 ( \19024 , \19021 , \19023 );
nand \U$18682 ( \19025 , \18532 , \18497 );
nand \U$18683 ( \19026 , \19024 , \19025 );
and \U$18684 ( \19027 , \19026 , \18529 );
not \U$18685 ( \19028 , \19026 );
not \U$18686 ( \19029 , \18529 );
and \U$18687 ( \19030 , \19028 , \19029 );
nor \U$18688 ( \19031 , \19027 , \19030 );
xor \U$18689 ( \19032 , \19020 , \19031 );
xor \U$18690 ( \19033 , \18041 , \17983 );
xnor \U$18691 ( \19034 , \19033 , \18007 );
and \U$18692 ( \19035 , \19032 , \19034 );
and \U$18693 ( \19036 , \19020 , \19031 );
or \U$18694 ( \19037 , \19035 , \19036 );
nand \U$18695 ( \19038 , \19018 , \19037 );
nand \U$18696 ( \19039 , \19014 , \19038 );
not \U$18697 ( \19040 , \19039 );
or \U$18698 ( \19041 , \18760 , \19040 );
not \U$18699 ( \19042 , \18758 );
not \U$18700 ( \19043 , \19039 );
not \U$18701 ( \19044 , \19043 );
or \U$18702 ( \19045 , \19042 , \19044 );
xor \U$18703 ( \19046 , \18653 , \18655 );
xor \U$18704 ( \19047 , \19046 , \18658 );
xor \U$18705 ( \19048 , \17775 , \17784 );
xor \U$18706 ( \19049 , \19048 , \17795 );
not \U$18707 ( \19050 , \1089 );
not \U$18708 ( \19051 , \18945 );
or \U$18709 ( \19052 , \19050 , \19051 );
nand \U$18710 ( \19053 , \16858 , \1147 );
nand \U$18711 ( \19054 , \19052 , \19053 );
not \U$18712 ( \19055 , \18926 );
not \U$18713 ( \19056 , \1264 );
or \U$18714 ( \19057 , \19055 , \19056 );
nand \U$18715 ( \19058 , \17770 , \1261 );
nand \U$18716 ( \19059 , \19057 , \19058 );
xor \U$18717 ( \19060 , \19054 , \19059 );
not \U$18718 ( \19061 , \1369 );
nand \U$18719 ( \19062 , \19061 , \1244 );
not \U$18720 ( \19063 , \17505 );
not \U$18721 ( \19064 , \19063 );
and \U$18722 ( \19065 , \19062 , \19064 );
not \U$18723 ( \19066 , \1369 );
not \U$18724 ( \19067 , \18913 );
or \U$18725 ( \19068 , \19066 , \19067 );
nand \U$18726 ( \19069 , \19068 , \1312 );
nor \U$18727 ( \19070 , \19065 , \19069 );
not \U$18728 ( \19071 , \1737 );
not \U$18729 ( \19072 , \17545 );
or \U$18730 ( \19073 , \19071 , \19072 );
not \U$18731 ( \19074 , RIbb2f340_7);
not \U$18732 ( \19075 , \16747 );
or \U$18733 ( \19076 , \19074 , \19075 );
not \U$18734 ( \19077 , \16747 );
nand \U$18735 ( \19078 , \19077 , \2700 );
nand \U$18736 ( \19079 , \19076 , \19078 );
nand \U$18737 ( \19080 , \19079 , \1701 );
nand \U$18738 ( \19081 , \19073 , \19080 );
and \U$18739 ( \19082 , \19070 , \19081 );
and \U$18740 ( \19083 , \19060 , \19082 );
and \U$18741 ( \19084 , \19054 , \19059 );
or \U$18742 ( \19085 , \19083 , \19084 );
xor \U$18743 ( \19086 , \17746 , \17760 );
xor \U$18744 ( \19087 , \19086 , \17772 );
xor \U$18745 ( \19088 , \19085 , \19087 );
not \U$18746 ( \19089 , \4712 );
not \U$18747 ( \19090 , \17627 );
or \U$18748 ( \19091 , \19089 , \19090 );
nand \U$18749 ( \19092 , \16902 , \5845 );
nand \U$18750 ( \19093 , \19091 , \19092 );
and \U$18751 ( \19094 , \19088 , \19093 );
and \U$18752 ( \19095 , \19085 , \19087 );
or \U$18753 ( \19096 , \19094 , \19095 );
xor \U$18754 ( \19097 , \19049 , \19096 );
not \U$18755 ( \19098 , \15738 );
not \U$18756 ( \19099 , \18745 );
or \U$18757 ( \19100 , \19098 , \19099 );
not \U$18758 ( \19101 , \15747 );
nand \U$18759 ( \19102 , \17403 , \19101 );
nand \U$18760 ( \19103 , \19100 , \19102 );
not \U$18761 ( \19104 , \19103 );
not \U$18762 ( \19105 , \12965 );
not \U$18763 ( \19106 , \18736 );
or \U$18764 ( \19107 , \19105 , \19106 );
nand \U$18765 ( \19108 , \17382 , \11176 );
nand \U$18766 ( \19109 , \19107 , \19108 );
not \U$18767 ( \19110 , \19109 );
or \U$18768 ( \19111 , \19104 , \19110 );
not \U$18769 ( \19112 , \19103 );
not \U$18770 ( \19113 , \19112 );
not \U$18771 ( \19114 , \19109 );
not \U$18772 ( \19115 , \19114 );
or \U$18773 ( \19116 , \19113 , \19115 );
not \U$18774 ( \19117 , \16533 );
not \U$18775 ( \19118 , \18724 );
or \U$18776 ( \19119 , \19117 , \19118 );
nand \U$18777 ( \19120 , \18991 , \18717 );
nand \U$18778 ( \19121 , \19119 , \19120 );
nand \U$18779 ( \19122 , \19116 , \19121 );
nand \U$18780 ( \19123 , \19111 , \19122 );
and \U$18781 ( \19124 , \19097 , \19123 );
and \U$18782 ( \19125 , \19049 , \19096 );
or \U$18783 ( \19126 , \19124 , \19125 );
xor \U$18784 ( \19127 , \19047 , \19126 );
xor \U$18785 ( \19128 , \18694 , \18715 );
xor \U$18786 ( \19129 , \19128 , \18752 );
and \U$18787 ( \19130 , \19127 , \19129 );
and \U$18788 ( \19131 , \19047 , \19126 );
or \U$18789 ( \19132 , \19130 , \19131 );
xor \U$18790 ( \19133 , \16365 , \16378 );
xor \U$18791 ( \19134 , \19133 , \16390 );
not \U$18792 ( \19135 , \19134 );
xor \U$18793 ( \19136 , \18705 , \18713 );
xnor \U$18794 ( \19137 , \19136 , \18699 );
not \U$18795 ( \19138 , \19137 );
or \U$18796 ( \19139 , \19135 , \19138 );
xor \U$18797 ( \19140 , \18680 , \18685 );
xor \U$18798 ( \19141 , \19140 , \18691 );
nand \U$18799 ( \19142 , \19139 , \19141 );
not \U$18800 ( \19143 , \19134 );
not \U$18801 ( \19144 , \19137 );
nand \U$18802 ( \19145 , \19143 , \19144 );
nand \U$18803 ( \19146 , \19142 , \19145 );
xor \U$18804 ( \19147 , \17947 , \17935 );
and \U$18805 ( \19148 , \19147 , \17918 );
not \U$18806 ( \19149 , \19147 );
and \U$18807 ( \19150 , \19149 , \17919 );
or \U$18808 ( \19151 , \19148 , \19150 );
xor \U$18809 ( \19152 , \18728 , \18738 );
xor \U$18810 ( \19153 , \19152 , \18749 );
or \U$18811 ( \19154 , \19151 , \19153 );
xor \U$18812 ( \19155 , \16851 , \16892 );
xor \U$18813 ( \19156 , \19155 , \16904 );
nand \U$18814 ( \19157 , \19154 , \19156 );
nand \U$18815 ( \19158 , \19151 , \19153 );
nand \U$18816 ( \19159 , \19157 , \19158 );
xor \U$18817 ( \19160 , \19146 , \19159 );
xor \U$18818 ( \19161 , \16356 , \16393 );
xor \U$18819 ( \19162 , \19161 , \16451 );
and \U$18820 ( \19163 , \19160 , \19162 );
and \U$18821 ( \19164 , \19146 , \19159 );
or \U$18822 ( \19165 , \19163 , \19164 );
xor \U$18823 ( \19166 , \19132 , \19165 );
xor \U$18824 ( \19167 , \16621 , \16454 );
xnor \U$18825 ( \19168 , \19167 , \16307 );
xor \U$18826 ( \19169 , \19166 , \19168 );
nand \U$18827 ( \19170 , \19045 , \19169 );
nand \U$18828 ( \19171 , \19041 , \19170 );
xor \U$18829 ( \19172 , \18649 , \18665 );
and \U$18830 ( \19173 , \19172 , \18756 );
and \U$18831 ( \19174 , \18649 , \18665 );
or \U$18832 ( \19175 , \19173 , \19174 );
xor \U$18833 ( \19176 , \18651 , \18661 );
and \U$18834 ( \19177 , \19176 , \18664 );
and \U$18835 ( \19178 , \18651 , \18661 );
or \U$18836 ( \19179 , \19177 , \19178 );
not \U$18837 ( \19180 , \1570 );
not \U$18838 ( \19181 , RIbb2f250_9);
not \U$18839 ( \19182 , \12934 );
or \U$18840 ( \19183 , \19181 , \19182 );
nand \U$18841 ( \19184 , \12933 , \1566 );
nand \U$18842 ( \19185 , \19183 , \19184 );
not \U$18843 ( \19186 , \19185 );
or \U$18844 ( \19187 , \19180 , \19186 );
nand \U$18845 ( \19188 , \18104 , \1533 );
nand \U$18846 ( \19189 , \19187 , \19188 );
not \U$18847 ( \19190 , \19189 );
not \U$18848 ( \19191 , \1428 );
not \U$18849 ( \19192 , \18095 );
or \U$18850 ( \19193 , \19191 , \19192 );
not \U$18851 ( \19194 , \1312 );
not \U$18852 ( \19195 , \16576 );
not \U$18853 ( \19196 , \19195 );
or \U$18854 ( \19197 , \19194 , \19196 );
nand \U$18855 ( \19198 , \16576 , \13990 );
nand \U$18856 ( \19199 , \19197 , \19198 );
nand \U$18857 ( \19200 , \19199 , \1375 );
nand \U$18858 ( \19201 , \19193 , \19200 );
not \U$18859 ( \19202 , \19201 );
and \U$18860 ( \19203 , \1312 , \16729 );
not \U$18861 ( \19204 , \19203 );
and \U$18862 ( \19205 , \19202 , \19204 );
and \U$18863 ( \19206 , \19201 , \19203 );
nor \U$18864 ( \19207 , \19205 , \19206 );
not \U$18865 ( \19208 , \19207 );
and \U$18866 ( \19209 , \19190 , \19208 );
and \U$18867 ( \19210 , \19189 , \19207 );
nor \U$18868 ( \19211 , \19209 , \19210 );
not \U$18869 ( \19212 , \1737 );
and \U$18870 ( \19213 , \18857 , RIbb2f340_7);
not \U$18871 ( \19214 , \18857 );
and \U$18872 ( \19215 , \19214 , \1692 );
or \U$18873 ( \19216 , \19213 , \19215 );
not \U$18874 ( \19217 , \19216 );
or \U$18875 ( \19218 , \19212 , \19217 );
nand \U$18876 ( \19219 , \18365 , \1702 );
nand \U$18877 ( \19220 , \19218 , \19219 );
not \U$18878 ( \19221 , \1147 );
not \U$18879 ( \19222 , RIbb2f430_5);
not \U$18880 ( \19223 , \15456 );
or \U$18881 ( \19224 , \19222 , \19223 );
nand \U$18882 ( \19225 , \13979 , \1980 );
nand \U$18883 ( \19226 , \19224 , \19225 );
not \U$18884 ( \19227 , \19226 );
or \U$18885 ( \19228 , \19221 , \19227 );
nand \U$18886 ( \19229 , \18357 , \1089 );
nand \U$18887 ( \19230 , \19228 , \19229 );
xor \U$18888 ( \19231 , \19220 , \19230 );
not \U$18889 ( \19232 , \1294 );
and \U$18890 ( \19233 , \17681 , \1288 );
not \U$18891 ( \19234 , \17681 );
and \U$18892 ( \19235 , \19234 , \1244 );
or \U$18893 ( \19236 , \19233 , \19235 );
not \U$18894 ( \19237 , \19236 );
or \U$18895 ( \19238 , \19232 , \19237 );
nand \U$18896 ( \19239 , \1264 , \16571 );
nand \U$18897 ( \19240 , \19238 , \19239 );
xor \U$18898 ( \19241 , \19231 , \19240 );
xor \U$18899 ( \19242 , \19211 , \19241 );
not \U$18900 ( \19243 , \19242 );
xor \U$18901 ( \19244 , \16584 , \16597 );
and \U$18902 ( \19245 , \19244 , \16615 );
and \U$18903 ( \19246 , \16584 , \16597 );
or \U$18904 ( \19247 , \19245 , \19246 );
not \U$18905 ( \19248 , \19247 );
or \U$18906 ( \19249 , \19243 , \19248 );
or \U$18907 ( \19250 , \19247 , \19242 );
nand \U$18908 ( \19251 , \19249 , \19250 );
xor \U$18909 ( \19252 , \18359 , \18369 );
and \U$18910 ( \19253 , \19252 , \18376 );
and \U$18911 ( \19254 , \18359 , \18369 );
or \U$18912 ( \19255 , \19253 , \19254 );
not \U$18913 ( \19256 , \16956 );
not \U$18914 ( \19257 , \16938 );
or \U$18915 ( \19258 , \19256 , \19257 );
nand \U$18916 ( \19259 , \19258 , \16926 );
not \U$18917 ( \19260 , \16956 );
nand \U$18918 ( \19261 , \19260 , \16937 );
nand \U$18919 ( \19262 , \19259 , \19261 );
xor \U$18920 ( \19263 , \19255 , \19262 );
not \U$18921 ( \19264 , \16470 );
not \U$18922 ( \19265 , \19264 );
not \U$18923 ( \19266 , \16489 );
or \U$18924 ( \19267 , \19265 , \19266 );
nand \U$18925 ( \19268 , \19267 , \16507 );
not \U$18926 ( \19269 , \16489 );
nand \U$18927 ( \19270 , \19269 , \16470 );
nand \U$18928 ( \19271 , \19268 , \19270 );
xor \U$18929 ( \19272 , \19263 , \19271 );
xor \U$18930 ( \19273 , \19251 , \19272 );
not \U$18931 ( \19274 , \16512 );
not \U$18932 ( \19275 , \16523 );
or \U$18933 ( \19276 , \19274 , \19275 );
nand \U$18934 ( \19277 , \19276 , \16616 );
not \U$18935 ( \19278 , \16523 );
nand \U$18936 ( \19279 , \19278 , \16513 );
nand \U$18937 ( \19280 , \19277 , \19279 );
xor \U$18938 ( \19281 , \19273 , \19280 );
xor \U$18939 ( \19282 , \19179 , \19281 );
xor \U$18940 ( \19283 , \18670 , \18674 );
and \U$18941 ( \19284 , \19283 , \18755 );
and \U$18942 ( \19285 , \18670 , \18674 );
or \U$18943 ( \19286 , \19284 , \19285 );
xor \U$18944 ( \19287 , \19282 , \19286 );
xor \U$18945 ( \19288 , \19175 , \19287 );
xor \U$18946 ( \19289 , \19132 , \19165 );
and \U$18947 ( \19290 , \19289 , \19168 );
and \U$18948 ( \19291 , \19132 , \19165 );
or \U$18949 ( \19292 , \19290 , \19291 );
xor \U$18950 ( \19293 , \19288 , \19292 );
xor \U$18951 ( \19294 , \19171 , \19293 );
xor \U$18952 ( \19295 , \17851 , \17951 );
xor \U$18953 ( \19296 , \19295 , \18044 );
not \U$18954 ( \19297 , \19121 );
not \U$18955 ( \19298 , \19112 );
or \U$18956 ( \19299 , \19297 , \19298 );
or \U$18957 ( \19300 , \19112 , \19121 );
nand \U$18958 ( \19301 , \19299 , \19300 );
and \U$18959 ( \19302 , \19301 , \19114 );
not \U$18960 ( \19303 , \19301 );
and \U$18961 ( \19304 , \19303 , \19109 );
nor \U$18962 ( \19305 , \19302 , \19304 );
not \U$18963 ( \19306 , \19305 );
not \U$18964 ( \19307 , \19306 );
xor \U$18965 ( \19308 , \17993 , \17998 );
xor \U$18966 ( \19309 , \19308 , \18004 );
not \U$18967 ( \19310 , \19309 );
or \U$18968 ( \19311 , \19307 , \19310 );
or \U$18969 ( \19312 , \19309 , \19306 );
xor \U$18970 ( \19313 , \19085 , \19087 );
xor \U$18971 ( \19314 , \19313 , \19093 );
nand \U$18972 ( \19315 , \19312 , \19314 );
nand \U$18973 ( \19316 , \19311 , \19315 );
not \U$18974 ( \19317 , \19316 );
xor \U$18975 ( \19318 , \18517 , \18508 );
xor \U$18976 ( \19319 , \19318 , \18526 );
not \U$18977 ( \19320 , \19319 );
not \U$18978 ( \19321 , \19320 );
xor \U$18979 ( \19322 , \18018 , \18038 );
xnor \U$18980 ( \19323 , \19322 , \18027 );
not \U$18981 ( \19324 , \19323 );
not \U$18982 ( \19325 , \19324 );
or \U$18983 ( \19326 , \19321 , \19325 );
not \U$18984 ( \19327 , \19319 );
not \U$18985 ( \19328 , \19323 );
or \U$18986 ( \19329 , \19327 , \19328 );
xor \U$18987 ( \19330 , \17963 , \17974 );
xor \U$18988 ( \19331 , \19330 , \17980 );
nand \U$18989 ( \19332 , \19329 , \19331 );
nand \U$18990 ( \19333 , \19326 , \19332 );
not \U$18991 ( \19334 , \19333 );
or \U$18992 ( \19335 , \19317 , \19334 );
or \U$18993 ( \19336 , \19333 , \19316 );
xor \U$18994 ( \19337 , \19049 , \19096 );
xor \U$18995 ( \19338 , \19337 , \19123 );
nand \U$18996 ( \19339 , \19336 , \19338 );
nand \U$18997 ( \19340 , \19335 , \19339 );
xor \U$18998 ( \19341 , \19296 , \19340 );
xor \U$18999 ( \19342 , \19146 , \19159 );
xor \U$19000 ( \19343 , \19342 , \19162 );
and \U$19001 ( \19344 , \19341 , \19343 );
and \U$19002 ( \19345 , \19296 , \19340 );
or \U$19003 ( \19346 , \19344 , \19345 );
xor \U$19004 ( \19347 , \19047 , \19126 );
xor \U$19005 ( \19348 , \19347 , \19129 );
not \U$19006 ( \19349 , \19141 );
and \U$19007 ( \19350 , \19134 , \19349 );
not \U$19008 ( \19351 , \19134 );
and \U$19009 ( \19352 , \19351 , \19141 );
nor \U$19010 ( \19353 , \19350 , \19352 );
and \U$19011 ( \19354 , \19353 , \19144 );
not \U$19012 ( \19355 , \19353 );
not \U$19013 ( \19356 , \19144 );
and \U$19014 ( \19357 , \19355 , \19356 );
nor \U$19015 ( \19358 , \19354 , \19357 );
xor \U$19016 ( \19359 , \18766 , \18768 );
xor \U$19017 ( \19360 , \19359 , \18810 );
xor \U$19018 ( \19361 , \18808 , \18795 );
xnor \U$19019 ( \19362 , \19361 , \18793 );
not \U$19020 ( \19363 , \19362 );
xor \U$19021 ( \19364 , \18863 , \18872 );
xor \U$19022 ( \19365 , \19364 , \18883 );
not \U$19023 ( \19366 , \19365 );
not \U$19024 ( \19367 , \19366 );
or \U$19025 ( \19368 , \19363 , \19367 );
not \U$19026 ( \19369 , \15181 );
not \U$19027 ( \19370 , \18996 );
or \U$19028 ( \19371 , \19369 , \19370 );
and \U$19029 ( \19372 , RIbb2dcc0_55, \1685 );
not \U$19030 ( \19373 , RIbb2dcc0_55);
and \U$19031 ( \19374 , \19373 , \1686 );
nor \U$19032 ( \19375 , \19372 , \19374 );
nand \U$19033 ( \19376 , \19375 , \14613 );
nand \U$19034 ( \19377 , \19371 , \19376 );
not \U$19035 ( \19378 , \9098 );
not \U$19036 ( \19379 , RIbb2e260_43);
not \U$19037 ( \19380 , \3516 );
or \U$19038 ( \19381 , \19379 , \19380 );
not \U$19039 ( \19382 , RIbb2e260_43);
nand \U$19040 ( \19383 , \19382 , \3341 );
nand \U$19041 ( \19384 , \19381 , \19383 );
not \U$19042 ( \19385 , \19384 );
or \U$19043 ( \19386 , \19378 , \19385 );
nand \U$19044 ( \19387 , \17497 , \9099 );
nand \U$19045 ( \19388 , \19386 , \19387 );
xor \U$19046 ( \19389 , \19377 , \19388 );
not \U$19047 ( \19390 , \10119 );
not \U$19048 ( \19391 , \18976 );
or \U$19049 ( \19392 , \19390 , \19391 );
and \U$19050 ( \19393 , \2114 , \9094 );
not \U$19051 ( \19394 , \2114 );
and \U$19052 ( \19395 , \19394 , RIbb2e170_45);
or \U$19053 ( \19396 , \19393 , \19395 );
nand \U$19054 ( \19397 , \19396 , \10117 );
nand \U$19055 ( \19398 , \19392 , \19397 );
and \U$19056 ( \19399 , \19389 , \19398 );
and \U$19057 ( \19400 , \19377 , \19388 );
or \U$19058 ( \19401 , \19399 , \19400 );
nand \U$19059 ( \19402 , \19368 , \19401 );
not \U$19060 ( \19403 , \19366 );
not \U$19061 ( \19404 , \19362 );
nand \U$19062 ( \19405 , \19403 , \19404 );
nand \U$19063 ( \19406 , \19402 , \19405 );
xor \U$19064 ( \19407 , \19360 , \19406 );
xor \U$19065 ( \19408 , \18957 , \18906 );
not \U$19066 ( \19409 , \18896 );
xnor \U$19067 ( \19410 , \19408 , \19409 );
not \U$19068 ( \19411 , \19410 );
xor \U$19069 ( \19412 , \18836 , \18823 );
xnor \U$19070 ( \19413 , \19412 , \18848 );
not \U$19071 ( \19414 , \19413 );
not \U$19072 ( \19415 , \15746 );
not \U$19073 ( \19416 , RIbb2dbd0_57);
not \U$19074 ( \19417 , \5003 );
or \U$19075 ( \19418 , \19416 , \19417 );
nand \U$19076 ( \19419 , \1548 , \15741 );
nand \U$19077 ( \19420 , \19418 , \19419 );
not \U$19078 ( \19421 , \19420 );
or \U$19079 ( \19422 , \19415 , \19421 );
nand \U$19080 ( \19423 , \17413 , \17100 );
nand \U$19081 ( \19424 , \19422 , \19423 );
not \U$19082 ( \19425 , \4791 );
not \U$19083 ( \19426 , \17423 );
or \U$19084 ( \19427 , \19425 , \19426 );
not \U$19085 ( \19428 , RIbb2e710_33);
not \U$19086 ( \19429 , \4085 );
not \U$19087 ( \19430 , \19429 );
or \U$19088 ( \19431 , \19428 , \19430 );
nand \U$19089 ( \19432 , \13551 , \18295 );
nand \U$19090 ( \19433 , \19431 , \19432 );
nand \U$19091 ( \19434 , \19433 , \3887 );
nand \U$19092 ( \19435 , \19427 , \19434 );
or \U$19093 ( \19436 , \19424 , \19435 );
not \U$19094 ( \19437 , \13295 );
not \U$19095 ( \19438 , RIbb2df90_49);
not \U$19096 ( \19439 , \4339 );
or \U$19097 ( \19440 , \19438 , \19439 );
nand \U$19098 ( \19441 , \17380 , \12278 );
nand \U$19099 ( \19442 , \19440 , \19441 );
not \U$19100 ( \19443 , \19442 );
or \U$19101 ( \19444 , \19437 , \19443 );
nand \U$19102 ( \19445 , \17372 , \16427 );
nand \U$19103 ( \19446 , \19444 , \19445 );
nand \U$19104 ( \19447 , \19436 , \19446 );
nand \U$19105 ( \19448 , \19435 , \19424 );
and \U$19106 ( \19449 , \19447 , \19448 );
nand \U$19107 ( \19450 , \19414 , \19449 );
not \U$19108 ( \19451 , \19450 );
or \U$19109 ( \19452 , \19411 , \19451 );
nand \U$19110 ( \19453 , \19447 , \19448 );
nand \U$19111 ( \19454 , \19453 , \19413 );
nand \U$19112 ( \19455 , \19452 , \19454 );
and \U$19113 ( \19456 , \19407 , \19455 );
and \U$19114 ( \19457 , \19360 , \19406 );
or \U$19115 ( \19458 , \19456 , \19457 );
nor \U$19116 ( \19459 , \19358 , \19458 );
xor \U$19117 ( \19460 , \19156 , \19153 );
xnor \U$19118 ( \19461 , \19460 , \19151 );
buf \U$19119 ( \19462 , \19461 );
or \U$19120 ( \19463 , \19459 , \19462 );
nand \U$19121 ( \19464 , \19458 , \19358 );
nand \U$19122 ( \19465 , \19463 , \19464 );
xor \U$19123 ( \19466 , \19348 , \19465 );
not \U$19124 ( \19467 , \17641 );
not \U$19125 ( \19468 , \19467 );
xnor \U$19126 ( \19469 , \17257 , \17251 );
not \U$19127 ( \19470 , \19469 );
or \U$19128 ( \19471 , \19468 , \19470 );
or \U$19129 ( \19472 , \19467 , \19469 );
nand \U$19130 ( \19473 , \19471 , \19472 );
and \U$19131 ( \19474 , \19466 , \19473 );
and \U$19132 ( \19475 , \19348 , \19465 );
or \U$19133 ( \19476 , \19474 , \19475 );
xor \U$19134 ( \19477 , \19346 , \19476 );
xor \U$19135 ( \19478 , \17249 , \17646 );
xor \U$19136 ( \19479 , \19478 , \18048 );
and \U$19137 ( \19480 , \19477 , \19479 );
and \U$19138 ( \19481 , \19346 , \19476 );
or \U$19139 ( \19482 , \19480 , \19481 );
xor \U$19140 ( \19483 , \19294 , \19482 );
xor \U$19141 ( \19484 , \18481 , \19483 );
xor \U$19142 ( \19485 , \18813 , \18964 );
xor \U$19143 ( \19486 , \19485 , \19009 );
not \U$19144 ( \19487 , \19486 );
not \U$19145 ( \19488 , \19487 );
xor \U$19146 ( \19489 , \17468 , \17499 );
not \U$19147 ( \19490 , \17481 );
and \U$19148 ( \19491 , \19489 , \19490 );
not \U$19149 ( \19492 , \19489 );
and \U$19150 ( \19493 , \19492 , \17481 );
nor \U$19151 ( \19494 , \19491 , \19493 );
not \U$19152 ( \19495 , \19494 );
not \U$19153 ( \19496 , \19495 );
xor \U$19154 ( \19497 , \17446 , \17415 );
xnor \U$19155 ( \19498 , \19497 , \17432 );
not \U$19156 ( \19499 , \19498 );
not \U$19157 ( \19500 , \19499 );
or \U$19158 ( \19501 , \19496 , \19500 );
not \U$19159 ( \19502 , \19498 );
not \U$19160 ( \19503 , \19494 );
or \U$19161 ( \19504 , \19502 , \19503 );
xor \U$19162 ( \19505 , \17357 , \17374 );
xor \U$19163 ( \19506 , \19505 , \17392 );
nand \U$19164 ( \19507 , \19504 , \19506 );
nand \U$19165 ( \19508 , \19501 , \19507 );
not \U$19166 ( \19509 , \19508 );
xor \U$19167 ( \19510 , \19006 , \18967 );
xnor \U$19168 ( \19511 , \19510 , \19003 );
not \U$19169 ( \19512 , \19511 );
or \U$19170 ( \19513 , \19509 , \19512 );
or \U$19171 ( \19514 , \19508 , \19511 );
xor \U$19172 ( \19515 , \17598 , \17613 );
xor \U$19173 ( \19516 , \19515 , \17629 );
not \U$19174 ( \19517 , \19516 );
xor \U$19175 ( \19518 , \18978 , \18993 );
xor \U$19176 ( \19519 , \19518 , \19000 );
not \U$19177 ( \19520 , \19519 );
or \U$19178 ( \19521 , \19517 , \19520 );
or \U$19179 ( \19522 , \19519 , \19516 );
not \U$19180 ( \19523 , \5845 );
not \U$19181 ( \19524 , \17620 );
or \U$19182 ( \19525 , \19523 , \19524 );
not \U$19183 ( \19526 , RIbb2e620_35);
not \U$19184 ( \19527 , \15605 );
or \U$19185 ( \19528 , \19526 , \19527 );
nand \U$19186 ( \19529 , \13732 , \3866 );
nand \U$19187 ( \19530 , \19528 , \19529 );
nand \U$19188 ( \19531 , \19530 , \4712 );
nand \U$19189 ( \19532 , \19525 , \19531 );
not \U$19190 ( \19533 , \915 );
not \U$19191 ( \19534 , RIbb2f070_13);
not \U$19192 ( \19535 , \18829 );
or \U$19193 ( \19536 , \19534 , \19535 );
nand \U$19194 ( \19537 , \13977 , \906 );
nand \U$19195 ( \19538 , \19536 , \19537 );
not \U$19196 ( \19539 , \19538 );
or \U$19197 ( \19540 , \19533 , \19539 );
not \U$19198 ( \19541 , RIbb2f070_13);
not \U$19199 ( \19542 , \18552 );
or \U$19200 ( \19543 , \19541 , \19542 );
nand \U$19201 ( \19544 , \13545 , \1656 );
nand \U$19202 ( \19545 , \19543 , \19544 );
nand \U$19203 ( \19546 , \998 , \19545 );
nand \U$19204 ( \19547 , \19540 , \19546 );
not \U$19205 ( \19548 , \19547 );
not \U$19206 ( \19549 , \1011 );
not \U$19207 ( \19550 , RIbb2f160_11);
not \U$19208 ( \19551 , \15031 );
or \U$19209 ( \19552 , \19550 , \19551 );
nand \U$19210 ( \19553 , \16782 , \1805 );
nand \U$19211 ( \19554 , \19552 , \19553 );
not \U$19212 ( \19555 , \19554 );
or \U$19213 ( \19556 , \19549 , \19555 );
not \U$19214 ( \19557 , RIbb2f160_11);
not \U$19215 ( \19558 , \16309 );
or \U$19216 ( \19559 , \19557 , \19558 );
nand \U$19217 ( \19560 , \14526 , \1048 );
nand \U$19218 ( \19561 , \19559 , \19560 );
nand \U$19219 ( \19562 , \19561 , \1077 );
nand \U$19220 ( \19563 , \19556 , \19562 );
not \U$19221 ( \19564 , \19563 );
or \U$19222 ( \19565 , \19548 , \19564 );
or \U$19223 ( \19566 , \19563 , \19547 );
not \U$19224 ( \19567 , \1445 );
and \U$19225 ( \19568 , RIbb2ef80_15, \18857 );
not \U$19226 ( \19569 , RIbb2ef80_15);
and \U$19227 ( \19570 , \19569 , \13210 );
or \U$19228 ( \19571 , \19568 , \19570 );
not \U$19229 ( \19572 , \19571 );
or \U$19230 ( \19573 , \19567 , \19572 );
and \U$19231 ( \19574 , RIbb2ef80_15, \14838 );
not \U$19232 ( \19575 , RIbb2ef80_15);
and \U$19233 ( \19576 , \19575 , \14843 );
or \U$19234 ( \19577 , \19574 , \19576 );
nand \U$19235 ( \19578 , \19577 , \1517 );
nand \U$19236 ( \19579 , \19573 , \19578 );
nand \U$19237 ( \19580 , \19566 , \19579 );
nand \U$19238 ( \19581 , \19565 , \19580 );
nor \U$19239 ( \19582 , \19532 , \19581 );
xor \U$19240 ( \19583 , \18928 , \18938 );
xor \U$19241 ( \19584 , \19583 , \18954 );
not \U$19242 ( \19585 , \19584 );
or \U$19243 ( \19586 , \19582 , \19585 );
nand \U$19244 ( \19587 , \19532 , \19581 );
nand \U$19245 ( \19588 , \19586 , \19587 );
nand \U$19246 ( \19589 , \19522 , \19588 );
nand \U$19247 ( \19590 , \19521 , \19589 );
nand \U$19248 ( \19591 , \19514 , \19590 );
nand \U$19249 ( \19592 , \19513 , \19591 );
not \U$19250 ( \19593 , \19592 );
not \U$19251 ( \19594 , \19593 );
or \U$19252 ( \19595 , \19488 , \19594 );
xor \U$19253 ( \19596 , \19054 , \19059 );
xor \U$19254 ( \19597 , \19596 , \19082 );
not \U$19255 ( \19598 , \1570 );
not \U$19256 ( \19599 , \18821 );
or \U$19257 ( \19600 , \19598 , \19599 );
not \U$19258 ( \19601 , RIbb2f250_9);
not \U$19259 ( \19602 , \15754 );
or \U$19260 ( \19603 , \19601 , \19602 );
nand \U$19261 ( \19604 , \16562 , \5064 );
nand \U$19262 ( \19605 , \19603 , \19604 );
nand \U$19263 ( \19606 , \19605 , \1533 );
nand \U$19264 ( \19607 , \19600 , \19606 );
not \U$19265 ( \19608 , \19607 );
not \U$19266 ( \19609 , \1077 );
not \U$19267 ( \19610 , \18833 );
or \U$19268 ( \19611 , \19609 , \19610 );
nand \U$19269 ( \19612 , \19561 , \1011 );
nand \U$19270 ( \19613 , \19611 , \19612 );
not \U$19271 ( \19614 , \19613 );
or \U$19272 ( \19615 , \19608 , \19614 );
or \U$19273 ( \19616 , \19613 , \19607 );
xor \U$19274 ( \19617 , \19070 , \19081 );
nand \U$19275 ( \19618 , \19616 , \19617 );
nand \U$19276 ( \19619 , \19615 , \19618 );
xor \U$19277 ( \19620 , \19597 , \19619 );
not \U$19278 ( \19621 , \915 );
not \U$19279 ( \19622 , \19545 );
or \U$19280 ( \19623 , \19621 , \19622 );
nand \U$19281 ( \19624 , \18861 , \998 );
nand \U$19282 ( \19625 , \19623 , \19624 );
not \U$19283 ( \19626 , \1445 );
not \U$19284 ( \19627 , \19577 );
or \U$19285 ( \19628 , \19626 , \19627 );
nand \U$19286 ( \19629 , \18846 , \1517 );
nand \U$19287 ( \19630 , \19628 , \19629 );
xor \U$19288 ( \19631 , \19625 , \19630 );
not \U$19289 ( \19632 , \2921 );
not \U$19290 ( \19633 , RIbb2e8f0_29);
not \U$19291 ( \19634 , \14041 );
or \U$19292 ( \19635 , \19633 , \19634 );
nand \U$19293 ( \19636 , \7308 , \4800 );
nand \U$19294 ( \19637 , \19635 , \19636 );
not \U$19295 ( \19638 , \19637 );
or \U$19296 ( \19639 , \19632 , \19638 );
nand \U$19297 ( \19640 , \18870 , \2925 );
nand \U$19298 ( \19641 , \19639 , \19640 );
and \U$19299 ( \19642 , \19631 , \19641 );
and \U$19300 ( \19643 , \19625 , \19630 );
or \U$19301 ( \19644 , \19642 , \19643 );
and \U$19302 ( \19645 , \19620 , \19644 );
and \U$19303 ( \19646 , \19597 , \19619 );
or \U$19304 ( \19647 , \19645 , \19646 );
not \U$19305 ( \19648 , \14067 );
and \U$19306 ( \19649 , RIbb2dea0_51, \1281 );
not \U$19307 ( \19650 , RIbb2dea0_51);
and \U$19308 ( \19651 , \19650 , \12036 );
or \U$19309 ( \19652 , \19649 , \19651 );
not \U$19310 ( \19653 , \19652 );
or \U$19311 ( \19654 , \19648 , \19653 );
nand \U$19312 ( \19655 , \17611 , \12692 );
nand \U$19313 ( \19656 , \19654 , \19655 );
not \U$19314 ( \19657 , \19656 );
not \U$19315 ( \19658 , \7104 );
not \U$19316 ( \19659 , \17578 );
or \U$19317 ( \19660 , \19658 , \19659 );
and \U$19318 ( \19661 , RIbb2e440_39, \6172 );
not \U$19319 ( \19662 , RIbb2e440_39);
and \U$19320 ( \19663 , \19662 , \13903 );
or \U$19321 ( \19664 , \19661 , \19663 );
nand \U$19322 ( \19665 , \19664 , \7103 );
nand \U$19323 ( \19666 , \19660 , \19665 );
not \U$19324 ( \19667 , \19666 );
or \U$19325 ( \19668 , \19657 , \19667 );
or \U$19326 ( \19669 , \19656 , \19666 );
not \U$19327 ( \19670 , \6242 );
not \U$19328 ( \19671 , \17596 );
or \U$19329 ( \19672 , \19670 , \19671 );
not \U$19330 ( \19673 , RIbb2e530_37);
not \U$19331 ( \19674 , \4021 );
or \U$19332 ( \19675 , \19673 , \19674 );
not \U$19333 ( \19676 , \3021 );
nand \U$19334 ( \19677 , \19676 , \6246 );
nand \U$19335 ( \19678 , \19675 , \19677 );
nand \U$19336 ( \19679 , \19678 , \6251 );
nand \U$19337 ( \19680 , \19672 , \19679 );
nand \U$19338 ( \19681 , \19669 , \19680 );
nand \U$19339 ( \19682 , \19668 , \19681 );
not \U$19340 ( \19683 , \16257 );
not \U$19341 ( \19684 , \17479 );
or \U$19342 ( \19685 , \19683 , \19684 );
and \U$19343 ( \19686 , RIbb2dae0_59, \1068 );
not \U$19344 ( \19687 , RIbb2dae0_59);
and \U$19345 ( \19688 , \19687 , \13610 );
nor \U$19346 ( \19689 , \19686 , \19688 );
nand \U$19347 ( \19690 , \19689 , \16271 );
nand \U$19348 ( \19691 , \19685 , \19690 );
not \U$19349 ( \19692 , \8353 );
not \U$19350 ( \19693 , \17459 );
or \U$19351 ( \19694 , \19692 , \19693 );
and \U$19352 ( \19695 , \7097 , \3139 );
not \U$19353 ( \19696 , \7097 );
and \U$19354 ( \19697 , \19696 , \17568 );
nor \U$19355 ( \19698 , \19695 , \19697 );
not \U$19356 ( \19699 , \19698 );
nand \U$19357 ( \19700 , \19699 , \8362 );
nand \U$19358 ( \19701 , \19694 , \19700 );
xor \U$19359 ( \19702 , \19691 , \19701 );
not \U$19360 ( \19703 , \17562 );
not \U$19361 ( \19704 , RIbb2ddb0_53);
not \U$19362 ( \19705 , \8862 );
or \U$19363 ( \19706 , \19704 , \19705 );
nand \U$19364 ( \19707 , \3053 , \16210 );
nand \U$19365 ( \19708 , \19706 , \19707 );
not \U$19366 ( \19709 , \19708 );
or \U$19367 ( \19710 , \19703 , \19709 );
nand \U$19368 ( \19711 , \17561 , \15688 );
nand \U$19369 ( \19712 , \19710 , \19711 );
and \U$19370 ( \19713 , \19702 , \19712 );
and \U$19371 ( \19714 , \19691 , \19701 );
or \U$19372 ( \19715 , \19713 , \19714 );
or \U$19373 ( \19716 , \19682 , \19715 );
not \U$19374 ( \19717 , \17275 );
not \U$19375 ( \19718 , RIbb2d900_63);
not \U$19376 ( \19719 , \8754 );
or \U$19377 ( \19720 , \19718 , \19719 );
not \U$19378 ( \19721 , RIbb2d900_63);
nand \U$19379 ( \19722 , \1508 , \19721 );
nand \U$19380 ( \19723 , \19720 , \19722 );
not \U$19381 ( \19724 , \19723 );
or \U$19382 ( \19725 , \19717 , \19724 );
nand \U$19383 ( \19726 , \17353 , RIbb2d888_64);
nand \U$19384 ( \19727 , \19725 , \19726 );
not \U$19385 ( \19728 , \19727 );
not \U$19386 ( \19729 , \11177 );
not \U$19387 ( \19730 , \17390 );
or \U$19388 ( \19731 , \19729 , \19730 );
not \U$19389 ( \19732 , RIbb2e080_47);
not \U$19390 ( \19733 , \1337 );
not \U$19391 ( \19734 , \19733 );
or \U$19392 ( \19735 , \19732 , \19734 );
nand \U$19393 ( \19736 , \1337 , \12971 );
nand \U$19394 ( \19737 , \19735 , \19736 );
nand \U$19395 ( \19738 , \19737 , \11176 );
nand \U$19396 ( \19739 , \19731 , \19738 );
not \U$19397 ( \19740 , \19739 );
or \U$19398 ( \19741 , \19728 , \19740 );
or \U$19399 ( \19742 , \19739 , \19727 );
not \U$19400 ( \19743 , \16533 );
not \U$19401 ( \19744 , \18984 );
or \U$19402 ( \19745 , \19743 , \19744 );
not \U$19403 ( \19746 , RIbb2d9f0_61);
not \U$19404 ( \19747 , \19746 );
not \U$19405 ( \19748 , \984 );
or \U$19406 ( \19749 , \19747 , \19748 );
or \U$19407 ( \19750 , \986 , \19746 );
nand \U$19408 ( \19751 , \19749 , \19750 );
nand \U$19409 ( \19752 , \19751 , \16541 );
nand \U$19410 ( \19753 , \19745 , \19752 );
nand \U$19411 ( \19754 , \19742 , \19753 );
nand \U$19412 ( \19755 , \19741 , \19754 );
nand \U$19413 ( \19756 , \19716 , \19755 );
nand \U$19414 ( \19757 , \19682 , \19715 );
nand \U$19415 ( \19758 , \19756 , \19757 );
xor \U$19416 ( \19759 , \19647 , \19758 );
not \U$19417 ( \19760 , \3382 );
not \U$19418 ( \19761 , \18904 );
or \U$19419 ( \19762 , \19760 , \19761 );
not \U$19420 ( \19763 , RIbb2ebc0_23);
not \U$19421 ( \19764 , \12819 );
or \U$19422 ( \19765 , \19763 , \19764 );
nand \U$19423 ( \19766 , \9277 , \3401 );
nand \U$19424 ( \19767 , \19765 , \19766 );
nand \U$19425 ( \19768 , \19767 , \3406 );
nand \U$19426 ( \19769 , \19762 , \19768 );
not \U$19427 ( \19770 , \2980 );
not \U$19428 ( \19771 , RIbb2ead0_25);
not \U$19429 ( \19772 , \12210 );
or \U$19430 ( \19773 , \19771 , \19772 );
nand \U$19431 ( \19774 , \14024 , \18636 );
nand \U$19432 ( \19775 , \19773 , \19774 );
not \U$19433 ( \19776 , \19775 );
or \U$19434 ( \19777 , \19770 , \19776 );
nand \U$19435 ( \19778 , \18894 , \2963 );
nand \U$19436 ( \19779 , \19777 , \19778 );
buf \U$19437 ( \19780 , \19779 );
nor \U$19438 ( \19781 , \19769 , \19780 );
not \U$19439 ( \19782 , \2078 );
not \U$19440 ( \19783 , \18775 );
or \U$19441 ( \19784 , \19782 , \19783 );
not \U$19442 ( \19785 , RIbb2ecb0_21);
not \U$19443 ( \19786 , \12744 );
or \U$19444 ( \19787 , \19785 , \19786 );
nand \U$19445 ( \19788 , \10301 , \5481 );
nand \U$19446 ( \19789 , \19787 , \19788 );
nand \U$19447 ( \19790 , \19789 , \2077 );
nand \U$19448 ( \19791 , \19784 , \19790 );
not \U$19449 ( \19792 , \19791 );
or \U$19450 ( \19793 , \19781 , \19792 );
nand \U$19451 ( \19794 , \19780 , \19769 );
nand \U$19452 ( \19795 , \19793 , \19794 );
not \U$19453 ( \19796 , \1147 );
not \U$19454 ( \19797 , \18952 );
or \U$19455 ( \19798 , \19796 , \19797 );
not \U$19456 ( \19799 , RIbb2f430_5);
not \U$19457 ( \19800 , \17750 );
or \U$19458 ( \19801 , \19799 , \19800 );
nand \U$19459 ( \19802 , \18923 , \1980 );
nand \U$19460 ( \19803 , \19801 , \19802 );
nand \U$19461 ( \19804 , \19803 , \1089 );
nand \U$19462 ( \19805 , \19798 , \19804 );
and \U$19463 ( \19806 , \1375 , \19064 );
xor \U$19464 ( \19807 , \19805 , \19806 );
nand \U$19465 ( \19808 , \1898 , \1256 );
and \U$19466 ( \19809 , \17506 , \19808 );
and \U$19467 ( \19810 , RIbb2f4a8_4, RIbb2f430_5);
nor \U$19468 ( \19811 , \19809 , \19810 );
and \U$19469 ( \19812 , \1253 , \19811 );
not \U$19470 ( \19813 , \1147 );
not \U$19471 ( \19814 , \19803 );
or \U$19472 ( \19815 , \19813 , \19814 );
not \U$19473 ( \19816 , RIbb2f430_5);
not \U$19474 ( \19817 , \18908 );
or \U$19475 ( \19818 , \19816 , \19817 );
nand \U$19476 ( \19819 , \17529 , \1980 );
nand \U$19477 ( \19820 , \19818 , \19819 );
nand \U$19478 ( \19821 , \19820 , \1089 );
nand \U$19479 ( \19822 , \19815 , \19821 );
and \U$19480 ( \19823 , \19812 , \19822 );
and \U$19481 ( \19824 , \19807 , \19823 );
and \U$19482 ( \19825 , \19805 , \19806 );
or \U$19483 ( \19826 , \19824 , \19825 );
not \U$19484 ( \19827 , \1701 );
not \U$19485 ( \19828 , RIbb2f340_7);
not \U$19486 ( \19829 , \16727 );
or \U$19487 ( \19830 , \19828 , \19829 );
buf \U$19488 ( \19831 , \16726 );
nand \U$19489 ( \19832 , \19831 , \2700 );
nand \U$19490 ( \19833 , \19830 , \19832 );
not \U$19491 ( \19834 , \19833 );
or \U$19492 ( \19835 , \19827 , \19834 );
nand \U$19493 ( \19836 , \19079 , \1737 );
nand \U$19494 ( \19837 , \19835 , \19836 );
not \U$19495 ( \19838 , \17745 );
not \U$19496 ( \19839 , \18913 );
or \U$19497 ( \19840 , \19838 , \19839 );
not \U$19498 ( \19841 , \17745 );
nand \U$19499 ( \19842 , \1243 , \19841 );
nand \U$19500 ( \19843 , \19840 , \19842 );
not \U$19501 ( \19844 , \19843 );
not \U$19502 ( \19845 , \1264 );
or \U$19503 ( \19846 , \19844 , \19845 );
nand \U$19504 ( \19847 , \1261 , \18915 );
nand \U$19505 ( \19848 , \19846 , \19847 );
xor \U$19506 ( \19849 , \19837 , \19848 );
not \U$19507 ( \19850 , \1570 );
not \U$19508 ( \19851 , \19605 );
or \U$19509 ( \19852 , \19850 , \19851 );
not \U$19510 ( \19853 , RIbb2f250_9);
not \U$19511 ( \19854 , \16844 );
or \U$19512 ( \19855 , \19853 , \19854 );
nand \U$19513 ( \19856 , \16575 , \1566 );
nand \U$19514 ( \19857 , \19855 , \19856 );
nand \U$19515 ( \19858 , \19857 , \1533 );
nand \U$19516 ( \19859 , \19852 , \19858 );
and \U$19517 ( \19860 , \19849 , \19859 );
and \U$19518 ( \19861 , \19837 , \19848 );
or \U$19519 ( \19862 , \19860 , \19861 );
xor \U$19520 ( \19863 , \19826 , \19862 );
not \U$19521 ( \19864 , \3445 );
not \U$19522 ( \19865 , RIbb2e9e0_27);
not \U$19523 ( \19866 , \8639 );
or \U$19524 ( \19867 , \19865 , \19866 );
not \U$19525 ( \19868 , \6936 );
buf \U$19526 ( \19869 , \19868 );
not \U$19527 ( \19870 , \19869 );
nand \U$19528 ( \19871 , \19870 , \3454 );
nand \U$19529 ( \19872 , \19867 , \19871 );
not \U$19530 ( \19873 , \19872 );
or \U$19531 ( \19874 , \19864 , \19873 );
nand \U$19532 ( \19875 , \18879 , \3465 );
nand \U$19533 ( \19876 , \19874 , \19875 );
and \U$19534 ( \19877 , \19863 , \19876 );
and \U$19535 ( \19878 , \19826 , \19862 );
or \U$19536 ( \19879 , \19877 , \19878 );
xor \U$19537 ( \19880 , \19795 , \19879 );
not \U$19538 ( \19881 , \3613 );
not \U$19539 ( \19882 , \18788 );
or \U$19540 ( \19883 , \19881 , \19882 );
and \U$19541 ( \19884 , RIbb2e800_31, \10555 );
not \U$19542 ( \19885 , RIbb2e800_31);
and \U$19543 ( \19886 , \19885 , \4697 );
or \U$19544 ( \19887 , \19884 , \19886 );
nand \U$19545 ( \19888 , \19887 , \2940 );
nand \U$19546 ( \19889 , \19883 , \19888 );
not \U$19547 ( \19890 , \836 );
not \U$19548 ( \19891 , \17444 );
or \U$19549 ( \19892 , \19890 , \19891 );
not \U$19550 ( \19893 , RIbb2ee90_17);
not \U$19551 ( \19894 , \12174 );
not \U$19552 ( \19895 , \19894 );
or \U$19553 ( \19896 , \19893 , \19895 );
nand \U$19554 ( \19897 , \12174 , \3057 );
nand \U$19555 ( \19898 , \19896 , \19897 );
nand \U$19556 ( \19899 , \19898 , \832 );
nand \U$19557 ( \19900 , \19892 , \19899 );
or \U$19558 ( \19901 , \19889 , \19900 );
not \U$19559 ( \19902 , \853 );
not \U$19560 ( \19903 , RIbb2eda0_19);
not \U$19561 ( \19904 , \17294 );
or \U$19562 ( \19905 , \19903 , \19904 );
not \U$19563 ( \19906 , RIbb2eda0_19);
nand \U$19564 ( \19907 , \19906 , \11142 );
nand \U$19565 ( \19908 , \19905 , \19907 );
not \U$19566 ( \19909 , \19908 );
or \U$19567 ( \19910 , \19902 , \19909 );
nand \U$19568 ( \19911 , \18806 , \854 );
nand \U$19569 ( \19912 , \19910 , \19911 );
nand \U$19570 ( \19913 , \19901 , \19912 );
nand \U$19571 ( \19914 , \19889 , \19900 );
nand \U$19572 ( \19915 , \19913 , \19914 );
and \U$19573 ( \19916 , \19880 , \19915 );
and \U$19574 ( \19917 , \19795 , \19879 );
or \U$19575 ( \19918 , \19916 , \19917 );
and \U$19576 ( \19919 , \19759 , \19918 );
and \U$19577 ( \19920 , \19647 , \19758 );
or \U$19578 ( \19921 , \19919 , \19920 );
nand \U$19579 ( \19922 , \19595 , \19921 );
not \U$19580 ( \19923 , \19487 );
nand \U$19581 ( \19924 , \19923 , \19592 );
nand \U$19582 ( \19925 , \19922 , \19924 );
xor \U$19583 ( \19926 , \19016 , \18763 );
xnor \U$19584 ( \19927 , \19926 , \19037 );
xor \U$19585 ( \19928 , \19925 , \19927 );
xor \U$19586 ( \19929 , \19296 , \19340 );
xor \U$19587 ( \19930 , \19929 , \19343 );
and \U$19588 ( \19931 , \19928 , \19930 );
and \U$19589 ( \19932 , \19925 , \19927 );
or \U$19590 ( \19933 , \19931 , \19932 );
not \U$19591 ( \19934 , \19043 );
not \U$19592 ( \19935 , \18757 );
or \U$19593 ( \19936 , \19934 , \19935 );
or \U$19594 ( \19937 , \19043 , \18757 );
nand \U$19595 ( \19938 , \19936 , \19937 );
and \U$19596 ( \19939 , \19938 , \19169 );
not \U$19597 ( \19940 , \19938 );
not \U$19598 ( \19941 , \19169 );
and \U$19599 ( \19942 , \19940 , \19941 );
nor \U$19600 ( \19943 , \19939 , \19942 );
xor \U$19601 ( \19944 , \19933 , \19943 );
xor \U$19602 ( \19945 , \19346 , \19476 );
xor \U$19603 ( \19946 , \19945 , \19479 );
and \U$19604 ( \19947 , \19944 , \19946 );
and \U$19605 ( \19948 , \19933 , \19943 );
or \U$19606 ( \19949 , \19947 , \19948 );
xnor \U$19607 ( \19950 , \19484 , \19949 );
xor \U$19608 ( \19951 , \19933 , \19943 );
xor \U$19609 ( \19952 , \19951 , \19946 );
xor \U$19610 ( \19953 , \17351 , \17503 );
xor \U$19611 ( \19954 , \19953 , \17638 );
xor \U$19612 ( \19955 , \18852 , \18886 );
xor \U$19613 ( \19956 , \19955 , \18961 );
not \U$19614 ( \19957 , \19956 );
xor \U$19615 ( \19958 , \17501 , \17450 );
xor \U$19616 ( \19959 , \19958 , \17395 );
not \U$19617 ( \19960 , \19959 );
or \U$19618 ( \19961 , \19957 , \19960 );
or \U$19619 ( \19962 , \19959 , \19956 );
xor \U$19620 ( \19963 , \17583 , \17632 );
xor \U$19621 ( \19964 , \19963 , \17635 );
nand \U$19622 ( \19965 , \19962 , \19964 );
nand \U$19623 ( \19966 , \19961 , \19965 );
xor \U$19624 ( \19967 , \19954 , \19966 );
not \U$19625 ( \19968 , \19331 );
not \U$19626 ( \19969 , \19323 );
or \U$19627 ( \19970 , \19968 , \19969 );
or \U$19628 ( \19971 , \19323 , \19331 );
nand \U$19629 ( \19972 , \19970 , \19971 );
and \U$19630 ( \19973 , \19972 , \19319 );
not \U$19631 ( \19974 , \19972 );
and \U$19632 ( \19975 , \19974 , \19320 );
nor \U$19633 ( \19976 , \19973 , \19975 );
not \U$19634 ( \19977 , \19976 );
xor \U$19635 ( \19978 , \19309 , \19305 );
xnor \U$19636 ( \19979 , \19978 , \19314 );
or \U$19637 ( \19980 , \19977 , \19979 );
xor \U$19638 ( \19981 , \19597 , \19619 );
xor \U$19639 ( \19982 , \19981 , \19644 );
not \U$19640 ( \19983 , \19982 );
xor \U$19641 ( \19984 , \17548 , \17565 );
xor \U$19642 ( \19985 , \19984 , \17580 );
not \U$19643 ( \19986 , \19985 );
or \U$19644 ( \19987 , \19983 , \19986 );
or \U$19645 ( \19988 , \19982 , \19985 );
not \U$19646 ( \19989 , \2939 );
not \U$19647 ( \19990 , RIbb2e800_31);
not \U$19648 ( \19991 , \6231 );
or \U$19649 ( \19992 , \19990 , \19991 );
not \U$19650 ( \19993 , RIbb2e800_31);
nand \U$19651 ( \19994 , \19993 , \8387 );
nand \U$19652 ( \19995 , \19992 , \19994 );
not \U$19653 ( \19996 , \19995 );
or \U$19654 ( \19997 , \19989 , \19996 );
nand \U$19655 ( \19998 , \19887 , \2941 );
nand \U$19656 ( \19999 , \19997 , \19998 );
buf \U$19657 ( \20000 , \19999 );
not \U$19658 ( \20001 , \20000 );
not \U$19659 ( \20002 , \2922 );
not \U$19660 ( \20003 , RIbb2e8f0_29);
not \U$19661 ( \20004 , \8338 );
or \U$19662 ( \20005 , \20003 , \20004 );
not \U$19663 ( \20006 , \13875 );
nand \U$19664 ( \20007 , \20006 , \3440 );
nand \U$19665 ( \20008 , \20005 , \20007 );
not \U$19666 ( \20009 , \20008 );
or \U$19667 ( \20010 , \20002 , \20009 );
nand \U$19668 ( \20011 , \19637 , \2925 );
nand \U$19669 ( \20012 , \20010 , \20011 );
not \U$19670 ( \20013 , \20012 );
or \U$19671 ( \20014 , \20001 , \20013 );
or \U$19672 ( \20015 , \20012 , \20000 );
not \U$19673 ( \20016 , \836 );
not \U$19674 ( \20017 , \19898 );
or \U$19675 ( \20018 , \20016 , \20017 );
not \U$19676 ( \20019 , RIbb2ee90_17);
not \U$19677 ( \20020 , \16865 );
or \U$19678 ( \20021 , \20019 , \20020 );
nand \U$19679 ( \20022 , \14635 , \822 );
nand \U$19680 ( \20023 , \20021 , \20022 );
nand \U$19681 ( \20024 , \20023 , \832 );
nand \U$19682 ( \20025 , \20018 , \20024 );
nand \U$19683 ( \20026 , \20015 , \20025 );
nand \U$19684 ( \20027 , \20014 , \20026 );
not \U$19685 ( \20028 , \20027 );
not \U$19686 ( \20029 , \854 );
not \U$19687 ( \20030 , \19908 );
or \U$19688 ( \20031 , \20029 , \20030 );
not \U$19689 ( \20032 , RIbb2eda0_19);
not \U$19690 ( \20033 , \17440 );
or \U$19691 ( \20034 , \20032 , \20033 );
not \U$19692 ( \20035 , RIbb2eda0_19);
nand \U$19693 ( \20036 , \20035 , \11578 );
nand \U$19694 ( \20037 , \20034 , \20036 );
nand \U$19695 ( \20038 , \20037 , \853 );
nand \U$19696 ( \20039 , \20031 , \20038 );
not \U$19697 ( \20040 , \3406 );
not \U$19698 ( \20041 , RIbb2ebc0_23);
not \U$19699 ( \20042 , \14550 );
or \U$19700 ( \20043 , \20041 , \20042 );
not \U$19701 ( \20044 , \9840 );
not \U$19702 ( \20045 , \20044 );
nand \U$19703 ( \20046 , \20045 , \3388 );
nand \U$19704 ( \20047 , \20043 , \20046 );
not \U$19705 ( \20048 , \20047 );
or \U$19706 ( \20049 , \20040 , \20048 );
nand \U$19707 ( \20050 , \19767 , \3383 );
nand \U$19708 ( \20051 , \20049 , \20050 );
xor \U$19709 ( \20052 , \20039 , \20051 );
not \U$19710 ( \20053 , \2078 );
not \U$19711 ( \20054 , \19789 );
or \U$19712 ( \20055 , \20053 , \20054 );
not \U$19713 ( \20056 , RIbb2ecb0_21);
not \U$19714 ( \20057 , \14563 );
or \U$19715 ( \20058 , \20056 , \20057 );
nand \U$19716 ( \20059 , \10764 , \2254 );
nand \U$19717 ( \20060 , \20058 , \20059 );
nand \U$19718 ( \20061 , \20060 , \2077 );
nand \U$19719 ( \20062 , \20055 , \20061 );
and \U$19720 ( \20063 , \20052 , \20062 );
and \U$19721 ( \20064 , \20039 , \20051 );
or \U$19722 ( \20065 , \20063 , \20064 );
not \U$19723 ( \20066 , \20065 );
or \U$19724 ( \20067 , \20028 , \20066 );
not \U$19725 ( \20068 , \20065 );
not \U$19726 ( \20069 , \20068 );
not \U$19727 ( \20070 , \20027 );
not \U$19728 ( \20071 , \20070 );
or \U$19729 ( \20072 , \20069 , \20071 );
not \U$19730 ( \20073 , \1737 );
not \U$19731 ( \20074 , \19833 );
or \U$19732 ( \20075 , \20073 , \20074 );
not \U$19733 ( \20076 , RIbb2f340_7);
not \U$19734 ( \20077 , \16710 );
or \U$19735 ( \20078 , \20076 , \20077 );
nand \U$19736 ( \20079 , \16553 , \1692 );
nand \U$19737 ( \20080 , \20078 , \20079 );
nand \U$19738 ( \20081 , \20080 , \1701 );
nand \U$19739 ( \20082 , \20075 , \20081 );
and \U$19740 ( \20083 , \17506 , \1253 );
not \U$19741 ( \20084 , \17506 );
and \U$19742 ( \20085 , \20084 , \1243 );
nor \U$19743 ( \20086 , \20083 , \20085 );
not \U$19744 ( \20087 , \20086 );
not \U$19745 ( \20088 , \1264 );
or \U$19746 ( \20089 , \20087 , \20088 );
nand \U$19747 ( \20090 , \19843 , \1261 );
nand \U$19748 ( \20091 , \20089 , \20090 );
xor \U$19749 ( \20092 , \20082 , \20091 );
not \U$19750 ( \20093 , \1570 );
not \U$19751 ( \20094 , \19857 );
or \U$19752 ( \20095 , \20093 , \20094 );
not \U$19753 ( \20096 , RIbb2f250_9);
not \U$19754 ( \20097 , \16747 );
or \U$19755 ( \20098 , \20096 , \20097 );
nand \U$19756 ( \20099 , \19077 , \1554 );
nand \U$19757 ( \20100 , \20098 , \20099 );
nand \U$19758 ( \20101 , \20100 , \1533 );
nand \U$19759 ( \20102 , \20095 , \20101 );
and \U$19760 ( \20103 , \20092 , \20102 );
and \U$19761 ( \20104 , \20082 , \20091 );
or \U$19762 ( \20105 , \20103 , \20104 );
not \U$19763 ( \20106 , \2963 );
not \U$19764 ( \20107 , \19775 );
or \U$19765 ( \20108 , \20106 , \20107 );
xor \U$19766 ( \20109 , \8630 , RIbb2ead0_25);
nand \U$19767 ( \20110 , \20109 , \2980 );
nand \U$19768 ( \20111 , \20108 , \20110 );
xor \U$19769 ( \20112 , \20105 , \20111 );
not \U$19770 ( \20113 , \3465 );
not \U$19771 ( \20114 , \19872 );
or \U$19772 ( \20115 , \20113 , \20114 );
not \U$19773 ( \20116 , RIbb2e9e0_27);
not \U$19774 ( \20117 , \17811 );
or \U$19775 ( \20118 , \20116 , \20117 );
nand \U$19776 ( \20119 , \14673 , \4598 );
nand \U$19777 ( \20120 , \20118 , \20119 );
nand \U$19778 ( \20121 , \20120 , \3445 );
nand \U$19779 ( \20122 , \20115 , \20121 );
and \U$19780 ( \20123 , \20112 , \20122 );
and \U$19781 ( \20124 , \20105 , \20111 );
or \U$19782 ( \20125 , \20123 , \20124 );
nand \U$19783 ( \20126 , \20072 , \20125 );
nand \U$19784 ( \20127 , \20067 , \20126 );
nand \U$19785 ( \20128 , \19988 , \20127 );
nand \U$19786 ( \20129 , \19987 , \20128 );
nand \U$19787 ( \20130 , \19980 , \20129 );
nand \U$19788 ( \20131 , \19977 , \19979 );
nand \U$19789 ( \20132 , \20130 , \20131 );
and \U$19790 ( \20133 , \19967 , \20132 );
and \U$19791 ( \20134 , \19954 , \19966 );
or \U$19792 ( \20135 , \20133 , \20134 );
xor \U$19793 ( \20136 , \19020 , \19031 );
xor \U$19794 ( \20137 , \20136 , \19034 );
xor \U$19795 ( \20138 , \19338 , \19316 );
xor \U$19796 ( \20139 , \20138 , \19333 );
xor \U$19797 ( \20140 , \20137 , \20139 );
not \U$19798 ( \20141 , \19461 );
not \U$19799 ( \20142 , \19358 );
or \U$19800 ( \20143 , \20141 , \20142 );
or \U$19801 ( \20144 , \19461 , \19358 );
nand \U$19802 ( \20145 , \20143 , \20144 );
and \U$19803 ( \20146 , \20145 , \19458 );
not \U$19804 ( \20147 , \20145 );
not \U$19805 ( \20148 , \19458 );
and \U$19806 ( \20149 , \20147 , \20148 );
nor \U$19807 ( \20150 , \20146 , \20149 );
and \U$19808 ( \20151 , \20140 , \20150 );
and \U$19809 ( \20152 , \20137 , \20139 );
or \U$19810 ( \20153 , \20151 , \20152 );
xor \U$19811 ( \20154 , \20135 , \20153 );
xor \U$19812 ( \20155 , \19348 , \19465 );
xor \U$19813 ( \20156 , \20155 , \19473 );
and \U$19814 ( \20157 , \20154 , \20156 );
and \U$19815 ( \20158 , \20135 , \20153 );
or \U$19816 ( \20159 , \20157 , \20158 );
or \U$19817 ( \20160 , \19952 , \20159 );
xor \U$19818 ( \20161 , \19921 , \19486 );
xor \U$19819 ( \20162 , \20161 , \19593 );
xor \U$19820 ( \20163 , \19647 , \19758 );
xor \U$19821 ( \20164 , \20163 , \19918 );
xor \U$19822 ( \20165 , \19912 , \19900 );
xnor \U$19823 ( \20166 , \20165 , \19889 );
not \U$19824 ( \20167 , \20166 );
not \U$19825 ( \20168 , \20167 );
not \U$19826 ( \20169 , \16271 );
and \U$19827 ( \20170 , RIbb2dae0_59, \1036 );
not \U$19828 ( \20171 , RIbb2dae0_59);
and \U$19829 ( \20172 , \20171 , \1559 );
nor \U$19830 ( \20173 , \20170 , \20172 );
not \U$19831 ( \20174 , \20173 );
or \U$19832 ( \20175 , \20169 , \20174 );
nand \U$19833 ( \20176 , \19689 , \16257 );
nand \U$19834 ( \20177 , \20175 , \20176 );
not \U$19835 ( \20178 , \20177 );
not \U$19836 ( \20179 , \20178 );
not \U$19837 ( \20180 , \19698 );
not \U$19838 ( \20181 , \8352 );
and \U$19839 ( \20182 , \20180 , \20181 );
not \U$19840 ( \20183 , RIbb2e350_41);
not \U$19841 ( \20184 , \3200 );
or \U$19842 ( \20185 , \20183 , \20184 );
nand \U$19843 ( \20186 , \3199 , \13400 );
nand \U$19844 ( \20187 , \20185 , \20186 );
and \U$19845 ( \20188 , \20187 , \8361 );
nor \U$19846 ( \20189 , \20182 , \20188 );
not \U$19847 ( \20190 , \20189 );
or \U$19848 ( \20191 , \20179 , \20190 );
not \U$19849 ( \20192 , \9098 );
and \U$19850 ( \20193 , RIbb2e260_43, \6107 );
not \U$19851 ( \20194 , RIbb2e260_43);
and \U$19852 ( \20195 , \20194 , \3166 );
or \U$19853 ( \20196 , \20193 , \20195 );
not \U$19854 ( \20197 , \20196 );
or \U$19855 ( \20198 , \20192 , \20197 );
nand \U$19856 ( \20199 , \19384 , \10451 );
nand \U$19857 ( \20200 , \20198 , \20199 );
nand \U$19858 ( \20201 , \20191 , \20200 );
not \U$19859 ( \20202 , \20189 );
nand \U$19860 ( \20203 , \20202 , \20177 );
nand \U$19861 ( \20204 , \20201 , \20203 );
not \U$19862 ( \20205 , \20204 );
or \U$19863 ( \20206 , \20168 , \20205 );
or \U$19864 ( \20207 , \20204 , \20167 );
xor \U$19865 ( \20208 , \19837 , \19848 );
xor \U$19866 ( \20209 , \20208 , \19859 );
not \U$19867 ( \20210 , \12692 );
not \U$19868 ( \20211 , \19652 );
or \U$19869 ( \20212 , \20210 , \20211 );
and \U$19870 ( \20213 , RIbb2dea0_51, \1169 );
not \U$19871 ( \20214 , RIbb2dea0_51);
not \U$19872 ( \20215 , \1169 );
and \U$19873 ( \20216 , \20214 , \20215 );
nor \U$19874 ( \20217 , \20213 , \20216 );
nand \U$19875 ( \20218 , \20217 , \14067 );
nand \U$19876 ( \20219 , \20212 , \20218 );
xor \U$19877 ( \20220 , \20209 , \20219 );
not \U$19878 ( \20221 , \6242 );
not \U$19879 ( \20222 , \19678 );
or \U$19880 ( \20223 , \20221 , \20222 );
not \U$19881 ( \20224 , RIbb2e530_37);
not \U$19882 ( \20225 , \17910 );
or \U$19883 ( \20226 , \20224 , \20225 );
nand \U$19884 ( \20227 , \3044 , \6246 );
nand \U$19885 ( \20228 , \20226 , \20227 );
nand \U$19886 ( \20229 , \20228 , \6251 );
nand \U$19887 ( \20230 , \20223 , \20229 );
and \U$19888 ( \20231 , \20220 , \20230 );
and \U$19889 ( \20232 , \20209 , \20219 );
or \U$19890 ( \20233 , \20231 , \20232 );
nand \U$19891 ( \20234 , \20207 , \20233 );
nand \U$19892 ( \20235 , \20206 , \20234 );
xor \U$19893 ( \20236 , \19795 , \19879 );
xor \U$19894 ( \20237 , \20236 , \19915 );
xor \U$19895 ( \20238 , \20235 , \20237 );
not \U$19896 ( \20239 , \10599 );
and \U$19897 ( \20240 , \2222 , \9094 );
not \U$19898 ( \20241 , \2222 );
and \U$19899 ( \20242 , \20241 , RIbb2e170_45);
or \U$19900 ( \20243 , \20240 , \20242 );
not \U$19901 ( \20244 , \20243 );
or \U$19902 ( \20245 , \20239 , \20244 );
nand \U$19903 ( \20246 , \19396 , \10119 );
nand \U$19904 ( \20247 , \20245 , \20246 );
not \U$19905 ( \20248 , RIbb2d888_64);
not \U$19906 ( \20249 , \19723 );
or \U$19907 ( \20250 , \20248 , \20249 );
not \U$19908 ( \20251 , RIbb2d900_63);
not \U$19909 ( \20252 , \1473 );
or \U$19910 ( \20253 , \20251 , \20252 );
not \U$19911 ( \20254 , RIbb2d900_63);
nand \U$19912 ( \20255 , \20254 , \1472 );
nand \U$19913 ( \20256 , \20253 , \20255 );
nand \U$19914 ( \20257 , \20256 , \17275 );
nand \U$19915 ( \20258 , \20250 , \20257 );
nor \U$19916 ( \20259 , \20247 , \20258 );
not \U$19917 ( \20260 , \14613 );
and \U$19918 ( \20261 , RIbb2dcc0_55, \1642 );
not \U$19919 ( \20262 , RIbb2dcc0_55);
and \U$19920 ( \20263 , \20262 , \3238 );
nor \U$19921 ( \20264 , \20261 , \20263 );
not \U$19922 ( \20265 , \20264 );
or \U$19923 ( \20266 , \20260 , \20265 );
nand \U$19924 ( \20267 , \19375 , \15181 );
nand \U$19925 ( \20268 , \20266 , \20267 );
not \U$19926 ( \20269 , \20268 );
or \U$19927 ( \20270 , \20259 , \20269 );
nand \U$19928 ( \20271 , \20258 , \20247 );
nand \U$19929 ( \20272 , \20270 , \20271 );
not \U$19930 ( \20273 , \8445 );
not \U$19931 ( \20274 , RIbb2e440_39);
not \U$19932 ( \20275 , \16898 );
or \U$19933 ( \20276 , \20274 , \20275 );
not \U$19934 ( \20277 , RIbb2e440_39);
nand \U$19935 ( \20278 , \20277 , \3653 );
nand \U$19936 ( \20279 , \20276 , \20278 );
not \U$19937 ( \20280 , \20279 );
or \U$19938 ( \20281 , \20273 , \20280 );
nand \U$19939 ( \20282 , \19664 , \8450 );
nand \U$19940 ( \20283 , \20281 , \20282 );
not \U$19941 ( \20284 , \20283 );
not \U$19942 ( \20285 , \5845 );
not \U$19943 ( \20286 , \19530 );
or \U$19944 ( \20287 , \20285 , \20286 );
not \U$19945 ( \20288 , RIbb2e620_35);
not \U$19946 ( \20289 , \12577 );
or \U$19947 ( \20290 , \20288 , \20289 );
nand \U$19948 ( \20291 , \13750 , \6002 );
nand \U$19949 ( \20292 , \20290 , \20291 );
nand \U$19950 ( \20293 , \20292 , \4712 );
nand \U$19951 ( \20294 , \20287 , \20293 );
not \U$19952 ( \20295 , \20294 );
or \U$19953 ( \20296 , \20284 , \20295 );
or \U$19954 ( \20297 , \20294 , \20283 );
not \U$19955 ( \20298 , \15688 );
not \U$19956 ( \20299 , \19708 );
or \U$19957 ( \20300 , \20298 , \20299 );
not \U$19958 ( \20301 , RIbb2ddb0_53);
not \U$19959 ( \20302 , \1110 );
or \U$19960 ( \20303 , \20301 , \20302 );
nand \U$19961 ( \20304 , \13463 , \1109 );
nand \U$19962 ( \20305 , \20303 , \20304 );
nand \U$19963 ( \20306 , \20305 , \17562 );
nand \U$19964 ( \20307 , \20300 , \20306 );
nand \U$19965 ( \20308 , \20297 , \20307 );
nand \U$19966 ( \20309 , \20296 , \20308 );
nand \U$19967 ( \20310 , \20272 , \20309 );
or \U$19968 ( \20311 , \20272 , \20309 );
not \U$19969 ( \20312 , \15738 );
not \U$19970 ( \20313 , \19420 );
or \U$19971 ( \20314 , \20312 , \20313 );
not \U$19972 ( \20315 , RIbb2dbd0_57);
not \U$19973 ( \20316 , \14819 );
or \U$19974 ( \20317 , \20315 , \20316 );
nand \U$19975 ( \20318 , \14818 , \17097 );
nand \U$19976 ( \20319 , \20317 , \20318 );
nand \U$19977 ( \20320 , \20319 , \16674 );
nand \U$19978 ( \20321 , \20314 , \20320 );
not \U$19979 ( \20322 , \20321 );
not \U$19980 ( \20323 , \11176 );
not \U$19981 ( \20324 , RIbb2e080_47);
not \U$19982 ( \20325 , \1851 );
not \U$19983 ( \20326 , \20325 );
or \U$19984 ( \20327 , \20324 , \20326 );
nand \U$19985 ( \20328 , \1851 , \10113 );
nand \U$19986 ( \20329 , \20327 , \20328 );
not \U$19987 ( \20330 , \20329 );
or \U$19988 ( \20331 , \20323 , \20330 );
nand \U$19989 ( \20332 , \19737 , \11177 );
nand \U$19990 ( \20333 , \20331 , \20332 );
not \U$19991 ( \20334 , \20333 );
or \U$19992 ( \20335 , \20322 , \20334 );
not \U$19993 ( \20336 , \20333 );
not \U$19994 ( \20337 , \20336 );
not \U$19995 ( \20338 , \20321 );
not \U$19996 ( \20339 , \20338 );
or \U$19997 ( \20340 , \20337 , \20339 );
not \U$19998 ( \20341 , \16533 );
not \U$19999 ( \20342 , \19751 );
or \U$20000 ( \20343 , \20341 , \20342 );
not \U$20001 ( \20344 , \19746 );
not \U$20002 ( \20345 , \950 );
or \U$20003 ( \20346 , \20344 , \20345 );
or \U$20004 ( \20347 , \950 , \19746 );
nand \U$20005 ( \20348 , \20346 , \20347 );
nand \U$20006 ( \20349 , \20348 , \16541 );
nand \U$20007 ( \20350 , \20343 , \20349 );
nand \U$20008 ( \20351 , \20340 , \20350 );
nand \U$20009 ( \20352 , \20335 , \20351 );
nand \U$20010 ( \20353 , \20311 , \20352 );
nand \U$20011 ( \20354 , \20310 , \20353 );
and \U$20012 ( \20355 , \20238 , \20354 );
and \U$20013 ( \20356 , \20235 , \20237 );
or \U$20014 ( \20357 , \20355 , \20356 );
xor \U$20015 ( \20358 , \20164 , \20357 );
xor \U$20016 ( \20359 , \19360 , \19406 );
xor \U$20017 ( \20360 , \20359 , \19455 );
and \U$20018 ( \20361 , \20358 , \20360 );
and \U$20019 ( \20362 , \20164 , \20357 );
or \U$20020 ( \20363 , \20361 , \20362 );
not \U$20021 ( \20364 , \20363 );
nand \U$20022 ( \20365 , \20162 , \20364 );
not \U$20023 ( \20366 , \20365 );
xor \U$20024 ( \20367 , \19954 , \19966 );
xor \U$20025 ( \20368 , \20367 , \20132 );
not \U$20026 ( \20369 , \20368 );
or \U$20027 ( \20370 , \20366 , \20369 );
not \U$20028 ( \20371 , \20162 );
nand \U$20029 ( \20372 , \20371 , \20363 );
nand \U$20030 ( \20373 , \20370 , \20372 );
xor \U$20031 ( \20374 , \19590 , \19508 );
xnor \U$20032 ( \20375 , \20374 , \19511 );
xor \U$20033 ( \20376 , \19607 , \19613 );
xor \U$20034 ( \20377 , \20376 , \19617 );
xor \U$20035 ( \20378 , \19625 , \19630 );
xor \U$20036 ( \20379 , \20378 , \19641 );
xor \U$20037 ( \20380 , \20377 , \20379 );
xor \U$20038 ( \20381 , \19805 , \19806 );
xor \U$20039 ( \20382 , \20381 , \19823 );
not \U$20040 ( \20383 , \4075 );
not \U$20041 ( \20384 , \19433 );
or \U$20042 ( \20385 , \20383 , \20384 );
not \U$20043 ( \20386 , RIbb2e710_33);
not \U$20044 ( \20387 , \4390 );
not \U$20045 ( \20388 , \20387 );
or \U$20046 ( \20389 , \20386 , \20388 );
not \U$20047 ( \20390 , \13559 );
nand \U$20048 ( \20391 , \20390 , \7390 );
nand \U$20049 ( \20392 , \20389 , \20391 );
nand \U$20050 ( \20393 , \20392 , \3886 );
nand \U$20051 ( \20394 , \20385 , \20393 );
xor \U$20052 ( \20395 , \20382 , \20394 );
not \U$20053 ( \20396 , \13295 );
not \U$20054 ( \20397 , RIbb2df90_49);
not \U$20055 ( \20398 , \1420 );
or \U$20056 ( \20399 , \20397 , \20398 );
nand \U$20057 ( \20400 , \3821 , \12278 );
nand \U$20058 ( \20401 , \20399 , \20400 );
not \U$20059 ( \20402 , \20401 );
or \U$20060 ( \20403 , \20396 , \20402 );
nand \U$20061 ( \20404 , \19442 , \12169 );
nand \U$20062 ( \20405 , \20403 , \20404 );
and \U$20063 ( \20406 , \20395 , \20405 );
and \U$20064 ( \20407 , \20382 , \20394 );
or \U$20065 ( \20408 , \20406 , \20407 );
and \U$20066 ( \20409 , \20380 , \20408 );
and \U$20067 ( \20410 , \20377 , \20379 );
or \U$20068 ( \20411 , \20409 , \20410 );
xor \U$20069 ( \20412 , \19755 , \19715 );
xor \U$20070 ( \20413 , \20412 , \19682 );
xor \U$20071 ( \20414 , \20411 , \20413 );
xor \U$20072 ( \20415 , \19666 , \19680 );
buf \U$20073 ( \20416 , \19656 );
and \U$20074 ( \20417 , \20415 , \20416 );
not \U$20075 ( \20418 , \20415 );
not \U$20076 ( \20419 , \20416 );
and \U$20077 ( \20420 , \20418 , \20419 );
nor \U$20078 ( \20421 , \20417 , \20420 );
not \U$20079 ( \20422 , \20421 );
not \U$20080 ( \20423 , \20422 );
xor \U$20081 ( \20424 , \19446 , \19424 );
xnor \U$20082 ( \20425 , \20424 , \19435 );
not \U$20083 ( \20426 , \20425 );
or \U$20084 ( \20427 , \20423 , \20426 );
xor \U$20085 ( \20428 , \19753 , \19739 );
not \U$20086 ( \20429 , \19727 );
and \U$20087 ( \20430 , \20428 , \20429 );
not \U$20088 ( \20431 , \20428 );
and \U$20089 ( \20432 , \20431 , \19727 );
nor \U$20090 ( \20433 , \20430 , \20432 );
not \U$20091 ( \20434 , \20433 );
nand \U$20092 ( \20435 , \20427 , \20434 );
not \U$20093 ( \20436 , \20422 );
not \U$20094 ( \20437 , \20425 );
nand \U$20095 ( \20438 , \20436 , \20437 );
nand \U$20096 ( \20439 , \20435 , \20438 );
and \U$20097 ( \20440 , \20414 , \20439 );
and \U$20098 ( \20441 , \20411 , \20413 );
or \U$20099 ( \20442 , \20440 , \20441 );
not \U$20100 ( \20443 , \20442 );
nand \U$20101 ( \20444 , \20375 , \20443 );
not \U$20102 ( \20445 , \20444 );
xor \U$20103 ( \20446 , \18906 , \19413 );
xor \U$20104 ( \20447 , \19409 , \18957 );
xnor \U$20105 ( \20448 , \20446 , \20447 );
and \U$20106 ( \20449 , \20448 , \19453 );
not \U$20107 ( \20450 , \20448 );
and \U$20108 ( \20451 , \20450 , \19449 );
nor \U$20109 ( \20452 , \20449 , \20451 );
not \U$20110 ( \20453 , \20452 );
xor \U$20111 ( \20454 , \19365 , \19401 );
xnor \U$20112 ( \20455 , \20454 , \19404 );
or \U$20113 ( \20456 , \20453 , \20455 );
not \U$20114 ( \20457 , \20453 );
not \U$20115 ( \20458 , \20455 );
or \U$20116 ( \20459 , \20457 , \20458 );
xor \U$20117 ( \20460 , \19779 , \19769 );
and \U$20118 ( \20461 , \20460 , \19792 );
not \U$20119 ( \20462 , \20460 );
and \U$20120 ( \20463 , \20462 , \19791 );
nor \U$20121 ( \20464 , \20461 , \20463 );
not \U$20122 ( \20465 , \20464 );
not \U$20123 ( \20466 , \20465 );
xor \U$20124 ( \20467 , \19584 , \19581 );
xnor \U$20125 ( \20468 , \20467 , \19532 );
not \U$20126 ( \20469 , \20468 );
not \U$20127 ( \20470 , \20469 );
or \U$20128 ( \20471 , \20466 , \20470 );
not \U$20129 ( \20472 , \20464 );
not \U$20130 ( \20473 , \20468 );
or \U$20131 ( \20474 , \20472 , \20473 );
xor \U$20132 ( \20475 , \19826 , \19862 );
xor \U$20133 ( \20476 , \20475 , \19876 );
nand \U$20134 ( \20477 , \20474 , \20476 );
nand \U$20135 ( \20478 , \20471 , \20477 );
nand \U$20136 ( \20479 , \20459 , \20478 );
nand \U$20137 ( \20480 , \20456 , \20479 );
not \U$20138 ( \20481 , \20480 );
or \U$20139 ( \20482 , \20445 , \20481 );
not \U$20140 ( \20483 , \20375 );
nand \U$20141 ( \20484 , \20483 , \20442 );
nand \U$20142 ( \20485 , \20482 , \20484 );
xor \U$20143 ( \20486 , \19956 , \19964 );
xnor \U$20144 ( \20487 , \20486 , \19959 );
not \U$20145 ( \20488 , \20487 );
not \U$20146 ( \20489 , \20488 );
xor \U$20147 ( \20490 , \19519 , \19516 );
not \U$20148 ( \20491 , \19588 );
and \U$20149 ( \20492 , \20490 , \20491 );
not \U$20150 ( \20493 , \20490 );
and \U$20151 ( \20494 , \20493 , \19588 );
nor \U$20152 ( \20495 , \20492 , \20494 );
not \U$20153 ( \20496 , \20495 );
not \U$20154 ( \20497 , \19506 );
not \U$20155 ( \20498 , \19494 );
or \U$20156 ( \20499 , \20497 , \20498 );
or \U$20157 ( \20500 , \19506 , \19494 );
nand \U$20158 ( \20501 , \20499 , \20500 );
and \U$20159 ( \20502 , \20501 , \19499 );
not \U$20160 ( \20503 , \20501 );
and \U$20161 ( \20504 , \20503 , \19498 );
nor \U$20162 ( \20505 , \20502 , \20504 );
nand \U$20163 ( \20506 , \20496 , \20505 );
not \U$20164 ( \20507 , \20505 );
not \U$20165 ( \20508 , \20507 );
not \U$20166 ( \20509 , \20495 );
or \U$20167 ( \20510 , \20508 , \20509 );
xor \U$20168 ( \20511 , \19547 , \19563 );
xor \U$20169 ( \20512 , \20511 , \19579 );
not \U$20170 ( \20513 , \1077 );
not \U$20171 ( \20514 , \19554 );
or \U$20172 ( \20515 , \20513 , \20514 );
not \U$20173 ( \20516 , RIbb2f160_11);
not \U$20174 ( \20517 , \16567 );
or \U$20175 ( \20518 , \20516 , \20517 );
nand \U$20176 ( \20519 , \16562 , \1043 );
nand \U$20177 ( \20520 , \20518 , \20519 );
nand \U$20178 ( \20521 , \20520 , \1011 );
nand \U$20179 ( \20522 , \20515 , \20521 );
not \U$20180 ( \20523 , \1517 );
not \U$20181 ( \20524 , \19571 );
or \U$20182 ( \20525 , \20523 , \20524 );
and \U$20183 ( \20526 , RIbb2ef80_15, \15054 );
not \U$20184 ( \20527 , RIbb2ef80_15);
and \U$20185 ( \20528 , \20527 , \13545 );
or \U$20186 ( \20529 , \20526 , \20528 );
nand \U$20187 ( \20530 , \20529 , \1444 );
nand \U$20188 ( \20531 , \20525 , \20530 );
xor \U$20189 ( \20532 , \20522 , \20531 );
not \U$20190 ( \20533 , \832 );
not \U$20191 ( \20534 , RIbb2ee90_17);
not \U$20192 ( \20535 , \12348 );
or \U$20193 ( \20536 , \20534 , \20535 );
nand \U$20194 ( \20537 , \14839 , \2240 );
nand \U$20195 ( \20538 , \20536 , \20537 );
not \U$20196 ( \20539 , \20538 );
or \U$20197 ( \20540 , \20533 , \20539 );
nand \U$20198 ( \20541 , \20023 , \836 );
nand \U$20199 ( \20542 , \20540 , \20541 );
and \U$20200 ( \20543 , \20532 , \20542 );
and \U$20201 ( \20544 , \20522 , \20531 );
or \U$20202 ( \20545 , \20543 , \20544 );
or \U$20203 ( \20546 , \20512 , \20545 );
and \U$20204 ( \20547 , \17506 , \1261 );
not \U$20205 ( \20548 , \1146 );
not \U$20206 ( \20549 , \19820 );
or \U$20207 ( \20550 , \20548 , \20549 );
not \U$20208 ( \20551 , RIbb2f430_5);
not \U$20209 ( \20552 , \17517 );
not \U$20210 ( \20553 , \20552 );
or \U$20211 ( \20554 , \20551 , \20553 );
nand \U$20212 ( \20555 , \17517 , \1980 );
nand \U$20213 ( \20556 , \20554 , \20555 );
nand \U$20214 ( \20557 , \20556 , \1089 );
nand \U$20215 ( \20558 , \20550 , \20557 );
xor \U$20216 ( \20559 , \20547 , \20558 );
not \U$20217 ( \20560 , \1701 );
not \U$20218 ( \20561 , RIbb2f340_7);
not \U$20219 ( \20562 , \17750 );
or \U$20220 ( \20563 , \20561 , \20562 );
nand \U$20221 ( \20564 , \16703 , \1734 );
nand \U$20222 ( \20565 , \20563 , \20564 );
not \U$20223 ( \20566 , \20565 );
or \U$20224 ( \20567 , \20560 , \20566 );
nand \U$20225 ( \20568 , \20080 , \1737 );
nand \U$20226 ( \20569 , \20567 , \20568 );
and \U$20227 ( \20570 , \20559 , \20569 );
and \U$20228 ( \20571 , \20547 , \20558 );
or \U$20229 ( \20572 , \20570 , \20571 );
xor \U$20230 ( \20573 , \19812 , \19822 );
xor \U$20231 ( \20574 , \20572 , \20573 );
not \U$20232 ( \20575 , \915 );
not \U$20233 ( \20576 , RIbb2f070_13);
not \U$20234 ( \20577 , \14526 );
not \U$20235 ( \20578 , \20577 );
or \U$20236 ( \20579 , \20576 , \20578 );
not \U$20237 ( \20580 , \18353 );
nand \U$20238 ( \20581 , \20580 , \1656 );
nand \U$20239 ( \20582 , \20579 , \20581 );
not \U$20240 ( \20583 , \20582 );
or \U$20241 ( \20584 , \20575 , \20583 );
nand \U$20242 ( \20585 , \19538 , \998 );
nand \U$20243 ( \20586 , \20584 , \20585 );
and \U$20244 ( \20587 , \20574 , \20586 );
and \U$20245 ( \20588 , \20572 , \20573 );
or \U$20246 ( \20589 , \20587 , \20588 );
nand \U$20247 ( \20590 , \20546 , \20589 );
nand \U$20248 ( \20591 , \20512 , \20545 );
nand \U$20249 ( \20592 , \20590 , \20591 );
xor \U$20250 ( \20593 , \19691 , \19701 );
xor \U$20251 ( \20594 , \20593 , \19712 );
xor \U$20252 ( \20595 , \20592 , \20594 );
xor \U$20253 ( \20596 , \19377 , \19388 );
xor \U$20254 ( \20597 , \20596 , \19398 );
and \U$20255 ( \20598 , \20595 , \20597 );
and \U$20256 ( \20599 , \20592 , \20594 );
or \U$20257 ( \20600 , \20598 , \20599 );
nand \U$20258 ( \20601 , \20510 , \20600 );
nand \U$20259 ( \20602 , \20506 , \20601 );
not \U$20260 ( \20603 , \20602 );
or \U$20261 ( \20604 , \20489 , \20603 );
not \U$20262 ( \20605 , \20487 );
not \U$20263 ( \20606 , \20602 );
not \U$20264 ( \20607 , \20606 );
or \U$20265 ( \20608 , \20605 , \20607 );
xor \U$20266 ( \20609 , \20129 , \19976 );
xnor \U$20267 ( \20610 , \20609 , \19979 );
nand \U$20268 ( \20611 , \20608 , \20610 );
nand \U$20269 ( \20612 , \20604 , \20611 );
or \U$20270 ( \20613 , \20485 , \20612 );
xor \U$20271 ( \20614 , \20137 , \20139 );
xor \U$20272 ( \20615 , \20614 , \20150 );
nand \U$20273 ( \20616 , \20613 , \20615 );
nand \U$20274 ( \20617 , \20612 , \20485 );
nand \U$20275 ( \20618 , \20616 , \20617 );
xor \U$20276 ( \20619 , \20373 , \20618 );
xor \U$20277 ( \20620 , \19925 , \19927 );
xor \U$20278 ( \20621 , \20620 , \19930 );
and \U$20279 ( \20622 , \20619 , \20621 );
and \U$20280 ( \20623 , \20373 , \20618 );
or \U$20281 ( \20624 , \20622 , \20623 );
buf \U$20282 ( \20625 , \20624 );
nand \U$20283 ( \20626 , \20160 , \20625 );
nand \U$20284 ( \20627 , \19952 , \20159 );
nand \U$20285 ( \20628 , \20626 , \20627 );
not \U$20286 ( \20629 , \20628 );
nand \U$20287 ( \20630 , \19950 , \20629 );
not \U$20288 ( \20631 , \20630 );
xor \U$20289 ( \20632 , \20159 , \20624 );
xnor \U$20290 ( \20633 , \20632 , \19952 );
xor \U$20291 ( \20634 , \20373 , \20618 );
xor \U$20292 ( \20635 , \20634 , \20621 );
not \U$20293 ( \20636 , \20635 );
xor \U$20294 ( \20637 , \19982 , \19985 );
xnor \U$20295 ( \20638 , \20637 , \20127 );
not \U$20296 ( \20639 , \20638 );
not \U$20297 ( \20640 , \854 );
not \U$20298 ( \20641 , \20037 );
or \U$20299 ( \20642 , \20640 , \20641 );
and \U$20300 ( \20643 , \12174 , \1776 );
not \U$20301 ( \20644 , \12174 );
and \U$20302 ( \20645 , \20644 , RIbb2eda0_19);
or \U$20303 ( \20646 , \20643 , \20645 );
nand \U$20304 ( \20647 , \20646 , \853 );
nand \U$20305 ( \20648 , \20642 , \20647 );
buf \U$20306 ( \20649 , \20648 );
not \U$20307 ( \20650 , \20649 );
not \U$20308 ( \20651 , \20650 );
not \U$20309 ( \20652 , \3886 );
not \U$20310 ( \20653 , RIbb2e710_33);
not \U$20311 ( \20654 , \6197 );
or \U$20312 ( \20655 , \20653 , \20654 );
nand \U$20313 ( \20656 , \9020 , \13352 );
nand \U$20314 ( \20657 , \20655 , \20656 );
not \U$20315 ( \20658 , \20657 );
or \U$20316 ( \20659 , \20652 , \20658 );
nand \U$20317 ( \20660 , \20392 , \4075 );
nand \U$20318 ( \20661 , \20659 , \20660 );
not \U$20319 ( \20662 , \20661 );
not \U$20320 ( \20663 , \20662 );
or \U$20321 ( \20664 , \20651 , \20663 );
not \U$20322 ( \20665 , \2078 );
not \U$20323 ( \20666 , \20060 );
or \U$20324 ( \20667 , \20665 , \20666 );
not \U$20325 ( \20668 , RIbb2ecb0_21);
not \U$20326 ( \20669 , \17294 );
or \U$20327 ( \20670 , \20668 , \20669 );
nand \U$20328 ( \20671 , \11142 , \2067 );
nand \U$20329 ( \20672 , \20670 , \20671 );
nand \U$20330 ( \20673 , \20672 , \2077 );
nand \U$20331 ( \20674 , \20667 , \20673 );
nand \U$20332 ( \20675 , \20664 , \20674 );
nand \U$20333 ( \20676 , \20661 , \20649 );
nand \U$20334 ( \20677 , \20675 , \20676 );
not \U$20335 ( \20678 , \2980 );
not \U$20336 ( \20679 , RIbb2ead0_25);
not \U$20337 ( \20680 , \12819 );
or \U$20338 ( \20681 , \20679 , \20680 );
not \U$20339 ( \20682 , RIbb2ead0_25);
nand \U$20340 ( \20683 , \20682 , \9277 );
nand \U$20341 ( \20684 , \20681 , \20683 );
not \U$20342 ( \20685 , \20684 );
or \U$20343 ( \20686 , \20678 , \20685 );
nand \U$20344 ( \20687 , \20109 , \2963 );
nand \U$20345 ( \20688 , \20686 , \20687 );
not \U$20346 ( \20689 , \3465 );
not \U$20347 ( \20690 , \20120 );
or \U$20348 ( \20691 , \20689 , \20690 );
not \U$20349 ( \20692 , \8318 );
not \U$20350 ( \20693 , \20692 );
xor \U$20351 ( \20694 , RIbb2e9e0_27, \20693 );
nand \U$20352 ( \20695 , \20694 , \3445 );
nand \U$20353 ( \20696 , \20691 , \20695 );
xor \U$20354 ( \20697 , \20688 , \20696 );
not \U$20355 ( \20698 , \3383 );
not \U$20356 ( \20699 , \20047 );
or \U$20357 ( \20700 , \20698 , \20699 );
not \U$20358 ( \20701 , RIbb2ebc0_23);
not \U$20359 ( \20702 , \15105 );
or \U$20360 ( \20703 , \20701 , \20702 );
nand \U$20361 ( \20704 , \10300 , \3396 );
nand \U$20362 ( \20705 , \20703 , \20704 );
nand \U$20363 ( \20706 , \20705 , \3406 );
nand \U$20364 ( \20707 , \20700 , \20706 );
and \U$20365 ( \20708 , \20697 , \20707 );
and \U$20366 ( \20709 , \20688 , \20696 );
or \U$20367 ( \20710 , \20708 , \20709 );
nor \U$20368 ( \20711 , \20677 , \20710 );
not \U$20369 ( \20712 , \1077 );
not \U$20370 ( \20713 , \20520 );
or \U$20371 ( \20714 , \20712 , \20713 );
not \U$20372 ( \20715 , RIbb2f160_11);
not \U$20373 ( \20716 , \16576 );
not \U$20374 ( \20717 , \20716 );
or \U$20375 ( \20718 , \20715 , \20717 );
nand \U$20376 ( \20719 , \16575 , \1048 );
nand \U$20377 ( \20720 , \20718 , \20719 );
nand \U$20378 ( \20721 , \20720 , \1011 );
nand \U$20379 ( \20722 , \20714 , \20721 );
not \U$20380 ( \20723 , \20722 );
not \U$20381 ( \20724 , \1533 );
not \U$20382 ( \20725 , RIbb2f250_9);
not \U$20383 ( \20726 , \16728 );
or \U$20384 ( \20727 , \20725 , \20726 );
nand \U$20385 ( \20728 , \19831 , \5064 );
nand \U$20386 ( \20729 , \20727 , \20728 );
not \U$20387 ( \20730 , \20729 );
or \U$20388 ( \20731 , \20724 , \20730 );
nand \U$20389 ( \20732 , \1570 , \20100 );
nand \U$20390 ( \20733 , \20731 , \20732 );
not \U$20391 ( \20734 , \20733 );
nand \U$20392 ( \20735 , \20723 , \20734 );
or \U$20393 ( \20736 , RIbb2f3b8_6, RIbb2f340_7);
nand \U$20394 ( \20737 , \20736 , \17506 );
and \U$20395 ( \20738 , RIbb2f3b8_6, RIbb2f340_7);
nor \U$20396 ( \20739 , \20738 , \1647 );
nand \U$20397 ( \20740 , \20737 , \20739 );
not \U$20398 ( \20741 , \20740 );
not \U$20399 ( \20742 , \1146 );
not \U$20400 ( \20743 , \20556 );
or \U$20401 ( \20744 , \20742 , \20743 );
and \U$20402 ( \20745 , RIbb2f430_5, \17506 );
not \U$20403 ( \20746 , RIbb2f430_5);
not \U$20404 ( \20747 , \17506 );
and \U$20405 ( \20748 , \20746 , \20747 );
nor \U$20406 ( \20749 , \20745 , \20748 );
nand \U$20407 ( \20750 , \20749 , \1089 );
nand \U$20408 ( \20751 , \20744 , \20750 );
nand \U$20409 ( \20752 , \20741 , \20751 );
not \U$20410 ( \20753 , \20752 );
and \U$20411 ( \20754 , \20735 , \20753 );
not \U$20412 ( \20755 , \20722 );
nor \U$20413 ( \20756 , \20755 , \20734 );
nor \U$20414 ( \20757 , \20754 , \20756 );
not \U$20415 ( \20758 , RIbb2e800_31);
not \U$20416 ( \20759 , \14041 );
or \U$20417 ( \20760 , \20758 , \20759 );
nand \U$20418 ( \20761 , \7308 , \9169 );
nand \U$20419 ( \20762 , \20760 , \20761 );
and \U$20420 ( \20763 , \2939 , \20762 );
not \U$20421 ( \20764 , RIbb2e800_31);
not \U$20422 ( \20765 , \6231 );
or \U$20423 ( \20766 , \20764 , \20765 );
nand \U$20424 ( \20767 , \20766 , \19994 );
and \U$20425 ( \20768 , \20767 , \3613 );
nor \U$20426 ( \20769 , \20763 , \20768 );
xor \U$20427 ( \20770 , \20757 , \20769 );
not \U$20428 ( \20771 , RIbb2e8f0_29);
not \U$20429 ( \20772 , \12791 );
not \U$20430 ( \20773 , \20772 );
or \U$20431 ( \20774 , \20771 , \20773 );
nand \U$20432 ( \20775 , \8638 , \2911 );
nand \U$20433 ( \20776 , \20774 , \20775 );
and \U$20434 ( \20777 , \20776 , \2922 );
not \U$20435 ( \20778 , \20008 );
nor \U$20436 ( \20779 , \20778 , \4460 );
nor \U$20437 ( \20780 , \20777 , \20779 );
and \U$20438 ( \20781 , \20770 , \20780 );
and \U$20439 ( \20782 , \20757 , \20769 );
or \U$20440 ( \20783 , \20781 , \20782 );
or \U$20441 ( \20784 , \20711 , \20783 );
nand \U$20442 ( \20785 , \20677 , \20710 );
nand \U$20443 ( \20786 , \20784 , \20785 );
xor \U$20444 ( \20787 , \20377 , \20379 );
xor \U$20445 ( \20788 , \20787 , \20408 );
xor \U$20446 ( \20789 , \20786 , \20788 );
xor \U$20447 ( \20790 , \20039 , \20051 );
xor \U$20448 ( \20791 , \20790 , \20062 );
buf \U$20449 ( \20792 , \6241 );
not \U$20450 ( \20793 , \20792 );
not \U$20451 ( \20794 , \20228 );
or \U$20452 ( \20795 , \20793 , \20794 );
not \U$20453 ( \20796 , RIbb2e530_37);
not \U$20454 ( \20797 , \3001 );
or \U$20455 ( \20798 , \20796 , \20797 );
nand \U$20456 ( \20799 , \3274 , \6246 );
nand \U$20457 ( \20800 , \20798 , \20799 );
nand \U$20458 ( \20801 , \20800 , \6251 );
nand \U$20459 ( \20802 , \20795 , \20801 );
not \U$20460 ( \20803 , \12774 );
xor \U$20461 ( \20804 , RIbb2dea0_51, \1384 );
not \U$20462 ( \20805 , \20804 );
or \U$20463 ( \20806 , \20803 , \20805 );
nand \U$20464 ( \20807 , \20217 , \12692 );
nand \U$20465 ( \20808 , \20806 , \20807 );
xor \U$20466 ( \20809 , \20802 , \20808 );
not \U$20467 ( \20810 , \7104 );
not \U$20468 ( \20811 , \20279 );
or \U$20469 ( \20812 , \20810 , \20811 );
and \U$20470 ( \20813 , RIbb2e440_39, \4015 );
not \U$20471 ( \20814 , RIbb2e440_39);
and \U$20472 ( \20815 , \20814 , \4022 );
or \U$20473 ( \20816 , \20813 , \20815 );
nand \U$20474 ( \20817 , \20816 , \7103 );
nand \U$20475 ( \20818 , \20812 , \20817 );
and \U$20476 ( \20819 , \20809 , \20818 );
and \U$20477 ( \20820 , \20802 , \20808 );
or \U$20478 ( \20821 , \20819 , \20820 );
xor \U$20479 ( \20822 , \20791 , \20821 );
xor \U$20480 ( \20823 , \20382 , \20394 );
xor \U$20481 ( \20824 , \20823 , \20405 );
and \U$20482 ( \20825 , \20822 , \20824 );
and \U$20483 ( \20826 , \20791 , \20821 );
or \U$20484 ( \20827 , \20825 , \20826 );
and \U$20485 ( \20828 , \20789 , \20827 );
and \U$20486 ( \20829 , \20786 , \20788 );
or \U$20487 ( \20830 , \20828 , \20829 );
not \U$20488 ( \20831 , \20830 );
not \U$20489 ( \20832 , \20831 );
or \U$20490 ( \20833 , \20639 , \20832 );
not \U$20491 ( \20834 , \8353 );
not \U$20492 ( \20835 , \20187 );
or \U$20493 ( \20836 , \20834 , \20835 );
not \U$20494 ( \20837 , RIbb2e350_41);
not \U$20495 ( \20838 , \3223 );
not \U$20496 ( \20839 , \20838 );
or \U$20497 ( \20840 , \20837 , \20839 );
nand \U$20498 ( \20841 , \13392 , \3223 );
nand \U$20499 ( \20842 , \20840 , \20841 );
nand \U$20500 ( \20843 , \20842 , \8362 );
nand \U$20501 ( \20844 , \20836 , \20843 );
not \U$20502 ( \20845 , \20844 );
not \U$20503 ( \20846 , \16271 );
xor \U$20504 ( \20847 , RIbb2dae0_59, \1547 );
not \U$20505 ( \20848 , \20847 );
or \U$20506 ( \20849 , \20846 , \20848 );
nand \U$20507 ( \20850 , \20173 , \16257 );
nand \U$20508 ( \20851 , \20849 , \20850 );
not \U$20509 ( \20852 , \20851 );
or \U$20510 ( \20853 , \20845 , \20852 );
not \U$20511 ( \20854 , \20851 );
not \U$20512 ( \20855 , \20854 );
not \U$20513 ( \20856 , \20844 );
not \U$20514 ( \20857 , \20856 );
or \U$20515 ( \20858 , \20855 , \20857 );
not \U$20516 ( \20859 , \13467 );
xor \U$20517 ( \20860 , RIbb2ddb0_53, \1280 );
not \U$20518 ( \20861 , \20860 );
or \U$20519 ( \20862 , \20859 , \20861 );
nand \U$20520 ( \20863 , \20305 , \14929 );
nand \U$20521 ( \20864 , \20862 , \20863 );
nand \U$20522 ( \20865 , \20858 , \20864 );
nand \U$20523 ( \20866 , \20853 , \20865 );
not \U$20524 ( \20867 , \20866 );
xor \U$20525 ( \20868 , \20025 , \19999 );
xnor \U$20526 ( \20869 , \20868 , \20012 );
not \U$20527 ( \20870 , \20869 );
not \U$20528 ( \20871 , \20870 );
or \U$20529 ( \20872 , \20867 , \20871 );
not \U$20530 ( \20873 , \20869 );
not \U$20531 ( \20874 , \20866 );
not \U$20532 ( \20875 , \20874 );
or \U$20533 ( \20876 , \20873 , \20875 );
xor \U$20534 ( \20877 , \20105 , \20111 );
xor \U$20535 ( \20878 , \20877 , \20122 );
nand \U$20536 ( \20879 , \20876 , \20878 );
nand \U$20537 ( \20880 , \20872 , \20879 );
not \U$20538 ( \20881 , \20070 );
not \U$20539 ( \20882 , \20125 );
or \U$20540 ( \20883 , \20881 , \20882 );
or \U$20541 ( \20884 , \20125 , \20070 );
nand \U$20542 ( \20885 , \20883 , \20884 );
xor \U$20543 ( \20886 , \20885 , \20065 );
xor \U$20544 ( \20887 , \20880 , \20886 );
not \U$20545 ( \20888 , \17275 );
not \U$20546 ( \20889 , RIbb2d900_63);
not \U$20547 ( \20890 , \985 );
or \U$20548 ( \20891 , \20889 , \20890 );
nand \U$20549 ( \20892 , \984 , \17262 );
nand \U$20550 ( \20893 , \20891 , \20892 );
not \U$20551 ( \20894 , \20893 );
or \U$20552 ( \20895 , \20888 , \20894 );
nand \U$20553 ( \20896 , \20256 , RIbb2d888_64);
nand \U$20554 ( \20897 , \20895 , \20896 );
not \U$20555 ( \20898 , \17397 );
not \U$20556 ( \20899 , \20319 );
or \U$20557 ( \20900 , \20898 , \20899 );
not \U$20558 ( \20901 , RIbb2dbd0_57);
not \U$20559 ( \20902 , \1686 );
or \U$20560 ( \20903 , \20901 , \20902 );
nand \U$20561 ( \20904 , \3363 , \14602 );
nand \U$20562 ( \20905 , \20903 , \20904 );
nand \U$20563 ( \20906 , \20905 , \16674 );
nand \U$20564 ( \20907 , \20900 , \20906 );
xor \U$20565 ( \20908 , \20897 , \20907 );
not \U$20566 ( \20909 , \11176 );
and \U$20567 ( \20910 , \2115 , RIbb2e080_47);
not \U$20568 ( \20911 , \2115 );
and \U$20569 ( \20912 , \20911 , \16171 );
or \U$20570 ( \20913 , \20910 , \20912 );
not \U$20571 ( \20914 , \20913 );
or \U$20572 ( \20915 , \20909 , \20914 );
nand \U$20573 ( \20916 , \20329 , \11177 );
nand \U$20574 ( \20917 , \20915 , \20916 );
and \U$20575 ( \20918 , \20908 , \20917 );
and \U$20576 ( \20919 , \20897 , \20907 );
or \U$20577 ( \20920 , \20918 , \20919 );
xor \U$20578 ( \20921 , \20082 , \20091 );
xor \U$20579 ( \20922 , \20921 , \20102 );
not \U$20580 ( \20923 , \16541 );
not \U$20581 ( \20924 , RIbb2d9f0_61);
not \U$20582 ( \20925 , \1070 );
or \U$20583 ( \20926 , \20924 , \20925 );
nand \U$20584 ( \20927 , \1886 , \19746 );
nand \U$20585 ( \20928 , \20926 , \20927 );
not \U$20586 ( \20929 , \20928 );
or \U$20587 ( \20930 , \20923 , \20929 );
nand \U$20588 ( \20931 , \20348 , \16533 );
nand \U$20589 ( \20932 , \20930 , \20931 );
xor \U$20590 ( \20933 , \20922 , \20932 );
not \U$20591 ( \20934 , \12167 );
not \U$20592 ( \20935 , RIbb2df90_49);
not \U$20593 ( \20936 , \3494 );
or \U$20594 ( \20937 , \20935 , \20936 );
not \U$20595 ( \20938 , \19733 );
nand \U$20596 ( \20939 , \20938 , \12278 );
nand \U$20597 ( \20940 , \20937 , \20939 );
not \U$20598 ( \20941 , \20940 );
or \U$20599 ( \20942 , \20934 , \20941 );
nand \U$20600 ( \20943 , \20401 , \12285 );
nand \U$20601 ( \20944 , \20942 , \20943 );
and \U$20602 ( \20945 , \20933 , \20944 );
and \U$20603 ( \20946 , \20922 , \20932 );
or \U$20604 ( \20947 , \20945 , \20946 );
xor \U$20605 ( \20948 , \20920 , \20947 );
not \U$20606 ( \20949 , \10117 );
not \U$20607 ( \20950 , RIbb2e170_45);
not \U$20608 ( \20951 , \3341 );
not \U$20609 ( \20952 , \20951 );
or \U$20610 ( \20953 , \20950 , \20952 );
nand \U$20611 ( \20954 , \3341 , \12003 );
nand \U$20612 ( \20955 , \20953 , \20954 );
not \U$20613 ( \20956 , \20955 );
or \U$20614 ( \20957 , \20949 , \20956 );
nand \U$20615 ( \20958 , \20243 , \10119 );
nand \U$20616 ( \20959 , \20957 , \20958 );
not \U$20617 ( \20960 , \10449 );
not \U$20618 ( \20961 , RIbb2e260_43);
not \U$20619 ( \20962 , \17568 );
or \U$20620 ( \20963 , \20961 , \20962 );
nand \U$20621 ( \20964 , \3146 , \10444 );
nand \U$20622 ( \20965 , \20963 , \20964 );
not \U$20623 ( \20966 , \20965 );
or \U$20624 ( \20967 , \20960 , \20966 );
nand \U$20625 ( \20968 , \20196 , \9099 );
nand \U$20626 ( \20969 , \20967 , \20968 );
nor \U$20627 ( \20970 , \20959 , \20969 );
not \U$20628 ( \20971 , \15181 );
not \U$20629 ( \20972 , \20264 );
or \U$20630 ( \20973 , \20971 , \20972 );
and \U$20631 ( \20974 , RIbb2dcc0_55, \7423 );
not \U$20632 ( \20975 , RIbb2dcc0_55);
and \U$20633 ( \20976 , \20975 , \1136 );
or \U$20634 ( \20977 , \20974 , \20976 );
nand \U$20635 ( \20978 , \20977 , \14613 );
nand \U$20636 ( \20979 , \20973 , \20978 );
not \U$20637 ( \20980 , \20979 );
or \U$20638 ( \20981 , \20970 , \20980 );
nand \U$20639 ( \20982 , \20959 , \20969 );
nand \U$20640 ( \20983 , \20981 , \20982 );
and \U$20641 ( \20984 , \20948 , \20983 );
and \U$20642 ( \20985 , \20920 , \20947 );
or \U$20643 ( \20986 , \20984 , \20985 );
and \U$20644 ( \20987 , \20887 , \20986 );
and \U$20645 ( \20988 , \20880 , \20886 );
or \U$20646 ( \20989 , \20987 , \20988 );
nand \U$20647 ( \20990 , \20833 , \20989 );
or \U$20648 ( \20991 , \20831 , \20638 );
nand \U$20649 ( \20992 , \20990 , \20991 );
xor \U$20650 ( \20993 , \20235 , \20237 );
xor \U$20651 ( \20994 , \20993 , \20354 );
not \U$20652 ( \20995 , \20994 );
xor \U$20653 ( \20996 , \20350 , \20336 );
xnor \U$20654 ( \20997 , \20996 , \20338 );
not \U$20655 ( \20998 , \20997 );
not \U$20656 ( \20999 , \20998 );
not \U$20657 ( \21000 , \20247 );
not \U$20658 ( \21001 , \20269 );
or \U$20659 ( \21002 , \21000 , \21001 );
or \U$20660 ( \21003 , \20247 , \20269 );
nand \U$20661 ( \21004 , \21002 , \21003 );
not \U$20662 ( \21005 , \20258 );
and \U$20663 ( \21006 , \21004 , \21005 );
not \U$20664 ( \21007 , \21004 );
and \U$20665 ( \21008 , \21007 , \20258 );
nor \U$20666 ( \21009 , \21006 , \21008 );
not \U$20667 ( \21010 , \21009 );
not \U$20668 ( \21011 , \21010 );
or \U$20669 ( \21012 , \20999 , \21011 );
not \U$20670 ( \21013 , \20997 );
not \U$20671 ( \21014 , \21009 );
or \U$20672 ( \21015 , \21013 , \21014 );
xor \U$20673 ( \21016 , \20177 , \20200 );
xor \U$20674 ( \21017 , \21016 , \20202 );
nand \U$20675 ( \21018 , \21015 , \21017 );
nand \U$20676 ( \21019 , \21012 , \21018 );
not \U$20677 ( \21020 , \21019 );
not \U$20678 ( \21021 , \20204 );
not \U$20679 ( \21022 , \21021 );
not \U$20680 ( \21023 , \20167 );
or \U$20681 ( \21024 , \21022 , \21023 );
nand \U$20682 ( \21025 , \20204 , \20166 );
nand \U$20683 ( \21026 , \21024 , \21025 );
not \U$20684 ( \21027 , \20233 );
and \U$20685 ( \21028 , \21026 , \21027 );
not \U$20686 ( \21029 , \21026 );
and \U$20687 ( \21030 , \21029 , \20233 );
nor \U$20688 ( \21031 , \21028 , \21030 );
not \U$20689 ( \21032 , \21031 );
not \U$20690 ( \21033 , \21032 );
or \U$20691 ( \21034 , \21020 , \21033 );
not \U$20692 ( \21035 , \21019 );
nand \U$20693 ( \21036 , \21035 , \21031 );
xor \U$20694 ( \21037 , \20592 , \20594 );
xor \U$20695 ( \21038 , \21037 , \20597 );
nand \U$20696 ( \21039 , \21036 , \21038 );
nand \U$20697 ( \21040 , \21034 , \21039 );
not \U$20698 ( \21041 , \21040 );
or \U$20699 ( \21042 , \20995 , \21041 );
or \U$20700 ( \21043 , \21040 , \20994 );
not \U$20701 ( \21044 , \20476 );
not \U$20702 ( \21045 , \20464 );
or \U$20703 ( \21046 , \21044 , \21045 );
or \U$20704 ( \21047 , \20464 , \20476 );
nand \U$20705 ( \21048 , \21046 , \21047 );
buf \U$20706 ( \21049 , \20468 );
and \U$20707 ( \21050 , \21048 , \21049 );
not \U$20708 ( \21051 , \21048 );
and \U$20709 ( \21052 , \21051 , \20469 );
nor \U$20710 ( \21053 , \21050 , \21052 );
not \U$20711 ( \21054 , \21053 );
not \U$20712 ( \21055 , \21054 );
xor \U$20713 ( \21056 , \20272 , \20352 );
xnor \U$20714 ( \21057 , \21056 , \20309 );
not \U$20715 ( \21058 , \21057 );
not \U$20716 ( \21059 , \21058 );
or \U$20717 ( \21060 , \21055 , \21059 );
not \U$20718 ( \21061 , \21053 );
not \U$20719 ( \21062 , \21057 );
or \U$20720 ( \21063 , \21061 , \21062 );
xor \U$20721 ( \21064 , \20209 , \20219 );
xor \U$20722 ( \21065 , \21064 , \20230 );
xor \U$20723 ( \21066 , \20572 , \20573 );
xor \U$20724 ( \21067 , \21066 , \20586 );
xor \U$20725 ( \21068 , \20547 , \20558 );
xor \U$20726 ( \21069 , \21068 , \20569 );
not \U$20727 ( \21070 , \1444 );
and \U$20728 ( \21071 , RIbb2ef80_15, \18829 );
not \U$20729 ( \21072 , RIbb2ef80_15);
and \U$20730 ( \21073 , \21072 , \13977 );
or \U$20731 ( \21074 , \21071 , \21073 );
not \U$20732 ( \21075 , \21074 );
or \U$20733 ( \21076 , \21070 , \21075 );
nand \U$20734 ( \21077 , \20529 , \1517 );
nand \U$20735 ( \21078 , \21076 , \21077 );
xor \U$20736 ( \21079 , \21069 , \21078 );
not \U$20737 ( \21080 , \836 );
not \U$20738 ( \21081 , \20538 );
or \U$20739 ( \21082 , \21080 , \21081 );
and \U$20740 ( \21083 , \13210 , \3057 );
not \U$20741 ( \21084 , \13210 );
and \U$20742 ( \21085 , \21084 , RIbb2ee90_17);
or \U$20743 ( \21086 , \21083 , \21085 );
nand \U$20744 ( \21087 , \832 , \21086 );
nand \U$20745 ( \21088 , \21082 , \21087 );
and \U$20746 ( \21089 , \21079 , \21088 );
and \U$20747 ( \21090 , \21069 , \21078 );
or \U$20748 ( \21091 , \21089 , \21090 );
xor \U$20749 ( \21092 , \21067 , \21091 );
not \U$20750 ( \21093 , \20292 );
not \U$20751 ( \21094 , \5845 );
or \U$20752 ( \21095 , \21093 , \21094 );
not \U$20753 ( \21096 , RIbb2e620_35);
not \U$20754 ( \21097 , \13756 );
or \U$20755 ( \21098 , \21096 , \21097 );
nand \U$20756 ( \21099 , \4324 , \6688 );
nand \U$20757 ( \21100 , \21098 , \21099 );
nand \U$20758 ( \21101 , \21100 , \4712 );
nand \U$20759 ( \21102 , \21095 , \21101 );
and \U$20760 ( \21103 , \21092 , \21102 );
and \U$20761 ( \21104 , \21067 , \21091 );
or \U$20762 ( \21105 , \21103 , \21104 );
xor \U$20763 ( \21106 , \21065 , \21105 );
not \U$20764 ( \21107 , \20294 );
not \U$20765 ( \21108 , \21107 );
not \U$20766 ( \21109 , \8450 );
not \U$20767 ( \21110 , \19664 );
or \U$20768 ( \21111 , \21109 , \21110 );
not \U$20769 ( \21112 , \8444 );
nand \U$20770 ( \21113 , \21112 , \20279 );
nand \U$20771 ( \21114 , \21111 , \21113 );
not \U$20772 ( \21115 , \21114 );
not \U$20773 ( \21116 , \20307 );
not \U$20774 ( \21117 , \21116 );
or \U$20775 ( \21118 , \21115 , \21117 );
or \U$20776 ( \21119 , \21116 , \20283 );
nand \U$20777 ( \21120 , \21118 , \21119 );
not \U$20778 ( \21121 , \21120 );
or \U$20779 ( \21122 , \21108 , \21121 );
or \U$20780 ( \21123 , \21120 , \21107 );
nand \U$20781 ( \21124 , \21122 , \21123 );
and \U$20782 ( \21125 , \21106 , \21124 );
and \U$20783 ( \21126 , \21065 , \21105 );
or \U$20784 ( \21127 , \21125 , \21126 );
nand \U$20785 ( \21128 , \21063 , \21127 );
nand \U$20786 ( \21129 , \21060 , \21128 );
nand \U$20787 ( \21130 , \21043 , \21129 );
nand \U$20788 ( \21131 , \21042 , \21130 );
xor \U$20789 ( \21132 , \20992 , \21131 );
xor \U$20790 ( \21133 , \20164 , \20357 );
xor \U$20791 ( \21134 , \21133 , \20360 );
and \U$20792 ( \21135 , \21132 , \21134 );
and \U$20793 ( \21136 , \20992 , \21131 );
or \U$20794 ( \21137 , \21135 , \21136 );
not \U$20795 ( \21138 , \20368 );
not \U$20796 ( \21139 , \21138 );
not \U$20797 ( \21140 , \20363 );
not \U$20798 ( \21141 , \20162 );
or \U$20799 ( \21142 , \21140 , \21141 );
or \U$20800 ( \21143 , \20162 , \20363 );
nand \U$20801 ( \21144 , \21142 , \21143 );
not \U$20802 ( \21145 , \21144 );
or \U$20803 ( \21146 , \21139 , \21145 );
or \U$20804 ( \21147 , \21144 , \21138 );
nand \U$20805 ( \21148 , \21146 , \21147 );
xor \U$20806 ( \21149 , \21137 , \21148 );
xor \U$20807 ( \21150 , \20478 , \20452 );
xor \U$20808 ( \21151 , \21150 , \20455 );
not \U$20809 ( \21152 , \21151 );
not \U$20810 ( \21153 , \21152 );
xor \U$20811 ( \21154 , \20411 , \20413 );
xor \U$20812 ( \21155 , \21154 , \20439 );
not \U$20813 ( \21156 , \21155 );
not \U$20814 ( \21157 , \21156 );
not \U$20815 ( \21158 , \21157 );
or \U$20816 ( \21159 , \21153 , \21158 );
not \U$20817 ( \21160 , \21156 );
not \U$20818 ( \21161 , \21151 );
or \U$20819 ( \21162 , \21160 , \21161 );
not \U$20820 ( \21163 , \20434 );
not \U$20821 ( \21164 , \20421 );
not \U$20822 ( \21165 , \21164 );
or \U$20823 ( \21166 , \21163 , \21165 );
nand \U$20824 ( \21167 , \20433 , \20421 );
nand \U$20825 ( \21168 , \21166 , \21167 );
and \U$20826 ( \21169 , \21168 , \20437 );
not \U$20827 ( \21170 , \21168 );
and \U$20828 ( \21171 , \21170 , \20425 );
nor \U$20829 ( \21172 , \21169 , \21171 );
not \U$20830 ( \21173 , \20545 );
not \U$20831 ( \21174 , \20589 );
not \U$20832 ( \21175 , \21174 );
or \U$20833 ( \21176 , \21173 , \21175 );
or \U$20834 ( \21177 , \20545 , \21174 );
nand \U$20835 ( \21178 , \21176 , \21177 );
xor \U$20836 ( \21179 , \20512 , \21178 );
not \U$20837 ( \21180 , \3886 );
not \U$20838 ( \21181 , RIbb2e710_33);
not \U$20839 ( \21182 , \6230 );
or \U$20840 ( \21183 , \21181 , \21182 );
nand \U$20841 ( \21184 , \6229 , \3882 );
nand \U$20842 ( \21185 , \21183 , \21184 );
not \U$20843 ( \21186 , \21185 );
or \U$20844 ( \21187 , \21180 , \21186 );
nand \U$20845 ( \21188 , \20657 , \4075 );
nand \U$20846 ( \21189 , \21187 , \21188 );
not \U$20847 ( \21190 , \3406 );
not \U$20848 ( \21191 , RIbb2ebc0_23);
not \U$20849 ( \21192 , \18802 );
or \U$20850 ( \21193 , \21191 , \21192 );
nand \U$20851 ( \21194 , \10764 , \3388 );
nand \U$20852 ( \21195 , \21193 , \21194 );
not \U$20853 ( \21196 , \21195 );
or \U$20854 ( \21197 , \21190 , \21196 );
nand \U$20855 ( \21198 , \20705 , \3382 );
nand \U$20856 ( \21199 , \21197 , \21198 );
xor \U$20857 ( \21200 , \21189 , \21199 );
not \U$20858 ( \21201 , \3445 );
and \U$20859 ( \21202 , \15786 , RIbb2e9e0_27);
not \U$20860 ( \21203 , \15786 );
and \U$20861 ( \21204 , \21203 , \3454 );
or \U$20862 ( \21205 , \21202 , \21204 );
not \U$20863 ( \21206 , \21205 );
or \U$20864 ( \21207 , \21201 , \21206 );
nand \U$20865 ( \21208 , \20694 , \3465 );
nand \U$20866 ( \21209 , \21207 , \21208 );
and \U$20867 ( \21210 , \21200 , \21209 );
and \U$20868 ( \21211 , \21189 , \21199 );
or \U$20869 ( \21212 , \21210 , \21211 );
not \U$20870 ( \21213 , \21212 );
not \U$20871 ( \21214 , \998 );
not \U$20872 ( \21215 , \20582 );
or \U$20873 ( \21216 , \21214 , \21215 );
not \U$20874 ( \21217 , RIbb2f070_13);
not \U$20875 ( \21218 , \15469 );
or \U$20876 ( \21219 , \21217 , \21218 );
nand \U$20877 ( \21220 , \15030 , \1656 );
nand \U$20878 ( \21221 , \21219 , \21220 );
nand \U$20879 ( \21222 , \21221 , \916 );
nand \U$20880 ( \21223 , \21216 , \21222 );
not \U$20881 ( \21224 , \854 );
not \U$20882 ( \21225 , \20646 );
or \U$20883 ( \21226 , \21224 , \21225 );
not \U$20884 ( \21227 , RIbb2eda0_19);
not \U$20885 ( \21228 , \17663 );
or \U$20886 ( \21229 , \21227 , \21228 );
nand \U$20887 ( \21230 , \12932 , \843 );
nand \U$20888 ( \21231 , \21229 , \21230 );
nand \U$20889 ( \21232 , \21231 , \853 );
nand \U$20890 ( \21233 , \21226 , \21232 );
xor \U$20891 ( \21234 , \21223 , \21233 );
not \U$20892 ( \21235 , \4714 );
not \U$20893 ( \21236 , \21100 );
or \U$20894 ( \21237 , \21235 , \21236 );
not \U$20895 ( \21238 , RIbb2e620_35);
not \U$20896 ( \21239 , \14536 );
or \U$20897 ( \21240 , \21238 , \21239 );
nand \U$20898 ( \21241 , \4390 , \3866 );
nand \U$20899 ( \21242 , \21240 , \21241 );
nand \U$20900 ( \21243 , \21242 , \4712 );
nand \U$20901 ( \21244 , \21237 , \21243 );
and \U$20902 ( \21245 , \21234 , \21244 );
and \U$20903 ( \21246 , \21223 , \21233 );
or \U$20904 ( \21247 , \21245 , \21246 );
not \U$20905 ( \21248 , \21247 );
nand \U$20906 ( \21249 , \21213 , \21248 );
not \U$20907 ( \21250 , \21249 );
not \U$20908 ( \21251 , \20740 );
not \U$20909 ( \21252 , \20751 );
or \U$20910 ( \21253 , \21251 , \21252 );
or \U$20911 ( \21254 , \20751 , \20740 );
nand \U$20912 ( \21255 , \21253 , \21254 );
not \U$20913 ( \21256 , \1737 );
not \U$20914 ( \21257 , \20565 );
or \U$20915 ( \21258 , \21256 , \21257 );
not \U$20916 ( \21259 , RIbb2f340_7);
not \U$20917 ( \21260 , \16819 );
or \U$20918 ( \21261 , \21259 , \21260 );
nand \U$20919 ( \21262 , \17529 , \1734 );
nand \U$20920 ( \21263 , \21261 , \21262 );
nand \U$20921 ( \21264 , \21263 , \1701 );
nand \U$20922 ( \21265 , \21258 , \21264 );
xor \U$20923 ( \21266 , \21255 , \21265 );
not \U$20924 ( \21267 , \1011 );
not \U$20925 ( \21268 , RIbb2f160_11);
not \U$20926 ( \21269 , \16747 );
or \U$20927 ( \21270 , \21268 , \21269 );
nand \U$20928 ( \21271 , \19077 , \1043 );
nand \U$20929 ( \21272 , \21270 , \21271 );
not \U$20930 ( \21273 , \21272 );
or \U$20931 ( \21274 , \21267 , \21273 );
nand \U$20932 ( \21275 , \20720 , \1077 );
nand \U$20933 ( \21276 , \21274 , \21275 );
and \U$20934 ( \21277 , \21266 , \21276 );
and \U$20935 ( \21278 , \21255 , \21265 );
or \U$20936 ( \21279 , \21277 , \21278 );
not \U$20937 ( \21280 , \2939 );
not \U$20938 ( \21281 , RIbb2e800_31);
not \U$20939 ( \21282 , \13875 );
or \U$20940 ( \21283 , \21281 , \21282 );
nand \U$20941 ( \21284 , \6604 , \3608 );
nand \U$20942 ( \21285 , \21283 , \21284 );
not \U$20943 ( \21286 , \21285 );
or \U$20944 ( \21287 , \21280 , \21286 );
nand \U$20945 ( \21288 , \20762 , \3613 );
nand \U$20946 ( \21289 , \21287 , \21288 );
xor \U$20947 ( \21290 , \21279 , \21289 );
not \U$20948 ( \21291 , \2922 );
not \U$20949 ( \21292 , RIbb2e8f0_29);
not \U$20950 ( \21293 , \13853 );
or \U$20951 ( \21294 , \21292 , \21293 );
not \U$20952 ( \21295 , \9070 );
nand \U$20953 ( \21296 , \21295 , \3265 );
nand \U$20954 ( \21297 , \21294 , \21296 );
not \U$20955 ( \21298 , \21297 );
or \U$20956 ( \21299 , \21291 , \21298 );
nand \U$20957 ( \21300 , \20776 , \2925 );
nand \U$20958 ( \21301 , \21299 , \21300 );
and \U$20959 ( \21302 , \21290 , \21301 );
and \U$20960 ( \21303 , \21279 , \21289 );
or \U$20961 ( \21304 , \21302 , \21303 );
not \U$20962 ( \21305 , \21304 );
or \U$20963 ( \21306 , \21250 , \21305 );
nand \U$20964 ( \21307 , \21212 , \21247 );
nand \U$20965 ( \21308 , \21306 , \21307 );
xor \U$20966 ( \21309 , \21179 , \21308 );
xor \U$20967 ( \21310 , \20522 , \20531 );
xor \U$20968 ( \21311 , \21310 , \20542 );
xor \U$20969 ( \21312 , \20688 , \20696 );
xor \U$20970 ( \21313 , \21312 , \20707 );
xor \U$20971 ( \21314 , \21311 , \21313 );
xor \U$20972 ( \21315 , \20752 , \20733 );
xnor \U$20973 ( \21316 , \21315 , \20722 );
not \U$20974 ( \21317 , \6251 );
not \U$20975 ( \21318 , RIbb2e530_37);
not \U$20976 ( \21319 , \3090 );
or \U$20977 ( \21320 , \21318 , \21319 );
nand \U$20978 ( \21321 , \3089 , \4708 );
nand \U$20979 ( \21322 , \21320 , \21321 );
not \U$20980 ( \21323 , \21322 );
or \U$20981 ( \21324 , \21317 , \21323 );
nand \U$20982 ( \21325 , \20800 , \6242 );
nand \U$20983 ( \21326 , \21324 , \21325 );
xor \U$20984 ( \21327 , \21316 , \21326 );
not \U$20985 ( \21328 , \7103 );
and \U$20986 ( \21329 , RIbb2e440_39, \3045 );
not \U$20987 ( \21330 , RIbb2e440_39);
and \U$20988 ( \21331 , \21330 , \3046 );
or \U$20989 ( \21332 , \21329 , \21331 );
not \U$20990 ( \21333 , \21332 );
or \U$20991 ( \21334 , \21328 , \21333 );
nand \U$20992 ( \21335 , \20816 , \8450 );
nand \U$20993 ( \21336 , \21334 , \21335 );
and \U$20994 ( \21337 , \21327 , \21336 );
and \U$20995 ( \21338 , \21316 , \21326 );
or \U$20996 ( \21339 , \21337 , \21338 );
and \U$20997 ( \21340 , \21314 , \21339 );
and \U$20998 ( \21341 , \21311 , \21313 );
or \U$20999 ( \21342 , \21340 , \21341 );
and \U$21000 ( \21343 , \21309 , \21342 );
and \U$21001 ( \21344 , \21179 , \21308 );
or \U$21002 ( \21345 , \21343 , \21344 );
xor \U$21003 ( \21346 , \21172 , \21345 );
xor \U$21004 ( \21347 , \20648 , \20674 );
xor \U$21005 ( \21348 , \21347 , \20662 );
not \U$21006 ( \21349 , \21348 );
not \U$21007 ( \21350 , \2077 );
and \U$21008 ( \21351 , \11578 , \2254 );
not \U$21009 ( \21352 , \11578 );
and \U$21010 ( \21353 , \21352 , RIbb2ecb0_21);
or \U$21011 ( \21354 , \21351 , \21353 );
not \U$21012 ( \21355 , \21354 );
or \U$21013 ( \21356 , \21350 , \21355 );
nand \U$21014 ( \21357 , \20672 , \2078 );
nand \U$21015 ( \21358 , \21356 , \21357 );
not \U$21016 ( \21359 , \21358 );
not \U$21017 ( \21360 , \21359 );
not \U$21018 ( \21361 , \2980 );
and \U$21019 ( \21362 , RIbb2ead0_25, \13498 );
not \U$21020 ( \21363 , RIbb2ead0_25);
and \U$21021 ( \21364 , \21363 , \9840 );
or \U$21022 ( \21365 , \21362 , \21364 );
not \U$21023 ( \21366 , \21365 );
or \U$21024 ( \21367 , \21361 , \21366 );
nand \U$21025 ( \21368 , \20684 , \2963 );
nand \U$21026 ( \21369 , \21367 , \21368 );
not \U$21027 ( \21370 , \21369 );
not \U$21028 ( \21371 , \21370 );
or \U$21029 ( \21372 , \21360 , \21371 );
not \U$21030 ( \21373 , \12167 );
not \U$21031 ( \21374 , RIbb2df90_49);
not \U$21032 ( \21375 , \14725 );
or \U$21033 ( \21376 , \21374 , \21375 );
nand \U$21034 ( \21377 , \1852 , \12278 );
nand \U$21035 ( \21378 , \21376 , \21377 );
not \U$21036 ( \21379 , \21378 );
or \U$21037 ( \21380 , \21373 , \21379 );
nand \U$21038 ( \21381 , \20940 , \14752 );
nand \U$21039 ( \21382 , \21380 , \21381 );
nand \U$21040 ( \21383 , \21372 , \21382 );
not \U$21041 ( \21384 , \21359 );
nand \U$21042 ( \21385 , \21384 , \21369 );
nand \U$21043 ( \21386 , \21383 , \21385 );
not \U$21044 ( \21387 , \21386 );
not \U$21045 ( \21388 , \21387 );
or \U$21046 ( \21389 , \21349 , \21388 );
xor \U$21047 ( \21390 , \20757 , \20769 );
xor \U$21048 ( \21391 , \21390 , \20780 );
not \U$21049 ( \21392 , \21391 );
nand \U$21050 ( \21393 , \21389 , \21392 );
not \U$21051 ( \21394 , \21348 );
nand \U$21052 ( \21395 , \21394 , \21386 );
nand \U$21053 ( \21396 , \21393 , \21395 );
xor \U$21054 ( \21397 , \20710 , \20677 );
not \U$21055 ( \21398 , \20783 );
xor \U$21056 ( \21399 , \21397 , \21398 );
xor \U$21057 ( \21400 , \21396 , \21399 );
not \U$21058 ( \21401 , \9098 );
not \U$21059 ( \21402 , RIbb2e260_43);
not \U$21060 ( \21403 , \16399 );
or \U$21061 ( \21404 , \21402 , \21403 );
nand \U$21062 ( \21405 , \3201 , \8347 );
nand \U$21063 ( \21406 , \21404 , \21405 );
not \U$21064 ( \21407 , \21406 );
or \U$21065 ( \21408 , \21401 , \21407 );
nand \U$21066 ( \21409 , \20965 , \9099 );
nand \U$21067 ( \21410 , \21408 , \21409 );
not \U$21068 ( \21411 , \10119 );
not \U$21069 ( \21412 , \20955 );
or \U$21070 ( \21413 , \21411 , \21412 );
and \U$21071 ( \21414 , RIbb2e170_45, \13414 );
not \U$21072 ( \21415 , RIbb2e170_45);
and \U$21073 ( \21416 , \21415 , \3166 );
or \U$21074 ( \21417 , \21414 , \21416 );
nand \U$21075 ( \21418 , \21417 , \10599 );
nand \U$21076 ( \21419 , \21413 , \21418 );
or \U$21077 ( \21420 , \21410 , \21419 );
not \U$21078 ( \21421 , \14613 );
and \U$21079 ( \21422 , RIbb2dcc0_55, \4766 );
not \U$21080 ( \21423 , RIbb2dcc0_55);
and \U$21081 ( \21424 , \21423 , \1111 );
or \U$21082 ( \21425 , \21422 , \21424 );
not \U$21083 ( \21426 , \21425 );
or \U$21084 ( \21427 , \21421 , \21426 );
nand \U$21085 ( \21428 , \20977 , \15181 );
nand \U$21086 ( \21429 , \21427 , \21428 );
nand \U$21087 ( \21430 , \21420 , \21429 );
nand \U$21088 ( \21431 , \21419 , \21410 );
nand \U$21089 ( \21432 , \21430 , \21431 );
not \U$21090 ( \21433 , \16674 );
not \U$21091 ( \21434 , RIbb2dbd0_57);
not \U$21092 ( \21435 , \3238 );
or \U$21093 ( \21436 , \21434 , \21435 );
nand \U$21094 ( \21437 , \1642 , \17097 );
nand \U$21095 ( \21438 , \21436 , \21437 );
not \U$21096 ( \21439 , \21438 );
or \U$21097 ( \21440 , \21433 , \21439 );
nand \U$21098 ( \21441 , \20905 , \15738 );
nand \U$21099 ( \21442 , \21440 , \21441 );
not \U$21100 ( \21443 , \16533 );
not \U$21101 ( \21444 , \20928 );
or \U$21102 ( \21445 , \21443 , \21444 );
not \U$21103 ( \21446 , RIbb2d9f0_61);
not \U$21104 ( \21447 , \18204 );
or \U$21105 ( \21448 , \21446 , \21447 );
not \U$21106 ( \21449 , RIbb2d9f0_61);
nand \U$21107 ( \21450 , \17410 , \21449 );
nand \U$21108 ( \21451 , \21448 , \21450 );
nand \U$21109 ( \21452 , \21451 , \18717 );
nand \U$21110 ( \21453 , \21445 , \21452 );
xor \U$21111 ( \21454 , \21442 , \21453 );
not \U$21112 ( \21455 , \11176 );
not \U$21113 ( \21456 , RIbb2e080_47);
not \U$21114 ( \21457 , \13289 );
or \U$21115 ( \21458 , \21456 , \21457 );
nand \U$21116 ( \21459 , \13290 , \10113 );
nand \U$21117 ( \21460 , \21458 , \21459 );
not \U$21118 ( \21461 , \21460 );
or \U$21119 ( \21462 , \21455 , \21461 );
nand \U$21120 ( \21463 , \20913 , \11177 );
nand \U$21121 ( \21464 , \21462 , \21463 );
and \U$21122 ( \21465 , \21454 , \21464 );
and \U$21123 ( \21466 , \21442 , \21453 );
or \U$21124 ( \21467 , \21465 , \21466 );
xor \U$21125 ( \21468 , \21432 , \21467 );
not \U$21126 ( \21469 , \17275 );
and \U$21127 ( \21470 , \950 , \19721 );
not \U$21128 ( \21471 , \950 );
and \U$21129 ( \21472 , \21471 , RIbb2d900_63);
or \U$21130 ( \21473 , \21470 , \21472 );
not \U$21131 ( \21474 , \21473 );
or \U$21132 ( \21475 , \21469 , \21474 );
nand \U$21133 ( \21476 , \20893 , RIbb2d888_64);
nand \U$21134 ( \21477 , \21475 , \21476 );
not \U$21135 ( \21478 , \13467 );
and \U$21136 ( \21479 , \1169 , \13463 );
not \U$21137 ( \21480 , \1169 );
and \U$21138 ( \21481 , \21480 , RIbb2ddb0_53);
or \U$21139 ( \21482 , \21479 , \21481 );
not \U$21140 ( \21483 , \21482 );
or \U$21141 ( \21484 , \21478 , \21483 );
nand \U$21142 ( \21485 , \20860 , \14930 );
nand \U$21143 ( \21486 , \21484 , \21485 );
xor \U$21144 ( \21487 , \21477 , \21486 );
not \U$21145 ( \21488 , \8362 );
not \U$21146 ( \21489 , RIbb2e350_41);
not \U$21147 ( \21490 , \3653 );
not \U$21148 ( \21491 , \21490 );
or \U$21149 ( \21492 , \21489 , \21491 );
nand \U$21150 ( \21493 , \3653 , \13400 );
nand \U$21151 ( \21494 , \21492 , \21493 );
not \U$21152 ( \21495 , \21494 );
or \U$21153 ( \21496 , \21488 , \21495 );
nand \U$21154 ( \21497 , \20842 , \8354 );
nand \U$21155 ( \21498 , \21496 , \21497 );
and \U$21156 ( \21499 , \21487 , \21498 );
and \U$21157 ( \21500 , \21477 , \21486 );
or \U$21158 ( \21501 , \21499 , \21500 );
and \U$21159 ( \21502 , \21468 , \21501 );
and \U$21160 ( \21503 , \21432 , \21467 );
or \U$21161 ( \21504 , \21502 , \21503 );
and \U$21162 ( \21505 , \21400 , \21504 );
and \U$21163 ( \21506 , \21396 , \21399 );
or \U$21164 ( \21507 , \21505 , \21506 );
and \U$21165 ( \21508 , \21346 , \21507 );
and \U$21166 ( \21509 , \21172 , \21345 );
or \U$21167 ( \21510 , \21508 , \21509 );
nand \U$21168 ( \21511 , \21162 , \21510 );
nand \U$21169 ( \21512 , \21159 , \21511 );
not \U$21170 ( \21513 , \20442 );
not \U$21171 ( \21514 , \20480 );
not \U$21172 ( \21515 , \21514 );
or \U$21173 ( \21516 , \21513 , \21515 );
nand \U$21174 ( \21517 , \20443 , \20480 );
nand \U$21175 ( \21518 , \21516 , \21517 );
not \U$21176 ( \21519 , \20375 );
xor \U$21177 ( \21520 , \21518 , \21519 );
xor \U$21178 ( \21521 , \21512 , \21520 );
not \U$21179 ( \21522 , \20488 );
not \U$21180 ( \21523 , \20606 );
or \U$21181 ( \21524 , \21522 , \21523 );
nand \U$21182 ( \21525 , \20487 , \20602 );
nand \U$21183 ( \21526 , \21524 , \21525 );
and \U$21184 ( \21527 , \21526 , \20610 );
not \U$21185 ( \21528 , \21526 );
not \U$21186 ( \21529 , \20610 );
and \U$21187 ( \21530 , \21528 , \21529 );
nor \U$21188 ( \21531 , \21527 , \21530 );
and \U$21189 ( \21532 , \21521 , \21531 );
and \U$21190 ( \21533 , \21512 , \21520 );
or \U$21191 ( \21534 , \21532 , \21533 );
and \U$21192 ( \21535 , \21149 , \21534 );
and \U$21193 ( \21536 , \21137 , \21148 );
or \U$21194 ( \21537 , \21535 , \21536 );
not \U$21195 ( \21538 , \21537 );
xor \U$21196 ( \21539 , \20135 , \20153 );
xor \U$21197 ( \21540 , \21539 , \20156 );
not \U$21198 ( \21541 , \21540 );
nand \U$21199 ( \21542 , \21538 , \21541 );
not \U$21200 ( \21543 , \21542 );
or \U$21201 ( \21544 , \20636 , \21543 );
nand \U$21202 ( \21545 , \21537 , \21540 );
nand \U$21203 ( \21546 , \21544 , \21545 );
not \U$21204 ( \21547 , \21546 );
nand \U$21205 ( \21548 , \20633 , \21547 );
not \U$21206 ( \21549 , \21548 );
not \U$21207 ( \21550 , \18481 );
not \U$21208 ( \21551 , \19483 );
not \U$21209 ( \21552 , \21551 );
not \U$21210 ( \21553 , \21552 );
or \U$21211 ( \21554 , \21550 , \21553 );
not \U$21212 ( \21555 , \18481 );
nand \U$21213 ( \21556 , \21555 , \21551 );
nand \U$21214 ( \21557 , \21556 , \19949 );
nand \U$21215 ( \21558 , \21554 , \21557 );
or \U$21216 ( \21559 , \18133 , \18079 );
nand \U$21217 ( \21560 , \21559 , \18085 );
nand \U$21218 ( \21561 , \18133 , \18079 );
nand \U$21219 ( \21562 , \21560 , \21561 );
xor \U$21220 ( \21563 , \18269 , \18303 );
and \U$21221 ( \21564 , \21563 , \18344 );
and \U$21222 ( \21565 , \18269 , \18303 );
or \U$21223 ( \21566 , \21564 , \21565 );
xor \U$21224 ( \21567 , \21562 , \21566 );
not \U$21225 ( \21568 , \2078 );
not \U$21226 ( \21569 , RIbb2ecb0_21);
not \U$21227 ( \21570 , \5955 );
not \U$21228 ( \21571 , \21570 );
or \U$21229 ( \21572 , \21569 , \21571 );
nand \U$21230 ( \21573 , \5955 , \2254 );
nand \U$21231 ( \21574 , \21572 , \21573 );
not \U$21232 ( \21575 , \21574 );
or \U$21233 ( \21576 , \21568 , \21575 );
nand \U$21234 ( \21577 , \17064 , \2077 );
nand \U$21235 ( \21578 , \21576 , \21577 );
not \U$21236 ( \21579 , \855 );
not \U$21237 ( \21580 , RIbb2eda0_19);
not \U$21238 ( \21581 , \9791 );
or \U$21239 ( \21582 , \21580 , \21581 );
nand \U$21240 ( \21583 , \19870 , \843 );
nand \U$21241 ( \21584 , \21582 , \21583 );
not \U$21242 ( \21585 , \21584 );
or \U$21243 ( \21586 , \21579 , \21585 );
nand \U$21244 ( \21587 , \17072 , \853 );
nand \U$21245 ( \21588 , \21586 , \21587 );
and \U$21246 ( \21589 , \21578 , \21588 );
not \U$21247 ( \21590 , \21578 );
not \U$21248 ( \21591 , \21588 );
and \U$21249 ( \21592 , \21590 , \21591 );
nor \U$21250 ( \21593 , \21589 , \21592 );
not \U$21251 ( \21594 , \3406 );
not \U$21252 ( \21595 , \18062 );
or \U$21253 ( \21596 , \21594 , \21595 );
not \U$21254 ( \21597 , RIbb2ebc0_23);
not \U$21255 ( \21598 , \4698 );
or \U$21256 ( \21599 , \21597 , \21598 );
nand \U$21257 ( \21600 , \15078 , \3396 );
nand \U$21258 ( \21601 , \21599 , \21600 );
nand \U$21259 ( \21602 , \21601 , \3383 );
nand \U$21260 ( \21603 , \21596 , \21602 );
not \U$21261 ( \21604 , \21603 );
and \U$21262 ( \21605 , \21593 , \21604 );
not \U$21263 ( \21606 , \21593 );
and \U$21264 ( \21607 , \21606 , \21603 );
nor \U$21265 ( \21608 , \21605 , \21607 );
not \U$21266 ( \21609 , \21608 );
not \U$21267 ( \21610 , \836 );
not \U$21268 ( \21611 , RIbb2ee90_17);
not \U$21269 ( \21612 , \12211 );
or \U$21270 ( \21613 , \21611 , \21612 );
not \U$21271 ( \21614 , \14025 );
nand \U$21272 ( \21615 , \21614 , \822 );
nand \U$21273 ( \21616 , \21613 , \21615 );
not \U$21274 ( \21617 , \21616 );
or \U$21275 ( \21618 , \21610 , \21617 );
nand \U$21276 ( \21619 , \17084 , \832 );
nand \U$21277 ( \21620 , \21618 , \21619 );
not \U$21278 ( \21621 , \1517 );
not \U$21279 ( \21622 , RIbb2ef80_15);
not \U$21280 ( \21623 , \9279 );
or \U$21281 ( \21624 , \21622 , \21623 );
nand \U$21282 ( \21625 , \16475 , \2356 );
nand \U$21283 ( \21626 , \21624 , \21625 );
not \U$21284 ( \21627 , \21626 );
or \U$21285 ( \21628 , \21621 , \21627 );
not \U$21286 ( \21629 , \1575 );
nand \U$21287 ( \21630 , \21629 , \17037 );
nand \U$21288 ( \21631 , \21628 , \21630 );
and \U$21289 ( \21632 , \21620 , \21631 );
not \U$21290 ( \21633 , \21620 );
not \U$21291 ( \21634 , \21631 );
and \U$21292 ( \21635 , \21633 , \21634 );
nor \U$21293 ( \21636 , \21632 , \21635 );
not \U$21294 ( \21637 , \916 );
not \U$21295 ( \21638 , \17052 );
or \U$21296 ( \21639 , \21637 , \21638 );
not \U$21297 ( \21640 , RIbb2f070_13);
not \U$21298 ( \21641 , \12744 );
or \U$21299 ( \21642 , \21640 , \21641 );
nand \U$21300 ( \21643 , \12235 , \906 );
nand \U$21301 ( \21644 , \21642 , \21643 );
nand \U$21302 ( \21645 , \21644 , \998 );
nand \U$21303 ( \21646 , \21639 , \21645 );
not \U$21304 ( \21647 , \21646 );
xor \U$21305 ( \21648 , \21636 , \21647 );
and \U$21306 ( \21649 , \21609 , \21648 );
not \U$21307 ( \21650 , \21609 );
not \U$21308 ( \21651 , \21648 );
and \U$21309 ( \21652 , \21650 , \21651 );
or \U$21310 ( \21653 , \21649 , \21652 );
not \U$21311 ( \21654 , \16256 );
not \U$21312 ( \21655 , \21654 );
not \U$21313 ( \21656 , \16270 );
not \U$21314 ( \21657 , \21656 );
or \U$21315 ( \21658 , \21655 , \21657 );
nand \U$21316 ( \21659 , \21658 , RIbb2dae0_59);
not \U$21317 ( \21660 , \18093 );
nor \U$21318 ( \21661 , \21660 , \1392 );
xor \U$21319 ( \21662 , \21659 , \21661 );
not \U$21320 ( \21663 , \1375 );
not \U$21321 ( \21664 , \1393 );
buf \U$21322 ( \21665 , \16567 );
not \U$21323 ( \21666 , \21665 );
or \U$21324 ( \21667 , \21664 , \21666 );
nand \U$21325 ( \21668 , \16566 , \1392 );
nand \U$21326 ( \21669 , \21667 , \21668 );
not \U$21327 ( \21670 , \21669 );
or \U$21328 ( \21671 , \21663 , \21670 );
nand \U$21329 ( \21672 , \1428 , \19199 );
nand \U$21330 ( \21673 , \21671 , \21672 );
xor \U$21331 ( \21674 , \21662 , \21673 );
not \U$21332 ( \21675 , \12965 );
and \U$21333 ( \21676 , \3368 , RIbb2e080_47);
not \U$21334 ( \21677 , \3368 );
and \U$21335 ( \21678 , \21677 , \16171 );
or \U$21336 ( \21679 , \21676 , \21678 );
not \U$21337 ( \21680 , \21679 );
or \U$21338 ( \21681 , \21675 , \21680 );
nand \U$21339 ( \21682 , \18117 , \11176 );
nand \U$21340 ( \21683 , \21681 , \21682 );
xor \U$21341 ( \21684 , \21674 , \21683 );
not \U$21342 ( \21685 , \2941 );
not \U$21343 ( \21686 , RIbb2e800_31);
not \U$21344 ( \21687 , \6173 );
or \U$21345 ( \21688 , \21686 , \21687 );
nand \U$21346 ( \21689 , \13903 , \2917 );
nand \U$21347 ( \21690 , \21688 , \21689 );
not \U$21348 ( \21691 , \21690 );
or \U$21349 ( \21692 , \21685 , \21691 );
nand \U$21350 ( \21693 , \18130 , \2940 );
nand \U$21351 ( \21694 , \21692 , \21693 );
xor \U$21352 ( \21695 , \21684 , \21694 );
buf \U$21353 ( \21696 , \21695 );
xor \U$21354 ( \21697 , \21653 , \21696 );
xor \U$21355 ( \21698 , \21567 , \21697 );
buf \U$21356 ( \21699 , \19241 );
not \U$21357 ( \21700 , \21699 );
nand \U$21358 ( \21701 , \21700 , \19211 );
not \U$21359 ( \21702 , \21701 );
not \U$21360 ( \21703 , \19247 );
or \U$21361 ( \21704 , \21702 , \21703 );
not \U$21362 ( \21705 , \19211 );
nand \U$21363 ( \21706 , \21705 , \21699 );
nand \U$21364 ( \21707 , \21704 , \21706 );
not \U$21365 ( \21708 , \17089 );
not \U$21366 ( \21709 , \17126 );
or \U$21367 ( \21710 , \21708 , \21709 );
or \U$21368 ( \21711 , \17126 , \17089 );
not \U$21369 ( \21712 , \17056 );
nand \U$21370 ( \21713 , \21711 , \21712 );
nand \U$21371 ( \21714 , \21710 , \21713 );
xor \U$21372 ( \21715 , \21707 , \21714 );
xor \U$21373 ( \21716 , \17166 , \17203 );
and \U$21374 ( \21717 , \21716 , \17240 );
and \U$21375 ( \21718 , \17166 , \17203 );
or \U$21376 ( \21719 , \21717 , \21718 );
xnor \U$21377 ( \21720 , \21715 , \21719 );
and \U$21378 ( \21721 , \21698 , \21720 );
not \U$21379 ( \21722 , \21698 );
not \U$21380 ( \21723 , \21720 );
and \U$21381 ( \21724 , \21722 , \21723 );
or \U$21382 ( \21725 , \21721 , \21724 );
xor \U$21383 ( \21726 , \18158 , \18199 );
and \U$21384 ( \21727 , \21726 , \18231 );
and \U$21385 ( \21728 , \18158 , \18199 );
or \U$21386 ( \21729 , \21727 , \21728 );
or \U$21387 ( \21730 , \18210 , \18230 );
nand \U$21388 ( \21731 , \21730 , \18220 );
nand \U$21389 ( \21732 , \18230 , \18210 );
nand \U$21390 ( \21733 , \21731 , \21732 );
not \U$21391 ( \21734 , \18168 );
not \U$21392 ( \21735 , \21734 );
not \U$21393 ( \21736 , \18190 );
or \U$21394 ( \21737 , \21735 , \21736 );
not \U$21395 ( \21738 , \18168 );
not \U$21396 ( \21739 , \18193 );
or \U$21397 ( \21740 , \21738 , \21739 );
nand \U$21398 ( \21741 , \21740 , \18180 );
nand \U$21399 ( \21742 , \21737 , \21741 );
xor \U$21400 ( \21743 , \21733 , \21742 );
xor \U$21401 ( \21744 , \18279 , \18289 );
and \U$21402 ( \21745 , \21744 , \18302 );
and \U$21403 ( \21746 , \18279 , \18289 );
or \U$21404 ( \21747 , \21745 , \21746 );
not \U$21405 ( \21748 , \21747 );
and \U$21406 ( \21749 , \21743 , \21748 );
not \U$21407 ( \21750 , \21743 );
and \U$21408 ( \21751 , \21750 , \21747 );
nor \U$21409 ( \21752 , \21749 , \21751 );
xor \U$21410 ( \21753 , \21729 , \21752 );
not \U$21411 ( \21754 , \1737 );
not \U$21412 ( \21755 , RIbb2f340_7);
not \U$21413 ( \21756 , \14843 );
not \U$21414 ( \21757 , \21756 );
or \U$21415 ( \21758 , \21755 , \21757 );
nand \U$21416 ( \21759 , \14844 , \1692 );
nand \U$21417 ( \21760 , \21758 , \21759 );
not \U$21418 ( \21761 , \21760 );
or \U$21419 ( \21762 , \21754 , \21761 );
nand \U$21420 ( \21763 , \19216 , \1702 );
nand \U$21421 ( \21764 , \21762 , \21763 );
xor \U$21422 ( \21765 , \19201 , \21764 );
not \U$21423 ( \21766 , \1264 );
not \U$21424 ( \21767 , \19236 );
or \U$21425 ( \21768 , \21766 , \21767 );
not \U$21426 ( \21769 , \1288 );
not \U$21427 ( \21770 , \14527 );
not \U$21428 ( \21771 , \21770 );
or \U$21429 ( \21772 , \21769 , \21771 );
nand \U$21430 ( \21773 , \15036 , \1244 );
nand \U$21431 ( \21774 , \21772 , \21773 );
nand \U$21432 ( \21775 , \21774 , \1294 );
nand \U$21433 ( \21776 , \21768 , \21775 );
xor \U$21434 ( \21777 , \21765 , \21776 );
not \U$21435 ( \21778 , \18342 );
not \U$21436 ( \21779 , \18325 );
or \U$21437 ( \21780 , \21778 , \21779 );
nand \U$21438 ( \21781 , \21780 , \18314 );
nand \U$21439 ( \21782 , \18339 , \18324 );
nand \U$21440 ( \21783 , \21781 , \21782 );
xor \U$21441 ( \21784 , \21777 , \21783 );
xor \U$21442 ( \21785 , \18247 , \18257 );
and \U$21443 ( \21786 , \21785 , \18268 );
and \U$21444 ( \21787 , \18247 , \18257 );
or \U$21445 ( \21788 , \21786 , \21787 );
xor \U$21446 ( \21789 , \21784 , \21788 );
xor \U$21447 ( \21790 , \21753 , \21789 );
buf \U$21448 ( \21791 , \21790 );
xnor \U$21449 ( \21792 , \21725 , \21791 );
not \U$21450 ( \21793 , \18134 );
not \U$21451 ( \21794 , \18141 );
not \U$21452 ( \21795 , \21794 );
or \U$21453 ( \21796 , \21793 , \21795 );
nand \U$21454 ( \21797 , \21796 , \18149 );
not \U$21455 ( \21798 , \18134 );
nand \U$21456 ( \21799 , \21798 , \18141 );
nand \U$21457 ( \21800 , \21797 , \21799 );
xor \U$21458 ( \21801 , \18232 , \18345 );
and \U$21459 ( \21802 , \21801 , \18464 );
and \U$21460 ( \21803 , \18232 , \18345 );
or \U$21461 ( \21804 , \21802 , \21803 );
xor \U$21462 ( \21805 , \21800 , \21804 );
xor \U$21463 ( \21806 , \18111 , \18121 );
and \U$21464 ( \21807 , \21806 , \18132 );
and \U$21465 ( \21808 , \18111 , \18121 );
or \U$21466 ( \21809 , \21807 , \21808 );
not \U$21467 ( \21810 , \1011 );
not \U$21468 ( \21811 , \18238 );
or \U$21469 ( \21812 , \21810 , \21811 );
not \U$21470 ( \21813 , RIbb2f160_11);
not \U$21471 ( \21814 , \12756 );
or \U$21472 ( \21815 , \21813 , \21814 );
nand \U$21473 ( \21816 , \11144 , \1043 );
nand \U$21474 ( \21817 , \21815 , \21816 );
nand \U$21475 ( \21818 , \21817 , \1077 );
nand \U$21476 ( \21819 , \21812 , \21818 );
not \U$21477 ( \21820 , \2925 );
not \U$21478 ( \21821 , RIbb2e8f0_29);
not \U$21479 ( \21822 , \3021 );
or \U$21480 ( \21823 , \21821 , \21822 );
nand \U$21481 ( \21824 , \10095 , \3440 );
nand \U$21482 ( \21825 , \21823 , \21824 );
not \U$21483 ( \21826 , \21825 );
or \U$21484 ( \21827 , \21820 , \21826 );
nand \U$21485 ( \21828 , \18255 , \2922 );
nand \U$21486 ( \21829 , \21827 , \21828 );
xor \U$21487 ( \21830 , \21819 , \21829 );
not \U$21488 ( \21831 , \10119 );
not \U$21489 ( \21832 , RIbb2e170_45);
not \U$21490 ( \21833 , \7424 );
or \U$21491 ( \21834 , \21832 , \21833 );
nand \U$21492 ( \21835 , \10673 , \9094 );
nand \U$21493 ( \21836 , \21834 , \21835 );
not \U$21494 ( \21837 , \21836 );
or \U$21495 ( \21838 , \21831 , \21837 );
nand \U$21496 ( \21839 , \18266 , \10117 );
nand \U$21497 ( \21840 , \21838 , \21839 );
xor \U$21498 ( \21841 , \21830 , \21840 );
xor \U$21499 ( \21842 , \21809 , \21841 );
not \U$21500 ( \21843 , \12285 );
and \U$21501 ( \21844 , \1549 , RIbb2df90_49);
not \U$21502 ( \21845 , \1549 );
and \U$21503 ( \21846 , \21845 , \12278 );
or \U$21504 ( \21847 , \21844 , \21846 );
not \U$21505 ( \21848 , \21847 );
or \U$21506 ( \21849 , \21843 , \21848 );
nand \U$21507 ( \21850 , \18287 , \12167 );
nand \U$21508 ( \21851 , \21849 , \21850 );
not \U$21509 ( \21852 , \4712 );
not \U$21510 ( \21853 , \18275 );
or \U$21511 ( \21854 , \21852 , \21853 );
not \U$21512 ( \21855 , RIbb2e620_35);
not \U$21513 ( \21856 , \3517 );
or \U$21514 ( \21857 , \21855 , \21856 );
nand \U$21515 ( \21858 , \12096 , \3866 );
nand \U$21516 ( \21859 , \21857 , \21858 );
nand \U$21517 ( \21860 , \5845 , \21859 );
nand \U$21518 ( \21861 , \21854 , \21860 );
not \U$21519 ( \21862 , \21861 );
xor \U$21520 ( \21863 , \21851 , \21862 );
not \U$21521 ( \21864 , \3887 );
nor \U$21522 ( \21865 , \21864 , \18297 );
not \U$21523 ( \21866 , RIbb2e710_33);
not \U$21524 ( \21867 , \6301 );
or \U$21525 ( \21868 , \21866 , \21867 );
nand \U$21526 ( \21869 , \3139 , \3877 );
nand \U$21527 ( \21870 , \21868 , \21869 );
not \U$21528 ( \21871 , \21870 );
nor \U$21529 ( \21872 , \21871 , \3871 );
nor \U$21530 ( \21873 , \21865 , \21872 );
not \U$21531 ( \21874 , \21873 );
not \U$21532 ( \21875 , \21874 );
xor \U$21533 ( \21876 , \21863 , \21875 );
xor \U$21534 ( \21877 , \21842 , \21876 );
not \U$21535 ( \21878 , \12692 );
not \U$21536 ( \21879 , RIbb2dea0_51);
not \U$21537 ( \21880 , \1070 );
or \U$21538 ( \21881 , \21879 , \21880 );
not \U$21539 ( \21882 , RIbb2dea0_51);
nand \U$21540 ( \21883 , \1886 , \21882 );
nand \U$21541 ( \21884 , \21881 , \21883 );
not \U$21542 ( \21885 , \21884 );
or \U$21543 ( \21886 , \21878 , \21885 );
nand \U$21544 ( \21887 , \18208 , \14067 );
nand \U$21545 ( \21888 , \21886 , \21887 );
not \U$21546 ( \21889 , \14930 );
not \U$21547 ( \21890 , RIbb2ddb0_53);
not \U$21548 ( \21891 , \992 );
or \U$21549 ( \21892 , \21890 , \21891 );
nand \U$21550 ( \21893 , \17474 , \12681 );
nand \U$21551 ( \21894 , \21892 , \21893 );
not \U$21552 ( \21895 , \21894 );
or \U$21553 ( \21896 , \21889 , \21895 );
nand \U$21554 ( \21897 , \18216 , \17563 );
nand \U$21555 ( \21898 , \21896 , \21897 );
xor \U$21556 ( \21899 , \21888 , \21898 );
not \U$21557 ( \21900 , \8361 );
not \U$21558 ( \21901 , \18226 );
or \U$21559 ( \21902 , \21900 , \21901 );
not \U$21560 ( \21903 , RIbb2e350_41);
not \U$21561 ( \21904 , \4339 );
or \U$21562 ( \21905 , \21903 , \21904 );
nand \U$21563 ( \21906 , \4340 , \7097 );
nand \U$21564 ( \21907 , \21905 , \21906 );
nand \U$21565 ( \21908 , \21907 , \8995 );
nand \U$21566 ( \21909 , \21902 , \21908 );
xnor \U$21567 ( \21910 , \21899 , \21909 );
not \U$21568 ( \21911 , \6251 );
not \U$21569 ( \21912 , \18185 );
or \U$21570 ( \21913 , \21911 , \21912 );
not \U$21571 ( \21914 , RIbb2e530_37);
not \U$21572 ( \21915 , \3310 );
or \U$21573 ( \21916 , \21914 , \21915 );
nand \U$21574 ( \21917 , \16235 , \6246 );
nand \U$21575 ( \21918 , \21916 , \21917 );
nand \U$21576 ( \21919 , \21918 , \6242 );
nand \U$21577 ( \21920 , \21913 , \21919 );
not \U$21578 ( \21921 , \14613 );
not \U$21579 ( \21922 , \18176 );
or \U$21580 ( \21923 , \21921 , \21922 );
and \U$21581 ( \21924 , RIbb2dcc0_55, \8754 );
not \U$21582 ( \21925 , RIbb2dcc0_55);
and \U$21583 ( \21926 , \21925 , \13308 );
or \U$21584 ( \21927 , \21924 , \21926 );
nand \U$21585 ( \21928 , \21927 , \15181 );
nand \U$21586 ( \21929 , \21923 , \21928 );
xor \U$21587 ( \21930 , \21920 , \21929 );
not \U$21588 ( \21931 , RIbb2e440_39);
not \U$21589 ( \21932 , \3575 );
or \U$21590 ( \21933 , \21931 , \21932 );
not \U$21591 ( \21934 , RIbb2e440_39);
nand \U$21592 ( \21935 , \21934 , \1338 );
nand \U$21593 ( \21936 , \21933 , \21935 );
not \U$21594 ( \21937 , \21936 );
not \U$21595 ( \21938 , \7104 );
or \U$21596 ( \21939 , \21937 , \21938 );
not \U$21597 ( \21940 , \18164 );
nand \U$21598 ( \21941 , \21940 , \8445 );
nand \U$21599 ( \21942 , \21939 , \21941 );
xor \U$21600 ( \21943 , \21930 , \21942 );
xor \U$21601 ( \21944 , \21910 , \21943 );
not \U$21602 ( \21945 , \15746 );
not \U$21603 ( \21946 , \18320 );
or \U$21604 ( \21947 , \21945 , \21946 );
and \U$21605 ( \21948 , \14602 , \812 );
not \U$21606 ( \21949 , \14602 );
and \U$21607 ( \21950 , \21949 , \811 );
nor \U$21608 ( \21951 , \21948 , \21950 );
nand \U$21609 ( \21952 , \21951 , \15738 );
nand \U$21610 ( \21953 , \21947 , \21952 );
not \U$21611 ( \21954 , \10451 );
not \U$21612 ( \21955 , RIbb2e260_43);
not \U$21613 ( \21956 , \12037 );
or \U$21614 ( \21957 , \21955 , \21956 );
nand \U$21615 ( \21958 , \3291 , \10444 );
nand \U$21616 ( \21959 , \21957 , \21958 );
not \U$21617 ( \21960 , \21959 );
or \U$21618 ( \21961 , \21954 , \21960 );
nand \U$21619 ( \21962 , \18312 , \10449 );
nand \U$21620 ( \21963 , \21961 , \21962 );
xor \U$21621 ( \21964 , \21953 , \21963 );
not \U$21622 ( \21965 , \3465 );
not \U$21623 ( \21966 , RIbb2e9e0_27);
not \U$21624 ( \21967 , \4411 );
or \U$21625 ( \21968 , \21966 , \21967 );
nand \U$21626 ( \21969 , \3275 , \4598 );
nand \U$21627 ( \21970 , \21968 , \21969 );
not \U$21628 ( \21971 , \21970 );
or \U$21629 ( \21972 , \21965 , \21971 );
nand \U$21630 ( \21973 , \18335 , \3445 );
nand \U$21631 ( \21974 , \21972 , \21973 );
xor \U$21632 ( \21975 , \21964 , \21974 );
xnor \U$21633 ( \21976 , \21944 , \21975 );
xor \U$21634 ( \21977 , \21877 , \21976 );
xor \U$21635 ( \21978 , \18406 , \18457 );
and \U$21636 ( \21979 , \21978 , \18463 );
and \U$21637 ( \21980 , \18406 , \18457 );
or \U$21638 ( \21981 , \21979 , \21980 );
xor \U$21639 ( \21982 , \21977 , \21981 );
xor \U$21640 ( \21983 , \21805 , \21982 );
xor \U$21641 ( \21984 , \21792 , \21983 );
buf \U$21642 ( \21985 , \18465 );
buf \U$21643 ( \21986 , \18154 );
or \U$21644 ( \21987 , \21985 , \21986 );
nand \U$21645 ( \21988 , \21987 , \18475 );
nand \U$21646 ( \21989 , \21985 , \21986 );
nand \U$21647 ( \21990 , \21988 , \21989 );
xor \U$21648 ( \21991 , \21984 , \21990 );
xor \U$21649 ( \21992 , \19171 , \19293 );
and \U$21650 ( \21993 , \21992 , \19482 );
and \U$21651 ( \21994 , \19171 , \19293 );
or \U$21652 ( \21995 , \21993 , \21994 );
xor \U$21653 ( \21996 , \21991 , \21995 );
xor \U$21654 ( \21997 , \19175 , \19287 );
and \U$21655 ( \21998 , \21997 , \19292 );
and \U$21656 ( \21999 , \19175 , \19287 );
or \U$21657 ( \22000 , \21998 , \21999 );
xor \U$21658 ( \22001 , \19179 , \19281 );
and \U$21659 ( \22002 , \22001 , \19286 );
and \U$21660 ( \22003 , \19179 , \19281 );
or \U$21661 ( \22004 , \22002 , \22003 );
xor \U$21662 ( \22005 , \19251 , \19272 );
and \U$21663 ( \22006 , \22005 , \19280 );
and \U$21664 ( \22007 , \19251 , \19272 );
or \U$21665 ( \22008 , \22006 , \22007 );
not \U$21666 ( \22009 , \17020 );
not \U$21667 ( \22010 , \17241 );
or \U$21668 ( \22011 , \22009 , \22010 );
or \U$21669 ( \22012 , \17020 , \17241 );
nand \U$21670 ( \22013 , \22012 , \17128 );
nand \U$21671 ( \22014 , \22011 , \22013 );
xor \U$21672 ( \22015 , \22008 , \22014 );
xor \U$21673 ( \22016 , \19220 , \19230 );
and \U$21674 ( \22017 , \22016 , \19240 );
and \U$21675 ( \22018 , \19220 , \19230 );
or \U$21676 ( \22019 , \22017 , \22018 );
not \U$21677 ( \22020 , \19203 );
nand \U$21678 ( \22021 , \22020 , \19201 );
not \U$21679 ( \22022 , \22021 );
not \U$21680 ( \22023 , \19189 );
or \U$21681 ( \22024 , \22022 , \22023 );
not \U$21682 ( \22025 , \19201 );
nand \U$21683 ( \22026 , \22025 , \19203 );
nand \U$21684 ( \22027 , \22024 , \22026 );
not \U$21685 ( \22028 , \22027 );
and \U$21686 ( \22029 , \22019 , \22028 );
not \U$21687 ( \22030 , \22019 );
and \U$21688 ( \22031 , \22030 , \22027 );
nor \U$21689 ( \22032 , \22029 , \22031 );
not \U$21690 ( \22033 , \22032 );
xor \U$21691 ( \22034 , \18056 , \18066 );
and \U$21692 ( \22035 , \22034 , \18078 );
and \U$21693 ( \22036 , \18056 , \18066 );
or \U$21694 ( \22037 , \22035 , \22036 );
not \U$21695 ( \22038 , \22037 );
and \U$21696 ( \22039 , \22033 , \22038 );
and \U$21697 ( \22040 , \22037 , \22032 );
nor \U$21698 ( \22041 , \22039 , \22040 );
not \U$21699 ( \22042 , \22041 );
not \U$21700 ( \22043 , \22042 );
xor \U$21701 ( \22044 , \19255 , \19262 );
and \U$21702 ( \22045 , \22044 , \19271 );
and \U$21703 ( \22046 , \19255 , \19262 );
or \U$21704 ( \22047 , \22045 , \22046 );
not \U$21705 ( \22048 , \22047 );
not \U$21706 ( \22049 , \22048 );
or \U$21707 ( \22050 , \22043 , \22049 );
nand \U$21708 ( \22051 , \22047 , \22041 );
nand \U$21709 ( \22052 , \22050 , \22051 );
xor \U$21710 ( \22053 , \17066 , \17076 );
and \U$21711 ( \22054 , \22053 , \17088 );
and \U$21712 ( \22055 , \17066 , \17076 );
or \U$21713 ( \22056 , \22054 , \22055 );
not \U$21714 ( \22057 , \1147 );
not \U$21715 ( \22058 , RIbb2f430_5);
not \U$21716 ( \22059 , \13986 );
or \U$21717 ( \22060 , \22058 , \22059 );
not \U$21718 ( \22061 , \15054 );
nand \U$21719 ( \22062 , \22061 , \1647 );
nand \U$21720 ( \22063 , \22060 , \22062 );
not \U$21721 ( \22064 , \22063 );
or \U$21722 ( \22065 , \22057 , \22064 );
nand \U$21723 ( \22066 , \19226 , \1089 );
nand \U$21724 ( \22067 , \22065 , \22066 );
not \U$21725 ( \22068 , \1570 );
not \U$21726 ( \22069 , RIbb2f250_9);
not \U$21727 ( \22070 , \12175 );
not \U$21728 ( \22071 , \22070 );
or \U$21729 ( \22072 , \22069 , \22071 );
buf \U$21730 ( \22073 , \12175 );
nand \U$21731 ( \22074 , \22073 , \1566 );
nand \U$21732 ( \22075 , \22072 , \22074 );
not \U$21733 ( \22076 , \22075 );
or \U$21734 ( \22077 , \22068 , \22076 );
nand \U$21735 ( \22078 , \19185 , \1533 );
nand \U$21736 ( \22079 , \22077 , \22078 );
xor \U$21737 ( \22080 , \22067 , \22079 );
not \U$21738 ( \22081 , \2963 );
and \U$21739 ( \22082 , RIbb2ead0_25, \4325 );
not \U$21740 ( \22083 , RIbb2ead0_25);
and \U$21741 ( \22084 , \22083 , \4324 );
or \U$21742 ( \22085 , \22082 , \22084 );
not \U$21743 ( \22086 , \22085 );
or \U$21744 ( \22087 , \22081 , \22086 );
nand \U$21745 ( \22088 , \18074 , \2980 );
nand \U$21746 ( \22089 , \22087 , \22088 );
xor \U$21747 ( \22090 , \22080 , \22089 );
xor \U$21748 ( \22091 , \22056 , \22090 );
not \U$21749 ( \22092 , \17032 );
not \U$21750 ( \22093 , \22092 );
not \U$21751 ( \22094 , \17055 );
or \U$21752 ( \22095 , \22093 , \22094 );
nand \U$21753 ( \22096 , \22095 , \17043 );
nand \U$21754 ( \22097 , \17054 , \17032 );
nand \U$21755 ( \22098 , \22096 , \22097 );
xor \U$21756 ( \22099 , \22091 , \22098 );
not \U$21757 ( \22100 , \22099 );
and \U$21758 ( \22101 , \22052 , \22100 );
not \U$21759 ( \22102 , \22052 );
and \U$21760 ( \22103 , \22102 , \22099 );
nor \U$21761 ( \22104 , \22101 , \22103 );
not \U$21762 ( \22105 , \22104 );
xor \U$21763 ( \22106 , \22015 , \22105 );
xor \U$21764 ( \22107 , \22004 , \22106 );
xor \U$21765 ( \22108 , \16625 , \17011 );
and \U$21766 ( \22109 , \22108 , \17246 );
and \U$21767 ( \22110 , \16625 , \17011 );
or \U$21768 ( \22111 , \22109 , \22110 );
xor \U$21769 ( \22112 , \22107 , \22111 );
xor \U$21770 ( \22113 , \22000 , \22112 );
not \U$21771 ( \22114 , \17247 );
not \U$21772 ( \22115 , \22114 );
not \U$21773 ( \22116 , \18479 );
or \U$21774 ( \22117 , \22115 , \22116 );
nand \U$21775 ( \22118 , \22117 , \18051 );
not \U$21776 ( \22119 , \22114 );
nand \U$21777 ( \22120 , \22119 , \18480 );
nand \U$21778 ( \22121 , \22118 , \22120 );
xor \U$21779 ( \22122 , \22113 , \22121 );
xor \U$21780 ( \22123 , \21996 , \22122 );
nor \U$21781 ( \22124 , \21558 , \22123 );
xor \U$21782 ( \22125 , \21792 , \21983 );
and \U$21783 ( \22126 , \22125 , \21990 );
and \U$21784 ( \22127 , \21792 , \21983 );
or \U$21785 ( \22128 , \22126 , \22127 );
xor \U$21786 ( \22129 , \22000 , \22112 );
and \U$21787 ( \22130 , \22129 , \22121 );
and \U$21788 ( \22131 , \22000 , \22112 );
or \U$21789 ( \22132 , \22130 , \22131 );
xor \U$21790 ( \22133 , \22128 , \22132 );
not \U$21791 ( \22134 , \21790 );
not \U$21792 ( \22135 , \22134 );
not \U$21793 ( \22136 , \21723 );
or \U$21794 ( \22137 , \22135 , \22136 );
not \U$21795 ( \22138 , \21720 );
not \U$21796 ( \22139 , \21790 );
or \U$21797 ( \22140 , \22138 , \22139 );
nand \U$21798 ( \22141 , \22140 , \21698 );
nand \U$21799 ( \22142 , \22137 , \22141 );
xor \U$21800 ( \22143 , \21800 , \21804 );
and \U$21801 ( \22144 , \22143 , \21982 );
and \U$21802 ( \22145 , \21800 , \21804 );
or \U$21803 ( \22146 , \22144 , \22145 );
xor \U$21804 ( \22147 , \22142 , \22146 );
not \U$21805 ( \22148 , \21975 );
not \U$21806 ( \22149 , \21943 );
or \U$21807 ( \22150 , \22148 , \22149 );
or \U$21808 ( \22151 , \21975 , \21943 );
not \U$21809 ( \22152 , \21910 );
nand \U$21810 ( \22153 , \22151 , \22152 );
nand \U$21811 ( \22154 , \22150 , \22153 );
not \U$21812 ( \22155 , \21942 );
not \U$21813 ( \22156 , \21920 );
or \U$21814 ( \22157 , \22155 , \22156 );
or \U$21815 ( \22158 , \21920 , \21942 );
nand \U$21816 ( \22159 , \22158 , \21929 );
nand \U$21817 ( \22160 , \22157 , \22159 );
not \U$21818 ( \22161 , \21861 );
not \U$21819 ( \22162 , \21874 );
or \U$21820 ( \22163 , \22161 , \22162 );
not \U$21821 ( \22164 , \21873 );
not \U$21822 ( \22165 , \21862 );
or \U$21823 ( \22166 , \22164 , \22165 );
nand \U$21824 ( \22167 , \22166 , \21851 );
nand \U$21825 ( \22168 , \22163 , \22167 );
and \U$21826 ( \22169 , \22160 , \22168 );
not \U$21827 ( \22170 , \22160 );
not \U$21828 ( \22171 , \22168 );
and \U$21829 ( \22172 , \22170 , \22171 );
nor \U$21830 ( \22173 , \22169 , \22172 );
xor \U$21831 ( \22174 , \21953 , \21963 );
and \U$21832 ( \22175 , \22174 , \21974 );
and \U$21833 ( \22176 , \21953 , \21963 );
or \U$21834 ( \22177 , \22175 , \22176 );
not \U$21835 ( \22178 , \22177 );
and \U$21836 ( \22179 , \22173 , \22178 );
not \U$21837 ( \22180 , \22173 );
and \U$21838 ( \22181 , \22180 , \22177 );
nor \U$21839 ( \22182 , \22179 , \22181 );
or \U$21840 ( \22183 , \22154 , \22182 );
nand \U$21841 ( \22184 , \22182 , \22154 );
nand \U$21842 ( \22185 , \22183 , \22184 );
xor \U$21843 ( \22186 , \21809 , \21841 );
and \U$21844 ( \22187 , \22186 , \21876 );
and \U$21845 ( \22188 , \21809 , \21841 );
or \U$21846 ( \22189 , \22187 , \22188 );
and \U$21847 ( \22190 , \22185 , \22189 );
not \U$21848 ( \22191 , \22185 );
not \U$21849 ( \22192 , \22189 );
and \U$21850 ( \22193 , \22191 , \22192 );
nor \U$21851 ( \22194 , \22190 , \22193 );
xor \U$21852 ( \22195 , \21877 , \21976 );
and \U$21853 ( \22196 , \22195 , \21981 );
and \U$21854 ( \22197 , \21877 , \21976 );
or \U$21855 ( \22198 , \22196 , \22197 );
xor \U$21856 ( \22199 , \22194 , \22198 );
xor \U$21857 ( \22200 , \21659 , \21661 );
and \U$21858 ( \22201 , \22200 , \21673 );
and \U$21859 ( \22202 , \21659 , \21661 );
or \U$21860 ( \22203 , \22201 , \22202 );
not \U$21861 ( \22204 , \853 );
not \U$21862 ( \22205 , \21584 );
or \U$21863 ( \22206 , \22204 , \22205 );
nand \U$21864 ( \22207 , \15801 , \854 );
nand \U$21865 ( \22208 , \22206 , \22207 );
xor \U$21866 ( \22209 , \22203 , \22208 );
not \U$21867 ( \22210 , \2077 );
not \U$21868 ( \22211 , \21574 );
or \U$21869 ( \22212 , \22210 , \22211 );
nand \U$21870 ( \22213 , \15843 , \2078 );
nand \U$21871 ( \22214 , \22212 , \22213 );
xor \U$21872 ( \22215 , \22209 , \22214 );
not \U$21873 ( \22216 , \15181 );
not \U$21874 ( \22217 , RIbb2dcc0_55);
not \U$21875 ( \22218 , \12969 );
or \U$21876 ( \22219 , \22217 , \22218 );
not \U$21877 ( \22220 , RIbb2dcc0_55);
nand \U$21878 ( \22221 , \22220 , \892 );
nand \U$21879 ( \22222 , \22219 , \22221 );
not \U$21880 ( \22223 , \22222 );
or \U$21881 ( \22224 , \22216 , \22223 );
nand \U$21882 ( \22225 , \21927 , \14613 );
nand \U$21883 ( \22226 , \22224 , \22225 );
not \U$21884 ( \22227 , \12692 );
and \U$21885 ( \22228 , RIbb2dea0_51, \951 );
not \U$21886 ( \22229 , RIbb2dea0_51);
and \U$21887 ( \22230 , \22229 , \956 );
or \U$21888 ( \22231 , \22228 , \22230 );
not \U$21889 ( \22232 , \22231 );
or \U$21890 ( \22233 , \22227 , \22232 );
nand \U$21891 ( \22234 , \21884 , \14067 );
nand \U$21892 ( \22235 , \22233 , \22234 );
xor \U$21893 ( \22236 , \22226 , \22235 );
not \U$21894 ( \22237 , \8361 );
not \U$21895 ( \22238 , \21907 );
or \U$21896 ( \22239 , \22237 , \22238 );
not \U$21897 ( \22240 , RIbb2e350_41);
not \U$21898 ( \22241 , \3990 );
or \U$21899 ( \22242 , \22240 , \22241 );
nand \U$21900 ( \22243 , \1169 , \9402 );
nand \U$21901 ( \22244 , \22242 , \22243 );
nand \U$21902 ( \22245 , \22244 , \8995 );
nand \U$21903 ( \22246 , \22239 , \22245 );
xnor \U$21904 ( \22247 , \22236 , \22246 );
xor \U$21905 ( \22248 , \22215 , \22247 );
not \U$21906 ( \22249 , \10599 );
not \U$21907 ( \22250 , \21836 );
or \U$21908 ( \22251 , \22249 , \22250 );
not \U$21909 ( \22252 , RIbb2e170_45);
not \U$21910 ( \22253 , \3238 );
or \U$21911 ( \22254 , \22252 , \22253 );
nand \U$21912 ( \22255 , \3243 , \9094 );
nand \U$21913 ( \22256 , \22254 , \22255 );
nand \U$21914 ( \22257 , \22256 , \10119 );
nand \U$21915 ( \22258 , \22251 , \22257 );
not \U$21916 ( \22259 , \22258 );
not \U$21917 ( \22260 , \3887 );
not \U$21918 ( \22261 , \21870 );
or \U$21919 ( \22262 , \22260 , \22261 );
not \U$21920 ( \22263 , \3871 );
not \U$21921 ( \22264 , RIbb2e710_33);
not \U$21922 ( \22265 , \13414 );
or \U$21923 ( \22266 , \22264 , \22265 );
nand \U$21924 ( \22267 , \6108 , \12019 );
nand \U$21925 ( \22268 , \22266 , \22267 );
nand \U$21926 ( \22269 , \22263 , \22268 );
nand \U$21927 ( \22270 , \22262 , \22269 );
not \U$21928 ( \22271 , \22270 );
not \U$21929 ( \22272 , \22271 );
or \U$21930 ( \22273 , \22259 , \22272 );
or \U$21931 ( \22274 , \22271 , \22258 );
nand \U$21932 ( \22275 , \22273 , \22274 );
not \U$21933 ( \22276 , \22275 );
not \U$21934 ( \22277 , \2940 );
not \U$21935 ( \22278 , \21690 );
or \U$21936 ( \22279 , \22277 , \22278 );
not \U$21937 ( \22280 , RIbb2e800_31);
not \U$21938 ( \22281 , \4638 );
or \U$21939 ( \22282 , \22280 , \22281 );
nand \U$21940 ( \22283 , \4637 , \11975 );
nand \U$21941 ( \22284 , \22282 , \22283 );
nand \U$21942 ( \22285 , \22284 , \3613 );
nand \U$21943 ( \22286 , \22279 , \22285 );
not \U$21944 ( \22287 , \22286 );
not \U$21945 ( \22288 , \22287 );
and \U$21946 ( \22289 , \22276 , \22288 );
and \U$21947 ( \22290 , \22275 , \22287 );
nor \U$21948 ( \22291 , \22289 , \22290 );
not \U$21949 ( \22292 , \22291 );
xnor \U$21950 ( \22293 , \22248 , \22292 );
not \U$21951 ( \22294 , \13295 );
not \U$21952 ( \22295 , \21847 );
or \U$21953 ( \22296 , \22294 , \22295 );
not \U$21954 ( \22297 , RIbb2df90_49);
not \U$21955 ( \22298 , \17407 );
or \U$21956 ( \22299 , \22297 , \22298 );
nand \U$21957 ( \22300 , \1560 , \12278 );
nand \U$21958 ( \22301 , \22299 , \22300 );
nand \U$21959 ( \22302 , \22301 , \16427 );
nand \U$21960 ( \22303 , \22296 , \22302 );
not \U$21961 ( \22304 , \7104 );
and \U$21962 ( \22305 , RIbb2e440_39, \17386 );
not \U$21963 ( \22306 , RIbb2e440_39);
and \U$21964 ( \22307 , \22306 , \3821 );
or \U$21965 ( \22308 , \22305 , \22307 );
not \U$21966 ( \22309 , \22308 );
or \U$21967 ( \22310 , \22304 , \22309 );
nand \U$21968 ( \22311 , \21936 , \7103 );
nand \U$21969 ( \22312 , \22310 , \22311 );
not \U$21970 ( \22313 , \22312 );
xnor \U$21971 ( \22314 , \22303 , \22313 );
and \U$21972 ( \22315 , \21918 , \6251 );
not \U$21973 ( \22316 , RIbb2e530_37);
not \U$21974 ( \22317 , \3807 );
or \U$21975 ( \22318 , \22316 , \22317 );
not \U$21976 ( \22319 , \20325 );
nand \U$21977 ( \22320 , \22319 , \4708 );
nand \U$21978 ( \22321 , \22318 , \22320 );
and \U$21979 ( \22322 , \22321 , \6242 );
nor \U$21980 ( \22323 , \22315 , \22322 );
and \U$21981 ( \22324 , \22314 , \22323 );
not \U$21982 ( \22325 , \22314 );
not \U$21983 ( \22326 , \22323 );
and \U$21984 ( \22327 , \22325 , \22326 );
or \U$21985 ( \22328 , \22324 , \22327 );
not \U$21986 ( \22329 , \17563 );
not \U$21987 ( \22330 , \21894 );
or \U$21988 ( \22331 , \22329 , \22330 );
not \U$21989 ( \22332 , RIbb2ddb0_53);
not \U$21990 ( \22333 , \1475 );
or \U$21991 ( \22334 , \22332 , \22333 );
nand \U$21992 ( \22335 , \1474 , \12681 );
nand \U$21993 ( \22336 , \22334 , \22335 );
nand \U$21994 ( \22337 , \22336 , \14930 );
nand \U$21995 ( \22338 , \22331 , \22337 );
not \U$21996 ( \22339 , \4712 );
not \U$21997 ( \22340 , \21859 );
or \U$21998 ( \22341 , \22339 , \22340 );
not \U$21999 ( \22342 , RIbb2e620_35);
not \U$22000 ( \22343 , \13289 );
or \U$22001 ( \22344 , \22342 , \22343 );
not \U$22002 ( \22345 , \2223 );
nand \U$22003 ( \22346 , \22345 , \6002 );
nand \U$22004 ( \22347 , \22344 , \22346 );
nand \U$22005 ( \22348 , \22347 , \5845 );
nand \U$22006 ( \22349 , \22341 , \22348 );
xor \U$22007 ( \22350 , \22338 , \22349 );
not \U$22008 ( \22351 , \11176 );
not \U$22009 ( \22352 , \21679 );
or \U$22010 ( \22353 , \22351 , \22352 );
not \U$22011 ( \22354 , RIbb2e080_47);
not \U$22012 ( \22355 , \5130 );
or \U$22013 ( \22356 , \22354 , \22355 );
not \U$22014 ( \22357 , RIbb2e080_47);
nand \U$22015 ( \22358 , \1730 , \22357 );
nand \U$22016 ( \22359 , \22356 , \22358 );
nand \U$22017 ( \22360 , \22359 , \12965 );
nand \U$22018 ( \22361 , \22353 , \22360 );
buf \U$22019 ( \22362 , \22361 );
xor \U$22020 ( \22363 , \22350 , \22362 );
xor \U$22021 ( \22364 , \22328 , \22363 );
not \U$22022 ( \22365 , \2963 );
and \U$22023 ( \22366 , RIbb2ead0_25, \4748 );
not \U$22024 ( \22367 , RIbb2ead0_25);
and \U$22025 ( \22368 , \22367 , \13750 );
or \U$22026 ( \22369 , \22366 , \22368 );
not \U$22027 ( \22370 , \22369 );
or \U$22028 ( \22371 , \22365 , \22370 );
nand \U$22029 ( \22372 , \22085 , \2980 );
nand \U$22030 ( \22373 , \22371 , \22372 );
not \U$22031 ( \22374 , \3445 );
not \U$22032 ( \22375 , \21970 );
or \U$22033 ( \22376 , \22374 , \22375 );
not \U$22034 ( \22377 , RIbb2e9e0_27);
not \U$22035 ( \22378 , \3045 );
or \U$22036 ( \22379 , \22377 , \22378 );
nand \U$22037 ( \22380 , \16185 , \3454 );
nand \U$22038 ( \22381 , \22379 , \22380 );
nand \U$22039 ( \22382 , \22381 , \3465 );
nand \U$22040 ( \22383 , \22376 , \22382 );
xor \U$22041 ( \22384 , \22373 , \22383 );
not \U$22042 ( \22385 , \10449 );
not \U$22043 ( \22386 , \21959 );
or \U$22044 ( \22387 , \22385 , \22386 );
not \U$22045 ( \22388 , RIbb2e260_43);
not \U$22046 ( \22389 , \3066 );
or \U$22047 ( \22390 , \22388 , \22389 );
not \U$22048 ( \22391 , \13707 );
nand \U$22049 ( \22392 , \22391 , \10444 );
nand \U$22050 ( \22393 , \22390 , \22392 );
nand \U$22051 ( \22394 , \22393 , \9099 );
nand \U$22052 ( \22395 , \22387 , \22394 );
xor \U$22053 ( \22396 , \22384 , \22395 );
xor \U$22054 ( \22397 , \22364 , \22396 );
xor \U$22055 ( \22398 , \22293 , \22397 );
or \U$22056 ( \22399 , \21719 , \21714 );
nand \U$22057 ( \22400 , \22399 , \21707 );
nand \U$22058 ( \22401 , \21719 , \21714 );
nand \U$22059 ( \22402 , \22400 , \22401 );
xor \U$22060 ( \22403 , \22398 , \22402 );
xor \U$22061 ( \22404 , \22199 , \22403 );
xnor \U$22062 ( \22405 , \22147 , \22404 );
not \U$22063 ( \22406 , \22405 );
xor \U$22064 ( \22407 , \22004 , \22106 );
and \U$22065 ( \22408 , \22407 , \22111 );
and \U$22066 ( \22409 , \22004 , \22106 );
or \U$22067 ( \22410 , \22408 , \22409 );
not \U$22068 ( \22411 , \22410 );
not \U$22069 ( \22412 , \22411 );
not \U$22070 ( \22413 , \22008 );
not \U$22071 ( \22414 , \22413 );
not \U$22072 ( \22415 , \22104 );
or \U$22073 ( \22416 , \22414 , \22415 );
nand \U$22074 ( \22417 , \22416 , \22014 );
nand \U$22075 ( \22418 , \22105 , \22008 );
and \U$22076 ( \22419 , \22417 , \22418 );
not \U$22077 ( \22420 , \22041 );
not \U$22078 ( \22421 , \22048 );
or \U$22079 ( \22422 , \22420 , \22421 );
nand \U$22080 ( \22423 , \22422 , \22099 );
nand \U$22081 ( \22424 , \22047 , \22042 );
nand \U$22082 ( \22425 , \22423 , \22424 );
xor \U$22083 ( \22426 , \19201 , \21764 );
and \U$22084 ( \22427 , \22426 , \21776 );
and \U$22085 ( \22428 , \19201 , \21764 );
or \U$22086 ( \22429 , \22427 , \22428 );
not \U$22087 ( \22430 , \2925 );
not \U$22088 ( \22431 , RIbb2e8f0_29);
not \U$22089 ( \22432 , \12707 );
or \U$22090 ( \22433 , \22431 , \22432 );
nand \U$22091 ( \22434 , \3654 , \3265 );
nand \U$22092 ( \22435 , \22433 , \22434 );
not \U$22093 ( \22436 , \22435 );
or \U$22094 ( \22437 , \22430 , \22436 );
nand \U$22095 ( \22438 , \21825 , \2922 );
nand \U$22096 ( \22439 , \22437 , \22438 );
xor \U$22097 ( \22440 , \22429 , \22439 );
xor \U$22098 ( \22441 , \22067 , \22079 );
and \U$22099 ( \22442 , \22441 , \22089 );
and \U$22100 ( \22443 , \22067 , \22079 );
or \U$22101 ( \22444 , \22442 , \22443 );
xor \U$22102 ( \22445 , \22440 , \22444 );
not \U$22103 ( \22446 , \22019 );
nand \U$22104 ( \22447 , \22446 , \22028 );
not \U$22105 ( \22448 , \22447 );
not \U$22106 ( \22449 , \22037 );
or \U$22107 ( \22450 , \22448 , \22449 );
nand \U$22108 ( \22451 , \22019 , \22027 );
nand \U$22109 ( \22452 , \22450 , \22451 );
xor \U$22110 ( \22453 , \22445 , \22452 );
xor \U$22111 ( \22454 , \22056 , \22090 );
and \U$22112 ( \22455 , \22454 , \22098 );
and \U$22113 ( \22456 , \22056 , \22090 );
or \U$22114 ( \22457 , \22455 , \22456 );
xor \U$22115 ( \22458 , \22453 , \22457 );
xor \U$22116 ( \22459 , \22425 , \22458 );
not \U$22117 ( \22460 , \3406 );
not \U$22118 ( \22461 , \21601 );
or \U$22119 ( \22462 , \22460 , \22461 );
nand \U$22120 ( \22463 , \15834 , \3383 );
nand \U$22121 ( \22464 , \22462 , \22463 );
not \U$22122 ( \22465 , \22464 );
not \U$22123 ( \22466 , \1264 );
not \U$22124 ( \22467 , \21774 );
or \U$22125 ( \22468 , \22466 , \22467 );
nand \U$22126 ( \22469 , \15460 , \1294 );
nand \U$22127 ( \22470 , \22468 , \22469 );
not \U$22128 ( \22471 , \22470 );
not \U$22129 ( \22472 , \15826 );
and \U$22130 ( \22473 , \22471 , \22472 );
and \U$22131 ( \22474 , \22470 , \15826 );
nor \U$22132 ( \22475 , \22473 , \22474 );
not \U$22133 ( \22476 , \22475 );
or \U$22134 ( \22477 , \22465 , \22476 );
or \U$22135 ( \22478 , \22475 , \22464 );
nand \U$22136 ( \22479 , \22477 , \22478 );
not \U$22137 ( \22480 , \21647 );
not \U$22138 ( \22481 , \21634 );
or \U$22139 ( \22482 , \22480 , \22481 );
nand \U$22140 ( \22483 , \22482 , \21620 );
not \U$22141 ( \22484 , \21634 );
nand \U$22142 ( \22485 , \22484 , \21646 );
nand \U$22143 ( \22486 , \22483 , \22485 );
xor \U$22144 ( \22487 , \22479 , \22486 );
not \U$22145 ( \22488 , \21604 );
not \U$22146 ( \22489 , \21591 );
or \U$22147 ( \22490 , \22488 , \22489 );
nand \U$22148 ( \22491 , \22490 , \21578 );
not \U$22149 ( \22492 , \21591 );
nand \U$22150 ( \22493 , \22492 , \21603 );
nand \U$22151 ( \22494 , \22491 , \22493 );
xor \U$22152 ( \22495 , \22487 , \22494 );
xor \U$22153 ( \22496 , \21777 , \21783 );
and \U$22154 ( \22497 , \22496 , \21788 );
and \U$22155 ( \22498 , \21777 , \21783 );
or \U$22156 ( \22499 , \22497 , \22498 );
xor \U$22157 ( \22500 , \22495 , \22499 );
not \U$22158 ( \22501 , \21747 );
not \U$22159 ( \22502 , \21742 );
or \U$22160 ( \22503 , \22501 , \22502 );
or \U$22161 ( \22504 , \21742 , \21747 );
nand \U$22162 ( \22505 , \22504 , \21733 );
nand \U$22163 ( \22506 , \22503 , \22505 );
xor \U$22164 ( \22507 , \22500 , \22506 );
xnor \U$22165 ( \22508 , \22459 , \22507 );
xor \U$22166 ( \22509 , \22419 , \22508 );
not \U$22167 ( \22510 , \21651 );
not \U$22168 ( \22511 , \21609 );
or \U$22169 ( \22512 , \22510 , \22511 );
not \U$22170 ( \22513 , \21608 );
not \U$22171 ( \22514 , \21648 );
or \U$22172 ( \22515 , \22513 , \22514 );
nand \U$22173 ( \22516 , \22515 , \21695 );
nand \U$22174 ( \22517 , \22512 , \22516 );
not \U$22175 ( \22518 , \1089 );
not \U$22176 ( \22519 , \22063 );
or \U$22177 ( \22520 , \22518 , \22519 );
nand \U$22178 ( \22521 , \15765 , \1147 );
nand \U$22179 ( \22522 , \22520 , \22521 );
not \U$22180 ( \22523 , \1376 );
not \U$22181 ( \22524 , \15476 );
or \U$22182 ( \22525 , \22523 , \22524 );
nand \U$22183 ( \22526 , \21669 , \1429 );
nand \U$22184 ( \22527 , \22525 , \22526 );
xor \U$22185 ( \22528 , \22522 , \22527 );
not \U$22186 ( \22529 , \1737 );
not \U$22187 ( \22530 , \15488 );
or \U$22188 ( \22531 , \22529 , \22530 );
nand \U$22189 ( \22532 , \21760 , \1702 );
nand \U$22190 ( \22533 , \22531 , \22532 );
xor \U$22191 ( \22534 , \22528 , \22533 );
xor \U$22192 ( \22535 , \21819 , \21829 );
and \U$22193 ( \22536 , \22535 , \21840 );
and \U$22194 ( \22537 , \21819 , \21829 );
or \U$22195 ( \22538 , \22536 , \22537 );
xor \U$22196 ( \22539 , \22534 , \22538 );
or \U$22197 ( \22540 , \21888 , \21909 );
nand \U$22198 ( \22541 , \22540 , \21898 );
nand \U$22199 ( \22542 , \21888 , \21909 );
nand \U$22200 ( \22543 , \22541 , \22542 );
xor \U$22201 ( \22544 , \22539 , \22543 );
xor \U$22202 ( \22545 , \22517 , \22544 );
not \U$22203 ( \22546 , \16674 );
not \U$22204 ( \22547 , \21951 );
or \U$22205 ( \22548 , \22546 , \22547 );
nand \U$22206 ( \22549 , \15738 , RIbb2dbd0_57);
nand \U$22207 ( \22550 , \22548 , \22549 );
not \U$22208 ( \22551 , \1570 );
not \U$22209 ( \22552 , RIbb2f250_9);
not \U$22210 ( \22553 , \11580 );
or \U$22211 ( \22554 , \22552 , \22553 );
not \U$22212 ( \22555 , \17440 );
nand \U$22213 ( \22556 , \22555 , \1566 );
nand \U$22214 ( \22557 , \22554 , \22556 );
not \U$22215 ( \22558 , \22557 );
or \U$22216 ( \22559 , \22551 , \22558 );
nand \U$22217 ( \22560 , \22075 , \1533 );
nand \U$22218 ( \22561 , \22559 , \22560 );
xor \U$22219 ( \22562 , \22550 , \22561 );
not \U$22220 ( \22563 , \1077 );
not \U$22221 ( \22564 , RIbb2f160_11);
not \U$22222 ( \22565 , \12249 );
or \U$22223 ( \22566 , \22564 , \22565 );
nand \U$22224 ( \22567 , \10764 , \1805 );
nand \U$22225 ( \22568 , \22566 , \22567 );
not \U$22226 ( \22569 , \22568 );
or \U$22227 ( \22570 , \22563 , \22569 );
nand \U$22228 ( \22571 , \21817 , \1011 );
nand \U$22229 ( \22572 , \22570 , \22571 );
xor \U$22230 ( \22573 , \22562 , \22572 );
xor \U$22231 ( \22574 , \21674 , \21683 );
and \U$22232 ( \22575 , \22574 , \21694 );
and \U$22233 ( \22576 , \21674 , \21683 );
or \U$22234 ( \22577 , \22575 , \22576 );
xor \U$22235 ( \22578 , \22573 , \22577 );
not \U$22236 ( \22579 , RIbb2f070_13);
not \U$22237 ( \22580 , \9841 );
not \U$22238 ( \22581 , \22580 );
or \U$22239 ( \22582 , \22579 , \22581 );
nand \U$22240 ( \22583 , \9841 , \906 );
nand \U$22241 ( \22584 , \22582 , \22583 );
and \U$22242 ( \22585 , \22584 , \998 );
not \U$22243 ( \22586 , \21644 );
nor \U$22244 ( \22587 , \22586 , \1654 );
nor \U$22245 ( \22588 , \22585 , \22587 );
not \U$22246 ( \22589 , \22588 );
not \U$22247 ( \22590 , \1445 );
not \U$22248 ( \22591 , \21626 );
or \U$22249 ( \22592 , \22590 , \22591 );
nand \U$22250 ( \22593 , \15790 , \1517 );
nand \U$22251 ( \22594 , \22592 , \22593 );
not \U$22252 ( \22595 , \22594 );
not \U$22253 ( \22596 , \832 );
not \U$22254 ( \22597 , \21616 );
or \U$22255 ( \22598 , \22596 , \22597 );
nand \U$22256 ( \22599 , \15778 , \836 );
nand \U$22257 ( \22600 , \22598 , \22599 );
not \U$22258 ( \22601 , \22600 );
not \U$22259 ( \22602 , \22601 );
or \U$22260 ( \22603 , \22595 , \22602 );
or \U$22261 ( \22604 , \22601 , \22594 );
nand \U$22262 ( \22605 , \22603 , \22604 );
not \U$22263 ( \22606 , \22605 );
or \U$22264 ( \22607 , \22589 , \22606 );
or \U$22265 ( \22608 , \22605 , \22588 );
nand \U$22266 ( \22609 , \22607 , \22608 );
xor \U$22267 ( \22610 , \22578 , \22609 );
xnor \U$22268 ( \22611 , \22545 , \22610 );
not \U$22269 ( \22612 , \22611 );
not \U$22270 ( \22613 , \21752 );
not \U$22271 ( \22614 , \22613 );
not \U$22272 ( \22615 , \21729 );
not \U$22273 ( \22616 , \22615 );
not \U$22274 ( \22617 , \22616 );
or \U$22275 ( \22618 , \22614 , \22617 );
not \U$22276 ( \22619 , \22615 );
not \U$22277 ( \22620 , \21752 );
or \U$22278 ( \22621 , \22619 , \22620 );
nand \U$22279 ( \22622 , \22621 , \21789 );
nand \U$22280 ( \22623 , \22618 , \22622 );
not \U$22281 ( \22624 , \22623 );
nand \U$22282 ( \22625 , \22612 , \22624 );
nand \U$22283 ( \22626 , \22611 , \22623 );
nand \U$22284 ( \22627 , \22625 , \22626 );
xor \U$22285 ( \22628 , \21562 , \21566 );
and \U$22286 ( \22629 , \22628 , \21697 );
and \U$22287 ( \22630 , \21562 , \21566 );
or \U$22288 ( \22631 , \22629 , \22630 );
not \U$22289 ( \22632 , \22631 );
and \U$22290 ( \22633 , \22627 , \22632 );
not \U$22291 ( \22634 , \22627 );
and \U$22292 ( \22635 , \22634 , \22631 );
nor \U$22293 ( \22636 , \22633 , \22635 );
xor \U$22294 ( \22637 , \22509 , \22636 );
not \U$22295 ( \22638 , \22637 );
not \U$22296 ( \22639 , \22638 );
or \U$22297 ( \22640 , \22412 , \22639 );
nand \U$22298 ( \22641 , \22637 , \22410 );
nand \U$22299 ( \22642 , \22640 , \22641 );
not \U$22300 ( \22643 , \22642 );
or \U$22301 ( \22644 , \22406 , \22643 );
or \U$22302 ( \22645 , \22642 , \22405 );
nand \U$22303 ( \22646 , \22644 , \22645 );
xor \U$22304 ( \22647 , \22133 , \22646 );
xor \U$22305 ( \22648 , \21991 , \21995 );
and \U$22306 ( \22649 , \22648 , \22122 );
and \U$22307 ( \22650 , \21991 , \21995 );
or \U$22308 ( \22651 , \22649 , \22650 );
nor \U$22309 ( \22652 , \22647 , \22651 );
nor \U$22310 ( \22653 , \20631 , \21549 , \22124 , \22652 );
not \U$22311 ( \22654 , \22653 );
xor \U$22312 ( \22655 , \21540 , \21537 );
xnor \U$22313 ( \22656 , \22655 , \20635 );
xor \U$22314 ( \22657 , \20485 , \20612 );
xor \U$22315 ( \22658 , \22657 , \20615 );
not \U$22316 ( \22659 , \22658 );
xor \U$22317 ( \22660 , \21137 , \21148 );
xor \U$22318 ( \22661 , \22660 , \21534 );
not \U$22319 ( \22662 , \22661 );
nand \U$22320 ( \22663 , \22659 , \22662 );
xor \U$22321 ( \22664 , \20600 , \20505 );
xor \U$22322 ( \22665 , \22664 , \20495 );
not \U$22323 ( \22666 , \22665 );
xor \U$22324 ( \22667 , \20830 , \20638 );
xor \U$22325 ( \22668 , \22667 , \20989 );
not \U$22326 ( \22669 , \22668 );
or \U$22327 ( \22670 , \22666 , \22669 );
xor \U$22328 ( \22671 , \20802 , \20808 );
xor \U$22329 ( \22672 , \22671 , \20818 );
not \U$22330 ( \22673 , \22672 );
and \U$22331 ( \22674 , \20864 , \20844 );
not \U$22332 ( \22675 , \20864 );
and \U$22333 ( \22676 , \22675 , \20856 );
nor \U$22334 ( \22677 , \22674 , \22676 );
xnor \U$22335 ( \22678 , \22677 , \20851 );
not \U$22336 ( \22679 , \22678 );
not \U$22337 ( \22680 , \22679 );
or \U$22338 ( \22681 , \22673 , \22680 );
or \U$22339 ( \22682 , \22679 , \22672 );
not \U$22340 ( \22683 , \12690 );
not \U$22341 ( \22684 , \1419 );
and \U$22342 ( \22685 , RIbb2dea0_51, \22684 );
not \U$22343 ( \22686 , RIbb2dea0_51);
and \U$22344 ( \22687 , \22686 , \1419 );
or \U$22345 ( \22688 , \22685 , \22687 );
not \U$22346 ( \22689 , \22688 );
or \U$22347 ( \22690 , \22683 , \22689 );
nand \U$22348 ( \22691 , \20804 , \12692 );
nand \U$22349 ( \22692 , \22690 , \22691 );
not \U$22350 ( \22693 , \22692 );
and \U$22351 ( \22694 , RIbb2dae0_59, \1729 );
not \U$22352 ( \22695 , RIbb2dae0_59);
and \U$22353 ( \22696 , \22695 , \3478 );
or \U$22354 ( \22697 , \22694 , \22696 );
and \U$22355 ( \22698 , \22697 , \16271 );
and \U$22356 ( \22699 , \20847 , \16257 );
nor \U$22357 ( \22700 , \22698 , \22699 );
nand \U$22358 ( \22701 , \22693 , \22700 );
not \U$22359 ( \22702 , \22701 );
not \U$22360 ( \22703 , \1570 );
not \U$22361 ( \22704 , \20729 );
or \U$22362 ( \22705 , \22703 , \22704 );
and \U$22363 ( \22706 , \16553 , \5064 );
not \U$22364 ( \22707 , \16553 );
and \U$22365 ( \22708 , \22707 , RIbb2f250_9);
or \U$22366 ( \22709 , \22706 , \22708 );
nand \U$22367 ( \22710 , \22709 , \1533 );
nand \U$22368 ( \22711 , \22705 , \22710 );
nor \U$22369 ( \22712 , \19063 , \1084 );
not \U$22370 ( \22713 , \1737 );
not \U$22371 ( \22714 , \21263 );
or \U$22372 ( \22715 , \22713 , \22714 );
not \U$22373 ( \22716 , RIbb2f340_7);
not \U$22374 ( \22717 , \20552 );
or \U$22375 ( \22718 , \22716 , \22717 );
nand \U$22376 ( \22719 , \17517 , \2700 );
nand \U$22377 ( \22720 , \22718 , \22719 );
nand \U$22378 ( \22721 , \22720 , \1701 );
nand \U$22379 ( \22722 , \22715 , \22721 );
xor \U$22380 ( \22723 , \22712 , \22722 );
not \U$22381 ( \22724 , \1533 );
not \U$22382 ( \22725 , RIbb2f250_9);
not \U$22383 ( \22726 , \17755 );
or \U$22384 ( \22727 , \22725 , \22726 );
nand \U$22385 ( \22728 , \16703 , \1524 );
nand \U$22386 ( \22729 , \22727 , \22728 );
not \U$22387 ( \22730 , \22729 );
or \U$22388 ( \22731 , \22724 , \22730 );
nand \U$22389 ( \22732 , \22709 , \1569 );
nand \U$22390 ( \22733 , \22731 , \22732 );
and \U$22391 ( \22734 , \22723 , \22733 );
and \U$22392 ( \22735 , \22712 , \22722 );
or \U$22393 ( \22736 , \22734 , \22735 );
xor \U$22394 ( \22737 , \22711 , \22736 );
not \U$22395 ( \22738 , \836 );
not \U$22396 ( \22739 , \21086 );
or \U$22397 ( \22740 , \22738 , \22739 );
not \U$22398 ( \22741 , RIbb2ee90_17);
not \U$22399 ( \22742 , \18552 );
or \U$22400 ( \22743 , \22741 , \22742 );
nand \U$22401 ( \22744 , \13545 , \3699 );
nand \U$22402 ( \22745 , \22743 , \22744 );
nand \U$22403 ( \22746 , \22745 , \831 );
nand \U$22404 ( \22747 , \22740 , \22746 );
and \U$22405 ( \22748 , \22737 , \22747 );
and \U$22406 ( \22749 , \22711 , \22736 );
or \U$22407 ( \22750 , \22748 , \22749 );
not \U$22408 ( \22751 , \22750 );
or \U$22409 ( \22752 , \22702 , \22751 );
not \U$22410 ( \22753 , \16271 );
not \U$22411 ( \22754 , \22697 );
or \U$22412 ( \22755 , \22753 , \22754 );
nand \U$22413 ( \22756 , \20847 , \16257 );
nand \U$22414 ( \22757 , \22755 , \22756 );
nand \U$22415 ( \22758 , \22757 , \22692 );
nand \U$22416 ( \22759 , \22752 , \22758 );
nand \U$22417 ( \22760 , \22682 , \22759 );
nand \U$22418 ( \22761 , \22681 , \22760 );
not \U$22419 ( \22762 , \22761 );
not \U$22420 ( \22763 , \20870 );
not \U$22421 ( \22764 , \20874 );
or \U$22422 ( \22765 , \22763 , \22764 );
nand \U$22423 ( \22766 , \20866 , \20869 );
nand \U$22424 ( \22767 , \22765 , \22766 );
not \U$22425 ( \22768 , \20878 );
and \U$22426 ( \22769 , \22767 , \22768 );
not \U$22427 ( \22770 , \22767 );
and \U$22428 ( \22771 , \22770 , \20878 );
nor \U$22429 ( \22772 , \22769 , \22771 );
not \U$22430 ( \22773 , \22772 );
not \U$22431 ( \22774 , \22773 );
or \U$22432 ( \22775 , \22762 , \22774 );
not \U$22433 ( \22776 , \22761 );
not \U$22434 ( \22777 , \22776 );
not \U$22435 ( \22778 , \22772 );
or \U$22436 ( \22779 , \22777 , \22778 );
xor \U$22437 ( \22780 , \20920 , \20947 );
xor \U$22438 ( \22781 , \22780 , \20983 );
nand \U$22439 ( \22782 , \22779 , \22781 );
nand \U$22440 ( \22783 , \22775 , \22782 );
not \U$22441 ( \22784 , \22783 );
xor \U$22442 ( \22785 , \20786 , \20788 );
xor \U$22443 ( \22786 , \22785 , \20827 );
not \U$22444 ( \22787 , \22786 );
or \U$22445 ( \22788 , \22784 , \22787 );
or \U$22446 ( \22789 , \22783 , \22786 );
xor \U$22447 ( \22790 , \20880 , \20886 );
xor \U$22448 ( \22791 , \22790 , \20986 );
nand \U$22449 ( \22792 , \22789 , \22791 );
nand \U$22450 ( \22793 , \22788 , \22792 );
nand \U$22451 ( \22794 , \22670 , \22793 );
not \U$22452 ( \22795 , \22665 );
not \U$22453 ( \22796 , \22668 );
nand \U$22454 ( \22797 , \22795 , \22796 );
nand \U$22455 ( \22798 , \22794 , \22797 );
xor \U$22456 ( \22799 , \20992 , \21131 );
xor \U$22457 ( \22800 , \22799 , \21134 );
xor \U$22458 ( \22801 , \22798 , \22800 );
xor \U$22459 ( \22802 , \20979 , \20969 );
xnor \U$22460 ( \22803 , \22802 , \20959 );
not \U$22461 ( \22804 , \22803 );
not \U$22462 ( \22805 , \22804 );
xor \U$22463 ( \22806 , \20897 , \20907 );
xor \U$22464 ( \22807 , \22806 , \20917 );
not \U$22465 ( \22808 , \22807 );
or \U$22466 ( \22809 , \22805 , \22808 );
not \U$22467 ( \22810 , \22803 );
not \U$22468 ( \22811 , \22807 );
not \U$22469 ( \22812 , \22811 );
or \U$22470 ( \22813 , \22810 , \22812 );
xor \U$22471 ( \22814 , \20922 , \20932 );
xor \U$22472 ( \22815 , \22814 , \20944 );
nand \U$22473 ( \22816 , \22813 , \22815 );
nand \U$22474 ( \22817 , \22809 , \22816 );
not \U$22475 ( \22818 , \22817 );
and \U$22476 ( \22819 , \21017 , \21009 );
not \U$22477 ( \22820 , \21017 );
and \U$22478 ( \22821 , \22820 , \21010 );
or \U$22479 ( \22822 , \22819 , \22821 );
xor \U$22480 ( \22823 , \20998 , \22822 );
not \U$22481 ( \22824 , \22823 );
or \U$22482 ( \22825 , \22818 , \22824 );
or \U$22483 ( \22826 , \22817 , \22823 );
xor \U$22484 ( \22827 , \20791 , \20821 );
xor \U$22485 ( \22828 , \22827 , \20824 );
nand \U$22486 ( \22829 , \22826 , \22828 );
nand \U$22487 ( \22830 , \22825 , \22829 );
not \U$22488 ( \22831 , \22830 );
xor \U$22489 ( \22832 , \21019 , \21031 );
xnor \U$22490 ( \22833 , \22832 , \21038 );
not \U$22491 ( \22834 , \22833 );
or \U$22492 ( \22835 , \22831 , \22834 );
or \U$22493 ( \22836 , \22830 , \22833 );
xor \U$22494 ( \22837 , \21127 , \21054 );
xnor \U$22495 ( \22838 , \22837 , \21057 );
nand \U$22496 ( \22839 , \22836 , \22838 );
nand \U$22497 ( \22840 , \22835 , \22839 );
xor \U$22498 ( \22841 , \21040 , \21129 );
and \U$22499 ( \22842 , \22841 , \20994 );
not \U$22500 ( \22843 , \22841 );
not \U$22501 ( \22844 , \20994 );
and \U$22502 ( \22845 , \22843 , \22844 );
nor \U$22503 ( \22846 , \22842 , \22845 );
or \U$22504 ( \22847 , \22840 , \22846 );
not \U$22505 ( \22848 , \21152 );
not \U$22506 ( \22849 , \21155 );
not \U$22507 ( \22850 , \22849 );
or \U$22508 ( \22851 , \22848 , \22850 );
nand \U$22509 ( \22852 , \21151 , \21155 );
nand \U$22510 ( \22853 , \22851 , \22852 );
and \U$22511 ( \22854 , \22853 , \21510 );
not \U$22512 ( \22855 , \22853 );
not \U$22513 ( \22856 , \21510 );
and \U$22514 ( \22857 , \22855 , \22856 );
nor \U$22515 ( \22858 , \22854 , \22857 );
nand \U$22516 ( \22859 , \22847 , \22858 );
nand \U$22517 ( \22860 , \22846 , \22840 );
nand \U$22518 ( \22861 , \22859 , \22860 );
and \U$22519 ( \22862 , \22801 , \22861 );
and \U$22520 ( \22863 , \22798 , \22800 );
or \U$22521 ( \22864 , \22862 , \22863 );
buf \U$22522 ( \22865 , \22864 );
and \U$22523 ( \22866 , \22663 , \22865 );
not \U$22524 ( \22867 , \22658 );
nor \U$22525 ( \22868 , \22867 , \22662 );
nor \U$22526 ( \22869 , \22866 , \22868 );
nand \U$22527 ( \22870 , \22656 , \22869 );
not \U$22528 ( \22871 , \22870 );
xor \U$22529 ( \22872 , \22846 , \22840 );
not \U$22530 ( \22873 , \22858 );
and \U$22531 ( \22874 , \22872 , \22873 );
not \U$22532 ( \22875 , \22872 );
and \U$22533 ( \22876 , \22875 , \22858 );
nor \U$22534 ( \22877 , \22874 , \22876 );
buf \U$22535 ( \22878 , \22877 );
not \U$22536 ( \22879 , \22878 );
xor \U$22537 ( \22880 , \21358 , \21370 );
xor \U$22538 ( \22881 , \22880 , \21382 );
not \U$22539 ( \22882 , \22881 );
not \U$22540 ( \22883 , \22882 );
xor \U$22541 ( \22884 , \21189 , \21199 );
xor \U$22542 ( \22885 , \22884 , \21209 );
not \U$22543 ( \22886 , \22885 );
or \U$22544 ( \22887 , \22883 , \22886 );
not \U$22545 ( \22888 , \22885 );
not \U$22546 ( \22889 , \22888 );
not \U$22547 ( \22890 , \22881 );
or \U$22548 ( \22891 , \22889 , \22890 );
not \U$22549 ( \22892 , \8362 );
not \U$22550 ( \22893 , RIbb2e350_41);
not \U$22551 ( \22894 , \19676 );
not \U$22552 ( \22895 , \22894 );
or \U$22553 ( \22896 , \22893 , \22895 );
nand \U$22554 ( \22897 , \3022 , \7097 );
nand \U$22555 ( \22898 , \22896 , \22897 );
not \U$22556 ( \22899 , \22898 );
or \U$22557 ( \22900 , \22892 , \22899 );
nand \U$22558 ( \22901 , \21494 , \8353 );
nand \U$22559 ( \22902 , \22900 , \22901 );
not \U$22560 ( \22903 , \14930 );
not \U$22561 ( \22904 , \21482 );
or \U$22562 ( \22905 , \22903 , \22904 );
not \U$22563 ( \22906 , RIbb2ddb0_53);
not \U$22564 ( \22907 , \4339 );
or \U$22565 ( \22908 , \22906 , \22907 );
nand \U$22566 ( \22909 , \4340 , \13463 );
nand \U$22567 ( \22910 , \22908 , \22909 );
nand \U$22568 ( \22911 , \22910 , \14920 );
nand \U$22569 ( \22912 , \22905 , \22911 );
xor \U$22570 ( \22913 , \22902 , \22912 );
not \U$22571 ( \22914 , \7104 );
not \U$22572 ( \22915 , \21332 );
or \U$22573 ( \22916 , \22914 , \22915 );
and \U$22574 ( \22917 , RIbb2e440_39, \13731 );
not \U$22575 ( \22918 , RIbb2e440_39);
and \U$22576 ( \22919 , \22918 , \3274 );
or \U$22577 ( \22920 , \22917 , \22919 );
nand \U$22578 ( \22921 , \22920 , \7103 );
nand \U$22579 ( \22922 , \22916 , \22921 );
and \U$22580 ( \22923 , \22913 , \22922 );
and \U$22581 ( \22924 , \22902 , \22912 );
or \U$22582 ( \22925 , \22923 , \22924 );
nand \U$22583 ( \22926 , \22891 , \22925 );
nand \U$22584 ( \22927 , \22887 , \22926 );
not \U$22585 ( \22928 , \22927 );
not \U$22586 ( \22929 , \9098 );
not \U$22587 ( \22930 , RIbb2e260_43);
not \U$22588 ( \22931 , \13835 );
or \U$22589 ( \22932 , \22930 , \22931 );
not \U$22590 ( \22933 , RIbb2e260_43);
nand \U$22591 ( \22934 , \22933 , \13903 );
nand \U$22592 ( \22935 , \22932 , \22934 );
not \U$22593 ( \22936 , \22935 );
or \U$22594 ( \22937 , \22929 , \22936 );
nand \U$22595 ( \22938 , \21406 , \9099 );
nand \U$22596 ( \22939 , \22937 , \22938 );
not \U$22597 ( \22940 , RIbb2d888_64);
not \U$22598 ( \22941 , \21473 );
or \U$22599 ( \22942 , \22940 , \22941 );
not \U$22600 ( \22943 , RIbb2d900_63);
not \U$22601 ( \22944 , \1069 );
or \U$22602 ( \22945 , \22943 , \22944 );
not \U$22603 ( \22946 , RIbb2d900_63);
nand \U$22604 ( \22947 , \16277 , \22946 );
nand \U$22605 ( \22948 , \22945 , \22947 );
nand \U$22606 ( \22949 , \22948 , \17275 );
nand \U$22607 ( \22950 , \22942 , \22949 );
nor \U$22608 ( \22951 , \22939 , \22950 );
buf \U$22609 ( \22952 , \14613 );
not \U$22610 ( \22953 , \22952 );
and \U$22611 ( \22954 , RIbb2dcc0_55, \15582 );
not \U$22612 ( \22955 , RIbb2dcc0_55);
and \U$22613 ( \22956 , \22955 , \1282 );
or \U$22614 ( \22957 , \22954 , \22956 );
not \U$22615 ( \22958 , \22957 );
or \U$22616 ( \22959 , \22953 , \22958 );
nand \U$22617 ( \22960 , \21425 , \15182 );
nand \U$22618 ( \22961 , \22959 , \22960 );
not \U$22619 ( \22962 , \22961 );
or \U$22620 ( \22963 , \22951 , \22962 );
nand \U$22621 ( \22964 , \22939 , \22950 );
nand \U$22622 ( \22965 , \22963 , \22964 );
not \U$22623 ( \22966 , \16674 );
not \U$22624 ( \22967 , RIbb2dbd0_57);
not \U$22625 ( \22968 , \7423 );
or \U$22626 ( \22969 , \22967 , \22968 );
nand \U$22627 ( \22970 , \3053 , \15741 );
nand \U$22628 ( \22971 , \22969 , \22970 );
not \U$22629 ( \22972 , \22971 );
or \U$22630 ( \22973 , \22966 , \22972 );
nand \U$22631 ( \22974 , \21438 , \15738 );
nand \U$22632 ( \22975 , \22973 , \22974 );
not \U$22633 ( \22976 , \10117 );
not \U$22634 ( \22977 , RIbb2e170_45);
buf \U$22635 ( \22978 , \17568 );
not \U$22636 ( \22979 , \22978 );
or \U$22637 ( \22980 , \22977 , \22979 );
nand \U$22638 ( \22981 , \3146 , \11065 );
nand \U$22639 ( \22982 , \22980 , \22981 );
not \U$22640 ( \22983 , \22982 );
or \U$22641 ( \22984 , \22976 , \22983 );
nand \U$22642 ( \22985 , \21417 , \10119 );
nand \U$22643 ( \22986 , \22984 , \22985 );
xor \U$22644 ( \22987 , \22975 , \22986 );
not \U$22645 ( \22988 , \11176 );
not \U$22646 ( \22989 , RIbb2e080_47);
not \U$22647 ( \22990 , \3520 );
or \U$22648 ( \22991 , \22989 , \22990 );
nand \U$22649 ( \22992 , \12096 , \10113 );
nand \U$22650 ( \22993 , \22991 , \22992 );
not \U$22651 ( \22994 , \22993 );
or \U$22652 ( \22995 , \22988 , \22994 );
nand \U$22653 ( \22996 , \12965 , \21460 );
nand \U$22654 ( \22997 , \22995 , \22996 );
and \U$22655 ( \22998 , \22987 , \22997 );
and \U$22656 ( \22999 , \22975 , \22986 );
or \U$22657 ( \23000 , \22998 , \22999 );
xor \U$22658 ( \23001 , \22965 , \23000 );
not \U$22659 ( \23002 , \12774 );
and \U$22660 ( \23003 , RIbb2dea0_51, \17207 );
not \U$22661 ( \23004 , RIbb2dea0_51);
and \U$22662 ( \23005 , \23004 , \1338 );
or \U$22663 ( \23006 , \23003 , \23005 );
not \U$22664 ( \23007 , \23006 );
or \U$22665 ( \23008 , \23002 , \23007 );
nand \U$22666 ( \23009 , \22688 , \12692 );
nand \U$22667 ( \23010 , \23008 , \23009 );
not \U$22668 ( \23011 , \6242 );
not \U$22669 ( \23012 , \21322 );
or \U$22670 ( \23013 , \23011 , \23012 );
not \U$22671 ( \23014 , RIbb2e530_37);
not \U$22672 ( \23015 , \19429 );
or \U$22673 ( \23016 , \23014 , \23015 );
nand \U$22674 ( \23017 , \4324 , \8701 );
nand \U$22675 ( \23018 , \23016 , \23017 );
nand \U$22676 ( \23019 , \23018 , \6251 );
nand \U$22677 ( \23020 , \23013 , \23019 );
xor \U$22678 ( \23021 , \23010 , \23020 );
not \U$22679 ( \23022 , \16271 );
and \U$22680 ( \23023 , RIbb2dae0_59, \3370 );
not \U$22681 ( \23024 , RIbb2dae0_59);
and \U$22682 ( \23025 , \23024 , \3363 );
or \U$22683 ( \23026 , \23023 , \23025 );
not \U$22684 ( \23027 , \23026 );
or \U$22685 ( \23028 , \23022 , \23027 );
nand \U$22686 ( \23029 , \22697 , \16257 );
nand \U$22687 ( \23030 , \23028 , \23029 );
and \U$22688 ( \23031 , \23021 , \23030 );
and \U$22689 ( \23032 , \23010 , \23020 );
or \U$22690 ( \23033 , \23031 , \23032 );
and \U$22691 ( \23034 , \23001 , \23033 );
and \U$22692 ( \23035 , \22965 , \23000 );
or \U$22693 ( \23036 , \23034 , \23035 );
not \U$22694 ( \23037 , \23036 );
or \U$22695 ( \23038 , \22928 , \23037 );
or \U$22696 ( \23039 , \22927 , \23036 );
and \U$22697 ( \23040 , \21212 , \21247 );
not \U$22698 ( \23041 , \21212 );
and \U$22699 ( \23042 , \23041 , \21248 );
nor \U$22700 ( \23043 , \23040 , \23042 );
not \U$22701 ( \23044 , \21304 );
and \U$22702 ( \23045 , \23043 , \23044 );
not \U$22703 ( \23046 , \23043 );
and \U$22704 ( \23047 , \23046 , \21304 );
nor \U$22705 ( \23048 , \23045 , \23047 );
not \U$22706 ( \23049 , \23048 );
nand \U$22707 ( \23050 , \23039 , \23049 );
nand \U$22708 ( \23051 , \23038 , \23050 );
not \U$22709 ( \23052 , \23051 );
xor \U$22710 ( \23053 , \21311 , \21313 );
xor \U$22711 ( \23054 , \23053 , \21339 );
not \U$22712 ( \23055 , \23054 );
not \U$22713 ( \23056 , \23055 );
not \U$22714 ( \23057 , \23056 );
not \U$22715 ( \23058 , \21387 );
not \U$22716 ( \23059 , \21348 );
not \U$22717 ( \23060 , \23059 );
or \U$22718 ( \23061 , \23058 , \23060 );
nand \U$22719 ( \23062 , \21386 , \21348 );
nand \U$22720 ( \23063 , \23061 , \23062 );
and \U$22721 ( \23064 , \23063 , \21391 );
not \U$22722 ( \23065 , \23063 );
and \U$22723 ( \23066 , \23065 , \21392 );
nor \U$22724 ( \23067 , \23064 , \23066 );
not \U$22725 ( \23068 , \23067 );
not \U$22726 ( \23069 , \23068 );
or \U$22727 ( \23070 , \23057 , \23069 );
or \U$22728 ( \23071 , \23056 , \23068 );
xor \U$22729 ( \23072 , \21477 , \21486 );
xor \U$22730 ( \23073 , \23072 , \21498 );
xor \U$22731 ( \23074 , \21316 , \21326 );
xor \U$22732 ( \23075 , \23074 , \21336 );
xor \U$22733 ( \23076 , \23073 , \23075 );
xor \U$22734 ( \23077 , \21442 , \21453 );
xor \U$22735 ( \23078 , \23077 , \21464 );
and \U$22736 ( \23079 , \23076 , \23078 );
and \U$22737 ( \23080 , \23073 , \23075 );
or \U$22738 ( \23081 , \23079 , \23080 );
nand \U$22739 ( \23082 , \23071 , \23081 );
nand \U$22740 ( \23083 , \23070 , \23082 );
not \U$22741 ( \23084 , \23083 );
or \U$22742 ( \23085 , \23052 , \23084 );
or \U$22743 ( \23086 , \23083 , \23051 );
xor \U$22744 ( \23087 , \21396 , \21399 );
xor \U$22745 ( \23088 , \23087 , \21504 );
nand \U$22746 ( \23089 , \23086 , \23088 );
nand \U$22747 ( \23090 , \23085 , \23089 );
xor \U$22748 ( \23091 , \21065 , \21105 );
xor \U$22749 ( \23092 , \23091 , \21124 );
xor \U$22750 ( \23093 , \21067 , \21091 );
xor \U$22751 ( \23094 , \23093 , \21102 );
not \U$22752 ( \23095 , \998 );
not \U$22753 ( \23096 , \21221 );
or \U$22754 ( \23097 , \23095 , \23096 );
buf \U$22755 ( \23098 , \15752 );
and \U$22756 ( \23099 , RIbb2f070_13, \23098 );
not \U$22757 ( \23100 , RIbb2f070_13);
and \U$22758 ( \23101 , \23100 , \16567 );
nor \U$22759 ( \23102 , \23099 , \23101 );
nand \U$22760 ( \23103 , \23102 , \915 );
nand \U$22761 ( \23104 , \23097 , \23103 );
not \U$22762 ( \23105 , \1444 );
and \U$22763 ( \23106 , RIbb2ef80_15, \18353 );
not \U$22764 ( \23107 , RIbb2ef80_15);
and \U$22765 ( \23108 , \23107 , \14526 );
or \U$22766 ( \23109 , \23106 , \23108 );
not \U$22767 ( \23110 , \23109 );
or \U$22768 ( \23111 , \23105 , \23110 );
nand \U$22769 ( \23112 , \21074 , \1517 );
nand \U$22770 ( \23113 , \23111 , \23112 );
xor \U$22771 ( \23114 , \23104 , \23113 );
not \U$22772 ( \23115 , \853 );
not \U$22773 ( \23116 , RIbb2eda0_19);
not \U$22774 ( \23117 , \13809 );
or \U$22775 ( \23118 , \23116 , \23117 );
nand \U$22776 ( \23119 , \12347 , \3251 );
nand \U$22777 ( \23120 , \23118 , \23119 );
not \U$22778 ( \23121 , \23120 );
or \U$22779 ( \23122 , \23115 , \23121 );
nand \U$22780 ( \23123 , \21231 , \854 );
nand \U$22781 ( \23124 , \23122 , \23123 );
and \U$22782 ( \23125 , \23114 , \23124 );
and \U$22783 ( \23126 , \23104 , \23113 );
or \U$22784 ( \23127 , \23125 , \23126 );
not \U$22785 ( \23128 , \23127 );
not \U$22786 ( \23129 , \3886 );
not \U$22787 ( \23130 , RIbb2e710_33);
not \U$22788 ( \23131 , \18564 );
or \U$22789 ( \23132 , \23130 , \23131 );
nand \U$22790 ( \23133 , \5954 , \2935 );
nand \U$22791 ( \23134 , \23132 , \23133 );
not \U$22792 ( \23135 , \23134 );
or \U$22793 ( \23136 , \23129 , \23135 );
nand \U$22794 ( \23137 , \21185 , \4791 );
nand \U$22795 ( \23138 , \23136 , \23137 );
not \U$22796 ( \23139 , \2925 );
not \U$22797 ( \23140 , \21297 );
or \U$22798 ( \23141 , \23139 , \23140 );
not \U$22799 ( \23142 , RIbb2e8f0_29);
not \U$22800 ( \23143 , \8319 );
or \U$22801 ( \23144 , \23142 , \23143 );
nand \U$22802 ( \23145 , \8318 , \2949 );
nand \U$22803 ( \23146 , \23144 , \23145 );
nand \U$22804 ( \23147 , \23146 , \2922 );
nand \U$22805 ( \23148 , \23141 , \23147 );
xor \U$22806 ( \23149 , \23138 , \23148 );
not \U$22807 ( \23150 , \3445 );
not \U$22808 ( \23151 , RIbb2e9e0_27);
not \U$22809 ( \23152 , \13919 );
or \U$22810 ( \23153 , \23151 , \23152 );
nand \U$22811 ( \23154 , \9278 , \11284 );
nand \U$22812 ( \23155 , \23153 , \23154 );
not \U$22813 ( \23156 , \23155 );
or \U$22814 ( \23157 , \23150 , \23156 );
nand \U$22815 ( \23158 , \21205 , \3465 );
nand \U$22816 ( \23159 , \23157 , \23158 );
and \U$22817 ( \23160 , \23149 , \23159 );
and \U$22818 ( \23161 , \23138 , \23148 );
or \U$22819 ( \23162 , \23160 , \23161 );
not \U$22820 ( \23163 , \23162 );
or \U$22821 ( \23164 , \23128 , \23163 );
or \U$22822 ( \23165 , \23162 , \23127 );
or \U$22823 ( \23166 , RIbb2f2c8_8, RIbb2f250_9);
nand \U$22824 ( \23167 , \23166 , \19064 );
and \U$22825 ( \23168 , RIbb2f2c8_8, RIbb2f250_9);
nor \U$22826 ( \23169 , \23168 , \1734 );
and \U$22827 ( \23170 , \23167 , \23169 );
not \U$22828 ( \23171 , \1737 );
not \U$22829 ( \23172 , \22720 );
or \U$22830 ( \23173 , \23171 , \23172 );
and \U$22831 ( \23174 , RIbb2f340_7, \17506 );
not \U$22832 ( \23175 , RIbb2f340_7);
and \U$22833 ( \23176 , \23175 , \19063 );
nor \U$22834 ( \23177 , \23174 , \23176 );
nand \U$22835 ( \23178 , \23177 , \1701 );
nand \U$22836 ( \23179 , \23173 , \23178 );
and \U$22837 ( \23180 , \23170 , \23179 );
not \U$22838 ( \23181 , \1077 );
not \U$22839 ( \23182 , \21272 );
or \U$22840 ( \23183 , \23181 , \23182 );
not \U$22841 ( \23184 , RIbb2f160_11);
not \U$22842 ( \23185 , \19831 );
not \U$22843 ( \23186 , \23185 );
or \U$22844 ( \23187 , \23184 , \23186 );
nand \U$22845 ( \23188 , \19831 , \1805 );
nand \U$22846 ( \23189 , \23187 , \23188 );
nand \U$22847 ( \23190 , \23189 , \1011 );
nand \U$22848 ( \23191 , \23183 , \23190 );
xor \U$22849 ( \23192 , \23180 , \23191 );
not \U$22850 ( \23193 , \998 );
not \U$22851 ( \23194 , \23102 );
or \U$22852 ( \23195 , \23193 , \23194 );
not \U$22853 ( \23196 , RIbb2f070_13);
not \U$22854 ( \23197 , \16575 );
not \U$22855 ( \23198 , \23197 );
or \U$22856 ( \23199 , \23196 , \23198 );
nand \U$22857 ( \23200 , \16575 , \1656 );
nand \U$22858 ( \23201 , \23199 , \23200 );
nand \U$22859 ( \23202 , \23201 , \915 );
nand \U$22860 ( \23203 , \23195 , \23202 );
and \U$22861 ( \23204 , \23192 , \23203 );
and \U$22862 ( \23205 , \23180 , \23191 );
or \U$22863 ( \23206 , \23204 , \23205 );
not \U$22864 ( \23207 , \2941 );
not \U$22865 ( \23208 , \21285 );
or \U$22866 ( \23209 , \23207 , \23208 );
not \U$22867 ( \23210 , RIbb2e800_31);
not \U$22868 ( \23211 , \19868 );
or \U$22869 ( \23212 , \23210 , \23211 );
nand \U$22870 ( \23213 , \6937 , \9169 );
nand \U$22871 ( \23214 , \23212 , \23213 );
nand \U$22872 ( \23215 , \23214 , \2939 );
nand \U$22873 ( \23216 , \23209 , \23215 );
xor \U$22874 ( \23217 , \23206 , \23216 );
not \U$22875 ( \23218 , \4712 );
not \U$22876 ( \23219 , RIbb2e620_35);
not \U$22877 ( \23220 , \6197 );
or \U$22878 ( \23221 , \23219 , \23220 );
nand \U$22879 ( \23222 , \9020 , \6688 );
nand \U$22880 ( \23223 , \23221 , \23222 );
not \U$22881 ( \23224 , \23223 );
or \U$22882 ( \23225 , \23218 , \23224 );
nand \U$22883 ( \23226 , \21242 , \5845 );
nand \U$22884 ( \23227 , \23225 , \23226 );
and \U$22885 ( \23228 , \23217 , \23227 );
and \U$22886 ( \23229 , \23206 , \23216 );
or \U$22887 ( \23230 , \23228 , \23229 );
nand \U$22888 ( \23231 , \23165 , \23230 );
nand \U$22889 ( \23232 , \23164 , \23231 );
xor \U$22890 ( \23233 , \23094 , \23232 );
xor \U$22891 ( \23234 , \21069 , \21078 );
xor \U$22892 ( \23235 , \23234 , \21088 );
xor \U$22893 ( \23236 , \21223 , \21233 );
xor \U$22894 ( \23237 , \23236 , \21244 );
xor \U$22895 ( \23238 , \23235 , \23237 );
not \U$22896 ( \23239 , \2078 );
not \U$22897 ( \23240 , \21354 );
or \U$22898 ( \23241 , \23239 , \23240 );
not \U$22899 ( \23242 , RIbb2ecb0_21);
not \U$22900 ( \23243 , \12174 );
not \U$22901 ( \23244 , \23243 );
or \U$22902 ( \23245 , \23242 , \23244 );
nand \U$22903 ( \23246 , \12174 , \5481 );
nand \U$22904 ( \23247 , \23245 , \23246 );
nand \U$22905 ( \23248 , \2077 , \23247 );
nand \U$22906 ( \23249 , \23241 , \23248 );
not \U$22907 ( \23250 , \3382 );
not \U$22908 ( \23251 , \21195 );
or \U$22909 ( \23252 , \23250 , \23251 );
not \U$22910 ( \23253 , RIbb2ebc0_23);
not \U$22911 ( \23254 , \11143 );
or \U$22912 ( \23255 , \23253 , \23254 );
nand \U$22913 ( \23256 , \11142 , \3401 );
nand \U$22914 ( \23257 , \23255 , \23256 );
nand \U$22915 ( \23258 , \23257 , \3406 );
nand \U$22916 ( \23259 , \23252 , \23258 );
xor \U$22917 ( \23260 , \23249 , \23259 );
not \U$22918 ( \23261 , \2980 );
and \U$22919 ( \23262 , RIbb2ead0_25, \12233 );
not \U$22920 ( \23263 , RIbb2ead0_25);
and \U$22921 ( \23264 , \23263 , \10300 );
or \U$22922 ( \23265 , \23262 , \23264 );
not \U$22923 ( \23266 , \23265 );
or \U$22924 ( \23267 , \23261 , \23266 );
nand \U$22925 ( \23268 , \21365 , \2963 );
nand \U$22926 ( \23269 , \23267 , \23268 );
and \U$22927 ( \23270 , \23260 , \23269 );
and \U$22928 ( \23271 , \23249 , \23259 );
or \U$22929 ( \23272 , \23270 , \23271 );
and \U$22930 ( \23273 , \23238 , \23272 );
and \U$22931 ( \23274 , \23235 , \23237 );
or \U$22932 ( \23275 , \23273 , \23274 );
and \U$22933 ( \23276 , \23233 , \23275 );
and \U$22934 ( \23277 , \23094 , \23232 );
or \U$22935 ( \23278 , \23276 , \23277 );
xor \U$22936 ( \23279 , \23092 , \23278 );
xor \U$22937 ( \23280 , \21179 , \21308 );
xor \U$22938 ( \23281 , \23280 , \21342 );
and \U$22939 ( \23282 , \23279 , \23281 );
and \U$22940 ( \23283 , \23092 , \23278 );
or \U$22941 ( \23284 , \23282 , \23283 );
xor \U$22942 ( \23285 , \23090 , \23284 );
xor \U$22943 ( \23286 , \21172 , \21345 );
xor \U$22944 ( \23287 , \23286 , \21507 );
and \U$22945 ( \23288 , \23285 , \23287 );
and \U$22946 ( \23289 , \23090 , \23284 );
or \U$22947 ( \23290 , \23288 , \23289 );
xor \U$22948 ( \23291 , \22665 , \22793 );
xnor \U$22949 ( \23292 , \23291 , \22796 );
xor \U$22950 ( \23293 , \23290 , \23292 );
xor \U$22951 ( \23294 , \21279 , \21289 );
xor \U$22952 ( \23295 , \23294 , \21301 );
not \U$22953 ( \23296 , \23295 );
not \U$22954 ( \23297 , \23296 );
xor \U$22955 ( \23298 , \22750 , \22757 );
xnor \U$22956 ( \23299 , \23298 , \22692 );
not \U$22957 ( \23300 , \23299 );
or \U$22958 ( \23301 , \23297 , \23300 );
xor \U$22959 ( \23302 , \21255 , \21265 );
xor \U$22960 ( \23303 , \23302 , \21276 );
not \U$22961 ( \23304 , \18717 );
not \U$22962 ( \23305 , RIbb2d9f0_61);
not \U$22963 ( \23306 , \5003 );
or \U$22964 ( \23307 , \23305 , \23306 );
nand \U$22965 ( \23308 , \1548 , \16254 );
nand \U$22966 ( \23309 , \23307 , \23308 );
not \U$22967 ( \23310 , \23309 );
or \U$22968 ( \23311 , \23304 , \23310 );
nand \U$22969 ( \23312 , \21451 , \16533 );
nand \U$22970 ( \23313 , \23311 , \23312 );
xor \U$22971 ( \23314 , \23303 , \23313 );
not \U$22972 ( \23315 , \12167 );
not \U$22973 ( \23316 , RIbb2df90_49);
not \U$22974 ( \23317 , \3310 );
or \U$22975 ( \23318 , \23316 , \23317 );
nand \U$22976 ( \23319 , \13280 , \12278 );
nand \U$22977 ( \23320 , \23318 , \23319 );
not \U$22978 ( \23321 , \23320 );
or \U$22979 ( \23322 , \23315 , \23321 );
nand \U$22980 ( \23323 , \21378 , \16427 );
nand \U$22981 ( \23324 , \23322 , \23323 );
and \U$22982 ( \23325 , \23314 , \23324 );
and \U$22983 ( \23326 , \23303 , \23313 );
or \U$22984 ( \23327 , \23325 , \23326 );
nand \U$22985 ( \23328 , \23301 , \23327 );
or \U$22986 ( \23329 , \23299 , \23296 );
nand \U$22987 ( \23330 , \23328 , \23329 );
xor \U$22988 ( \23331 , \21432 , \21467 );
xor \U$22989 ( \23332 , \23331 , \21501 );
xor \U$22990 ( \23333 , \23330 , \23332 );
not \U$22991 ( \23334 , \22804 );
not \U$22992 ( \23335 , \22811 );
or \U$22993 ( \23336 , \23334 , \23335 );
nand \U$22994 ( \23337 , \22803 , \22807 );
nand \U$22995 ( \23338 , \23336 , \23337 );
and \U$22996 ( \23339 , \23338 , \22815 );
not \U$22997 ( \23340 , \23338 );
not \U$22998 ( \23341 , \22815 );
and \U$22999 ( \23342 , \23340 , \23341 );
nor \U$23000 ( \23343 , \23339 , \23342 );
and \U$23001 ( \23344 , \23333 , \23343 );
and \U$23002 ( \23345 , \23330 , \23332 );
or \U$23003 ( \23346 , \23344 , \23345 );
not \U$23004 ( \23347 , \23346 );
not \U$23005 ( \23348 , \23347 );
xor \U$23006 ( \23349 , \22761 , \22773 );
xnor \U$23007 ( \23350 , \23349 , \22781 );
not \U$23008 ( \23351 , \23350 );
or \U$23009 ( \23352 , \23348 , \23351 );
not \U$23010 ( \23353 , \22823 );
not \U$23011 ( \23354 , \23353 );
xor \U$23012 ( \23355 , \22828 , \22817 );
not \U$23013 ( \23356 , \23355 );
or \U$23014 ( \23357 , \23354 , \23356 );
or \U$23015 ( \23358 , \23355 , \23353 );
nand \U$23016 ( \23359 , \23357 , \23358 );
nand \U$23017 ( \23360 , \23352 , \23359 );
not \U$23018 ( \23361 , \23350 );
not \U$23019 ( \23362 , \23347 );
nand \U$23020 ( \23363 , \23361 , \23362 );
nand \U$23021 ( \23364 , \23360 , \23363 );
xor \U$23022 ( \23365 , \22786 , \22783 );
xor \U$23023 ( \23366 , \23365 , \22791 );
xor \U$23024 ( \23367 , \23364 , \23366 );
xor \U$23025 ( \23368 , \22830 , \22833 );
xor \U$23026 ( \23369 , \23368 , \22838 );
and \U$23027 ( \23370 , \23367 , \23369 );
and \U$23028 ( \23371 , \23364 , \23366 );
or \U$23029 ( \23372 , \23370 , \23371 );
xor \U$23030 ( \23373 , \23293 , \23372 );
or \U$23031 ( \23374 , \22879 , \23373 );
not \U$23032 ( \23375 , \831 );
not \U$23033 ( \23376 , RIbb2ee90_17);
not \U$23034 ( \23377 , \18829 );
or \U$23035 ( \23378 , \23376 , \23377 );
nand \U$23036 ( \23379 , \13977 , \3699 );
nand \U$23037 ( \23380 , \23378 , \23379 );
not \U$23038 ( \23381 , \23380 );
or \U$23039 ( \23382 , \23375 , \23381 );
nand \U$23040 ( \23383 , \22745 , \836 );
nand \U$23041 ( \23384 , \23382 , \23383 );
not \U$23042 ( \23385 , \1444 );
and \U$23043 ( \23386 , RIbb2ef80_15, \15471 );
not \U$23044 ( \23387 , RIbb2ef80_15);
and \U$23045 ( \23388 , \23387 , \15470 );
or \U$23046 ( \23389 , \23386 , \23388 );
not \U$23047 ( \23390 , \23389 );
or \U$23048 ( \23391 , \23385 , \23390 );
nand \U$23049 ( \23392 , \23109 , \1517 );
nand \U$23050 ( \23393 , \23391 , \23392 );
xor \U$23051 ( \23394 , \23384 , \23393 );
not \U$23052 ( \23395 , \3613 );
not \U$23053 ( \23396 , \23214 );
or \U$23054 ( \23397 , \23395 , \23396 );
not \U$23055 ( \23398 , RIbb2e800_31);
not \U$23056 ( \23399 , \7296 );
not \U$23057 ( \23400 , \23399 );
or \U$23058 ( \23401 , \23398 , \23400 );
nand \U$23059 ( \23402 , \7296 , \4096 );
nand \U$23060 ( \23403 , \23401 , \23402 );
nand \U$23061 ( \23404 , \23403 , \2939 );
nand \U$23062 ( \23405 , \23397 , \23404 );
and \U$23063 ( \23406 , \23394 , \23405 );
and \U$23064 ( \23407 , \23384 , \23393 );
or \U$23065 ( \23408 , \23406 , \23407 );
not \U$23066 ( \23409 , \23408 );
xor \U$23067 ( \23410 , \22711 , \22736 );
xor \U$23068 ( \23411 , \23410 , \22747 );
not \U$23069 ( \23412 , \23411 );
nand \U$23070 ( \23413 , \23409 , \23412 );
not \U$23071 ( \23414 , \2078 );
not \U$23072 ( \23415 , \23247 );
or \U$23073 ( \23416 , \23414 , \23415 );
not \U$23074 ( \23417 , RIbb2ecb0_21);
not \U$23075 ( \23418 , \17663 );
or \U$23076 ( \23419 , \23417 , \23418 );
nand \U$23077 ( \23420 , \12932 , \849 );
nand \U$23078 ( \23421 , \23419 , \23420 );
nand \U$23079 ( \23422 , \23421 , \2077 );
nand \U$23080 ( \23423 , \23416 , \23422 );
not \U$23081 ( \23424 , \854 );
not \U$23082 ( \23425 , \23120 );
or \U$23083 ( \23426 , \23424 , \23425 );
not \U$23084 ( \23427 , RIbb2eda0_19);
not \U$23085 ( \23428 , \14624 );
or \U$23086 ( \23429 , \23427 , \23428 );
nand \U$23087 ( \23430 , \13210 , \3251 );
nand \U$23088 ( \23431 , \23429 , \23430 );
nand \U$23089 ( \23432 , \23431 , \853 );
nand \U$23090 ( \23433 , \23426 , \23432 );
or \U$23091 ( \23434 , \23423 , \23433 );
xor \U$23092 ( \23435 , \22712 , \22722 );
xor \U$23093 ( \23436 , \23435 , \22733 );
nand \U$23094 ( \23437 , \23434 , \23436 );
nand \U$23095 ( \23438 , \23423 , \23433 );
nand \U$23096 ( \23439 , \23437 , \23438 );
and \U$23097 ( \23440 , \23413 , \23439 );
not \U$23098 ( \23441 , \23408 );
nor \U$23099 ( \23442 , \23441 , \23412 );
nor \U$23100 ( \23443 , \23440 , \23442 );
not \U$23101 ( \23444 , \23443 );
xor \U$23102 ( \23445 , \21429 , \21419 );
xnor \U$23103 ( \23446 , \23445 , \21410 );
not \U$23104 ( \23447 , \23446 );
or \U$23105 ( \23448 , \23444 , \23447 );
xor \U$23106 ( \23449 , \23104 , \23113 );
xor \U$23107 ( \23450 , \23449 , \23124 );
not \U$23108 ( \23451 , \23450 );
not \U$23109 ( \23452 , \23451 );
not \U$23110 ( \23453 , \3382 );
not \U$23111 ( \23454 , \23257 );
or \U$23112 ( \23455 , \23453 , \23454 );
and \U$23113 ( \23456 , \11578 , \3401 );
not \U$23114 ( \23457 , \11578 );
and \U$23115 ( \23458 , \23457 , RIbb2ebc0_23);
or \U$23116 ( \23459 , \23456 , \23458 );
nand \U$23117 ( \23460 , \23459 , \3406 );
nand \U$23118 ( \23461 , \23455 , \23460 );
not \U$23119 ( \23462 , \23461 );
not \U$23120 ( \23463 , \4075 );
not \U$23121 ( \23464 , \23134 );
or \U$23122 ( \23465 , \23463 , \23464 );
not \U$23123 ( \23466 , RIbb2e710_33);
not \U$23124 ( \23467 , \8337 );
or \U$23125 ( \23468 , \23466 , \23467 );
nand \U$23126 ( \23469 , \15796 , \16803 );
nand \U$23127 ( \23470 , \23468 , \23469 );
nand \U$23128 ( \23471 , \23470 , \3886 );
nand \U$23129 ( \23472 , \23465 , \23471 );
not \U$23130 ( \23473 , \23472 );
or \U$23131 ( \23474 , \23462 , \23473 );
or \U$23132 ( \23475 , \23461 , \23472 );
not \U$23133 ( \23476 , \6241 );
not \U$23134 ( \23477 , \23018 );
or \U$23135 ( \23478 , \23476 , \23477 );
not \U$23136 ( \23479 , RIbb2e530_37);
not \U$23137 ( \23480 , \13559 );
or \U$23138 ( \23481 , \23479 , \23480 );
nand \U$23139 ( \23482 , \4390 , \4708 );
nand \U$23140 ( \23483 , \23481 , \23482 );
nand \U$23141 ( \23484 , \23483 , \6251 );
nand \U$23142 ( \23485 , \23478 , \23484 );
nand \U$23143 ( \23486 , \23475 , \23485 );
nand \U$23144 ( \23487 , \23474 , \23486 );
not \U$23145 ( \23488 , \23487 );
not \U$23146 ( \23489 , \23488 );
or \U$23147 ( \23490 , \23452 , \23489 );
xor \U$23148 ( \23491 , \23170 , \23179 );
not \U$23149 ( \23492 , \1570 );
not \U$23150 ( \23493 , \22729 );
or \U$23151 ( \23494 , \23492 , \23493 );
not \U$23152 ( \23495 , RIbb2f250_9);
not \U$23153 ( \23496 , \16819 );
or \U$23154 ( \23497 , \23495 , \23496 );
nand \U$23155 ( \23498 , \17529 , \1566 );
nand \U$23156 ( \23499 , \23497 , \23498 );
nand \U$23157 ( \23500 , \23499 , \1533 );
nand \U$23158 ( \23501 , \23494 , \23500 );
xor \U$23159 ( \23502 , \23491 , \23501 );
not \U$23160 ( \23503 , \1077 );
not \U$23161 ( \23504 , \23189 );
or \U$23162 ( \23505 , \23503 , \23504 );
not \U$23163 ( \23506 , RIbb2f160_11);
not \U$23164 ( \23507 , \16710 );
or \U$23165 ( \23508 , \23506 , \23507 );
nand \U$23166 ( \23509 , \16553 , \1805 );
nand \U$23167 ( \23510 , \23508 , \23509 );
nand \U$23168 ( \23511 , \23510 , \1011 );
nand \U$23169 ( \23512 , \23505 , \23511 );
and \U$23170 ( \23513 , \23502 , \23512 );
and \U$23171 ( \23514 , \23491 , \23501 );
or \U$23172 ( \23515 , \23513 , \23514 );
not \U$23173 ( \23516 , \3465 );
not \U$23174 ( \23517 , \23155 );
or \U$23175 ( \23518 , \23516 , \23517 );
not \U$23176 ( \23519 , RIbb2e9e0_27);
not \U$23177 ( \23520 , \14550 );
or \U$23178 ( \23521 , \23519 , \23520 );
nand \U$23179 ( \23522 , \9841 , \3454 );
nand \U$23180 ( \23523 , \23521 , \23522 );
nand \U$23181 ( \23524 , \23523 , \3445 );
nand \U$23182 ( \23525 , \23518 , \23524 );
xor \U$23183 ( \23526 , \23515 , \23525 );
not \U$23184 ( \23527 , \2922 );
not \U$23185 ( \23528 , RIbb2e8f0_29);
not \U$23186 ( \23529 , \8630 );
not \U$23187 ( \23530 , \23529 );
or \U$23188 ( \23531 , \23528 , \23530 );
nand \U$23189 ( \23532 , \13866 , \3265 );
nand \U$23190 ( \23533 , \23531 , \23532 );
not \U$23191 ( \23534 , \23533 );
or \U$23192 ( \23535 , \23527 , \23534 );
nand \U$23193 ( \23536 , \23146 , \2925 );
nand \U$23194 ( \23537 , \23535 , \23536 );
and \U$23195 ( \23538 , \23526 , \23537 );
and \U$23196 ( \23539 , \23515 , \23525 );
or \U$23197 ( \23540 , \23538 , \23539 );
nand \U$23198 ( \23541 , \23490 , \23540 );
not \U$23199 ( \23542 , \23488 );
nand \U$23200 ( \23543 , \23542 , \23450 );
nand \U$23201 ( \23544 , \23541 , \23543 );
nand \U$23202 ( \23545 , \23448 , \23544 );
not \U$23203 ( \23546 , \23446 );
not \U$23204 ( \23547 , \23443 );
nand \U$23205 ( \23548 , \23546 , \23547 );
nand \U$23206 ( \23549 , \23545 , \23548 );
not \U$23207 ( \23550 , \23549 );
not \U$23208 ( \23551 , \22678 );
not \U$23209 ( \23552 , \22759 );
and \U$23210 ( \23553 , \23551 , \23552 );
and \U$23211 ( \23554 , \22759 , \22678 );
nor \U$23212 ( \23555 , \23553 , \23554 );
not \U$23213 ( \23556 , \22672 );
and \U$23214 ( \23557 , \23555 , \23556 );
not \U$23215 ( \23558 , \23555 );
and \U$23216 ( \23559 , \23558 , \22672 );
nor \U$23217 ( \23560 , \23557 , \23559 );
not \U$23218 ( \23561 , \23560 );
nand \U$23219 ( \23562 , \23550 , \23561 );
not \U$23220 ( \23563 , \23562 );
xor \U$23221 ( \23564 , \23235 , \23237 );
xor \U$23222 ( \23565 , \23564 , \23272 );
buf \U$23223 ( \23566 , \23565 );
not \U$23224 ( \23567 , \23566 );
xor \U$23225 ( \23568 , \23249 , \23259 );
xor \U$23226 ( \23569 , \23568 , \23269 );
not \U$23227 ( \23570 , \23569 );
not \U$23228 ( \23571 , \8354 );
not \U$23229 ( \23572 , \22898 );
or \U$23230 ( \23573 , \23571 , \23572 );
not \U$23231 ( \23574 , RIbb2e350_41);
not \U$23232 ( \23575 , \4028 );
or \U$23233 ( \23576 , \23574 , \23575 );
nand \U$23234 ( \23577 , \3044 , \13392 );
nand \U$23235 ( \23578 , \23576 , \23577 );
nand \U$23236 ( \23579 , \23578 , \8362 );
nand \U$23237 ( \23580 , \23573 , \23579 );
not \U$23238 ( \23581 , \8450 );
not \U$23239 ( \23582 , \22920 );
or \U$23240 ( \23583 , \23581 , \23582 );
xor \U$23241 ( \23584 , RIbb2e440_39, \3089 );
nand \U$23242 ( \23585 , \23584 , \7103 );
nand \U$23243 ( \23586 , \23583 , \23585 );
xor \U$23244 ( \23587 , \23580 , \23586 );
not \U$23245 ( \23588 , \17563 );
not \U$23246 ( \23589 , RIbb2ddb0_53);
not \U$23247 ( \23590 , \22684 );
or \U$23248 ( \23591 , \23589 , \23590 );
nand \U$23249 ( \23592 , \1419 , \13463 );
nand \U$23250 ( \23593 , \23591 , \23592 );
not \U$23251 ( \23594 , \23593 );
or \U$23252 ( \23595 , \23588 , \23594 );
nand \U$23253 ( \23596 , \22910 , \14930 );
nand \U$23254 ( \23597 , \23595 , \23596 );
and \U$23255 ( \23598 , \23587 , \23597 );
and \U$23256 ( \23599 , \23580 , \23586 );
or \U$23257 ( \23600 , \23598 , \23599 );
not \U$23258 ( \23601 , \23600 );
or \U$23259 ( \23602 , \23570 , \23601 );
or \U$23260 ( \23603 , \23600 , \23569 );
xor \U$23261 ( \23604 , \23180 , \23191 );
xor \U$23262 ( \23605 , \23604 , \23203 );
not \U$23263 ( \23606 , \17275 );
not \U$23264 ( \23607 , RIbb2d900_63);
not \U$23265 ( \23608 , \16207 );
or \U$23266 ( \23609 , \23607 , \23608 );
nand \U$23267 ( \23610 , \1037 , \17270 );
nand \U$23268 ( \23611 , \23609 , \23610 );
not \U$23269 ( \23612 , \23611 );
or \U$23270 ( \23613 , \23606 , \23612 );
nand \U$23271 ( \23614 , \22948 , RIbb2d888_64);
nand \U$23272 ( \23615 , \23613 , \23614 );
xor \U$23273 ( \23616 , \23605 , \23615 );
not \U$23274 ( \23617 , \12692 );
not \U$23275 ( \23618 , \23006 );
or \U$23276 ( \23619 , \23617 , \23618 );
not \U$23277 ( \23620 , RIbb2dea0_51);
not \U$23278 ( \23621 , \20325 );
or \U$23279 ( \23622 , \23620 , \23621 );
not \U$23280 ( \23623 , RIbb2dea0_51);
nand \U$23281 ( \23624 , \23623 , \1851 );
nand \U$23282 ( \23625 , \23622 , \23624 );
nand \U$23283 ( \23626 , \23625 , \12774 );
nand \U$23284 ( \23627 , \23619 , \23626 );
and \U$23285 ( \23628 , \23616 , \23627 );
and \U$23286 ( \23629 , \23605 , \23615 );
or \U$23287 ( \23630 , \23628 , \23629 );
nand \U$23288 ( \23631 , \23603 , \23630 );
nand \U$23289 ( \23632 , \23602 , \23631 );
not \U$23290 ( \23633 , \23632 );
or \U$23291 ( \23634 , \23567 , \23633 );
or \U$23292 ( \23635 , \23632 , \23566 );
not \U$23293 ( \23636 , \4714 );
not \U$23294 ( \23637 , \23223 );
or \U$23295 ( \23638 , \23636 , \23637 );
not \U$23296 ( \23639 , \4713 );
not \U$23297 ( \23640 , RIbb2e620_35);
not \U$23298 ( \23641 , \6230 );
or \U$23299 ( \23642 , \23640 , \23641 );
nand \U$23300 ( \23643 , \6229 , \6002 );
nand \U$23301 ( \23644 , \23642 , \23643 );
nand \U$23302 ( \23645 , \23639 , \23644 );
nand \U$23303 ( \23646 , \23638 , \23645 );
not \U$23304 ( \23647 , \23646 );
not \U$23305 ( \23648 , \23647 );
not \U$23306 ( \23649 , \2963 );
not \U$23307 ( \23650 , \23265 );
or \U$23308 ( \23651 , \23649 , \23650 );
and \U$23309 ( \23652 , RIbb2ead0_25, \18802 );
not \U$23310 ( \23653 , RIbb2ead0_25);
and \U$23311 ( \23654 , \23653 , \13525 );
or \U$23312 ( \23655 , \23652 , \23654 );
nand \U$23313 ( \23656 , \23655 , \2980 );
nand \U$23314 ( \23657 , \23651 , \23656 );
not \U$23315 ( \23658 , \23657 );
not \U$23316 ( \23659 , \23658 );
or \U$23317 ( \23660 , \23648 , \23659 );
not \U$23318 ( \23661 , \16533 );
not \U$23319 ( \23662 , \23309 );
or \U$23320 ( \23663 , \23661 , \23662 );
not \U$23321 ( \23664 , RIbb2d9f0_61);
not \U$23322 ( \23665 , \14819 );
or \U$23323 ( \23666 , \23664 , \23665 );
nand \U$23324 ( \23667 , \14818 , \19746 );
nand \U$23325 ( \23668 , \23666 , \23667 );
nand \U$23326 ( \23669 , \23668 , \16541 );
nand \U$23327 ( \23670 , \23663 , \23669 );
nand \U$23328 ( \23671 , \23660 , \23670 );
not \U$23329 ( \23672 , \23658 );
nand \U$23330 ( \23673 , \23672 , \23646 );
nand \U$23331 ( \23674 , \23671 , \23673 );
xor \U$23332 ( \23675 , \23206 , \23216 );
xor \U$23333 ( \23676 , \23675 , \23227 );
xor \U$23334 ( \23677 , \23674 , \23676 );
not \U$23335 ( \23678 , \9098 );
not \U$23336 ( \23679 , RIbb2e260_43);
not \U$23337 ( \23680 , \21490 );
or \U$23338 ( \23681 , \23679 , \23680 );
nand \U$23339 ( \23682 , \3653 , \8347 );
nand \U$23340 ( \23683 , \23681 , \23682 );
not \U$23341 ( \23684 , \23683 );
or \U$23342 ( \23685 , \23678 , \23684 );
nand \U$23343 ( \23686 , \22935 , \10451 );
nand \U$23344 ( \23687 , \23685 , \23686 );
not \U$23345 ( \23688 , \15181 );
not \U$23346 ( \23689 , \22957 );
or \U$23347 ( \23690 , \23688 , \23689 );
and \U$23348 ( \23691 , RIbb2dcc0_55, \3990 );
not \U$23349 ( \23692 , RIbb2dcc0_55);
and \U$23350 ( \23693 , \23692 , \1169 );
or \U$23351 ( \23694 , \23691 , \23693 );
nand \U$23352 ( \23695 , \23694 , \14613 );
nand \U$23353 ( \23696 , \23690 , \23695 );
xor \U$23354 ( \23697 , \23687 , \23696 );
not \U$23355 ( \23698 , \10119 );
not \U$23356 ( \23699 , \22982 );
or \U$23357 ( \23700 , \23698 , \23699 );
not \U$23358 ( \23701 , RIbb2e170_45);
not \U$23359 ( \23702 , \16399 );
or \U$23360 ( \23703 , \23701 , \23702 );
nand \U$23361 ( \23704 , \16400 , \12003 );
nand \U$23362 ( \23705 , \23703 , \23704 );
nand \U$23363 ( \23706 , \23705 , \10117 );
nand \U$23364 ( \23707 , \23700 , \23706 );
and \U$23365 ( \23708 , \23697 , \23707 );
and \U$23366 ( \23709 , \23687 , \23696 );
or \U$23367 ( \23710 , \23708 , \23709 );
and \U$23368 ( \23711 , \23677 , \23710 );
and \U$23369 ( \23712 , \23674 , \23676 );
or \U$23370 ( \23713 , \23711 , \23712 );
nand \U$23371 ( \23714 , \23635 , \23713 );
nand \U$23372 ( \23715 , \23634 , \23714 );
not \U$23373 ( \23716 , \23715 );
or \U$23374 ( \23717 , \23563 , \23716 );
not \U$23375 ( \23718 , \23561 );
nand \U$23376 ( \23719 , \23718 , \23549 );
nand \U$23377 ( \23720 , \23717 , \23719 );
xor \U$23378 ( \23721 , \23092 , \23278 );
xor \U$23379 ( \23722 , \23721 , \23281 );
xor \U$23380 ( \23723 , \23720 , \23722 );
xor \U$23381 ( \23724 , \23094 , \23232 );
xor \U$23382 ( \23725 , \23724 , \23275 );
nand \U$23383 ( \23726 , \22885 , \22882 );
and \U$23384 ( \23727 , \22926 , \23726 );
and \U$23385 ( \23728 , \23048 , \23727 );
not \U$23386 ( \23729 , \23048 );
and \U$23387 ( \23730 , \23729 , \22927 );
nor \U$23388 ( \23731 , \23728 , \23730 );
and \U$23389 ( \23732 , \23731 , \23036 );
not \U$23390 ( \23733 , \23731 );
not \U$23391 ( \23734 , \23036 );
and \U$23392 ( \23735 , \23733 , \23734 );
nor \U$23393 ( \23736 , \23732 , \23735 );
xor \U$23394 ( \23737 , \23725 , \23736 );
xnor \U$23395 ( \23738 , \23230 , \23127 );
not \U$23396 ( \23739 , \23162 );
and \U$23397 ( \23740 , \23738 , \23739 );
not \U$23398 ( \23741 , \23738 );
and \U$23399 ( \23742 , \23741 , \23162 );
nor \U$23400 ( \23743 , \23740 , \23742 );
xor \U$23401 ( \23744 , \23295 , \23299 );
xnor \U$23402 ( \23745 , \23744 , \23327 );
xor \U$23403 ( \23746 , \23743 , \23745 );
xor \U$23404 ( \23747 , \23138 , \23148 );
xor \U$23405 ( \23748 , \23747 , \23159 );
not \U$23406 ( \23749 , \19101 );
not \U$23407 ( \23750 , RIbb2dbd0_57);
not \U$23408 ( \23751 , \4766 );
or \U$23409 ( \23752 , \23750 , \23751 );
nand \U$23410 ( \23753 , \4769 , \15741 );
nand \U$23411 ( \23754 , \23752 , \23753 );
not \U$23412 ( \23755 , \23754 );
or \U$23413 ( \23756 , \23749 , \23755 );
nand \U$23414 ( \23757 , \15738 , \22971 );
nand \U$23415 ( \23758 , \23756 , \23757 );
not \U$23416 ( \23759 , \23758 );
not \U$23417 ( \23760 , \11176 );
not \U$23418 ( \23761 , RIbb2e080_47);
not \U$23419 ( \23762 , \3168 );
or \U$23420 ( \23763 , \23761 , \23762 );
nand \U$23421 ( \23764 , \3951 , \12971 );
nand \U$23422 ( \23765 , \23763 , \23764 );
not \U$23423 ( \23766 , \23765 );
or \U$23424 ( \23767 , \23760 , \23766 );
nand \U$23425 ( \23768 , \22993 , \12965 );
nand \U$23426 ( \23769 , \23767 , \23768 );
not \U$23427 ( \23770 , \23769 );
or \U$23428 ( \23771 , \23759 , \23770 );
or \U$23429 ( \23772 , \23769 , \23758 );
not \U$23430 ( \23773 , \12167 );
not \U$23431 ( \23774 , RIbb2df90_49);
not \U$23432 ( \23775 , \2223 );
or \U$23433 ( \23776 , \23774 , \23775 );
nand \U$23434 ( \23777 , \13290 , \12278 );
nand \U$23435 ( \23778 , \23776 , \23777 );
not \U$23436 ( \23779 , \23778 );
or \U$23437 ( \23780 , \23773 , \23779 );
nand \U$23438 ( \23781 , \23320 , \12284 );
nand \U$23439 ( \23782 , \23780 , \23781 );
nand \U$23440 ( \23783 , \23772 , \23782 );
nand \U$23441 ( \23784 , \23771 , \23783 );
xor \U$23442 ( \23785 , \23748 , \23784 );
xor \U$23443 ( \23786 , \22975 , \22986 );
xor \U$23444 ( \23787 , \23786 , \22997 );
and \U$23445 ( \23788 , \23785 , \23787 );
and \U$23446 ( \23789 , \23748 , \23784 );
or \U$23447 ( \23790 , \23788 , \23789 );
and \U$23448 ( \23791 , \23746 , \23790 );
and \U$23449 ( \23792 , \23743 , \23745 );
or \U$23450 ( \23793 , \23791 , \23792 );
and \U$23451 ( \23794 , \23737 , \23793 );
and \U$23452 ( \23795 , \23725 , \23736 );
or \U$23453 ( \23796 , \23794 , \23795 );
and \U$23454 ( \23797 , \23723 , \23796 );
and \U$23455 ( \23798 , \23720 , \23722 );
or \U$23456 ( \23799 , \23797 , \23798 );
not \U$23457 ( \23800 , \23799 );
xor \U$23458 ( \23801 , \23090 , \23284 );
xor \U$23459 ( \23802 , \23801 , \23287 );
not \U$23460 ( \23803 , \23802 );
or \U$23461 ( \23804 , \23800 , \23803 );
not \U$23462 ( \23805 , \23799 );
not \U$23463 ( \23806 , \23805 );
not \U$23464 ( \23807 , \23802 );
not \U$23465 ( \23808 , \23807 );
or \U$23466 ( \23809 , \23806 , \23808 );
xor \U$23467 ( \23810 , \23364 , \23366 );
xor \U$23468 ( \23811 , \23810 , \23369 );
nand \U$23469 ( \23812 , \23809 , \23811 );
nand \U$23470 ( \23813 , \23804 , \23812 );
buf \U$23471 ( \23814 , \23813 );
nand \U$23472 ( \23815 , \23374 , \23814 );
not \U$23473 ( \23816 , \22878 );
nand \U$23474 ( \23817 , \23816 , \23373 );
nand \U$23475 ( \23818 , \23815 , \23817 );
not \U$23476 ( \23819 , \23818 );
xor \U$23477 ( \23820 , \21512 , \21520 );
xor \U$23478 ( \23821 , \23820 , \21531 );
xor \U$23479 ( \23822 , \22798 , \22800 );
xor \U$23480 ( \23823 , \23822 , \22861 );
xor \U$23481 ( \23824 , \23821 , \23823 );
xor \U$23482 ( \23825 , \23290 , \23292 );
and \U$23483 ( \23826 , \23825 , \23372 );
and \U$23484 ( \23827 , \23290 , \23292 );
or \U$23485 ( \23828 , \23826 , \23827 );
xor \U$23486 ( \23829 , \23824 , \23828 );
not \U$23487 ( \23830 , \23829 );
or \U$23488 ( \23831 , \23819 , \23830 );
xor \U$23489 ( \23832 , \22877 , \23813 );
xnor \U$23490 ( \23833 , \23832 , \23373 );
not \U$23491 ( \23834 , \23799 );
not \U$23492 ( \23835 , \23807 );
or \U$23493 ( \23836 , \23834 , \23835 );
nand \U$23494 ( \23837 , \23802 , \23805 );
nand \U$23495 ( \23838 , \23836 , \23837 );
and \U$23496 ( \23839 , \23838 , \23811 );
not \U$23497 ( \23840 , \23838 );
not \U$23498 ( \23841 , \23811 );
and \U$23499 ( \23842 , \23840 , \23841 );
nor \U$23500 ( \23843 , \23839 , \23842 );
not \U$23501 ( \23844 , \23843 );
xor \U$23502 ( \23845 , \23515 , \23525 );
xor \U$23503 ( \23846 , \23845 , \23537 );
xor \U$23504 ( \23847 , \23461 , \23472 );
xor \U$23505 ( \23848 , \23847 , \23485 );
xor \U$23506 ( \23849 , \23846 , \23848 );
not \U$23507 ( \23850 , \16675 );
not \U$23508 ( \23851 , RIbb2dbd0_57);
not \U$23509 ( \23852 , \12037 );
or \U$23510 ( \23853 , \23851 , \23852 );
nand \U$23511 ( \23854 , \12036 , \17411 );
nand \U$23512 ( \23855 , \23853 , \23854 );
not \U$23513 ( \23856 , \23855 );
or \U$23514 ( \23857 , \23850 , \23856 );
nand \U$23515 ( \23858 , \23754 , \17100 );
nand \U$23516 ( \23859 , \23857 , \23858 );
not \U$23517 ( \23860 , \11176 );
not \U$23518 ( \23861 , \17568 );
xor \U$23519 ( \23862 , RIbb2e080_47, \23861 );
not \U$23520 ( \23863 , \23862 );
or \U$23521 ( \23864 , \23860 , \23863 );
nand \U$23522 ( \23865 , \23765 , \12965 );
nand \U$23523 ( \23866 , \23864 , \23865 );
or \U$23524 ( \23867 , \23859 , \23866 );
not \U$23525 ( \23868 , \10599 );
not \U$23526 ( \23869 , RIbb2e170_45);
not \U$23527 ( \23870 , \3225 );
or \U$23528 ( \23871 , \23869 , \23870 );
nand \U$23529 ( \23872 , \3224 , \12003 );
nand \U$23530 ( \23873 , \23871 , \23872 );
not \U$23531 ( \23874 , \23873 );
or \U$23532 ( \23875 , \23868 , \23874 );
nand \U$23533 ( \23876 , \23705 , \10119 );
nand \U$23534 ( \23877 , \23875 , \23876 );
nand \U$23535 ( \23878 , \23867 , \23877 );
nand \U$23536 ( \23879 , \23866 , \23859 );
nand \U$23537 ( \23880 , \23878 , \23879 );
and \U$23538 ( \23881 , \23849 , \23880 );
and \U$23539 ( \23882 , \23846 , \23848 );
or \U$23540 ( \23883 , \23881 , \23882 );
not \U$23541 ( \23884 , \23883 );
not \U$23542 ( \23885 , \3886 );
not \U$23543 ( \23886 , RIbb2e710_33);
not \U$23544 ( \23887 , \19868 );
or \U$23545 ( \23888 , \23886 , \23887 );
nand \U$23546 ( \23889 , \8637 , \12019 );
nand \U$23547 ( \23890 , \23888 , \23889 );
not \U$23548 ( \23891 , \23890 );
or \U$23549 ( \23892 , \23885 , \23891 );
nand \U$23550 ( \23893 , \23470 , \4790 );
nand \U$23551 ( \23894 , \23892 , \23893 );
not \U$23552 ( \23895 , \4712 );
not \U$23553 ( \23896 , RIbb2e620_35);
not \U$23554 ( \23897 , \18564 );
or \U$23555 ( \23898 , \23896 , \23897 );
nand \U$23556 ( \23899 , \5954 , \3866 );
nand \U$23557 ( \23900 , \23898 , \23899 );
not \U$23558 ( \23901 , \23900 );
or \U$23559 ( \23902 , \23895 , \23901 );
nand \U$23560 ( \23903 , \23644 , \4714 );
nand \U$23561 ( \23904 , \23902 , \23903 );
xor \U$23562 ( \23905 , \23894 , \23904 );
not \U$23563 ( \23906 , \2980 );
not \U$23564 ( \23907 , RIbb2ead0_25);
not \U$23565 ( \23908 , \12260 );
or \U$23566 ( \23909 , \23907 , \23908 );
not \U$23567 ( \23910 , \11143 );
nand \U$23568 ( \23911 , \23910 , \18636 );
nand \U$23569 ( \23912 , \23909 , \23911 );
not \U$23570 ( \23913 , \23912 );
or \U$23571 ( \23914 , \23906 , \23913 );
nand \U$23572 ( \23915 , \23655 , \2963 );
nand \U$23573 ( \23916 , \23914 , \23915 );
and \U$23574 ( \23917 , \23905 , \23916 );
and \U$23575 ( \23918 , \23894 , \23904 );
or \U$23576 ( \23919 , \23917 , \23918 );
not \U$23577 ( \23920 , \23919 );
not \U$23578 ( \23921 , \3382 );
not \U$23579 ( \23922 , \23459 );
or \U$23580 ( \23923 , \23921 , \23922 );
not \U$23581 ( \23924 , RIbb2ebc0_23);
not \U$23582 ( \23925 , \23243 );
or \U$23583 ( \23926 , \23924 , \23925 );
nand \U$23584 ( \23927 , \12174 , \3396 );
nand \U$23585 ( \23928 , \23926 , \23927 );
nand \U$23586 ( \23929 , \23928 , \3406 );
nand \U$23587 ( \23930 , \23923 , \23929 );
not \U$23588 ( \23931 , \20792 );
not \U$23589 ( \23932 , \23483 );
or \U$23590 ( \23933 , \23931 , \23932 );
not \U$23591 ( \23934 , RIbb2e530_37);
not \U$23592 ( \23935 , \4696 );
or \U$23593 ( \23936 , \23934 , \23935 );
nand \U$23594 ( \23937 , \4695 , \4708 );
nand \U$23595 ( \23938 , \23936 , \23937 );
nand \U$23596 ( \23939 , \23938 , \6251 );
nand \U$23597 ( \23940 , \23933 , \23939 );
xor \U$23598 ( \23941 , \23930 , \23940 );
not \U$23599 ( \23942 , \3465 );
not \U$23600 ( \23943 , \23523 );
or \U$23601 ( \23944 , \23942 , \23943 );
not \U$23602 ( \23945 , RIbb2e9e0_27);
not \U$23603 ( \23946 , \15106 );
or \U$23604 ( \23947 , \23945 , \23946 );
nand \U$23605 ( \23948 , \10301 , \4598 );
nand \U$23606 ( \23949 , \23947 , \23948 );
nand \U$23607 ( \23950 , \23949 , \3445 );
nand \U$23608 ( \23951 , \23944 , \23950 );
and \U$23609 ( \23952 , \23941 , \23951 );
and \U$23610 ( \23953 , \23930 , \23940 );
or \U$23611 ( \23954 , \23952 , \23953 );
not \U$23612 ( \23955 , \23954 );
or \U$23613 ( \23956 , \23920 , \23955 );
or \U$23614 ( \23957 , \23954 , \23919 );
not \U$23615 ( \23958 , \2939 );
not \U$23616 ( \23959 , RIbb2e800_31);
not \U$23617 ( \23960 , \8318 );
not \U$23618 ( \23961 , \23960 );
or \U$23619 ( \23962 , \23959 , \23961 );
nand \U$23620 ( \23963 , \8318 , \8810 );
nand \U$23621 ( \23964 , \23962 , \23963 );
not \U$23622 ( \23965 , \23964 );
or \U$23623 ( \23966 , \23958 , \23965 );
nand \U$23624 ( \23967 , \23403 , \3613 );
nand \U$23625 ( \23968 , \23966 , \23967 );
not \U$23626 ( \23969 , \23968 );
not \U$23627 ( \23970 , \2925 );
not \U$23628 ( \23971 , \23533 );
or \U$23629 ( \23972 , \23970 , \23971 );
not \U$23630 ( \23973 , RIbb2e8f0_29);
not \U$23631 ( \23974 , \12819 );
or \U$23632 ( \23975 , \23973 , \23974 );
nand \U$23633 ( \23976 , \9277 , \2911 );
nand \U$23634 ( \23977 , \23975 , \23976 );
nand \U$23635 ( \23978 , \23977 , \2922 );
nand \U$23636 ( \23979 , \23972 , \23978 );
not \U$23637 ( \23980 , \23979 );
or \U$23638 ( \23981 , \23969 , \23980 );
or \U$23639 ( \23982 , \23979 , \23968 );
not \U$23640 ( \23983 , \1531 );
not \U$23641 ( \23984 , RIbb2f250_9);
not \U$23642 ( \23985 , \17744 );
or \U$23643 ( \23986 , \23984 , \23985 );
nand \U$23644 ( \23987 , \17517 , \1554 );
nand \U$23645 ( \23988 , \23986 , \23987 );
not \U$23646 ( \23989 , \23988 );
or \U$23647 ( \23990 , \23983 , \23989 );
not \U$23648 ( \23991 , RIbb2f250_9);
not \U$23649 ( \23992 , \19063 );
or \U$23650 ( \23993 , \23991 , \23992 );
nand \U$23651 ( \23994 , \17506 , \1554 );
nand \U$23652 ( \23995 , \23993 , \23994 );
nand \U$23653 ( \23996 , \23995 , \1532 );
nand \U$23654 ( \23997 , \23990 , \23996 );
nand \U$23655 ( \23998 , \1805 , \1525 );
and \U$23656 ( \23999 , \19064 , \23998 );
not \U$23657 ( \24000 , RIbb2f160_11);
not \U$23658 ( \24001 , RIbb2f1d8_10);
or \U$23659 ( \24002 , \24000 , \24001 );
nand \U$23660 ( \24003 , \24002 , RIbb2f250_9);
nor \U$23661 ( \24004 , \23999 , \24003 );
and \U$23662 ( \24005 , \23997 , \24004 );
not \U$23663 ( \24006 , \998 );
not \U$23664 ( \24007 , RIbb2f070_13);
not \U$23665 ( \24008 , \16746 );
or \U$23666 ( \24009 , \24007 , \24008 );
not \U$23667 ( \24010 , \16746 );
nand \U$23668 ( \24011 , \24010 , \1656 );
nand \U$23669 ( \24012 , \24009 , \24011 );
not \U$23670 ( \24013 , \24012 );
or \U$23671 ( \24014 , \24006 , \24013 );
not \U$23672 ( \24015 , RIbb2f070_13);
not \U$23673 ( \24016 , \16727 );
or \U$23674 ( \24017 , \24015 , \24016 );
nand \U$23675 ( \24018 , \1656 , \16726 );
nand \U$23676 ( \24019 , \24017 , \24018 );
nand \U$23677 ( \24020 , \24019 , \915 );
nand \U$23678 ( \24021 , \24014 , \24020 );
xor \U$23679 ( \24022 , \24005 , \24021 );
not \U$23680 ( \24023 , \1517 );
not \U$23681 ( \24024 , RIbb2ef80_15);
not \U$23682 ( \24025 , \16561 );
or \U$23683 ( \24026 , \24024 , \24025 );
not \U$23684 ( \24027 , RIbb2ef80_15);
nand \U$23685 ( \24028 , \24027 , \15752 );
nand \U$23686 ( \24029 , \24026 , \24028 );
not \U$23687 ( \24030 , \24029 );
or \U$23688 ( \24031 , \24023 , \24030 );
and \U$23689 ( \24032 , RIbb2ef80_15, \23197 );
not \U$23690 ( \24033 , RIbb2ef80_15);
and \U$23691 ( \24034 , \24033 , \16575 );
or \U$23692 ( \24035 , \24032 , \24034 );
nand \U$23693 ( \24036 , \24035 , \1444 );
nand \U$23694 ( \24037 , \24031 , \24036 );
and \U$23695 ( \24038 , \24022 , \24037 );
and \U$23696 ( \24039 , \24005 , \24021 );
or \U$23697 ( \24040 , \24038 , \24039 );
nand \U$23698 ( \24041 , \23982 , \24040 );
nand \U$23699 ( \24042 , \23981 , \24041 );
nand \U$23700 ( \24043 , \23957 , \24042 );
nand \U$23701 ( \24044 , \23956 , \24043 );
not \U$23702 ( \24045 , \24044 );
xor \U$23703 ( \24046 , \23450 , \23487 );
xnor \U$23704 ( \24047 , \24046 , \23540 );
nand \U$23705 ( \24048 , \24045 , \24047 );
not \U$23706 ( \24049 , \24048 );
or \U$23707 ( \24050 , \23884 , \24049 );
not \U$23708 ( \24051 , \24047 );
nand \U$23709 ( \24052 , \24051 , \24044 );
nand \U$23710 ( \24053 , \24050 , \24052 );
not \U$23711 ( \24054 , \24053 );
xor \U$23712 ( \24055 , \23073 , \23075 );
xor \U$23713 ( \24056 , \24055 , \23078 );
not \U$23714 ( \24057 , \24056 );
xor \U$23715 ( \24058 , \22902 , \22912 );
xor \U$23716 ( \24059 , \24058 , \22922 );
xor \U$23717 ( \24060 , \22950 , \22939 );
and \U$23718 ( \24061 , \24060 , \22961 );
not \U$23719 ( \24062 , \24060 );
and \U$23720 ( \24063 , \24062 , \22962 );
nor \U$23721 ( \24064 , \24061 , \24063 );
or \U$23722 ( \24065 , \24059 , \24064 );
xor \U$23723 ( \24066 , \23412 , \23408 );
xnor \U$23724 ( \24067 , \24066 , \23439 );
nand \U$23725 ( \24068 , \24065 , \24067 );
nand \U$23726 ( \24069 , \24059 , \24064 );
nand \U$23727 ( \24070 , \24068 , \24069 );
not \U$23728 ( \24071 , \24070 );
nand \U$23729 ( \24072 , \24057 , \24071 );
not \U$23730 ( \24073 , \24072 );
or \U$23731 ( \24074 , \24054 , \24073 );
nand \U$23732 ( \24075 , \24056 , \24070 );
nand \U$23733 ( \24076 , \24074 , \24075 );
not \U$23734 ( \24077 , \24076 );
not \U$23735 ( \24078 , \24077 );
and \U$23736 ( \24079 , \23549 , \23561 );
not \U$23737 ( \24080 , \23549 );
and \U$23738 ( \24081 , \24080 , \23560 );
nor \U$23739 ( \24082 , \24079 , \24081 );
xor \U$23740 ( \24083 , \23715 , \24082 );
not \U$23741 ( \24084 , \24083 );
or \U$23742 ( \24085 , \24078 , \24084 );
xor \U$23743 ( \24086 , \23384 , \23393 );
xor \U$23744 ( \24087 , \24086 , \23405 );
not \U$23745 ( \24088 , \24087 );
xor \U$23746 ( \24089 , \23436 , \23433 );
xnor \U$23747 ( \24090 , \24089 , \23423 );
nand \U$23748 ( \24091 , \24088 , \24090 );
not \U$23749 ( \24092 , \24091 );
xor \U$23750 ( \24093 , \23491 , \23501 );
xor \U$23751 ( \24094 , \24093 , \23512 );
not \U$23752 ( \24095 , \16533 );
not \U$23753 ( \24096 , \23668 );
or \U$23754 ( \24097 , \24095 , \24096 );
not \U$23755 ( \24098 , RIbb2d9f0_61);
not \U$23756 ( \24099 , \3368 );
or \U$23757 ( \24100 , \24098 , \24099 );
nand \U$23758 ( \24101 , \3369 , \16254 );
nand \U$23759 ( \24102 , \24100 , \24101 );
nand \U$23760 ( \24103 , \24102 , \16541 );
nand \U$23761 ( \24104 , \24097 , \24103 );
xor \U$23762 ( \24105 , \24094 , \24104 );
not \U$23763 ( \24106 , \12284 );
not \U$23764 ( \24107 , \23778 );
or \U$23765 ( \24108 , \24106 , \24107 );
not \U$23766 ( \24109 , RIbb2df90_49);
not \U$23767 ( \24110 , \20951 );
or \U$23768 ( \24111 , \24109 , \24110 );
nand \U$23769 ( \24112 , \12096 , \12278 );
nand \U$23770 ( \24113 , \24111 , \24112 );
nand \U$23771 ( \24114 , \24113 , \12167 );
nand \U$23772 ( \24115 , \24108 , \24114 );
and \U$23773 ( \24116 , \24105 , \24115 );
and \U$23774 ( \24117 , \24094 , \24104 );
or \U$23775 ( \24118 , \24116 , \24117 );
not \U$23776 ( \24119 , \24118 );
or \U$23777 ( \24120 , \24092 , \24119 );
or \U$23778 ( \24121 , \24088 , \24090 );
nand \U$23779 ( \24122 , \24120 , \24121 );
not \U$23780 ( \24123 , \8362 );
not \U$23781 ( \24124 , RIbb2e350_41);
not \U$23782 ( \24125 , \13731 );
or \U$23783 ( \24126 , \24124 , \24125 );
nand \U$23784 ( \24127 , \3274 , \9402 );
nand \U$23785 ( \24128 , \24126 , \24127 );
not \U$23786 ( \24129 , \24128 );
or \U$23787 ( \24130 , \24123 , \24129 );
nand \U$23788 ( \24131 , \23578 , \8354 );
nand \U$23789 ( \24132 , \24130 , \24131 );
not \U$23790 ( \24133 , \24132 );
not \U$23791 ( \24134 , \24133 );
not \U$23792 ( \24135 , \9099 );
not \U$23793 ( \24136 , \23683 );
or \U$23794 ( \24137 , \24135 , \24136 );
not \U$23795 ( \24138 , RIbb2e260_43);
not \U$23796 ( \24139 , \22894 );
or \U$23797 ( \24140 , \24138 , \24139 );
nand \U$23798 ( \24141 , \4020 , \10444 );
nand \U$23799 ( \24142 , \24140 , \24141 );
nand \U$23800 ( \24143 , \24142 , \9098 );
nand \U$23801 ( \24144 , \24137 , \24143 );
not \U$23802 ( \24145 , \24144 );
not \U$23803 ( \24146 , \24145 );
or \U$23804 ( \24147 , \24134 , \24146 );
not \U$23805 ( \24148 , \14613 );
not \U$23806 ( \24149 , RIbb2dcc0_55);
not \U$23807 ( \24150 , \13619 );
or \U$23808 ( \24151 , \24149 , \24150 );
nand \U$23809 ( \24152 , \1386 , \17959 );
nand \U$23810 ( \24153 , \24151 , \24152 );
not \U$23811 ( \24154 , \24153 );
or \U$23812 ( \24155 , \24148 , \24154 );
nand \U$23813 ( \24156 , \23694 , \15181 );
nand \U$23814 ( \24157 , \24155 , \24156 );
nand \U$23815 ( \24158 , \24147 , \24157 );
nand \U$23816 ( \24159 , \24132 , \24144 );
nand \U$23817 ( \24160 , \24158 , \24159 );
not \U$23818 ( \24161 , \24160 );
not \U$23819 ( \24162 , \12690 );
and \U$23820 ( \24163 , RIbb2dea0_51, \9983 );
not \U$23821 ( \24164 , RIbb2dea0_51);
and \U$23822 ( \24165 , \24164 , \2114 );
or \U$23823 ( \24166 , \24163 , \24165 );
not \U$23824 ( \24167 , \24166 );
or \U$23825 ( \24168 , \24162 , \24167 );
nand \U$23826 ( \24169 , \23625 , \12692 );
nand \U$23827 ( \24170 , \24168 , \24169 );
not \U$23828 ( \24171 , \24170 );
not \U$23829 ( \24172 , \8450 );
not \U$23830 ( \24173 , \23584 );
or \U$23831 ( \24174 , \24172 , \24173 );
and \U$23832 ( \24175 , RIbb2e440_39, \13756 );
not \U$23833 ( \24176 , RIbb2e440_39);
and \U$23834 ( \24177 , \24176 , \4324 );
or \U$23835 ( \24178 , \24175 , \24177 );
nand \U$23836 ( \24179 , \24178 , \7102 );
nand \U$23837 ( \24180 , \24174 , \24179 );
not \U$23838 ( \24181 , \24180 );
not \U$23839 ( \24182 , \24181 );
not \U$23840 ( \24183 , \24182 );
or \U$23841 ( \24184 , \24171 , \24183 );
not \U$23842 ( \24185 , \24170 );
not \U$23843 ( \24186 , \24185 );
not \U$23844 ( \24187 , \24181 );
or \U$23845 ( \24188 , \24186 , \24187 );
not \U$23846 ( \24189 , \14929 );
not \U$23847 ( \24190 , \23593 );
or \U$23848 ( \24191 , \24189 , \24190 );
not \U$23849 ( \24192 , RIbb2ddb0_53);
not \U$23850 ( \24193 , \19733 );
or \U$23851 ( \24194 , \24192 , \24193 );
nand \U$23852 ( \24195 , \1337 , \12681 );
nand \U$23853 ( \24196 , \24194 , \24195 );
nand \U$23854 ( \24197 , \24196 , \13467 );
nand \U$23855 ( \24198 , \24191 , \24197 );
nand \U$23856 ( \24199 , \24188 , \24198 );
nand \U$23857 ( \24200 , \24184 , \24199 );
not \U$23858 ( \24201 , \24200 );
or \U$23859 ( \24202 , \24161 , \24201 );
or \U$23860 ( \24203 , \24160 , \24200 );
xor \U$23861 ( \24204 , \23657 , \23646 );
xnor \U$23862 ( \24205 , \24204 , \23670 );
not \U$23863 ( \24206 , \24205 );
nand \U$23864 ( \24207 , \24203 , \24206 );
nand \U$23865 ( \24208 , \24202 , \24207 );
xor \U$23866 ( \24209 , \24122 , \24208 );
xor \U$23867 ( \24210 , \23748 , \23784 );
xor \U$23868 ( \24211 , \24210 , \23787 );
and \U$23869 ( \24212 , \24209 , \24211 );
and \U$23870 ( \24213 , \24122 , \24208 );
or \U$23871 ( \24214 , \24212 , \24213 );
xor \U$23872 ( \24215 , \23446 , \23547 );
xnor \U$23873 ( \24216 , \24215 , \23544 );
nor \U$23874 ( \24217 , \24214 , \24216 );
xor \U$23875 ( \24218 , \23565 , \23713 );
xnor \U$23876 ( \24219 , \24218 , \23632 );
or \U$23877 ( \24220 , \24217 , \24219 );
nand \U$23878 ( \24221 , \24214 , \24216 );
nand \U$23879 ( \24222 , \24220 , \24221 );
nand \U$23880 ( \24223 , \24085 , \24222 );
or \U$23881 ( \24224 , \24083 , \24077 );
nand \U$23882 ( \24225 , \24223 , \24224 );
xor \U$23883 ( \24226 , \23720 , \23722 );
xor \U$23884 ( \24227 , \24226 , \23796 );
xor \U$23885 ( \24228 , \24225 , \24227 );
not \U$23886 ( \24229 , \23067 );
not \U$23887 ( \24230 , \24229 );
not \U$23888 ( \24231 , \23055 );
or \U$23889 ( \24232 , \24230 , \24231 );
nand \U$23890 ( \24233 , \23067 , \23054 );
nand \U$23891 ( \24234 , \24232 , \24233 );
and \U$23892 ( \24235 , \24234 , \23081 );
not \U$23893 ( \24236 , \24234 );
not \U$23894 ( \24237 , \23081 );
and \U$23895 ( \24238 , \24236 , \24237 );
nor \U$23896 ( \24239 , \24235 , \24238 );
xor \U$23897 ( \24240 , \23330 , \23332 );
xor \U$23898 ( \24241 , \24240 , \23343 );
xor \U$23899 ( \24242 , \24239 , \24241 );
xor \U$23900 ( \24243 , \22881 , \22885 );
xnor \U$23901 ( \24244 , \24243 , \22925 );
not \U$23902 ( \24245 , \998 );
not \U$23903 ( \24246 , \23201 );
or \U$23904 ( \24247 , \24245 , \24246 );
nand \U$23905 ( \24248 , \915 , \24012 );
nand \U$23906 ( \24249 , \24247 , \24248 );
and \U$23907 ( \24250 , \19064 , \1737 );
not \U$23908 ( \24251 , \1569 );
not \U$23909 ( \24252 , \23499 );
or \U$23910 ( \24253 , \24251 , \24252 );
nand \U$23911 ( \24254 , \23988 , \1532 );
nand \U$23912 ( \24255 , \24253 , \24254 );
xor \U$23913 ( \24256 , \24250 , \24255 );
not \U$23914 ( \24257 , \1011 );
not \U$23915 ( \24258 , RIbb2f160_11);
not \U$23916 ( \24259 , \17755 );
or \U$23917 ( \24260 , \24258 , \24259 );
nand \U$23918 ( \24261 , \16703 , \1043 );
nand \U$23919 ( \24262 , \24260 , \24261 );
not \U$23920 ( \24263 , \24262 );
or \U$23921 ( \24264 , \24257 , \24263 );
nand \U$23922 ( \24265 , \23510 , \1077 );
nand \U$23923 ( \24266 , \24264 , \24265 );
and \U$23924 ( \24267 , \24256 , \24266 );
and \U$23925 ( \24268 , \24250 , \24255 );
or \U$23926 ( \24269 , \24267 , \24268 );
xor \U$23927 ( \24270 , \24249 , \24269 );
not \U$23928 ( \24271 , \853 );
not \U$23929 ( \24272 , RIbb2eda0_19);
not \U$23930 ( \24273 , \13986 );
or \U$23931 ( \24274 , \24272 , \24273 );
nand \U$23932 ( \24275 , \13545 , \5277 );
nand \U$23933 ( \24276 , \24274 , \24275 );
not \U$23934 ( \24277 , \24276 );
or \U$23935 ( \24278 , \24271 , \24277 );
nand \U$23936 ( \24279 , \23431 , \854 );
nand \U$23937 ( \24280 , \24278 , \24279 );
and \U$23938 ( \24281 , \24270 , \24280 );
and \U$23939 ( \24282 , \24249 , \24269 );
or \U$23940 ( \24283 , \24281 , \24282 );
not \U$23941 ( \24284 , \2078 );
not \U$23942 ( \24285 , \23421 );
or \U$23943 ( \24286 , \24284 , \24285 );
not \U$23944 ( \24287 , RIbb2ecb0_21);
not \U$23945 ( \24288 , \13809 );
or \U$23946 ( \24289 , \24287 , \24288 );
not \U$23947 ( \24290 , \12346 );
not \U$23948 ( \24291 , \24290 );
nand \U$23949 ( \24292 , \24291 , \5481 );
nand \U$23950 ( \24293 , \24289 , \24292 );
nand \U$23951 ( \24294 , \24293 , \2077 );
nand \U$23952 ( \24295 , \24286 , \24294 );
not \U$23953 ( \24296 , \24295 );
not \U$23954 ( \24297 , \24296 );
not \U$23955 ( \24298 , \836 );
not \U$23956 ( \24299 , \23380 );
or \U$23957 ( \24300 , \24298 , \24299 );
not \U$23958 ( \24301 , RIbb2ee90_17);
not \U$23959 ( \24302 , \16309 );
or \U$23960 ( \24303 , \24301 , \24302 );
nand \U$23961 ( \24304 , \14526 , \822 );
nand \U$23962 ( \24305 , \24303 , \24304 );
nand \U$23963 ( \24306 , \831 , \24305 );
nand \U$23964 ( \24307 , \24300 , \24306 );
not \U$23965 ( \24308 , \24307 );
not \U$23966 ( \24309 , \24308 );
or \U$23967 ( \24310 , \24297 , \24309 );
not \U$23968 ( \24311 , \1517 );
not \U$23969 ( \24312 , \23389 );
or \U$23970 ( \24313 , \24311 , \24312 );
nand \U$23971 ( \24314 , \1445 , \24029 );
nand \U$23972 ( \24315 , \24313 , \24314 );
nand \U$23973 ( \24316 , \24310 , \24315 );
nand \U$23974 ( \24317 , \24295 , \24307 );
nand \U$23975 ( \24318 , \24316 , \24317 );
xor \U$23976 ( \24319 , \24283 , \24318 );
not \U$23977 ( \24320 , \16271 );
and \U$23978 ( \24321 , RIbb2dae0_59, \3238 );
not \U$23979 ( \24322 , RIbb2dae0_59);
and \U$23980 ( \24323 , \24322 , \8856 );
or \U$23981 ( \24324 , \24321 , \24323 );
not \U$23982 ( \24325 , \24324 );
or \U$23983 ( \24326 , \24320 , \24325 );
nand \U$23984 ( \24327 , \23026 , \17470 );
nand \U$23985 ( \24328 , \24326 , \24327 );
and \U$23986 ( \24329 , \24319 , \24328 );
and \U$23987 ( \24330 , \24283 , \24318 );
or \U$23988 ( \24331 , \24329 , \24330 );
xor \U$23989 ( \24332 , \23303 , \23313 );
xor \U$23990 ( \24333 , \24332 , \23324 );
xor \U$23991 ( \24334 , \24331 , \24333 );
xor \U$23992 ( \24335 , \23010 , \23020 );
xor \U$23993 ( \24336 , \24335 , \23030 );
and \U$23994 ( \24337 , \24334 , \24336 );
and \U$23995 ( \24338 , \24331 , \24333 );
or \U$23996 ( \24339 , \24337 , \24338 );
xor \U$23997 ( \24340 , \24244 , \24339 );
xor \U$23998 ( \24341 , \22965 , \23000 );
xor \U$23999 ( \24342 , \24341 , \23033 );
and \U$24000 ( \24343 , \24340 , \24342 );
and \U$24001 ( \24344 , \24244 , \24339 );
or \U$24002 ( \24345 , \24343 , \24344 );
xor \U$24003 ( \24346 , \24242 , \24345 );
xor \U$24004 ( \24347 , \23725 , \23736 );
xor \U$24005 ( \24348 , \24347 , \23793 );
or \U$24006 ( \24349 , \24346 , \24348 );
xor \U$24007 ( \24350 , \23674 , \23676 );
xor \U$24008 ( \24351 , \24350 , \23710 );
xor \U$24009 ( \24352 , \23569 , \23630 );
xor \U$24010 ( \24353 , \24352 , \23600 );
xor \U$24011 ( \24354 , \24351 , \24353 );
xor \U$24012 ( \24355 , \23605 , \23615 );
xor \U$24013 ( \24356 , \24355 , \23627 );
xor \U$24014 ( \24357 , \24250 , \24255 );
xor \U$24015 ( \24358 , \24357 , \24266 );
not \U$24016 ( \24359 , \2078 );
not \U$24017 ( \24360 , \24293 );
or \U$24018 ( \24361 , \24359 , \24360 );
not \U$24019 ( \24362 , RIbb2ecb0_21);
not \U$24020 ( \24363 , \14624 );
or \U$24021 ( \24364 , \24362 , \24363 );
nand \U$24022 ( \24365 , \13210 , \849 );
nand \U$24023 ( \24366 , \24364 , \24365 );
nand \U$24024 ( \24367 , \24366 , \2077 );
nand \U$24025 ( \24368 , \24361 , \24367 );
xor \U$24026 ( \24369 , \24358 , \24368 );
not \U$24027 ( \24370 , \24276 );
not \U$24028 ( \24371 , \854 );
or \U$24029 ( \24372 , \24370 , \24371 );
not \U$24030 ( \24373 , RIbb2eda0_19);
not \U$24031 ( \24374 , \16317 );
or \U$24032 ( \24375 , \24373 , \24374 );
nand \U$24033 ( \24376 , \13977 , \1776 );
nand \U$24034 ( \24377 , \24375 , \24376 );
nand \U$24035 ( \24378 , \24377 , \853 );
nand \U$24036 ( \24379 , \24372 , \24378 );
and \U$24037 ( \24380 , \24369 , \24379 );
and \U$24038 ( \24381 , \24358 , \24368 );
or \U$24039 ( \24382 , \24380 , \24381 );
not \U$24040 ( \24383 , RIbb2d888_64);
not \U$24041 ( \24384 , \23611 );
or \U$24042 ( \24385 , \24383 , \24384 );
not \U$24043 ( \24386 , RIbb2d900_63);
not \U$24044 ( \24387 , \15629 );
or \U$24045 ( \24388 , \24386 , \24387 );
nand \U$24046 ( \24389 , \1548 , \17270 );
nand \U$24047 ( \24390 , \24388 , \24389 );
nand \U$24048 ( \24391 , \24390 , \17275 );
nand \U$24049 ( \24392 , \24385 , \24391 );
xor \U$24050 ( \24393 , \24382 , \24392 );
not \U$24051 ( \24394 , \17470 );
not \U$24052 ( \24395 , \24324 );
or \U$24053 ( \24396 , \24394 , \24395 );
and \U$24054 ( \24397 , RIbb2dae0_59, \7423 );
not \U$24055 ( \24398 , RIbb2dae0_59);
not \U$24056 ( \24399 , \7423 );
and \U$24057 ( \24400 , \24398 , \24399 );
or \U$24058 ( \24401 , \24397 , \24400 );
nand \U$24059 ( \24402 , \24401 , \16271 );
nand \U$24060 ( \24403 , \24396 , \24402 );
and \U$24061 ( \24404 , \24393 , \24403 );
and \U$24062 ( \24405 , \24382 , \24392 );
or \U$24063 ( \24406 , \24404 , \24405 );
xor \U$24064 ( \24407 , \24356 , \24406 );
xor \U$24065 ( \24408 , \23782 , \23769 );
xor \U$24066 ( \24409 , \24408 , \23758 );
and \U$24067 ( \24410 , \24407 , \24409 );
and \U$24068 ( \24411 , \24356 , \24406 );
or \U$24069 ( \24412 , \24410 , \24411 );
and \U$24070 ( \24413 , \24354 , \24412 );
and \U$24071 ( \24414 , \24351 , \24353 );
or \U$24072 ( \24415 , \24413 , \24414 );
xor \U$24073 ( \24416 , \23743 , \23745 );
xor \U$24074 ( \24417 , \24416 , \23790 );
xor \U$24075 ( \24418 , \24415 , \24417 );
xor \U$24076 ( \24419 , \23687 , \23696 );
xor \U$24077 ( \24420 , \24419 , \23707 );
xor \U$24078 ( \24421 , \23580 , \23586 );
xor \U$24079 ( \24422 , \24421 , \23597 );
xor \U$24080 ( \24423 , \24420 , \24422 );
xor \U$24081 ( \24424 , \24249 , \24269 );
xor \U$24082 ( \24425 , \24424 , \24280 );
not \U$24083 ( \24426 , \3382 );
not \U$24084 ( \24427 , \23928 );
or \U$24085 ( \24428 , \24426 , \24427 );
not \U$24086 ( \24429 , RIbb2ebc0_23);
not \U$24087 ( \24430 , \12321 );
not \U$24088 ( \24431 , \24430 );
or \U$24089 ( \24432 , \24429 , \24431 );
nand \U$24090 ( \24433 , \12321 , \3388 );
nand \U$24091 ( \24434 , \24432 , \24433 );
nand \U$24092 ( \24435 , \24434 , \3406 );
nand \U$24093 ( \24436 , \24428 , \24435 );
not \U$24094 ( \24437 , \24436 );
not \U$24095 ( \24438 , \3613 );
not \U$24096 ( \24439 , \23964 );
or \U$24097 ( \24440 , \24438 , \24439 );
and \U$24098 ( \24441 , \8630 , \4096 );
not \U$24099 ( \24442 , \8630 );
and \U$24100 ( \24443 , \24442 , RIbb2e800_31);
or \U$24101 ( \24444 , \24441 , \24443 );
nand \U$24102 ( \24445 , \24444 , \2939 );
nand \U$24103 ( \24446 , \24440 , \24445 );
not \U$24104 ( \24447 , \24446 );
nand \U$24105 ( \24448 , \24437 , \24447 );
not \U$24106 ( \24449 , \24448 );
not \U$24107 ( \24450 , \836 );
not \U$24108 ( \24451 , \24305 );
or \U$24109 ( \24452 , \24450 , \24451 );
not \U$24110 ( \24453 , RIbb2ee90_17);
not \U$24111 ( \24454 , \15031 );
or \U$24112 ( \24455 , \24453 , \24454 );
nand \U$24113 ( \24456 , \15470 , \2240 );
nand \U$24114 ( \24457 , \24455 , \24456 );
nand \U$24115 ( \24458 , \24457 , \831 );
nand \U$24116 ( \24459 , \24452 , \24458 );
not \U$24117 ( \24460 , \24459 );
or \U$24118 ( \24461 , \24449 , \24460 );
nand \U$24119 ( \24462 , \24446 , \24436 );
nand \U$24120 ( \24463 , \24461 , \24462 );
xor \U$24121 ( \24464 , \24425 , \24463 );
not \U$24122 ( \24465 , \2925 );
not \U$24123 ( \24466 , \23977 );
or \U$24124 ( \24467 , \24465 , \24466 );
not \U$24125 ( \24468 , RIbb2e8f0_29);
not \U$24126 ( \24469 , \13498 );
or \U$24127 ( \24470 , \24468 , \24469 );
nand \U$24128 ( \24471 , \9840 , \3800 );
nand \U$24129 ( \24472 , \24470 , \24471 );
nand \U$24130 ( \24473 , \24472 , \2921 );
nand \U$24131 ( \24474 , \24467 , \24473 );
not \U$24132 ( \24475 , \2963 );
not \U$24133 ( \24476 , \23912 );
or \U$24134 ( \24477 , \24475 , \24476 );
not \U$24135 ( \24478 , RIbb2ead0_25);
not \U$24136 ( \24479 , \11579 );
or \U$24137 ( \24480 , \24478 , \24479 );
not \U$24138 ( \24481 , RIbb2ead0_25);
nand \U$24139 ( \24482 , \24481 , \11578 );
nand \U$24140 ( \24483 , \24480 , \24482 );
nand \U$24141 ( \24484 , \24483 , \2980 );
nand \U$24142 ( \24485 , \24477 , \24484 );
xor \U$24143 ( \24486 , \24474 , \24485 );
not \U$24144 ( \24487 , \3465 );
not \U$24145 ( \24488 , \23949 );
or \U$24146 ( \24489 , \24487 , \24488 );
not \U$24147 ( \24490 , RIbb2e9e0_27);
not \U$24148 ( \24491 , \12249 );
or \U$24149 ( \24492 , \24490 , \24491 );
nand \U$24150 ( \24493 , \13526 , \3462 );
nand \U$24151 ( \24494 , \24492 , \24493 );
nand \U$24152 ( \24495 , \24494 , \3445 );
nand \U$24153 ( \24496 , \24489 , \24495 );
and \U$24154 ( \24497 , \24486 , \24496 );
and \U$24155 ( \24498 , \24474 , \24485 );
or \U$24156 ( \24499 , \24497 , \24498 );
and \U$24157 ( \24500 , \24464 , \24499 );
and \U$24158 ( \24501 , \24425 , \24463 );
or \U$24159 ( \24502 , \24500 , \24501 );
and \U$24160 ( \24503 , \24423 , \24502 );
and \U$24161 ( \24504 , \24420 , \24422 );
or \U$24162 ( \24505 , \24503 , \24504 );
xor \U$24163 ( \24506 , \24331 , \24333 );
xor \U$24164 ( \24507 , \24506 , \24336 );
xor \U$24165 ( \24508 , \24505 , \24507 );
xor \U$24166 ( \24509 , \24064 , \24059 );
xor \U$24167 ( \24510 , \24509 , \24067 );
and \U$24168 ( \24511 , \24508 , \24510 );
and \U$24169 ( \24512 , \24505 , \24507 );
or \U$24170 ( \24513 , \24511 , \24512 );
and \U$24171 ( \24514 , \24418 , \24513 );
and \U$24172 ( \24515 , \24415 , \24417 );
or \U$24173 ( \24516 , \24514 , \24515 );
nand \U$24174 ( \24517 , \24349 , \24516 );
nand \U$24175 ( \24518 , \24346 , \24348 );
nand \U$24176 ( \24519 , \24517 , \24518 );
and \U$24177 ( \24520 , \24228 , \24519 );
and \U$24178 ( \24521 , \24225 , \24227 );
or \U$24179 ( \24522 , \24520 , \24521 );
xor \U$24180 ( \24523 , \24239 , \24241 );
and \U$24181 ( \24524 , \24523 , \24345 );
and \U$24182 ( \24525 , \24239 , \24241 );
or \U$24183 ( \24526 , \24524 , \24525 );
xor \U$24184 ( \24527 , \23083 , \23051 );
buf \U$24185 ( \24528 , \23088 );
and \U$24186 ( \24529 , \24527 , \24528 );
not \U$24187 ( \24530 , \24527 );
not \U$24188 ( \24531 , \24528 );
and \U$24189 ( \24532 , \24530 , \24531 );
nor \U$24190 ( \24533 , \24529 , \24532 );
buf \U$24191 ( \24534 , \24533 );
or \U$24192 ( \24535 , \24526 , \24534 );
xor \U$24193 ( \24536 , \23361 , \23362 );
xor \U$24194 ( \24537 , \24536 , \23359 );
nand \U$24195 ( \24538 , \24535 , \24537 );
nand \U$24196 ( \24539 , \24526 , \24534 );
nand \U$24197 ( \24540 , \24538 , \24539 );
or \U$24198 ( \24541 , \24522 , \24540 );
not \U$24199 ( \24542 , \24541 );
or \U$24200 ( \24543 , \23844 , \24542 );
nand \U$24201 ( \24544 , \24522 , \24540 );
nand \U$24202 ( \24545 , \24543 , \24544 );
nand \U$24203 ( \24546 , \23833 , \24545 );
nand \U$24204 ( \24547 , \23831 , \24546 );
not \U$24205 ( \24548 , \23829 );
not \U$24206 ( \24549 , \23818 );
nand \U$24207 ( \24550 , \24548 , \24549 );
nand \U$24208 ( \24551 , \24547 , \24550 );
xor \U$24209 ( \24552 , \22658 , \22864 );
xor \U$24210 ( \24553 , \24552 , \22661 );
xor \U$24211 ( \24554 , \23821 , \23823 );
and \U$24212 ( \24555 , \24554 , \23828 );
and \U$24213 ( \24556 , \23821 , \23823 );
or \U$24214 ( \24557 , \24555 , \24556 );
nor \U$24215 ( \24558 , \24553 , \24557 );
or \U$24216 ( \24559 , \24551 , \24558 );
nand \U$24217 ( \24560 , \24553 , \24557 );
nand \U$24218 ( \24561 , \24559 , \24560 );
not \U$24219 ( \24562 , \24561 );
or \U$24220 ( \24563 , \22871 , \24562 );
not \U$24221 ( \24564 , \22656 );
not \U$24222 ( \24565 , \22869 );
nand \U$24223 ( \24566 , \24564 , \24565 );
nand \U$24224 ( \24567 , \24563 , \24566 );
not \U$24225 ( \24568 , \24567 );
or \U$24226 ( \24569 , \22654 , \24568 );
buf \U$24227 ( \24570 , \22647 );
nand \U$24228 ( \24571 , \24570 , \22651 );
nand \U$24229 ( \24572 , \24569 , \24571 );
nor \U$24230 ( \24573 , \21547 , \20633 );
not \U$24231 ( \24574 , \24573 );
not \U$24232 ( \24575 , \20630 );
or \U$24233 ( \24576 , \24574 , \24575 );
not \U$24234 ( \24577 , \19950 );
nand \U$24235 ( \24578 , \24577 , \20628 );
nand \U$24236 ( \24579 , \24576 , \24578 );
not \U$24237 ( \24580 , \22124 );
nand \U$24238 ( \24581 , \24579 , \24580 );
buf \U$24239 ( \24582 , \22123 );
nand \U$24240 ( \24583 , \24582 , \21558 );
and \U$24241 ( \24584 , \24581 , \24583 );
not \U$24242 ( \24585 , \22652 );
not \U$24243 ( \24586 , \24585 );
nor \U$24244 ( \24587 , \24584 , \24586 );
nor \U$24245 ( \24588 , \24572 , \24587 );
xor \U$24246 ( \24589 , \22293 , \22397 );
and \U$24247 ( \24590 , \24589 , \22402 );
and \U$24248 ( \24591 , \22293 , \22397 );
or \U$24249 ( \24592 , \24590 , \24591 );
not \U$24250 ( \24593 , \13295 );
not \U$24251 ( \24594 , \22301 );
or \U$24252 ( \24595 , \24593 , \24594 );
nand \U$24253 ( \24596 , \15665 , \12169 );
nand \U$24254 ( \24597 , \24595 , \24596 );
not \U$24255 ( \24598 , \6242 );
not \U$24256 ( \24599 , \15647 );
or \U$24257 ( \24600 , \24598 , \24599 );
nand \U$24258 ( \24601 , \22321 , \6251 );
nand \U$24259 ( \24602 , \24600 , \24601 );
not \U$24260 ( \24603 , \24602 );
and \U$24261 ( \24604 , \24597 , \24603 );
not \U$24262 ( \24605 , \24597 );
and \U$24263 ( \24606 , \24605 , \24602 );
or \U$24264 ( \24607 , \24604 , \24606 );
not \U$24265 ( \24608 , \7103 );
not \U$24266 ( \24609 , \22308 );
or \U$24267 ( \24610 , \24608 , \24609 );
nand \U$24268 ( \24611 , \15674 , \8450 );
nand \U$24269 ( \24612 , \24610 , \24611 );
not \U$24270 ( \24613 , \24612 );
and \U$24271 ( \24614 , \24607 , \24613 );
not \U$24272 ( \24615 , \24607 );
and \U$24273 ( \24616 , \24615 , \24612 );
nor \U$24274 ( \24617 , \24614 , \24616 );
not \U$24275 ( \24618 , \24617 );
not \U$24276 ( \24619 , \14613 );
not \U$24277 ( \24620 , \22222 );
or \U$24278 ( \24621 , \24619 , \24620 );
nand \U$24279 ( \24622 , \15178 , \15181 );
nand \U$24280 ( \24623 , \24621 , \24622 );
not \U$24281 ( \24624 , \12774 );
not \U$24282 ( \24625 , \22231 );
or \U$24283 ( \24626 , \24624 , \24625 );
nand \U$24284 ( \24627 , \15560 , \12692 );
nand \U$24285 ( \24628 , \24626 , \24627 );
xor \U$24286 ( \24629 , \24623 , \24628 );
not \U$24287 ( \24630 , \8362 );
not \U$24288 ( \24631 , \22244 );
or \U$24289 ( \24632 , \24630 , \24631 );
nand \U$24290 ( \24633 , \15585 , \8354 );
nand \U$24291 ( \24634 , \24632 , \24633 );
xor \U$24292 ( \24635 , \24629 , \24634 );
not \U$24293 ( \24636 , \24635 );
or \U$24294 ( \24637 , \24618 , \24636 );
or \U$24295 ( \24638 , \24617 , \24635 );
nand \U$24296 ( \24639 , \24637 , \24638 );
not \U$24297 ( \24640 , \9098 );
not \U$24298 ( \24641 , \22393 );
or \U$24299 ( \24642 , \24640 , \24641 );
nand \U$24300 ( \24643 , \15433 , \9099 );
nand \U$24301 ( \24644 , \24642 , \24643 );
not \U$24302 ( \24645 , \3445 );
not \U$24303 ( \24646 , \22381 );
or \U$24304 ( \24647 , \24645 , \24646 );
nand \U$24305 ( \24648 , \15446 , \3465 );
nand \U$24306 ( \24649 , \24647 , \24648 );
xor \U$24307 ( \24650 , \24644 , \24649 );
not \U$24308 ( \24651 , \2980 );
not \U$24309 ( \24652 , \22369 );
or \U$24310 ( \24653 , \24651 , \24652 );
not \U$24311 ( \24654 , \16353 );
nand \U$24312 ( \24655 , \24654 , \15609 );
nand \U$24313 ( \24656 , \24653 , \24655 );
xnor \U$24314 ( \24657 , \24650 , \24656 );
and \U$24315 ( \24658 , \24639 , \24657 );
not \U$24316 ( \24659 , \24639 );
not \U$24317 ( \24660 , \24657 );
and \U$24318 ( \24661 , \24659 , \24660 );
nor \U$24319 ( \24662 , \24658 , \24661 );
not \U$24320 ( \24663 , \24662 );
not \U$24321 ( \24664 , \24663 );
not \U$24322 ( \24665 , \22323 );
not \U$24323 ( \24666 , \22313 );
or \U$24324 ( \24667 , \24665 , \24666 );
nand \U$24325 ( \24668 , \24667 , \22303 );
nand \U$24326 ( \24669 , \22326 , \22312 );
nand \U$24327 ( \24670 , \24668 , \24669 );
not \U$24328 ( \24671 , \11176 );
not \U$24329 ( \24672 , \22359 );
or \U$24330 ( \24673 , \24671 , \24672 );
nand \U$24331 ( \24674 , \15634 , \11177 );
nand \U$24332 ( \24675 , \24673 , \24674 );
not \U$24333 ( \24676 , \4712 );
not \U$24334 ( \24677 , \22347 );
or \U$24335 ( \24678 , \24676 , \24677 );
nand \U$24336 ( \24679 , \15622 , \5845 );
nand \U$24337 ( \24680 , \24678 , \24679 );
xor \U$24338 ( \24681 , \24675 , \24680 );
not \U$24339 ( \24682 , \13467 );
not \U$24340 ( \24683 , \22336 );
or \U$24341 ( \24684 , \24682 , \24683 );
nand \U$24342 ( \24685 , \15685 , \14930 );
nand \U$24343 ( \24686 , \24684 , \24685 );
xor \U$24344 ( \24687 , \24681 , \24686 );
xor \U$24345 ( \24688 , \24670 , \24687 );
not \U$24346 ( \24689 , \2941 );
not \U$24347 ( \24690 , \15402 );
or \U$24348 ( \24691 , \24689 , \24690 );
nand \U$24349 ( \24692 , \22284 , \2939 );
nand \U$24350 ( \24693 , \24691 , \24692 );
not \U$24351 ( \24694 , \10599 );
not \U$24352 ( \24695 , \22256 );
or \U$24353 ( \24696 , \24694 , \24695 );
nand \U$24354 ( \24697 , \15539 , \10119 );
nand \U$24355 ( \24698 , \24696 , \24697 );
xor \U$24356 ( \24699 , \24693 , \24698 );
not \U$24357 ( \24700 , \4791 );
not \U$24358 ( \24701 , \15549 );
or \U$24359 ( \24702 , \24700 , \24701 );
nand \U$24360 ( \24703 , \22268 , \3887 );
nand \U$24361 ( \24704 , \24702 , \24703 );
xor \U$24362 ( \24705 , \24699 , \24704 );
xor \U$24363 ( \24706 , \24688 , \24705 );
not \U$24364 ( \24707 , \24706 );
not \U$24365 ( \24708 , \24707 );
or \U$24366 ( \24709 , \24664 , \24708 );
nand \U$24367 ( \24710 , \24662 , \24706 );
nand \U$24368 ( \24711 , \24709 , \24710 );
xor \U$24369 ( \24712 , \22445 , \22452 );
and \U$24370 ( \24713 , \24712 , \22457 );
and \U$24371 ( \24714 , \22445 , \22452 );
or \U$24372 ( \24715 , \24713 , \24714 );
and \U$24373 ( \24716 , \24711 , \24715 );
not \U$24374 ( \24717 , \24711 );
not \U$24375 ( \24718 , \24715 );
and \U$24376 ( \24719 , \24717 , \24718 );
nor \U$24377 ( \24720 , \24716 , \24719 );
xor \U$24378 ( \24721 , \15826 , \15836 );
xor \U$24379 ( \24722 , \24721 , \15847 );
not \U$24380 ( \24723 , \832 );
not \U$24381 ( \24724 , \15778 );
or \U$24382 ( \24725 , \24723 , \24724 );
nand \U$24383 ( \24726 , \24725 , \15781 );
xor \U$24384 ( \24727 , \15805 , \24726 );
xor \U$24385 ( \24728 , \24727 , \15792 );
xor \U$24386 ( \24729 , \24722 , \24728 );
not \U$24387 ( \24730 , \916 );
not \U$24388 ( \24731 , \22584 );
or \U$24389 ( \24732 , \24730 , \24731 );
nand \U$24390 ( \24733 , \15130 , \998 );
nand \U$24391 ( \24734 , \24732 , \24733 );
not \U$24392 ( \24735 , \1011 );
not \U$24393 ( \24736 , \22568 );
or \U$24394 ( \24737 , \24735 , \24736 );
nand \U$24395 ( \24738 , \15109 , \1077 );
nand \U$24396 ( \24739 , \24737 , \24738 );
xor \U$24397 ( \24740 , \24734 , \24739 );
not \U$24398 ( \24741 , \1570 );
not \U$24399 ( \24742 , \15192 );
or \U$24400 ( \24743 , \24741 , \24742 );
nand \U$24401 ( \24744 , \22557 , \1533 );
nand \U$24402 ( \24745 , \24743 , \24744 );
and \U$24403 ( \24746 , \24740 , \24745 );
not \U$24404 ( \24747 , \24740 );
not \U$24405 ( \24748 , \24745 );
and \U$24406 ( \24749 , \24747 , \24748 );
nor \U$24407 ( \24750 , \24746 , \24749 );
xor \U$24408 ( \24751 , \24729 , \24750 );
not \U$24409 ( \24752 , \22247 );
not \U$24410 ( \24753 , \22291 );
or \U$24411 ( \24754 , \24752 , \24753 );
nand \U$24412 ( \24755 , \24754 , \22215 );
not \U$24413 ( \24756 , \22247 );
nand \U$24414 ( \24757 , \24756 , \22292 );
nand \U$24415 ( \24758 , \24755 , \24757 );
xor \U$24416 ( \24759 , \24751 , \24758 );
or \U$24417 ( \24760 , \22235 , \22246 );
nand \U$24418 ( \24761 , \24760 , \22226 );
nand \U$24419 ( \24762 , \22235 , \22246 );
nand \U$24420 ( \24763 , \24761 , \24762 );
or \U$24421 ( \24764 , \22349 , \22361 );
nand \U$24422 ( \24765 , \24764 , \22338 );
nand \U$24423 ( \24766 , \22349 , \22361 );
nand \U$24424 ( \24767 , \24765 , \24766 );
xor \U$24425 ( \24768 , \24763 , \24767 );
not \U$24426 ( \24769 , \22286 );
not \U$24427 ( \24770 , \24769 );
not \U$24428 ( \24771 , \22271 );
or \U$24429 ( \24772 , \24770 , \24771 );
nand \U$24430 ( \24773 , \24772 , \22258 );
nand \U$24431 ( \24774 , \22270 , \22286 );
and \U$24432 ( \24775 , \24773 , \24774 );
xnor \U$24433 ( \24776 , \24768 , \24775 );
xor \U$24434 ( \24777 , \24759 , \24776 );
not \U$24435 ( \24778 , \24777 );
and \U$24436 ( \24779 , \24720 , \24778 );
not \U$24437 ( \24780 , \24720 );
and \U$24438 ( \24781 , \24780 , \24777 );
nor \U$24439 ( \24782 , \24779 , \24781 );
xnor \U$24440 ( \24783 , \24592 , \24782 );
xor \U$24441 ( \24784 , \22194 , \22198 );
and \U$24442 ( \24785 , \24784 , \22403 );
and \U$24443 ( \24786 , \22194 , \22198 );
or \U$24444 ( \24787 , \24785 , \24786 );
or \U$24445 ( \24788 , \24783 , \24787 );
or \U$24446 ( \24789 , \22623 , \22631 );
nand \U$24447 ( \24790 , \24789 , \22612 );
nand \U$24448 ( \24791 , \22623 , \22631 );
nand \U$24449 ( \24792 , \24790 , \24791 );
nand \U$24450 ( \24793 , \24788 , \24792 );
nand \U$24451 ( \24794 , \24787 , \24783 );
nand \U$24452 ( \24795 , \24793 , \24794 );
xor \U$24453 ( \24796 , \22429 , \22439 );
and \U$24454 ( \24797 , \24796 , \22444 );
and \U$24455 ( \24798 , \22429 , \22439 );
or \U$24456 ( \24799 , \24797 , \24798 );
xor \U$24457 ( \24800 , \15750 , \15757 );
xor \U$24458 ( \24801 , \24800 , \15769 );
xor \U$24459 ( \24802 , \22522 , \22527 );
and \U$24460 ( \24803 , \24802 , \22533 );
and \U$24461 ( \24804 , \22522 , \22527 );
or \U$24462 ( \24805 , \24803 , \24804 );
xor \U$24463 ( \24806 , \24801 , \24805 );
not \U$24464 ( \24807 , \2922 );
not \U$24465 ( \24808 , \22435 );
or \U$24466 ( \24809 , \24807 , \24808 );
nand \U$24467 ( \24810 , \15418 , \2925 );
nand \U$24468 ( \24811 , \24809 , \24810 );
xor \U$24469 ( \24812 , \24806 , \24811 );
xor \U$24470 ( \24813 , \24799 , \24812 );
xor \U$24471 ( \24814 , \22479 , \22486 );
and \U$24472 ( \24815 , \24814 , \22494 );
and \U$24473 ( \24816 , \22479 , \22486 );
or \U$24474 ( \24817 , \24815 , \24816 );
xor \U$24475 ( \24818 , \24813 , \24817 );
xor \U$24476 ( \24819 , \22495 , \22499 );
and \U$24477 ( \24820 , \24819 , \22506 );
and \U$24478 ( \24821 , \22495 , \22499 );
or \U$24479 ( \24822 , \24820 , \24821 );
xor \U$24480 ( \24823 , \24818 , \24822 );
not \U$24481 ( \24824 , \22610 );
not \U$24482 ( \24825 , \22544 );
or \U$24483 ( \24826 , \24824 , \24825 );
or \U$24484 ( \24827 , \22610 , \22544 );
nand \U$24485 ( \24828 , \24827 , \22517 );
nand \U$24486 ( \24829 , \24826 , \24828 );
and \U$24487 ( \24830 , \24823 , \24829 );
and \U$24488 ( \24831 , \24818 , \24822 );
or \U$24489 ( \24832 , \24830 , \24831 );
xor \U$24490 ( \24833 , \15543 , \15553 );
xor \U$24491 ( \24834 , \24833 , \15565 );
xor \U$24492 ( \24835 , \15669 , \15678 );
xnor \U$24493 ( \24836 , \24835 , \15691 );
xor \U$24494 ( \24837 , \14848 , \15406 );
xor \U$24495 ( \24838 , \24837 , \15422 );
and \U$24496 ( \24839 , \24836 , \24838 );
not \U$24497 ( \24840 , \24836 );
not \U$24498 ( \24841 , \24838 );
and \U$24499 ( \24842 , \24840 , \24841 );
nor \U$24500 ( \24843 , \24839 , \24842 );
xnor \U$24501 ( \24844 , \24834 , \24843 );
not \U$24502 ( \24845 , \22470 );
nand \U$24503 ( \24846 , \24845 , \15826 );
not \U$24504 ( \24847 , \24846 );
not \U$24505 ( \24848 , \22464 );
or \U$24506 ( \24849 , \24847 , \24848 );
not \U$24507 ( \24850 , \15826 );
nand \U$24508 ( \24851 , \24850 , \22470 );
nand \U$24509 ( \24852 , \24849 , \24851 );
xor \U$24510 ( \24853 , \22203 , \22208 );
and \U$24511 ( \24854 , \24853 , \22214 );
and \U$24512 ( \24855 , \22203 , \22208 );
or \U$24513 ( \24856 , \24854 , \24855 );
xor \U$24514 ( \24857 , \24852 , \24856 );
not \U$24515 ( \24858 , \22600 );
not \U$24516 ( \24859 , \22588 );
not \U$24517 ( \24860 , \24859 );
or \U$24518 ( \24861 , \24858 , \24860 );
not \U$24519 ( \24862 , \22601 );
not \U$24520 ( \24863 , \22588 );
or \U$24521 ( \24864 , \24862 , \24863 );
nand \U$24522 ( \24865 , \24864 , \22594 );
nand \U$24523 ( \24866 , \24861 , \24865 );
xor \U$24524 ( \24867 , \24857 , \24866 );
not \U$24525 ( \24868 , \24867 );
xor \U$24526 ( \24869 , \15464 , \15478 );
xor \U$24527 ( \24870 , \24869 , \15490 );
xor \U$24528 ( \24871 , \22550 , \22561 );
and \U$24529 ( \24872 , \24871 , \22572 );
and \U$24530 ( \24873 , \22550 , \22561 );
or \U$24531 ( \24874 , \24872 , \24873 );
xor \U$24532 ( \24875 , \24870 , \24874 );
not \U$24533 ( \24876 , \22373 );
not \U$24534 ( \24877 , \22395 );
or \U$24535 ( \24878 , \24876 , \24877 );
or \U$24536 ( \24879 , \22395 , \22373 );
nand \U$24537 ( \24880 , \24879 , \22383 );
nand \U$24538 ( \24881 , \24878 , \24880 );
xnor \U$24539 ( \24882 , \24875 , \24881 );
not \U$24540 ( \24883 , \24882 );
not \U$24541 ( \24884 , \24883 );
or \U$24542 ( \24885 , \24868 , \24884 );
not \U$24543 ( \24886 , \24867 );
not \U$24544 ( \24887 , \24886 );
not \U$24545 ( \24888 , \24882 );
or \U$24546 ( \24889 , \24887 , \24888 );
not \U$24547 ( \24890 , \22573 );
not \U$24548 ( \24891 , \22609 );
or \U$24549 ( \24892 , \24890 , \24891 );
or \U$24550 ( \24893 , \22609 , \22573 );
nand \U$24551 ( \24894 , \24893 , \22577 );
nand \U$24552 ( \24895 , \24892 , \24894 );
nand \U$24553 ( \24896 , \24889 , \24895 );
nand \U$24554 ( \24897 , \24885 , \24896 );
xor \U$24555 ( \24898 , \24844 , \24897 );
xor \U$24556 ( \24899 , \24751 , \24758 );
and \U$24557 ( \24900 , \24899 , \24776 );
and \U$24558 ( \24901 , \24751 , \24758 );
or \U$24559 ( \24902 , \24900 , \24901 );
xor \U$24560 ( \24903 , \24898 , \24902 );
xor \U$24561 ( \24904 , \24832 , \24903 );
xor \U$24562 ( \24905 , \24867 , \24895 );
xor \U$24563 ( \24906 , \24905 , \24883 );
not \U$24564 ( \24907 , \22189 );
not \U$24565 ( \24908 , \22154 );
or \U$24566 ( \24909 , \24907 , \24908 );
or \U$24567 ( \24910 , \22154 , \22189 );
not \U$24568 ( \24911 , \22182 );
nand \U$24569 ( \24912 , \24910 , \24911 );
nand \U$24570 ( \24913 , \24909 , \24912 );
xor \U$24571 ( \24914 , \24906 , \24913 );
xor \U$24572 ( \24915 , \22534 , \22538 );
and \U$24573 ( \24916 , \24915 , \22543 );
and \U$24574 ( \24917 , \22534 , \22538 );
or \U$24575 ( \24918 , \24916 , \24917 );
not \U$24576 ( \24919 , \22168 );
not \U$24577 ( \24920 , \22177 );
or \U$24578 ( \24921 , \24919 , \24920 );
not \U$24579 ( \24922 , \22178 );
not \U$24580 ( \24923 , \22171 );
or \U$24581 ( \24924 , \24922 , \24923 );
nand \U$24582 ( \24925 , \24924 , \22160 );
nand \U$24583 ( \24926 , \24921 , \24925 );
xor \U$24584 ( \24927 , \24918 , \24926 );
xor \U$24585 ( \24928 , \22328 , \22363 );
and \U$24586 ( \24929 , \24928 , \22396 );
and \U$24587 ( \24930 , \22328 , \22363 );
or \U$24588 ( \24931 , \24929 , \24930 );
xor \U$24589 ( \24932 , \24927 , \24931 );
and \U$24590 ( \24933 , \24914 , \24932 );
and \U$24591 ( \24934 , \24906 , \24913 );
or \U$24592 ( \24935 , \24933 , \24934 );
xor \U$24593 ( \24936 , \24904 , \24935 );
not \U$24594 ( \24937 , \22458 );
not \U$24595 ( \24938 , \24937 );
not \U$24596 ( \24939 , \22507 );
not \U$24597 ( \24940 , \24939 );
or \U$24598 ( \24941 , \24938 , \24940 );
buf \U$24599 ( \24942 , \22425 );
nand \U$24600 ( \24943 , \24941 , \24942 );
not \U$24601 ( \24944 , \24937 );
nand \U$24602 ( \24945 , \24944 , \22507 );
nand \U$24603 ( \24946 , \24943 , \24945 );
xor \U$24604 ( \24947 , \24818 , \24822 );
xor \U$24605 ( \24948 , \24947 , \24829 );
xor \U$24606 ( \24949 , \24946 , \24948 );
xor \U$24607 ( \24950 , \24906 , \24913 );
xor \U$24608 ( \24951 , \24950 , \24932 );
and \U$24609 ( \24952 , \24949 , \24951 );
and \U$24610 ( \24953 , \24946 , \24948 );
or \U$24611 ( \24954 , \24952 , \24953 );
xor \U$24612 ( \24955 , \24936 , \24954 );
xor \U$24613 ( \24956 , \15772 , \15808 );
xor \U$24614 ( \24957 , \24956 , \15850 );
xor \U$24615 ( \24958 , \15033 , \15045 );
xor \U$24616 ( \24959 , \24958 , \15059 );
not \U$24617 ( \24960 , \24745 );
not \U$24618 ( \24961 , \24734 );
or \U$24619 ( \24962 , \24960 , \24961 );
or \U$24620 ( \24963 , \24745 , \24734 );
nand \U$24621 ( \24964 , \24963 , \24739 );
nand \U$24622 ( \24965 , \24962 , \24964 );
xor \U$24623 ( \24966 , \24959 , \24965 );
not \U$24624 ( \24967 , \24675 );
not \U$24625 ( \24968 , \24679 );
not \U$24626 ( \24969 , \22347 );
nor \U$24627 ( \24970 , \24969 , \4713 );
nor \U$24628 ( \24971 , \24968 , \24970 );
nand \U$24629 ( \24972 , \24967 , \24971 );
not \U$24630 ( \24973 , \24972 );
not \U$24631 ( \24974 , \24686 );
or \U$24632 ( \24975 , \24973 , \24974 );
nand \U$24633 ( \24976 , \24680 , \24675 );
nand \U$24634 ( \24977 , \24975 , \24976 );
xor \U$24635 ( \24978 , \24966 , \24977 );
xor \U$24636 ( \24979 , \24957 , \24978 );
nor \U$24637 ( \24980 , \24763 , \24767 );
or \U$24638 ( \24981 , \24980 , \24775 );
nand \U$24639 ( \24982 , \24767 , \24763 );
nand \U$24640 ( \24983 , \24981 , \24982 );
xor \U$24641 ( \24984 , \24979 , \24983 );
not \U$24642 ( \24985 , \24874 );
not \U$24643 ( \24986 , \24881 );
or \U$24644 ( \24987 , \24985 , \24986 );
or \U$24645 ( \24988 , \24881 , \24874 );
nand \U$24646 ( \24989 , \24988 , \24870 );
nand \U$24647 ( \24990 , \24987 , \24989 );
xor \U$24648 ( \24991 , \24722 , \24728 );
and \U$24649 ( \24992 , \24991 , \24750 );
and \U$24650 ( \24993 , \24722 , \24728 );
or \U$24651 ( \24994 , \24992 , \24993 );
xor \U$24652 ( \24995 , \24990 , \24994 );
not \U$24653 ( \24996 , \24634 );
not \U$24654 ( \24997 , \24628 );
or \U$24655 ( \24998 , \24996 , \24997 );
or \U$24656 ( \24999 , \24628 , \24634 );
nand \U$24657 ( \25000 , \24999 , \24623 );
nand \U$24658 ( \25001 , \24998 , \25000 );
not \U$24659 ( \25002 , \24602 );
not \U$24660 ( \25003 , \24612 );
or \U$24661 ( \25004 , \25002 , \25003 );
not \U$24662 ( \25005 , \24613 );
not \U$24663 ( \25006 , \24603 );
or \U$24664 ( \25007 , \25005 , \25006 );
nand \U$24665 ( \25008 , \25007 , \24597 );
nand \U$24666 ( \25009 , \25004 , \25008 );
xor \U$24667 ( \25010 , \25001 , \25009 );
buf \U$24668 ( \25011 , \24644 );
or \U$24669 ( \25012 , \24656 , \25011 );
nand \U$24670 ( \25013 , \25012 , \24649 );
nand \U$24671 ( \25014 , \24656 , \25011 );
nand \U$24672 ( \25015 , \25013 , \25014 );
xor \U$24673 ( \25016 , \25010 , \25015 );
xor \U$24674 ( \25017 , \24995 , \25016 );
xor \U$24675 ( \25018 , \24984 , \25017 );
xor \U$24676 ( \25019 , \24918 , \24926 );
and \U$24677 ( \25020 , \25019 , \24931 );
and \U$24678 ( \25021 , \24918 , \24926 );
or \U$24679 ( \25022 , \25020 , \25021 );
xor \U$24680 ( \25023 , \25018 , \25022 );
not \U$24681 ( \25024 , \24777 );
not \U$24682 ( \25025 , \24720 );
or \U$24683 ( \25026 , \25024 , \25025 );
or \U$24684 ( \25027 , \24720 , \24777 );
nand \U$24685 ( \25028 , \25027 , \24592 );
nand \U$24686 ( \25029 , \25026 , \25028 );
xor \U$24687 ( \25030 , \25023 , \25029 );
not \U$24688 ( \25031 , \24617 );
not \U$24689 ( \25032 , \25031 );
not \U$24690 ( \25033 , \24660 );
or \U$24691 ( \25034 , \25032 , \25033 );
not \U$24692 ( \25035 , \24657 );
not \U$24693 ( \25036 , \24617 );
or \U$24694 ( \25037 , \25035 , \25036 );
nand \U$24695 ( \25038 , \25037 , \24635 );
nand \U$24696 ( \25039 , \25034 , \25038 );
not \U$24697 ( \25040 , \24670 );
not \U$24698 ( \25041 , \24705 );
or \U$24699 ( \25042 , \25040 , \25041 );
or \U$24700 ( \25043 , \24670 , \24705 );
nand \U$24701 ( \25044 , \25043 , \24687 );
nand \U$24702 ( \25045 , \25042 , \25044 );
xor \U$24703 ( \25046 , \15173 , \15184 );
xor \U$24704 ( \25047 , \25046 , \15196 );
xor \U$24705 ( \25048 , \15113 , \15122 );
xor \U$24706 ( \25049 , \25048 , \15134 );
xor \U$24707 ( \25050 , \25047 , \25049 );
xor \U$24708 ( \25051 , \24693 , \24698 );
and \U$24709 ( \25052 , \25051 , \24704 );
and \U$24710 ( \25053 , \24693 , \24698 );
or \U$24711 ( \25054 , \25052 , \25053 );
xor \U$24712 ( \25055 , \25050 , \25054 );
not \U$24713 ( \25056 , \25055 );
and \U$24714 ( \25057 , \25045 , \25056 );
not \U$24715 ( \25058 , \25045 );
and \U$24716 ( \25059 , \25058 , \25055 );
nor \U$24717 ( \25060 , \25057 , \25059 );
xnor \U$24718 ( \25061 , \25039 , \25060 );
not \U$24719 ( \25062 , \24662 );
not \U$24720 ( \25063 , \25062 );
not \U$24721 ( \25064 , \24706 );
or \U$24722 ( \25065 , \25063 , \25064 );
or \U$24723 ( \25066 , \24706 , \25062 );
nand \U$24724 ( \25067 , \25066 , \24715 );
nand \U$24725 ( \25068 , \25065 , \25067 );
xor \U$24726 ( \25069 , \25061 , \25068 );
xor \U$24727 ( \25070 , \15084 , \15072 );
xor \U$24728 ( \25071 , \25070 , \15097 );
xor \U$24729 ( \25072 , \24801 , \24805 );
and \U$24730 ( \25073 , \25072 , \24811 );
and \U$24731 ( \25074 , \24801 , \24805 );
or \U$24732 ( \25075 , \25073 , \25074 );
xor \U$24733 ( \25076 , \25071 , \25075 );
xor \U$24734 ( \25077 , \15437 , \15450 );
xor \U$24735 ( \25078 , \25077 , \15493 );
xor \U$24736 ( \25079 , \25076 , \25078 );
xor \U$24737 ( \25080 , \15638 , \15649 );
xor \U$24738 ( \25081 , \25080 , \15626 );
xor \U$24739 ( \25082 , \15613 , \15589 );
xor \U$24740 ( \25083 , \25082 , \15600 );
xor \U$24741 ( \25084 , \25081 , \25083 );
xor \U$24742 ( \25085 , \24852 , \24856 );
and \U$24743 ( \25086 , \25085 , \24866 );
and \U$24744 ( \25087 , \24852 , \24856 );
or \U$24745 ( \25088 , \25086 , \25087 );
xor \U$24746 ( \25089 , \25084 , \25088 );
xor \U$24747 ( \25090 , \25079 , \25089 );
xor \U$24748 ( \25091 , \24799 , \24812 );
and \U$24749 ( \25092 , \25091 , \24817 );
and \U$24750 ( \25093 , \24799 , \24812 );
or \U$24751 ( \25094 , \25092 , \25093 );
xor \U$24752 ( \25095 , \25090 , \25094 );
xor \U$24753 ( \25096 , \25069 , \25095 );
xor \U$24754 ( \25097 , \25030 , \25096 );
xor \U$24755 ( \25098 , \24955 , \25097 );
xor \U$24756 ( \25099 , \24795 , \25098 );
xor \U$24757 ( \25100 , \24946 , \24948 );
xor \U$24758 ( \25101 , \25100 , \24951 );
buf \U$24759 ( \25102 , \25101 );
not \U$24760 ( \25103 , \25102 );
buf \U$24761 ( \25104 , \22142 );
not \U$24762 ( \25105 , \25104 );
buf \U$24763 ( \25106 , \22404 );
not \U$24764 ( \25107 , \25106 );
or \U$24765 ( \25108 , \25105 , \25107 );
or \U$24766 ( \25109 , \25106 , \25104 );
buf \U$24767 ( \25110 , \22146 );
nand \U$24768 ( \25111 , \25109 , \25110 );
nand \U$24769 ( \25112 , \25108 , \25111 );
not \U$24770 ( \25113 , \25112 );
or \U$24771 ( \25114 , \25103 , \25113 );
or \U$24772 ( \25115 , \25112 , \25102 );
xor \U$24773 ( \25116 , \22419 , \22508 );
and \U$24774 ( \25117 , \25116 , \22636 );
and \U$24775 ( \25118 , \22419 , \22508 );
or \U$24776 ( \25119 , \25117 , \25118 );
not \U$24777 ( \25120 , \25119 );
nand \U$24778 ( \25121 , \25115 , \25120 );
nand \U$24779 ( \25122 , \25114 , \25121 );
xnor \U$24780 ( \25123 , \25099 , \25122 );
xor \U$24781 ( \25124 , \24792 , \24787 );
xnor \U$24782 ( \25125 , \25124 , \24783 );
not \U$24783 ( \25126 , \22638 );
nand \U$24784 ( \25127 , \25126 , \22405 );
buf \U$24785 ( \25128 , \22410 );
and \U$24786 ( \25129 , \25127 , \25128 );
nor \U$24787 ( \25130 , \22405 , \22637 );
nor \U$24788 ( \25131 , \25129 , \25130 );
xor \U$24789 ( \25132 , \25125 , \25131 );
not \U$24790 ( \25133 , \25119 );
not \U$24791 ( \25134 , \25101 );
or \U$24792 ( \25135 , \25133 , \25134 );
or \U$24793 ( \25136 , \25119 , \25101 );
nand \U$24794 ( \25137 , \25135 , \25136 );
not \U$24795 ( \25138 , \25112 );
and \U$24796 ( \25139 , \25137 , \25138 );
not \U$24797 ( \25140 , \25137 );
and \U$24798 ( \25141 , \25140 , \25112 );
nor \U$24799 ( \25142 , \25139 , \25141 );
and \U$24800 ( \25143 , \25132 , \25142 );
and \U$24801 ( \25144 , \25125 , \25131 );
or \U$24802 ( \25145 , \25143 , \25144 );
nand \U$24803 ( \25146 , \25123 , \25145 );
xor \U$24804 ( \25147 , \25125 , \25131 );
xor \U$24805 ( \25148 , \25147 , \25142 );
xor \U$24806 ( \25149 , \22128 , \22132 );
and \U$24807 ( \25150 , \25149 , \22646 );
and \U$24808 ( \25151 , \22128 , \22132 );
or \U$24809 ( \25152 , \25150 , \25151 );
not \U$24810 ( \25153 , \25152 );
nand \U$24811 ( \25154 , \25148 , \25153 );
and \U$24812 ( \25155 , \25146 , \25154 );
xor \U$24813 ( \25156 , \15698 , \15499 );
xnor \U$24814 ( \25157 , \25156 , \15502 );
not \U$24815 ( \25158 , \25157 );
xnor \U$24816 ( \25159 , \15712 , \15855 );
and \U$24817 ( \25160 , \25159 , \15719 );
not \U$24818 ( \25161 , \25159 );
and \U$24819 ( \25162 , \25161 , \15858 );
nor \U$24820 ( \25163 , \25160 , \25162 );
not \U$24821 ( \25164 , \25163 );
not \U$24822 ( \25165 , \25164 );
xor \U$24823 ( \25166 , \15385 , \15369 );
xor \U$24824 ( \25167 , \25166 , \15497 );
not \U$24825 ( \25168 , \25167 );
not \U$24826 ( \25169 , \25168 );
or \U$24827 ( \25170 , \25165 , \25169 );
not \U$24828 ( \25171 , \25167 );
not \U$24829 ( \25172 , \25163 );
or \U$24830 ( \25173 , \25171 , \25172 );
not \U$24831 ( \25174 , \15373 );
not \U$24832 ( \25175 , \25174 );
not \U$24833 ( \25176 , \15377 );
or \U$24834 ( \25177 , \25175 , \25176 );
nand \U$24835 ( \25178 , \15376 , \15373 );
nand \U$24836 ( \25179 , \25177 , \25178 );
and \U$24837 ( \25180 , \25179 , \15383 );
not \U$24838 ( \25181 , \25179 );
not \U$24839 ( \25182 , \15383 );
and \U$24840 ( \25183 , \25181 , \25182 );
nor \U$24841 ( \25184 , \25180 , \25183 );
buf \U$24842 ( \25185 , \25184 );
not \U$24843 ( \25186 , \25185 );
not \U$24844 ( \25187 , \25186 );
not \U$24845 ( \25188 , \15724 );
not \U$24846 ( \25189 , \15733 );
or \U$24847 ( \25190 , \25188 , \25189 );
nand \U$24848 ( \25191 , \15732 , \15723 );
nand \U$24849 ( \25192 , \25190 , \25191 );
not \U$24850 ( \25193 , \15853 );
and \U$24851 ( \25194 , \25192 , \25193 );
not \U$24852 ( \25195 , \25192 );
and \U$24853 ( \25196 , \25195 , \15853 );
nor \U$24854 ( \25197 , \25194 , \25196 );
buf \U$24855 ( \25198 , \25197 );
not \U$24856 ( \25199 , \25198 );
or \U$24857 ( \25200 , \25187 , \25199 );
xor \U$24858 ( \25201 , \25081 , \25083 );
and \U$24859 ( \25202 , \25201 , \25088 );
and \U$24860 ( \25203 , \25081 , \25083 );
or \U$24861 ( \25204 , \25202 , \25203 );
nand \U$24862 ( \25205 , \25200 , \25204 );
not \U$24863 ( \25206 , \25198 );
nand \U$24864 ( \25207 , \25206 , \25185 );
nand \U$24865 ( \25208 , \25205 , \25207 );
nand \U$24866 ( \25209 , \25173 , \25208 );
nand \U$24867 ( \25210 , \25170 , \25209 );
buf \U$24868 ( \25211 , \25210 );
xor \U$24869 ( \25212 , \25158 , \25211 );
xor \U$24870 ( \25213 , \15710 , \15860 );
xor \U$24871 ( \25214 , \25213 , \15863 );
xor \U$24872 ( \25215 , \25212 , \25214 );
xor \U$24873 ( \25216 , \24844 , \24897 );
and \U$24874 ( \25217 , \25216 , \24902 );
and \U$24875 ( \25218 , \24844 , \24897 );
or \U$24876 ( \25219 , \25217 , \25218 );
not \U$24877 ( \25220 , \15495 );
xor \U$24878 ( \25221 , \15390 , \15424 );
not \U$24879 ( \25222 , \25221 );
or \U$24880 ( \25223 , \25220 , \25222 );
or \U$24881 ( \25224 , \25221 , \15495 );
nand \U$24882 ( \25225 , \25223 , \25224 );
xor \U$24883 ( \25226 , \24957 , \24978 );
and \U$24884 ( \25227 , \25226 , \24983 );
and \U$24885 ( \25228 , \24957 , \24978 );
or \U$24886 ( \25229 , \25227 , \25228 );
xor \U$24887 ( \25230 , \25225 , \25229 );
nand \U$24888 ( \25231 , \24705 , \24670 );
nand \U$24889 ( \25232 , \25044 , \25231 );
or \U$24890 ( \25233 , \25232 , \25039 );
nand \U$24891 ( \25234 , \25233 , \25055 );
nand \U$24892 ( \25235 , \25232 , \25039 );
nand \U$24893 ( \25236 , \25234 , \25235 );
xor \U$24894 ( \25237 , \25230 , \25236 );
or \U$24895 ( \25238 , \25219 , \25237 );
xor \U$24896 ( \25239 , \24984 , \25017 );
and \U$24897 ( \25240 , \25239 , \25022 );
and \U$24898 ( \25241 , \24984 , \25017 );
or \U$24899 ( \25242 , \25240 , \25241 );
nand \U$24900 ( \25243 , \25238 , \25242 );
nand \U$24901 ( \25244 , \25237 , \25219 );
nand \U$24902 ( \25245 , \25243 , \25244 );
xor \U$24903 ( \25246 , \25225 , \25229 );
and \U$24904 ( \25247 , \25246 , \25236 );
and \U$24905 ( \25248 , \25225 , \25229 );
or \U$24906 ( \25249 , \25247 , \25248 );
xor \U$24907 ( \25250 , \15014 , \15016 );
xor \U$24908 ( \25251 , \25250 , \15140 );
xor \U$24909 ( \25252 , \15157 , \15202 );
xor \U$24910 ( \25253 , \25252 , \15205 );
xor \U$24911 ( \25254 , \25251 , \25253 );
xor \U$24912 ( \25255 , \15062 , \15099 );
xor \U$24913 ( \25256 , \25255 , \15137 );
xor \U$24914 ( \25257 , \15159 , \15162 );
xor \U$24915 ( \25258 , \25257 , \15199 );
xor \U$24916 ( \25259 , \25256 , \25258 );
xor \U$24917 ( \25260 , \25047 , \25049 );
and \U$24918 ( \25261 , \25260 , \25054 );
and \U$24919 ( \25262 , \25047 , \25049 );
or \U$24920 ( \25263 , \25261 , \25262 );
and \U$24921 ( \25264 , \25259 , \25263 );
and \U$24922 ( \25265 , \25256 , \25258 );
or \U$24923 ( \25266 , \25264 , \25265 );
xor \U$24924 ( \25267 , \25254 , \25266 );
xor \U$24925 ( \25268 , \25249 , \25267 );
xor \U$24926 ( \25269 , \25256 , \25258 );
xor \U$24927 ( \25270 , \25269 , \25263 );
xor \U$24928 ( \25271 , \24990 , \24994 );
and \U$24929 ( \25272 , \25271 , \25016 );
and \U$24930 ( \25273 , \24990 , \24994 );
or \U$24931 ( \25274 , \25272 , \25273 );
xor \U$24932 ( \25275 , \25270 , \25274 );
xor \U$24933 ( \25276 , \24959 , \24965 );
and \U$24934 ( \25277 , \25276 , \24977 );
and \U$24935 ( \25278 , \24959 , \24965 );
or \U$24936 ( \25279 , \25277 , \25278 );
not \U$24937 ( \25280 , \25009 );
not \U$24938 ( \25281 , \25001 );
or \U$24939 ( \25282 , \25280 , \25281 );
or \U$24940 ( \25283 , \25001 , \25009 );
nand \U$24941 ( \25284 , \25283 , \25015 );
nand \U$24942 ( \25285 , \25282 , \25284 );
xor \U$24943 ( \25286 , \25279 , \25285 );
not \U$24944 ( \25287 , \15694 );
not \U$24945 ( \25288 , \15657 );
or \U$24946 ( \25289 , \25287 , \25288 );
not \U$24947 ( \25290 , \15694 );
nand \U$24948 ( \25291 , \25290 , \15652 );
nand \U$24949 ( \25292 , \25289 , \25291 );
buf \U$24950 ( \25293 , \15615 );
and \U$24951 ( \25294 , \25292 , \25293 );
not \U$24952 ( \25295 , \25292 );
not \U$24953 ( \25296 , \25293 );
and \U$24954 ( \25297 , \25295 , \25296 );
nor \U$24955 ( \25298 , \25294 , \25297 );
xor \U$24956 ( \25299 , \25286 , \25298 );
and \U$24957 ( \25300 , \25275 , \25299 );
and \U$24958 ( \25301 , \25270 , \25274 );
or \U$24959 ( \25302 , \25300 , \25301 );
xor \U$24960 ( \25303 , \25268 , \25302 );
xor \U$24961 ( \25304 , \25245 , \25303 );
xor \U$24962 ( \25305 , \25270 , \25274 );
xor \U$24963 ( \25306 , \25305 , \25299 );
not \U$24964 ( \25307 , \25306 );
or \U$24965 ( \25308 , \24834 , \24836 );
nand \U$24966 ( \25309 , \25308 , \24841 );
nand \U$24967 ( \25310 , \24834 , \24836 );
nand \U$24968 ( \25311 , \25309 , \25310 );
not \U$24969 ( \25312 , \15516 );
not \U$24970 ( \25313 , \15528 );
or \U$24971 ( \25314 , \25312 , \25313 );
nand \U$24972 ( \25315 , \15517 , \15527 );
nand \U$24973 ( \25316 , \25314 , \25315 );
and \U$24974 ( \25317 , \25316 , \15568 );
not \U$24975 ( \25318 , \25316 );
not \U$24976 ( \25319 , \15568 );
and \U$24977 ( \25320 , \25318 , \25319 );
nor \U$24978 ( \25321 , \25317 , \25320 );
xor \U$24979 ( \25322 , \25311 , \25321 );
xor \U$24980 ( \25323 , \25071 , \25075 );
and \U$24981 ( \25324 , \25323 , \25078 );
and \U$24982 ( \25325 , \25071 , \25075 );
or \U$24983 ( \25326 , \25324 , \25325 );
xor \U$24984 ( \25327 , \25322 , \25326 );
not \U$24985 ( \25328 , \25327 );
not \U$24986 ( \25329 , \25328 );
not \U$24987 ( \25330 , \25184 );
not \U$24988 ( \25331 , \25197 );
or \U$24989 ( \25332 , \25330 , \25331 );
or \U$24990 ( \25333 , \25184 , \25197 );
nand \U$24991 ( \25334 , \25332 , \25333 );
not \U$24992 ( \25335 , \25204 );
and \U$24993 ( \25336 , \25334 , \25335 );
not \U$24994 ( \25337 , \25334 );
and \U$24995 ( \25338 , \25337 , \25204 );
nor \U$24996 ( \25339 , \25336 , \25338 );
not \U$24997 ( \25340 , \25339 );
not \U$24998 ( \25341 , \25340 );
or \U$24999 ( \25342 , \25329 , \25341 );
nand \U$25000 ( \25343 , \25339 , \25327 );
nand \U$25001 ( \25344 , \25342 , \25343 );
xor \U$25002 ( \25345 , \25079 , \25089 );
and \U$25003 ( \25346 , \25345 , \25094 );
and \U$25004 ( \25347 , \25079 , \25089 );
or \U$25005 ( \25348 , \25346 , \25347 );
not \U$25006 ( \25349 , \25348 );
and \U$25007 ( \25350 , \25344 , \25349 );
not \U$25008 ( \25351 , \25344 );
and \U$25009 ( \25352 , \25351 , \25348 );
nor \U$25010 ( \25353 , \25350 , \25352 );
nand \U$25011 ( \25354 , \25307 , \25353 );
not \U$25012 ( \25355 , \25354 );
xor \U$25013 ( \25356 , \25061 , \25068 );
and \U$25014 ( \25357 , \25356 , \25095 );
and \U$25015 ( \25358 , \25061 , \25068 );
or \U$25016 ( \25359 , \25357 , \25358 );
not \U$25017 ( \25360 , \25359 );
or \U$25018 ( \25361 , \25355 , \25360 );
not \U$25019 ( \25362 , \25353 );
nand \U$25020 ( \25363 , \25362 , \25306 );
nand \U$25021 ( \25364 , \25361 , \25363 );
and \U$25022 ( \25365 , \25304 , \25364 );
and \U$25023 ( \25366 , \25245 , \25303 );
or \U$25024 ( \25367 , \25365 , \25366 );
xor \U$25025 ( \25368 , \25215 , \25367 );
xor \U$25026 ( \25369 , \25249 , \25267 );
and \U$25027 ( \25370 , \25369 , \25302 );
and \U$25028 ( \25371 , \25249 , \25267 );
or \U$25029 ( \25372 , \25370 , \25371 );
xor \U$25030 ( \25373 , \25251 , \25253 );
and \U$25031 ( \25374 , \25373 , \25266 );
and \U$25032 ( \25375 , \25251 , \25253 );
or \U$25033 ( \25376 , \25374 , \25375 );
xor \U$25034 ( \25377 , \15152 , \15154 );
xor \U$25035 ( \25378 , \25377 , \15208 );
xor \U$25036 ( \25379 , \25376 , \25378 );
or \U$25037 ( \25380 , \25285 , \25298 );
nand \U$25038 ( \25381 , \25380 , \25279 );
nand \U$25039 ( \25382 , \25298 , \25285 );
nand \U$25040 ( \25383 , \25381 , \25382 );
not \U$25041 ( \25384 , \25383 );
not \U$25042 ( \25385 , \15570 );
not \U$25043 ( \25386 , \15696 );
not \U$25044 ( \25387 , \25386 );
or \U$25045 ( \25388 , \25385 , \25387 );
not \U$25046 ( \25389 , \15570 );
nand \U$25047 ( \25390 , \25389 , \15696 );
nand \U$25048 ( \25391 , \25388 , \25390 );
not \U$25049 ( \25392 , \15574 );
and \U$25050 ( \25393 , \25391 , \25392 );
not \U$25051 ( \25394 , \25391 );
and \U$25052 ( \25395 , \25394 , \15574 );
nor \U$25053 ( \25396 , \25393 , \25395 );
not \U$25054 ( \25397 , \25396 );
not \U$25055 ( \25398 , \25397 );
or \U$25056 ( \25399 , \25384 , \25398 );
not \U$25057 ( \25400 , \25383 );
not \U$25058 ( \25401 , \25400 );
not \U$25059 ( \25402 , \25396 );
or \U$25060 ( \25403 , \25401 , \25402 );
xor \U$25061 ( \25404 , \25311 , \25321 );
and \U$25062 ( \25405 , \25404 , \25326 );
and \U$25063 ( \25406 , \25311 , \25321 );
or \U$25064 ( \25407 , \25405 , \25406 );
nand \U$25065 ( \25408 , \25403 , \25407 );
nand \U$25066 ( \25409 , \25399 , \25408 );
xor \U$25067 ( \25410 , \25379 , \25409 );
xor \U$25068 ( \25411 , \25372 , \25410 );
and \U$25069 ( \25412 , \25400 , \25397 );
not \U$25070 ( \25413 , \25400 );
and \U$25071 ( \25414 , \25413 , \25396 );
or \U$25072 ( \25415 , \25412 , \25414 );
xor \U$25073 ( \25416 , \25415 , \25407 );
not \U$25074 ( \25417 , \25416 );
not \U$25075 ( \25418 , \25167 );
not \U$25076 ( \25419 , \25164 );
or \U$25077 ( \25420 , \25418 , \25419 );
nand \U$25078 ( \25421 , \25163 , \25168 );
nand \U$25079 ( \25422 , \25420 , \25421 );
buf \U$25080 ( \25423 , \25208 );
and \U$25081 ( \25424 , \25422 , \25423 );
not \U$25082 ( \25425 , \25422 );
not \U$25083 ( \25426 , \25423 );
and \U$25084 ( \25427 , \25425 , \25426 );
nor \U$25085 ( \25428 , \25424 , \25427 );
not \U$25086 ( \25429 , \25428 );
or \U$25087 ( \25430 , \25417 , \25429 );
or \U$25088 ( \25431 , \25428 , \25416 );
buf \U$25089 ( \25432 , \25339 );
not \U$25090 ( \25433 , \25327 );
nand \U$25091 ( \25434 , \25432 , \25433 );
not \U$25092 ( \25435 , \25434 );
not \U$25093 ( \25436 , \25348 );
or \U$25094 ( \25437 , \25435 , \25436 );
or \U$25095 ( \25438 , \25433 , \25432 );
nand \U$25096 ( \25439 , \25437 , \25438 );
nand \U$25097 ( \25440 , \25431 , \25439 );
nand \U$25098 ( \25441 , \25430 , \25440 );
xor \U$25099 ( \25442 , \25411 , \25441 );
and \U$25100 ( \25443 , \25368 , \25442 );
and \U$25101 ( \25444 , \25215 , \25367 );
or \U$25102 ( \25445 , \25443 , \25444 );
xor \U$25103 ( \25446 , \15708 , \15866 );
xor \U$25104 ( \25447 , \25446 , \15869 );
nor \U$25105 ( \25448 , \25378 , \25409 );
not \U$25106 ( \25449 , \25376 );
or \U$25107 ( \25450 , \25448 , \25449 );
nand \U$25108 ( \25451 , \25409 , \25378 );
nand \U$25109 ( \25452 , \25450 , \25451 );
xor \U$25110 ( \25453 , \15364 , \15366 );
xor \U$25111 ( \25454 , \25453 , \15700 );
xor \U$25112 ( \25455 , \25452 , \25454 );
not \U$25113 ( \25456 , \25210 );
not \U$25114 ( \25457 , \25158 );
or \U$25115 ( \25458 , \25456 , \25457 );
not \U$25116 ( \25459 , \25157 );
not \U$25117 ( \25460 , \25210 );
not \U$25118 ( \25461 , \25460 );
or \U$25119 ( \25462 , \25459 , \25461 );
nand \U$25120 ( \25463 , \25462 , \25214 );
nand \U$25121 ( \25464 , \25458 , \25463 );
xor \U$25122 ( \25465 , \25455 , \25464 );
xor \U$25123 ( \25466 , \25447 , \25465 );
xor \U$25124 ( \25467 , \25372 , \25410 );
and \U$25125 ( \25468 , \25467 , \25441 );
and \U$25126 ( \25469 , \25372 , \25410 );
or \U$25127 ( \25470 , \25468 , \25469 );
xor \U$25128 ( \25471 , \25466 , \25470 );
nor \U$25129 ( \25472 , \25445 , \25471 );
not \U$25130 ( \25473 , \25472 );
xor \U$25131 ( \25474 , \25215 , \25367 );
xor \U$25132 ( \25475 , \25474 , \25442 );
not \U$25133 ( \25476 , \25475 );
xnor \U$25134 ( \25477 , \25439 , \25416 );
buf \U$25135 ( \25478 , \25428 );
not \U$25136 ( \25479 , \25478 );
and \U$25137 ( \25480 , \25477 , \25479 );
not \U$25138 ( \25481 , \25477 );
and \U$25139 ( \25482 , \25481 , \25478 );
nor \U$25140 ( \25483 , \25480 , \25482 );
not \U$25141 ( \25484 , \25483 );
xor \U$25142 ( \25485 , \25245 , \25303 );
xor \U$25143 ( \25486 , \25485 , \25364 );
not \U$25144 ( \25487 , \25486 );
or \U$25145 ( \25488 , \25484 , \25487 );
or \U$25146 ( \25489 , \25486 , \25483 );
xor \U$25147 ( \25490 , \25237 , \25242 );
xor \U$25148 ( \25491 , \25490 , \25219 );
not \U$25149 ( \25492 , \25491 );
xor \U$25150 ( \25493 , \25023 , \25029 );
and \U$25151 ( \25494 , \25493 , \25096 );
and \U$25152 ( \25495 , \25023 , \25029 );
or \U$25153 ( \25496 , \25494 , \25495 );
not \U$25154 ( \25497 , \25496 );
or \U$25155 ( \25498 , \25492 , \25497 );
or \U$25156 ( \25499 , \25491 , \25496 );
xor \U$25157 ( \25500 , \24832 , \24903 );
and \U$25158 ( \25501 , \25500 , \24935 );
and \U$25159 ( \25502 , \24832 , \24903 );
or \U$25160 ( \25503 , \25501 , \25502 );
nand \U$25161 ( \25504 , \25499 , \25503 );
nand \U$25162 ( \25505 , \25498 , \25504 );
nand \U$25163 ( \25506 , \25489 , \25505 );
nand \U$25164 ( \25507 , \25488 , \25506 );
not \U$25165 ( \25508 , \25507 );
nand \U$25166 ( \25509 , \25476 , \25508 );
nand \U$25167 ( \25510 , \25473 , \25509 );
xor \U$25168 ( \25511 , \15879 , \15877 );
xnor \U$25169 ( \25512 , \25511 , \15883 );
xor \U$25170 ( \25513 , \15217 , \15214 );
xnor \U$25171 ( \25514 , \25513 , \15008 );
xor \U$25172 ( \25515 , \25452 , \25454 );
and \U$25173 ( \25516 , \25515 , \25464 );
and \U$25174 ( \25517 , \25452 , \25454 );
or \U$25175 ( \25518 , \25516 , \25517 );
not \U$25176 ( \25519 , \25518 );
xor \U$25177 ( \25520 , \25514 , \25519 );
xor \U$25178 ( \25521 , \15361 , \15704 );
xor \U$25179 ( \25522 , \25521 , \15872 );
and \U$25180 ( \25523 , \25520 , \25522 );
and \U$25181 ( \25524 , \25514 , \25519 );
or \U$25182 ( \25525 , \25523 , \25524 );
nand \U$25183 ( \25526 , \25512 , \25525 );
xor \U$25184 ( \25527 , \25514 , \25519 );
xor \U$25185 ( \25528 , \25527 , \25522 );
not \U$25186 ( \25529 , \25447 );
not \U$25187 ( \25530 , \25465 );
nand \U$25188 ( \25531 , \25529 , \25530 );
and \U$25189 ( \25532 , \25531 , \25470 );
not \U$25190 ( \25533 , \25447 );
nor \U$25191 ( \25534 , \25533 , \25530 );
nor \U$25192 ( \25535 , \25532 , \25534 );
nand \U$25193 ( \25536 , \25528 , \25535 );
nand \U$25194 ( \25537 , \25526 , \25536 );
nor \U$25195 ( \25538 , \25510 , \25537 );
not \U$25196 ( \25539 , \24795 );
not \U$25197 ( \25540 , \25098 );
nand \U$25198 ( \25541 , \25539 , \25540 );
not \U$25199 ( \25542 , \25541 );
not \U$25200 ( \25543 , \25122 );
or \U$25201 ( \25544 , \25542 , \25543 );
not \U$25202 ( \25545 , \25540 );
nand \U$25203 ( \25546 , \25545 , \24795 );
nand \U$25204 ( \25547 , \25544 , \25546 );
not \U$25205 ( \25548 , \25547 );
buf \U$25206 ( \25549 , \25362 );
not \U$25207 ( \25550 , \25549 );
xnor \U$25208 ( \25551 , \25359 , \25306 );
not \U$25209 ( \25552 , \25551 );
or \U$25210 ( \25553 , \25550 , \25552 );
or \U$25211 ( \25554 , \25551 , \25549 );
nand \U$25212 ( \25555 , \25553 , \25554 );
xor \U$25213 ( \25556 , \25503 , \25491 );
xnor \U$25214 ( \25557 , \25556 , \25496 );
xor \U$25215 ( \25558 , \25555 , \25557 );
xor \U$25216 ( \25559 , \24936 , \24954 );
and \U$25217 ( \25560 , \25559 , \25097 );
and \U$25218 ( \25561 , \24936 , \24954 );
or \U$25219 ( \25562 , \25560 , \25561 );
xnor \U$25220 ( \25563 , \25558 , \25562 );
not \U$25221 ( \25564 , \25563 );
nand \U$25222 ( \25565 , \25548 , \25564 );
xnor \U$25223 ( \25566 , \25486 , \25483 );
xnor \U$25224 ( \25567 , \25566 , \25505 );
not \U$25225 ( \25568 , \25555 );
not \U$25226 ( \25569 , \25568 );
not \U$25227 ( \25570 , \25557 );
or \U$25228 ( \25571 , \25569 , \25570 );
nand \U$25229 ( \25572 , \25571 , \25562 );
not \U$25230 ( \25573 , \25557 );
nand \U$25231 ( \25574 , \25573 , \25555 );
nand \U$25232 ( \25575 , \25572 , \25574 );
nor \U$25233 ( \25576 , \25567 , \25575 );
not \U$25234 ( \25577 , \25576 );
and \U$25235 ( \25578 , \25155 , \25538 , \25565 , \25577 );
not \U$25236 ( \25579 , \25578 );
or \U$25237 ( \25580 , \24588 , \25579 );
not \U$25238 ( \25581 , \25565 );
not \U$25239 ( \25582 , \25148 );
nand \U$25240 ( \25583 , \25582 , \25152 );
not \U$25241 ( \25584 , \25146 );
or \U$25242 ( \25585 , \25583 , \25584 );
or \U$25243 ( \25586 , \25123 , \25145 );
nand \U$25244 ( \25587 , \25585 , \25586 );
not \U$25245 ( \25588 , \25587 );
or \U$25246 ( \25589 , \25581 , \25588 );
nand \U$25247 ( \25590 , \25563 , \25547 );
nand \U$25248 ( \25591 , \25567 , \25575 );
and \U$25249 ( \25592 , \25590 , \25591 );
nand \U$25250 ( \25593 , \25589 , \25592 );
nand \U$25251 ( \25594 , \25538 , \25577 );
not \U$25252 ( \25595 , \25594 );
and \U$25253 ( \25596 , \25593 , \25595 );
not \U$25254 ( \25597 , \25536 );
nand \U$25255 ( \25598 , \25475 , \25507 );
or \U$25256 ( \25599 , \25472 , \25598 );
nand \U$25257 ( \25600 , \25471 , \25445 );
nand \U$25258 ( \25601 , \25599 , \25600 );
not \U$25259 ( \25602 , \25601 );
or \U$25260 ( \25603 , \25597 , \25602 );
or \U$25261 ( \25604 , \25528 , \25535 );
nand \U$25262 ( \25605 , \25603 , \25604 );
not \U$25263 ( \25606 , \25605 );
buf \U$25264 ( \25607 , \25526 );
not \U$25265 ( \25608 , \25607 );
or \U$25266 ( \25609 , \25606 , \25608 );
not \U$25267 ( \25610 , \25512 );
not \U$25268 ( \25611 , \25525 );
nand \U$25269 ( \25612 , \25610 , \25611 );
nand \U$25270 ( \25613 , \25609 , \25612 );
nor \U$25271 ( \25614 , \25596 , \25613 );
nand \U$25272 ( \25615 , \25580 , \25614 );
not \U$25273 ( \25616 , \17275 );
not \U$25274 ( \25617 , RIbb2d900_63);
not \U$25275 ( \25618 , \19733 );
or \U$25276 ( \25619 , \25617 , \25618 );
nand \U$25277 ( \25620 , \1337 , \20254 );
nand \U$25278 ( \25621 , \25619 , \25620 );
not \U$25279 ( \25622 , \25621 );
or \U$25280 ( \25623 , \25616 , \25622 );
and \U$25281 ( \25624 , RIbb2d900_63, \22684 );
not \U$25282 ( \25625 , RIbb2d900_63);
and \U$25283 ( \25626 , \25625 , \1419 );
or \U$25284 ( \25627 , \25624 , \25626 );
nand \U$25285 ( \25628 , \25627 , RIbb2d888_64);
nand \U$25286 ( \25629 , \25623 , \25628 );
not \U$25287 ( \25630 , \17397 );
not \U$25288 ( \25631 , RIbb2dbd0_57);
not \U$25289 ( \25632 , \6107 );
or \U$25290 ( \25633 , \25631 , \25632 );
nand \U$25291 ( \25634 , \3167 , \17411 );
nand \U$25292 ( \25635 , \25633 , \25634 );
not \U$25293 ( \25636 , \25635 );
or \U$25294 ( \25637 , \25630 , \25636 );
not \U$25295 ( \25638 , RIbb2dbd0_57);
not \U$25296 ( \25639 , \22978 );
or \U$25297 ( \25640 , \25638 , \25639 );
nand \U$25298 ( \25641 , \3146 , \17411 );
nand \U$25299 ( \25642 , \25640 , \25641 );
nand \U$25300 ( \25643 , \25642 , \16675 );
nand \U$25301 ( \25644 , \25637 , \25643 );
or \U$25302 ( \25645 , \25629 , \25644 );
not \U$25303 ( \25646 , \15181 );
not \U$25304 ( \25647 , RIbb2dcc0_55);
not \U$25305 ( \25648 , \14791 );
or \U$25306 ( \25649 , \25647 , \25648 );
not \U$25307 ( \25650 , RIbb2dcc0_55);
nand \U$25308 ( \25651 , \25650 , \4637 );
nand \U$25309 ( \25652 , \25649 , \25651 );
not \U$25310 ( \25653 , \25652 );
or \U$25311 ( \25654 , \25646 , \25653 );
and \U$25312 ( \25655 , RIbb2dcc0_55, \13835 );
not \U$25313 ( \25656 , RIbb2dcc0_55);
and \U$25314 ( \25657 , \25656 , \6171 );
or \U$25315 ( \25658 , \25655 , \25657 );
nand \U$25316 ( \25659 , \25658 , \14613 );
nand \U$25317 ( \25660 , \25654 , \25659 );
nand \U$25318 ( \25661 , \25645 , \25660 );
nand \U$25319 ( \25662 , \25629 , \25644 );
nand \U$25320 ( \25663 , \25661 , \25662 );
not \U$25321 ( \25664 , \17470 );
and \U$25322 ( \25665 , RIbb2dae0_59, \2223 );
not \U$25323 ( \25666 , RIbb2dae0_59);
and \U$25324 ( \25667 , \25666 , \3320 );
or \U$25325 ( \25668 , \25665 , \25667 );
not \U$25326 ( \25669 , \25668 );
or \U$25327 ( \25670 , \25664 , \25669 );
not \U$25328 ( \25671 , RIbb2dae0_59);
not \U$25329 ( \25672 , \3520 );
or \U$25330 ( \25673 , \25671 , \25672 );
not \U$25331 ( \25674 , \3342 );
not \U$25332 ( \25675 , RIbb2dae0_59);
nand \U$25333 ( \25676 , \25674 , \25675 );
nand \U$25334 ( \25677 , \25673 , \25676 );
nand \U$25335 ( \25678 , \25677 , \16271 );
nand \U$25336 ( \25679 , \25670 , \25678 );
not \U$25337 ( \25680 , \25679 );
not \U$25338 ( \25681 , \25680 );
and \U$25339 ( \25682 , \21882 , \12596 );
not \U$25340 ( \25683 , \21882 );
and \U$25341 ( \25684 , \25683 , \4028 );
nor \U$25342 ( \25685 , \25682 , \25684 );
not \U$25343 ( \25686 , \25685 );
not \U$25344 ( \25687 , \12692 );
not \U$25345 ( \25688 , \25687 );
and \U$25346 ( \25689 , \25686 , \25688 );
not \U$25347 ( \25690 , \12774 );
and \U$25348 ( \25691 , RIbb2dea0_51, \13731 );
not \U$25349 ( \25692 , RIbb2dea0_51);
and \U$25350 ( \25693 , \25692 , \3275 );
nor \U$25351 ( \25694 , \25691 , \25693 );
nor \U$25352 ( \25695 , \25690 , \25694 );
nor \U$25353 ( \25696 , \25689 , \25695 );
not \U$25354 ( \25697 , \25696 );
or \U$25355 ( \25698 , \25681 , \25697 );
not \U$25356 ( \25699 , \14930 );
not \U$25357 ( \25700 , RIbb2ddb0_53);
not \U$25358 ( \25701 , \7018 );
or \U$25359 ( \25702 , \25700 , \25701 );
not \U$25360 ( \25703 , \16898 );
nand \U$25361 ( \25704 , \25703 , \13463 );
nand \U$25362 ( \25705 , \25702 , \25704 );
not \U$25363 ( \25706 , \25705 );
or \U$25364 ( \25707 , \25699 , \25706 );
not \U$25365 ( \25708 , RIbb2ddb0_53);
not \U$25366 ( \25709 , \3023 );
or \U$25367 ( \25710 , \25708 , \25709 );
nand \U$25368 ( \25711 , \8491 , \13463 );
nand \U$25369 ( \25712 , \25710 , \25711 );
nand \U$25370 ( \25713 , \25712 , \17563 );
nand \U$25371 ( \25714 , \25707 , \25713 );
nand \U$25372 ( \25715 , \25698 , \25714 );
not \U$25373 ( \25716 , \25696 );
nand \U$25374 ( \25717 , \25716 , \25679 );
nand \U$25375 ( \25718 , \25715 , \25717 );
xor \U$25376 ( \25719 , \25663 , \25718 );
not \U$25377 ( \25720 , \5845 );
not \U$25378 ( \25721 , RIbb2e620_35);
not \U$25379 ( \25722 , \18802 );
or \U$25380 ( \25723 , \25721 , \25722 );
nand \U$25381 ( \25724 , \13526 , \6002 );
nand \U$25382 ( \25725 , \25723 , \25724 );
not \U$25383 ( \25726 , \25725 );
or \U$25384 ( \25727 , \25720 , \25726 );
not \U$25385 ( \25728 , RIbb2e620_35);
not \U$25386 ( \25729 , \12260 );
or \U$25387 ( \25730 , \25728 , \25729 );
nand \U$25388 ( \25731 , \12755 , \3866 );
nand \U$25389 ( \25732 , \25730 , \25731 );
nand \U$25390 ( \25733 , \25732 , \4712 );
nand \U$25391 ( \25734 , \25727 , \25733 );
not \U$25392 ( \25735 , \12169 );
not \U$25393 ( \25736 , RIbb2df90_49);
not \U$25394 ( \25737 , \4752 );
or \U$25395 ( \25738 , \25736 , \25737 );
nand \U$25396 ( \25739 , \3089 , \12278 );
nand \U$25397 ( \25740 , \25738 , \25739 );
not \U$25398 ( \25741 , \25740 );
or \U$25399 ( \25742 , \25735 , \25741 );
not \U$25400 ( \25743 , RIbb2df90_49);
not \U$25401 ( \25744 , \13756 );
or \U$25402 ( \25745 , \25743 , \25744 );
not \U$25403 ( \25746 , RIbb2df90_49);
nand \U$25404 ( \25747 , \25746 , \4086 );
nand \U$25405 ( \25748 , \25745 , \25747 );
nand \U$25406 ( \25749 , \25748 , \12167 );
nand \U$25407 ( \25750 , \25742 , \25749 );
xor \U$25408 ( \25751 , \25734 , \25750 );
not \U$25409 ( \25752 , \16533 );
not \U$25410 ( \25753 , RIbb2d9f0_61);
not \U$25411 ( \25754 , \1853 );
or \U$25412 ( \25755 , \25753 , \25754 );
nand \U$25413 ( \25756 , \4610 , \19746 );
nand \U$25414 ( \25757 , \25755 , \25756 );
not \U$25415 ( \25758 , \25757 );
or \U$25416 ( \25759 , \25752 , \25758 );
not \U$25417 ( \25760 , RIbb2d9f0_61);
not \U$25418 ( \25761 , \4449 );
or \U$25419 ( \25762 , \25760 , \25761 );
nand \U$25420 ( \25763 , \16235 , \19746 );
nand \U$25421 ( \25764 , \25762 , \25763 );
nand \U$25422 ( \25765 , \25764 , \18717 );
nand \U$25423 ( \25766 , \25759 , \25765 );
and \U$25424 ( \25767 , \25751 , \25766 );
and \U$25425 ( \25768 , \25734 , \25750 );
or \U$25426 ( \25769 , \25767 , \25768 );
xor \U$25427 ( \25770 , \25719 , \25769 );
not \U$25428 ( \25771 , \823 );
not \U$25429 ( \25772 , \1776 );
or \U$25430 ( \25773 , \25771 , \25772 );
nand \U$25431 ( \25774 , \25773 , \19064 );
and \U$25432 ( \25775 , RIbb2ee18_18, RIbb2eda0_19);
nor \U$25433 ( \25776 , \25775 , \3057 );
and \U$25434 ( \25777 , \25774 , \25776 );
not \U$25435 ( \25778 , \835 );
not \U$25436 ( \25779 , RIbb2ee90_17);
not \U$25437 ( \25780 , \17744 );
or \U$25438 ( \25781 , \25779 , \25780 );
nand \U$25439 ( \25782 , \17517 , \3057 );
nand \U$25440 ( \25783 , \25781 , \25782 );
not \U$25441 ( \25784 , \25783 );
or \U$25442 ( \25785 , \25778 , \25784 );
and \U$25443 ( \25786 , RIbb2ee90_17, \17506 );
not \U$25444 ( \25787 , RIbb2ee90_17);
and \U$25445 ( \25788 , \25787 , \19063 );
nor \U$25446 ( \25789 , \25786 , \25788 );
nand \U$25447 ( \25790 , \25789 , \830 );
nand \U$25448 ( \25791 , \25785 , \25790 );
xor \U$25449 ( \25792 , \25777 , \25791 );
not \U$25450 ( \25793 , \854 );
not \U$25451 ( \25794 , RIbb2eda0_19);
not \U$25452 ( \25795 , \17755 );
or \U$25453 ( \25796 , \25794 , \25795 );
nand \U$25454 ( \25797 , \1776 , \18923 );
nand \U$25455 ( \25798 , \25796 , \25797 );
not \U$25456 ( \25799 , \25798 );
or \U$25457 ( \25800 , \25793 , \25799 );
not \U$25458 ( \25801 , RIbb2eda0_19);
not \U$25459 ( \25802 , \16820 );
or \U$25460 ( \25803 , \25801 , \25802 );
nand \U$25461 ( \25804 , \17529 , \1776 );
nand \U$25462 ( \25805 , \25803 , \25804 );
nand \U$25463 ( \25806 , \25805 , \853 );
nand \U$25464 ( \25807 , \25800 , \25806 );
xor \U$25465 ( \25808 , \25792 , \25807 );
not \U$25466 ( \25809 , \3382 );
not \U$25467 ( \25810 , RIbb2ebc0_23);
not \U$25468 ( \25811 , \16844 );
or \U$25469 ( \25812 , \25810 , \25811 );
nand \U$25470 ( \25813 , \16575 , \3401 );
nand \U$25471 ( \25814 , \25812 , \25813 );
not \U$25472 ( \25815 , \25814 );
or \U$25473 ( \25816 , \25809 , \25815 );
not \U$25474 ( \25817 , RIbb2ebc0_23);
not \U$25475 ( \25818 , \16747 );
or \U$25476 ( \25819 , \25817 , \25818 );
nand \U$25477 ( \25820 , \16856 , \3396 );
nand \U$25478 ( \25821 , \25819 , \25820 );
not \U$25479 ( \25822 , \16947 );
nand \U$25480 ( \25823 , \25821 , \25822 );
nand \U$25481 ( \25824 , \25816 , \25823 );
and \U$25482 ( \25825 , \25808 , \25824 );
and \U$25483 ( \25826 , \25792 , \25807 );
or \U$25484 ( \25827 , \25825 , \25826 );
not \U$25485 ( \25828 , \7103 );
and \U$25486 ( \25829 , RIbb2e440_39, \23529 );
not \U$25487 ( \25830 , RIbb2e440_39);
and \U$25488 ( \25831 , \25830 , \13866 );
or \U$25489 ( \25832 , \25829 , \25831 );
not \U$25490 ( \25833 , \25832 );
or \U$25491 ( \25834 , \25828 , \25833 );
and \U$25492 ( \25835 , RIbb2e440_39, \20692 );
not \U$25493 ( \25836 , RIbb2e440_39);
and \U$25494 ( \25837 , \25836 , \14024 );
or \U$25495 ( \25838 , \25835 , \25837 );
nand \U$25496 ( \25839 , \25838 , \7104 );
nand \U$25497 ( \25840 , \25834 , \25839 );
xor \U$25498 ( \25841 , \25827 , \25840 );
not \U$25499 ( \25842 , \8353 );
not \U$25500 ( \25843 , RIbb2e350_41);
not \U$25501 ( \25844 , \19868 );
not \U$25502 ( \25845 , \25844 );
not \U$25503 ( \25846 , \25845 );
or \U$25504 ( \25847 , \25843 , \25846 );
nand \U$25505 ( \25848 , \11534 , \8357 );
nand \U$25506 ( \25849 , \25847 , \25848 );
not \U$25507 ( \25850 , \25849 );
or \U$25508 ( \25851 , \25842 , \25850 );
not \U$25509 ( \25852 , RIbb2e350_41);
not \U$25510 ( \25853 , \13853 );
or \U$25511 ( \25854 , \25852 , \25853 );
nand \U$25512 ( \25855 , \14673 , \7097 );
nand \U$25513 ( \25856 , \25854 , \25855 );
nand \U$25514 ( \25857 , \25856 , \8362 );
nand \U$25515 ( \25858 , \25851 , \25857 );
xnor \U$25516 ( \25859 , \25841 , \25858 );
not \U$25517 ( \25860 , \25859 );
not \U$25518 ( \25861 , \10119 );
not \U$25519 ( \25862 , RIbb2e170_45);
not \U$25520 ( \25863 , \9021 );
or \U$25521 ( \25864 , \25862 , \25863 );
nand \U$25522 ( \25865 , \9020 , \9094 );
nand \U$25523 ( \25866 , \25864 , \25865 );
not \U$25524 ( \25867 , \25866 );
or \U$25525 ( \25868 , \25861 , \25867 );
not \U$25526 ( \25869 , RIbb2e170_45);
not \U$25527 ( \25870 , \9108 );
or \U$25528 ( \25871 , \25869 , \25870 );
nand \U$25529 ( \25872 , \6229 , \13372 );
nand \U$25530 ( \25873 , \25871 , \25872 );
nand \U$25531 ( \25874 , \25873 , \10117 );
nand \U$25532 ( \25875 , \25868 , \25874 );
not \U$25533 ( \25876 , \9098 );
not \U$25534 ( \25877 , RIbb2e260_43);
not \U$25535 ( \25878 , \8338 );
or \U$25536 ( \25879 , \25877 , \25878 );
nand \U$25537 ( \25880 , \15796 , \10444 );
nand \U$25538 ( \25881 , \25879 , \25880 );
not \U$25539 ( \25882 , \25881 );
or \U$25540 ( \25883 , \25876 , \25882 );
not \U$25541 ( \25884 , RIbb2e260_43);
not \U$25542 ( \25885 , \14041 );
or \U$25543 ( \25886 , \25884 , \25885 );
nand \U$25544 ( \25887 , \7308 , \8347 );
nand \U$25545 ( \25888 , \25886 , \25887 );
nand \U$25546 ( \25889 , \25888 , \10451 );
nand \U$25547 ( \25890 , \25883 , \25889 );
xor \U$25548 ( \25891 , \25875 , \25890 );
not \U$25549 ( \25892 , \11177 );
not \U$25550 ( \25893 , RIbb2e080_47);
not \U$25551 ( \25894 , \13552 );
or \U$25552 ( \25895 , \25893 , \25894 );
nand \U$25553 ( \25896 , \4086 , \10113 );
nand \U$25554 ( \25897 , \25895 , \25896 );
not \U$25555 ( \25898 , \25897 );
or \U$25556 ( \25899 , \25892 , \25898 );
not \U$25557 ( \25900 , RIbb2e080_47);
not \U$25558 ( \25901 , \13560 );
or \U$25559 ( \25902 , \25900 , \25901 );
nand \U$25560 ( \25903 , \4391 , \12971 );
nand \U$25561 ( \25904 , \25902 , \25903 );
nand \U$25562 ( \25905 , \25904 , \11176 );
nand \U$25563 ( \25906 , \25899 , \25905 );
xor \U$25564 ( \25907 , \25891 , \25906 );
not \U$25565 ( \25908 , \25907 );
or \U$25566 ( \25909 , \25860 , \25908 );
or \U$25567 ( \25910 , \25907 , \25859 );
nand \U$25568 ( \25911 , \25909 , \25910 );
not \U$25569 ( \25912 , \4712 );
not \U$25570 ( \25913 , \25725 );
or \U$25571 ( \25914 , \25912 , \25913 );
not \U$25572 ( \25915 , RIbb2e620_35);
not \U$25573 ( \25916 , \15106 );
or \U$25574 ( \25917 , \25915 , \25916 );
nand \U$25575 ( \25918 , \10301 , \3866 );
nand \U$25576 ( \25919 , \25917 , \25918 );
nand \U$25577 ( \25920 , \25919 , \4714 );
nand \U$25578 ( \25921 , \25914 , \25920 );
not \U$25579 ( \25922 , \6241 );
not \U$25580 ( \25923 , RIbb2e530_37);
not \U$25581 ( \25924 , \18578 );
or \U$25582 ( \25925 , \25923 , \25924 );
nand \U$25583 ( \25926 , \9278 , \4708 );
nand \U$25584 ( \25927 , \25925 , \25926 );
not \U$25585 ( \25928 , \25927 );
or \U$25586 ( \25929 , \25922 , \25928 );
not \U$25587 ( \25930 , \6252 );
not \U$25588 ( \25931 , RIbb2e530_37);
not \U$25589 ( \25932 , \20044 );
or \U$25590 ( \25933 , \25931 , \25932 );
nand \U$25591 ( \25934 , \20045 , \6246 );
nand \U$25592 ( \25935 , \25933 , \25934 );
nand \U$25593 ( \25936 , \25930 , \25935 );
nand \U$25594 ( \25937 , \25929 , \25936 );
not \U$25595 ( \25938 , \25937 );
xor \U$25596 ( \25939 , \25921 , \25938 );
not \U$25597 ( \25940 , \14752 );
not \U$25598 ( \25941 , RIbb2df90_49);
buf \U$25599 ( \25942 , \3001 );
not \U$25600 ( \25943 , \25942 );
or \U$25601 ( \25944 , \25941 , \25943 );
nand \U$25602 ( \25945 , \3002 , \12278 );
nand \U$25603 ( \25946 , \25944 , \25945 );
not \U$25604 ( \25947 , \25946 );
or \U$25605 ( \25948 , \25940 , \25947 );
nand \U$25606 ( \25949 , \25740 , \13295 );
nand \U$25607 ( \25950 , \25948 , \25949 );
xor \U$25608 ( \25951 , \25939 , \25950 );
not \U$25609 ( \25952 , \25951 );
and \U$25610 ( \25953 , \25911 , \25952 );
not \U$25611 ( \25954 , \25911 );
and \U$25612 ( \25955 , \25954 , \25951 );
nor \U$25613 ( \25956 , \25953 , \25955 );
not \U$25614 ( \25957 , \25956 );
and \U$25615 ( \25958 , \25770 , \25957 );
not \U$25616 ( \25959 , \25770 );
and \U$25617 ( \25960 , \25959 , \25956 );
nor \U$25618 ( \25961 , \25958 , \25960 );
xor \U$25619 ( \25962 , \25734 , \25750 );
xor \U$25620 ( \25963 , \25962 , \25766 );
not \U$25621 ( \25964 , \2940 );
not \U$25622 ( \25965 , RIbb2e800_31);
not \U$25623 ( \25966 , \17315 );
or \U$25624 ( \25967 , \25965 , \25966 );
nand \U$25625 ( \25968 , \13989 , \2917 );
nand \U$25626 ( \25969 , \25967 , \25968 );
not \U$25627 ( \25970 , \25969 );
or \U$25628 ( \25971 , \25964 , \25970 );
not \U$25629 ( \25972 , RIbb2e800_31);
not \U$25630 ( \25973 , \14624 );
or \U$25631 ( \25974 , \25972 , \25973 );
nand \U$25632 ( \25975 , \13474 , \8810 );
nand \U$25633 ( \25976 , \25974 , \25975 );
nand \U$25634 ( \25977 , \25976 , \3613 );
nand \U$25635 ( \25978 , \25971 , \25977 );
not \U$25636 ( \25979 , \25978 );
not \U$25637 ( \25980 , \3886 );
not \U$25638 ( \25981 , RIbb2e710_33);
not \U$25639 ( \25982 , \14840 );
or \U$25640 ( \25983 , \25981 , \25982 );
not \U$25641 ( \25984 , \21756 );
nand \U$25642 ( \25985 , \25984 , \2935 );
nand \U$25643 ( \25986 , \25983 , \25985 );
not \U$25644 ( \25987 , \25986 );
or \U$25645 ( \25988 , \25980 , \25987 );
not \U$25646 ( \25989 , RIbb2e710_33);
not \U$25647 ( \25990 , \12323 );
or \U$25648 ( \25991 , \25989 , \25990 );
nand \U$25649 ( \25992 , \12933 , \6058 );
nand \U$25650 ( \25993 , \25991 , \25992 );
nand \U$25651 ( \25994 , \25993 , \4791 );
nand \U$25652 ( \25995 , \25988 , \25994 );
not \U$25653 ( \25996 , \25995 );
or \U$25654 ( \25997 , \25979 , \25996 );
or \U$25655 ( \25998 , \25995 , \25978 );
not \U$25656 ( \25999 , \3465 );
not \U$25657 ( \26000 , RIbb2e9e0_27);
not \U$25658 ( \26001 , \15469 );
or \U$25659 ( \26002 , \26000 , \26001 );
nand \U$25660 ( \26003 , \15030 , \3454 );
nand \U$25661 ( \26004 , \26002 , \26003 );
not \U$25662 ( \26005 , \26004 );
or \U$25663 ( \26006 , \25999 , \26005 );
not \U$25664 ( \26007 , RIbb2e9e0_27);
not \U$25665 ( \26008 , \16561 );
or \U$25666 ( \26009 , \26007 , \26008 );
not \U$25667 ( \26010 , RIbb2e9e0_27);
nand \U$25668 ( \26011 , \26010 , \16562 );
nand \U$25669 ( \26012 , \26009 , \26011 );
nand \U$25670 ( \26013 , \26012 , \3445 );
nand \U$25671 ( \26014 , \26006 , \26013 );
nand \U$25672 ( \26015 , \25998 , \26014 );
nand \U$25673 ( \26016 , \25997 , \26015 );
not \U$25674 ( \26017 , \26016 );
not \U$25675 ( \26018 , \12692 );
not \U$25676 ( \26019 , \25694 );
not \U$25677 ( \26020 , \26019 );
or \U$25678 ( \26021 , \26018 , \26020 );
and \U$25679 ( \26022 , RIbb2dea0_51, \4749 );
not \U$25680 ( \26023 , RIbb2dea0_51);
and \U$25681 ( \26024 , \26023 , \10458 );
or \U$25682 ( \26025 , \26022 , \26024 );
nand \U$25683 ( \26026 , \26025 , \12774 );
nand \U$25684 ( \26027 , \26021 , \26026 );
not \U$25685 ( \26028 , \26027 );
or \U$25686 ( \26029 , \26017 , \26028 );
or \U$25687 ( \26030 , \26027 , \26016 );
not \U$25688 ( \26031 , \3381 );
not \U$25689 ( \26032 , RIbb2ebc0_23);
not \U$25690 ( \26033 , \23185 );
or \U$25691 ( \26034 , \26032 , \26033 );
nand \U$25692 ( \26035 , \16829 , \3388 );
nand \U$25693 ( \26036 , \26034 , \26035 );
not \U$25694 ( \26037 , \26036 );
or \U$25695 ( \26038 , \26031 , \26037 );
not \U$25696 ( \26039 , \16710 );
and \U$25697 ( \26040 , \3388 , \26039 );
not \U$25698 ( \26041 , \3388 );
and \U$25699 ( \26042 , \26041 , \16710 );
nor \U$25700 ( \26043 , \26040 , \26042 );
not \U$25701 ( \26044 , \26043 );
nand \U$25702 ( \26045 , \26044 , \25822 );
nand \U$25703 ( \26046 , \26038 , \26045 );
and \U$25704 ( \26047 , \17506 , \854 );
not \U$25705 ( \26048 , \2078 );
not \U$25706 ( \26049 , RIbb2ecb0_21);
not \U$25707 ( \26050 , \17529 );
not \U$25708 ( \26051 , \26050 );
or \U$25709 ( \26052 , \26049 , \26051 );
nand \U$25710 ( \26053 , \17529 , \849 );
nand \U$25711 ( \26054 , \26052 , \26053 );
not \U$25712 ( \26055 , \26054 );
or \U$25713 ( \26056 , \26048 , \26055 );
not \U$25714 ( \26057 , RIbb2ecb0_21);
not \U$25715 ( \26058 , \17745 );
or \U$25716 ( \26059 , \26057 , \26058 );
nand \U$25717 ( \26060 , \17517 , \2249 );
nand \U$25718 ( \26061 , \26059 , \26060 );
nand \U$25719 ( \26062 , \26061 , \2077 );
nand \U$25720 ( \26063 , \26056 , \26062 );
xor \U$25721 ( \26064 , \26047 , \26063 );
not \U$25722 ( \26065 , \3406 );
not \U$25723 ( \26066 , RIbb2ebc0_23);
not \U$25724 ( \26067 , \18924 );
or \U$25725 ( \26068 , \26066 , \26067 );
nand \U$25726 ( \26069 , \16704 , \3388 );
nand \U$25727 ( \26070 , \26068 , \26069 );
not \U$25728 ( \26071 , \26070 );
or \U$25729 ( \26072 , \26065 , \26071 );
not \U$25730 ( \26073 , \3381 );
or \U$25731 ( \26074 , \26043 , \26073 );
nand \U$25732 ( \26075 , \26072 , \26074 );
and \U$25733 ( \26076 , \26064 , \26075 );
and \U$25734 ( \26077 , \26047 , \26063 );
or \U$25735 ( \26078 , \26076 , \26077 );
xor \U$25736 ( \26079 , \26046 , \26078 );
not \U$25737 ( \26080 , \2925 );
not \U$25738 ( \26081 , RIbb2e8f0_29);
not \U$25739 ( \26082 , \13978 );
or \U$25740 ( \26083 , \26081 , \26082 );
nand \U$25741 ( \26084 , \16320 , \6970 );
nand \U$25742 ( \26085 , \26083 , \26084 );
not \U$25743 ( \26086 , \26085 );
or \U$25744 ( \26087 , \26080 , \26086 );
not \U$25745 ( \26088 , RIbb2e8f0_29);
not \U$25746 ( \26089 , \20577 );
or \U$25747 ( \26090 , \26088 , \26089 );
nand \U$25748 ( \26091 , \14526 , \2911 );
nand \U$25749 ( \26092 , \26090 , \26091 );
nand \U$25750 ( \26093 , \26092 , \2921 );
nand \U$25751 ( \26094 , \26087 , \26093 );
and \U$25752 ( \26095 , \26079 , \26094 );
and \U$25753 ( \26096 , \26046 , \26078 );
or \U$25754 ( \26097 , \26095 , \26096 );
nand \U$25755 ( \26098 , \26030 , \26097 );
nand \U$25756 ( \26099 , \26029 , \26098 );
xor \U$25757 ( \26100 , \25963 , \26099 );
xor \U$25758 ( \26101 , \25696 , \25714 );
xor \U$25759 ( \26102 , \26101 , \25680 );
and \U$25760 ( \26103 , \26100 , \26102 );
and \U$25761 ( \26104 , \25963 , \26099 );
or \U$25762 ( \26105 , \26103 , \26104 );
not \U$25763 ( \26106 , \26105 );
and \U$25764 ( \26107 , \25961 , \26106 );
not \U$25765 ( \26108 , \25961 );
and \U$25766 ( \26109 , \26108 , \26105 );
nor \U$25767 ( \26110 , \26107 , \26109 );
not \U$25768 ( \26111 , \16271 );
and \U$25769 ( \26112 , RIbb2dae0_59, \6107 );
not \U$25770 ( \26113 , RIbb2dae0_59);
and \U$25771 ( \26114 , \26113 , \3951 );
or \U$25772 ( \26115 , \26112 , \26114 );
not \U$25773 ( \26116 , \26115 );
or \U$25774 ( \26117 , \26111 , \26116 );
nand \U$25775 ( \26118 , \25677 , \17470 );
nand \U$25776 ( \26119 , \26117 , \26118 );
or \U$25777 ( \26120 , RIbb2ed28_20, RIbb2ecb0_21);
nand \U$25778 ( \26121 , \26120 , \17506 );
and \U$25779 ( \26122 , RIbb2ed28_20, RIbb2ecb0_21);
nor \U$25780 ( \26123 , \26122 , \5277 );
and \U$25781 ( \26124 , \26121 , \26123 );
not \U$25782 ( \26125 , \854 );
not \U$25783 ( \26126 , RIbb2eda0_19);
not \U$25784 ( \26127 , \17745 );
or \U$25785 ( \26128 , \26126 , \26127 );
buf \U$25786 ( \26129 , \17516 );
nand \U$25787 ( \26130 , \26129 , \843 );
nand \U$25788 ( \26131 , \26128 , \26130 );
not \U$25789 ( \26132 , \26131 );
or \U$25790 ( \26133 , \26125 , \26132 );
and \U$25791 ( \26134 , RIbb2eda0_19, \17506 );
not \U$25792 ( \26135 , RIbb2eda0_19);
and \U$25793 ( \26136 , \26135 , \20747 );
nor \U$25794 ( \26137 , \26134 , \26136 );
nand \U$25795 ( \26138 , \26137 , \852 );
nand \U$25796 ( \26139 , \26133 , \26138 );
and \U$25797 ( \26140 , \26124 , \26139 );
not \U$25798 ( \26141 , \3382 );
not \U$25799 ( \26142 , \25821 );
or \U$25800 ( \26143 , \26141 , \26142 );
nand \U$25801 ( \26144 , \26036 , \3406 );
nand \U$25802 ( \26145 , \26143 , \26144 );
xor \U$25803 ( \26146 , \26140 , \26145 );
not \U$25804 ( \26147 , \2963 );
not \U$25805 ( \26148 , RIbb2ead0_25);
not \U$25806 ( \26149 , \15755 );
or \U$25807 ( \26150 , \26148 , \26149 );
not \U$25808 ( \26151 , RIbb2ead0_25);
nand \U$25809 ( \26152 , \26151 , \15753 );
nand \U$25810 ( \26153 , \26150 , \26152 );
not \U$25811 ( \26154 , \26153 );
or \U$25812 ( \26155 , \26147 , \26154 );
and \U$25813 ( \26156 , RIbb2ead0_25, \16844 );
not \U$25814 ( \26157 , RIbb2ead0_25);
and \U$25815 ( \26158 , \26157 , \16575 );
or \U$25816 ( \26159 , \26156 , \26158 );
nand \U$25817 ( \26160 , \26159 , \2980 );
nand \U$25818 ( \26161 , \26155 , \26160 );
xnor \U$25819 ( \26162 , \26146 , \26161 );
xor \U$25820 ( \26163 , \26119 , \26162 );
not \U$25821 ( \26164 , \13467 );
not \U$25822 ( \26165 , RIbb2ddb0_53);
not \U$25823 ( \26166 , \13738 );
or \U$25824 ( \26167 , \26165 , \26166 );
nand \U$25825 ( \26168 , \16185 , \13463 );
nand \U$25826 ( \26169 , \26167 , \26168 );
not \U$25827 ( \26170 , \26169 );
or \U$25828 ( \26171 , \26164 , \26170 );
nand \U$25829 ( \26172 , \25712 , \14930 );
nand \U$25830 ( \26173 , \26171 , \26172 );
xor \U$25831 ( \26174 , \26163 , \26173 );
not \U$25832 ( \26175 , \26174 );
xor \U$25833 ( \26176 , \26097 , \26016 );
xnor \U$25834 ( \26177 , \26176 , \26027 );
not \U$25835 ( \26178 , \26177 );
or \U$25836 ( \26179 , \26175 , \26178 );
xor \U$25837 ( \26180 , \26047 , \26063 );
xor \U$25838 ( \26181 , \26180 , \26075 );
not \U$25839 ( \26182 , \3613 );
not \U$25840 ( \26183 , \25969 );
or \U$25841 ( \26184 , \26182 , \26183 );
not \U$25842 ( \26185 , RIbb2e800_31);
not \U$25843 ( \26186 , \14503 );
or \U$25844 ( \26187 , \26185 , \26186 );
nand \U$25845 ( \26188 , \16320 , \9169 );
nand \U$25846 ( \26189 , \26187 , \26188 );
nand \U$25847 ( \26190 , \26189 , \2939 );
nand \U$25848 ( \26191 , \26184 , \26190 );
xor \U$25849 ( \26192 , \26181 , \26191 );
not \U$25850 ( \26193 , \4075 );
not \U$25851 ( \26194 , \25986 );
or \U$25852 ( \26195 , \26193 , \26194 );
not \U$25853 ( \26196 , RIbb2e710_33);
not \U$25854 ( \26197 , \13475 );
or \U$25855 ( \26198 , \26196 , \26197 );
nand \U$25856 ( \26199 , \13474 , \2935 );
nand \U$25857 ( \26200 , \26198 , \26199 );
nand \U$25858 ( \26201 , \26200 , \3886 );
nand \U$25859 ( \26202 , \26195 , \26201 );
and \U$25860 ( \26203 , \26192 , \26202 );
and \U$25861 ( \26204 , \26181 , \26191 );
or \U$25862 ( \26205 , \26203 , \26204 );
xor \U$25863 ( \26206 , \25978 , \26014 );
and \U$25864 ( \26207 , \26206 , \25995 );
not \U$25865 ( \26208 , \26206 );
not \U$25866 ( \26209 , \25995 );
and \U$25867 ( \26210 , \26208 , \26209 );
nor \U$25868 ( \26211 , \26207 , \26210 );
xor \U$25869 ( \26212 , \26205 , \26211 );
not \U$25870 ( \26213 , \12965 );
not \U$25871 ( \26214 , RIbb2e080_47);
not \U$25872 ( \26215 , \21570 );
or \U$25873 ( \26216 , \26214 , \26215 );
nand \U$25874 ( \26217 , \7308 , \15632 );
nand \U$25875 ( \26218 , \26216 , \26217 );
not \U$25876 ( \26219 , \26218 );
or \U$25877 ( \26220 , \26213 , \26219 );
not \U$25878 ( \26221 , RIbb2e080_47);
not \U$25879 ( \26222 , \13875 );
or \U$25880 ( \26223 , \26221 , \26222 );
nand \U$25881 ( \26224 , \6603 , \16163 );
nand \U$25882 ( \26225 , \26223 , \26224 );
nand \U$25883 ( \26226 , \26225 , \11176 );
nand \U$25884 ( \26227 , \26220 , \26226 );
not \U$25885 ( \26228 , \10119 );
not \U$25886 ( \26229 , RIbb2e170_45);
not \U$25887 ( \26230 , \19869 );
or \U$25888 ( \26231 , \26229 , \26230 );
not \U$25889 ( \26232 , \15066 );
nand \U$25890 ( \26233 , \26232 , \11065 );
nand \U$25891 ( \26234 , \26231 , \26233 );
not \U$25892 ( \26235 , \26234 );
or \U$25893 ( \26236 , \26228 , \26235 );
not \U$25894 ( \26237 , RIbb2e170_45);
not \U$25895 ( \26238 , \9070 );
or \U$25896 ( \26239 , \26237 , \26238 );
nand \U$25897 ( \26240 , \7296 , \9094 );
nand \U$25898 ( \26241 , \26239 , \26240 );
nand \U$25899 ( \26242 , \26241 , \10599 );
nand \U$25900 ( \26243 , \26236 , \26242 );
buf \U$25901 ( \26244 , \26243 );
nor \U$25902 ( \26245 , \26227 , \26244 );
not \U$25903 ( \26246 , RIbb2e260_43);
not \U$25904 ( \26247 , \8319 );
or \U$25905 ( \26248 , \26246 , \26247 );
nand \U$25906 ( \26249 , \14024 , \10444 );
nand \U$25907 ( \26250 , \26248 , \26249 );
and \U$25908 ( \26251 , \9099 , \26250 );
not \U$25909 ( \26252 , RIbb2e260_43);
not \U$25910 ( \26253 , \13863 );
or \U$25911 ( \26254 , \26252 , \26253 );
not \U$25912 ( \26255 , RIbb2e260_43);
nand \U$25913 ( \26256 , \13866 , \26255 );
nand \U$25914 ( \26257 , \26254 , \26256 );
and \U$25915 ( \26258 , \26257 , \9098 );
nor \U$25916 ( \26259 , \26251 , \26258 );
or \U$25917 ( \26260 , \26245 , \26259 );
nand \U$25918 ( \26261 , \26227 , \26244 );
nand \U$25919 ( \26262 , \26260 , \26261 );
and \U$25920 ( \26263 , \26212 , \26262 );
and \U$25921 ( \26264 , \26205 , \26211 );
or \U$25922 ( \26265 , \26263 , \26264 );
nand \U$25923 ( \26266 , \26179 , \26265 );
not \U$25924 ( \26267 , \26177 );
not \U$25925 ( \26268 , \26174 );
nand \U$25926 ( \26269 , \26267 , \26268 );
nand \U$25927 ( \26270 , \26266 , \26269 );
xor \U$25928 ( \26271 , \25963 , \26099 );
xor \U$25929 ( \26272 , \26271 , \26102 );
xor \U$25930 ( \26273 , \26270 , \26272 );
not \U$25931 ( \26274 , \16674 );
not \U$25932 ( \26275 , RIbb2dbd0_57);
not \U$25933 ( \26276 , \21490 );
or \U$25934 ( \26277 , \26275 , \26276 );
not \U$25935 ( \26278 , RIbb2dbd0_57);
nand \U$25936 ( \26279 , \26278 , \3653 );
nand \U$25937 ( \26280 , \26277 , \26279 );
not \U$25938 ( \26281 , \26280 );
or \U$25939 ( \26282 , \26274 , \26281 );
not \U$25940 ( \26283 , RIbb2dbd0_57);
not \U$25941 ( \26284 , \6172 );
or \U$25942 ( \26285 , \26283 , \26284 );
not \U$25943 ( \26286 , RIbb2dbd0_57);
nand \U$25944 ( \26287 , \26286 , \3224 );
nand \U$25945 ( \26288 , \26285 , \26287 );
nand \U$25946 ( \26289 , \26288 , \17100 );
nand \U$25947 ( \26290 , \26282 , \26289 );
buf \U$25948 ( \26291 , \26290 );
not \U$25949 ( \26292 , \26291 );
not \U$25950 ( \26293 , \8353 );
not \U$25951 ( \26294 , RIbb2e350_41);
not \U$25952 ( \26295 , \13916 );
or \U$25953 ( \26296 , \26294 , \26295 );
nand \U$25954 ( \26297 , \13920 , \13400 );
nand \U$25955 ( \26298 , \26296 , \26297 );
not \U$25956 ( \26299 , \26298 );
or \U$25957 ( \26300 , \26293 , \26299 );
not \U$25958 ( \26301 , RIbb2e350_41);
not \U$25959 ( \26302 , \10306 );
or \U$25960 ( \26303 , \26301 , \26302 );
nand \U$25961 ( \26304 , \9841 , \8357 );
nand \U$25962 ( \26305 , \26303 , \26304 );
nand \U$25963 ( \26306 , \26305 , \8362 );
nand \U$25964 ( \26307 , \26300 , \26306 );
not \U$25965 ( \26308 , \26307 );
or \U$25966 ( \26309 , \26292 , \26308 );
not \U$25967 ( \26310 , \26307 );
not \U$25968 ( \26311 , \26310 );
not \U$25969 ( \26312 , \26290 );
not \U$25970 ( \26313 , \26312 );
or \U$25971 ( \26314 , \26311 , \26313 );
not \U$25972 ( \26315 , \6251 );
not \U$25973 ( \26316 , RIbb2e530_37);
not \U$25974 ( \26317 , \11580 );
or \U$25975 ( \26318 , \26316 , \26317 );
nand \U$25976 ( \26319 , \14885 , \7473 );
nand \U$25977 ( \26320 , \26318 , \26319 );
not \U$25978 ( \26321 , \26320 );
or \U$25979 ( \26322 , \26315 , \26321 );
not \U$25980 ( \26323 , RIbb2e530_37);
not \U$25981 ( \26324 , \12257 );
or \U$25982 ( \26325 , \26323 , \26324 );
nand \U$25983 ( \26326 , \11142 , \8701 );
nand \U$25984 ( \26327 , \26325 , \26326 );
nand \U$25985 ( \26328 , \26327 , \20792 );
nand \U$25986 ( \26329 , \26322 , \26328 );
nand \U$25987 ( \26330 , \26314 , \26329 );
nand \U$25988 ( \26331 , \26309 , \26330 );
not \U$25989 ( \26332 , \26331 );
not \U$25990 ( \26333 , \16271 );
and \U$25991 ( \26334 , RIbb2dae0_59, \4637 );
not \U$25992 ( \26335 , RIbb2dae0_59);
and \U$25993 ( \26336 , \26335 , \14791 );
nor \U$25994 ( \26337 , \26334 , \26336 );
not \U$25995 ( \26338 , \26337 );
or \U$25996 ( \26339 , \26333 , \26338 );
and \U$25997 ( \26340 , RIbb2dae0_59, \15397 );
not \U$25998 ( \26341 , RIbb2dae0_59);
and \U$25999 ( \26342 , \26341 , \3140 );
nor \U$26000 ( \26343 , \26340 , \26342 );
nand \U$26001 ( \26344 , \26343 , \16257 );
nand \U$26002 ( \26345 , \26339 , \26344 );
not \U$26003 ( \26346 , \26345 );
not \U$26004 ( \26347 , \17275 );
not \U$26005 ( \26348 , RIbb2d900_63);
not \U$26006 ( \26349 , \3319 );
or \U$26007 ( \26350 , \26348 , \26349 );
nand \U$26008 ( \26351 , \2222 , \17262 );
nand \U$26009 ( \26352 , \26350 , \26351 );
not \U$26010 ( \26353 , \26352 );
or \U$26011 ( \26354 , \26347 , \26353 );
not \U$26012 ( \26355 , RIbb2d900_63);
not \U$26013 ( \26356 , \3563 );
or \U$26014 ( \26357 , \26355 , \26356 );
nand \U$26015 ( \26358 , \3309 , \17262 );
nand \U$26016 ( \26359 , \26357 , \26358 );
nand \U$26017 ( \26360 , \26359 , RIbb2d888_64);
nand \U$26018 ( \26361 , \26354 , \26360 );
not \U$26019 ( \26362 , \26361 );
or \U$26020 ( \26363 , \26346 , \26362 );
or \U$26021 ( \26364 , \26361 , \26345 );
not \U$26022 ( \26365 , \14930 );
not \U$26023 ( \26366 , RIbb2ddb0_53);
not \U$26024 ( \26367 , \13731 );
or \U$26025 ( \26368 , \26366 , \26367 );
nand \U$26026 ( \26369 , \3002 , \13463 );
nand \U$26027 ( \26370 , \26368 , \26369 );
not \U$26028 ( \26371 , \26370 );
or \U$26029 ( \26372 , \26365 , \26371 );
not \U$26030 ( \26373 , RIbb2ddb0_53);
not \U$26031 ( \26374 , \4748 );
or \U$26032 ( \26375 , \26373 , \26374 );
nand \U$26033 ( \26376 , \3089 , \13463 );
nand \U$26034 ( \26377 , \26375 , \26376 );
nand \U$26035 ( \26378 , \26377 , \17563 );
nand \U$26036 ( \26379 , \26372 , \26378 );
nand \U$26037 ( \26380 , \26364 , \26379 );
nand \U$26038 ( \26381 , \26363 , \26380 );
not \U$26039 ( \26382 , \26381 );
or \U$26040 ( \26383 , \26332 , \26382 );
or \U$26041 ( \26384 , \26381 , \26331 );
xor \U$26042 ( \26385 , \26124 , \26139 );
not \U$26043 ( \26386 , \2078 );
not \U$26044 ( \26387 , RIbb2ecb0_21);
not \U$26045 ( \26388 , \18924 );
or \U$26046 ( \26389 , \26387 , \26388 );
nand \U$26047 ( \26390 , \18920 , \2254 );
nand \U$26048 ( \26391 , \26389 , \26390 );
not \U$26049 ( \26392 , \26391 );
or \U$26050 ( \26393 , \26386 , \26392 );
nand \U$26051 ( \26394 , \26054 , \2077 );
nand \U$26052 ( \26395 , \26393 , \26394 );
xor \U$26053 ( \26396 , \26385 , \26395 );
not \U$26054 ( \26397 , \2963 );
not \U$26055 ( \26398 , \26159 );
or \U$26056 ( \26399 , \26397 , \26398 );
and \U$26057 ( \26400 , RIbb2ead0_25, \16747 );
not \U$26058 ( \26401 , RIbb2ead0_25);
and \U$26059 ( \26402 , \26401 , \19077 );
or \U$26060 ( \26403 , \26400 , \26402 );
nand \U$26061 ( \26404 , \26403 , \2979 );
nand \U$26062 ( \26405 , \26399 , \26404 );
xor \U$26063 ( \26406 , \26396 , \26405 );
not \U$26064 ( \26407 , \8362 );
not \U$26065 ( \26408 , \26298 );
or \U$26066 ( \26409 , \26407 , \26408 );
not \U$26067 ( \26410 , RIbb2e350_41);
not \U$26068 ( \26411 , \13863 );
or \U$26069 ( \26412 , \26410 , \26411 );
nand \U$26070 ( \26413 , \13866 , \9402 );
nand \U$26071 ( \26414 , \26412 , \26413 );
nand \U$26072 ( \26415 , \26414 , \8354 );
nand \U$26073 ( \26416 , \26409 , \26415 );
xor \U$26074 ( \26417 , \26406 , \26416 );
not \U$26075 ( \26418 , \10451 );
not \U$26076 ( \26419 , RIbb2e260_43);
not \U$26077 ( \26420 , \17811 );
or \U$26078 ( \26421 , \26419 , \26420 );
not \U$26079 ( \26422 , \13850 );
nand \U$26080 ( \26423 , \26422 , \9847 );
nand \U$26081 ( \26424 , \26421 , \26423 );
not \U$26082 ( \26425 , \26424 );
or \U$26083 ( \26426 , \26418 , \26425 );
nand \U$26084 ( \26427 , \26250 , \9098 );
nand \U$26085 ( \26428 , \26426 , \26427 );
xor \U$26086 ( \26429 , \26417 , \26428 );
nand \U$26087 ( \26430 , \26384 , \26429 );
nand \U$26088 ( \26431 , \26383 , \26430 );
not \U$26089 ( \26432 , \26431 );
not \U$26090 ( \26433 , \26432 );
not \U$26091 ( \26434 , \11176 );
not \U$26092 ( \26435 , \26218 );
or \U$26093 ( \26436 , \26434 , \26435 );
not \U$26094 ( \26437 , RIbb2e080_47);
not \U$26095 ( \26438 , \17341 );
or \U$26096 ( \26439 , \26437 , \26438 );
nand \U$26097 ( \26440 , \7111 , \12971 );
nand \U$26098 ( \26441 , \26439 , \26440 );
nand \U$26099 ( \26442 , \26441 , \12965 );
nand \U$26100 ( \26443 , \26436 , \26442 );
not \U$26101 ( \26444 , \26443 );
not \U$26102 ( \26445 , \13295 );
not \U$26103 ( \26446 , RIbb2df90_49);
not \U$26104 ( \26447 , \9021 );
or \U$26105 ( \26448 , \26446 , \26447 );
nand \U$26106 ( \26449 , \6198 , \12278 );
nand \U$26107 ( \26450 , \26448 , \26449 );
not \U$26108 ( \26451 , \26450 );
or \U$26109 ( \26452 , \26445 , \26451 );
not \U$26110 ( \26453 , RIbb2df90_49);
not \U$26111 ( \26454 , \13559 );
or \U$26112 ( \26455 , \26453 , \26454 );
nand \U$26113 ( \26456 , \6269 , \12278 );
nand \U$26114 ( \26457 , \26455 , \26456 );
nand \U$26115 ( \26458 , \26457 , \12284 );
nand \U$26116 ( \26459 , \26452 , \26458 );
not \U$26117 ( \26460 , \26459 );
or \U$26118 ( \26461 , \26444 , \26460 );
or \U$26119 ( \26462 , \26459 , \26443 );
not \U$26120 ( \26463 , \10119 );
not \U$26121 ( \26464 , RIbb2e170_45);
not \U$26122 ( \26465 , \8338 );
or \U$26123 ( \26466 , \26464 , \26465 );
not \U$26124 ( \26467 , \8338 );
nand \U$26125 ( \26468 , \26467 , \17970 );
nand \U$26126 ( \26469 , \26466 , \26468 );
not \U$26127 ( \26470 , \26469 );
or \U$26128 ( \26471 , \26463 , \26470 );
nand \U$26129 ( \26472 , \26234 , \10117 );
nand \U$26130 ( \26473 , \26471 , \26472 );
nand \U$26131 ( \26474 , \26462 , \26473 );
nand \U$26132 ( \26475 , \26461 , \26474 );
xor \U$26133 ( \26476 , \26406 , \26416 );
and \U$26134 ( \26477 , \26476 , \26428 );
and \U$26135 ( \26478 , \26406 , \26416 );
or \U$26136 ( \26479 , \26477 , \26478 );
xor \U$26137 ( \26480 , \26475 , \26479 );
not \U$26138 ( \26481 , \17100 );
not \U$26139 ( \26482 , RIbb2dbd0_57);
not \U$26140 ( \26483 , \4638 );
or \U$26141 ( \26484 , \26482 , \26483 );
nand \U$26142 ( \26485 , \3202 , \16671 );
nand \U$26143 ( \26486 , \26484 , \26485 );
not \U$26144 ( \26487 , \26486 );
or \U$26145 ( \26488 , \26481 , \26487 );
nand \U$26146 ( \26489 , \26288 , \19101 );
nand \U$26147 ( \26490 , \26488 , \26489 );
not \U$26148 ( \26491 , \26490 );
not \U$26149 ( \26492 , RIbb2d888_64);
not \U$26150 ( \26493 , RIbb2d900_63);
not \U$26151 ( \26494 , \4609 );
or \U$26152 ( \26495 , \26493 , \26494 );
nand \U$26153 ( \26496 , \1852 , \17262 );
nand \U$26154 ( \26497 , \26495 , \26496 );
not \U$26155 ( \26498 , \26497 );
or \U$26156 ( \26499 , \26492 , \26498 );
nand \U$26157 ( \26500 , \26359 , \17275 );
nand \U$26158 ( \26501 , \26499 , \26500 );
not \U$26159 ( \26502 , \26501 );
or \U$26160 ( \26503 , \26491 , \26502 );
or \U$26161 ( \26504 , \26490 , \26501 );
not \U$26162 ( \26505 , \5845 );
not \U$26163 ( \26506 , RIbb2e620_35);
not \U$26164 ( \26507 , \11580 );
or \U$26165 ( \26508 , \26506 , \26507 );
nand \U$26166 ( \26509 , \22555 , \3866 );
nand \U$26167 ( \26510 , \26508 , \26509 );
not \U$26168 ( \26511 , \26510 );
or \U$26169 ( \26512 , \26505 , \26511 );
not \U$26170 ( \26513 , RIbb2e620_35);
not \U$26171 ( \26514 , \23243 );
or \U$26172 ( \26515 , \26513 , \26514 );
nand \U$26173 ( \26516 , \12174 , \6002 );
nand \U$26174 ( \26517 , \26515 , \26516 );
nand \U$26175 ( \26518 , \26517 , \4712 );
nand \U$26176 ( \26519 , \26512 , \26518 );
nand \U$26177 ( \26520 , \26504 , \26519 );
nand \U$26178 ( \26521 , \26503 , \26520 );
not \U$26179 ( \26522 , \26521 );
and \U$26180 ( \26523 , \26480 , \26522 );
not \U$26181 ( \26524 , \26480 );
and \U$26182 ( \26525 , \26524 , \26521 );
nor \U$26183 ( \26526 , \26523 , \26525 );
not \U$26184 ( \26527 , \26526 );
or \U$26185 ( \26528 , \26433 , \26527 );
not \U$26186 ( \26529 , \4714 );
not \U$26187 ( \26530 , \26517 );
or \U$26188 ( \26531 , \26529 , \26530 );
not \U$26189 ( \26532 , RIbb2e620_35);
not \U$26190 ( \26533 , \16865 );
or \U$26191 ( \26534 , \26532 , \26533 );
nand \U$26192 ( \26535 , \12932 , \6002 );
nand \U$26193 ( \26536 , \26534 , \26535 );
nand \U$26194 ( \26537 , \26536 , \4712 );
nand \U$26195 ( \26538 , \26531 , \26537 );
not \U$26196 ( \26539 , \26538 );
not \U$26197 ( \26540 , \2925 );
not \U$26198 ( \26541 , \26092 );
or \U$26199 ( \26542 , \26540 , \26541 );
not \U$26200 ( \26543 , RIbb2e8f0_29);
not \U$26201 ( \26544 , \15471 );
or \U$26202 ( \26545 , \26543 , \26544 );
nand \U$26203 ( \26546 , \17682 , \6970 );
nand \U$26204 ( \26547 , \26545 , \26546 );
nand \U$26205 ( \26548 , \26547 , \2921 );
nand \U$26206 ( \26549 , \26542 , \26548 );
not \U$26207 ( \26550 , \26549 );
nand \U$26208 ( \26551 , \26539 , \26550 );
not \U$26209 ( \26552 , \26551 );
not \U$26210 ( \26553 , \16427 );
not \U$26211 ( \26554 , \26450 );
or \U$26212 ( \26555 , \26553 , \26554 );
not \U$26213 ( \26556 , RIbb2df90_49);
not \U$26214 ( \26557 , \17341 );
or \U$26215 ( \26558 , \26556 , \26557 );
nand \U$26216 ( \26559 , \7111 , \12278 );
nand \U$26217 ( \26560 , \26558 , \26559 );
nand \U$26218 ( \26561 , \26560 , \12167 );
nand \U$26219 ( \26562 , \26555 , \26561 );
not \U$26220 ( \26563 , \26562 );
or \U$26221 ( \26564 , \26552 , \26563 );
nand \U$26222 ( \26565 , \26538 , \26549 );
nand \U$26223 ( \26566 , \26564 , \26565 );
or \U$26224 ( \26567 , RIbb2ec38_22, RIbb2ebc0_23);
nand \U$26225 ( \26568 , \26567 , \19064 );
and \U$26226 ( \26569 , RIbb2ec38_22, RIbb2ebc0_23);
nor \U$26227 ( \26570 , \26569 , \849 );
and \U$26228 ( \26571 , \26568 , \26570 );
not \U$26229 ( \26572 , \2078 );
not \U$26230 ( \26573 , \26061 );
or \U$26231 ( \26574 , \26572 , \26573 );
and \U$26232 ( \26575 , RIbb2ecb0_21, \17506 );
not \U$26233 ( \26576 , RIbb2ecb0_21);
and \U$26234 ( \26577 , \26576 , \18929 );
nor \U$26235 ( \26578 , \26575 , \26577 );
nand \U$26236 ( \26579 , \26578 , \2076 );
nand \U$26237 ( \26580 , \26574 , \26579 );
xor \U$26238 ( \26581 , \26571 , \26580 );
not \U$26239 ( \26582 , \3381 );
not \U$26240 ( \26583 , \26070 );
or \U$26241 ( \26584 , \26582 , \26583 );
not \U$26242 ( \26585 , RIbb2ebc0_23);
not \U$26243 ( \26586 , \26050 );
or \U$26244 ( \26587 , \26585 , \26586 );
nand \U$26245 ( \26588 , \16818 , \3401 );
nand \U$26246 ( \26589 , \26587 , \26588 );
nand \U$26247 ( \26590 , \26589 , \3406 );
nand \U$26248 ( \26591 , \26584 , \26590 );
xor \U$26249 ( \26592 , \26581 , \26591 );
not \U$26250 ( \26593 , \3445 );
not \U$26251 ( \26594 , RIbb2e9e0_27);
not \U$26252 ( \26595 , \16747 );
or \U$26253 ( \26596 , \26594 , \26595 );
nand \U$26254 ( \26597 , \16751 , \3454 );
nand \U$26255 ( \26598 , \26596 , \26597 );
not \U$26256 ( \26599 , \26598 );
or \U$26257 ( \26600 , \26593 , \26599 );
not \U$26258 ( \26601 , RIbb2e9e0_27);
not \U$26259 ( \26602 , \16844 );
or \U$26260 ( \26603 , \26601 , \26602 );
nand \U$26261 ( \26604 , \16576 , \11284 );
nand \U$26262 ( \26605 , \26603 , \26604 );
nand \U$26263 ( \26606 , \26605 , \3465 );
nand \U$26264 ( \26607 , \26600 , \26606 );
and \U$26265 ( \26608 , \26592 , \26607 );
and \U$26266 ( \26609 , \26581 , \26591 );
or \U$26267 ( \26610 , \26608 , \26609 );
not \U$26268 ( \26611 , \7103 );
and \U$26269 ( \26612 , RIbb2e440_39, \12249 );
not \U$26270 ( \26613 , RIbb2e440_39);
and \U$26271 ( \26614 , \26613 , \10764 );
or \U$26272 ( \26615 , \26612 , \26614 );
not \U$26273 ( \26616 , \26615 );
or \U$26274 ( \26617 , \26611 , \26616 );
and \U$26275 ( \26618 , RIbb2e440_39, \12234 );
not \U$26276 ( \26619 , RIbb2e440_39);
and \U$26277 ( \26620 , \26619 , \10301 );
or \U$26278 ( \26621 , \26618 , \26620 );
nand \U$26279 ( \26622 , \26621 , \8450 );
nand \U$26280 ( \26623 , \26617 , \26622 );
xor \U$26281 ( \26624 , \26610 , \26623 );
not \U$26282 ( \26625 , \12692 );
and \U$26283 ( \26626 , RIbb2dea0_51, \4325 );
not \U$26284 ( \26627 , RIbb2dea0_51);
and \U$26285 ( \26628 , \26627 , \13551 );
or \U$26286 ( \26629 , \26626 , \26628 );
not \U$26287 ( \26630 , \26629 );
or \U$26288 ( \26631 , \26625 , \26630 );
not \U$26289 ( \26632 , RIbb2dea0_51);
not \U$26290 ( \26633 , \13559 );
or \U$26291 ( \26634 , \26632 , \26633 );
or \U$26292 ( \26635 , \20387 , RIbb2dea0_51);
nand \U$26293 ( \26636 , \26634 , \26635 );
nand \U$26294 ( \26637 , \14067 , \26636 );
nand \U$26295 ( \26638 , \26631 , \26637 );
and \U$26296 ( \26639 , \26624 , \26638 );
and \U$26297 ( \26640 , \26610 , \26623 );
or \U$26298 ( \26641 , \26639 , \26640 );
xor \U$26299 ( \26642 , \26566 , \26641 );
and \U$26300 ( \26643 , \26571 , \26580 );
not \U$26301 ( \26644 , \2979 );
and \U$26302 ( \26645 , RIbb2ead0_25, \19831 );
not \U$26303 ( \26646 , RIbb2ead0_25);
and \U$26304 ( \26647 , \26646 , \23185 );
nor \U$26305 ( \26648 , \26645 , \26647 );
not \U$26306 ( \26649 , \26648 );
or \U$26307 ( \26650 , \26644 , \26649 );
nand \U$26308 ( \26651 , \26403 , \2963 );
nand \U$26309 ( \26652 , \26650 , \26651 );
xor \U$26310 ( \26653 , \26643 , \26652 );
not \U$26311 ( \26654 , \3465 );
not \U$26312 ( \26655 , \26012 );
or \U$26313 ( \26656 , \26654 , \26655 );
nand \U$26314 ( \26657 , \26605 , \3445 );
nand \U$26315 ( \26658 , \26656 , \26657 );
xor \U$26316 ( \26659 , \26653 , \26658 );
not \U$26317 ( \26660 , \16533 );
not \U$26318 ( \26661 , RIbb2d9f0_61);
not \U$26319 ( \26662 , \3516 );
or \U$26320 ( \26663 , \26661 , \26662 );
nand \U$26321 ( \26664 , \3341 , \16537 );
nand \U$26322 ( \26665 , \26663 , \26664 );
not \U$26323 ( \26666 , \26665 );
or \U$26324 ( \26667 , \26660 , \26666 );
not \U$26325 ( \26668 , RIbb2d9f0_61);
not \U$26326 ( \26669 , \6107 );
or \U$26327 ( \26670 , \26668 , \26669 );
nand \U$26328 ( \26671 , \6108 , \19746 );
nand \U$26329 ( \26672 , \26670 , \26671 );
nand \U$26330 ( \26673 , \26672 , \18717 );
nand \U$26331 ( \26674 , \26667 , \26673 );
xor \U$26332 ( \26675 , \26659 , \26674 );
not \U$26333 ( \26676 , \15182 );
and \U$26334 ( \26677 , RIbb2dcc0_55, \22894 );
not \U$26335 ( \26678 , RIbb2dcc0_55);
and \U$26336 ( \26679 , \26678 , \4022 );
or \U$26337 ( \26680 , \26677 , \26679 );
not \U$26338 ( \26681 , \26680 );
or \U$26339 ( \26682 , \26676 , \26681 );
not \U$26340 ( \26683 , RIbb2dcc0_55);
not \U$26341 ( \26684 , \13738 );
or \U$26342 ( \26685 , \26683 , \26684 );
not \U$26343 ( \26686 , RIbb2dcc0_55);
nand \U$26344 ( \26687 , \26686 , \12596 );
nand \U$26345 ( \26688 , \26685 , \26687 );
nand \U$26346 ( \26689 , \26688 , \14613 );
nand \U$26347 ( \26690 , \26682 , \26689 );
and \U$26348 ( \26691 , \26675 , \26690 );
and \U$26349 ( \26692 , \26659 , \26674 );
or \U$26350 ( \26693 , \26691 , \26692 );
and \U$26351 ( \26694 , \26642 , \26693 );
and \U$26352 ( \26695 , \26566 , \26641 );
or \U$26353 ( \26696 , \26694 , \26695 );
nand \U$26354 ( \26697 , \26528 , \26696 );
not \U$26355 ( \26698 , \26432 );
not \U$26356 ( \26699 , \26526 );
nand \U$26357 ( \26700 , \26698 , \26699 );
nand \U$26358 ( \26701 , \26697 , \26700 );
and \U$26359 ( \26702 , \26273 , \26701 );
and \U$26360 ( \26703 , \26270 , \26272 );
or \U$26361 ( \26704 , \26702 , \26703 );
xor \U$26362 ( \26705 , \26110 , \26704 );
and \U$26363 ( \26706 , \25777 , \25791 );
not \U$26364 ( \26707 , \2078 );
not \U$26365 ( \26708 , RIbb2ecb0_21);
not \U$26366 ( \26709 , \16747 );
or \U$26367 ( \26710 , \26708 , \26709 );
nand \U$26368 ( \26711 , \16856 , \2067 );
nand \U$26369 ( \26712 , \26710 , \26711 );
not \U$26370 ( \26713 , \26712 );
or \U$26371 ( \26714 , \26707 , \26713 );
not \U$26372 ( \26715 , RIbb2ecb0_21);
not \U$26373 ( \26716 , \23185 );
or \U$26374 ( \26717 , \26715 , \26716 );
nand \U$26375 ( \26718 , \16829 , \2254 );
nand \U$26376 ( \26719 , \26717 , \26718 );
nand \U$26377 ( \26720 , \26719 , \2077 );
nand \U$26378 ( \26721 , \26714 , \26720 );
xor \U$26379 ( \26722 , \26706 , \26721 );
not \U$26380 ( \26723 , \3382 );
not \U$26381 ( \26724 , RIbb2ebc0_23);
not \U$26382 ( \26725 , \16561 );
or \U$26383 ( \26726 , \26724 , \26725 );
nand \U$26384 ( \26727 , \23098 , \3396 );
nand \U$26385 ( \26728 , \26726 , \26727 );
not \U$26386 ( \26729 , \26728 );
or \U$26387 ( \26730 , \26723 , \26729 );
nand \U$26388 ( \26731 , \25814 , \3406 );
nand \U$26389 ( \26732 , \26730 , \26731 );
xor \U$26390 ( \26733 , \26722 , \26732 );
not \U$26391 ( \26734 , RIbb2d888_64);
not \U$26392 ( \26735 , RIbb2d900_63);
not \U$26393 ( \26736 , \1385 );
or \U$26394 ( \26737 , \26735 , \26736 );
nand \U$26395 ( \26738 , \1384 , \20254 );
nand \U$26396 ( \26739 , \26737 , \26738 );
not \U$26397 ( \26740 , \26739 );
or \U$26398 ( \26741 , \26734 , \26740 );
nand \U$26399 ( \26742 , \25627 , \17275 );
nand \U$26400 ( \26743 , \26741 , \26742 );
xor \U$26401 ( \26744 , \26733 , \26743 );
not \U$26402 ( \26745 , \14930 );
not \U$26403 ( \26746 , RIbb2ddb0_53);
not \U$26404 ( \26747 , \6172 );
or \U$26405 ( \26748 , \26746 , \26747 );
not \U$26406 ( \26749 , \6172 );
not \U$26407 ( \26750 , RIbb2ddb0_53);
nand \U$26408 ( \26751 , \26749 , \26750 );
nand \U$26409 ( \26752 , \26748 , \26751 );
not \U$26410 ( \26753 , \26752 );
or \U$26411 ( \26754 , \26745 , \26753 );
nand \U$26412 ( \26755 , \25705 , \17562 );
nand \U$26413 ( \26756 , \26754 , \26755 );
xor \U$26414 ( \26757 , \26744 , \26756 );
not \U$26415 ( \26758 , \2078 );
not \U$26416 ( \26759 , \26719 );
or \U$26417 ( \26760 , \26758 , \26759 );
not \U$26418 ( \26761 , RIbb2ecb0_21);
not \U$26419 ( \26762 , \16710 );
or \U$26420 ( \26763 , \26761 , \26762 );
nand \U$26421 ( \26764 , \16706 , \849 );
nand \U$26422 ( \26765 , \26763 , \26764 );
nand \U$26423 ( \26766 , \26765 , \2077 );
nand \U$26424 ( \26767 , \26760 , \26766 );
and \U$26425 ( \26768 , \17506 , \835 );
not \U$26426 ( \26769 , \854 );
not \U$26427 ( \26770 , \25805 );
or \U$26428 ( \26771 , \26769 , \26770 );
nand \U$26429 ( \26772 , \853 , \26131 );
nand \U$26430 ( \26773 , \26771 , \26772 );
xor \U$26431 ( \26774 , \26768 , \26773 );
not \U$26432 ( \26775 , \2078 );
not \U$26433 ( \26776 , \26765 );
or \U$26434 ( \26777 , \26775 , \26776 );
nand \U$26435 ( \26778 , \26391 , \2077 );
nand \U$26436 ( \26779 , \26777 , \26778 );
and \U$26437 ( \26780 , \26774 , \26779 );
and \U$26438 ( \26781 , \26768 , \26773 );
or \U$26439 ( \26782 , \26780 , \26781 );
xor \U$26440 ( \26783 , \26767 , \26782 );
not \U$26441 ( \26784 , \3465 );
not \U$26442 ( \26785 , RIbb2e9e0_27);
not \U$26443 ( \26786 , \16317 );
or \U$26444 ( \26787 , \26785 , \26786 );
nand \U$26445 ( \26788 , \14506 , \3454 );
nand \U$26446 ( \26789 , \26787 , \26788 );
not \U$26447 ( \26790 , \26789 );
or \U$26448 ( \26791 , \26784 , \26790 );
not \U$26449 ( \26792 , RIbb2e9e0_27);
not \U$26450 ( \26793 , \16309 );
or \U$26451 ( \26794 , \26792 , \26793 );
nand \U$26452 ( \26795 , \14527 , \6065 );
nand \U$26453 ( \26796 , \26794 , \26795 );
nand \U$26454 ( \26797 , \26796 , \3445 );
nand \U$26455 ( \26798 , \26791 , \26797 );
and \U$26456 ( \26799 , \26783 , \26798 );
and \U$26457 ( \26800 , \26767 , \26782 );
or \U$26458 ( \26801 , \26799 , \26800 );
not \U$26459 ( \26802 , \16271 );
not \U$26460 ( \26803 , \25668 );
or \U$26461 ( \26804 , \26802 , \26803 );
not \U$26462 ( \26805 , RIbb2dae0_59);
not \U$26463 ( \26806 , \2115 );
or \U$26464 ( \26807 , \26805 , \26806 );
nand \U$26465 ( \26808 , \16235 , \17024 );
nand \U$26466 ( \26809 , \26807 , \26808 );
nand \U$26467 ( \26810 , \26809 , \16257 );
nand \U$26468 ( \26811 , \26804 , \26810 );
xor \U$26469 ( \26812 , \26801 , \26811 );
not \U$26470 ( \26813 , \12692 );
and \U$26471 ( \26814 , RIbb2dea0_51, \4021 );
not \U$26472 ( \26815 , RIbb2dea0_51);
and \U$26473 ( \26816 , \26815 , \4016 );
or \U$26474 ( \26817 , \26814 , \26816 );
not \U$26475 ( \26818 , \26817 );
or \U$26476 ( \26819 , \26813 , \26818 );
not \U$26477 ( \26820 , \25685 );
nand \U$26478 ( \26821 , \26820 , \12774 );
nand \U$26479 ( \26822 , \26819 , \26821 );
xor \U$26480 ( \26823 , \26812 , \26822 );
xor \U$26481 ( \26824 , \26757 , \26823 );
not \U$26482 ( \26825 , \16541 );
not \U$26483 ( \26826 , \25757 );
or \U$26484 ( \26827 , \26825 , \26826 );
not \U$26485 ( \26828 , RIbb2d9f0_61);
not \U$26486 ( \26829 , \17207 );
or \U$26487 ( \26830 , \26828 , \26829 );
not \U$26488 ( \26831 , \17207 );
nand \U$26489 ( \26832 , \26831 , \19746 );
nand \U$26490 ( \26833 , \26830 , \26832 );
buf \U$26491 ( \26834 , \16533 );
nand \U$26492 ( \26835 , \26833 , \26834 );
nand \U$26493 ( \26836 , \26827 , \26835 );
not \U$26494 ( \26837 , \15738 );
not \U$26495 ( \26838 , RIbb2dbd0_57);
not \U$26496 ( \26839 , \12097 );
or \U$26497 ( \26840 , \26838 , \26839 );
nand \U$26498 ( \26841 , \3521 , \14602 );
nand \U$26499 ( \26842 , \26840 , \26841 );
not \U$26500 ( \26843 , \26842 );
or \U$26501 ( \26844 , \26837 , \26843 );
nand \U$26502 ( \26845 , \25635 , \15746 );
nand \U$26503 ( \26846 , \26844 , \26845 );
xor \U$26504 ( \26847 , \26836 , \26846 );
not \U$26505 ( \26848 , \15181 );
and \U$26506 ( \26849 , RIbb2dcc0_55, \3141 );
not \U$26507 ( \26850 , RIbb2dcc0_55);
not \U$26508 ( \26851 , \22978 );
and \U$26509 ( \26852 , \26850 , \26851 );
or \U$26510 ( \26853 , \26849 , \26852 );
not \U$26511 ( \26854 , \26853 );
or \U$26512 ( \26855 , \26848 , \26854 );
nand \U$26513 ( \26856 , \25652 , \14613 );
nand \U$26514 ( \26857 , \26855 , \26856 );
xor \U$26515 ( \26858 , \26847 , \26857 );
xor \U$26516 ( \26859 , \26824 , \26858 );
xor \U$26517 ( \26860 , \25660 , \25629 );
xnor \U$26518 ( \26861 , \26860 , \25644 );
not \U$26519 ( \26862 , \26861 );
not \U$26520 ( \26863 , \26862 );
xor \U$26521 ( \26864 , \26768 , \26773 );
xor \U$26522 ( \26865 , \26864 , \26779 );
not \U$26523 ( \26866 , \2922 );
not \U$26524 ( \26867 , \26085 );
or \U$26525 ( \26868 , \26866 , \26867 );
not \U$26526 ( \26869 , RIbb2e8f0_29);
not \U$26527 ( \26870 , \13546 );
or \U$26528 ( \26871 , \26869 , \26870 );
not \U$26529 ( \26872 , \13986 );
nand \U$26530 ( \26873 , \26872 , \3440 );
nand \U$26531 ( \26874 , \26871 , \26873 );
nand \U$26532 ( \26875 , \26874 , \2925 );
nand \U$26533 ( \26876 , \26868 , \26875 );
xor \U$26534 ( \26877 , \26865 , \26876 );
not \U$26535 ( \26878 , \3445 );
not \U$26536 ( \26879 , \26004 );
or \U$26537 ( \26880 , \26878 , \26879 );
nand \U$26538 ( \26881 , \26796 , \3465 );
nand \U$26539 ( \26882 , \26880 , \26881 );
xor \U$26540 ( \26883 , \26877 , \26882 );
not \U$26541 ( \26884 , \3613 );
not \U$26542 ( \26885 , RIbb2e800_31);
not \U$26543 ( \26886 , \12348 );
or \U$26544 ( \26887 , \26885 , \26886 );
nand \U$26545 ( \26888 , \16765 , \3608 );
nand \U$26546 ( \26889 , \26887 , \26888 );
not \U$26547 ( \26890 , \26889 );
or \U$26548 ( \26891 , \26884 , \26890 );
nand \U$26549 ( \26892 , \25976 , \2940 );
nand \U$26550 ( \26893 , \26891 , \26892 );
not \U$26551 ( \26894 , \4075 );
not \U$26552 ( \26895 , RIbb2e710_33);
not \U$26553 ( \26896 , \22070 );
or \U$26554 ( \26897 , \26895 , \26896 );
nand \U$26555 ( \26898 , \12175 , \2935 );
nand \U$26556 ( \26899 , \26897 , \26898 );
not \U$26557 ( \26900 , \26899 );
or \U$26558 ( \26901 , \26894 , \26900 );
nand \U$26559 ( \26902 , \25993 , \3887 );
nand \U$26560 ( \26903 , \26901 , \26902 );
xor \U$26561 ( \26904 , \26893 , \26903 );
not \U$26562 ( \26905 , \11177 );
not \U$26563 ( \26906 , RIbb2e080_47);
not \U$26564 ( \26907 , \10556 );
or \U$26565 ( \26908 , \26906 , \26907 );
not \U$26566 ( \26909 , \18624 );
nand \U$26567 ( \26910 , \26909 , \12971 );
nand \U$26568 ( \26911 , \26908 , \26910 );
not \U$26569 ( \26912 , \26911 );
or \U$26570 ( \26913 , \26905 , \26912 );
nand \U$26571 ( \26914 , \26441 , \11176 );
nand \U$26572 ( \26915 , \26913 , \26914 );
xor \U$26573 ( \26916 , \26904 , \26915 );
xor \U$26574 ( \26917 , \26883 , \26916 );
xor \U$26575 ( \26918 , \26643 , \26652 );
and \U$26576 ( \26919 , \26918 , \26658 );
and \U$26577 ( \26920 , \26643 , \26652 );
or \U$26578 ( \26921 , \26919 , \26920 );
not \U$26579 ( \26922 , \7104 );
and \U$26580 ( \26923 , RIbb2e440_39, \14550 );
not \U$26581 ( \26924 , RIbb2e440_39);
and \U$26582 ( \26925 , \26924 , \20045 );
or \U$26583 ( \26926 , \26923 , \26925 );
not \U$26584 ( \26927 , \26926 );
or \U$26585 ( \26928 , \26922 , \26927 );
buf \U$26586 ( \26929 , \26621 );
nand \U$26587 ( \26930 , \26929 , \8445 );
nand \U$26588 ( \26931 , \26928 , \26930 );
xor \U$26589 ( \26932 , \26921 , \26931 );
not \U$26590 ( \26933 , \6242 );
not \U$26591 ( \26934 , RIbb2e530_37);
not \U$26592 ( \26935 , \12249 );
or \U$26593 ( \26936 , \26934 , \26935 );
not \U$26594 ( \26937 , \12249 );
nand \U$26595 ( \26938 , \26937 , \6246 );
nand \U$26596 ( \26939 , \26936 , \26938 );
not \U$26597 ( \26940 , \26939 );
or \U$26598 ( \26941 , \26933 , \26940 );
nand \U$26599 ( \26942 , \26327 , \6251 );
nand \U$26600 ( \26943 , \26941 , \26942 );
and \U$26601 ( \26944 , \26932 , \26943 );
and \U$26602 ( \26945 , \26921 , \26931 );
or \U$26603 ( \26946 , \26944 , \26945 );
and \U$26604 ( \26947 , \26917 , \26946 );
and \U$26605 ( \26948 , \26883 , \26916 );
or \U$26606 ( \26949 , \26947 , \26948 );
not \U$26607 ( \26950 , \26949 );
or \U$26608 ( \26951 , \26863 , \26950 );
or \U$26609 ( \26952 , \26949 , \26862 );
xor \U$26610 ( \26953 , \26767 , \26782 );
xor \U$26611 ( \26954 , \26953 , \26798 );
xor \U$26612 ( \26955 , \26865 , \26876 );
and \U$26613 ( \26956 , \26955 , \26882 );
and \U$26614 ( \26957 , \26865 , \26876 );
or \U$26615 ( \26958 , \26956 , \26957 );
xor \U$26616 ( \26959 , \26954 , \26958 );
not \U$26617 ( \26960 , \2925 );
not \U$26618 ( \26961 , RIbb2e8f0_29);
not \U$26619 ( \26962 , \18857 );
or \U$26620 ( \26963 , \26961 , \26962 );
buf \U$26621 ( \26964 , \13210 );
nand \U$26622 ( \26965 , \26964 , \3800 );
nand \U$26623 ( \26966 , \26963 , \26965 );
not \U$26624 ( \26967 , \26966 );
or \U$26625 ( \26968 , \26960 , \26967 );
nand \U$26626 ( \26969 , \2921 , \26874 );
nand \U$26627 ( \26970 , \26968 , \26969 );
not \U$26628 ( \26971 , \2963 );
and \U$26629 ( \26972 , RIbb2ead0_25, \16783 );
not \U$26630 ( \26973 , RIbb2ead0_25);
and \U$26631 ( \26974 , \26973 , \15474 );
or \U$26632 ( \26975 , \26972 , \26974 );
not \U$26633 ( \26976 , \26975 );
or \U$26634 ( \26977 , \26971 , \26976 );
nand \U$26635 ( \26978 , \26153 , \2980 );
nand \U$26636 ( \26979 , \26977 , \26978 );
xor \U$26637 ( \26980 , \26970 , \26979 );
not \U$26638 ( \26981 , \3613 );
not \U$26639 ( \26982 , RIbb2e800_31);
not \U$26640 ( \26983 , \14636 );
or \U$26641 ( \26984 , \26982 , \26983 );
not \U$26642 ( \26985 , \18842 );
nand \U$26643 ( \26986 , \26985 , \9169 );
nand \U$26644 ( \26987 , \26984 , \26986 );
not \U$26645 ( \26988 , \26987 );
or \U$26646 ( \26989 , \26981 , \26988 );
nand \U$26647 ( \26990 , \26889 , \2940 );
nand \U$26648 ( \26991 , \26989 , \26990 );
xor \U$26649 ( \26992 , \26980 , \26991 );
xor \U$26650 ( \26993 , \26959 , \26992 );
nand \U$26651 ( \26994 , \26952 , \26993 );
nand \U$26652 ( \26995 , \26951 , \26994 );
xor \U$26653 ( \26996 , \26859 , \26995 );
xor \U$26654 ( \26997 , \26893 , \26903 );
and \U$26655 ( \26998 , \26997 , \26915 );
and \U$26656 ( \26999 , \26893 , \26903 );
or \U$26657 ( \27000 , \26998 , \26999 );
xor \U$26658 ( \27001 , \26385 , \26395 );
and \U$26659 ( \27002 , \27001 , \26405 );
and \U$26660 ( \27003 , \26385 , \26395 );
or \U$26661 ( \27004 , \27002 , \27003 );
not \U$26662 ( \27005 , \7103 );
not \U$26663 ( \27006 , \26926 );
or \U$26664 ( \27007 , \27005 , \27006 );
and \U$26665 ( \27008 , RIbb2e440_39, \13916 );
not \U$26666 ( \27009 , RIbb2e440_39);
and \U$26667 ( \27010 , \27009 , \9278 );
or \U$26668 ( \27011 , \27008 , \27010 );
nand \U$26669 ( \27012 , \27011 , \7104 );
nand \U$26670 ( \27013 , \27007 , \27012 );
xor \U$26671 ( \27014 , \27004 , \27013 );
not \U$26672 ( \27015 , \8353 );
not \U$26673 ( \27016 , RIbb2e350_41);
not \U$26674 ( \27017 , \12211 );
or \U$26675 ( \27018 , \27016 , \27017 );
nand \U$26676 ( \27019 , \12214 , \9402 );
nand \U$26677 ( \27020 , \27018 , \27019 );
not \U$26678 ( \27021 , \27020 );
or \U$26679 ( \27022 , \27015 , \27021 );
nand \U$26680 ( \27023 , \26414 , \8361 );
nand \U$26681 ( \27024 , \27022 , \27023 );
and \U$26682 ( \27025 , \27014 , \27024 );
and \U$26683 ( \27026 , \27004 , \27013 );
or \U$26684 ( \27027 , \27025 , \27026 );
xor \U$26685 ( \27028 , \27000 , \27027 );
not \U$26686 ( \27029 , \9098 );
not \U$26687 ( \27030 , \26424 );
or \U$26688 ( \27031 , \27029 , \27030 );
not \U$26689 ( \27032 , RIbb2e260_43);
not \U$26690 ( \27033 , \15066 );
or \U$26691 ( \27034 , \27032 , \27033 );
nand \U$26692 ( \27035 , \25844 , \8347 );
nand \U$26693 ( \27036 , \27034 , \27035 );
nand \U$26694 ( \27037 , \27036 , \10451 );
nand \U$26695 ( \27038 , \27031 , \27037 );
not \U$26696 ( \27039 , \12167 );
not \U$26697 ( \27040 , \26457 );
or \U$26698 ( \27041 , \27039 , \27040 );
nand \U$26699 ( \27042 , \25748 , \12284 );
nand \U$26700 ( \27043 , \27041 , \27042 );
xor \U$26701 ( \27044 , \27038 , \27043 );
not \U$26702 ( \27045 , \10119 );
not \U$26703 ( \27046 , RIbb2e170_45);
not \U$26704 ( \27047 , \18564 );
or \U$26705 ( \27048 , \27046 , \27047 );
nand \U$26706 ( \27049 , \7308 , \13372 );
nand \U$26707 ( \27050 , \27048 , \27049 );
not \U$26708 ( \27051 , \27050 );
or \U$26709 ( \27052 , \27045 , \27051 );
nand \U$26710 ( \27053 , \26469 , \10599 );
nand \U$26711 ( \27054 , \27052 , \27053 );
and \U$26712 ( \27055 , \27044 , \27054 );
and \U$26713 ( \27056 , \27038 , \27043 );
or \U$26714 ( \27057 , \27055 , \27056 );
xor \U$26715 ( \27058 , \27028 , \27057 );
not \U$26716 ( \27059 , \26475 );
not \U$26717 ( \27060 , \26521 );
or \U$26718 ( \27061 , \27059 , \27060 );
not \U$26719 ( \27062 , \26475 );
not \U$26720 ( \27063 , \27062 );
not \U$26721 ( \27064 , \26522 );
or \U$26722 ( \27065 , \27063 , \27064 );
nand \U$26723 ( \27066 , \27065 , \26479 );
nand \U$26724 ( \27067 , \27061 , \27066 );
xor \U$26725 ( \27068 , \27058 , \27067 );
xor \U$26726 ( \27069 , \27004 , \27013 );
xor \U$26727 ( \27070 , \27069 , \27024 );
xor \U$26728 ( \27071 , \27038 , \27043 );
xor \U$26729 ( \27072 , \27071 , \27054 );
xor \U$26730 ( \27073 , \27070 , \27072 );
not \U$26731 ( \27074 , \15688 );
not \U$26732 ( \27075 , \26169 );
or \U$26733 ( \27076 , \27074 , \27075 );
nand \U$26734 ( \27077 , \26370 , \17562 );
nand \U$26735 ( \27078 , \27076 , \27077 );
not \U$26736 ( \27079 , \22952 );
not \U$26737 ( \27080 , \26680 );
or \U$26738 ( \27081 , \27079 , \27080 );
not \U$26739 ( \27082 , RIbb2dcc0_55);
not \U$26740 ( \27083 , \7018 );
or \U$26741 ( \27084 , \27082 , \27083 );
or \U$26742 ( \27085 , \21490 , RIbb2dcc0_55);
nand \U$26743 ( \27086 , \27084 , \27085 );
nand \U$26744 ( \27087 , \27086 , \15181 );
nand \U$26745 ( \27088 , \27081 , \27087 );
or \U$26746 ( \27089 , \27078 , \27088 );
not \U$26747 ( \27090 , \16533 );
not \U$26748 ( \27091 , RIbb2d9f0_61);
not \U$26749 ( \27092 , \13289 );
or \U$26750 ( \27093 , \27091 , \27092 );
not \U$26751 ( \27094 , \13286 );
nand \U$26752 ( \27095 , \27094 , \16537 );
nand \U$26753 ( \27096 , \27093 , \27095 );
not \U$26754 ( \27097 , \27096 );
or \U$26755 ( \27098 , \27090 , \27097 );
nand \U$26756 ( \27099 , \26665 , \16541 );
nand \U$26757 ( \27100 , \27098 , \27099 );
nand \U$26758 ( \27101 , \27089 , \27100 );
nand \U$26759 ( \27102 , \27078 , \27088 );
nand \U$26760 ( \27103 , \27101 , \27102 );
and \U$26761 ( \27104 , \27073 , \27103 );
and \U$26762 ( \27105 , \27070 , \27072 );
or \U$26763 ( \27106 , \27104 , \27105 );
and \U$26764 ( \27107 , \27068 , \27106 );
and \U$26765 ( \27108 , \27058 , \27067 );
or \U$26766 ( \27109 , \27107 , \27108 );
xor \U$26767 ( \27110 , \26996 , \27109 );
xor \U$26768 ( \27111 , \26705 , \27110 );
xor \U$26769 ( \27112 , \26883 , \26916 );
xor \U$26770 ( \27113 , \27112 , \26946 );
xor \U$26771 ( \27114 , \27070 , \27072 );
xor \U$26772 ( \27115 , \27114 , \27103 );
xor \U$26773 ( \27116 , \27113 , \27115 );
xor \U$26774 ( \27117 , \26921 , \26931 );
xor \U$26775 ( \27118 , \27117 , \26943 );
xor \U$26776 ( \27119 , \26459 , \26473 );
xor \U$26777 ( \27120 , \27119 , \26443 );
xor \U$26778 ( \27121 , \27118 , \27120 );
xor \U$26779 ( \27122 , \26519 , \26490 );
xor \U$26780 ( \27123 , \27122 , \26501 );
and \U$26781 ( \27124 , \27121 , \27123 );
and \U$26782 ( \27125 , \27118 , \27120 );
or \U$26783 ( \27126 , \27124 , \27125 );
xnor \U$26784 ( \27127 , \27116 , \27126 );
buf \U$26785 ( \27128 , \27127 );
not \U$26786 ( \27129 , \27128 );
xor \U$26787 ( \27130 , \26046 , \26078 );
xor \U$26788 ( \27131 , \27130 , \26094 );
not \U$26789 ( \27132 , \16257 );
not \U$26790 ( \27133 , \26115 );
or \U$26791 ( \27134 , \27132 , \27133 );
nand \U$26792 ( \27135 , \26343 , \16271 );
nand \U$26793 ( \27136 , \27134 , \27135 );
xor \U$26794 ( \27137 , \27131 , \27136 );
not \U$26795 ( \27138 , \12692 );
not \U$26796 ( \27139 , \26025 );
or \U$26797 ( \27140 , \27138 , \27139 );
nand \U$26798 ( \27141 , \26629 , \14067 );
nand \U$26799 ( \27142 , \27140 , \27141 );
xor \U$26800 ( \27143 , \27137 , \27142 );
xor \U$26801 ( \27144 , \27100 , \27078 );
xor \U$26802 ( \27145 , \27144 , \27088 );
xor \U$26803 ( \27146 , \27143 , \27145 );
xor \U$26804 ( \27147 , \26581 , \26591 );
xor \U$26805 ( \27148 , \27147 , \26607 );
not \U$26806 ( \27149 , \12692 );
not \U$26807 ( \27150 , \26636 );
or \U$26808 ( \27151 , \27149 , \27150 );
and \U$26809 ( \27152 , RIbb2dea0_51, \18624 );
not \U$26810 ( \27153 , RIbb2dea0_51);
and \U$26811 ( \27154 , \27153 , \18623 );
or \U$26812 ( \27155 , \27152 , \27154 );
nand \U$26813 ( \27156 , \27155 , \12774 );
nand \U$26814 ( \27157 , \27151 , \27156 );
xor \U$26815 ( \27158 , \27148 , \27157 );
not \U$26816 ( \27159 , \26257 );
not \U$26817 ( \27160 , \9099 );
or \U$26818 ( \27161 , \27159 , \27160 );
not \U$26819 ( \27162 , RIbb2e260_43);
not \U$26820 ( \27163 , \13919 );
or \U$26821 ( \27164 , \27162 , \27163 );
not \U$26822 ( \27165 , \18578 );
nand \U$26823 ( \27166 , \27165 , \9847 );
nand \U$26824 ( \27167 , \27164 , \27166 );
nand \U$26825 ( \27168 , \27167 , \10449 );
nand \U$26826 ( \27169 , \27161 , \27168 );
and \U$26827 ( \27170 , \27158 , \27169 );
and \U$26828 ( \27171 , \27148 , \27157 );
or \U$26829 ( \27172 , \27170 , \27171 );
not \U$26830 ( \27173 , \2941 );
not \U$26831 ( \27174 , \26189 );
or \U$26832 ( \27175 , \27173 , \27174 );
not \U$26833 ( \27176 , RIbb2e800_31);
not \U$26834 ( \27177 , \16309 );
or \U$26835 ( \27178 , \27176 , \27177 );
nand \U$26836 ( \27179 , \14526 , \9169 );
nand \U$26837 ( \27180 , \27178 , \27179 );
nand \U$26838 ( \27181 , \27180 , \2939 );
nand \U$26839 ( \27182 , \27175 , \27181 );
not \U$26840 ( \27183 , \2925 );
not \U$26841 ( \27184 , \26547 );
or \U$26842 ( \27185 , \27183 , \27184 );
not \U$26843 ( \27186 , RIbb2e8f0_29);
not \U$26844 ( \27187 , \16563 );
or \U$26845 ( \27188 , \27186 , \27187 );
nand \U$26846 ( \27189 , \23098 , \3800 );
nand \U$26847 ( \27190 , \27188 , \27189 );
nand \U$26848 ( \27191 , \27190 , \2922 );
nand \U$26849 ( \27192 , \27185 , \27191 );
xor \U$26850 ( \27193 , \27182 , \27192 );
not \U$26851 ( \27194 , \4714 );
not \U$26852 ( \27195 , \26536 );
or \U$26853 ( \27196 , \27194 , \27195 );
and \U$26854 ( \27197 , RIbb2e620_35, \14838 );
not \U$26855 ( \27198 , RIbb2e620_35);
not \U$26856 ( \27199 , \13809 );
and \U$26857 ( \27200 , \27198 , \27199 );
or \U$26858 ( \27201 , \27197 , \27200 );
nand \U$26859 ( \27202 , \27201 , \4712 );
nand \U$26860 ( \27203 , \27196 , \27202 );
and \U$26861 ( \27204 , \27193 , \27203 );
and \U$26862 ( \27205 , \27182 , \27192 );
or \U$26863 ( \27206 , \27204 , \27205 );
buf \U$26864 ( \27207 , \27206 );
or \U$26865 ( \27208 , \27172 , \27207 );
not \U$26866 ( \27209 , \2963 );
not \U$26867 ( \27210 , \26648 );
or \U$26868 ( \27211 , \27209 , \27210 );
and \U$26869 ( \27212 , RIbb2ead0_25, \16710 );
not \U$26870 ( \27213 , RIbb2ead0_25);
and \U$26871 ( \27214 , \27213 , \16706 );
or \U$26872 ( \27215 , \27212 , \27214 );
nand \U$26873 ( \27216 , \27215 , \2980 );
nand \U$26874 ( \27217 , \27211 , \27216 );
and \U$26875 ( \27218 , \17506 , \2078 );
not \U$26876 ( \27219 , \3381 );
not \U$26877 ( \27220 , \26589 );
or \U$26878 ( \27221 , \27219 , \27220 );
not \U$26879 ( \27222 , RIbb2ebc0_23);
not \U$26880 ( \27223 , \20552 );
or \U$26881 ( \27224 , \27222 , \27223 );
not \U$26882 ( \27225 , \17744 );
nand \U$26883 ( \27226 , \27225 , \3401 );
nand \U$26884 ( \27227 , \27224 , \27226 );
nand \U$26885 ( \27228 , \27227 , \3405 );
nand \U$26886 ( \27229 , \27221 , \27228 );
xor \U$26887 ( \27230 , \27218 , \27229 );
not \U$26888 ( \27231 , \2962 );
not \U$26889 ( \27232 , \27215 );
or \U$26890 ( \27233 , \27231 , \27232 );
not \U$26891 ( \27234 , \16704 );
and \U$26892 ( \27235 , RIbb2ead0_25, \27234 );
not \U$26893 ( \27236 , RIbb2ead0_25);
not \U$26894 ( \27237 , \17755 );
and \U$26895 ( \27238 , \27236 , \27237 );
or \U$26896 ( \27239 , \27235 , \27238 );
nand \U$26897 ( \27240 , \27239 , \2979 );
nand \U$26898 ( \27241 , \27233 , \27240 );
and \U$26899 ( \27242 , \27230 , \27241 );
and \U$26900 ( \27243 , \27218 , \27229 );
or \U$26901 ( \27244 , \27242 , \27243 );
xor \U$26902 ( \27245 , \27217 , \27244 );
not \U$26903 ( \27246 , \4791 );
not \U$26904 ( \27247 , \26200 );
or \U$26905 ( \27248 , \27246 , \27247 );
not \U$26906 ( \27249 , RIbb2e710_33);
not \U$26907 ( \27250 , \15054 );
or \U$26908 ( \27251 , \27249 , \27250 );
nand \U$26909 ( \27252 , \26872 , \7390 );
nand \U$26910 ( \27253 , \27251 , \27252 );
nand \U$26911 ( \27254 , \27253 , \3886 );
nand \U$26912 ( \27255 , \27248 , \27254 );
and \U$26913 ( \27256 , \27245 , \27255 );
and \U$26914 ( \27257 , \27217 , \27244 );
or \U$26915 ( \27258 , \27256 , \27257 );
nand \U$26916 ( \27259 , \27208 , \27258 );
nand \U$26917 ( \27260 , \27172 , \27207 );
nand \U$26918 ( \27261 , \27259 , \27260 );
and \U$26919 ( \27262 , \27146 , \27261 );
and \U$26920 ( \27263 , \27143 , \27145 );
or \U$26921 ( \27264 , \27262 , \27263 );
not \U$26922 ( \27265 , \27264 );
not \U$26923 ( \27266 , \27265 );
not \U$26924 ( \27267 , \4712 );
not \U$26925 ( \27268 , \26510 );
or \U$26926 ( \27269 , \27267 , \27268 );
nand \U$26927 ( \27270 , \25732 , \5845 );
nand \U$26928 ( \27271 , \27269 , \27270 );
not \U$26929 ( \27272 , \16675 );
not \U$26930 ( \27273 , \26486 );
or \U$26931 ( \27274 , \27272 , \27273 );
nand \U$26932 ( \27275 , \25642 , \17397 );
nand \U$26933 ( \27276 , \27274 , \27275 );
xor \U$26934 ( \27277 , \27271 , \27276 );
not \U$26935 ( \27278 , \6242 );
not \U$26936 ( \27279 , RIbb2e530_37);
not \U$26937 ( \27280 , \12744 );
or \U$26938 ( \27281 , \27279 , \27280 );
nand \U$26939 ( \27282 , \10301 , \8701 );
nand \U$26940 ( \27283 , \27281 , \27282 );
not \U$26941 ( \27284 , \27283 );
or \U$26942 ( \27285 , \27278 , \27284 );
nand \U$26943 ( \27286 , \26939 , \6251 );
nand \U$26944 ( \27287 , \27285 , \27286 );
xor \U$26945 ( \27288 , \27277 , \27287 );
xor \U$26946 ( \27289 , \27131 , \27136 );
and \U$26947 ( \27290 , \27289 , \27142 );
and \U$26948 ( \27291 , \27131 , \27136 );
or \U$26949 ( \27292 , \27290 , \27291 );
xor \U$26950 ( \27293 , \27288 , \27292 );
not \U$26951 ( \27294 , \15182 );
not \U$26952 ( \27295 , \25658 );
or \U$26953 ( \27296 , \27294 , \27295 );
nand \U$26954 ( \27297 , \27086 , \22952 );
nand \U$26955 ( \27298 , \27296 , \27297 );
not \U$26956 ( \27299 , \17275 );
not \U$26957 ( \27300 , \26497 );
or \U$26958 ( \27301 , \27299 , \27300 );
nand \U$26959 ( \27302 , \25621 , RIbb2d888_64);
nand \U$26960 ( \27303 , \27301 , \27302 );
xor \U$26961 ( \27304 , \27298 , \27303 );
not \U$26962 ( \27305 , \16541 );
not \U$26963 ( \27306 , \27096 );
or \U$26964 ( \27307 , \27305 , \27306 );
nand \U$26965 ( \27308 , \25764 , \26834 );
nand \U$26966 ( \27309 , \27307 , \27308 );
xor \U$26967 ( \27310 , \27304 , \27309 );
xnor \U$26968 ( \27311 , \27293 , \27310 );
not \U$26969 ( \27312 , \27311 );
not \U$26970 ( \27313 , \27312 );
or \U$26971 ( \27314 , \27266 , \27313 );
nand \U$26972 ( \27315 , \27311 , \27264 );
nand \U$26973 ( \27316 , \27314 , \27315 );
not \U$26974 ( \27317 , \26174 );
not \U$26975 ( \27318 , \26267 );
or \U$26976 ( \27319 , \27317 , \27318 );
nand \U$26977 ( \27320 , \26268 , \26177 );
nand \U$26978 ( \27321 , \27319 , \27320 );
xor \U$26979 ( \27322 , \27321 , \26265 );
not \U$26980 ( \27323 , \27322 );
and \U$26981 ( \27324 , \27316 , \27323 );
not \U$26982 ( \27325 , \27316 );
and \U$26983 ( \27326 , \27325 , \27322 );
nor \U$26984 ( \27327 , \27324 , \27326 );
not \U$26985 ( \27328 , \27327 );
or \U$26986 ( \27329 , \27129 , \27328 );
xor \U$26987 ( \27330 , \26331 , \26381 );
xor \U$26988 ( \27331 , \27330 , \26429 );
xor \U$26989 ( \27332 , \27118 , \27120 );
xor \U$26990 ( \27333 , \27332 , \27123 );
xor \U$26991 ( \27334 , \27331 , \27333 );
xor \U$26992 ( \27335 , \27143 , \27145 );
xor \U$26993 ( \27336 , \27335 , \27261 );
and \U$26994 ( \27337 , \27334 , \27336 );
and \U$26995 ( \27338 , \27331 , \27333 );
or \U$26996 ( \27339 , \27337 , \27338 );
nand \U$26997 ( \27340 , \27329 , \27339 );
or \U$26998 ( \27341 , \27327 , \27128 );
nand \U$26999 ( \27342 , \27340 , \27341 );
not \U$27000 ( \27343 , \27342 );
xor \U$27001 ( \27344 , \26861 , \26993 );
xor \U$27002 ( \27345 , \27344 , \26949 );
not \U$27003 ( \27346 , \27113 );
not \U$27004 ( \27347 , \27115 );
or \U$27005 ( \27348 , \27346 , \27347 );
or \U$27006 ( \27349 , \27115 , \27113 );
nand \U$27007 ( \27350 , \27349 , \27126 );
nand \U$27008 ( \27351 , \27348 , \27350 );
xor \U$27009 ( \27352 , \27345 , \27351 );
xor \U$27010 ( \27353 , \27058 , \27067 );
xor \U$27011 ( \27354 , \27353 , \27106 );
xnor \U$27012 ( \27355 , \27352 , \27354 );
not \U$27013 ( \27356 , \27355 );
xor \U$27014 ( \27357 , \26205 , \26211 );
xor \U$27015 ( \27358 , \27357 , \26262 );
not \U$27016 ( \27359 , \26259 );
not \U$27017 ( \27360 , \26243 );
or \U$27018 ( \27361 , \27359 , \27360 );
or \U$27019 ( \27362 , \26243 , \26259 );
nand \U$27020 ( \27363 , \27361 , \27362 );
not \U$27021 ( \27364 , \26227 );
and \U$27022 ( \27365 , \27363 , \27364 );
not \U$27023 ( \27366 , \27363 );
and \U$27024 ( \27367 , \27366 , \26227 );
nor \U$27025 ( \27368 , \27365 , \27367 );
not \U$27026 ( \27369 , \27368 );
not \U$27027 ( \27370 , \27369 );
not \U$27028 ( \27371 , \26307 );
not \U$27029 ( \27372 , \26329 );
not \U$27030 ( \27373 , \27372 );
or \U$27031 ( \27374 , \27371 , \27373 );
nand \U$27032 ( \27375 , \26310 , \26329 );
nand \U$27033 ( \27376 , \27374 , \27375 );
xor \U$27034 ( \27377 , \27376 , \26291 );
not \U$27035 ( \27378 , \27377 );
or \U$27036 ( \27379 , \27370 , \27378 );
or \U$27037 ( \27380 , \27369 , \27377 );
not \U$27038 ( \27381 , \6242 );
not \U$27039 ( \27382 , \26320 );
or \U$27040 ( \27383 , \27381 , \27382 );
not \U$27041 ( \27384 , RIbb2e530_37);
not \U$27042 ( \27385 , \22070 );
or \U$27043 ( \27386 , \27384 , \27385 );
nand \U$27044 ( \27387 , \12175 , \6246 );
nand \U$27045 ( \27388 , \27386 , \27387 );
nand \U$27046 ( \27389 , \27388 , \6251 );
nand \U$27047 ( \27390 , \27383 , \27389 );
not \U$27048 ( \27391 , \17100 );
not \U$27049 ( \27392 , \26280 );
or \U$27050 ( \27393 , \27391 , \27392 );
and \U$27051 ( \27394 , \14602 , \15443 );
not \U$27052 ( \27395 , \14602 );
and \U$27053 ( \27396 , \27395 , \19676 );
nor \U$27054 ( \27397 , \27394 , \27396 );
nand \U$27055 ( \27398 , \27397 , \16675 );
nand \U$27056 ( \27399 , \27393 , \27398 );
xor \U$27057 ( \27400 , \27390 , \27399 );
not \U$27058 ( \27401 , \18717 );
not \U$27059 ( \27402 , RIbb2d9f0_61);
not \U$27060 ( \27403 , \17568 );
or \U$27061 ( \27404 , \27402 , \27403 );
nand \U$27062 ( \27405 , \9707 , \21449 );
nand \U$27063 ( \27406 , \27404 , \27405 );
not \U$27064 ( \27407 , \27406 );
or \U$27065 ( \27408 , \27401 , \27407 );
nand \U$27066 ( \27409 , \26672 , \26834 );
nand \U$27067 ( \27410 , \27408 , \27409 );
and \U$27068 ( \27411 , \27400 , \27410 );
and \U$27069 ( \27412 , \27390 , \27399 );
or \U$27070 ( \27413 , \27411 , \27412 );
nand \U$27071 ( \27414 , \27380 , \27413 );
nand \U$27072 ( \27415 , \27379 , \27414 );
xor \U$27073 ( \27416 , \27358 , \27415 );
not \U$27074 ( \27417 , \26361 );
xor \U$27075 ( \27418 , \26345 , \27417 );
xor \U$27076 ( \27419 , \27418 , \26379 );
not \U$27077 ( \27420 , \27419 );
not \U$27078 ( \27421 , \27420 );
not \U$27079 ( \27422 , \27421 );
not \U$27080 ( \27423 , \27422 );
xor \U$27081 ( \27424 , \26659 , \26674 );
xor \U$27082 ( \27425 , \27424 , \26690 );
not \U$27083 ( \27426 , \27425 );
or \U$27084 ( \27427 , \27423 , \27426 );
not \U$27085 ( \27428 , \27425 );
not \U$27086 ( \27429 , \27428 );
not \U$27087 ( \27430 , \27421 );
or \U$27088 ( \27431 , \27429 , \27430 );
xor \U$27089 ( \27432 , \27217 , \27244 );
xor \U$27090 ( \27433 , \27432 , \27255 );
not \U$27091 ( \27434 , \16271 );
and \U$27092 ( \27435 , RIbb2dae0_59, \3905 );
not \U$27093 ( \27436 , RIbb2dae0_59);
not \U$27094 ( \27437 , \6173 );
and \U$27095 ( \27438 , \27436 , \27437 );
or \U$27096 ( \27439 , \27435 , \27438 );
not \U$27097 ( \27440 , \27439 );
or \U$27098 ( \27441 , \27434 , \27440 );
nand \U$27099 ( \27442 , \26337 , \17470 );
nand \U$27100 ( \27443 , \27441 , \27442 );
xor \U$27101 ( \27444 , \27433 , \27443 );
xor \U$27102 ( \27445 , \27218 , \27229 );
xor \U$27103 ( \27446 , \27445 , \27241 );
not \U$27104 ( \27447 , \3886 );
not \U$27105 ( \27448 , RIbb2e710_33);
not \U$27106 ( \27449 , \14506 );
not \U$27107 ( \27450 , \27449 );
or \U$27108 ( \27451 , \27448 , \27450 );
nand \U$27109 ( \27452 , \13977 , \6844 );
nand \U$27110 ( \27453 , \27451 , \27452 );
not \U$27111 ( \27454 , \27453 );
or \U$27112 ( \27455 , \27447 , \27454 );
nand \U$27113 ( \27456 , \27253 , \4075 );
nand \U$27114 ( \27457 , \27455 , \27456 );
xor \U$27115 ( \27458 , \27446 , \27457 );
not \U$27116 ( \27459 , \6241 );
not \U$27117 ( \27460 , \27388 );
or \U$27118 ( \27461 , \27459 , \27460 );
and \U$27119 ( \27462 , \16865 , RIbb2e530_37);
not \U$27120 ( \27463 , \16865 );
and \U$27121 ( \27464 , \27463 , \4708 );
or \U$27122 ( \27465 , \27462 , \27464 );
nand \U$27123 ( \27466 , \27465 , \6251 );
nand \U$27124 ( \27467 , \27461 , \27466 );
and \U$27125 ( \27468 , \27458 , \27467 );
and \U$27126 ( \27469 , \27446 , \27457 );
or \U$27127 ( \27470 , \27468 , \27469 );
and \U$27128 ( \27471 , \27444 , \27470 );
and \U$27129 ( \27472 , \27433 , \27443 );
or \U$27130 ( \27473 , \27471 , \27472 );
nand \U$27131 ( \27474 , \27431 , \27473 );
nand \U$27132 ( \27475 , \27427 , \27474 );
and \U$27133 ( \27476 , \27416 , \27475 );
and \U$27134 ( \27477 , \27358 , \27415 );
or \U$27135 ( \27478 , \27476 , \27477 );
not \U$27136 ( \27479 , \27478 );
not \U$27137 ( \27480 , \26432 );
not \U$27138 ( \27481 , \26696 );
or \U$27139 ( \27482 , \27480 , \27481 );
or \U$27140 ( \27483 , \26432 , \26696 );
nand \U$27141 ( \27484 , \27482 , \27483 );
and \U$27142 ( \27485 , \27484 , \26526 );
not \U$27143 ( \27486 , \27484 );
and \U$27144 ( \27487 , \27486 , \26699 );
nor \U$27145 ( \27488 , \27485 , \27487 );
not \U$27146 ( \27489 , \27488 );
not \U$27147 ( \27490 , \27489 );
or \U$27148 ( \27491 , \27479 , \27490 );
or \U$27149 ( \27492 , \27478 , \27489 );
not \U$27150 ( \27493 , \11176 );
not \U$27151 ( \27494 , RIbb2e080_47);
not \U$27152 ( \27495 , \19868 );
or \U$27153 ( \27496 , \27494 , \27495 );
nand \U$27154 ( \27497 , \8637 , \10113 );
nand \U$27155 ( \27498 , \27496 , \27497 );
not \U$27156 ( \27499 , \27498 );
or \U$27157 ( \27500 , \27493 , \27499 );
nand \U$27158 ( \27501 , \26225 , \11177 );
nand \U$27159 ( \27502 , \27500 , \27501 );
not \U$27160 ( \27503 , \10119 );
not \U$27161 ( \27504 , \26241 );
or \U$27162 ( \27505 , \27503 , \27504 );
not \U$27163 ( \27506 , RIbb2e170_45);
not \U$27164 ( \27507 , \8318 );
not \U$27165 ( \27508 , \27507 );
or \U$27166 ( \27509 , \27506 , \27508 );
nand \U$27167 ( \27510 , \14024 , \9094 );
nand \U$27168 ( \27511 , \27509 , \27510 );
nand \U$27169 ( \27512 , \27511 , \10117 );
nand \U$27170 ( \27513 , \27505 , \27512 );
xor \U$27171 ( \27514 , \27502 , \27513 );
not \U$27172 ( \27515 , \26560 );
not \U$27173 ( \27516 , \16427 );
or \U$27174 ( \27517 , \27515 , \27516 );
not \U$27175 ( \27518 , RIbb2df90_49);
not \U$27176 ( \27519 , \21570 );
or \U$27177 ( \27520 , \27518 , \27519 );
not \U$27178 ( \27521 , \18564 );
nand \U$27179 ( \27522 , \27521 , \12278 );
nand \U$27180 ( \27523 , \27520 , \27522 );
nand \U$27181 ( \27524 , \27523 , \13295 );
nand \U$27182 ( \27525 , \27517 , \27524 );
and \U$27183 ( \27526 , \27514 , \27525 );
and \U$27184 ( \27527 , \27502 , \27513 );
or \U$27185 ( \27528 , \27526 , \27527 );
not \U$27186 ( \27529 , \27528 );
buf \U$27187 ( \27530 , \26562 );
not \U$27188 ( \27531 , \27530 );
not \U$27189 ( \27532 , \26538 );
not \U$27190 ( \27533 , \26550 );
and \U$27191 ( \27534 , \27532 , \27533 );
and \U$27192 ( \27535 , \26538 , \26550 );
nor \U$27193 ( \27536 , \27534 , \27535 );
not \U$27194 ( \27537 , \27536 );
and \U$27195 ( \27538 , \27531 , \27537 );
and \U$27196 ( \27539 , \27530 , \27536 );
nor \U$27197 ( \27540 , \27538 , \27539 );
nand \U$27198 ( \27541 , \27529 , \27540 );
not \U$27199 ( \27542 , \27541 );
xor \U$27200 ( \27543 , \26181 , \26191 );
xor \U$27201 ( \27544 , \27543 , \26202 );
not \U$27202 ( \27545 , \27544 );
or \U$27203 ( \27546 , \27542 , \27545 );
not \U$27204 ( \27547 , \27540 );
xor \U$27205 ( \27548 , \27502 , \27513 );
and \U$27206 ( \27549 , \27548 , \27525 );
and \U$27207 ( \27550 , \27502 , \27513 );
or \U$27208 ( \27551 , \27549 , \27550 );
nand \U$27209 ( \27552 , \27547 , \27551 );
nand \U$27210 ( \27553 , \27546 , \27552 );
xor \U$27211 ( \27554 , \26566 , \26641 );
xor \U$27212 ( \27555 , \27554 , \26693 );
xor \U$27213 ( \27556 , \27553 , \27555 );
xor \U$27214 ( \27557 , \26610 , \26623 );
xor \U$27215 ( \27558 , \27557 , \26638 );
or \U$27216 ( \27559 , RIbb2eb48_24, RIbb2ead0_25);
nand \U$27217 ( \27560 , \27559 , \19064 );
and \U$27218 ( \27561 , RIbb2eb48_24, RIbb2ead0_25);
nor \U$27219 ( \27562 , \27561 , \2073 );
and \U$27220 ( \27563 , \27560 , \27562 );
not \U$27221 ( \27564 , \3381 );
not \U$27222 ( \27565 , \27227 );
or \U$27223 ( \27566 , \27564 , \27565 );
or \U$27224 ( \27567 , \17506 , \3388 );
or \U$27225 ( \27568 , \18929 , RIbb2ebc0_23);
nand \U$27226 ( \27569 , \27567 , \27568 );
nand \U$27227 ( \27570 , \27569 , \3405 );
nand \U$27228 ( \27571 , \27566 , \27570 );
and \U$27229 ( \27572 , \27563 , \27571 );
not \U$27230 ( \27573 , \3465 );
not \U$27231 ( \27574 , \26598 );
or \U$27232 ( \27575 , \27573 , \27574 );
not \U$27233 ( \27576 , RIbb2e9e0_27);
not \U$27234 ( \27577 , \19831 );
not \U$27235 ( \27578 , \27577 );
or \U$27236 ( \27579 , \27576 , \27578 );
nand \U$27237 ( \27580 , \16829 , \3454 );
nand \U$27238 ( \27581 , \27579 , \27580 );
nand \U$27239 ( \27582 , \27581 , \3445 );
nand \U$27240 ( \27583 , \27575 , \27582 );
xor \U$27241 ( \27584 , \27572 , \27583 );
not \U$27242 ( \27585 , \2925 );
not \U$27243 ( \27586 , \27190 );
or \U$27244 ( \27587 , \27585 , \27586 );
not \U$27245 ( \27588 , RIbb2e8f0_29);
not \U$27246 ( \27589 , \16844 );
or \U$27247 ( \27590 , \27588 , \27589 );
nand \U$27248 ( \27591 , \16576 , \3800 );
nand \U$27249 ( \27592 , \27590 , \27591 );
nand \U$27250 ( \27593 , \27592 , \2922 );
nand \U$27251 ( \27594 , \27587 , \27593 );
and \U$27252 ( \27595 , \27584 , \27594 );
and \U$27253 ( \27596 , \27572 , \27583 );
or \U$27254 ( \27597 , \27595 , \27596 );
not \U$27255 ( \27598 , \8354 );
not \U$27256 ( \27599 , \26305 );
or \U$27257 ( \27600 , \27598 , \27599 );
and \U$27258 ( \27601 , RIbb2e350_41, \12234 );
not \U$27259 ( \27602 , RIbb2e350_41);
and \U$27260 ( \27603 , \27602 , \12235 );
nor \U$27261 ( \27604 , \27601 , \27603 );
not \U$27262 ( \27605 , \27604 );
nand \U$27263 ( \27606 , \27605 , \8362 );
nand \U$27264 ( \27607 , \27600 , \27606 );
xor \U$27265 ( \27608 , \27597 , \27607 );
not \U$27266 ( \27609 , \7103 );
not \U$27267 ( \27610 , RIbb2e440_39);
not \U$27268 ( \27611 , \15188 );
or \U$27269 ( \27612 , \27610 , \27611 );
not \U$27270 ( \27613 , RIbb2e440_39);
nand \U$27271 ( \27614 , \27613 , \13692 );
nand \U$27272 ( \27615 , \27612 , \27614 );
not \U$27273 ( \27616 , \27615 );
or \U$27274 ( \27617 , \27609 , \27616 );
nand \U$27275 ( \27618 , \26615 , \8450 );
nand \U$27276 ( \27619 , \27617 , \27618 );
and \U$27277 ( \27620 , \27608 , \27619 );
and \U$27278 ( \27621 , \27597 , \27607 );
or \U$27279 ( \27622 , \27620 , \27621 );
xor \U$27280 ( \27623 , \27558 , \27622 );
not \U$27281 ( \27624 , \15688 );
not \U$27282 ( \27625 , \26377 );
or \U$27283 ( \27626 , \27624 , \27625 );
not \U$27284 ( \27627 , RIbb2ddb0_53);
not \U$27285 ( \27628 , \19429 );
or \U$27286 ( \27629 , \27627 , \27628 );
nand \U$27287 ( \27630 , \4086 , \12681 );
nand \U$27288 ( \27631 , \27629 , \27630 );
nand \U$27289 ( \27632 , \27631 , \17562 );
nand \U$27290 ( \27633 , \27626 , \27632 );
not \U$27291 ( \27634 , \22952 );
and \U$27292 ( \27635 , RIbb2dcc0_55, \13731 );
not \U$27293 ( \27636 , RIbb2dcc0_55);
and \U$27294 ( \27637 , \27636 , \3274 );
or \U$27295 ( \27638 , \27635 , \27637 );
not \U$27296 ( \27639 , \27638 );
or \U$27297 ( \27640 , \27634 , \27639 );
nand \U$27298 ( \27641 , \26688 , \15181 );
nand \U$27299 ( \27642 , \27640 , \27641 );
xor \U$27300 ( \27643 , \27633 , \27642 );
not \U$27301 ( \27644 , \17275 );
and \U$27302 ( \27645 , RIbb2d900_63, \12097 );
not \U$27303 ( \27646 , RIbb2d900_63);
and \U$27304 ( \27647 , \27646 , \3521 );
or \U$27305 ( \27648 , \27645 , \27647 );
not \U$27306 ( \27649 , \27648 );
or \U$27307 ( \27650 , \27644 , \27649 );
nand \U$27308 ( \27651 , \26352 , RIbb2d888_64);
nand \U$27309 ( \27652 , \27650 , \27651 );
and \U$27310 ( \27653 , \27643 , \27652 );
and \U$27311 ( \27654 , \27633 , \27642 );
or \U$27312 ( \27655 , \27653 , \27654 );
and \U$27313 ( \27656 , \27623 , \27655 );
and \U$27314 ( \27657 , \27558 , \27622 );
or \U$27315 ( \27658 , \27656 , \27657 );
and \U$27316 ( \27659 , \27556 , \27658 );
and \U$27317 ( \27660 , \27553 , \27555 );
or \U$27318 ( \27661 , \27659 , \27660 );
buf \U$27319 ( \27662 , \27661 );
nand \U$27320 ( \27663 , \27492 , \27662 );
nand \U$27321 ( \27664 , \27491 , \27663 );
not \U$27322 ( \27665 , \27664 );
nand \U$27323 ( \27666 , \27356 , \27665 );
not \U$27324 ( \27667 , \27666 );
or \U$27325 ( \27668 , \27343 , \27667 );
not \U$27326 ( \27669 , \27356 );
nand \U$27327 ( \27670 , \27669 , \27664 );
nand \U$27328 ( \27671 , \27668 , \27670 );
xor \U$27329 ( \27672 , \27111 , \27671 );
not \U$27330 ( \27673 , \27345 );
or \U$27331 ( \27674 , \27354 , \27673 );
nand \U$27332 ( \27675 , \27674 , \27351 );
nand \U$27333 ( \27676 , \27354 , \27673 );
nand \U$27334 ( \27677 , \27675 , \27676 );
xor \U$27335 ( \27678 , \26954 , \26958 );
and \U$27336 ( \27679 , \27678 , \26992 );
and \U$27337 ( \27680 , \26954 , \26958 );
or \U$27338 ( \27681 , \27679 , \27680 );
nor \U$27339 ( \27682 , \27057 , \27000 );
not \U$27340 ( \27683 , \27027 );
or \U$27341 ( \27684 , \27682 , \27683 );
nand \U$27342 ( \27685 , \27057 , \27000 );
nand \U$27343 ( \27686 , \27684 , \27685 );
xor \U$27344 ( \27687 , \27681 , \27686 );
not \U$27345 ( \27688 , \26145 );
not \U$27346 ( \27689 , \26161 );
or \U$27347 ( \27690 , \27688 , \27689 );
or \U$27348 ( \27691 , \26161 , \26145 );
nand \U$27349 ( \27692 , \27691 , \26140 );
nand \U$27350 ( \27693 , \27690 , \27692 );
not \U$27351 ( \27694 , \8450 );
not \U$27352 ( \27695 , \25832 );
or \U$27353 ( \27696 , \27694 , \27695 );
nand \U$27354 ( \27697 , \27011 , \8445 );
nand \U$27355 ( \27698 , \27696 , \27697 );
xor \U$27356 ( \27699 , \27693 , \27698 );
not \U$27357 ( \27700 , \6242 );
not \U$27358 ( \27701 , \25935 );
or \U$27359 ( \27702 , \27700 , \27701 );
nand \U$27360 ( \27703 , \27283 , \6251 );
nand \U$27361 ( \27704 , \27702 , \27703 );
xnor \U$27362 ( \27705 , \27699 , \27704 );
not \U$27363 ( \27706 , \27705 );
not \U$27364 ( \27707 , \4075 );
not \U$27365 ( \27708 , RIbb2e710_33);
not \U$27366 ( \27709 , \14886 );
or \U$27367 ( \27710 , \27708 , \27709 );
nand \U$27368 ( \27711 , \14885 , \6058 );
nand \U$27369 ( \27712 , \27710 , \27711 );
not \U$27370 ( \27713 , \27712 );
or \U$27371 ( \27714 , \27707 , \27713 );
nand \U$27372 ( \27715 , \26899 , \3886 );
nand \U$27373 ( \27716 , \27714 , \27715 );
not \U$27374 ( \27717 , \27716 );
not \U$27375 ( \27718 , \10599 );
not \U$27376 ( \27719 , \27050 );
or \U$27377 ( \27720 , \27718 , \27719 );
nand \U$27378 ( \27721 , \25873 , \10119 );
nand \U$27379 ( \27722 , \27720 , \27721 );
not \U$27380 ( \27723 , \27722 );
not \U$27381 ( \27724 , \27723 );
or \U$27382 ( \27725 , \27717 , \27724 );
or \U$27383 ( \27726 , \27716 , \27723 );
nand \U$27384 ( \27727 , \27725 , \27726 );
not \U$27385 ( \27728 , \11176 );
not \U$27386 ( \27729 , \26911 );
or \U$27387 ( \27730 , \27728 , \27729 );
nand \U$27388 ( \27731 , \25904 , \12965 );
nand \U$27389 ( \27732 , \27730 , \27731 );
not \U$27390 ( \27733 , \27732 );
and \U$27391 ( \27734 , \27727 , \27733 );
not \U$27392 ( \27735 , \27727 );
and \U$27393 ( \27736 , \27735 , \27732 );
nor \U$27394 ( \27737 , \27734 , \27736 );
not \U$27395 ( \27738 , \27737 );
or \U$27396 ( \27739 , \27706 , \27738 );
xor \U$27397 ( \27740 , \25792 , \25807 );
xor \U$27398 ( \27741 , \27740 , \25824 );
not \U$27399 ( \27742 , \9099 );
not \U$27400 ( \27743 , \25881 );
or \U$27401 ( \27744 , \27742 , \27743 );
nand \U$27402 ( \27745 , \27036 , \9098 );
nand \U$27403 ( \27746 , \27744 , \27745 );
xor \U$27404 ( \27747 , \27741 , \27746 );
not \U$27405 ( \27748 , \8362 );
not \U$27406 ( \27749 , \27020 );
or \U$27407 ( \27750 , \27748 , \27749 );
not \U$27408 ( \27751 , \25856 );
or \U$27409 ( \27752 , \27751 , \8355 );
nand \U$27410 ( \27753 , \27750 , \27752 );
xor \U$27411 ( \27754 , \27747 , \27753 );
nand \U$27412 ( \27755 , \27739 , \27754 );
not \U$27413 ( \27756 , \27737 );
not \U$27414 ( \27757 , \27705 );
nand \U$27415 ( \27758 , \27756 , \27757 );
nand \U$27416 ( \27759 , \27755 , \27758 );
xor \U$27417 ( \27760 , \27687 , \27759 );
xor \U$27418 ( \27761 , \26970 , \26979 );
and \U$27419 ( \27762 , \27761 , \26991 );
and \U$27420 ( \27763 , \26970 , \26979 );
or \U$27421 ( \27764 , \27762 , \27763 );
not \U$27422 ( \27765 , \2922 );
not \U$27423 ( \27766 , \26966 );
or \U$27424 ( \27767 , \27765 , \27766 );
not \U$27425 ( \27768 , RIbb2e8f0_29);
not \U$27426 ( \27769 , \14838 );
or \U$27427 ( \27770 , \27768 , \27769 );
nand \U$27428 ( \27771 , \12347 , \3265 );
nand \U$27429 ( \27772 , \27770 , \27771 );
nand \U$27430 ( \27773 , \27772 , \2925 );
nand \U$27431 ( \27774 , \27767 , \27773 );
not \U$27432 ( \27775 , \3613 );
not \U$27433 ( \27776 , RIbb2e800_31);
not \U$27434 ( \27777 , \13680 );
or \U$27435 ( \27778 , \27776 , \27777 );
nand \U$27436 ( \27779 , \12838 , \2917 );
nand \U$27437 ( \27780 , \27778 , \27779 );
not \U$27438 ( \27781 , \27780 );
or \U$27439 ( \27782 , \27775 , \27781 );
nand \U$27440 ( \27783 , \26987 , \2939 );
nand \U$27441 ( \27784 , \27782 , \27783 );
xor \U$27442 ( \27785 , \27774 , \27784 );
not \U$27443 ( \27786 , \4791 );
not \U$27444 ( \27787 , RIbb2e710_33);
not \U$27445 ( \27788 , \17294 );
or \U$27446 ( \27789 , \27787 , \27788 );
nand \U$27447 ( \27790 , \12261 , \6844 );
nand \U$27448 ( \27791 , \27789 , \27790 );
not \U$27449 ( \27792 , \27791 );
or \U$27450 ( \27793 , \27786 , \27792 );
nand \U$27451 ( \27794 , \27712 , \3886 );
nand \U$27452 ( \27795 , \27793 , \27794 );
xor \U$27453 ( \27796 , \27785 , \27795 );
xor \U$27454 ( \27797 , \27764 , \27796 );
or \U$27455 ( \27798 , \27704 , \27698 );
nand \U$27456 ( \27799 , \27798 , \27693 );
nand \U$27457 ( \27800 , \27704 , \27698 );
nand \U$27458 ( \27801 , \27799 , \27800 );
xor \U$27459 ( \27802 , \27797 , \27801 );
and \U$27460 ( \27803 , \17506 , \1517 );
not \U$27461 ( \27804 , \835 );
not \U$27462 ( \27805 , RIbb2ee90_17);
not \U$27463 ( \27806 , \16819 );
or \U$27464 ( \27807 , \27805 , \27806 );
nand \U$27465 ( \27808 , \17529 , \3057 );
nand \U$27466 ( \27809 , \27807 , \27808 );
not \U$27467 ( \27810 , \27809 );
or \U$27468 ( \27811 , \27804 , \27810 );
nand \U$27469 ( \27812 , \25783 , \831 );
nand \U$27470 ( \27813 , \27811 , \27812 );
xor \U$27471 ( \27814 , \27803 , \27813 );
not \U$27472 ( \27815 , \853 );
not \U$27473 ( \27816 , \25798 );
or \U$27474 ( \27817 , \27815 , \27816 );
not \U$27475 ( \27818 , RIbb2eda0_19);
not \U$27476 ( \27819 , \16554 );
or \U$27477 ( \27820 , \27818 , \27819 );
nand \U$27478 ( \27821 , \16706 , \5277 );
nand \U$27479 ( \27822 , \27820 , \27821 );
nand \U$27480 ( \27823 , \27822 , \854 );
nand \U$27481 ( \27824 , \27817 , \27823 );
xor \U$27482 ( \27825 , \27814 , \27824 );
not \U$27483 ( \27826 , \3445 );
not \U$27484 ( \27827 , \26789 );
or \U$27485 ( \27828 , \27826 , \27827 );
not \U$27486 ( \27829 , RIbb2e9e0_27);
not \U$27487 ( \27830 , \13546 );
or \U$27488 ( \27831 , \27829 , \27830 );
nand \U$27489 ( \27832 , \13545 , \3454 );
nand \U$27490 ( \27833 , \27831 , \27832 );
nand \U$27491 ( \27834 , \27833 , \3465 );
nand \U$27492 ( \27835 , \27828 , \27834 );
xor \U$27493 ( \27836 , \27825 , \27835 );
not \U$27494 ( \27837 , \2963 );
and \U$27495 ( \27838 , RIbb2ead0_25, \21770 );
not \U$27496 ( \27839 , RIbb2ead0_25);
and \U$27497 ( \27840 , \27839 , \15036 );
or \U$27498 ( \27841 , \27838 , \27840 );
not \U$27499 ( \27842 , \27841 );
or \U$27500 ( \27843 , \27837 , \27842 );
nand \U$27501 ( \27844 , \26975 , \2980 );
nand \U$27502 ( \27845 , \27843 , \27844 );
xor \U$27503 ( \27846 , \27836 , \27845 );
xor \U$27504 ( \27847 , \27741 , \27746 );
and \U$27505 ( \27848 , \27847 , \27753 );
and \U$27506 ( \27849 , \27741 , \27746 );
or \U$27507 ( \27850 , \27848 , \27849 );
xor \U$27508 ( \27851 , \27846 , \27850 );
nor \U$27509 ( \27852 , \27732 , \27716 );
or \U$27510 ( \27853 , \27852 , \27723 );
nand \U$27511 ( \27854 , \27732 , \27716 );
nand \U$27512 ( \27855 , \27853 , \27854 );
xor \U$27513 ( \27856 , \27851 , \27855 );
xor \U$27514 ( \27857 , \27802 , \27856 );
xor \U$27515 ( \27858 , \27271 , \27276 );
and \U$27516 ( \27859 , \27858 , \27287 );
and \U$27517 ( \27860 , \27271 , \27276 );
or \U$27518 ( \27861 , \27859 , \27860 );
not \U$27519 ( \27862 , \26173 );
not \U$27520 ( \27863 , \26119 );
or \U$27521 ( \27864 , \27862 , \27863 );
or \U$27522 ( \27865 , \26119 , \26173 );
not \U$27523 ( \27866 , \26162 );
nand \U$27524 ( \27867 , \27865 , \27866 );
nand \U$27525 ( \27868 , \27864 , \27867 );
xor \U$27526 ( \27869 , \27861 , \27868 );
xor \U$27527 ( \27870 , \27298 , \27303 );
and \U$27528 ( \27871 , \27870 , \27309 );
and \U$27529 ( \27872 , \27298 , \27303 );
or \U$27530 ( \27873 , \27871 , \27872 );
and \U$27531 ( \27874 , \27869 , \27873 );
and \U$27532 ( \27875 , \27861 , \27868 );
or \U$27533 ( \27876 , \27874 , \27875 );
xor \U$27534 ( \27877 , \27857 , \27876 );
xor \U$27535 ( \27878 , \27760 , \27877 );
not \U$27536 ( \27879 , \27288 );
not \U$27537 ( \27880 , \27310 );
or \U$27538 ( \27881 , \27879 , \27880 );
or \U$27539 ( \27882 , \27310 , \27288 );
nand \U$27540 ( \27883 , \27882 , \27292 );
nand \U$27541 ( \27884 , \27881 , \27883 );
not \U$27542 ( \27885 , \27884 );
xor \U$27543 ( \27886 , \27861 , \27868 );
xor \U$27544 ( \27887 , \27886 , \27873 );
not \U$27545 ( \27888 , \27887 );
or \U$27546 ( \27889 , \27885 , \27888 );
or \U$27547 ( \27890 , \27887 , \27884 );
not \U$27548 ( \27891 , \27754 );
not \U$27549 ( \27892 , \27737 );
or \U$27550 ( \27893 , \27891 , \27892 );
or \U$27551 ( \27894 , \27737 , \27754 );
nand \U$27552 ( \27895 , \27893 , \27894 );
and \U$27553 ( \27896 , \27895 , \27705 );
not \U$27554 ( \27897 , \27895 );
and \U$27555 ( \27898 , \27897 , \27757 );
nor \U$27556 ( \27899 , \27896 , \27898 );
not \U$27557 ( \27900 , \27899 );
nand \U$27558 ( \27901 , \27890 , \27900 );
nand \U$27559 ( \27902 , \27889 , \27901 );
xor \U$27560 ( \27903 , \27878 , \27902 );
xor \U$27561 ( \27904 , \27677 , \27903 );
not \U$27562 ( \27905 , \27900 );
xor \U$27563 ( \27906 , \27861 , \27868 );
xnor \U$27564 ( \27907 , \27906 , \27873 );
not \U$27565 ( \27908 , \27907 );
or \U$27566 ( \27909 , \27905 , \27908 );
nand \U$27567 ( \27910 , \27899 , \27887 );
nand \U$27568 ( \27911 , \27909 , \27910 );
xor \U$27569 ( \27912 , \27911 , \27884 );
not \U$27570 ( \27913 , \27264 );
not \U$27571 ( \27914 , \27312 );
or \U$27572 ( \27915 , \27913 , \27914 );
or \U$27573 ( \27916 , \27312 , \27264 );
nand \U$27574 ( \27917 , \27916 , \27322 );
nand \U$27575 ( \27918 , \27915 , \27917 );
xor \U$27576 ( \27919 , \27912 , \27918 );
xor \U$27577 ( \27920 , \26270 , \26272 );
xor \U$27578 ( \27921 , \27920 , \26701 );
and \U$27579 ( \27922 , \27919 , \27921 );
and \U$27580 ( \27923 , \27912 , \27918 );
or \U$27581 ( \27924 , \27922 , \27923 );
xor \U$27582 ( \27925 , \27904 , \27924 );
and \U$27583 ( \27926 , \27672 , \27925 );
and \U$27584 ( \27927 , \27111 , \27671 );
or \U$27585 ( \27928 , \27926 , \27927 );
not \U$27586 ( \27929 , \27928 );
not \U$27587 ( \27930 , \17275 );
not \U$27588 ( \27931 , \26739 );
or \U$27589 ( \27932 , \27930 , \27931 );
not \U$27590 ( \27933 , RIbb2d900_63);
not \U$27591 ( \27934 , \17369 );
or \U$27592 ( \27935 , \27933 , \27934 );
nand \U$27593 ( \27936 , \1169 , \17262 );
nand \U$27594 ( \27937 , \27935 , \27936 );
nand \U$27595 ( \27938 , \27937 , RIbb2d888_64);
nand \U$27596 ( \27939 , \27932 , \27938 );
not \U$27597 ( \27940 , \11177 );
not \U$27598 ( \27941 , RIbb2e080_47);
not \U$27599 ( \27942 , \3090 );
or \U$27600 ( \27943 , \27941 , \27942 );
nand \U$27601 ( \27944 , \3089 , \10113 );
nand \U$27602 ( \27945 , \27943 , \27944 );
not \U$27603 ( \27946 , \27945 );
or \U$27604 ( \27947 , \27940 , \27946 );
nand \U$27605 ( \27948 , \25897 , \11176 );
nand \U$27606 ( \27949 , \27947 , \27948 );
xor \U$27607 ( \27950 , \27939 , \27949 );
not \U$27608 ( \27951 , \14613 );
not \U$27609 ( \27952 , \26853 );
or \U$27610 ( \27953 , \27951 , \27952 );
not \U$27611 ( \27954 , \15181 );
not \U$27612 ( \27955 , \27954 );
and \U$27613 ( \27956 , RIbb2dcc0_55, \3952 );
not \U$27614 ( \27957 , RIbb2dcc0_55);
and \U$27615 ( \27958 , \27957 , \3951 );
or \U$27616 ( \27959 , \27956 , \27958 );
nand \U$27617 ( \27960 , \27955 , \27959 );
nand \U$27618 ( \27961 , \27953 , \27960 );
xor \U$27619 ( \27962 , \27950 , \27961 );
not \U$27620 ( \27963 , \5845 );
not \U$27621 ( \27964 , RIbb2e620_35);
not \U$27622 ( \27965 , \22580 );
or \U$27623 ( \27966 , \27964 , \27965 );
nand \U$27624 ( \27967 , \9841 , \6688 );
nand \U$27625 ( \27968 , \27966 , \27967 );
not \U$27626 ( \27969 , \27968 );
or \U$27627 ( \27970 , \27963 , \27969 );
nand \U$27628 ( \27971 , \25919 , \4712 );
nand \U$27629 ( \27972 , \27970 , \27971 );
not \U$27630 ( \27973 , \19101 );
not \U$27631 ( \27974 , \26842 );
or \U$27632 ( \27975 , \27973 , \27974 );
not \U$27633 ( \27976 , RIbb2dbd0_57);
not \U$27634 ( \27977 , \13286 );
or \U$27635 ( \27978 , \27976 , \27977 );
nand \U$27636 ( \27979 , \13290 , \17411 );
nand \U$27637 ( \27980 , \27978 , \27979 );
nand \U$27638 ( \27981 , \27980 , \17100 );
nand \U$27639 ( \27982 , \27975 , \27981 );
xor \U$27640 ( \27983 , \27972 , \27982 );
not \U$27641 ( \27984 , \12167 );
not \U$27642 ( \27985 , \25946 );
or \U$27643 ( \27986 , \27984 , \27985 );
not \U$27644 ( \27987 , RIbb2df90_49);
not \U$27645 ( \27988 , \13738 );
or \U$27646 ( \27989 , \27987 , \27988 );
nand \U$27647 ( \27990 , \16185 , \12278 );
nand \U$27648 ( \27991 , \27989 , \27990 );
nand \U$27649 ( \27992 , \12285 , \27991 );
nand \U$27650 ( \27993 , \27986 , \27992 );
xor \U$27651 ( \27994 , \27983 , \27993 );
xor \U$27652 ( \27995 , \27962 , \27994 );
not \U$27653 ( \27996 , \2077 );
not \U$27654 ( \27997 , \26712 );
or \U$27655 ( \27998 , \27996 , \27997 );
not \U$27656 ( \27999 , RIbb2ecb0_21);
not \U$27657 ( \28000 , \23197 );
or \U$27658 ( \28001 , \27999 , \28000 );
nand \U$27659 ( \28002 , \16575 , \849 );
nand \U$27660 ( \28003 , \28001 , \28002 );
nand \U$27661 ( \28004 , \28003 , \2078 );
nand \U$27662 ( \28005 , \27998 , \28004 );
xor \U$27663 ( \28006 , \27803 , \27813 );
and \U$27664 ( \28007 , \28006 , \27824 );
and \U$27665 ( \28008 , \27803 , \27813 );
or \U$27666 ( \28009 , \28007 , \28008 );
xor \U$27667 ( \28010 , \28005 , \28009 );
not \U$27668 ( \28011 , \2925 );
not \U$27669 ( \28012 , RIbb2e8f0_29);
not \U$27670 ( \28013 , \16865 );
or \U$27671 ( \28014 , \28012 , \28013 );
nand \U$27672 ( \28015 , \12932 , \4800 );
nand \U$27673 ( \28016 , \28014 , \28015 );
not \U$27674 ( \28017 , \28016 );
or \U$27675 ( \28018 , \28011 , \28017 );
nand \U$27676 ( \28019 , \27772 , \2922 );
nand \U$27677 ( \28020 , \28018 , \28019 );
xor \U$27678 ( \28021 , \28010 , \28020 );
xor \U$27679 ( \28022 , \27825 , \27835 );
and \U$27680 ( \28023 , \28022 , \27845 );
and \U$27681 ( \28024 , \27825 , \27835 );
or \U$27682 ( \28025 , \28023 , \28024 );
xor \U$27683 ( \28026 , \28021 , \28025 );
not \U$27684 ( \28027 , \14067 );
not \U$27685 ( \28028 , \26817 );
or \U$27686 ( \28029 , \28027 , \28028 );
not \U$27687 ( \28030 , RIbb2dea0_51);
not \U$27688 ( \28031 , \16898 );
or \U$27689 ( \28032 , \28030 , \28031 );
not \U$27690 ( \28033 , RIbb2dea0_51);
nand \U$27691 ( \28034 , \28033 , \25703 );
nand \U$27692 ( \28035 , \28032 , \28034 );
nand \U$27693 ( \28036 , \28035 , \12692 );
nand \U$27694 ( \28037 , \28029 , \28036 );
xor \U$27695 ( \28038 , \28026 , \28037 );
buf \U$27696 ( \28039 , \28038 );
and \U$27697 ( \28040 , \27995 , \28039 );
not \U$27698 ( \28041 , \27995 );
not \U$27699 ( \28042 , \28039 );
and \U$27700 ( \28043 , \28041 , \28042 );
nor \U$27701 ( \28044 , \28040 , \28043 );
xor \U$27702 ( \28045 , \26757 , \26823 );
and \U$27703 ( \28046 , \28045 , \26858 );
and \U$27704 ( \28047 , \26757 , \26823 );
or \U$27705 ( \28048 , \28046 , \28047 );
xor \U$27706 ( \28049 , \26706 , \26721 );
and \U$27707 ( \28050 , \28049 , \26732 );
and \U$27708 ( \28051 , \26706 , \26721 );
or \U$27709 ( \28052 , \28050 , \28051 );
not \U$27710 ( \28053 , \8445 );
not \U$27711 ( \28054 , \25838 );
or \U$27712 ( \28055 , \28053 , \28054 );
and \U$27713 ( \28056 , RIbb2e440_39, \14672 );
not \U$27714 ( \28057 , RIbb2e440_39);
and \U$27715 ( \28058 , \28057 , \7296 );
or \U$27716 ( \28059 , \28056 , \28058 );
nand \U$27717 ( \28060 , \28059 , \7104 );
nand \U$27718 ( \28061 , \28055 , \28060 );
xor \U$27719 ( \28062 , \28052 , \28061 );
not \U$27720 ( \28063 , \6251 );
not \U$27721 ( \28064 , \25927 );
or \U$27722 ( \28065 , \28063 , \28064 );
not \U$27723 ( \28066 , RIbb2e530_37);
not \U$27724 ( \28067 , \13863 );
or \U$27725 ( \28068 , \28066 , \28067 );
nand \U$27726 ( \28069 , \8630 , \6246 );
nand \U$27727 ( \28070 , \28068 , \28069 );
nand \U$27728 ( \28071 , \28070 , \6242 );
nand \U$27729 ( \28072 , \28065 , \28071 );
xor \U$27730 ( \28073 , \28062 , \28072 );
not \U$27731 ( \28074 , \1517 );
and \U$27732 ( \28075 , RIbb2ef80_15, \20552 );
not \U$27733 ( \28076 , RIbb2ef80_15);
and \U$27734 ( \28077 , \28076 , \26129 );
or \U$27735 ( \28078 , \28075 , \28077 );
not \U$27736 ( \28079 , \28078 );
or \U$27737 ( \28080 , \28074 , \28079 );
and \U$27738 ( \28081 , RIbb2ef80_15, \19064 );
not \U$27739 ( \28082 , RIbb2ef80_15);
and \U$27740 ( \28083 , \28082 , \20747 );
nor \U$27741 ( \28084 , \28081 , \28083 );
nand \U$27742 ( \28085 , \28084 , \1444 );
nand \U$27743 ( \28086 , \28080 , \28085 );
not \U$27744 ( \28087 , \1441 );
not \U$27745 ( \28088 , \816 );
or \U$27746 ( \28089 , \28087 , \28088 );
nand \U$27747 ( \28090 , \28089 , \17506 );
and \U$27748 ( \28091 , RIbb2ef08_16, RIbb2ee90_17);
nor \U$27749 ( \28092 , \28091 , \2356 );
and \U$27750 ( \28093 , \28090 , \28092 );
xor \U$27751 ( \28094 , \28086 , \28093 );
not \U$27752 ( \28095 , \835 );
not \U$27753 ( \28096 , RIbb2ee90_17);
not \U$27754 ( \28097 , \17756 );
or \U$27755 ( \28098 , \28096 , \28097 );
nand \U$27756 ( \28099 , \27237 , \859 );
nand \U$27757 ( \28100 , \28098 , \28099 );
not \U$27758 ( \28101 , \28100 );
or \U$27759 ( \28102 , \28095 , \28101 );
nand \U$27760 ( \28103 , \27809 , \831 );
nand \U$27761 ( \28104 , \28102 , \28103 );
xor \U$27762 ( \28105 , \28094 , \28104 );
not \U$27763 ( \28106 , \854 );
and \U$27764 ( \28107 , \19831 , \843 );
not \U$27765 ( \28108 , \19831 );
and \U$27766 ( \28109 , \28108 , RIbb2eda0_19);
or \U$27767 ( \28110 , \28107 , \28109 );
not \U$27768 ( \28111 , \28110 );
or \U$27769 ( \28112 , \28106 , \28111 );
nand \U$27770 ( \28113 , \27822 , \853 );
nand \U$27771 ( \28114 , \28112 , \28113 );
xor \U$27772 ( \28115 , \28105 , \28114 );
not \U$27773 ( \28116 , \8362 );
not \U$27774 ( \28117 , \25849 );
or \U$27775 ( \28118 , \28116 , \28117 );
and \U$27776 ( \28119 , RIbb2e350_41, \15797 );
not \U$27777 ( \28120 , RIbb2e350_41);
and \U$27778 ( \28121 , \28120 , \6604 );
nor \U$27779 ( \28122 , \28119 , \28121 );
not \U$27780 ( \28123 , \28122 );
nand \U$27781 ( \28124 , \28123 , \8354 );
nand \U$27782 ( \28125 , \28118 , \28124 );
xor \U$27783 ( \28126 , \28115 , \28125 );
not \U$27784 ( \28127 , \3887 );
not \U$27785 ( \28128 , \27791 );
or \U$27786 ( \28129 , \28127 , \28128 );
not \U$27787 ( \28130 , RIbb2e710_33);
not \U$27788 ( \28131 , \14563 );
or \U$27789 ( \28132 , \28130 , \28131 );
nand \U$27790 ( \28133 , \10764 , \7390 );
nand \U$27791 ( \28134 , \28132 , \28133 );
nand \U$27792 ( \28135 , \28134 , \4075 );
nand \U$27793 ( \28136 , \28129 , \28135 );
xor \U$27794 ( \28137 , \28126 , \28136 );
xor \U$27795 ( \28138 , \28073 , \28137 );
or \U$27796 ( \28139 , \26846 , \26857 );
nand \U$27797 ( \28140 , \28139 , \26836 );
nand \U$27798 ( \28141 , \26846 , \26857 );
nand \U$27799 ( \28142 , \28140 , \28141 );
xor \U$27800 ( \28143 , \28138 , \28142 );
xnor \U$27801 ( \28144 , \28048 , \28143 );
xnor \U$27802 ( \28145 , \28044 , \28144 );
xor \U$27803 ( \28146 , \26859 , \26995 );
and \U$27804 ( \28147 , \28146 , \27109 );
and \U$27805 ( \28148 , \26859 , \26995 );
or \U$27806 ( \28149 , \28147 , \28148 );
xor \U$27807 ( \28150 , \28145 , \28149 );
xor \U$27808 ( \28151 , \27760 , \27877 );
and \U$27809 ( \28152 , \28151 , \27902 );
and \U$27810 ( \28153 , \27760 , \27877 );
or \U$27811 ( \28154 , \28152 , \28153 );
xor \U$27812 ( \28155 , \28150 , \28154 );
xor \U$27813 ( \28156 , \27677 , \27903 );
and \U$27814 ( \28157 , \28156 , \27924 );
and \U$27815 ( \28158 , \27677 , \27903 );
or \U$27816 ( \28159 , \28157 , \28158 );
xor \U$27817 ( \28160 , \28155 , \28159 );
xor \U$27818 ( \28161 , \26801 , \26811 );
and \U$27819 ( \28162 , \28161 , \26822 );
and \U$27820 ( \28163 , \26801 , \26811 );
or \U$27821 ( \28164 , \28162 , \28163 );
not \U$27822 ( \28165 , \16271 );
not \U$27823 ( \28166 , \26809 );
or \U$27824 ( \28167 , \28165 , \28166 );
not \U$27825 ( \28168 , \14725 );
xor \U$27826 ( \28169 , RIbb2dae0_59, \28168 );
nand \U$27827 ( \28170 , \28169 , \17470 );
nand \U$27828 ( \28171 , \28167 , \28170 );
not \U$27829 ( \28172 , \16541 );
not \U$27830 ( \28173 , \26833 );
or \U$27831 ( \28174 , \28172 , \28173 );
not \U$27832 ( \28175 , RIbb2d9f0_61);
not \U$27833 ( \28176 , \17386 );
or \U$27834 ( \28177 , \28175 , \28176 );
not \U$27835 ( \28178 , \22684 );
nand \U$27836 ( \28179 , \28178 , \19746 );
nand \U$27837 ( \28180 , \28177 , \28179 );
nand \U$27838 ( \28181 , \28180 , \16533 );
nand \U$27839 ( \28182 , \28174 , \28181 );
xor \U$27840 ( \28183 , \28171 , \28182 );
not \U$27841 ( \28184 , \13467 );
not \U$27842 ( \28185 , \26752 );
or \U$27843 ( \28186 , \28184 , \28185 );
and \U$27844 ( \28187 , \16400 , \12681 );
not \U$27845 ( \28188 , \16400 );
and \U$27846 ( \28189 , \28188 , RIbb2ddb0_53);
or \U$27847 ( \28190 , \28187 , \28189 );
nand \U$27848 ( \28191 , \28190 , \14930 );
nand \U$27849 ( \28192 , \28186 , \28191 );
xor \U$27850 ( \28193 , \28183 , \28192 );
not \U$27851 ( \28194 , \3613 );
not \U$27852 ( \28195 , RIbb2e800_31);
not \U$27853 ( \28196 , \14886 );
or \U$27854 ( \28197 , \28195 , \28196 );
nand \U$27855 ( \28198 , \14885 , \2917 );
nand \U$27856 ( \28199 , \28197 , \28198 );
not \U$27857 ( \28200 , \28199 );
or \U$27858 ( \28201 , \28194 , \28200 );
nand \U$27859 ( \28202 , \27780 , \2939 );
nand \U$27860 ( \28203 , \28201 , \28202 );
not \U$27861 ( \28204 , \10119 );
not \U$27862 ( \28205 , RIbb2e170_45);
not \U$27863 ( \28206 , \13560 );
or \U$27864 ( \28207 , \28205 , \28206 );
nand \U$27865 ( \28208 , \8375 , \12003 );
nand \U$27866 ( \28209 , \28207 , \28208 );
not \U$27867 ( \28210 , \28209 );
or \U$27868 ( \28211 , \28204 , \28210 );
nand \U$27869 ( \28212 , \25866 , \10599 );
nand \U$27870 ( \28213 , \28211 , \28212 );
xor \U$27871 ( \28214 , \28203 , \28213 );
not \U$27872 ( \28215 , \9099 );
not \U$27873 ( \28216 , RIbb2e260_43);
not \U$27874 ( \28217 , \17341 );
or \U$27875 ( \28218 , \28216 , \28217 );
nand \U$27876 ( \28219 , \7111 , \8347 );
nand \U$27877 ( \28220 , \28218 , \28219 );
not \U$27878 ( \28221 , \28220 );
or \U$27879 ( \28222 , \28215 , \28221 );
nand \U$27880 ( \28223 , \25888 , \9098 );
nand \U$27881 ( \28224 , \28222 , \28223 );
xor \U$27882 ( \28225 , \28214 , \28224 );
and \U$27883 ( \28226 , \28193 , \28225 );
not \U$27884 ( \28227 , \28193 );
not \U$27885 ( \28228 , \28225 );
and \U$27886 ( \28229 , \28227 , \28228 );
nor \U$27887 ( \28230 , \28226 , \28229 );
xor \U$27888 ( \28231 , \28164 , \28230 );
xor \U$27889 ( \28232 , \27681 , \27686 );
and \U$27890 ( \28233 , \28232 , \27759 );
and \U$27891 ( \28234 , \27681 , \27686 );
or \U$27892 ( \28235 , \28233 , \28234 );
xor \U$27893 ( \28236 , \28231 , \28235 );
xor \U$27894 ( \28237 , \25663 , \25718 );
and \U$27895 ( \28238 , \28237 , \25769 );
and \U$27896 ( \28239 , \25663 , \25718 );
or \U$27897 ( \28240 , \28238 , \28239 );
not \U$27898 ( \28241 , \28240 );
xor \U$27899 ( \28242 , \27846 , \27850 );
and \U$27900 ( \28243 , \28242 , \27855 );
and \U$27901 ( \28244 , \27846 , \27850 );
or \U$27902 ( \28245 , \28243 , \28244 );
not \U$27903 ( \28246 , \28245 );
xor \U$27904 ( \28247 , \27764 , \27796 );
and \U$27905 ( \28248 , \28247 , \27801 );
and \U$27906 ( \28249 , \27764 , \27796 );
or \U$27907 ( \28250 , \28248 , \28249 );
not \U$27908 ( \28251 , \28250 );
not \U$27909 ( \28252 , \28251 );
and \U$27910 ( \28253 , \28246 , \28252 );
and \U$27911 ( \28254 , \28245 , \28251 );
nor \U$27912 ( \28255 , \28253 , \28254 );
not \U$27913 ( \28256 , \28255 );
or \U$27914 ( \28257 , \28241 , \28256 );
or \U$27915 ( \28258 , \28255 , \28240 );
nand \U$27916 ( \28259 , \28257 , \28258 );
xor \U$27917 ( \28260 , \28236 , \28259 );
not \U$27918 ( \28261 , \25956 );
not \U$27919 ( \28262 , \25770 );
or \U$27920 ( \28263 , \28261 , \28262 );
or \U$27921 ( \28264 , \25770 , \25956 );
nand \U$27922 ( \28265 , \28264 , \26105 );
nand \U$27923 ( \28266 , \28263 , \28265 );
xor \U$27924 ( \28267 , \27802 , \27856 );
and \U$27925 ( \28268 , \28267 , \27876 );
and \U$27926 ( \28269 , \27802 , \27856 );
or \U$27927 ( \28270 , \28268 , \28269 );
xor \U$27928 ( \28271 , \28266 , \28270 );
not \U$27929 ( \28272 , \2980 );
not \U$27930 ( \28273 , \27841 );
or \U$27931 ( \28274 , \28272 , \28273 );
and \U$27932 ( \28275 , RIbb2ead0_25, \14503 );
not \U$27933 ( \28276 , RIbb2ead0_25);
and \U$27934 ( \28277 , \28276 , \16320 );
or \U$27935 ( \28278 , \28275 , \28277 );
nand \U$27936 ( \28279 , \28278 , \2963 );
nand \U$27937 ( \28280 , \28274 , \28279 );
not \U$27938 ( \28281 , \3382 );
not \U$27939 ( \28282 , RIbb2ebc0_23);
not \U$27940 ( \28283 , \17681 );
or \U$27941 ( \28284 , \28282 , \28283 );
nand \U$27942 ( \28285 , \16782 , \3388 );
nand \U$27943 ( \28286 , \28284 , \28285 );
not \U$27944 ( \28287 , \28286 );
or \U$27945 ( \28288 , \28281 , \28287 );
nand \U$27946 ( \28289 , \26728 , \3406 );
nand \U$27947 ( \28290 , \28288 , \28289 );
not \U$27948 ( \28291 , \3465 );
not \U$27949 ( \28292 , RIbb2e9e0_27);
not \U$27950 ( \28293 , \18857 );
or \U$27951 ( \28294 , \28292 , \28293 );
nand \U$27952 ( \28295 , \13210 , \3454 );
nand \U$27953 ( \28296 , \28294 , \28295 );
not \U$27954 ( \28297 , \28296 );
or \U$27955 ( \28298 , \28291 , \28297 );
nand \U$27956 ( \28299 , \27833 , \3445 );
nand \U$27957 ( \28300 , \28298 , \28299 );
xor \U$27958 ( \28301 , \28290 , \28300 );
xor \U$27959 ( \28302 , \28280 , \28301 );
xor \U$27960 ( \28303 , \25875 , \25890 );
and \U$27961 ( \28304 , \28303 , \25906 );
and \U$27962 ( \28305 , \25875 , \25890 );
or \U$27963 ( \28306 , \28304 , \28305 );
xor \U$27964 ( \28307 , \28302 , \28306 );
buf \U$27965 ( \28308 , \25840 );
or \U$27966 ( \28309 , \28308 , \25858 );
nand \U$27967 ( \28310 , \28309 , \25827 );
nand \U$27968 ( \28311 , \25858 , \28308 );
nand \U$27969 ( \28312 , \28310 , \28311 );
xor \U$27970 ( \28313 , \28307 , \28312 );
not \U$27971 ( \28314 , \25907 );
not \U$27972 ( \28315 , \25952 );
or \U$27973 ( \28316 , \28314 , \28315 );
not \U$27974 ( \28317 , \25907 );
not \U$27975 ( \28318 , \28317 );
not \U$27976 ( \28319 , \25951 );
or \U$27977 ( \28320 , \28318 , \28319 );
not \U$27978 ( \28321 , \25859 );
nand \U$27979 ( \28322 , \28320 , \28321 );
nand \U$27980 ( \28323 , \28316 , \28322 );
not \U$27981 ( \28324 , \28323 );
xor \U$27982 ( \28325 , \28313 , \28324 );
xor \U$27983 ( \28326 , \27774 , \27784 );
and \U$27984 ( \28327 , \28326 , \27795 );
and \U$27985 ( \28328 , \27774 , \27784 );
or \U$27986 ( \28329 , \28327 , \28328 );
not \U$27987 ( \28330 , \25938 );
not \U$27988 ( \28331 , \28330 );
not \U$27989 ( \28332 , \25921 );
or \U$27990 ( \28333 , \28331 , \28332 );
not \U$27991 ( \28334 , \25938 );
not \U$27992 ( \28335 , \25921 );
not \U$27993 ( \28336 , \28335 );
or \U$27994 ( \28337 , \28334 , \28336 );
nand \U$27995 ( \28338 , \28337 , \25950 );
nand \U$27996 ( \28339 , \28333 , \28338 );
buf \U$27997 ( \28340 , \28339 );
xor \U$27998 ( \28341 , \28329 , \28340 );
xor \U$27999 ( \28342 , \26733 , \26743 );
and \U$28000 ( \28343 , \28342 , \26756 );
and \U$28001 ( \28344 , \26733 , \26743 );
or \U$28002 ( \28345 , \28343 , \28344 );
xnor \U$28003 ( \28346 , \28341 , \28345 );
xnor \U$28004 ( \28347 , \28325 , \28346 );
not \U$28005 ( \28348 , \28347 );
buf \U$28006 ( \28349 , \28348 );
xor \U$28007 ( \28350 , \28271 , \28349 );
xor \U$28008 ( \28351 , \28260 , \28350 );
xor \U$28009 ( \28352 , \26110 , \26704 );
and \U$28010 ( \28353 , \28352 , \27110 );
and \U$28011 ( \28354 , \26110 , \26704 );
or \U$28012 ( \28355 , \28353 , \28354 );
xor \U$28013 ( \28356 , \28351 , \28355 );
xor \U$28014 ( \28357 , \28160 , \28356 );
not \U$28015 ( \28358 , \28357 );
or \U$28016 ( \28359 , \27929 , \28358 );
xor \U$28017 ( \28360 , \27111 , \27671 );
xor \U$28018 ( \28361 , \28360 , \27925 );
xor \U$28019 ( \28362 , \27912 , \27918 );
xor \U$28020 ( \28363 , \28362 , \27921 );
not \U$28021 ( \28364 , \28363 );
not \U$28022 ( \28365 , \27355 );
not \U$28023 ( \28366 , \27665 );
and \U$28024 ( \28367 , \28365 , \28366 );
and \U$28025 ( \28368 , \27355 , \27665 );
nor \U$28026 ( \28369 , \28367 , \28368 );
xor \U$28027 ( \28370 , \28369 , \27342 );
nand \U$28028 ( \28371 , \28364 , \28370 );
not \U$28029 ( \28372 , \28371 );
xnor \U$28030 ( \28373 , \27206 , \27258 );
xnor \U$28031 ( \28374 , \27172 , \28373 );
xor \U$28032 ( \28375 , \27182 , \27192 );
xor \U$28033 ( \28376 , \28375 , \27203 );
not \U$28034 ( \28377 , \2939 );
not \U$28035 ( \28378 , RIbb2e800_31);
not \U$28036 ( \28379 , \17681 );
or \U$28037 ( \28380 , \28378 , \28379 );
nand \U$28038 ( \28381 , \17682 , \2917 );
nand \U$28039 ( \28382 , \28380 , \28381 );
not \U$28040 ( \28383 , \28382 );
or \U$28041 ( \28384 , \28377 , \28383 );
nand \U$28042 ( \28385 , \27180 , \2941 );
nand \U$28043 ( \28386 , \28384 , \28385 );
not \U$28044 ( \28387 , \28386 );
not \U$28045 ( \28388 , \4714 );
not \U$28046 ( \28389 , \27201 );
or \U$28047 ( \28390 , \28388 , \28389 );
buf \U$28048 ( \28391 , \13210 );
and \U$28049 ( \28392 , RIbb2e620_35, \28391 );
not \U$28050 ( \28393 , RIbb2e620_35);
and \U$28051 ( \28394 , \28393 , \13211 );
nor \U$28052 ( \28395 , \28392 , \28394 );
nand \U$28053 ( \28396 , \28395 , \4712 );
nand \U$28054 ( \28397 , \28390 , \28396 );
not \U$28055 ( \28398 , \28397 );
nand \U$28056 ( \28399 , \28387 , \28398 );
not \U$28057 ( \28400 , \28399 );
not \U$28058 ( \28401 , \14752 );
not \U$28059 ( \28402 , \27523 );
or \U$28060 ( \28403 , \28401 , \28402 );
not \U$28061 ( \28404 , RIbb2df90_49);
not \U$28062 ( \28405 , \13876 );
or \U$28063 ( \28406 , \28404 , \28405 );
nand \U$28064 ( \28407 , \6604 , \12278 );
nand \U$28065 ( \28408 , \28406 , \28407 );
nand \U$28066 ( \28409 , \28408 , \12167 );
nand \U$28067 ( \28410 , \28403 , \28409 );
not \U$28068 ( \28411 , \28410 );
or \U$28069 ( \28412 , \28400 , \28411 );
not \U$28070 ( \28413 , \28398 );
nand \U$28071 ( \28414 , \28413 , \28386 );
nand \U$28072 ( \28415 , \28412 , \28414 );
xor \U$28073 ( \28416 , \28376 , \28415 );
xor \U$28074 ( \28417 , \27563 , \27571 );
not \U$28075 ( \28418 , \2963 );
not \U$28076 ( \28419 , \27239 );
or \U$28077 ( \28420 , \28418 , \28419 );
and \U$28078 ( \28421 , RIbb2ead0_25, \16819 );
not \U$28079 ( \28422 , RIbb2ead0_25);
and \U$28080 ( \28423 , \28422 , \16818 );
or \U$28081 ( \28424 , \28421 , \28423 );
nand \U$28082 ( \28425 , \28424 , \2979 );
nand \U$28083 ( \28426 , \28420 , \28425 );
xor \U$28084 ( \28427 , \28417 , \28426 );
not \U$28085 ( \28428 , \3465 );
not \U$28086 ( \28429 , \27581 );
or \U$28087 ( \28430 , \28428 , \28429 );
not \U$28088 ( \28431 , RIbb2e9e0_27);
not \U$28089 ( \28432 , \16554 );
or \U$28090 ( \28433 , \28431 , \28432 );
nand \U$28091 ( \28434 , \16706 , \3462 );
nand \U$28092 ( \28435 , \28433 , \28434 );
nand \U$28093 ( \28436 , \28435 , \3445 );
nand \U$28094 ( \28437 , \28430 , \28436 );
and \U$28095 ( \28438 , \28427 , \28437 );
and \U$28096 ( \28439 , \28417 , \28426 );
or \U$28097 ( \28440 , \28438 , \28439 );
not \U$28098 ( \28441 , RIbb2e350_41);
not \U$28099 ( \28442 , \14563 );
or \U$28100 ( \28443 , \28441 , \28442 );
nand \U$28101 ( \28444 , \13526 , \7097 );
nand \U$28102 ( \28445 , \28443 , \28444 );
not \U$28103 ( \28446 , \28445 );
or \U$28104 ( \28447 , \28446 , \8363 );
or \U$28105 ( \28448 , \27604 , \8352 );
nand \U$28106 ( \28449 , \28447 , \28448 );
xor \U$28107 ( \28450 , \28440 , \28449 );
and \U$28108 ( \28451 , \8450 , \27615 );
and \U$28109 ( \28452 , RIbb2e440_39, \11580 );
not \U$28110 ( \28453 , RIbb2e440_39);
and \U$28111 ( \28454 , \28453 , \14885 );
or \U$28112 ( \28455 , \28452 , \28454 );
and \U$28113 ( \28456 , \28455 , \7103 );
nor \U$28114 ( \28457 , \28451 , \28456 );
not \U$28115 ( \28458 , \28457 );
and \U$28116 ( \28459 , \28450 , \28458 );
and \U$28117 ( \28460 , \28440 , \28449 );
or \U$28118 ( \28461 , \28459 , \28460 );
and \U$28119 ( \28462 , \28416 , \28461 );
and \U$28120 ( \28463 , \28376 , \28415 );
or \U$28121 ( \28464 , \28462 , \28463 );
or \U$28122 ( \28465 , \28374 , \28464 );
xor \U$28123 ( \28466 , \27544 , \27551 );
xor \U$28124 ( \28467 , \28466 , \27547 );
nand \U$28125 ( \28468 , \28465 , \28467 );
not \U$28126 ( \28469 , \27172 );
not \U$28127 ( \28470 , \28373 );
and \U$28128 ( \28471 , \28469 , \28470 );
and \U$28129 ( \28472 , \27172 , \28373 );
nor \U$28130 ( \28473 , \28471 , \28472 );
not \U$28131 ( \28474 , \28473 );
nand \U$28132 ( \28475 , \28474 , \28464 );
nand \U$28133 ( \28476 , \28468 , \28475 );
xor \U$28134 ( \28477 , \27553 , \27555 );
xor \U$28135 ( \28478 , \28477 , \27658 );
xor \U$28136 ( \28479 , \28476 , \28478 );
xor \U$28137 ( \28480 , \27358 , \27415 );
xor \U$28138 ( \28481 , \28480 , \27475 );
and \U$28139 ( \28482 , \28479 , \28481 );
and \U$28140 ( \28483 , \28476 , \28478 );
or \U$28141 ( \28484 , \28482 , \28483 );
not \U$28142 ( \28485 , \28484 );
not \U$28143 ( \28486 , \28485 );
xnor \U$28144 ( \28487 , \27661 , \27488 );
not \U$28145 ( \28488 , \27478 );
and \U$28146 ( \28489 , \28487 , \28488 );
not \U$28147 ( \28490 , \28487 );
and \U$28148 ( \28491 , \28490 , \27478 );
nor \U$28149 ( \28492 , \28489 , \28491 );
not \U$28150 ( \28493 , \28492 );
or \U$28151 ( \28494 , \28486 , \28493 );
not \U$28152 ( \28495 , \9098 );
not \U$28153 ( \28496 , RIbb2e260_43);
not \U$28154 ( \28497 , \20044 );
or \U$28155 ( \28498 , \28496 , \28497 );
nand \U$28156 ( \28499 , \9840 , \26255 );
nand \U$28157 ( \28500 , \28498 , \28499 );
not \U$28158 ( \28501 , \28500 );
or \U$28159 ( \28502 , \28495 , \28501 );
nand \U$28160 ( \28503 , \27167 , \9099 );
nand \U$28161 ( \28504 , \28502 , \28503 );
not \U$28162 ( \28505 , \28504 );
not \U$28163 ( \28506 , \28505 );
not \U$28164 ( \28507 , \11176 );
not \U$28165 ( \28508 , RIbb2e080_47);
not \U$28166 ( \28509 , \13850 );
or \U$28167 ( \28510 , \28508 , \28509 );
nand \U$28168 ( \28511 , \7296 , \10113 );
nand \U$28169 ( \28512 , \28510 , \28511 );
not \U$28170 ( \28513 , \28512 );
or \U$28171 ( \28514 , \28507 , \28513 );
nand \U$28172 ( \28515 , \27498 , \11177 );
nand \U$28173 ( \28516 , \28514 , \28515 );
not \U$28174 ( \28517 , \28516 );
not \U$28175 ( \28518 , \28517 );
or \U$28176 ( \28519 , \28506 , \28518 );
not \U$28177 ( \28520 , \10599 );
and \U$28178 ( \28521 , \23529 , RIbb2e170_45);
not \U$28179 ( \28522 , \23529 );
and \U$28180 ( \28523 , \28522 , \9094 );
or \U$28181 ( \28524 , \28521 , \28523 );
not \U$28182 ( \28525 , \28524 );
or \U$28183 ( \28526 , \28520 , \28525 );
nand \U$28184 ( \28527 , \27511 , \10119 );
nand \U$28185 ( \28528 , \28526 , \28527 );
nand \U$28186 ( \28529 , \28519 , \28528 );
not \U$28187 ( \28530 , \28505 );
nand \U$28188 ( \28531 , \28530 , \28516 );
nand \U$28189 ( \28532 , \28529 , \28531 );
xor \U$28190 ( \28533 , \27148 , \27157 );
xor \U$28191 ( \28534 , \28533 , \27169 );
xor \U$28192 ( \28535 , \28532 , \28534 );
xor \U$28193 ( \28536 , \27502 , \27513 );
xor \U$28194 ( \28537 , \28536 , \27525 );
and \U$28195 ( \28538 , \28535 , \28537 );
and \U$28196 ( \28539 , \28532 , \28534 );
or \U$28197 ( \28540 , \28538 , \28539 );
xor \U$28198 ( \28541 , \27597 , \27607 );
xor \U$28199 ( \28542 , \28541 , \27619 );
not \U$28200 ( \28543 , \12692 );
not \U$28201 ( \28544 , \27155 );
or \U$28202 ( \28545 , \28543 , \28544 );
and \U$28203 ( \28546 , RIbb2dea0_51, \9108 );
not \U$28204 ( \28547 , RIbb2dea0_51);
and \U$28205 ( \28548 , \28547 , \8387 );
or \U$28206 ( \28549 , \28546 , \28548 );
nand \U$28207 ( \28550 , \28549 , \12774 );
nand \U$28208 ( \28551 , \28545 , \28550 );
not \U$28209 ( \28552 , \28551 );
not \U$28210 ( \28553 , \28552 );
not \U$28211 ( \28554 , \15746 );
and \U$28212 ( \28555 , RIbb2dbd0_57, \16185 );
not \U$28213 ( \28556 , RIbb2dbd0_57);
and \U$28214 ( \28557 , \28556 , \17910 );
nor \U$28215 ( \28558 , \28555 , \28557 );
not \U$28216 ( \28559 , \28558 );
or \U$28217 ( \28560 , \28554 , \28559 );
nand \U$28218 ( \28561 , \27397 , \17397 );
nand \U$28219 ( \28562 , \28560 , \28561 );
not \U$28220 ( \28563 , \28562 );
not \U$28221 ( \28564 , \28563 );
or \U$28222 ( \28565 , \28553 , \28564 );
not \U$28223 ( \28566 , \14930 );
not \U$28224 ( \28567 , \27631 );
or \U$28225 ( \28568 , \28566 , \28567 );
not \U$28226 ( \28569 , RIbb2ddb0_53);
not \U$28227 ( \28570 , \4392 );
or \U$28228 ( \28571 , \28569 , \28570 );
nand \U$28229 ( \28572 , \8375 , \26750 );
nand \U$28230 ( \28573 , \28571 , \28572 );
nand \U$28231 ( \28574 , \28573 , \14920 );
nand \U$28232 ( \28575 , \28568 , \28574 );
nand \U$28233 ( \28576 , \28565 , \28575 );
not \U$28234 ( \28577 , \28552 );
nand \U$28235 ( \28578 , \28577 , \28562 );
nand \U$28236 ( \28579 , \28576 , \28578 );
xor \U$28237 ( \28580 , \28542 , \28579 );
xor \U$28238 ( \28581 , \27572 , \27583 );
xor \U$28239 ( \28582 , \28581 , \27594 );
not \U$28240 ( \28583 , \14613 );
and \U$28241 ( \28584 , RIbb2dcc0_55, \12577 );
not \U$28242 ( \28585 , RIbb2dcc0_55);
and \U$28243 ( \28586 , \28585 , \10458 );
or \U$28244 ( \28587 , \28584 , \28586 );
not \U$28245 ( \28588 , \28587 );
or \U$28246 ( \28589 , \28583 , \28588 );
nand \U$28247 ( \28590 , \27638 , \15181 );
nand \U$28248 ( \28591 , \28589 , \28590 );
xor \U$28249 ( \28592 , \28582 , \28591 );
not \U$28250 ( \28593 , \16541 );
not \U$28251 ( \28594 , RIbb2d9f0_61);
not \U$28252 ( \28595 , \4639 );
or \U$28253 ( \28596 , \28594 , \28595 );
nand \U$28254 ( \28597 , \4640 , \16537 );
nand \U$28255 ( \28598 , \28596 , \28597 );
not \U$28256 ( \28599 , \28598 );
or \U$28257 ( \28600 , \28593 , \28599 );
nand \U$28258 ( \28601 , \27406 , \26834 );
nand \U$28259 ( \28602 , \28600 , \28601 );
and \U$28260 ( \28603 , \28592 , \28602 );
and \U$28261 ( \28604 , \28582 , \28591 );
or \U$28262 ( \28605 , \28603 , \28604 );
and \U$28263 ( \28606 , \28580 , \28605 );
and \U$28264 ( \28607 , \28542 , \28579 );
or \U$28265 ( \28608 , \28606 , \28607 );
xor \U$28266 ( \28609 , \28540 , \28608 );
xor \U$28267 ( \28610 , \27390 , \27399 );
xor \U$28268 ( \28611 , \28610 , \27410 );
xor \U$28269 ( \28612 , \27633 , \27642 );
xor \U$28270 ( \28613 , \28612 , \27652 );
xor \U$28271 ( \28614 , \28611 , \28613 );
and \U$28272 ( \28615 , \17506 , \3381 );
not \U$28273 ( \28616 , \2962 );
not \U$28274 ( \28617 , \28424 );
or \U$28275 ( \28618 , \28616 , \28617 );
and \U$28276 ( \28619 , RIbb2ead0_25, \17745 );
not \U$28277 ( \28620 , RIbb2ead0_25);
not \U$28278 ( \28621 , \17745 );
and \U$28279 ( \28622 , \28620 , \28621 );
or \U$28280 ( \28623 , \28619 , \28622 );
nand \U$28281 ( \28624 , \28623 , \2979 );
nand \U$28282 ( \28625 , \28618 , \28624 );
xor \U$28283 ( \28626 , \28615 , \28625 );
not \U$28284 ( \28627 , \3444 );
not \U$28285 ( \28628 , RIbb2e9e0_27);
not \U$28286 ( \28629 , \18924 );
or \U$28287 ( \28630 , \28628 , \28629 );
nand \U$28288 ( \28631 , \18923 , \3454 );
nand \U$28289 ( \28632 , \28630 , \28631 );
not \U$28290 ( \28633 , \28632 );
or \U$28291 ( \28634 , \28627 , \28633 );
nand \U$28292 ( \28635 , \28435 , \3465 );
nand \U$28293 ( \28636 , \28634 , \28635 );
and \U$28294 ( \28637 , \28626 , \28636 );
and \U$28295 ( \28638 , \28615 , \28625 );
or \U$28296 ( \28639 , \28637 , \28638 );
not \U$28297 ( \28640 , \2922 );
not \U$28298 ( \28641 , RIbb2e8f0_29);
not \U$28299 ( \28642 , \16751 );
not \U$28300 ( \28643 , \28642 );
or \U$28301 ( \28644 , \28641 , \28643 );
not \U$28302 ( \28645 , \16747 );
nand \U$28303 ( \28646 , \28645 , \2949 );
nand \U$28304 ( \28647 , \28644 , \28646 );
not \U$28305 ( \28648 , \28647 );
or \U$28306 ( \28649 , \28640 , \28648 );
nand \U$28307 ( \28650 , \27592 , \2925 );
nand \U$28308 ( \28651 , \28649 , \28650 );
xor \U$28309 ( \28652 , \28639 , \28651 );
not \U$28310 ( \28653 , \6250 );
not \U$28311 ( \28654 , RIbb2e530_37);
not \U$28312 ( \28655 , \13809 );
or \U$28313 ( \28656 , \28654 , \28655 );
nand \U$28314 ( \28657 , \16765 , \8701 );
nand \U$28315 ( \28658 , \28656 , \28657 );
not \U$28316 ( \28659 , \28658 );
or \U$28317 ( \28660 , \28653 , \28659 );
nand \U$28318 ( \28661 , \27465 , \20792 );
nand \U$28319 ( \28662 , \28660 , \28661 );
and \U$28320 ( \28663 , \28652 , \28662 );
and \U$28321 ( \28664 , \28639 , \28651 );
or \U$28322 ( \28665 , \28663 , \28664 );
not \U$28323 ( \28666 , \17275 );
not \U$28324 ( \28667 , RIbb2d900_63);
not \U$28325 ( \28668 , \3168 );
or \U$28326 ( \28669 , \28667 , \28668 );
not \U$28327 ( \28670 , \6107 );
nand \U$28328 ( \28671 , \28670 , \17262 );
nand \U$28329 ( \28672 , \28669 , \28671 );
not \U$28330 ( \28673 , \28672 );
or \U$28331 ( \28674 , \28666 , \28673 );
nand \U$28332 ( \28675 , \27648 , RIbb2d888_64);
nand \U$28333 ( \28676 , \28674 , \28675 );
xor \U$28334 ( \28677 , \28665 , \28676 );
not \U$28335 ( \28678 , \16271 );
and \U$28336 ( \28679 , RIbb2dae0_59, \12707 );
not \U$28337 ( \28680 , RIbb2dae0_59);
and \U$28338 ( \28681 , \28680 , \7021 );
or \U$28339 ( \28682 , \28679 , \28681 );
not \U$28340 ( \28683 , \28682 );
or \U$28341 ( \28684 , \28678 , \28683 );
nand \U$28342 ( \28685 , \27439 , \16257 );
nand \U$28343 ( \28686 , \28684 , \28685 );
and \U$28344 ( \28687 , \28677 , \28686 );
and \U$28345 ( \28688 , \28665 , \28676 );
or \U$28346 ( \28689 , \28687 , \28688 );
and \U$28347 ( \28690 , \28614 , \28689 );
and \U$28348 ( \28691 , \28611 , \28613 );
or \U$28349 ( \28692 , \28690 , \28691 );
and \U$28350 ( \28693 , \28609 , \28692 );
and \U$28351 ( \28694 , \28540 , \28608 );
or \U$28352 ( \28695 , \28693 , \28694 );
not \U$28353 ( \28696 , \28695 );
xor \U$28354 ( \28697 , \27558 , \27622 );
xor \U$28355 ( \28698 , \28697 , \27655 );
not \U$28356 ( \28699 , \27413 );
not \U$28357 ( \28700 , \28699 );
not \U$28358 ( \28701 , \27377 );
not \U$28359 ( \28702 , \27368 );
or \U$28360 ( \28703 , \28701 , \28702 );
or \U$28361 ( \28704 , \27377 , \27368 );
nand \U$28362 ( \28705 , \28703 , \28704 );
not \U$28363 ( \28706 , \28705 );
or \U$28364 ( \28707 , \28700 , \28706 );
or \U$28365 ( \28708 , \28699 , \28705 );
nand \U$28366 ( \28709 , \28707 , \28708 );
xor \U$28367 ( \28710 , \28698 , \28709 );
xor \U$28368 ( \28711 , \28417 , \28426 );
xor \U$28369 ( \28712 , \28711 , \28437 );
not \U$28370 ( \28713 , \11176 );
not \U$28371 ( \28714 , RIbb2e080_47);
not \U$28372 ( \28715 , \8319 );
or \U$28373 ( \28716 , \28714 , \28715 );
nand \U$28374 ( \28717 , \9818 , \16171 );
nand \U$28375 ( \28718 , \28716 , \28717 );
not \U$28376 ( \28719 , \28718 );
or \U$28377 ( \28720 , \28713 , \28719 );
nand \U$28378 ( \28721 , \28512 , \12965 );
nand \U$28379 ( \28722 , \28720 , \28721 );
xor \U$28380 ( \28723 , \28712 , \28722 );
not \U$28381 ( \28724 , \13295 );
not \U$28382 ( \28725 , RIbb2df90_49);
not \U$28383 ( \28726 , \11535 );
or \U$28384 ( \28727 , \28725 , \28726 );
not \U$28385 ( \28728 , \9791 );
nand \U$28386 ( \28729 , \28728 , \12278 );
nand \U$28387 ( \28730 , \28727 , \28729 );
not \U$28388 ( \28731 , \28730 );
or \U$28389 ( \28732 , \28724 , \28731 );
nand \U$28390 ( \28733 , \28408 , \16427 );
nand \U$28391 ( \28734 , \28732 , \28733 );
and \U$28392 ( \28735 , \28723 , \28734 );
and \U$28393 ( \28736 , \28712 , \28722 );
or \U$28394 ( \28737 , \28735 , \28736 );
not \U$28395 ( \28738 , \28737 );
not \U$28396 ( \28739 , \2941 );
not \U$28397 ( \28740 , \28382 );
or \U$28398 ( \28741 , \28739 , \28740 );
not \U$28399 ( \28742 , RIbb2e800_31);
not \U$28400 ( \28743 , \16563 );
or \U$28401 ( \28744 , \28742 , \28743 );
nand \U$28402 ( \28745 , \15753 , \8810 );
nand \U$28403 ( \28746 , \28744 , \28745 );
nand \U$28404 ( \28747 , \2939 , \28746 );
nand \U$28405 ( \28748 , \28741 , \28747 );
not \U$28406 ( \28749 , \3886 );
not \U$28407 ( \28750 , RIbb2e710_33);
not \U$28408 ( \28751 , \18353 );
or \U$28409 ( \28752 , \28750 , \28751 );
nand \U$28410 ( \28753 , \20580 , \2935 );
nand \U$28411 ( \28754 , \28752 , \28753 );
not \U$28412 ( \28755 , \28754 );
or \U$28413 ( \28756 , \28749 , \28755 );
nand \U$28414 ( \28757 , \27453 , \4075 );
nand \U$28415 ( \28758 , \28756 , \28757 );
xor \U$28416 ( \28759 , \28748 , \28758 );
not \U$28417 ( \28760 , \4712 );
not \U$28418 ( \28761 , RIbb2e620_35);
not \U$28419 ( \28762 , \15054 );
or \U$28420 ( \28763 , \28761 , \28762 );
nand \U$28421 ( \28764 , \15055 , \6688 );
nand \U$28422 ( \28765 , \28763 , \28764 );
not \U$28423 ( \28766 , \28765 );
or \U$28424 ( \28767 , \28760 , \28766 );
nand \U$28425 ( \28768 , \28395 , \4714 );
nand \U$28426 ( \28769 , \28767 , \28768 );
and \U$28427 ( \28770 , \28759 , \28769 );
and \U$28428 ( \28771 , \28748 , \28758 );
or \U$28429 ( \28772 , \28770 , \28771 );
not \U$28430 ( \28773 , \28772 );
and \U$28431 ( \28774 , \28386 , \28398 );
not \U$28432 ( \28775 , \28386 );
and \U$28433 ( \28776 , \28775 , \28397 );
nor \U$28434 ( \28777 , \28774 , \28776 );
not \U$28435 ( \28778 , \28777 );
not \U$28436 ( \28779 , \28410 );
and \U$28437 ( \28780 , \28778 , \28779 );
and \U$28438 ( \28781 , \28410 , \28777 );
nor \U$28439 ( \28782 , \28780 , \28781 );
nand \U$28440 ( \28783 , \28773 , \28782 );
not \U$28441 ( \28784 , \28783 );
or \U$28442 ( \28785 , \28738 , \28784 );
not \U$28443 ( \28786 , \28782 );
nand \U$28444 ( \28787 , \28786 , \28772 );
nand \U$28445 ( \28788 , \28785 , \28787 );
xor \U$28446 ( \28789 , \27433 , \27443 );
xor \U$28447 ( \28790 , \28789 , \27470 );
nor \U$28448 ( \28791 , \28788 , \28790 );
not \U$28449 ( \28792 , \9098 );
not \U$28450 ( \28793 , RIbb2e260_43);
not \U$28451 ( \28794 , \12234 );
or \U$28452 ( \28795 , \28793 , \28794 );
nand \U$28453 ( \28796 , \10300 , \17231 );
nand \U$28454 ( \28797 , \28795 , \28796 );
not \U$28455 ( \28798 , \28797 );
or \U$28456 ( \28799 , \28792 , \28798 );
nand \U$28457 ( \28800 , \28500 , \10451 );
nand \U$28458 ( \28801 , \28799 , \28800 );
not \U$28459 ( \28802 , \28801 );
not \U$28460 ( \28803 , \8362 );
not \U$28461 ( \28804 , RIbb2e350_41);
not \U$28462 ( \28805 , \12260 );
or \U$28463 ( \28806 , \28804 , \28805 );
nand \U$28464 ( \28807 , \12261 , \8357 );
nand \U$28465 ( \28808 , \28806 , \28807 );
not \U$28466 ( \28809 , \28808 );
or \U$28467 ( \28810 , \28803 , \28809 );
nand \U$28468 ( \28811 , \28445 , \8353 );
nand \U$28469 ( \28812 , \28810 , \28811 );
not \U$28470 ( \28813 , \28812 );
or \U$28471 ( \28814 , \28802 , \28813 );
or \U$28472 ( \28815 , \28801 , \28812 );
not \U$28473 ( \28816 , \10599 );
not \U$28474 ( \28817 , RIbb2e170_45);
not \U$28475 ( \28818 , \13916 );
or \U$28476 ( \28819 , \28817 , \28818 );
nand \U$28477 ( \28820 , \16475 , \13372 );
nand \U$28478 ( \28821 , \28819 , \28820 );
not \U$28479 ( \28822 , \28821 );
or \U$28480 ( \28823 , \28816 , \28822 );
nand \U$28481 ( \28824 , \28524 , \10119 );
nand \U$28482 ( \28825 , \28823 , \28824 );
nand \U$28483 ( \28826 , \28815 , \28825 );
nand \U$28484 ( \28827 , \28814 , \28826 );
not \U$28485 ( \28828 , \28827 );
xor \U$28486 ( \28829 , \27446 , \27457 );
xor \U$28487 ( \28830 , \28829 , \27467 );
not \U$28488 ( \28831 , \28830 );
nand \U$28489 ( \28832 , \28828 , \28831 );
or \U$28490 ( \28833 , RIbb2ea58_26, RIbb2e9e0_27);
nand \U$28491 ( \28834 , \28833 , \19064 );
and \U$28492 ( \28835 , RIbb2ea58_26, RIbb2e9e0_27);
nor \U$28493 ( \28836 , \28835 , \18636 );
and \U$28494 ( \28837 , \28834 , \28836 );
not \U$28495 ( \28838 , \2962 );
not \U$28496 ( \28839 , \28623 );
or \U$28497 ( \28840 , \28838 , \28839 );
and \U$28498 ( \28841 , RIbb2ead0_25, \17506 );
not \U$28499 ( \28842 , RIbb2ead0_25);
and \U$28500 ( \28843 , \28842 , \18929 );
nor \U$28501 ( \28844 , \28841 , \28843 );
nand \U$28502 ( \28845 , \28844 , \2979 );
nand \U$28503 ( \28846 , \28840 , \28845 );
and \U$28504 ( \28847 , \28837 , \28846 );
not \U$28505 ( \28848 , \2924 );
not \U$28506 ( \28849 , \28647 );
or \U$28507 ( \28850 , \28848 , \28849 );
not \U$28508 ( \28851 , RIbb2e8f0_29);
not \U$28509 ( \28852 , \23185 );
or \U$28510 ( \28853 , \28851 , \28852 );
nand \U$28511 ( \28854 , \16829 , \3440 );
nand \U$28512 ( \28855 , \28853 , \28854 );
nand \U$28513 ( \28856 , \28855 , \2921 );
nand \U$28514 ( \28857 , \28850 , \28856 );
xor \U$28515 ( \28858 , \28847 , \28857 );
not \U$28516 ( \28859 , \3613 );
not \U$28517 ( \28860 , \28746 );
or \U$28518 ( \28861 , \28859 , \28860 );
not \U$28519 ( \28862 , RIbb2e800_31);
not \U$28520 ( \28863 , \19195 );
or \U$28521 ( \28864 , \28862 , \28863 );
nand \U$28522 ( \28865 , \16576 , \2917 );
nand \U$28523 ( \28866 , \28864 , \28865 );
nand \U$28524 ( \28867 , \28866 , \2939 );
nand \U$28525 ( \28868 , \28861 , \28867 );
and \U$28526 ( \28869 , \28858 , \28868 );
and \U$28527 ( \28870 , \28847 , \28857 );
or \U$28528 ( \28871 , \28869 , \28870 );
not \U$28529 ( \28872 , \7104 );
not \U$28530 ( \28873 , \28455 );
or \U$28531 ( \28874 , \28872 , \28873 );
and \U$28532 ( \28875 , RIbb2e440_39, \22070 );
not \U$28533 ( \28876 , RIbb2e440_39);
and \U$28534 ( \28877 , \28876 , \12175 );
or \U$28535 ( \28878 , \28875 , \28877 );
nand \U$28536 ( \28879 , \28878 , \7103 );
nand \U$28537 ( \28880 , \28874 , \28879 );
xor \U$28538 ( \28881 , \28871 , \28880 );
not \U$28539 ( \28882 , \17562 );
not \U$28540 ( \28883 , RIbb2ddb0_53);
not \U$28541 ( \28884 , \10556 );
or \U$28542 ( \28885 , \28883 , \28884 );
nand \U$28543 ( \28886 , \4699 , \16210 );
nand \U$28544 ( \28887 , \28885 , \28886 );
not \U$28545 ( \28888 , \28887 );
or \U$28546 ( \28889 , \28882 , \28888 );
nand \U$28547 ( \28890 , \28573 , \14930 );
nand \U$28548 ( \28891 , \28889 , \28890 );
and \U$28549 ( \28892 , \28881 , \28891 );
and \U$28550 ( \28893 , \28871 , \28880 );
or \U$28551 ( \28894 , \28892 , \28893 );
nand \U$28552 ( \28895 , \28832 , \28894 );
not \U$28553 ( \28896 , \28831 );
nand \U$28554 ( \28897 , \28827 , \28896 );
nand \U$28555 ( \28898 , \28895 , \28897 );
not \U$28556 ( \28899 , \28898 );
or \U$28557 ( \28900 , \28791 , \28899 );
nand \U$28558 ( \28901 , \28788 , \28790 );
nand \U$28559 ( \28902 , \28900 , \28901 );
and \U$28560 ( \28903 , \28710 , \28902 );
and \U$28561 ( \28904 , \28698 , \28709 );
or \U$28562 ( \28905 , \28903 , \28904 );
not \U$28563 ( \28906 , \28905 );
or \U$28564 ( \28907 , \28696 , \28906 );
or \U$28565 ( \28908 , \28905 , \28695 );
xor \U$28566 ( \28909 , \27331 , \27333 );
xor \U$28567 ( \28910 , \28909 , \27336 );
nand \U$28568 ( \28911 , \28908 , \28910 );
nand \U$28569 ( \28912 , \28907 , \28911 );
nand \U$28570 ( \28913 , \28494 , \28912 );
not \U$28571 ( \28914 , \28485 );
not \U$28572 ( \28915 , \28492 );
nand \U$28573 ( \28916 , \28914 , \28915 );
nand \U$28574 ( \28917 , \28913 , \28916 );
not \U$28575 ( \28918 , \28917 );
or \U$28576 ( \28919 , \28372 , \28918 );
not \U$28577 ( \28920 , \28370 );
nand \U$28578 ( \28921 , \28920 , \28363 );
nand \U$28579 ( \28922 , \28919 , \28921 );
nand \U$28580 ( \28923 , \28361 , \28922 );
nand \U$28581 ( \28924 , \28359 , \28923 );
xor \U$28582 ( \28925 , \28145 , \28149 );
and \U$28583 ( \28926 , \28925 , \28154 );
and \U$28584 ( \28927 , \28145 , \28149 );
or \U$28585 ( \28928 , \28926 , \28927 );
xor \U$28586 ( \28929 , \28260 , \28350 );
and \U$28587 ( \28930 , \28929 , \28355 );
and \U$28588 ( \28931 , \28260 , \28350 );
or \U$28589 ( \28932 , \28930 , \28931 );
xor \U$28590 ( \28933 , \28928 , \28932 );
xor \U$28591 ( \28934 , \28203 , \28213 );
and \U$28592 ( \28935 , \28934 , \28224 );
and \U$28593 ( \28936 , \28203 , \28213 );
or \U$28594 ( \28937 , \28935 , \28936 );
xor \U$28595 ( \28938 , \28094 , \28104 );
and \U$28596 ( \28939 , \28938 , \28114 );
and \U$28597 ( \28940 , \28094 , \28104 );
or \U$28598 ( \28941 , \28939 , \28940 );
not \U$28599 ( \28942 , \4712 );
not \U$28600 ( \28943 , \27968 );
or \U$28601 ( \28944 , \28942 , \28943 );
not \U$28602 ( \28945 , RIbb2e620_35);
not \U$28603 ( \28946 , \13916 );
or \U$28604 ( \28947 , \28945 , \28946 );
nand \U$28605 ( \28948 , \9278 , \11338 );
nand \U$28606 ( \28949 , \28947 , \28948 );
nand \U$28607 ( \28950 , \28949 , \5845 );
nand \U$28608 ( \28951 , \28944 , \28950 );
xor \U$28609 ( \28952 , \28941 , \28951 );
not \U$28610 ( \28953 , \14752 );
not \U$28611 ( \28954 , RIbb2df90_49);
not \U$28612 ( \28955 , \3021 );
or \U$28613 ( \28956 , \28954 , \28955 );
nand \U$28614 ( \28957 , \4020 , \12278 );
nand \U$28615 ( \28958 , \28956 , \28957 );
not \U$28616 ( \28959 , \28958 );
or \U$28617 ( \28960 , \28953 , \28959 );
nand \U$28618 ( \28961 , \27991 , \13295 );
nand \U$28619 ( \28962 , \28960 , \28961 );
xor \U$28620 ( \28963 , \28952 , \28962 );
xor \U$28621 ( \28964 , \28937 , \28963 );
xor \U$28622 ( \28965 , \28171 , \28182 );
and \U$28623 ( \28966 , \28965 , \28192 );
and \U$28624 ( \28967 , \28171 , \28182 );
or \U$28625 ( \28968 , \28966 , \28967 );
xor \U$28626 ( \28969 , \28964 , \28968 );
not \U$28627 ( \28970 , \27994 );
not \U$28628 ( \28971 , \27962 );
or \U$28629 ( \28972 , \28970 , \28971 );
or \U$28630 ( \28973 , \27962 , \27994 );
nand \U$28631 ( \28974 , \28973 , \28038 );
nand \U$28632 ( \28975 , \28972 , \28974 );
xor \U$28633 ( \28976 , \28969 , \28975 );
nand \U$28634 ( \28977 , \28086 , \28093 );
not \U$28635 ( \28978 , \854 );
and \U$28636 ( \28979 , \16747 , RIbb2eda0_19);
not \U$28637 ( \28980 , \16747 );
and \U$28638 ( \28981 , \28980 , \5277 );
or \U$28639 ( \28982 , \28979 , \28981 );
not \U$28640 ( \28983 , \28982 );
or \U$28641 ( \28984 , \28978 , \28983 );
nand \U$28642 ( \28985 , \28110 , \853 );
nand \U$28643 ( \28986 , \28984 , \28985 );
xor \U$28644 ( \28987 , \28977 , \28986 );
not \U$28645 ( \28988 , \28003 );
not \U$28646 ( \28989 , \2077 );
or \U$28647 ( \28990 , \28988 , \28989 );
and \U$28648 ( \28991 , RIbb2ecb0_21, \16561 );
not \U$28649 ( \28992 , RIbb2ecb0_21);
and \U$28650 ( \28993 , \28992 , \16566 );
nor \U$28651 ( \28994 , \28991 , \28993 );
or \U$28652 ( \28995 , \28994 , \7768 );
nand \U$28653 ( \28996 , \28990 , \28995 );
xnor \U$28654 ( \28997 , \28987 , \28996 );
not \U$28655 ( \28998 , \17470 );
and \U$28656 ( \28999 , RIbb2dae0_59, \17207 );
not \U$28657 ( \29000 , RIbb2dae0_59);
and \U$28658 ( \29001 , \29000 , \26831 );
or \U$28659 ( \29002 , \28999 , \29001 );
not \U$28660 ( \29003 , \29002 );
or \U$28661 ( \29004 , \28998 , \29003 );
nand \U$28662 ( \29005 , \28169 , \16271 );
nand \U$28663 ( \29006 , \29004 , \29005 );
xor \U$28664 ( \29007 , \28997 , \29006 );
not \U$28665 ( \29008 , \12774 );
not \U$28666 ( \29009 , \28035 );
or \U$28667 ( \29010 , \29008 , \29009 );
and \U$28668 ( \29011 , RIbb2dea0_51, \13836 );
not \U$28669 ( \29012 , RIbb2dea0_51);
and \U$28670 ( \29013 , \29012 , \3228 );
or \U$28671 ( \29014 , \29011 , \29013 );
nand \U$28672 ( \29015 , \29014 , \12692 );
nand \U$28673 ( \29016 , \29010 , \29015 );
xor \U$28674 ( \29017 , \29007 , \29016 );
not \U$28675 ( \29018 , \12965 );
not \U$28676 ( \29019 , RIbb2e080_47);
not \U$28677 ( \29020 , \25942 );
or \U$28678 ( \29021 , \29019 , \29020 );
nand \U$28679 ( \29022 , \13732 , \10113 );
nand \U$28680 ( \29023 , \29021 , \29022 );
not \U$28681 ( \29024 , \29023 );
or \U$28682 ( \29025 , \29018 , \29024 );
nand \U$28683 ( \29026 , \27945 , \11176 );
nand \U$28684 ( \29027 , \29025 , \29026 );
not \U$28685 ( \29028 , \17563 );
not \U$28686 ( \29029 , \28190 );
or \U$28687 ( \29030 , \29028 , \29029 );
not \U$28688 ( \29031 , RIbb2ddb0_53);
not \U$28689 ( \29032 , \3141 );
or \U$28690 ( \29033 , \29031 , \29032 );
nand \U$28691 ( \29034 , \26851 , \16210 );
nand \U$28692 ( \29035 , \29033 , \29034 );
nand \U$28693 ( \29036 , \14930 , \29035 );
nand \U$28694 ( \29037 , \29030 , \29036 );
xor \U$28695 ( \29038 , \29027 , \29037 );
not \U$28696 ( \29039 , \19101 );
not \U$28697 ( \29040 , \27980 );
or \U$28698 ( \29041 , \29039 , \29040 );
not \U$28699 ( \29042 , RIbb2dbd0_57);
not \U$28700 ( \29043 , \4449 );
or \U$28701 ( \29044 , \29042 , \29043 );
nand \U$28702 ( \29045 , \9984 , \17097 );
nand \U$28703 ( \29046 , \29044 , \29045 );
nand \U$28704 ( \29047 , \29046 , \17397 );
nand \U$28705 ( \29048 , \29041 , \29047 );
xor \U$28706 ( \29049 , \29038 , \29048 );
xor \U$28707 ( \29050 , \29017 , \29049 );
xor \U$28708 ( \29051 , \28302 , \28306 );
and \U$28709 ( \29052 , \29051 , \28312 );
and \U$28710 ( \29053 , \28302 , \28306 );
or \U$28711 ( \29054 , \29052 , \29053 );
xor \U$28712 ( \29055 , \29050 , \29054 );
xor \U$28713 ( \29056 , \28976 , \29055 );
xor \U$28714 ( \29057 , \28231 , \28235 );
and \U$28715 ( \29058 , \29057 , \28259 );
and \U$28716 ( \29059 , \28231 , \28235 );
or \U$28717 ( \29060 , \29058 , \29059 );
xor \U$28718 ( \29061 , \29056 , \29060 );
not \U$28719 ( \29062 , \28348 );
not \U$28720 ( \29063 , \28266 );
or \U$28721 ( \29064 , \29062 , \29063 );
not \U$28722 ( \29065 , \28347 );
not \U$28723 ( \29066 , \28266 );
not \U$28724 ( \29067 , \29066 );
or \U$28725 ( \29068 , \29065 , \29067 );
nand \U$28726 ( \29069 , \29068 , \28270 );
nand \U$28727 ( \29070 , \29064 , \29069 );
xor \U$28728 ( \29071 , \29061 , \29070 );
not \U$28729 ( \29072 , \28346 );
not \U$28730 ( \29073 , \29072 );
not \U$28731 ( \29074 , \28323 );
or \U$28732 ( \29075 , \29073 , \29074 );
not \U$28733 ( \29076 , \28346 );
not \U$28734 ( \29077 , \28324 );
or \U$28735 ( \29078 , \29076 , \29077 );
buf \U$28736 ( \29079 , \28313 );
nand \U$28737 ( \29080 , \29078 , \29079 );
nand \U$28738 ( \29081 , \29075 , \29080 );
or \U$28739 ( \29082 , \28339 , \28329 );
nand \U$28740 ( \29083 , \29082 , \28345 );
nand \U$28741 ( \29084 , \28329 , \28340 );
and \U$28742 ( \29085 , \29083 , \29084 );
not \U$28743 ( \29086 , \28225 );
not \U$28744 ( \29087 , \28193 );
or \U$28745 ( \29088 , \29086 , \29087 );
or \U$28746 ( \29089 , \28193 , \28225 );
nand \U$28747 ( \29090 , \29089 , \28164 );
nand \U$28748 ( \29091 , \29088 , \29090 );
xor \U$28749 ( \29092 , \29085 , \29091 );
not \U$28750 ( \29093 , \27939 );
not \U$28751 ( \29094 , \27949 );
or \U$28752 ( \29095 , \29093 , \29094 );
or \U$28753 ( \29096 , \27949 , \27939 );
nand \U$28754 ( \29097 , \29096 , \27961 );
nand \U$28755 ( \29098 , \29095 , \29097 );
not \U$28756 ( \29099 , \20792 );
not \U$28757 ( \29100 , RIbb2e530_37);
not \U$28758 ( \29101 , \12210 );
or \U$28759 ( \29102 , \29100 , \29101 );
nand \U$28760 ( \29103 , \8318 , \6246 );
nand \U$28761 ( \29104 , \29102 , \29103 );
not \U$28762 ( \29105 , \29104 );
or \U$28763 ( \29106 , \29099 , \29105 );
nand \U$28764 ( \29107 , \28070 , \6251 );
nand \U$28765 ( \29108 , \29106 , \29107 );
not \U$28766 ( \29109 , \7104 );
and \U$28767 ( \29110 , RIbb2e440_39, \19868 );
not \U$28768 ( \29111 , RIbb2e440_39);
and \U$28769 ( \29112 , \29111 , \25844 );
or \U$28770 ( \29113 , \29110 , \29112 );
not \U$28771 ( \29114 , \29113 );
or \U$28772 ( \29115 , \29109 , \29114 );
nand \U$28773 ( \29116 , \28059 , \7102 );
nand \U$28774 ( \29117 , \29115 , \29116 );
not \U$28775 ( \29118 , \29117 );
and \U$28776 ( \29119 , \29108 , \29118 );
not \U$28777 ( \29120 , \29108 );
and \U$28778 ( \29121 , \29120 , \29117 );
or \U$28779 ( \29122 , \29119 , \29121 );
not \U$28780 ( \29123 , \28122 );
not \U$28781 ( \29124 , \8363 );
and \U$28782 ( \29125 , \29123 , \29124 );
not \U$28783 ( \29126 , RIbb2e350_41);
not \U$28784 ( \29127 , \18564 );
or \U$28785 ( \29128 , \29126 , \29127 );
nand \U$28786 ( \29129 , \7308 , \9402 );
nand \U$28787 ( \29130 , \29128 , \29129 );
and \U$28788 ( \29131 , \29130 , \8354 );
nor \U$28789 ( \29132 , \29125 , \29131 );
buf \U$28790 ( \29133 , \29132 );
and \U$28791 ( \29134 , \29122 , \29133 );
not \U$28792 ( \29135 , \29122 );
not \U$28793 ( \29136 , \29133 );
and \U$28794 ( \29137 , \29135 , \29136 );
nor \U$28795 ( \29138 , \29134 , \29137 );
xor \U$28796 ( \29139 , \29098 , \29138 );
and \U$28797 ( \29140 , \9098 , \28220 );
not \U$28798 ( \29141 , RIbb2e260_43);
not \U$28799 ( \29142 , \10555 );
or \U$28800 ( \29143 , \29141 , \29142 );
nand \U$28801 ( \29144 , \9020 , \17231 );
nand \U$28802 ( \29145 , \29143 , \29144 );
and \U$28803 ( \29146 , \29145 , \9099 );
nor \U$28804 ( \29147 , \29140 , \29146 );
not \U$28805 ( \29148 , \29147 );
not \U$28806 ( \29149 , \4075 );
not \U$28807 ( \29150 , RIbb2e710_33);
not \U$28808 ( \29151 , \12233 );
or \U$28809 ( \29152 , \29150 , \29151 );
nand \U$28810 ( \29153 , \10301 , \2935 );
nand \U$28811 ( \29154 , \29152 , \29153 );
not \U$28812 ( \29155 , \29154 );
or \U$28813 ( \29156 , \29149 , \29155 );
nand \U$28814 ( \29157 , \28134 , \3886 );
nand \U$28815 ( \29158 , \29156 , \29157 );
not \U$28816 ( \29159 , \29158 );
or \U$28817 ( \29160 , \29148 , \29159 );
or \U$28818 ( \29161 , \29147 , \29158 );
nand \U$28819 ( \29162 , \29160 , \29161 );
not \U$28820 ( \29163 , \29162 );
not \U$28821 ( \29164 , \2939 );
not \U$28822 ( \29165 , \28199 );
or \U$28823 ( \29166 , \29164 , \29165 );
not \U$28824 ( \29167 , RIbb2e800_31);
not \U$28825 ( \29168 , \12260 );
or \U$28826 ( \29169 , \29167 , \29168 );
nand \U$28827 ( \29170 , \12261 , \9169 );
nand \U$28828 ( \29171 , \29169 , \29170 );
nand \U$28829 ( \29172 , \29171 , \3613 );
nand \U$28830 ( \29173 , \29166 , \29172 );
not \U$28831 ( \29174 , \29173 );
not \U$28832 ( \29175 , \29174 );
and \U$28833 ( \29176 , \29163 , \29175 );
and \U$28834 ( \29177 , \29162 , \29174 );
nor \U$28835 ( \29178 , \29176 , \29177 );
not \U$28836 ( \29179 , \29178 );
xor \U$28837 ( \29180 , \29139 , \29179 );
xor \U$28838 ( \29181 , \29092 , \29180 );
xor \U$28839 ( \29182 , \29081 , \29181 );
not \U$28840 ( \29183 , \28143 );
not \U$28841 ( \29184 , \28044 );
or \U$28842 ( \29185 , \29183 , \29184 );
or \U$28843 ( \29186 , \28044 , \28143 );
nand \U$28844 ( \29187 , \29186 , \28048 );
nand \U$28845 ( \29188 , \29185 , \29187 );
xor \U$28846 ( \29189 , \29182 , \29188 );
not \U$28847 ( \29190 , RIbb2d888_64);
not \U$28848 ( \29191 , RIbb2d900_63);
not \U$28849 ( \29192 , \15582 );
or \U$28850 ( \29193 , \29191 , \29192 );
nand \U$28851 ( \29194 , \12036 , \17270 );
nand \U$28852 ( \29195 , \29193 , \29194 );
not \U$28853 ( \29196 , \29195 );
or \U$28854 ( \29197 , \29190 , \29196 );
nand \U$28855 ( \29198 , \27937 , \17275 );
nand \U$28856 ( \29199 , \29197 , \29198 );
not \U$28857 ( \29200 , \16533 );
not \U$28858 ( \29201 , RIbb2d9f0_61);
not \U$28859 ( \29202 , \13619 );
or \U$28860 ( \29203 , \29201 , \29202 );
nand \U$28861 ( \29204 , \1386 , \16254 );
nand \U$28862 ( \29205 , \29203 , \29204 );
not \U$28863 ( \29206 , \29205 );
or \U$28864 ( \29207 , \29200 , \29206 );
nand \U$28865 ( \29208 , \16541 , \28180 );
nand \U$28866 ( \29209 , \29207 , \29208 );
xor \U$28867 ( \29210 , \29199 , \29209 );
not \U$28868 ( \29211 , \14613 );
not \U$28869 ( \29212 , \27959 );
or \U$28870 ( \29213 , \29211 , \29212 );
and \U$28871 ( \29214 , RIbb2dcc0_55, \3517 );
not \U$28872 ( \29215 , RIbb2dcc0_55);
and \U$28873 ( \29216 , \29215 , \3343 );
or \U$28874 ( \29217 , \29214 , \29216 );
nand \U$28875 ( \29218 , \29217 , \15181 );
nand \U$28876 ( \29219 , \29213 , \29218 );
xor \U$28877 ( \29220 , \29210 , \29219 );
xor \U$28878 ( \29221 , \27972 , \27982 );
and \U$28879 ( \29222 , \29221 , \27993 );
and \U$28880 ( \29223 , \27972 , \27982 );
or \U$28881 ( \29224 , \29222 , \29223 );
xor \U$28882 ( \29225 , \29220 , \29224 );
xor \U$28883 ( \29226 , \28021 , \28025 );
and \U$28884 ( \29227 , \29226 , \28037 );
and \U$28885 ( \29228 , \28021 , \28025 );
or \U$28886 ( \29229 , \29227 , \29228 );
xor \U$28887 ( \29230 , \29225 , \29229 );
not \U$28888 ( \29231 , \28300 );
not \U$28889 ( \29232 , \28290 );
or \U$28890 ( \29233 , \29231 , \29232 );
or \U$28891 ( \29234 , \28290 , \28300 );
nand \U$28892 ( \29235 , \29234 , \28280 );
nand \U$28893 ( \29236 , \29233 , \29235 );
not \U$28894 ( \29237 , \28020 );
not \U$28895 ( \29238 , \28005 );
nand \U$28896 ( \29239 , \29237 , \29238 );
and \U$28897 ( \29240 , \29239 , \28009 );
not \U$28898 ( \29241 , \28020 );
nor \U$28899 ( \29242 , \29241 , \29238 );
nor \U$28900 ( \29243 , \29240 , \29242 );
xor \U$28901 ( \29244 , \29236 , \29243 );
not \U$28902 ( \29245 , \29244 );
xor \U$28903 ( \29246 , \28115 , \28125 );
and \U$28904 ( \29247 , \29246 , \28136 );
and \U$28905 ( \29248 , \28115 , \28125 );
or \U$28906 ( \29249 , \29247 , \29248 );
not \U$28907 ( \29250 , \29249 );
or \U$28908 ( \29251 , \29245 , \29250 );
or \U$28909 ( \29252 , \29249 , \29244 );
nand \U$28910 ( \29253 , \29251 , \29252 );
and \U$28911 ( \29254 , \17506 , \997 );
not \U$28912 ( \29255 , \1517 );
and \U$28913 ( \29256 , RIbb2ef80_15, \16819 );
not \U$28914 ( \29257 , RIbb2ef80_15);
and \U$28915 ( \29258 , \29257 , \17529 );
or \U$28916 ( \29259 , \29256 , \29258 );
not \U$28917 ( \29260 , \29259 );
or \U$28918 ( \29261 , \29255 , \29260 );
nand \U$28919 ( \29262 , \28078 , \1444 );
nand \U$28920 ( \29263 , \29261 , \29262 );
xor \U$28921 ( \29264 , \29254 , \29263 );
not \U$28922 ( \29265 , \831 );
not \U$28923 ( \29266 , \28100 );
or \U$28924 ( \29267 , \29265 , \29266 );
not \U$28925 ( \29268 , RIbb2ee90_17);
not \U$28926 ( \29269 , \16554 );
or \U$28927 ( \29270 , \29268 , \29269 );
not \U$28928 ( \29271 , \16554 );
nand \U$28929 ( \29272 , \29271 , \816 );
nand \U$28930 ( \29273 , \29270 , \29272 );
nand \U$28931 ( \29274 , \29273 , \835 );
nand \U$28932 ( \29275 , \29267 , \29274 );
xor \U$28933 ( \29276 , \29264 , \29275 );
not \U$28934 ( \29277 , \3406 );
not \U$28935 ( \29278 , \28286 );
or \U$28936 ( \29279 , \29277 , \29278 );
not \U$28937 ( \29280 , RIbb2ebc0_23);
not \U$28938 ( \29281 , \18353 );
or \U$28939 ( \29282 , \29280 , \29281 );
nand \U$28940 ( \29283 , \14526 , \3401 );
nand \U$28941 ( \29284 , \29282 , \29283 );
nand \U$28942 ( \29285 , \29284 , \3382 );
nand \U$28943 ( \29286 , \29279 , \29285 );
xor \U$28944 ( \29287 , \29276 , \29286 );
not \U$28945 ( \29288 , \2925 );
not \U$28946 ( \29289 , RIbb2e8f0_29);
not \U$28947 ( \29290 , \13680 );
or \U$28948 ( \29291 , \29289 , \29290 );
nand \U$28949 ( \29292 , \12175 , \3440 );
nand \U$28950 ( \29293 , \29291 , \29292 );
not \U$28951 ( \29294 , \29293 );
or \U$28952 ( \29295 , \29288 , \29294 );
nand \U$28953 ( \29296 , \28016 , \2921 );
nand \U$28954 ( \29297 , \29295 , \29296 );
xor \U$28955 ( \29298 , \29287 , \29297 );
not \U$28956 ( \29299 , \10119 );
not \U$28957 ( \29300 , RIbb2e170_45);
not \U$28958 ( \29301 , \13552 );
or \U$28959 ( \29302 , \29300 , \29301 );
nand \U$28960 ( \29303 , \13551 , \17970 );
nand \U$28961 ( \29304 , \29302 , \29303 );
not \U$28962 ( \29305 , \29304 );
or \U$28963 ( \29306 , \29299 , \29305 );
nand \U$28964 ( \29307 , \10117 , \28209 );
nand \U$28965 ( \29308 , \29306 , \29307 );
not \U$28966 ( \29309 , \3445 );
not \U$28967 ( \29310 , \28296 );
or \U$28968 ( \29311 , \29309 , \29310 );
not \U$28969 ( \29312 , RIbb2e9e0_27);
not \U$28970 ( \29313 , \14838 );
or \U$28971 ( \29314 , \29312 , \29313 );
nand \U$28972 ( \29315 , \12347 , \3454 );
nand \U$28973 ( \29316 , \29314 , \29315 );
nand \U$28974 ( \29317 , \29316 , \3465 );
nand \U$28975 ( \29318 , \29311 , \29317 );
not \U$28976 ( \29319 , \29318 );
not \U$28977 ( \29320 , \2980 );
not \U$28978 ( \29321 , \28278 );
or \U$28979 ( \29322 , \29320 , \29321 );
xor \U$28980 ( \29323 , RIbb2ead0_25, \13545 );
nand \U$28981 ( \29324 , \29323 , \2963 );
nand \U$28982 ( \29325 , \29322 , \29324 );
not \U$28983 ( \29326 , \29325 );
not \U$28984 ( \29327 , \29326 );
or \U$28985 ( \29328 , \29319 , \29327 );
or \U$28986 ( \29329 , \29318 , \29326 );
nand \U$28987 ( \29330 , \29328 , \29329 );
xor \U$28988 ( \29331 , \29308 , \29330 );
xor \U$28989 ( \29332 , \29298 , \29331 );
xor \U$28990 ( \29333 , \28052 , \28061 );
and \U$28991 ( \29334 , \29333 , \28072 );
and \U$28992 ( \29335 , \28052 , \28061 );
or \U$28993 ( \29336 , \29334 , \29335 );
xor \U$28994 ( \29337 , \29332 , \29336 );
xor \U$28995 ( \29338 , \29253 , \29337 );
xor \U$28996 ( \29339 , \28073 , \28137 );
and \U$28997 ( \29340 , \29339 , \28142 );
and \U$28998 ( \29341 , \28073 , \28137 );
or \U$28999 ( \29342 , \29340 , \29341 );
xor \U$29000 ( \29343 , \29338 , \29342 );
xor \U$29001 ( \29344 , \29230 , \29343 );
not \U$29002 ( \29345 , \28240 );
nand \U$29003 ( \29346 , \29345 , \28251 );
and \U$29004 ( \29347 , \29346 , \28245 );
and \U$29005 ( \29348 , \28240 , \28250 );
nor \U$29006 ( \29349 , \29347 , \29348 );
not \U$29007 ( \29350 , \29349 );
xnor \U$29008 ( \29351 , \29344 , \29350 );
xor \U$29009 ( \29352 , \29189 , \29351 );
xnor \U$29010 ( \29353 , \29071 , \29352 );
xor \U$29011 ( \29354 , \28933 , \29353 );
not \U$29012 ( \29355 , \29354 );
xor \U$29013 ( \29356 , \28155 , \28159 );
and \U$29014 ( \29357 , \29356 , \28356 );
and \U$29015 ( \29358 , \28155 , \28159 );
or \U$29016 ( \29359 , \29357 , \29358 );
not \U$29017 ( \29360 , \29359 );
nand \U$29018 ( \29361 , \29355 , \29360 );
not \U$29019 ( \29362 , \28357 );
not \U$29020 ( \29363 , \27928 );
nand \U$29021 ( \29364 , \29362 , \29363 );
nand \U$29022 ( \29365 , \28924 , \29361 , \29364 );
not \U$29023 ( \29366 , \836 );
not \U$29024 ( \29367 , RIbb2ee90_17);
not \U$29025 ( \29368 , \23185 );
or \U$29026 ( \29369 , \29367 , \29368 );
nand \U$29027 ( \29370 , \16829 , \816 );
nand \U$29028 ( \29371 , \29369 , \29370 );
not \U$29029 ( \29372 , \29371 );
or \U$29030 ( \29373 , \29366 , \29372 );
nand \U$29031 ( \29374 , \831 , \29273 );
nand \U$29032 ( \29375 , \29373 , \29374 );
xor \U$29033 ( \29376 , \29254 , \29263 );
and \U$29034 ( \29377 , \29376 , \29275 );
and \U$29035 ( \29378 , \29254 , \29263 );
or \U$29036 ( \29379 , \29377 , \29378 );
xor \U$29037 ( \29380 , \29375 , \29379 );
not \U$29038 ( \29381 , \3445 );
not \U$29039 ( \29382 , \29316 );
or \U$29040 ( \29383 , \29381 , \29382 );
not \U$29041 ( \29384 , RIbb2e9e0_27);
not \U$29042 ( \29385 , \12322 );
or \U$29043 ( \29386 , \29384 , \29385 );
nand \U$29044 ( \29387 , \12932 , \11284 );
nand \U$29045 ( \29388 , \29386 , \29387 );
nand \U$29046 ( \29389 , \29388 , \3465 );
nand \U$29047 ( \29390 , \29383 , \29389 );
xor \U$29048 ( \29391 , \29380 , \29390 );
not \U$29049 ( \29392 , \17470 );
and \U$29050 ( \29393 , RIbb2dae0_59, \17386 );
not \U$29051 ( \29394 , RIbb2dae0_59);
and \U$29052 ( \29395 , \29394 , \3821 );
or \U$29053 ( \29396 , \29393 , \29395 );
not \U$29054 ( \29397 , \29396 );
or \U$29055 ( \29398 , \29392 , \29397 );
not \U$29056 ( \29399 , \16271 );
not \U$29057 ( \29400 , \29399 );
nand \U$29058 ( \29401 , \29400 , \29002 );
nand \U$29059 ( \29402 , \29398 , \29401 );
xor \U$29060 ( \29403 , \29391 , \29402 );
not \U$29061 ( \29404 , \12692 );
and \U$29062 ( \29405 , RIbb2dea0_51, \4638 );
not \U$29063 ( \29406 , RIbb2dea0_51);
and \U$29064 ( \29407 , \29406 , \4637 );
or \U$29065 ( \29408 , \29405 , \29407 );
not \U$29066 ( \29409 , \29408 );
or \U$29067 ( \29410 , \29404 , \29409 );
nand \U$29068 ( \29411 , \29014 , \12774 );
nand \U$29069 ( \29412 , \29410 , \29411 );
xnor \U$29070 ( \29413 , \29403 , \29412 );
not \U$29071 ( \29414 , \29236 );
nand \U$29072 ( \29415 , \29414 , \29243 );
not \U$29073 ( \29416 , \29415 );
not \U$29074 ( \29417 , \29249 );
or \U$29075 ( \29418 , \29416 , \29417 );
not \U$29076 ( \29419 , \29243 );
nand \U$29077 ( \29420 , \29419 , \29236 );
nand \U$29078 ( \29421 , \29418 , \29420 );
xor \U$29079 ( \29422 , \29413 , \29421 );
xor \U$29080 ( \29423 , \29298 , \29331 );
and \U$29081 ( \29424 , \29423 , \29336 );
and \U$29082 ( \29425 , \29298 , \29331 );
or \U$29083 ( \29426 , \29424 , \29425 );
xor \U$29084 ( \29427 , \29422 , \29426 );
xor \U$29085 ( \29428 , \29253 , \29337 );
and \U$29086 ( \29429 , \29428 , \29342 );
and \U$29087 ( \29430 , \29253 , \29337 );
or \U$29088 ( \29431 , \29429 , \29430 );
not \U$29089 ( \29432 , \29431 );
xor \U$29090 ( \29433 , \29427 , \29432 );
not \U$29091 ( \29434 , \29091 );
nand \U$29092 ( \29435 , \29434 , \29180 );
not \U$29093 ( \29436 , \29085 );
and \U$29094 ( \29437 , \29435 , \29436 );
not \U$29095 ( \29438 , \29091 );
nor \U$29096 ( \29439 , \29438 , \29180 );
nor \U$29097 ( \29440 , \29437 , \29439 );
xor \U$29098 ( \29441 , \29433 , \29440 );
not \U$29099 ( \29442 , \29441 );
not \U$29100 ( \29443 , \29230 );
not \U$29101 ( \29444 , \29350 );
or \U$29102 ( \29445 , \29443 , \29444 );
not \U$29103 ( \29446 , \29230 );
not \U$29104 ( \29447 , \29446 );
not \U$29105 ( \29448 , \29349 );
or \U$29106 ( \29449 , \29447 , \29448 );
nand \U$29107 ( \29450 , \29449 , \29343 );
nand \U$29108 ( \29451 , \29445 , \29450 );
not \U$29109 ( \29452 , \29224 );
not \U$29110 ( \29453 , \29220 );
or \U$29111 ( \29454 , \29452 , \29453 );
or \U$29112 ( \29455 , \29220 , \29224 );
nand \U$29113 ( \29456 , \29455 , \29229 );
nand \U$29114 ( \29457 , \29454 , \29456 );
xor \U$29115 ( \29458 , \29017 , \29049 );
and \U$29116 ( \29459 , \29458 , \29054 );
and \U$29117 ( \29460 , \29017 , \29049 );
or \U$29118 ( \29461 , \29459 , \29460 );
xor \U$29119 ( \29462 , \29457 , \29461 );
not \U$29120 ( \29463 , \5845 );
not \U$29121 ( \29464 , RIbb2e620_35);
not \U$29122 ( \29465 , \10175 );
or \U$29123 ( \29466 , \29464 , \29465 );
not \U$29124 ( \29467 , \13863 );
nand \U$29125 ( \29468 , \29467 , \3866 );
nand \U$29126 ( \29469 , \29466 , \29468 );
not \U$29127 ( \29470 , \29469 );
or \U$29128 ( \29471 , \29463 , \29470 );
nand \U$29129 ( \29472 , \28949 , \4712 );
nand \U$29130 ( \29473 , \29471 , \29472 );
not \U$29131 ( \29474 , \17275 );
not \U$29132 ( \29475 , \29195 );
or \U$29133 ( \29476 , \29474 , \29475 );
not \U$29134 ( \29477 , RIbb2d900_63);
not \U$29135 ( \29478 , \13707 );
or \U$29136 ( \29479 , \29477 , \29478 );
nand \U$29137 ( \29480 , \17262 , \1111 );
nand \U$29138 ( \29481 , \29479 , \29480 );
nand \U$29139 ( \29482 , \29481 , RIbb2d888_64);
nand \U$29140 ( \29483 , \29476 , \29482 );
xor \U$29141 ( \29484 , \29473 , \29483 );
not \U$29142 ( \29485 , \12167 );
not \U$29143 ( \29486 , \28958 );
or \U$29144 ( \29487 , \29485 , \29486 );
not \U$29145 ( \29488 , RIbb2df90_49);
not \U$29146 ( \29489 , \16898 );
or \U$29147 ( \29490 , \29488 , \29489 );
nand \U$29148 ( \29491 , \25703 , \12278 );
nand \U$29149 ( \29492 , \29490 , \29491 );
nand \U$29150 ( \29493 , \29492 , \16427 );
nand \U$29151 ( \29494 , \29487 , \29493 );
xor \U$29152 ( \29495 , \29484 , \29494 );
not \U$29153 ( \29496 , \16541 );
not \U$29154 ( \29497 , \29205 );
or \U$29155 ( \29498 , \29496 , \29497 );
not \U$29156 ( \29499 , RIbb2d9f0_61);
not \U$29157 ( \29500 , \20215 );
or \U$29158 ( \29501 , \29499 , \29500 );
nand \U$29159 ( \29502 , \1169 , \16254 );
nand \U$29160 ( \29503 , \29501 , \29502 );
nand \U$29161 ( \29504 , \29503 , \16533 );
nand \U$29162 ( \29505 , \29498 , \29504 );
not \U$29163 ( \29506 , \14930 );
and \U$29164 ( \29507 , \4219 , RIbb2ddb0_53);
not \U$29165 ( \29508 , \4219 );
and \U$29166 ( \29509 , \29508 , \13463 );
or \U$29167 ( \29510 , \29507 , \29509 );
not \U$29168 ( \29511 , \29510 );
or \U$29169 ( \29512 , \29506 , \29511 );
nand \U$29170 ( \29513 , \29035 , \17563 );
nand \U$29171 ( \29514 , \29512 , \29513 );
xor \U$29172 ( \29515 , \29505 , \29514 );
not \U$29173 ( \29516 , \15182 );
and \U$29174 ( \29517 , RIbb2dcc0_55, \2223 );
not \U$29175 ( \29518 , RIbb2dcc0_55);
and \U$29176 ( \29519 , \29518 , \2222 );
or \U$29177 ( \29520 , \29517 , \29519 );
not \U$29178 ( \29521 , \29520 );
or \U$29179 ( \29522 , \29516 , \29521 );
nand \U$29180 ( \29523 , \29217 , \22952 );
nand \U$29181 ( \29524 , \29522 , \29523 );
xor \U$29182 ( \29525 , \29515 , \29524 );
xor \U$29183 ( \29526 , \29495 , \29525 );
not \U$29184 ( \29527 , \19101 );
not \U$29185 ( \29528 , \29046 );
or \U$29186 ( \29529 , \29527 , \29528 );
not \U$29187 ( \29530 , RIbb2dbd0_57);
not \U$29188 ( \29531 , \3807 );
or \U$29189 ( \29532 , \29530 , \29531 );
nand \U$29190 ( \29533 , \1852 , \14602 );
nand \U$29191 ( \29534 , \29532 , \29533 );
nand \U$29192 ( \29535 , \29534 , \17100 );
nand \U$29193 ( \29536 , \29529 , \29535 );
not \U$29194 ( \29537 , \10119 );
not \U$29195 ( \29538 , RIbb2e170_45);
not \U$29196 ( \29539 , \4748 );
or \U$29197 ( \29540 , \29538 , \29539 );
nand \U$29198 ( \29541 , \3089 , \12003 );
nand \U$29199 ( \29542 , \29540 , \29541 );
not \U$29200 ( \29543 , \29542 );
or \U$29201 ( \29544 , \29537 , \29543 );
nand \U$29202 ( \29545 , \29304 , \10599 );
nand \U$29203 ( \29546 , \29544 , \29545 );
xor \U$29204 ( \29547 , \29536 , \29546 );
not \U$29205 ( \29548 , \11176 );
not \U$29206 ( \29549 , \29023 );
or \U$29207 ( \29550 , \29548 , \29549 );
not \U$29208 ( \29551 , RIbb2e080_47);
not \U$29209 ( \29552 , \3045 );
or \U$29210 ( \29553 , \29551 , \29552 );
nand \U$29211 ( \29554 , \14912 , \16163 );
nand \U$29212 ( \29555 , \29553 , \29554 );
nand \U$29213 ( \29556 , \29555 , \12965 );
nand \U$29214 ( \29557 , \29550 , \29556 );
xor \U$29215 ( \29558 , \29547 , \29557 );
xnor \U$29216 ( \29559 , \29526 , \29558 );
not \U$29217 ( \29560 , \29559 );
xnor \U$29218 ( \29561 , \29462 , \29560 );
and \U$29219 ( \29562 , \29451 , \29561 );
not \U$29220 ( \29563 , \29451 );
not \U$29221 ( \29564 , \29561 );
and \U$29222 ( \29565 , \29563 , \29564 );
nor \U$29223 ( \29566 , \29562 , \29565 );
not \U$29224 ( \29567 , \29566 );
xor \U$29225 ( \29568 , \29442 , \29567 );
xor \U$29226 ( \29569 , \29081 , \29181 );
and \U$29227 ( \29570 , \29569 , \29188 );
and \U$29228 ( \29571 , \29081 , \29181 );
or \U$29229 ( \29572 , \29570 , \29571 );
not \U$29230 ( \29573 , \29284 );
not \U$29231 ( \29574 , \3406 );
or \U$29232 ( \29575 , \29573 , \29574 );
not \U$29233 ( \29576 , RIbb2ebc0_23);
not \U$29234 ( \29577 , \18829 );
or \U$29235 ( \29578 , \29576 , \29577 );
nand \U$29236 ( \29579 , \13977 , \3388 );
nand \U$29237 ( \29580 , \29578 , \29579 );
nand \U$29238 ( \29581 , \29580 , \3381 );
nand \U$29239 ( \29582 , \29575 , \29581 );
not \U$29240 ( \29583 , \29582 );
not \U$29241 ( \29584 , \2963 );
not \U$29242 ( \29585 , RIbb2ead0_25);
not \U$29243 ( \29586 , \14624 );
or \U$29244 ( \29587 , \29585 , \29586 );
nand \U$29245 ( \29588 , \13210 , \18636 );
nand \U$29246 ( \29589 , \29587 , \29588 );
not \U$29247 ( \29590 , \29589 );
or \U$29248 ( \29591 , \29584 , \29590 );
nand \U$29249 ( \29592 , \29323 , \2979 );
nand \U$29250 ( \29593 , \29591 , \29592 );
not \U$29251 ( \29594 , \29593 );
not \U$29252 ( \29595 , \29594 );
or \U$29253 ( \29596 , \29583 , \29595 );
or \U$29254 ( \29597 , \29594 , \29582 );
nand \U$29255 ( \29598 , \29596 , \29597 );
not \U$29256 ( \29599 , \2078 );
not \U$29257 ( \29600 , RIbb2ecb0_21);
not \U$29258 ( \29601 , \16783 );
or \U$29259 ( \29602 , \29600 , \29601 );
nand \U$29260 ( \29603 , \15470 , \2249 );
nand \U$29261 ( \29604 , \29602 , \29603 );
not \U$29262 ( \29605 , \29604 );
or \U$29263 ( \29606 , \29599 , \29605 );
not \U$29264 ( \29607 , \28994 );
nand \U$29265 ( \29608 , \29607 , \2077 );
nand \U$29266 ( \29609 , \29606 , \29608 );
and \U$29267 ( \29610 , \29598 , \29609 );
not \U$29268 ( \29611 , \29598 );
not \U$29269 ( \29612 , \29609 );
and \U$29270 ( \29613 , \29611 , \29612 );
nor \U$29271 ( \29614 , \29610 , \29613 );
not \U$29272 ( \29615 , \29318 );
nand \U$29273 ( \29616 , \29615 , \29326 );
not \U$29274 ( \29617 , \29616 );
not \U$29275 ( \29618 , \29308 );
or \U$29276 ( \29619 , \29617 , \29618 );
nand \U$29277 ( \29620 , \29325 , \29318 );
nand \U$29278 ( \29621 , \29619 , \29620 );
xor \U$29279 ( \29622 , \29614 , \29621 );
xor \U$29280 ( \29623 , \28941 , \28951 );
and \U$29281 ( \29624 , \29623 , \28962 );
and \U$29282 ( \29625 , \28941 , \28951 );
or \U$29283 ( \29626 , \29624 , \29625 );
xor \U$29284 ( \29627 , \29622 , \29626 );
not \U$29285 ( \29628 , \29138 );
not \U$29286 ( \29629 , \29628 );
not \U$29287 ( \29630 , \29179 );
or \U$29288 ( \29631 , \29629 , \29630 );
not \U$29289 ( \29632 , \29178 );
not \U$29290 ( \29633 , \29138 );
or \U$29291 ( \29634 , \29632 , \29633 );
nand \U$29292 ( \29635 , \29634 , \29098 );
nand \U$29293 ( \29636 , \29631 , \29635 );
xor \U$29294 ( \29637 , \29627 , \29636 );
xor \U$29295 ( \29638 , \28937 , \28963 );
and \U$29296 ( \29639 , \29638 , \28968 );
and \U$29297 ( \29640 , \28937 , \28963 );
or \U$29298 ( \29641 , \29639 , \29640 );
xor \U$29299 ( \29642 , \29637 , \29641 );
not \U$29300 ( \29643 , \28975 );
not \U$29301 ( \29644 , \29643 );
not \U$29302 ( \29645 , \28969 );
not \U$29303 ( \29646 , \29645 );
or \U$29304 ( \29647 , \29644 , \29646 );
nand \U$29305 ( \29648 , \29647 , \29055 );
not \U$29306 ( \29649 , \29645 );
nand \U$29307 ( \29650 , \29649 , \28975 );
nand \U$29308 ( \29651 , \29648 , \29650 );
and \U$29309 ( \29652 , \29642 , \29651 );
not \U$29310 ( \29653 , \29642 );
not \U$29311 ( \29654 , \29651 );
and \U$29312 ( \29655 , \29653 , \29654 );
or \U$29313 ( \29656 , \29652 , \29655 );
xor \U$29314 ( \29657 , \29276 , \29286 );
and \U$29315 ( \29658 , \29657 , \29297 );
and \U$29316 ( \29659 , \29276 , \29286 );
or \U$29317 ( \29660 , \29658 , \29659 );
not \U$29318 ( \29661 , \29118 );
not \U$29319 ( \29662 , \29132 );
or \U$29320 ( \29663 , \29661 , \29662 );
nand \U$29321 ( \29664 , \29663 , \29108 );
not \U$29322 ( \29665 , \29132 );
nand \U$29323 ( \29666 , \29665 , \29117 );
nand \U$29324 ( \29667 , \29664 , \29666 );
xor \U$29325 ( \29668 , \29660 , \29667 );
nor \U$29326 ( \29669 , \29173 , \29158 );
or \U$29327 ( \29670 , \29669 , \29147 );
nand \U$29328 ( \29671 , \29158 , \29173 );
nand \U$29329 ( \29672 , \29670 , \29671 );
xor \U$29330 ( \29673 , \29668 , \29672 );
or \U$29331 ( \29674 , RIbb2eff8_14, RIbb2ef80_15);
nand \U$29332 ( \29675 , \29674 , \19064 );
and \U$29333 ( \29676 , RIbb2eff8_14, RIbb2ef80_15);
nor \U$29334 ( \29677 , \29676 , \906 );
and \U$29335 ( \29678 , \29675 , \29677 );
not \U$29336 ( \29679 , \997 );
not \U$29337 ( \29680 , RIbb2f070_13);
not \U$29338 ( \29681 , \17745 );
or \U$29339 ( \29682 , \29680 , \29681 );
nand \U$29340 ( \29683 , \27225 , \1656 );
nand \U$29341 ( \29684 , \29682 , \29683 );
not \U$29342 ( \29685 , \29684 );
or \U$29343 ( \29686 , \29679 , \29685 );
and \U$29344 ( \29687 , RIbb2f070_13, \17506 );
not \U$29345 ( \29688 , RIbb2f070_13);
and \U$29346 ( \29689 , \29688 , \19063 );
nor \U$29347 ( \29690 , \29687 , \29689 );
nand \U$29348 ( \29691 , \29690 , \915 );
nand \U$29349 ( \29692 , \29686 , \29691 );
xor \U$29350 ( \29693 , \29678 , \29692 );
not \U$29351 ( \29694 , \1517 );
and \U$29352 ( \29695 , RIbb2ef80_15, \17756 );
not \U$29353 ( \29696 , RIbb2ef80_15);
and \U$29354 ( \29697 , \29696 , \17751 );
or \U$29355 ( \29698 , \29695 , \29697 );
not \U$29356 ( \29699 , \29698 );
or \U$29357 ( \29700 , \29694 , \29699 );
nand \U$29358 ( \29701 , \29259 , \1444 );
nand \U$29359 ( \29702 , \29700 , \29701 );
xor \U$29360 ( \29703 , \29693 , \29702 );
not \U$29361 ( \29704 , \854 );
not \U$29362 ( \29705 , RIbb2eda0_19);
not \U$29363 ( \29706 , \23197 );
or \U$29364 ( \29707 , \29705 , \29706 );
nand \U$29365 ( \29708 , \16575 , \843 );
nand \U$29366 ( \29709 , \29707 , \29708 );
not \U$29367 ( \29710 , \29709 );
or \U$29368 ( \29711 , \29704 , \29710 );
nand \U$29369 ( \29712 , \28982 , \853 );
nand \U$29370 ( \29713 , \29711 , \29712 );
xor \U$29371 ( \29714 , \29703 , \29713 );
or \U$29372 ( \29715 , \28996 , \28986 );
not \U$29373 ( \29716 , \28977 );
nand \U$29374 ( \29717 , \29715 , \29716 );
nand \U$29375 ( \29718 , \28996 , \28986 );
and \U$29376 ( \29719 , \29717 , \29718 );
xor \U$29377 ( \29720 , \29714 , \29719 );
not \U$29378 ( \29721 , \6241 );
not \U$29379 ( \29722 , RIbb2e530_37);
not \U$29380 ( \29723 , \7298 );
or \U$29381 ( \29724 , \29722 , \29723 );
nand \U$29382 ( \29725 , \14673 , \6246 );
nand \U$29383 ( \29726 , \29724 , \29725 );
not \U$29384 ( \29727 , \29726 );
or \U$29385 ( \29728 , \29721 , \29727 );
nand \U$29386 ( \29729 , \29104 , \6251 );
nand \U$29387 ( \29730 , \29728 , \29729 );
xnor \U$29388 ( \29731 , \29720 , \29730 );
xor \U$29389 ( \29732 , \29199 , \29209 );
and \U$29390 ( \29733 , \29732 , \29219 );
and \U$29391 ( \29734 , \29199 , \29209 );
or \U$29392 ( \29735 , \29733 , \29734 );
xor \U$29393 ( \29736 , \29731 , \29735 );
xor \U$29394 ( \29737 , \28997 , \29006 );
and \U$29395 ( \29738 , \29737 , \29016 );
and \U$29396 ( \29739 , \28997 , \29006 );
or \U$29397 ( \29740 , \29738 , \29739 );
xor \U$29398 ( \29741 , \29736 , \29740 );
xor \U$29399 ( \29742 , \29673 , \29741 );
not \U$29400 ( \29743 , \8450 );
and \U$29401 ( \29744 , RIbb2e440_39, \15797 );
not \U$29402 ( \29745 , RIbb2e440_39);
and \U$29403 ( \29746 , \29745 , \15796 );
or \U$29404 ( \29747 , \29744 , \29746 );
not \U$29405 ( \29748 , \29747 );
or \U$29406 ( \29749 , \29743 , \29748 );
nand \U$29407 ( \29750 , \29113 , \7103 );
nand \U$29408 ( \29751 , \29749 , \29750 );
not \U$29409 ( \29752 , \29751 );
not \U$29410 ( \29753 , \10449 );
not \U$29411 ( \29754 , \29145 );
or \U$29412 ( \29755 , \29753 , \29754 );
not \U$29413 ( \29756 , RIbb2e260_43);
not \U$29414 ( \29757 , \4392 );
or \U$29415 ( \29758 , \29756 , \29757 );
nand \U$29416 ( \29759 , \20390 , \8347 );
nand \U$29417 ( \29760 , \29758 , \29759 );
nand \U$29418 ( \29761 , \29760 , \10451 );
nand \U$29419 ( \29762 , \29755 , \29761 );
not \U$29420 ( \29763 , \29762 );
not \U$29421 ( \29764 , \29763 );
or \U$29422 ( \29765 , \29752 , \29764 );
not \U$29423 ( \29766 , \29751 );
nand \U$29424 ( \29767 , \29766 , \29762 );
nand \U$29425 ( \29768 , \29765 , \29767 );
not \U$29426 ( \29769 , \8362 );
not \U$29427 ( \29770 , \29130 );
or \U$29428 ( \29771 , \29769 , \29770 );
and \U$29429 ( \29772 , \9108 , RIbb2e350_41);
not \U$29430 ( \29773 , \9108 );
and \U$29431 ( \29774 , \29773 , \7097 );
or \U$29432 ( \29775 , \29772 , \29774 );
nand \U$29433 ( \29776 , \29775 , \8353 );
nand \U$29434 ( \29777 , \29771 , \29776 );
xor \U$29435 ( \29778 , \29768 , \29777 );
not \U$29436 ( \29779 , \2925 );
not \U$29437 ( \29780 , RIbb2e8f0_29);
not \U$29438 ( \29781 , \11579 );
or \U$29439 ( \29782 , \29780 , \29781 );
nand \U$29440 ( \29783 , \14885 , \3440 );
nand \U$29441 ( \29784 , \29782 , \29783 );
not \U$29442 ( \29785 , \29784 );
or \U$29443 ( \29786 , \29779 , \29785 );
nand \U$29444 ( \29787 , \29293 , \2921 );
nand \U$29445 ( \29788 , \29786 , \29787 );
not \U$29446 ( \29789 , \4075 );
not \U$29447 ( \29790 , RIbb2e710_33);
not \U$29448 ( \29791 , \20044 );
or \U$29449 ( \29792 , \29790 , \29791 );
nand \U$29450 ( \29793 , \9841 , \3882 );
nand \U$29451 ( \29794 , \29792 , \29793 );
not \U$29452 ( \29795 , \29794 );
or \U$29453 ( \29796 , \29789 , \29795 );
nand \U$29454 ( \29797 , \29154 , \3886 );
nand \U$29455 ( \29798 , \29796 , \29797 );
xor \U$29456 ( \29799 , \29788 , \29798 );
not \U$29457 ( \29800 , \2940 );
not \U$29458 ( \29801 , \29171 );
or \U$29459 ( \29802 , \29800 , \29801 );
not \U$29460 ( \29803 , RIbb2e800_31);
not \U$29461 ( \29804 , \14563 );
or \U$29462 ( \29805 , \29803 , \29804 );
nand \U$29463 ( \29806 , \10764 , \8810 );
nand \U$29464 ( \29807 , \29805 , \29806 );
nand \U$29465 ( \29808 , \29807 , \2941 );
nand \U$29466 ( \29809 , \29802 , \29808 );
xnor \U$29467 ( \29810 , \29799 , \29809 );
xnor \U$29468 ( \29811 , \29778 , \29810 );
not \U$29469 ( \29812 , \29027 );
not \U$29470 ( \29813 , \29048 );
or \U$29471 ( \29814 , \29812 , \29813 );
or \U$29472 ( \29815 , \29048 , \29027 );
nand \U$29473 ( \29816 , \29815 , \29037 );
nand \U$29474 ( \29817 , \29814 , \29816 );
not \U$29475 ( \29818 , \29817 );
and \U$29476 ( \29819 , \29811 , \29818 );
not \U$29477 ( \29820 , \29811 );
and \U$29478 ( \29821 , \29820 , \29817 );
nor \U$29479 ( \29822 , \29819 , \29821 );
not \U$29480 ( \29823 , \29822 );
xnor \U$29481 ( \29824 , \29742 , \29823 );
xor \U$29482 ( \29825 , \29656 , \29824 );
xor \U$29483 ( \29826 , \29572 , \29825 );
xor \U$29484 ( \29827 , \29056 , \29060 );
and \U$29485 ( \29828 , \29827 , \29070 );
and \U$29486 ( \29829 , \29056 , \29060 );
or \U$29487 ( \29830 , \29828 , \29829 );
xor \U$29488 ( \29831 , \29826 , \29830 );
xor \U$29489 ( \29832 , \29568 , \29831 );
not \U$29490 ( \29833 , \29189 );
buf \U$29491 ( \29834 , \29351 );
nand \U$29492 ( \29835 , \29833 , \29834 );
not \U$29493 ( \29836 , \29835 );
not \U$29494 ( \29837 , \29071 );
or \U$29495 ( \29838 , \29836 , \29837 );
or \U$29496 ( \29839 , \29833 , \29834 );
nand \U$29497 ( \29840 , \29838 , \29839 );
xor \U$29498 ( \29841 , \29832 , \29840 );
xor \U$29499 ( \29842 , \28928 , \28932 );
and \U$29500 ( \29843 , \29842 , \29353 );
and \U$29501 ( \29844 , \28928 , \28932 );
or \U$29502 ( \29845 , \29843 , \29844 );
nand \U$29503 ( \29846 , \29841 , \29845 );
nand \U$29504 ( \29847 , \29354 , \29359 );
and \U$29505 ( \29848 , \29846 , \29847 );
and \U$29506 ( \29849 , \29365 , \29848 );
buf \U$29507 ( \29850 , \29841 );
nor \U$29508 ( \29851 , \29850 , \29845 );
nor \U$29509 ( \29852 , \29849 , \29851 );
not \U$29510 ( \29853 , \29852 );
xor \U$29511 ( \29854 , \29614 , \29621 );
and \U$29512 ( \29855 , \29854 , \29626 );
and \U$29513 ( \29856 , \29614 , \29621 );
or \U$29514 ( \29857 , \29855 , \29856 );
not \U$29515 ( \29858 , \29857 );
not \U$29516 ( \29859 , \29809 );
not \U$29517 ( \29860 , \29788 );
or \U$29518 ( \29861 , \29859 , \29860 );
or \U$29519 ( \29862 , \29809 , \29788 );
nand \U$29520 ( \29863 , \29862 , \29798 );
nand \U$29521 ( \29864 , \29861 , \29863 );
not \U$29522 ( \29865 , \29777 );
not \U$29523 ( \29866 , \29865 );
not \U$29524 ( \29867 , \29766 );
or \U$29525 ( \29868 , \29866 , \29867 );
nand \U$29526 ( \29869 , \29868 , \29762 );
nand \U$29527 ( \29870 , \29751 , \29777 );
nand \U$29528 ( \29871 , \29869 , \29870 );
xor \U$29529 ( \29872 , \29864 , \29871 );
or \U$29530 ( \29873 , \29730 , \29714 );
not \U$29531 ( \29874 , \29719 );
nand \U$29532 ( \29875 , \29873 , \29874 );
nand \U$29533 ( \29876 , \29730 , \29714 );
nand \U$29534 ( \29877 , \29875 , \29876 );
not \U$29535 ( \29878 , \29877 );
and \U$29536 ( \29879 , \29872 , \29878 );
not \U$29537 ( \29880 , \29872 );
and \U$29538 ( \29881 , \29880 , \29877 );
nor \U$29539 ( \29882 , \29879 , \29881 );
not \U$29540 ( \29883 , \29882 );
not \U$29541 ( \29884 , \29883 );
or \U$29542 ( \29885 , \29858 , \29884 );
not \U$29543 ( \29886 , \29857 );
not \U$29544 ( \29887 , \29886 );
not \U$29545 ( \29888 , \29882 );
or \U$29546 ( \29889 , \29887 , \29888 );
and \U$29547 ( \29890 , \17506 , \1077 );
not \U$29548 ( \29891 , \998 );
not \U$29549 ( \29892 , RIbb2f070_13);
not \U$29550 ( \29893 , \16819 );
or \U$29551 ( \29894 , \29892 , \29893 );
nand \U$29552 ( \29895 , \17529 , \906 );
nand \U$29553 ( \29896 , \29894 , \29895 );
not \U$29554 ( \29897 , \29896 );
or \U$29555 ( \29898 , \29891 , \29897 );
nand \U$29556 ( \29899 , \29684 , \915 );
nand \U$29557 ( \29900 , \29898 , \29899 );
xor \U$29558 ( \29901 , \29890 , \29900 );
not \U$29559 ( \29902 , \1517 );
and \U$29560 ( \29903 , RIbb2ef80_15, \16554 );
not \U$29561 ( \29904 , RIbb2ef80_15);
and \U$29562 ( \29905 , \29904 , \29271 );
or \U$29563 ( \29906 , \29903 , \29905 );
not \U$29564 ( \29907 , \29906 );
or \U$29565 ( \29908 , \29902 , \29907 );
nand \U$29566 ( \29909 , \29698 , \1444 );
nand \U$29567 ( \29910 , \29908 , \29909 );
xor \U$29568 ( \29911 , \29901 , \29910 );
not \U$29569 ( \29912 , \2963 );
and \U$29570 ( \29913 , RIbb2ead0_25, \12348 );
not \U$29571 ( \29914 , RIbb2ead0_25);
and \U$29572 ( \29915 , \29914 , \12347 );
or \U$29573 ( \29916 , \29913 , \29915 );
not \U$29574 ( \29917 , \29916 );
or \U$29575 ( \29918 , \29912 , \29917 );
nand \U$29576 ( \29919 , \29589 , \2980 );
nand \U$29577 ( \29920 , \29918 , \29919 );
xor \U$29578 ( \29921 , \29911 , \29920 );
not \U$29579 ( \29922 , \3465 );
and \U$29580 ( \29923 , \12174 , \6065 );
not \U$29581 ( \29924 , \12174 );
and \U$29582 ( \29925 , \29924 , RIbb2e9e0_27);
or \U$29583 ( \29926 , \29923 , \29925 );
not \U$29584 ( \29927 , \29926 );
or \U$29585 ( \29928 , \29922 , \29927 );
nand \U$29586 ( \29929 , \29388 , \3445 );
nand \U$29587 ( \29930 , \29928 , \29929 );
xor \U$29588 ( \29931 , \29921 , \29930 );
not \U$29589 ( \29932 , \3406 );
not \U$29590 ( \29933 , \29580 );
or \U$29591 ( \29934 , \29932 , \29933 );
not \U$29592 ( \29935 , RIbb2ebc0_23);
not \U$29593 ( \29936 , \13986 );
or \U$29594 ( \29937 , \29935 , \29936 );
not \U$29595 ( \29938 , \18552 );
nand \U$29596 ( \29939 , \29938 , \3388 );
nand \U$29597 ( \29940 , \29937 , \29939 );
nand \U$29598 ( \29941 , \29940 , \3382 );
nand \U$29599 ( \29942 , \29934 , \29941 );
not \U$29600 ( \29943 , \2077 );
not \U$29601 ( \29944 , \29604 );
or \U$29602 ( \29945 , \29943 , \29944 );
not \U$29603 ( \29946 , \7768 );
and \U$29604 ( \29947 , \20577 , RIbb2ecb0_21);
not \U$29605 ( \29948 , \20577 );
and \U$29606 ( \29949 , \29948 , \2249 );
or \U$29607 ( \29950 , \29947 , \29949 );
nand \U$29608 ( \29951 , \29946 , \29950 );
nand \U$29609 ( \29952 , \29945 , \29951 );
not \U$29610 ( \29953 , \29952 );
xor \U$29611 ( \29954 , \29942 , \29953 );
not \U$29612 ( \29955 , \3887 );
not \U$29613 ( \29956 , \29794 );
or \U$29614 ( \29957 , \29955 , \29956 );
not \U$29615 ( \29958 , RIbb2e710_33);
not \U$29616 ( \29959 , \9277 );
not \U$29617 ( \29960 , \29959 );
or \U$29618 ( \29961 , \29958 , \29960 );
nand \U$29619 ( \29962 , \9277 , \2935 );
nand \U$29620 ( \29963 , \29961 , \29962 );
nand \U$29621 ( \29964 , \29963 , \4075 );
nand \U$29622 ( \29965 , \29957 , \29964 );
xnor \U$29623 ( \29966 , \29954 , \29965 );
xor \U$29624 ( \29967 , \29931 , \29966 );
xor \U$29625 ( \29968 , \29473 , \29483 );
and \U$29626 ( \29969 , \29968 , \29494 );
and \U$29627 ( \29970 , \29473 , \29483 );
or \U$29628 ( \29971 , \29969 , \29970 );
xor \U$29629 ( \29972 , \29967 , \29971 );
nand \U$29630 ( \29973 , \29889 , \29972 );
nand \U$29631 ( \29974 , \29885 , \29973 );
not \U$29632 ( \29975 , \29974 );
xor \U$29633 ( \29976 , \29693 , \29702 );
and \U$29634 ( \29977 , \29976 , \29713 );
and \U$29635 ( \29978 , \29693 , \29702 );
or \U$29636 ( \29979 , \29977 , \29978 );
not \U$29637 ( \29980 , \4712 );
not \U$29638 ( \29981 , \29469 );
or \U$29639 ( \29982 , \29980 , \29981 );
not \U$29640 ( \29983 , RIbb2e620_35);
not \U$29641 ( \29984 , \20692 );
or \U$29642 ( \29985 , \29983 , \29984 );
nand \U$29643 ( \29986 , \8318 , \6002 );
nand \U$29644 ( \29987 , \29985 , \29986 );
nand \U$29645 ( \29988 , \29987 , \5845 );
nand \U$29646 ( \29989 , \29982 , \29988 );
xor \U$29647 ( \29990 , \29979 , \29989 );
not \U$29648 ( \29991 , RIbb2d888_64);
not \U$29649 ( \29992 , RIbb2d900_63);
not \U$29650 ( \29993 , \7423 );
or \U$29651 ( \29994 , \29992 , \29993 );
nand \U$29652 ( \29995 , \24399 , \17262 );
nand \U$29653 ( \29996 , \29994 , \29995 );
not \U$29654 ( \29997 , \29996 );
or \U$29655 ( \29998 , \29991 , \29997 );
nand \U$29656 ( \29999 , \29481 , \17275 );
nand \U$29657 ( \30000 , \29998 , \29999 );
and \U$29658 ( \30001 , \29990 , \30000 );
and \U$29659 ( \30002 , \29979 , \29989 );
or \U$29660 ( \30003 , \30001 , \30002 );
not \U$29661 ( \30004 , \15738 );
not \U$29662 ( \30005 , RIbb2dbd0_57);
not \U$29663 ( \30006 , \22684 );
or \U$29664 ( \30007 , \30005 , \30006 );
nand \U$29665 ( \30008 , \1419 , \16671 );
nand \U$29666 ( \30009 , \30007 , \30008 );
not \U$29667 ( \30010 , \30009 );
or \U$29668 ( \30011 , \30004 , \30010 );
not \U$29669 ( \30012 , RIbb2dbd0_57);
not \U$29670 ( \30013 , \19733 );
or \U$29671 ( \30014 , \30012 , \30013 );
nand \U$29672 ( \30015 , \1337 , \15741 );
nand \U$29673 ( \30016 , \30014 , \30015 );
nand \U$29674 ( \30017 , \30016 , \15746 );
nand \U$29675 ( \30018 , \30011 , \30017 );
not \U$29676 ( \30019 , \11176 );
not \U$29677 ( \30020 , \11959 );
not \U$29678 ( \30021 , \4020 );
or \U$29679 ( \30022 , \30020 , \30021 );
or \U$29680 ( \30023 , \3022 , \12971 );
nand \U$29681 ( \30024 , \30022 , \30023 );
not \U$29682 ( \30025 , \30024 );
or \U$29683 ( \30026 , \30019 , \30025 );
not \U$29684 ( \30027 , RIbb2e080_47);
not \U$29685 ( \30028 , \21490 );
or \U$29686 ( \30029 , \30027 , \30028 );
nand \U$29687 ( \30030 , \3653 , \10113 );
nand \U$29688 ( \30031 , \30029 , \30030 );
nand \U$29689 ( \30032 , \30031 , \11177 );
nand \U$29690 ( \30033 , \30026 , \30032 );
xor \U$29691 ( \30034 , \30018 , \30033 );
not \U$29692 ( \30035 , \10599 );
not \U$29693 ( \30036 , RIbb2e170_45);
not \U$29694 ( \30037 , \15605 );
or \U$29695 ( \30038 , \30036 , \30037 );
nand \U$29696 ( \30039 , \13732 , \11065 );
nand \U$29697 ( \30040 , \30038 , \30039 );
not \U$29698 ( \30041 , \30040 );
or \U$29699 ( \30042 , \30035 , \30041 );
not \U$29700 ( \30043 , RIbb2e170_45);
not \U$29701 ( \30044 , \17910 );
or \U$29702 ( \30045 , \30043 , \30044 );
nand \U$29703 ( \30046 , \3044 , \12003 );
nand \U$29704 ( \30047 , \30045 , \30046 );
nand \U$29705 ( \30048 , \30047 , \10119 );
nand \U$29706 ( \30049 , \30042 , \30048 );
xor \U$29707 ( \30050 , \30034 , \30049 );
xor \U$29708 ( \30051 , \30003 , \30050 );
and \U$29709 ( \30052 , \29678 , \29692 );
not \U$29710 ( \30053 , \831 );
not \U$29711 ( \30054 , \29371 );
or \U$29712 ( \30055 , \30053 , \30054 );
not \U$29713 ( \30056 , RIbb2ee90_17);
not \U$29714 ( \30057 , \16746 );
or \U$29715 ( \30058 , \30056 , \30057 );
nand \U$29716 ( \30059 , \24010 , \3057 );
nand \U$29717 ( \30060 , \30058 , \30059 );
nand \U$29718 ( \30061 , \30060 , \836 );
nand \U$29719 ( \30062 , \30055 , \30061 );
xor \U$29720 ( \30063 , \30052 , \30062 );
not \U$29721 ( \30064 , \854 );
and \U$29722 ( \30065 , \1776 , \16567 );
not \U$29723 ( \30066 , \1776 );
and \U$29724 ( \30067 , \30066 , \23098 );
nor \U$29725 ( \30068 , \30065 , \30067 );
not \U$29726 ( \30069 , \30068 );
or \U$29727 ( \30070 , \30064 , \30069 );
nand \U$29728 ( \30071 , \29709 , \853 );
nand \U$29729 ( \30072 , \30070 , \30071 );
and \U$29730 ( \30073 , \30063 , \30072 );
and \U$29731 ( \30074 , \30052 , \30062 );
or \U$29732 ( \30075 , \30073 , \30074 );
not \U$29733 ( \30076 , \16541 );
not \U$29734 ( \30077 , RIbb2d9f0_61);
not \U$29735 ( \30078 , \12037 );
or \U$29736 ( \30079 , \30077 , \30078 );
nand \U$29737 ( \30080 , \12036 , \19746 );
nand \U$29738 ( \30081 , \30079 , \30080 );
not \U$29739 ( \30082 , \30081 );
or \U$29740 ( \30083 , \30076 , \30082 );
not \U$29741 ( \30084 , RIbb2d9f0_61);
not \U$29742 ( \30085 , \13707 );
or \U$29743 ( \30086 , \30084 , \30085 );
nand \U$29744 ( \30087 , \1111 , \16254 );
nand \U$29745 ( \30088 , \30086 , \30087 );
nand \U$29746 ( \30089 , \30088 , \16533 );
nand \U$29747 ( \30090 , \30083 , \30089 );
xor \U$29748 ( \30091 , \30075 , \30090 );
not \U$29749 ( \30092 , \12167 );
not \U$29750 ( \30093 , RIbb2df90_49);
not \U$29751 ( \30094 , \6172 );
or \U$29752 ( \30095 , \30093 , \30094 );
nand \U$29753 ( \30096 , \26749 , \12278 );
nand \U$29754 ( \30097 , \30095 , \30096 );
not \U$29755 ( \30098 , \30097 );
or \U$29756 ( \30099 , \30092 , \30098 );
not \U$29757 ( \30100 , RIbb2df90_49);
not \U$29758 ( \30101 , \3200 );
or \U$29759 ( \30102 , \30100 , \30101 );
nand \U$29760 ( \30103 , \3201 , \12278 );
nand \U$29761 ( \30104 , \30102 , \30103 );
nand \U$29762 ( \30105 , \30104 , \16427 );
nand \U$29763 ( \30106 , \30099 , \30105 );
xor \U$29764 ( \30107 , \30091 , \30106 );
xor \U$29765 ( \30108 , \30051 , \30107 );
not \U$29766 ( \30109 , \3146 );
not \U$29767 ( \30110 , \21882 );
and \U$29768 ( \30111 , \30109 , \30110 );
not \U$29769 ( \30112 , \15398 );
and \U$29770 ( \30113 , \30112 , \21882 );
nor \U$29771 ( \30114 , \30111 , \30113 );
not \U$29772 ( \30115 , \30114 );
not \U$29773 ( \30116 , \25687 );
and \U$29774 ( \30117 , \30115 , \30116 );
and \U$29775 ( \30118 , \29408 , \12774 );
nor \U$29776 ( \30119 , \30117 , \30118 );
not \U$29777 ( \30120 , \30119 );
not \U$29778 ( \30121 , \30120 );
not \U$29779 ( \30122 , \29594 );
not \U$29780 ( \30123 , \30122 );
not \U$29781 ( \30124 , \29582 );
or \U$29782 ( \30125 , \30123 , \30124 );
or \U$29783 ( \30126 , \29582 , \30122 );
nand \U$29784 ( \30127 , \30126 , \29609 );
nand \U$29785 ( \30128 , \30125 , \30127 );
not \U$29786 ( \30129 , \30128 );
or \U$29787 ( \30130 , \30121 , \30129 );
not \U$29788 ( \30131 , \30128 );
not \U$29789 ( \30132 , \30131 );
not \U$29790 ( \30133 , \30119 );
or \U$29791 ( \30134 , \30132 , \30133 );
xor \U$29792 ( \30135 , \29375 , \29379 );
and \U$29793 ( \30136 , \30135 , \29390 );
and \U$29794 ( \30137 , \29375 , \29379 );
or \U$29795 ( \30138 , \30136 , \30137 );
nand \U$29796 ( \30139 , \30134 , \30138 );
nand \U$29797 ( \30140 , \30130 , \30139 );
not \U$29798 ( \30141 , \17275 );
not \U$29799 ( \30142 , \29996 );
or \U$29800 ( \30143 , \30141 , \30142 );
not \U$29801 ( \30144 , RIbb2d900_63);
not \U$29802 ( \30145 , \3238 );
or \U$29803 ( \30146 , \30144 , \30145 );
nand \U$29804 ( \30147 , \1642 , \17262 );
nand \U$29805 ( \30148 , \30146 , \30147 );
nand \U$29806 ( \30149 , \30148 , RIbb2d888_64);
nand \U$29807 ( \30150 , \30143 , \30149 );
not \U$29808 ( \30151 , \16271 );
and \U$29809 ( \30152 , RIbb2dae0_59, \4339 );
not \U$29810 ( \30153 , RIbb2dae0_59);
and \U$29811 ( \30154 , \30153 , \1386 );
or \U$29812 ( \30155 , \30152 , \30154 );
not \U$29813 ( \30156 , \30155 );
or \U$29814 ( \30157 , \30151 , \30156 );
not \U$29815 ( \30158 , \3990 );
xor \U$29816 ( \30159 , RIbb2dae0_59, \30158 );
nand \U$29817 ( \30160 , \30159 , \17470 );
nand \U$29818 ( \30161 , \30157 , \30160 );
xor \U$29819 ( \30162 , \30150 , \30161 );
not \U$29820 ( \30163 , \12692 );
and \U$29821 ( \30164 , RIbb2dea0_51, \13414 );
not \U$29822 ( \30165 , RIbb2dea0_51);
and \U$29823 ( \30166 , \30165 , \3167 );
or \U$29824 ( \30167 , \30164 , \30166 );
not \U$29825 ( \30168 , \30167 );
or \U$29826 ( \30169 , \30163 , \30168 );
not \U$29827 ( \30170 , \30114 );
nand \U$29828 ( \30171 , \30170 , \14067 );
nand \U$29829 ( \30172 , \30169 , \30171 );
xor \U$29830 ( \30173 , \30162 , \30172 );
xor \U$29831 ( \30174 , \30140 , \30173 );
not \U$29832 ( \30175 , \9099 );
not \U$29833 ( \30176 , RIbb2e260_43);
not \U$29834 ( \30177 , \3090 );
or \U$29835 ( \30178 , \30176 , \30177 );
nand \U$29836 ( \30179 , \3089 , \8347 );
nand \U$29837 ( \30180 , \30178 , \30179 );
not \U$29838 ( \30181 , \30180 );
or \U$29839 ( \30182 , \30175 , \30181 );
not \U$29840 ( \30183 , RIbb2e260_43);
not \U$29841 ( \30184 , \13552 );
or \U$29842 ( \30185 , \30183 , \30184 );
nand \U$29843 ( \30186 , \13551 , \8347 );
nand \U$29844 ( \30187 , \30185 , \30186 );
nand \U$29845 ( \30188 , \30187 , \9098 );
nand \U$29846 ( \30189 , \30182 , \30188 );
not \U$29847 ( \30190 , \14920 );
not \U$29848 ( \30191 , RIbb2ddb0_53);
not \U$29849 ( \30192 , \20951 );
or \U$29850 ( \30193 , \30191 , \30192 );
not \U$29851 ( \30194 , \3516 );
nand \U$29852 ( \30195 , \30194 , \12681 );
nand \U$29853 ( \30196 , \30193 , \30195 );
not \U$29854 ( \30197 , \30196 );
or \U$29855 ( \30198 , \30190 , \30197 );
not \U$29856 ( \30199 , RIbb2ddb0_53);
not \U$29857 ( \30200 , \3319 );
or \U$29858 ( \30201 , \30199 , \30200 );
nand \U$29859 ( \30202 , \2222 , \13463 );
nand \U$29860 ( \30203 , \30201 , \30202 );
nand \U$29861 ( \30204 , \30203 , \14930 );
nand \U$29862 ( \30205 , \30198 , \30204 );
xor \U$29863 ( \30206 , \30189 , \30205 );
not \U$29864 ( \30207 , \14613 );
not \U$29865 ( \30208 , RIbb2dcc0_55);
not \U$29866 ( \30209 , \3309 );
not \U$29867 ( \30210 , \30209 );
or \U$29868 ( \30211 , \30208 , \30210 );
not \U$29869 ( \30212 , RIbb2dcc0_55);
nand \U$29870 ( \30213 , \30212 , \2114 );
nand \U$29871 ( \30214 , \30211 , \30213 );
not \U$29872 ( \30215 , \30214 );
or \U$29873 ( \30216 , \30207 , \30215 );
and \U$29874 ( \30217 , RIbb2dcc0_55, \20325 );
not \U$29875 ( \30218 , RIbb2dcc0_55);
and \U$29876 ( \30219 , \30218 , \1851 );
or \U$29877 ( \30220 , \30217 , \30219 );
nand \U$29878 ( \30221 , \30220 , \15181 );
nand \U$29879 ( \30222 , \30216 , \30221 );
xor \U$29880 ( \30223 , \30206 , \30222 );
xor \U$29881 ( \30224 , \30174 , \30223 );
not \U$29882 ( \30225 , \30224 );
and \U$29883 ( \30226 , \30108 , \30225 );
not \U$29884 ( \30227 , \30108 );
and \U$29885 ( \30228 , \30227 , \30224 );
nor \U$29886 ( \30229 , \30226 , \30228 );
not \U$29887 ( \30230 , \30229 );
or \U$29888 ( \30231 , \29975 , \30230 );
or \U$29889 ( \30232 , \30229 , \29974 );
nand \U$29890 ( \30233 , \30231 , \30232 );
xor \U$29891 ( \30234 , \30138 , \30128 );
xor \U$29892 ( \30235 , \30234 , \30119 );
not \U$29893 ( \30236 , \30235 );
not \U$29894 ( \30237 , \30236 );
xor \U$29895 ( \30238 , \29660 , \29667 );
and \U$29896 ( \30239 , \30238 , \29672 );
and \U$29897 ( \30240 , \29660 , \29667 );
or \U$29898 ( \30241 , \30239 , \30240 );
not \U$29899 ( \30242 , \30241 );
not \U$29900 ( \30243 , \30242 );
or \U$29901 ( \30244 , \30237 , \30243 );
nand \U$29902 ( \30245 , \30241 , \30235 );
nand \U$29903 ( \30246 , \30244 , \30245 );
xor \U$29904 ( \30247 , \29731 , \29735 );
and \U$29905 ( \30248 , \30247 , \29740 );
and \U$29906 ( \30249 , \29731 , \29735 );
or \U$29907 ( \30250 , \30248 , \30249 );
xnor \U$29908 ( \30251 , \30246 , \30250 );
not \U$29909 ( \30252 , \30251 );
not \U$29910 ( \30253 , \30252 );
xor \U$29911 ( \30254 , \29857 , \29972 );
xnor \U$29912 ( \30255 , \30254 , \29883 );
not \U$29913 ( \30256 , \30255 );
not \U$29914 ( \30257 , \30256 );
or \U$29915 ( \30258 , \30253 , \30257 );
not \U$29916 ( \30259 , \30255 );
not \U$29917 ( \30260 , \30251 );
or \U$29918 ( \30261 , \30259 , \30260 );
xor \U$29919 ( \30262 , \29627 , \29636 );
and \U$29920 ( \30263 , \30262 , \29641 );
and \U$29921 ( \30264 , \29627 , \29636 );
or \U$29922 ( \30265 , \30263 , \30264 );
nand \U$29923 ( \30266 , \30261 , \30265 );
nand \U$29924 ( \30267 , \30258 , \30266 );
xor \U$29925 ( \30268 , \30233 , \30267 );
not \U$29926 ( \30269 , \30235 );
not \U$29927 ( \30270 , \30242 );
or \U$29928 ( \30271 , \30269 , \30270 );
nand \U$29929 ( \30272 , \30271 , \30250 );
not \U$29930 ( \30273 , \30242 );
nand \U$29931 ( \30274 , \30273 , \30236 );
nand \U$29932 ( \30275 , \30272 , \30274 );
not \U$29933 ( \30276 , \1517 );
and \U$29934 ( \30277 , RIbb2ef80_15, \27577 );
not \U$29935 ( \30278 , RIbb2ef80_15);
and \U$29936 ( \30279 , \30278 , \16829 );
or \U$29937 ( \30280 , \30277 , \30279 );
not \U$29938 ( \30281 , \30280 );
or \U$29939 ( \30282 , \30276 , \30281 );
nand \U$29940 ( \30283 , \29906 , \1444 );
nand \U$29941 ( \30284 , \30282 , \30283 );
xor \U$29942 ( \30285 , \29890 , \29900 );
and \U$29943 ( \30286 , \30285 , \29910 );
and \U$29944 ( \30287 , \29890 , \29900 );
or \U$29945 ( \30288 , \30286 , \30287 );
xor \U$29946 ( \30289 , \30284 , \30288 );
not \U$29947 ( \30290 , \3406 );
not \U$29948 ( \30291 , \29940 );
or \U$29949 ( \30292 , \30290 , \30291 );
not \U$29950 ( \30293 , RIbb2ebc0_23);
not \U$29951 ( \30294 , \14624 );
or \U$29952 ( \30295 , \30293 , \30294 );
nand \U$29953 ( \30296 , \13210 , \3388 );
nand \U$29954 ( \30297 , \30295 , \30296 );
nand \U$29955 ( \30298 , \30297 , \3382 );
nand \U$29956 ( \30299 , \30292 , \30298 );
xor \U$29957 ( \30300 , \30289 , \30299 );
xor \U$29958 ( \30301 , \29911 , \29920 );
and \U$29959 ( \30302 , \30301 , \29930 );
and \U$29960 ( \30303 , \29911 , \29920 );
or \U$29961 ( \30304 , \30302 , \30303 );
xor \U$29962 ( \30305 , \30300 , \30304 );
nor \U$29963 ( \30306 , \29965 , \29942 );
or \U$29964 ( \30307 , \30306 , \29953 );
nand \U$29965 ( \30308 , \29965 , \29942 );
nand \U$29966 ( \30309 , \30307 , \30308 );
xor \U$29967 ( \30310 , \30305 , \30309 );
nor \U$29968 ( \30311 , \29871 , \29864 );
or \U$29969 ( \30312 , \29878 , \30311 );
nand \U$29970 ( \30313 , \29864 , \29871 );
nand \U$29971 ( \30314 , \30312 , \30313 );
xor \U$29972 ( \30315 , \30310 , \30314 );
not \U$29973 ( \30316 , \854 );
not \U$29974 ( \30317 , RIbb2eda0_19);
not \U$29975 ( \30318 , \15469 );
or \U$29976 ( \30319 , \30317 , \30318 );
nand \U$29977 ( \30320 , \15030 , \1776 );
nand \U$29978 ( \30321 , \30319 , \30320 );
not \U$29979 ( \30322 , \30321 );
or \U$29980 ( \30323 , \30316 , \30322 );
nand \U$29981 ( \30324 , \853 , \30068 );
nand \U$29982 ( \30325 , \30323 , \30324 );
not \U$29983 ( \30326 , \2980 );
not \U$29984 ( \30327 , \29916 );
or \U$29985 ( \30328 , \30326 , \30327 );
and \U$29986 ( \30329 , RIbb2ead0_25, \17663 );
not \U$29987 ( \30330 , RIbb2ead0_25);
and \U$29988 ( \30331 , \30330 , \12932 );
or \U$29989 ( \30332 , \30329 , \30331 );
nand \U$29990 ( \30333 , \30332 , \2963 );
nand \U$29991 ( \30334 , \30328 , \30333 );
xor \U$29992 ( \30335 , \30325 , \30334 );
not \U$29993 ( \30336 , \2077 );
not \U$29994 ( \30337 , \29950 );
or \U$29995 ( \30338 , \30336 , \30337 );
not \U$29996 ( \30339 , RIbb2ecb0_21);
not \U$29997 ( \30340 , \13978 );
or \U$29998 ( \30341 , \30339 , \30340 );
nand \U$29999 ( \30342 , \16320 , \5481 );
nand \U$30000 ( \30343 , \30341 , \30342 );
nand \U$30001 ( \30344 , \30343 , \2078 );
nand \U$30002 ( \30345 , \30338 , \30344 );
xor \U$30003 ( \30346 , \30335 , \30345 );
not \U$30004 ( \30347 , \2940 );
not \U$30005 ( \30348 , \29807 );
or \U$30006 ( \30349 , \30347 , \30348 );
not \U$30007 ( \30350 , RIbb2e800_31);
not \U$30008 ( \30351 , \15105 );
or \U$30009 ( \30352 , \30350 , \30351 );
nand \U$30010 ( \30353 , \2917 , \10300 );
nand \U$30011 ( \30354 , \30352 , \30353 );
nand \U$30012 ( \30355 , \30354 , \3613 );
nand \U$30013 ( \30356 , \30349 , \30355 );
not \U$30014 ( \30357 , \2921 );
not \U$30015 ( \30358 , \29784 );
or \U$30016 ( \30359 , \30357 , \30358 );
not \U$30017 ( \30360 , RIbb2e8f0_29);
not \U$30018 ( \30361 , \11143 );
or \U$30019 ( \30362 , \30360 , \30361 );
nand \U$30020 ( \30363 , \11142 , \2949 );
nand \U$30021 ( \30364 , \30362 , \30363 );
nand \U$30022 ( \30365 , \30364 , \2925 );
nand \U$30023 ( \30366 , \30359 , \30365 );
xor \U$30024 ( \30367 , \30356 , \30366 );
not \U$30025 ( \30368 , \9099 );
not \U$30026 ( \30369 , \30187 );
or \U$30027 ( \30370 , \30368 , \30369 );
nand \U$30028 ( \30371 , \29760 , \9098 );
nand \U$30029 ( \30372 , \30370 , \30371 );
and \U$30030 ( \30373 , \30367 , \30372 );
and \U$30031 ( \30374 , \30356 , \30366 );
or \U$30032 ( \30375 , \30373 , \30374 );
xor \U$30033 ( \30376 , \30346 , \30375 );
not \U$30034 ( \30377 , \7103 );
not \U$30035 ( \30378 , \29747 );
or \U$30036 ( \30379 , \30377 , \30378 );
xor \U$30037 ( \30380 , RIbb2e440_39, \5954 );
nand \U$30038 ( \30381 , \30380 , \8450 );
nand \U$30039 ( \30382 , \30379 , \30381 );
not \U$30040 ( \30383 , \8353 );
not \U$30041 ( \30384 , RIbb2e350_41);
not \U$30042 ( \30385 , \9021 );
or \U$30043 ( \30386 , \30384 , \30385 );
not \U$30044 ( \30387 , \10555 );
nand \U$30045 ( \30388 , \30387 , \9402 );
nand \U$30046 ( \30389 , \30386 , \30388 );
not \U$30047 ( \30390 , \30389 );
or \U$30048 ( \30391 , \30383 , \30390 );
nand \U$30049 ( \30392 , \29775 , \8362 );
nand \U$30050 ( \30393 , \30391 , \30392 );
xor \U$30051 ( \30394 , \30382 , \30393 );
not \U$30052 ( \30395 , \6251 );
not \U$30053 ( \30396 , \29726 );
or \U$30054 ( \30397 , \30395 , \30396 );
not \U$30055 ( \30398 , RIbb2e530_37);
not \U$30056 ( \30399 , \12790 );
or \U$30057 ( \30400 , \30398 , \30399 );
nand \U$30058 ( \30401 , \25844 , \6246 );
nand \U$30059 ( \30402 , \30400 , \30401 );
nand \U$30060 ( \30403 , \30402 , \6242 );
nand \U$30061 ( \30404 , \30397 , \30403 );
and \U$30062 ( \30405 , \30394 , \30404 );
and \U$30063 ( \30406 , \30382 , \30393 );
or \U$30064 ( \30407 , \30405 , \30406 );
xor \U$30065 ( \30408 , \30376 , \30407 );
xor \U$30066 ( \30409 , \30315 , \30408 );
xor \U$30067 ( \30410 , \30275 , \30409 );
not \U$30068 ( \30411 , \29966 );
not \U$30069 ( \30412 , \29971 );
or \U$30070 ( \30413 , \30411 , \30412 );
or \U$30071 ( \30414 , \29971 , \29966 );
nand \U$30072 ( \30415 , \30414 , \29931 );
nand \U$30073 ( \30416 , \30413 , \30415 );
xor \U$30074 ( \30417 , \29979 , \29989 );
xor \U$30075 ( \30418 , \30417 , \30000 );
not \U$30076 ( \30419 , \29536 );
not \U$30077 ( \30420 , \29557 );
or \U$30078 ( \30421 , \30419 , \30420 );
or \U$30079 ( \30422 , \29557 , \29536 );
nand \U$30080 ( \30423 , \30422 , \29546 );
nand \U$30081 ( \30424 , \30421 , \30423 );
xor \U$30082 ( \30425 , \30418 , \30424 );
xor \U$30083 ( \30426 , \29505 , \29514 );
and \U$30084 ( \30427 , \30426 , \29524 );
and \U$30085 ( \30428 , \29505 , \29514 );
or \U$30086 ( \30429 , \30427 , \30428 );
and \U$30087 ( \30430 , \30425 , \30429 );
and \U$30088 ( \30431 , \30418 , \30424 );
or \U$30089 ( \30432 , \30430 , \30431 );
xor \U$30090 ( \30433 , \30416 , \30432 );
not \U$30091 ( \30434 , \14613 );
not \U$30092 ( \30435 , \29520 );
or \U$30093 ( \30436 , \30434 , \30435 );
nand \U$30094 ( \30437 , \30214 , \15181 );
nand \U$30095 ( \30438 , \30436 , \30437 );
not \U$30096 ( \30439 , \30438 );
not \U$30097 ( \30440 , \10599 );
not \U$30098 ( \30441 , \29542 );
or \U$30099 ( \30442 , \30440 , \30441 );
nand \U$30100 ( \30443 , \30040 , \10119 );
nand \U$30101 ( \30444 , \30442 , \30443 );
not \U$30102 ( \30445 , \30444 );
or \U$30103 ( \30446 , \30439 , \30445 );
or \U$30104 ( \30447 , \30444 , \30438 );
not \U$30105 ( \30448 , \16533 );
not \U$30106 ( \30449 , \30081 );
or \U$30107 ( \30450 , \30448 , \30449 );
nand \U$30108 ( \30451 , \29503 , \16541 );
nand \U$30109 ( \30452 , \30450 , \30451 );
nand \U$30110 ( \30453 , \30447 , \30452 );
nand \U$30111 ( \30454 , \30446 , \30453 );
xor \U$30112 ( \30455 , \30052 , \30062 );
xor \U$30113 ( \30456 , \30455 , \30072 );
not \U$30114 ( \30457 , \17563 );
not \U$30115 ( \30458 , \29510 );
or \U$30116 ( \30459 , \30457 , \30458 );
nand \U$30117 ( \30460 , \30196 , \15688 );
nand \U$30118 ( \30461 , \30459 , \30460 );
xor \U$30119 ( \30462 , \30456 , \30461 );
not \U$30120 ( \30463 , \16271 );
not \U$30121 ( \30464 , \29396 );
or \U$30122 ( \30465 , \30463 , \30464 );
nand \U$30123 ( \30466 , \30155 , \17470 );
nand \U$30124 ( \30467 , \30465 , \30466 );
and \U$30125 ( \30468 , \30462 , \30467 );
and \U$30126 ( \30469 , \30456 , \30461 );
or \U$30127 ( \30470 , \30468 , \30469 );
xor \U$30128 ( \30471 , \30454 , \30470 );
not \U$30129 ( \30472 , \11176 );
not \U$30130 ( \30473 , \29555 );
or \U$30131 ( \30474 , \30472 , \30473 );
nand \U$30132 ( \30475 , \30024 , \12965 );
nand \U$30133 ( \30476 , \30474 , \30475 );
not \U$30134 ( \30477 , \16674 );
not \U$30135 ( \30478 , \29534 );
or \U$30136 ( \30479 , \30477 , \30478 );
nand \U$30137 ( \30480 , \30016 , \17100 );
nand \U$30138 ( \30481 , \30479 , \30480 );
nor \U$30139 ( \30482 , \30476 , \30481 );
not \U$30140 ( \30483 , \12167 );
not \U$30141 ( \30484 , \29492 );
or \U$30142 ( \30485 , \30483 , \30484 );
nand \U$30143 ( \30486 , \30097 , \14752 );
nand \U$30144 ( \30487 , \30485 , \30486 );
not \U$30145 ( \30488 , \30487 );
or \U$30146 ( \30489 , \30482 , \30488 );
nand \U$30147 ( \30490 , \30481 , \30476 );
nand \U$30148 ( \30491 , \30489 , \30490 );
xor \U$30149 ( \30492 , \30471 , \30491 );
xor \U$30150 ( \30493 , \30433 , \30492 );
xor \U$30151 ( \30494 , \30410 , \30493 );
xor \U$30152 ( \30495 , \30268 , \30494 );
not \U$30153 ( \30496 , \29642 );
not \U$30154 ( \30497 , \30496 );
not \U$30155 ( \30498 , \29824 );
or \U$30156 ( \30499 , \30497 , \30498 );
not \U$30157 ( \30500 , \29654 );
nand \U$30158 ( \30501 , \30499 , \30500 );
not \U$30159 ( \30502 , \29824 );
nand \U$30160 ( \30503 , \30502 , \29642 );
nand \U$30161 ( \30504 , \30501 , \30503 );
not \U$30162 ( \30505 , \29823 );
not \U$30163 ( \30506 , \29673 );
or \U$30164 ( \30507 , \30505 , \30506 );
not \U$30165 ( \30508 , \29673 );
not \U$30166 ( \30509 , \30508 );
not \U$30167 ( \30510 , \29822 );
or \U$30168 ( \30511 , \30509 , \30510 );
nand \U$30169 ( \30512 , \30511 , \29741 );
nand \U$30170 ( \30513 , \30507 , \30512 );
not \U$30171 ( \30514 , \29560 );
not \U$30172 ( \30515 , \29457 );
or \U$30173 ( \30516 , \30514 , \30515 );
not \U$30174 ( \30517 , \29457 );
not \U$30175 ( \30518 , \30517 );
not \U$30176 ( \30519 , \29559 );
or \U$30177 ( \30520 , \30518 , \30519 );
nand \U$30178 ( \30521 , \30520 , \29461 );
nand \U$30179 ( \30522 , \30516 , \30521 );
xor \U$30180 ( \30523 , \30513 , \30522 );
not \U$30181 ( \30524 , \29810 );
or \U$30182 ( \30525 , \30524 , \29817 );
nand \U$30183 ( \30526 , \30525 , \29778 );
nand \U$30184 ( \30527 , \29817 , \30524 );
nand \U$30185 ( \30528 , \30526 , \30527 );
not \U$30186 ( \30529 , \29495 );
not \U$30187 ( \30530 , \29525 );
or \U$30188 ( \30531 , \30529 , \30530 );
or \U$30189 ( \30532 , \29525 , \29495 );
nand \U$30190 ( \30533 , \30532 , \29558 );
nand \U$30191 ( \30534 , \30531 , \30533 );
xor \U$30192 ( \30535 , \30528 , \30534 );
xor \U$30193 ( \30536 , \30382 , \30393 );
xor \U$30194 ( \30537 , \30536 , \30404 );
xor \U$30195 ( \30538 , \30356 , \30366 );
xor \U$30196 ( \30539 , \30538 , \30372 );
not \U$30197 ( \30540 , \30539 );
and \U$30198 ( \30541 , \30537 , \30540 );
not \U$30199 ( \30542 , \30537 );
and \U$30200 ( \30543 , \30542 , \30539 );
nor \U$30201 ( \30544 , \30541 , \30543 );
not \U$30202 ( \30545 , \29412 );
not \U$30203 ( \30546 , \29402 );
or \U$30204 ( \30547 , \30545 , \30546 );
or \U$30205 ( \30548 , \29412 , \29402 );
nand \U$30206 ( \30549 , \30548 , \29391 );
nand \U$30207 ( \30550 , \30547 , \30549 );
xor \U$30208 ( \30551 , \30544 , \30550 );
xnor \U$30209 ( \30552 , \30535 , \30551 );
xor \U$30210 ( \30553 , \30523 , \30552 );
xor \U$30211 ( \30554 , \30504 , \30553 );
not \U$30212 ( \30555 , \29442 );
not \U$30213 ( \30556 , \29564 );
or \U$30214 ( \30557 , \30555 , \30556 );
not \U$30215 ( \30558 , \29561 );
not \U$30216 ( \30559 , \29441 );
or \U$30217 ( \30560 , \30558 , \30559 );
nand \U$30218 ( \30561 , \30560 , \29451 );
nand \U$30219 ( \30562 , \30557 , \30561 );
and \U$30220 ( \30563 , \30554 , \30562 );
and \U$30221 ( \30564 , \30504 , \30553 );
or \U$30222 ( \30565 , \30563 , \30564 );
xor \U$30223 ( \30566 , \30495 , \30565 );
xor \U$30224 ( \30567 , \30418 , \30424 );
xor \U$30225 ( \30568 , \30567 , \30429 );
not \U$30226 ( \30569 , \29413 );
not \U$30227 ( \30570 , \30569 );
not \U$30228 ( \30571 , \29426 );
or \U$30229 ( \30572 , \30570 , \30571 );
or \U$30230 ( \30573 , \29426 , \30569 );
nand \U$30231 ( \30574 , \30573 , \29421 );
nand \U$30232 ( \30575 , \30572 , \30574 );
xor \U$30233 ( \30576 , \30568 , \30575 );
xor \U$30234 ( \30577 , \30456 , \30461 );
xor \U$30235 ( \30578 , \30577 , \30467 );
not \U$30236 ( \30579 , \30578 );
not \U$30237 ( \30580 , \30579 );
not \U$30238 ( \30581 , \30452 );
xor \U$30239 ( \30582 , \30438 , \30581 );
xor \U$30240 ( \30583 , \30582 , \30444 );
not \U$30241 ( \30584 , \30583 );
not \U$30242 ( \30585 , \30584 );
or \U$30243 ( \30586 , \30580 , \30585 );
nand \U$30244 ( \30587 , \30583 , \30578 );
nand \U$30245 ( \30588 , \30586 , \30587 );
xor \U$30246 ( \30589 , \30481 , \30488 );
xnor \U$30247 ( \30590 , \30589 , \30476 );
buf \U$30248 ( \30591 , \30590 );
xor \U$30249 ( \30592 , \30588 , \30591 );
xor \U$30250 ( \30593 , \30576 , \30592 );
not \U$30251 ( \30594 , \30593 );
not \U$30252 ( \30595 , \30594 );
not \U$30253 ( \30596 , \30595 );
not \U$30254 ( \30597 , \30265 );
not \U$30255 ( \30598 , \30251 );
or \U$30256 ( \30599 , \30597 , \30598 );
or \U$30257 ( \30600 , \30265 , \30251 );
nand \U$30258 ( \30601 , \30599 , \30600 );
buf \U$30259 ( \30602 , \30255 );
and \U$30260 ( \30603 , \30601 , \30602 );
not \U$30261 ( \30604 , \30601 );
not \U$30262 ( \30605 , \30602 );
and \U$30263 ( \30606 , \30604 , \30605 );
nor \U$30264 ( \30607 , \30603 , \30606 );
not \U$30265 ( \30608 , \30607 );
not \U$30266 ( \30609 , \30608 );
or \U$30267 ( \30610 , \30596 , \30609 );
xor \U$30268 ( \30611 , \29427 , \29432 );
and \U$30269 ( \30612 , \30611 , \29440 );
and \U$30270 ( \30613 , \29427 , \29432 );
or \U$30271 ( \30614 , \30612 , \30613 );
not \U$30272 ( \30615 , \30614 );
nand \U$30273 ( \30616 , \30607 , \30594 );
nand \U$30274 ( \30617 , \30615 , \30616 );
nand \U$30275 ( \30618 , \30610 , \30617 );
not \U$30276 ( \30619 , \30618 );
xor \U$30277 ( \30620 , \30513 , \30522 );
and \U$30278 ( \30621 , \30620 , \30552 );
and \U$30279 ( \30622 , \30513 , \30522 );
or \U$30280 ( \30623 , \30621 , \30622 );
not \U$30281 ( \30624 , \30623 );
not \U$30282 ( \30625 , \30528 );
not \U$30283 ( \30626 , \30551 );
not \U$30284 ( \30627 , \30626 );
or \U$30285 ( \30628 , \30625 , \30627 );
not \U$30286 ( \30629 , \30528 );
nand \U$30287 ( \30630 , \30629 , \30551 );
nand \U$30288 ( \30631 , \30630 , \30534 );
nand \U$30289 ( \30632 , \30628 , \30631 );
not \U$30290 ( \30633 , \30632 );
not \U$30291 ( \30634 , \30539 );
not \U$30292 ( \30635 , \30537 );
or \U$30293 ( \30636 , \30634 , \30635 );
or \U$30294 ( \30637 , \30537 , \30539 );
nand \U$30295 ( \30638 , \30637 , \30550 );
nand \U$30296 ( \30639 , \30636 , \30638 );
not \U$30297 ( \30640 , RIbb2f0e8_12);
not \U$30298 ( \30641 , \30640 );
not \U$30299 ( \30642 , \1656 );
or \U$30300 ( \30643 , \30641 , \30642 );
nand \U$30301 ( \30644 , \30643 , \17506 );
and \U$30302 ( \30645 , RIbb2f0e8_12, RIbb2f070_13);
nor \U$30303 ( \30646 , \30645 , \1805 );
and \U$30304 ( \30647 , \30644 , \30646 );
not \U$30305 ( \30648 , \1077 );
not \U$30306 ( \30649 , RIbb2f160_11);
not \U$30307 ( \30650 , \17744 );
or \U$30308 ( \30651 , \30649 , \30650 );
nand \U$30309 ( \30652 , \17517 , \1805 );
nand \U$30310 ( \30653 , \30651 , \30652 );
not \U$30311 ( \30654 , \30653 );
or \U$30312 ( \30655 , \30648 , \30654 );
not \U$30313 ( \30656 , RIbb2f160_11);
not \U$30314 ( \30657 , \19063 );
or \U$30315 ( \30658 , \30656 , \30657 );
nand \U$30316 ( \30659 , \19064 , \1043 );
nand \U$30317 ( \30660 , \30658 , \30659 );
nand \U$30318 ( \30661 , \30660 , \1010 );
nand \U$30319 ( \30662 , \30655 , \30661 );
xor \U$30320 ( \30663 , \30647 , \30662 );
not \U$30321 ( \30664 , \998 );
and \U$30322 ( \30665 , \16703 , \3421 );
not \U$30323 ( \30666 , \16703 );
and \U$30324 ( \30667 , \30666 , RIbb2f070_13);
or \U$30325 ( \30668 , \30665 , \30667 );
not \U$30326 ( \30669 , \30668 );
or \U$30327 ( \30670 , \30664 , \30669 );
nand \U$30328 ( \30671 , \29896 , \915 );
nand \U$30329 ( \30672 , \30670 , \30671 );
xor \U$30330 ( \30673 , \30663 , \30672 );
not \U$30331 ( \30674 , \831 );
not \U$30332 ( \30675 , \30060 );
or \U$30333 ( \30676 , \30674 , \30675 );
not \U$30334 ( \30677 , RIbb2ee90_17);
not \U$30335 ( \30678 , \15823 );
or \U$30336 ( \30679 , \30677 , \30678 );
nand \U$30337 ( \30680 , \16575 , \3057 );
nand \U$30338 ( \30681 , \30679 , \30680 );
nand \U$30339 ( \30682 , \30681 , \835 );
nand \U$30340 ( \30683 , \30676 , \30682 );
xor \U$30341 ( \30684 , \30673 , \30683 );
not \U$30342 ( \30685 , \4714 );
not \U$30343 ( \30686 , RIbb2e620_35);
not \U$30344 ( \30687 , \7297 );
or \U$30345 ( \30688 , \30686 , \30687 );
nand \U$30346 ( \30689 , \7296 , \11338 );
nand \U$30347 ( \30690 , \30688 , \30689 );
not \U$30348 ( \30691 , \30690 );
or \U$30349 ( \30692 , \30685 , \30691 );
nand \U$30350 ( \30693 , \29987 , \4712 );
nand \U$30351 ( \30694 , \30692 , \30693 );
xor \U$30352 ( \30695 , \30684 , \30694 );
not \U$30353 ( \30696 , \6251 );
not \U$30354 ( \30697 , \30402 );
or \U$30355 ( \30698 , \30696 , \30697 );
not \U$30356 ( \30699 , RIbb2e530_37);
not \U$30357 ( \30700 , \13875 );
or \U$30358 ( \30701 , \30699 , \30700 );
nand \U$30359 ( \30702 , \6603 , \8701 );
nand \U$30360 ( \30703 , \30701 , \30702 );
nand \U$30361 ( \30704 , \30703 , \20792 );
nand \U$30362 ( \30705 , \30698 , \30704 );
xor \U$30363 ( \30706 , \30695 , \30705 );
not \U$30364 ( \30707 , \2939 );
not \U$30365 ( \30708 , \30354 );
or \U$30366 ( \30709 , \30707 , \30708 );
not \U$30367 ( \30710 , RIbb2e800_31);
not \U$30368 ( \30711 , \13498 );
or \U$30369 ( \30712 , \30710 , \30711 );
nand \U$30370 ( \30713 , \9840 , \8810 );
nand \U$30371 ( \30714 , \30712 , \30713 );
nand \U$30372 ( \30715 , \30714 , \2941 );
nand \U$30373 ( \30716 , \30709 , \30715 );
not \U$30374 ( \30717 , \3465 );
not \U$30375 ( \30718 , RIbb2e9e0_27);
not \U$30376 ( \30719 , \17440 );
or \U$30377 ( \30720 , \30718 , \30719 );
nand \U$30378 ( \30721 , \11578 , \3454 );
nand \U$30379 ( \30722 , \30720 , \30721 );
not \U$30380 ( \30723 , \30722 );
or \U$30381 ( \30724 , \30717 , \30723 );
nand \U$30382 ( \30725 , \29926 , \3445 );
nand \U$30383 ( \30726 , \30724 , \30725 );
xor \U$30384 ( \30727 , \30716 , \30726 );
not \U$30385 ( \30728 , \2922 );
not \U$30386 ( \30729 , \30364 );
or \U$30387 ( \30730 , \30728 , \30729 );
not \U$30388 ( \30731 , RIbb2e8f0_29);
not \U$30389 ( \30732 , \18802 );
or \U$30390 ( \30733 , \30731 , \30732 );
nand \U$30391 ( \30734 , \13526 , \3265 );
nand \U$30392 ( \30735 , \30733 , \30734 );
nand \U$30393 ( \30736 , \30735 , \2925 );
nand \U$30394 ( \30737 , \30730 , \30736 );
xnor \U$30395 ( \30738 , \30727 , \30737 );
xor \U$30396 ( \30739 , \30706 , \30738 );
not \U$30397 ( \30740 , \4075 );
and \U$30398 ( \30741 , \8630 , \2935 );
not \U$30399 ( \30742 , \8630 );
and \U$30400 ( \30743 , \30742 , RIbb2e710_33);
or \U$30401 ( \30744 , \30741 , \30743 );
not \U$30402 ( \30745 , \30744 );
or \U$30403 ( \30746 , \30740 , \30745 );
nand \U$30404 ( \30747 , \29963 , \3886 );
nand \U$30405 ( \30748 , \30746 , \30747 );
not \U$30406 ( \30749 , \30748 );
not \U$30407 ( \30750 , \8362 );
not \U$30408 ( \30751 , \30389 );
or \U$30409 ( \30752 , \30750 , \30751 );
not \U$30410 ( \30753 , RIbb2e350_41);
not \U$30411 ( \30754 , \4392 );
or \U$30412 ( \30755 , \30753 , \30754 );
nand \U$30413 ( \30756 , \20390 , \9402 );
nand \U$30414 ( \30757 , \30755 , \30756 );
nand \U$30415 ( \30758 , \30757 , \8354 );
nand \U$30416 ( \30759 , \30752 , \30758 );
not \U$30417 ( \30760 , \30759 );
not \U$30418 ( \30761 , \30760 );
or \U$30419 ( \30762 , \30749 , \30761 );
not \U$30420 ( \30763 , \30748 );
nand \U$30421 ( \30764 , \30759 , \30763 );
nand \U$30422 ( \30765 , \30762 , \30764 );
not \U$30423 ( \30766 , \7102 );
not \U$30424 ( \30767 , \30380 );
or \U$30425 ( \30768 , \30766 , \30767 );
not \U$30426 ( \30769 , RIbb2e440_39);
not \U$30427 ( \30770 , \6230 );
or \U$30428 ( \30771 , \30769 , \30770 );
nand \U$30429 ( \30772 , \6229 , \10908 );
nand \U$30430 ( \30773 , \30771 , \30772 );
nand \U$30431 ( \30774 , \30773 , \7104 );
nand \U$30432 ( \30775 , \30768 , \30774 );
buf \U$30433 ( \30776 , \30775 );
not \U$30434 ( \30777 , \30776 );
and \U$30435 ( \30778 , \30765 , \30777 );
not \U$30436 ( \30779 , \30765 );
and \U$30437 ( \30780 , \30779 , \30776 );
nor \U$30438 ( \30781 , \30778 , \30780 );
xnor \U$30439 ( \30782 , \30739 , \30781 );
xor \U$30440 ( \30783 , \30639 , \30782 );
not \U$30441 ( \30784 , \30584 );
not \U$30442 ( \30785 , \30590 );
or \U$30443 ( \30786 , \30784 , \30785 );
or \U$30444 ( \30787 , \30584 , \30590 );
nand \U$30445 ( \30788 , \30787 , \30578 );
nand \U$30446 ( \30789 , \30786 , \30788 );
xor \U$30447 ( \30790 , \30783 , \30789 );
not \U$30448 ( \30791 , \30790 );
or \U$30449 ( \30792 , \30633 , \30791 );
or \U$30450 ( \30793 , \30632 , \30790 );
nand \U$30451 ( \30794 , \30792 , \30793 );
not \U$30452 ( \30795 , \30568 );
not \U$30453 ( \30796 , \30592 );
or \U$30454 ( \30797 , \30795 , \30796 );
or \U$30455 ( \30798 , \30568 , \30592 );
nand \U$30456 ( \30799 , \30798 , \30575 );
nand \U$30457 ( \30800 , \30797 , \30799 );
not \U$30458 ( \30801 , \30800 );
and \U$30459 ( \30802 , \30794 , \30801 );
not \U$30460 ( \30803 , \30794 );
and \U$30461 ( \30804 , \30803 , \30800 );
nor \U$30462 ( \30805 , \30802 , \30804 );
not \U$30463 ( \30806 , \30805 );
and \U$30464 ( \30807 , \30624 , \30806 );
and \U$30465 ( \30808 , \30623 , \30805 );
nor \U$30466 ( \30809 , \30807 , \30808 );
not \U$30467 ( \30810 , \30809 );
or \U$30468 ( \30811 , \30619 , \30810 );
or \U$30469 ( \30812 , \30618 , \30809 );
nand \U$30470 ( \30813 , \30811 , \30812 );
xor \U$30471 ( \30814 , \30566 , \30813 );
xor \U$30472 ( \30815 , \30593 , \30614 );
xnor \U$30473 ( \30816 , \30815 , \30608 );
xor \U$30474 ( \30817 , \29572 , \29825 );
and \U$30475 ( \30818 , \30817 , \29830 );
and \U$30476 ( \30819 , \29572 , \29825 );
or \U$30477 ( \30820 , \30818 , \30819 );
xor \U$30478 ( \30821 , \30816 , \30820 );
xor \U$30479 ( \30822 , \30504 , \30553 );
xor \U$30480 ( \30823 , \30822 , \30562 );
and \U$30481 ( \30824 , \30821 , \30823 );
and \U$30482 ( \30825 , \30816 , \30820 );
or \U$30483 ( \30826 , \30824 , \30825 );
nor \U$30484 ( \30827 , \30814 , \30826 );
not \U$30485 ( \30828 , \30827 );
xor \U$30486 ( \30829 , \30816 , \30820 );
xor \U$30487 ( \30830 , \30829 , \30823 );
not \U$30488 ( \30831 , \30830 );
xor \U$30489 ( \30832 , \29568 , \29831 );
and \U$30490 ( \30833 , \30832 , \29840 );
and \U$30491 ( \30834 , \29568 , \29831 );
or \U$30492 ( \30835 , \30833 , \30834 );
not \U$30493 ( \30836 , \30835 );
nand \U$30494 ( \30837 , \30831 , \30836 );
nand \U$30495 ( \30838 , \30828 , \30837 );
not \U$30496 ( \30839 , \3465 );
not \U$30497 ( \30840 , RIbb2e9e0_27);
not \U$30498 ( \30841 , \12257 );
or \U$30499 ( \30842 , \30840 , \30841 );
nand \U$30500 ( \30843 , \11142 , \3454 );
nand \U$30501 ( \30844 , \30842 , \30843 );
not \U$30502 ( \30845 , \30844 );
or \U$30503 ( \30846 , \30839 , \30845 );
nand \U$30504 ( \30847 , \30722 , \3445 );
nand \U$30505 ( \30848 , \30846 , \30847 );
not \U$30506 ( \30849 , \3886 );
not \U$30507 ( \30850 , \30744 );
or \U$30508 ( \30851 , \30849 , \30850 );
not \U$30509 ( \30852 , RIbb2e710_33);
not \U$30510 ( \30853 , \23960 );
or \U$30511 ( \30854 , \30852 , \30853 );
nand \U$30512 ( \30855 , \8318 , \18295 );
nand \U$30513 ( \30856 , \30854 , \30855 );
nand \U$30514 ( \30857 , \30856 , \4791 );
nand \U$30515 ( \30858 , \30851 , \30857 );
xor \U$30516 ( \30859 , \30848 , \30858 );
not \U$30517 ( \30860 , \2921 );
not \U$30518 ( \30861 , \30735 );
or \U$30519 ( \30862 , \30860 , \30861 );
not \U$30520 ( \30863 , RIbb2e8f0_29);
not \U$30521 ( \30864 , \13929 );
or \U$30522 ( \30865 , \30863 , \30864 );
nand \U$30523 ( \30866 , \10300 , \3440 );
nand \U$30524 ( \30867 , \30865 , \30866 );
nand \U$30525 ( \30868 , \30867 , \2925 );
nand \U$30526 ( \30869 , \30862 , \30868 );
xor \U$30527 ( \30870 , \30859 , \30869 );
xor \U$30528 ( \30871 , \30325 , \30334 );
and \U$30529 ( \30872 , \30871 , \30345 );
and \U$30530 ( \30873 , \30325 , \30334 );
or \U$30531 ( \30874 , \30872 , \30873 );
not \U$30532 ( \30875 , \16271 );
not \U$30533 ( \30876 , \30159 );
or \U$30534 ( \30877 , \30875 , \30876 );
and \U$30535 ( \30878 , RIbb2dae0_59, \15582 );
not \U$30536 ( \30879 , RIbb2dae0_59);
and \U$30537 ( \30880 , \30879 , \1280 );
or \U$30538 ( \30881 , \30878 , \30880 );
nand \U$30539 ( \30882 , \30881 , \17470 );
nand \U$30540 ( \30883 , \30877 , \30882 );
xor \U$30541 ( \30884 , \30874 , \30883 );
not \U$30542 ( \30885 , \14067 );
not \U$30543 ( \30886 , \30167 );
or \U$30544 ( \30887 , \30885 , \30886 );
and \U$30545 ( \30888 , RIbb2dea0_51, \20951 );
not \U$30546 ( \30889 , RIbb2dea0_51);
and \U$30547 ( \30890 , \30889 , \3341 );
or \U$30548 ( \30891 , \30888 , \30890 );
nand \U$30549 ( \30892 , \30891 , \12692 );
nand \U$30550 ( \30893 , \30887 , \30892 );
xor \U$30551 ( \30894 , \30884 , \30893 );
xor \U$30552 ( \30895 , \30870 , \30894 );
not \U$30553 ( \30896 , \11177 );
not \U$30554 ( \30897 , RIbb2e080_47);
not \U$30555 ( \30898 , \13835 );
or \U$30556 ( \30899 , \30897 , \30898 );
nand \U$30557 ( \30900 , \6171 , \16171 );
nand \U$30558 ( \30901 , \30899 , \30900 );
not \U$30559 ( \30902 , \30901 );
or \U$30560 ( \30903 , \30896 , \30902 );
nand \U$30561 ( \30904 , \30031 , \11176 );
nand \U$30562 ( \30905 , \30903 , \30904 );
not \U$30563 ( \30906 , \12167 );
not \U$30564 ( \30907 , \30104 );
or \U$30565 ( \30908 , \30906 , \30907 );
not \U$30566 ( \30909 , RIbb2df90_49);
not \U$30567 ( \30910 , \15398 );
or \U$30568 ( \30911 , \30909 , \30910 );
nand \U$30569 ( \30912 , \3146 , \12278 );
nand \U$30570 ( \30913 , \30911 , \30912 );
nand \U$30571 ( \30914 , \30913 , \14752 );
nand \U$30572 ( \30915 , \30908 , \30914 );
xor \U$30573 ( \30916 , \30905 , \30915 );
not \U$30574 ( \30917 , \15738 );
not \U$30575 ( \30918 , RIbb2dbd0_57);
not \U$30576 ( \30919 , \1385 );
or \U$30577 ( \30920 , \30918 , \30919 );
nand \U$30578 ( \30921 , \1386 , \17411 );
nand \U$30579 ( \30922 , \30920 , \30921 );
not \U$30580 ( \30923 , \30922 );
or \U$30581 ( \30924 , \30917 , \30923 );
nand \U$30582 ( \30925 , \30009 , \19101 );
nand \U$30583 ( \30926 , \30924 , \30925 );
xor \U$30584 ( \30927 , \30916 , \30926 );
xnor \U$30585 ( \30928 , \30895 , \30927 );
not \U$30586 ( \30929 , \30928 );
and \U$30587 ( \30930 , \30647 , \30662 );
not \U$30588 ( \30931 , \1517 );
not \U$30589 ( \30932 , RIbb2ef80_15);
not \U$30590 ( \30933 , \16747 );
or \U$30591 ( \30934 , \30932 , \30933 );
not \U$30592 ( \30935 , RIbb2ef80_15);
nand \U$30593 ( \30936 , \30935 , \19077 );
nand \U$30594 ( \30937 , \30934 , \30936 );
not \U$30595 ( \30938 , \30937 );
or \U$30596 ( \30939 , \30931 , \30938 );
nand \U$30597 ( \30940 , \30280 , \1444 );
nand \U$30598 ( \30941 , \30939 , \30940 );
xor \U$30599 ( \30942 , \30930 , \30941 );
not \U$30600 ( \30943 , \836 );
and \U$30601 ( \30944 , RIbb2ee90_17, \16562 );
not \U$30602 ( \30945 , RIbb2ee90_17);
and \U$30603 ( \30946 , \30945 , \15754 );
nor \U$30604 ( \30947 , \30944 , \30946 );
not \U$30605 ( \30948 , \30947 );
or \U$30606 ( \30949 , \30943 , \30948 );
nand \U$30607 ( \30950 , \30681 , \831 );
nand \U$30608 ( \30951 , \30949 , \30950 );
xor \U$30609 ( \30952 , \30942 , \30951 );
not \U$30610 ( \30953 , RIbb2d888_64);
not \U$30611 ( \30954 , RIbb2d900_63);
not \U$30612 ( \30955 , \3368 );
or \U$30613 ( \30956 , \30954 , \30955 );
nand \U$30614 ( \30957 , \1687 , \22946 );
nand \U$30615 ( \30958 , \30956 , \30957 );
not \U$30616 ( \30959 , \30958 );
or \U$30617 ( \30960 , \30953 , \30959 );
nand \U$30618 ( \30961 , \30148 , \17275 );
nand \U$30619 ( \30962 , \30960 , \30961 );
xor \U$30620 ( \30963 , \30952 , \30962 );
not \U$30621 ( \30964 , \15688 );
not \U$30622 ( \30965 , RIbb2ddb0_53);
not \U$30623 ( \30966 , \3310 );
or \U$30624 ( \30967 , \30965 , \30966 );
nand \U$30625 ( \30968 , \3309 , \16210 );
nand \U$30626 ( \30969 , \30967 , \30968 );
not \U$30627 ( \30970 , \30969 );
or \U$30628 ( \30971 , \30964 , \30970 );
nand \U$30629 ( \30972 , \30203 , \17562 );
nand \U$30630 ( \30973 , \30971 , \30972 );
xor \U$30631 ( \30974 , \30963 , \30973 );
not \U$30632 ( \30975 , \10117 );
not \U$30633 ( \30976 , \30047 );
or \U$30634 ( \30977 , \30975 , \30976 );
not \U$30635 ( \30978 , RIbb2e170_45);
not \U$30636 ( \30979 , \3021 );
or \U$30637 ( \30980 , \30978 , \30979 );
not \U$30638 ( \30981 , \3021 );
nand \U$30639 ( \30982 , \30981 , \12003 );
nand \U$30640 ( \30983 , \30980 , \30982 );
nand \U$30641 ( \30984 , \30983 , \10119 );
nand \U$30642 ( \30985 , \30977 , \30984 );
not \U$30643 ( \30986 , \15181 );
and \U$30644 ( \30987 , RIbb2dcc0_55, \19733 );
not \U$30645 ( \30988 , RIbb2dcc0_55);
and \U$30646 ( \30989 , \30988 , \1337 );
or \U$30647 ( \30990 , \30987 , \30989 );
not \U$30648 ( \30991 , \30990 );
or \U$30649 ( \30992 , \30986 , \30991 );
nand \U$30650 ( \30993 , \30220 , \14613 );
nand \U$30651 ( \30994 , \30992 , \30993 );
xor \U$30652 ( \30995 , \30985 , \30994 );
not \U$30653 ( \30996 , \9098 );
not \U$30654 ( \30997 , \30180 );
or \U$30655 ( \30998 , \30996 , \30997 );
not \U$30656 ( \30999 , RIbb2e260_43);
not \U$30657 ( \31000 , \25942 );
or \U$30658 ( \31001 , \30999 , \31000 );
nand \U$30659 ( \31002 , \13732 , \13772 );
nand \U$30660 ( \31003 , \31001 , \31002 );
nand \U$30661 ( \31004 , \31003 , \9099 );
nand \U$30662 ( \31005 , \30998 , \31004 );
xor \U$30663 ( \31006 , \30995 , \31005 );
xor \U$30664 ( \31007 , \30974 , \31006 );
xor \U$30665 ( \31008 , \30300 , \30304 );
and \U$30666 ( \31009 , \31008 , \30309 );
and \U$30667 ( \31010 , \30300 , \30304 );
or \U$30668 ( \31011 , \31009 , \31010 );
not \U$30669 ( \31012 , \31011 );
xor \U$30670 ( \31013 , \31007 , \31012 );
not \U$30671 ( \31014 , \31013 );
not \U$30672 ( \31015 , \31014 );
or \U$30673 ( \31016 , \30929 , \31015 );
not \U$30674 ( \31017 , \30928 );
nand \U$30675 ( \31018 , \31017 , \31013 );
nand \U$30676 ( \31019 , \31016 , \31018 );
xor \U$30677 ( \31020 , \30310 , \30314 );
and \U$30678 ( \31021 , \31020 , \30408 );
and \U$30679 ( \31022 , \30310 , \30314 );
or \U$30680 ( \31023 , \31021 , \31022 );
buf \U$30681 ( \31024 , \31023 );
not \U$30682 ( \31025 , \31024 );
and \U$30683 ( \31026 , \31019 , \31025 );
not \U$30684 ( \31027 , \31019 );
and \U$30685 ( \31028 , \31027 , \31024 );
nor \U$30686 ( \31029 , \31026 , \31028 );
xor \U$30687 ( \31030 , \30275 , \30409 );
and \U$30688 ( \31031 , \31030 , \30493 );
and \U$30689 ( \31032 , \30275 , \30409 );
or \U$30690 ( \31033 , \31031 , \31032 );
xor \U$30691 ( \31034 , \31029 , \31033 );
not \U$30692 ( \31035 , \30632 );
not \U$30693 ( \31036 , \31035 );
not \U$30694 ( \31037 , \30790 );
or \U$30695 ( \31038 , \31036 , \31037 );
nand \U$30696 ( \31039 , \31038 , \30800 );
not \U$30697 ( \31040 , \30790 );
not \U$30698 ( \31041 , \31035 );
nand \U$30699 ( \31042 , \31040 , \31041 );
nand \U$30700 ( \31043 , \31039 , \31042 );
xnor \U$30701 ( \31044 , \31034 , \31043 );
not \U$30702 ( \31045 , \30748 );
not \U$30703 ( \31046 , \30775 );
or \U$30704 ( \31047 , \31045 , \31046 );
not \U$30705 ( \31048 , \30775 );
not \U$30706 ( \31049 , \31048 );
not \U$30707 ( \31050 , \30763 );
or \U$30708 ( \31051 , \31049 , \31050 );
nand \U$30709 ( \31052 , \31051 , \30759 );
nand \U$30710 ( \31053 , \31047 , \31052 );
not \U$30711 ( \31054 , \31053 );
xor \U$30712 ( \31055 , \30284 , \30288 );
and \U$30713 ( \31056 , \31055 , \30299 );
and \U$30714 ( \31057 , \30284 , \30288 );
or \U$30715 ( \31058 , \31056 , \31057 );
not \U$30716 ( \31059 , \31058 );
not \U$30717 ( \31060 , \31059 );
and \U$30718 ( \31061 , \31054 , \31060 );
and \U$30719 ( \31062 , \31053 , \31059 );
nor \U$30720 ( \31063 , \31061 , \31062 );
not \U$30721 ( \31064 , \30737 );
not \U$30722 ( \31065 , \30716 );
or \U$30723 ( \31066 , \31064 , \31065 );
or \U$30724 ( \31067 , \30716 , \30737 );
nand \U$30725 ( \31068 , \31067 , \30726 );
nand \U$30726 ( \31069 , \31066 , \31068 );
xnor \U$30727 ( \31070 , \31063 , \31069 );
xor \U$30728 ( \31071 , \30346 , \30375 );
and \U$30729 ( \31072 , \31071 , \30407 );
and \U$30730 ( \31073 , \30346 , \30375 );
or \U$30731 ( \31074 , \31072 , \31073 );
xor \U$30732 ( \31075 , \31070 , \31074 );
not \U$30733 ( \31076 , \30738 );
not \U$30734 ( \31077 , \30781 );
or \U$30735 ( \31078 , \31076 , \31077 );
nand \U$30736 ( \31079 , \31078 , \30706 );
or \U$30737 ( \31080 , \30781 , \30738 );
nand \U$30738 ( \31081 , \31079 , \31080 );
xor \U$30739 ( \31082 , \31075 , \31081 );
not \U$30740 ( \31083 , \30639 );
not \U$30741 ( \31084 , \31083 );
not \U$30742 ( \31085 , \30782 );
or \U$30743 ( \31086 , \31084 , \31085 );
nand \U$30744 ( \31087 , \31086 , \30789 );
or \U$30745 ( \31088 , \30782 , \31083 );
nand \U$30746 ( \31089 , \31087 , \31088 );
xor \U$30747 ( \31090 , \31082 , \31089 );
xor \U$30748 ( \31091 , \30416 , \30432 );
and \U$30749 ( \31092 , \31091 , \30492 );
and \U$30750 ( \31093 , \30416 , \30432 );
or \U$30751 ( \31094 , \31092 , \31093 );
xor \U$30752 ( \31095 , \31090 , \31094 );
and \U$30753 ( \31096 , \17506 , \1531 );
not \U$30754 ( \31097 , \1077 );
and \U$30755 ( \31098 , \18908 , RIbb2f160_11);
not \U$30756 ( \31099 , \18908 );
and \U$30757 ( \31100 , \31099 , \1805 );
or \U$30758 ( \31101 , \31098 , \31100 );
not \U$30759 ( \31102 , \31101 );
or \U$30760 ( \31103 , \31097 , \31102 );
nand \U$30761 ( \31104 , \30653 , \1010 );
nand \U$30762 ( \31105 , \31103 , \31104 );
xor \U$30763 ( \31106 , \31096 , \31105 );
not \U$30764 ( \31107 , \915 );
not \U$30765 ( \31108 , \30668 );
or \U$30766 ( \31109 , \31107 , \31108 );
and \U$30767 ( \31110 , \16553 , \1656 );
not \U$30768 ( \31111 , \16553 );
and \U$30769 ( \31112 , \31111 , RIbb2f070_13);
or \U$30770 ( \31113 , \31110 , \31112 );
nand \U$30771 ( \31114 , \31113 , \997 );
nand \U$30772 ( \31115 , \31109 , \31114 );
xor \U$30773 ( \31116 , \31106 , \31115 );
not \U$30774 ( \31117 , \3406 );
not \U$30775 ( \31118 , \30297 );
or \U$30776 ( \31119 , \31117 , \31118 );
not \U$30777 ( \31120 , RIbb2ebc0_23);
not \U$30778 ( \31121 , \24290 );
or \U$30779 ( \31122 , \31120 , \31121 );
not \U$30780 ( \31123 , RIbb2ebc0_23);
nand \U$30781 ( \31124 , \31123 , \12346 );
nand \U$30782 ( \31125 , \31122 , \31124 );
nand \U$30783 ( \31126 , \31125 , \3381 );
nand \U$30784 ( \31127 , \31119 , \31126 );
xor \U$30785 ( \31128 , \31116 , \31127 );
not \U$30786 ( \31129 , \2077 );
not \U$30787 ( \31130 , \30343 );
or \U$30788 ( \31131 , \31129 , \31130 );
not \U$30789 ( \31132 , RIbb2ecb0_21);
not \U$30790 ( \31133 , \18552 );
or \U$30791 ( \31134 , \31132 , \31133 );
nand \U$30792 ( \31135 , \13545 , \2067 );
nand \U$30793 ( \31136 , \31134 , \31135 );
nand \U$30794 ( \31137 , \31136 , \2078 );
nand \U$30795 ( \31138 , \31131 , \31137 );
xor \U$30796 ( \31139 , \31128 , \31138 );
xor \U$30797 ( \31140 , \30684 , \30694 );
and \U$30798 ( \31141 , \31140 , \30705 );
and \U$30799 ( \31142 , \30684 , \30694 );
or \U$30800 ( \31143 , \31141 , \31142 );
xor \U$30801 ( \31144 , \31139 , \31143 );
not \U$30802 ( \31145 , \853 );
not \U$30803 ( \31146 , \30321 );
or \U$30804 ( \31147 , \31145 , \31146 );
and \U$30805 ( \31148 , \14526 , \1776 );
not \U$30806 ( \31149 , \14526 );
and \U$30807 ( \31150 , \31149 , RIbb2eda0_19);
or \U$30808 ( \31151 , \31148 , \31150 );
nand \U$30809 ( \31152 , \31151 , \854 );
nand \U$30810 ( \31153 , \31147 , \31152 );
not \U$30811 ( \31154 , \2963 );
xor \U$30812 ( \31155 , \12174 , RIbb2ead0_25);
not \U$30813 ( \31156 , \31155 );
or \U$30814 ( \31157 , \31154 , \31156 );
nand \U$30815 ( \31158 , \30332 , \2980 );
nand \U$30816 ( \31159 , \31157 , \31158 );
xor \U$30817 ( \31160 , \31153 , \31159 );
not \U$30818 ( \31161 , \2939 );
not \U$30819 ( \31162 , \30714 );
or \U$30820 ( \31163 , \31161 , \31162 );
not \U$30821 ( \31164 , RIbb2e800_31);
not \U$30822 ( \31165 , \29959 );
or \U$30823 ( \31166 , \31164 , \31165 );
nand \U$30824 ( \31167 , \9277 , \11975 );
nand \U$30825 ( \31168 , \31166 , \31167 );
nand \U$30826 ( \31169 , \31168 , \2941 );
nand \U$30827 ( \31170 , \31163 , \31169 );
xor \U$30828 ( \31171 , \31160 , \31170 );
xor \U$30829 ( \31172 , \31144 , \31171 );
not \U$30830 ( \31173 , \30491 );
not \U$30831 ( \31174 , \30454 );
or \U$30832 ( \31175 , \31173 , \31174 );
or \U$30833 ( \31176 , \30454 , \30491 );
nand \U$30834 ( \31177 , \31176 , \30470 );
nand \U$30835 ( \31178 , \31175 , \31177 );
xor \U$30836 ( \31179 , \31172 , \31178 );
xor \U$30837 ( \31180 , \30140 , \30173 );
and \U$30838 ( \31181 , \31180 , \30223 );
and \U$30839 ( \31182 , \30140 , \30173 );
or \U$30840 ( \31183 , \31181 , \31182 );
xor \U$30841 ( \31184 , \31179 , \31183 );
xor \U$30842 ( \31185 , \30003 , \30050 );
and \U$30843 ( \31186 , \31185 , \30107 );
and \U$30844 ( \31187 , \30003 , \30050 );
or \U$30845 ( \31188 , \31186 , \31187 );
xor \U$30846 ( \31189 , \30018 , \30033 );
and \U$30847 ( \31190 , \31189 , \30049 );
and \U$30848 ( \31191 , \30018 , \30033 );
or \U$30849 ( \31192 , \31190 , \31191 );
xor \U$30850 ( \31193 , \30075 , \30090 );
and \U$30851 ( \31194 , \31193 , \30106 );
and \U$30852 ( \31195 , \30075 , \30090 );
or \U$30853 ( \31196 , \31194 , \31195 );
xor \U$30854 ( \31197 , \31192 , \31196 );
or \U$30855 ( \31198 , \30205 , \30222 );
nand \U$30856 ( \31199 , \31198 , \30189 );
nand \U$30857 ( \31200 , \30205 , \30222 );
nand \U$30858 ( \31201 , \31199 , \31200 );
xor \U$30859 ( \31202 , \31197 , \31201 );
xor \U$30860 ( \31203 , \31188 , \31202 );
not \U$30861 ( \31204 , \7103 );
not \U$30862 ( \31205 , \30773 );
or \U$30863 ( \31206 , \31204 , \31205 );
not \U$30864 ( \31207 , RIbb2e440_39);
not \U$30865 ( \31208 , \10555 );
or \U$30866 ( \31209 , \31207 , \31208 );
nand \U$30867 ( \31210 , \18623 , \10908 );
nand \U$30868 ( \31211 , \31209 , \31210 );
nand \U$30869 ( \31212 , \31211 , \8450 );
nand \U$30870 ( \31213 , \31206 , \31212 );
not \U$30871 ( \31214 , \6251 );
not \U$30872 ( \31215 , \30703 );
or \U$30873 ( \31216 , \31214 , \31215 );
not \U$30874 ( \31217 , RIbb2e530_37);
not \U$30875 ( \31218 , \18564 );
or \U$30876 ( \31219 , \31217 , \31218 );
nand \U$30877 ( \31220 , \7308 , \6246 );
nand \U$30878 ( \31221 , \31219 , \31220 );
nand \U$30879 ( \31222 , \31221 , \20792 );
nand \U$30880 ( \31223 , \31216 , \31222 );
xor \U$30881 ( \31224 , \31213 , \31223 );
not \U$30882 ( \31225 , \8353 );
not \U$30883 ( \31226 , RIbb2e350_41);
not \U$30884 ( \31227 , \4087 );
or \U$30885 ( \31228 , \31226 , \31227 );
nand \U$30886 ( \31229 , \4086 , \9402 );
nand \U$30887 ( \31230 , \31228 , \31229 );
not \U$30888 ( \31231 , \31230 );
or \U$30889 ( \31232 , \31225 , \31231 );
nand \U$30890 ( \31233 , \30757 , \8362 );
nand \U$30891 ( \31234 , \31232 , \31233 );
xor \U$30892 ( \31235 , \31224 , \31234 );
xor \U$30893 ( \31236 , \30663 , \30672 );
and \U$30894 ( \31237 , \31236 , \30683 );
and \U$30895 ( \31238 , \30663 , \30672 );
or \U$30896 ( \31239 , \31237 , \31238 );
not \U$30897 ( \31240 , \4712 );
not \U$30898 ( \31241 , \30690 );
or \U$30899 ( \31242 , \31240 , \31241 );
not \U$30900 ( \31243 , RIbb2e620_35);
not \U$30901 ( \31244 , \25845 );
or \U$30902 ( \31245 , \31243 , \31244 );
nand \U$30903 ( \31246 , \26232 , \6002 );
nand \U$30904 ( \31247 , \31245 , \31246 );
nand \U$30905 ( \31248 , \31247 , \5845 );
nand \U$30906 ( \31249 , \31242 , \31248 );
xor \U$30907 ( \31250 , \31239 , \31249 );
not \U$30908 ( \31251 , \16533 );
not \U$30909 ( \31252 , RIbb2d9f0_61);
not \U$30910 ( \31253 , \7423 );
or \U$30911 ( \31254 , \31252 , \31253 );
nand \U$30912 ( \31255 , \1136 , \16254 );
nand \U$30913 ( \31256 , \31254 , \31255 );
not \U$30914 ( \31257 , \31256 );
or \U$30915 ( \31258 , \31251 , \31257 );
nand \U$30916 ( \31259 , \30088 , \16541 );
nand \U$30917 ( \31260 , \31258 , \31259 );
xor \U$30918 ( \31261 , \31250 , \31260 );
xor \U$30919 ( \31262 , \31235 , \31261 );
xor \U$30920 ( \31263 , \30150 , \30161 );
and \U$30921 ( \31264 , \31263 , \30172 );
and \U$30922 ( \31265 , \30150 , \30161 );
or \U$30923 ( \31266 , \31264 , \31265 );
xor \U$30924 ( \31267 , \31262 , \31266 );
xor \U$30925 ( \31268 , \31203 , \31267 );
xor \U$30926 ( \31269 , \31184 , \31268 );
not \U$30927 ( \31270 , \29974 );
not \U$30928 ( \31271 , \30108 );
nand \U$30929 ( \31272 , \31271 , \30225 );
not \U$30930 ( \31273 , \31272 );
or \U$30931 ( \31274 , \31270 , \31273 );
not \U$30932 ( \31275 , \30225 );
nand \U$30933 ( \31276 , \31275 , \30108 );
nand \U$30934 ( \31277 , \31274 , \31276 );
xor \U$30935 ( \31278 , \31269 , \31277 );
xor \U$30936 ( \31279 , \31095 , \31278 );
xor \U$30937 ( \31280 , \30233 , \30267 );
and \U$30938 ( \31281 , \31280 , \30494 );
and \U$30939 ( \31282 , \30233 , \30267 );
or \U$30940 ( \31283 , \31281 , \31282 );
xor \U$30941 ( \31284 , \31279 , \31283 );
xor \U$30942 ( \31285 , \31044 , \31284 );
not \U$30943 ( \31286 , \30623 );
buf \U$30944 ( \31287 , \30805 );
nand \U$30945 ( \31288 , \31286 , \31287 );
not \U$30946 ( \31289 , \31288 );
not \U$30947 ( \31290 , \30618 );
or \U$30948 ( \31291 , \31289 , \31290 );
not \U$30949 ( \31292 , \31287 );
buf \U$30950 ( \31293 , \30623 );
nand \U$30951 ( \31294 , \31292 , \31293 );
nand \U$30952 ( \31295 , \31291 , \31294 );
xor \U$30953 ( \31296 , \31285 , \31295 );
not \U$30954 ( \31297 , \31296 );
xor \U$30955 ( \31298 , \30495 , \30565 );
and \U$30956 ( \31299 , \31298 , \30813 );
and \U$30957 ( \31300 , \30495 , \30565 );
or \U$30958 ( \31301 , \31299 , \31300 );
not \U$30959 ( \31302 , \31301 );
nand \U$30960 ( \31303 , \31297 , \31302 );
xor \U$30961 ( \31304 , \31044 , \31284 );
and \U$30962 ( \31305 , \31304 , \31295 );
and \U$30963 ( \31306 , \31044 , \31284 );
or \U$30964 ( \31307 , \31305 , \31306 );
not \U$30965 ( \31308 , \31307 );
xor \U$30966 ( \31309 , \30930 , \30941 );
and \U$30967 ( \31310 , \31309 , \30951 );
and \U$30968 ( \31311 , \30930 , \30941 );
or \U$30969 ( \31312 , \31310 , \31311 );
not \U$30970 ( \31313 , \18717 );
not \U$30971 ( \31314 , \31256 );
or \U$30972 ( \31315 , \31313 , \31314 );
not \U$30973 ( \31316 , RIbb2d9f0_61);
not \U$30974 ( \31317 , \3238 );
or \U$30975 ( \31318 , \31316 , \31317 );
nand \U$30976 ( \31319 , \1642 , \21449 );
nand \U$30977 ( \31320 , \31318 , \31319 );
nand \U$30978 ( \31321 , \31320 , \16533 );
nand \U$30979 ( \31322 , \31315 , \31321 );
xor \U$30980 ( \31323 , \31312 , \31322 );
not \U$30981 ( \31324 , \14752 );
not \U$30982 ( \31325 , RIbb2df90_49);
not \U$30983 ( \31326 , \13414 );
or \U$30984 ( \31327 , \31325 , \31326 );
nand \U$30985 ( \31328 , \3166 , \12278 );
nand \U$30986 ( \31329 , \31327 , \31328 );
not \U$30987 ( \31330 , \31329 );
or \U$30988 ( \31331 , \31324 , \31330 );
nand \U$30989 ( \31332 , \30913 , \13295 );
nand \U$30990 ( \31333 , \31331 , \31332 );
xor \U$30991 ( \31334 , \31323 , \31333 );
not \U$30992 ( \31335 , \30883 );
not \U$30993 ( \31336 , \30893 );
or \U$30994 ( \31337 , \31335 , \31336 );
or \U$30995 ( \31338 , \30893 , \30883 );
nand \U$30996 ( \31339 , \31338 , \30874 );
nand \U$30997 ( \31340 , \31337 , \31339 );
xor \U$30998 ( \31341 , \31334 , \31340 );
not \U$30999 ( \31342 , \12774 );
not \U$31000 ( \31343 , \30891 );
or \U$31001 ( \31344 , \31342 , \31343 );
xor \U$31002 ( \31345 , RIbb2dea0_51, \2222 );
nand \U$31003 ( \31346 , \31345 , \12692 );
nand \U$31004 ( \31347 , \31344 , \31346 );
not \U$31005 ( \31348 , \17562 );
not \U$31006 ( \31349 , \30969 );
or \U$31007 ( \31350 , \31348 , \31349 );
and \U$31008 ( \31351 , \14725 , RIbb2ddb0_53);
not \U$31009 ( \31352 , \14725 );
and \U$31010 ( \31353 , \31352 , \16210 );
or \U$31011 ( \31354 , \31351 , \31353 );
nand \U$31012 ( \31355 , \31354 , \14930 );
nand \U$31013 ( \31356 , \31350 , \31355 );
not \U$31014 ( \31357 , \31356 );
xor \U$31015 ( \31358 , \31347 , \31357 );
not \U$31016 ( \31359 , \16271 );
not \U$31017 ( \31360 , \30881 );
or \U$31018 ( \31361 , \31359 , \31360 );
xnor \U$31019 ( \31362 , RIbb2dae0_59, \1110 );
nand \U$31020 ( \31363 , \31362 , \16257 );
nand \U$31021 ( \31364 , \31361 , \31363 );
xnor \U$31022 ( \31365 , \31358 , \31364 );
xor \U$31023 ( \31366 , \31341 , \31365 );
xor \U$31024 ( \31367 , \31096 , \31105 );
and \U$31025 ( \31368 , \31367 , \31115 );
and \U$31026 ( \31369 , \31096 , \31105 );
or \U$31027 ( \31370 , \31368 , \31369 );
not \U$31028 ( \31371 , \1444 );
not \U$31029 ( \31372 , \30937 );
or \U$31030 ( \31373 , \31371 , \31372 );
nand \U$31031 ( \31374 , \24035 , \1517 );
nand \U$31032 ( \31375 , \31373 , \31374 );
xor \U$31033 ( \31376 , \31370 , \31375 );
not \U$31034 ( \31377 , \2078 );
not \U$31035 ( \31378 , \24366 );
or \U$31036 ( \31379 , \31377 , \31378 );
nand \U$31037 ( \31380 , \31136 , \2077 );
nand \U$31038 ( \31381 , \31379 , \31380 );
xor \U$31039 ( \31382 , \31376 , \31381 );
xor \U$31040 ( \31383 , \31116 , \31127 );
and \U$31041 ( \31384 , \31383 , \31138 );
and \U$31042 ( \31385 , \31116 , \31127 );
or \U$31043 ( \31386 , \31384 , \31385 );
xor \U$31044 ( \31387 , \31382 , \31386 );
not \U$31045 ( \31388 , RIbb2d888_64);
not \U$31046 ( \31389 , RIbb2d900_63);
not \U$31047 ( \31390 , \3479 );
or \U$31048 ( \31391 , \31389 , \31390 );
nand \U$31049 ( \31392 , \1730 , \20254 );
nand \U$31050 ( \31393 , \31391 , \31392 );
not \U$31051 ( \31394 , \31393 );
or \U$31052 ( \31395 , \31388 , \31394 );
nand \U$31053 ( \31396 , \30958 , \17275 );
nand \U$31054 ( \31397 , \31395 , \31396 );
xor \U$31055 ( \31398 , \31387 , \31397 );
xor \U$31056 ( \31399 , \31139 , \31143 );
and \U$31057 ( \31400 , \31399 , \31171 );
and \U$31058 ( \31401 , \31139 , \31143 );
or \U$31059 ( \31402 , \31400 , \31401 );
xor \U$31060 ( \31403 , \31398 , \31402 );
not \U$31061 ( \31404 , \8353 );
not \U$31062 ( \31405 , RIbb2e350_41);
not \U$31063 ( \31406 , \3090 );
or \U$31064 ( \31407 , \31405 , \31406 );
nand \U$31065 ( \31408 , \3089 , \9402 );
nand \U$31066 ( \31409 , \31407 , \31408 );
not \U$31067 ( \31410 , \31409 );
or \U$31068 ( \31411 , \31404 , \31410 );
nand \U$31069 ( \31412 , \31230 , \8361 );
nand \U$31070 ( \31413 , \31411 , \31412 );
not \U$31071 ( \31414 , \31413 );
not \U$31072 ( \31415 , \9099 );
not \U$31073 ( \31416 , RIbb2e260_43);
not \U$31074 ( \31417 , \4028 );
or \U$31075 ( \31418 , \31416 , \31417 );
nand \U$31076 ( \31419 , \16180 , \8347 );
nand \U$31077 ( \31420 , \31418 , \31419 );
not \U$31078 ( \31421 , \31420 );
or \U$31079 ( \31422 , \31415 , \31421 );
nand \U$31080 ( \31423 , \31003 , \9098 );
nand \U$31081 ( \31424 , \31422 , \31423 );
xor \U$31082 ( \31425 , \31414 , \31424 );
not \U$31083 ( \31426 , \15181 );
and \U$31084 ( \31427 , RIbb2dcc0_55, \17386 );
not \U$31085 ( \31428 , RIbb2dcc0_55);
and \U$31086 ( \31429 , \31428 , \1419 );
or \U$31087 ( \31430 , \31427 , \31429 );
not \U$31088 ( \31431 , \31430 );
or \U$31089 ( \31432 , \31426 , \31431 );
nand \U$31090 ( \31433 , \30990 , \14613 );
nand \U$31091 ( \31434 , \31432 , \31433 );
not \U$31092 ( \31435 , \31434 );
xor \U$31093 ( \31436 , \31425 , \31435 );
xor \U$31094 ( \31437 , \31403 , \31436 );
xor \U$31095 ( \31438 , \31366 , \31437 );
xor \U$31096 ( \31439 , \31070 , \31074 );
and \U$31097 ( \31440 , \31439 , \31081 );
and \U$31098 ( \31441 , \31070 , \31074 );
or \U$31099 ( \31442 , \31440 , \31441 );
xor \U$31100 ( \31443 , \31438 , \31442 );
xor \U$31101 ( \31444 , \31082 , \31089 );
and \U$31102 ( \31445 , \31444 , \31094 );
and \U$31103 ( \31446 , \31082 , \31089 );
or \U$31104 ( \31447 , \31445 , \31446 );
xor \U$31105 ( \31448 , \31443 , \31447 );
xor \U$31106 ( \31449 , \31188 , \31202 );
and \U$31107 ( \31450 , \31449 , \31267 );
and \U$31108 ( \31451 , \31188 , \31202 );
or \U$31109 ( \31452 , \31450 , \31451 );
not \U$31110 ( \31453 , \31452 );
xor \U$31111 ( \31454 , \31172 , \31178 );
and \U$31112 ( \31455 , \31454 , \31183 );
and \U$31113 ( \31456 , \31172 , \31178 );
or \U$31114 ( \31457 , \31455 , \31456 );
not \U$31115 ( \31458 , \31125 );
not \U$31116 ( \31459 , \3406 );
or \U$31117 ( \31460 , \31458 , \31459 );
nand \U$31118 ( \31461 , \24434 , \3382 );
nand \U$31119 ( \31462 , \31460 , \31461 );
not \U$31120 ( \31463 , \854 );
not \U$31121 ( \31464 , \24377 );
or \U$31122 ( \31465 , \31463 , \31464 );
nand \U$31123 ( \31466 , \31151 , \853 );
nand \U$31124 ( \31467 , \31465 , \31466 );
xor \U$31125 ( \31468 , \31462 , \31467 );
not \U$31126 ( \31469 , \836 );
not \U$31127 ( \31470 , \24457 );
or \U$31128 ( \31471 , \31469 , \31470 );
nand \U$31129 ( \31472 , \831 , \30947 );
nand \U$31130 ( \31473 , \31471 , \31472 );
xor \U$31131 ( \31474 , \31468 , \31473 );
not \U$31132 ( \31475 , \31153 );
not \U$31133 ( \31476 , \31170 );
or \U$31134 ( \31477 , \31475 , \31476 );
or \U$31135 ( \31478 , \31170 , \31153 );
nand \U$31136 ( \31479 , \31478 , \31159 );
nand \U$31137 ( \31480 , \31477 , \31479 );
xor \U$31138 ( \31481 , \31474 , \31480 );
not \U$31139 ( \31482 , \30858 );
not \U$31140 ( \31483 , \30869 );
or \U$31141 ( \31484 , \31482 , \31483 );
or \U$31142 ( \31485 , \30858 , \30869 );
nand \U$31143 ( \31486 , \31485 , \30848 );
nand \U$31144 ( \31487 , \31484 , \31486 );
xnor \U$31145 ( \31488 , \31481 , \31487 );
not \U$31146 ( \31489 , \31488 );
not \U$31147 ( \31490 , \31489 );
not \U$31148 ( \31491 , \31069 );
not \U$31149 ( \31492 , \31053 );
or \U$31150 ( \31493 , \31491 , \31492 );
or \U$31151 ( \31494 , \31069 , \31053 );
nand \U$31152 ( \31495 , \31494 , \31058 );
nand \U$31153 ( \31496 , \31493 , \31495 );
not \U$31154 ( \31497 , \31496 );
not \U$31155 ( \31498 , \31497 );
or \U$31156 ( \31499 , \31490 , \31498 );
or \U$31157 ( \31500 , \31497 , \31489 );
nand \U$31158 ( \31501 , \31499 , \31500 );
or \U$31159 ( \31502 , \31201 , \31192 );
nand \U$31160 ( \31503 , \31502 , \31196 );
nand \U$31161 ( \31504 , \31201 , \31192 );
nand \U$31162 ( \31505 , \31503 , \31504 );
xor \U$31163 ( \31506 , \31501 , \31505 );
not \U$31164 ( \31507 , \31506 );
and \U$31165 ( \31508 , \31457 , \31507 );
not \U$31166 ( \31509 , \31457 );
and \U$31167 ( \31510 , \31509 , \31506 );
nor \U$31168 ( \31511 , \31508 , \31510 );
not \U$31169 ( \31512 , \31511 );
or \U$31170 ( \31513 , \31453 , \31512 );
or \U$31171 ( \31514 , \31511 , \31452 );
nand \U$31172 ( \31515 , \31513 , \31514 );
xor \U$31173 ( \31516 , \31448 , \31515 );
xor \U$31174 ( \31517 , \31095 , \31278 );
and \U$31175 ( \31518 , \31517 , \31283 );
and \U$31176 ( \31519 , \31095 , \31278 );
or \U$31177 ( \31520 , \31518 , \31519 );
xor \U$31178 ( \31521 , \31516 , \31520 );
or \U$31179 ( \31522 , \30974 , \31006 );
nand \U$31180 ( \31523 , \31522 , \31011 );
nand \U$31181 ( \31524 , \31006 , \30974 );
nand \U$31182 ( \31525 , \31523 , \31524 );
xor \U$31183 ( \31526 , \31213 , \31223 );
and \U$31184 ( \31527 , \31526 , \31234 );
and \U$31185 ( \31528 , \31213 , \31223 );
or \U$31186 ( \31529 , \31527 , \31528 );
xor \U$31187 ( \31530 , \31239 , \31249 );
and \U$31188 ( \31531 , \31530 , \31260 );
and \U$31189 ( \31532 , \31239 , \31249 );
or \U$31190 ( \31533 , \31531 , \31532 );
xor \U$31191 ( \31534 , \31529 , \31533 );
xor \U$31192 ( \31535 , \30905 , \30915 );
and \U$31193 ( \31536 , \31535 , \30926 );
and \U$31194 ( \31537 , \30905 , \30915 );
or \U$31195 ( \31538 , \31536 , \31537 );
xor \U$31196 ( \31539 , \31534 , \31538 );
xor \U$31197 ( \31540 , \31525 , \31539 );
buf \U$31198 ( \31541 , \30870 );
or \U$31199 ( \31542 , \30927 , \31541 );
nand \U$31200 ( \31543 , \31542 , \30894 );
nand \U$31201 ( \31544 , \30927 , \31541 );
nand \U$31202 ( \31545 , \31543 , \31544 );
xor \U$31203 ( \31546 , \31540 , \31545 );
not \U$31204 ( \31547 , \31017 );
not \U$31205 ( \31548 , \31023 );
or \U$31206 ( \31549 , \31547 , \31548 );
or \U$31207 ( \31550 , \31023 , \31017 );
nand \U$31208 ( \31551 , \31550 , \31014 );
nand \U$31209 ( \31552 , \31549 , \31551 );
xor \U$31210 ( \31553 , \31546 , \31552 );
not \U$31211 ( \31554 , \31235 );
not \U$31212 ( \31555 , \31266 );
or \U$31213 ( \31556 , \31554 , \31555 );
or \U$31214 ( \31557 , \31235 , \31266 );
nand \U$31215 ( \31558 , \31557 , \31261 );
nand \U$31216 ( \31559 , \31556 , \31558 );
not \U$31217 ( \31560 , \2921 );
not \U$31218 ( \31561 , \30867 );
or \U$31219 ( \31562 , \31560 , \31561 );
nand \U$31220 ( \31563 , \24472 , \2925 );
nand \U$31221 ( \31564 , \31562 , \31563 );
not \U$31222 ( \31565 , \3613 );
not \U$31223 ( \31566 , \24444 );
or \U$31224 ( \31567 , \31565 , \31566 );
nand \U$31225 ( \31568 , \31168 , \2940 );
nand \U$31226 ( \31569 , \31567 , \31568 );
xor \U$31227 ( \31570 , \31564 , \31569 );
not \U$31228 ( \31571 , \3445 );
not \U$31229 ( \31572 , \30844 );
or \U$31230 ( \31573 , \31571 , \31572 );
nand \U$31231 ( \31574 , \24494 , \3465 );
nand \U$31232 ( \31575 , \31573 , \31574 );
xor \U$31233 ( \31576 , \31570 , \31575 );
not \U$31234 ( \31577 , \2963 );
not \U$31235 ( \31578 , \24483 );
or \U$31236 ( \31579 , \31577 , \31578 );
nand \U$31237 ( \31580 , \31155 , \2980 );
nand \U$31238 ( \31581 , \31579 , \31580 );
not \U$31239 ( \31582 , \4075 );
not \U$31240 ( \31583 , RIbb2e710_33);
not \U$31241 ( \31584 , \23399 );
or \U$31242 ( \31585 , \31583 , \31584 );
nand \U$31243 ( \31586 , \7296 , \4785 );
nand \U$31244 ( \31587 , \31585 , \31586 );
not \U$31245 ( \31588 , \31587 );
or \U$31246 ( \31589 , \31582 , \31588 );
nand \U$31247 ( \31590 , \30856 , \3886 );
nand \U$31248 ( \31591 , \31589 , \31590 );
xor \U$31249 ( \31592 , \31581 , \31591 );
not \U$31250 ( \31593 , \7104 );
not \U$31251 ( \31594 , RIbb2e440_39);
not \U$31252 ( \31595 , \13559 );
or \U$31253 ( \31596 , \31594 , \31595 );
not \U$31254 ( \31597 , RIbb2e440_39);
nand \U$31255 ( \31598 , \31597 , \4390 );
nand \U$31256 ( \31599 , \31596 , \31598 );
not \U$31257 ( \31600 , \31599 );
or \U$31258 ( \31601 , \31593 , \31600 );
nand \U$31259 ( \31602 , \31211 , \8445 );
nand \U$31260 ( \31603 , \31601 , \31602 );
not \U$31261 ( \31604 , \31603 );
and \U$31262 ( \31605 , \31592 , \31604 );
not \U$31263 ( \31606 , \31592 );
and \U$31264 ( \31607 , \31606 , \31603 );
nor \U$31265 ( \31608 , \31605 , \31607 );
xor \U$31266 ( \31609 , \31576 , \31608 );
not \U$31267 ( \31610 , \10119 );
not \U$31268 ( \31611 , RIbb2e170_45);
not \U$31269 ( \31612 , \21490 );
or \U$31270 ( \31613 , \31611 , \31612 );
nand \U$31271 ( \31614 , \3653 , \12003 );
nand \U$31272 ( \31615 , \31613 , \31614 );
not \U$31273 ( \31616 , \31615 );
or \U$31274 ( \31617 , \31610 , \31616 );
nand \U$31275 ( \31618 , \30983 , \10117 );
nand \U$31276 ( \31619 , \31617 , \31618 );
not \U$31277 ( \31620 , \11176 );
not \U$31278 ( \31621 , \30901 );
or \U$31279 ( \31622 , \31620 , \31621 );
not \U$31280 ( \31623 , RIbb2e080_47);
not \U$31281 ( \31624 , \3200 );
or \U$31282 ( \31625 , \31623 , \31624 );
nand \U$31283 ( \31626 , \4637 , \16171 );
nand \U$31284 ( \31627 , \31625 , \31626 );
nand \U$31285 ( \31628 , \31627 , \11177 );
nand \U$31286 ( \31629 , \31622 , \31628 );
and \U$31287 ( \31630 , \31619 , \31629 );
not \U$31288 ( \31631 , \31619 );
not \U$31289 ( \31632 , \31629 );
and \U$31290 ( \31633 , \31631 , \31632 );
nor \U$31291 ( \31634 , \31630 , \31633 );
not \U$31292 ( \31635 , \16674 );
not \U$31293 ( \31636 , \30922 );
or \U$31294 ( \31637 , \31635 , \31636 );
not \U$31295 ( \31638 , RIbb2dbd0_57);
not \U$31296 ( \31639 , \20215 );
or \U$31297 ( \31640 , \31638 , \31639 );
nand \U$31298 ( \31641 , \1169 , \17097 );
nand \U$31299 ( \31642 , \31640 , \31641 );
nand \U$31300 ( \31643 , \31642 , \15738 );
nand \U$31301 ( \31644 , \31637 , \31643 );
not \U$31302 ( \31645 , \31644 );
and \U$31303 ( \31646 , \31634 , \31645 );
not \U$31304 ( \31647 , \31634 );
and \U$31305 ( \31648 , \31647 , \31644 );
nor \U$31306 ( \31649 , \31646 , \31648 );
xor \U$31307 ( \31650 , \31609 , \31649 );
xor \U$31308 ( \31651 , \31559 , \31650 );
xor \U$31309 ( \31652 , \30952 , \30962 );
and \U$31310 ( \31653 , \31652 , \30973 );
and \U$31311 ( \31654 , \30952 , \30962 );
or \U$31312 ( \31655 , \31653 , \31654 );
xor \U$31313 ( \31656 , \30985 , \30994 );
and \U$31314 ( \31657 , \31656 , \31005 );
and \U$31315 ( \31658 , \30985 , \30994 );
or \U$31316 ( \31659 , \31657 , \31658 );
xor \U$31317 ( \31660 , \31655 , \31659 );
xor \U$31318 ( \31661 , \23997 , \24004 );
not \U$31319 ( \31662 , \1077 );
not \U$31320 ( \31663 , \24262 );
or \U$31321 ( \31664 , \31662 , \31663 );
nand \U$31322 ( \31665 , \31101 , \1011 );
nand \U$31323 ( \31666 , \31664 , \31665 );
xor \U$31324 ( \31667 , \31661 , \31666 );
not \U$31325 ( \31668 , \998 );
not \U$31326 ( \31669 , \24019 );
or \U$31327 ( \31670 , \31668 , \31669 );
nand \U$31328 ( \31671 , \31113 , \915 );
nand \U$31329 ( \31672 , \31670 , \31671 );
xor \U$31330 ( \31673 , \31667 , \31672 );
not \U$31331 ( \31674 , \20792 );
and \U$31332 ( \31675 , \6229 , \7473 );
not \U$31333 ( \31676 , \6229 );
and \U$31334 ( \31677 , \31676 , RIbb2e530_37);
or \U$31335 ( \31678 , \31675 , \31677 );
not \U$31336 ( \31679 , \31678 );
or \U$31337 ( \31680 , \31674 , \31679 );
nand \U$31338 ( \31681 , \31221 , \6251 );
nand \U$31339 ( \31682 , \31680 , \31681 );
xor \U$31340 ( \31683 , \31673 , \31682 );
not \U$31341 ( \31684 , \4712 );
not \U$31342 ( \31685 , \31247 );
or \U$31343 ( \31686 , \31684 , \31685 );
not \U$31344 ( \31687 , RIbb2e620_35);
not \U$31345 ( \31688 , \8338 );
or \U$31346 ( \31689 , \31687 , \31688 );
nand \U$31347 ( \31690 , \15796 , \5840 );
nand \U$31348 ( \31691 , \31689 , \31690 );
nand \U$31349 ( \31692 , \31691 , \5845 );
nand \U$31350 ( \31693 , \31686 , \31692 );
xor \U$31351 ( \31694 , \31683 , \31693 );
xor \U$31352 ( \31695 , \31660 , \31694 );
xor \U$31353 ( \31696 , \31651 , \31695 );
xor \U$31354 ( \31697 , \31553 , \31696 );
not \U$31355 ( \31698 , \31697 );
xor \U$31356 ( \31699 , \31184 , \31268 );
and \U$31357 ( \31700 , \31699 , \31277 );
and \U$31358 ( \31701 , \31184 , \31268 );
or \U$31359 ( \31702 , \31700 , \31701 );
not \U$31360 ( \31703 , \31702 );
not \U$31361 ( \31704 , \31703 );
or \U$31362 ( \31705 , \31698 , \31704 );
or \U$31363 ( \31706 , \31697 , \31703 );
nand \U$31364 ( \31707 , \31705 , \31706 );
nand \U$31365 ( \31708 , \31039 , \31042 , \31029 );
not \U$31366 ( \31709 , \31708 );
not \U$31367 ( \31710 , \31033 );
or \U$31368 ( \31711 , \31709 , \31710 );
not \U$31369 ( \31712 , \31029 );
nand \U$31370 ( \31713 , \31712 , \31043 );
nand \U$31371 ( \31714 , \31711 , \31713 );
not \U$31372 ( \31715 , \31714 );
and \U$31373 ( \31716 , \31707 , \31715 );
not \U$31374 ( \31717 , \31707 );
and \U$31375 ( \31718 , \31717 , \31714 );
nor \U$31376 ( \31719 , \31716 , \31718 );
xor \U$31377 ( \31720 , \31521 , \31719 );
nand \U$31378 ( \31721 , \31308 , \31720 );
nand \U$31379 ( \31722 , \31303 , \31721 );
nor \U$31380 ( \31723 , \30838 , \31722 );
not \U$31381 ( \31724 , \31723 );
or \U$31382 ( \31725 , \29853 , \31724 );
nand \U$31383 ( \31726 , \30830 , \30835 );
nor \U$31384 ( \31727 , \30827 , \31726 );
nand \U$31385 ( \31728 , \31296 , \31301 );
nand \U$31386 ( \31729 , \30814 , \30826 );
nand \U$31387 ( \31730 , \31728 , \31729 );
nor \U$31388 ( \31731 , \31727 , \31730 );
or \U$31389 ( \31732 , \31731 , \31722 );
not \U$31390 ( \31733 , \31720 );
nand \U$31391 ( \31734 , \31733 , \31307 );
nand \U$31392 ( \31735 , \31732 , \31734 );
not \U$31393 ( \31736 , \31735 );
nand \U$31394 ( \31737 , \31725 , \31736 );
xor \U$31395 ( \31738 , \24358 , \24368 );
xor \U$31396 ( \31739 , \31738 , \24379 );
not \U$31397 ( \31740 , \31629 );
not \U$31398 ( \31741 , \31644 );
or \U$31399 ( \31742 , \31740 , \31741 );
or \U$31400 ( \31743 , \31644 , \31629 );
nand \U$31401 ( \31744 , \31743 , \31619 );
nand \U$31402 ( \31745 , \31742 , \31744 );
xor \U$31403 ( \31746 , \31739 , \31745 );
xor \U$31404 ( \31747 , \31312 , \31322 );
and \U$31405 ( \31748 , \31747 , \31333 );
and \U$31406 ( \31749 , \31312 , \31322 );
or \U$31407 ( \31750 , \31748 , \31749 );
and \U$31408 ( \31751 , \31746 , \31750 );
and \U$31409 ( \31752 , \31739 , \31745 );
or \U$31410 ( \31753 , \31751 , \31752 );
not \U$31411 ( \31754 , \31753 );
xor \U$31412 ( \31755 , \24436 , \24459 );
xor \U$31413 ( \31756 , \31755 , \24447 );
not \U$31414 ( \31757 , \31756 );
not \U$31415 ( \31758 , \31757 );
not \U$31416 ( \31759 , \31603 );
not \U$31417 ( \31760 , \31591 );
or \U$31418 ( \31761 , \31759 , \31760 );
or \U$31419 ( \31762 , \31591 , \31603 );
nand \U$31420 ( \31763 , \31762 , \31581 );
nand \U$31421 ( \31764 , \31761 , \31763 );
not \U$31422 ( \31765 , \31764 );
or \U$31423 ( \31766 , \31758 , \31765 );
or \U$31424 ( \31767 , \31757 , \31764 );
xor \U$31425 ( \31768 , \31673 , \31682 );
and \U$31426 ( \31769 , \31768 , \31693 );
and \U$31427 ( \31770 , \31673 , \31682 );
or \U$31428 ( \31771 , \31769 , \31770 );
nand \U$31429 ( \31772 , \31767 , \31771 );
nand \U$31430 ( \31773 , \31766 , \31772 );
not \U$31431 ( \31774 , \31773 );
xor \U$31432 ( \31775 , \31462 , \31467 );
and \U$31433 ( \31776 , \31775 , \31473 );
and \U$31434 ( \31777 , \31462 , \31467 );
or \U$31435 ( \31778 , \31776 , \31777 );
xor \U$31436 ( \31779 , \31370 , \31375 );
and \U$31437 ( \31780 , \31779 , \31381 );
and \U$31438 ( \31781 , \31370 , \31375 );
or \U$31439 ( \31782 , \31780 , \31781 );
xor \U$31440 ( \31783 , \31778 , \31782 );
xor \U$31441 ( \31784 , \31564 , \31569 );
and \U$31442 ( \31785 , \31784 , \31575 );
and \U$31443 ( \31786 , \31564 , \31569 );
or \U$31444 ( \31787 , \31785 , \31786 );
and \U$31445 ( \31788 , \31783 , \31787 );
and \U$31446 ( \31789 , \31778 , \31782 );
or \U$31447 ( \31790 , \31788 , \31789 );
not \U$31448 ( \31791 , \31790 );
nand \U$31449 ( \31792 , \31774 , \31791 );
not \U$31450 ( \31793 , \31792 );
or \U$31451 ( \31794 , \31754 , \31793 );
nand \U$31452 ( \31795 , \31773 , \31790 );
nand \U$31453 ( \31796 , \31794 , \31795 );
xor \U$31454 ( \31797 , \24425 , \24463 );
xor \U$31455 ( \31798 , \31797 , \24499 );
and \U$31456 ( \31799 , \24296 , \24308 );
not \U$31457 ( \31800 , \24296 );
and \U$31458 ( \31801 , \31800 , \24307 );
nor \U$31459 ( \31802 , \31799 , \31801 );
and \U$31460 ( \31803 , \31802 , \24315 );
not \U$31461 ( \31804 , \31802 );
not \U$31462 ( \31805 , \24315 );
and \U$31463 ( \31806 , \31804 , \31805 );
nor \U$31464 ( \31807 , \31803 , \31806 );
xor \U$31465 ( \31808 , \23930 , \23940 );
xor \U$31466 ( \31809 , \31808 , \23951 );
xor \U$31467 ( \31810 , \31807 , \31809 );
not \U$31468 ( \31811 , \8450 );
not \U$31469 ( \31812 , \24178 );
or \U$31470 ( \31813 , \31811 , \31812 );
nand \U$31471 ( \31814 , \31599 , \8445 );
nand \U$31472 ( \31815 , \31813 , \31814 );
not \U$31473 ( \31816 , \4791 );
not \U$31474 ( \31817 , \23890 );
or \U$31475 ( \31818 , \31816 , \31817 );
nand \U$31476 ( \31819 , \31587 , \3886 );
nand \U$31477 ( \31820 , \31818 , \31819 );
buf \U$31478 ( \31821 , \31820 );
nor \U$31479 ( \31822 , \31815 , \31821 );
not \U$31480 ( \31823 , \6241 );
not \U$31481 ( \31824 , \23938 );
or \U$31482 ( \31825 , \31823 , \31824 );
nand \U$31483 ( \31826 , \31678 , \6250 );
nand \U$31484 ( \31827 , \31825 , \31826 );
not \U$31485 ( \31828 , \31827 );
or \U$31486 ( \31829 , \31822 , \31828 );
nand \U$31487 ( \31830 , \31815 , \31821 );
nand \U$31488 ( \31831 , \31829 , \31830 );
xor \U$31489 ( \31832 , \31810 , \31831 );
xor \U$31490 ( \31833 , \31798 , \31832 );
nor \U$31491 ( \31834 , \31347 , \31364 );
or \U$31492 ( \31835 , \31834 , \31357 );
nand \U$31493 ( \31836 , \31347 , \31364 );
nand \U$31494 ( \31837 , \31835 , \31836 );
not \U$31495 ( \31838 , \31837 );
not \U$31496 ( \31839 , \31838 );
and \U$31497 ( \31840 , \31820 , \31827 );
not \U$31498 ( \31841 , \31820 );
and \U$31499 ( \31842 , \31841 , \31828 );
nor \U$31500 ( \31843 , \31840 , \31842 );
and \U$31501 ( \31844 , \24178 , \8450 );
not \U$31502 ( \31845 , \31599 );
nor \U$31503 ( \31846 , \31845 , \8444 );
nor \U$31504 ( \31847 , \31844 , \31846 );
and \U$31505 ( \31848 , \31843 , \31847 );
not \U$31506 ( \31849 , \31843 );
and \U$31507 ( \31850 , \31849 , \31815 );
nor \U$31508 ( \31851 , \31848 , \31850 );
buf \U$31509 ( \31852 , \31851 );
not \U$31510 ( \31853 , \31852 );
or \U$31511 ( \31854 , \31839 , \31853 );
xor \U$31512 ( \31855 , \31661 , \31666 );
and \U$31513 ( \31856 , \31855 , \31672 );
and \U$31514 ( \31857 , \31661 , \31666 );
or \U$31515 ( \31858 , \31856 , \31857 );
not \U$31516 ( \31859 , \5845 );
not \U$31517 ( \31860 , \23900 );
or \U$31518 ( \31861 , \31859 , \31860 );
nand \U$31519 ( \31862 , \31691 , \4712 );
nand \U$31520 ( \31863 , \31861 , \31862 );
xor \U$31521 ( \31864 , \31858 , \31863 );
not \U$31522 ( \31865 , \16533 );
not \U$31523 ( \31866 , \24102 );
or \U$31524 ( \31867 , \31865 , \31866 );
nand \U$31525 ( \31868 , \31320 , \16541 );
nand \U$31526 ( \31869 , \31867 , \31868 );
xor \U$31527 ( \31870 , \31864 , \31869 );
nand \U$31528 ( \31871 , \31854 , \31870 );
not \U$31529 ( \31872 , \31852 );
not \U$31530 ( \31873 , \31838 );
nand \U$31531 ( \31874 , \31872 , \31873 );
nand \U$31532 ( \31875 , \31871 , \31874 );
and \U$31533 ( \31876 , \31833 , \31875 );
and \U$31534 ( \31877 , \31798 , \31832 );
or \U$31535 ( \31878 , \31876 , \31877 );
buf \U$31536 ( \31879 , \31878 );
xor \U$31537 ( \31880 , \31796 , \31879 );
not \U$31538 ( \31881 , \24087 );
not \U$31539 ( \31882 , \24090 );
or \U$31540 ( \31883 , \31881 , \31882 );
or \U$31541 ( \31884 , \24087 , \24090 );
nand \U$31542 ( \31885 , \31883 , \31884 );
xor \U$31543 ( \31886 , \24118 , \31885 );
not \U$31544 ( \31887 , \9098 );
not \U$31545 ( \31888 , \31420 );
or \U$31546 ( \31889 , \31887 , \31888 );
nand \U$31547 ( \31890 , \24142 , \10451 );
nand \U$31548 ( \31891 , \31889 , \31890 );
not \U$31549 ( \31892 , \31891 );
not \U$31550 ( \31893 , \10119 );
not \U$31551 ( \31894 , \23873 );
or \U$31552 ( \31895 , \31893 , \31894 );
nand \U$31553 ( \31896 , \31615 , \10117 );
nand \U$31554 ( \31897 , \31895 , \31896 );
not \U$31555 ( \31898 , \31897 );
or \U$31556 ( \31899 , \31892 , \31898 );
or \U$31557 ( \31900 , \31891 , \31897 );
not \U$31558 ( \31901 , \14613 );
not \U$31559 ( \31902 , \31430 );
or \U$31560 ( \31903 , \31901 , \31902 );
nand \U$31561 ( \31904 , \24153 , \15181 );
nand \U$31562 ( \31905 , \31903 , \31904 );
nand \U$31563 ( \31906 , \31900 , \31905 );
nand \U$31564 ( \31907 , \31899 , \31906 );
not \U$31565 ( \31908 , \31907 );
xor \U$31566 ( \31909 , \23894 , \23904 );
xor \U$31567 ( \31910 , \31909 , \23916 );
not \U$31568 ( \31911 , \31910 );
or \U$31569 ( \31912 , \31908 , \31911 );
or \U$31570 ( \31913 , \31907 , \31910 );
xor \U$31571 ( \31914 , \24040 , \23968 );
xnor \U$31572 ( \31915 , \31914 , \23979 );
not \U$31573 ( \31916 , \31915 );
nand \U$31574 ( \31917 , \31913 , \31916 );
nand \U$31575 ( \31918 , \31912 , \31917 );
xor \U$31576 ( \31919 , \31886 , \31918 );
not \U$31577 ( \31920 , \23919 );
not \U$31578 ( \31921 , \31920 );
xor \U$31579 ( \31922 , \24042 , \23954 );
not \U$31580 ( \31923 , \31922 );
or \U$31581 ( \31924 , \31921 , \31923 );
or \U$31582 ( \31925 , \31922 , \31920 );
nand \U$31583 ( \31926 , \31924 , \31925 );
xor \U$31584 ( \31927 , \31919 , \31926 );
xor \U$31585 ( \31928 , \31880 , \31927 );
xor \U$31586 ( \31929 , \31798 , \31832 );
xor \U$31587 ( \31930 , \31929 , \31875 );
buf \U$31588 ( \31931 , \31930 );
not \U$31589 ( \31932 , \31931 );
xor \U$31590 ( \31933 , \24474 , \24485 );
xor \U$31591 ( \31934 , \31933 , \24496 );
not \U$31592 ( \31935 , \31934 );
not \U$31593 ( \31936 , \31935 );
not \U$31594 ( \31937 , \31414 );
not \U$31595 ( \31938 , \31435 );
or \U$31596 ( \31939 , \31937 , \31938 );
nand \U$31597 ( \31940 , \31939 , \31424 );
nand \U$31598 ( \31941 , \31434 , \31413 );
nand \U$31599 ( \31942 , \31940 , \31941 );
not \U$31600 ( \31943 , \31942 );
not \U$31601 ( \31944 , \31943 );
or \U$31602 ( \31945 , \31936 , \31944 );
xor \U$31603 ( \31946 , \24005 , \24021 );
xor \U$31604 ( \31947 , \31946 , \24037 );
not \U$31605 ( \31948 , \17275 );
not \U$31606 ( \31949 , \31393 );
or \U$31607 ( \31950 , \31948 , \31949 );
nand \U$31608 ( \31951 , \24390 , RIbb2d888_64);
nand \U$31609 ( \31952 , \31950 , \31951 );
xor \U$31610 ( \31953 , \31947 , \31952 );
not \U$31611 ( \31954 , \12692 );
not \U$31612 ( \31955 , \24166 );
or \U$31613 ( \31956 , \31954 , \31955 );
nand \U$31614 ( \31957 , \31345 , \14067 );
nand \U$31615 ( \31958 , \31956 , \31957 );
xor \U$31616 ( \31959 , \31953 , \31958 );
nand \U$31617 ( \31960 , \31945 , \31959 );
nand \U$31618 ( \31961 , \31942 , \31934 );
nand \U$31619 ( \31962 , \31960 , \31961 );
xor \U$31620 ( \31963 , \31897 , \31905 );
and \U$31621 ( \31964 , \31963 , \31891 );
not \U$31622 ( \31965 , \31963 );
not \U$31623 ( \31966 , \31891 );
and \U$31624 ( \31967 , \31965 , \31966 );
nor \U$31625 ( \31968 , \31964 , \31967 );
not \U$31626 ( \31969 , \31968 );
not \U$31627 ( \31970 , \11177 );
not \U$31628 ( \31971 , \23862 );
or \U$31629 ( \31972 , \31970 , \31971 );
nand \U$31630 ( \31973 , \31627 , \11176 );
nand \U$31631 ( \31974 , \31972 , \31973 );
not \U$31632 ( \31975 , \12284 );
not \U$31633 ( \31976 , \24113 );
or \U$31634 ( \31977 , \31975 , \31976 );
nand \U$31635 ( \31978 , \31329 , \13295 );
nand \U$31636 ( \31979 , \31977 , \31978 );
xor \U$31637 ( \31980 , \31974 , \31979 );
not \U$31638 ( \31981 , \15738 );
not \U$31639 ( \31982 , \23855 );
or \U$31640 ( \31983 , \31981 , \31982 );
nand \U$31641 ( \31984 , \31642 , \16674 );
nand \U$31642 ( \31985 , \31983 , \31984 );
xor \U$31643 ( \31986 , \31980 , \31985 );
not \U$31644 ( \31987 , \31986 );
or \U$31645 ( \31988 , \31969 , \31987 );
or \U$31646 ( \31989 , \31986 , \31968 );
xor \U$31647 ( \31990 , \31382 , \31386 );
and \U$31648 ( \31991 , \31990 , \31397 );
and \U$31649 ( \31992 , \31382 , \31386 );
or \U$31650 ( \31993 , \31991 , \31992 );
nand \U$31651 ( \31994 , \31989 , \31993 );
nand \U$31652 ( \31995 , \31988 , \31994 );
xor \U$31653 ( \31996 , \31962 , \31995 );
xor \U$31654 ( \31997 , \31947 , \31952 );
and \U$31655 ( \31998 , \31997 , \31958 );
and \U$31656 ( \31999 , \31947 , \31952 );
or \U$31657 ( \32000 , \31998 , \31999 );
xor \U$31658 ( \32001 , \31974 , \31979 );
and \U$31659 ( \32002 , \32001 , \31985 );
and \U$31660 ( \32003 , \31974 , \31979 );
or \U$31661 ( \32004 , \32002 , \32003 );
xor \U$31662 ( \32005 , \32000 , \32004 );
not \U$31663 ( \32006 , \16271 );
not \U$31664 ( \32007 , \31362 );
or \U$31665 ( \32008 , \32006 , \32007 );
nand \U$31666 ( \32009 , \24401 , \16257 );
nand \U$31667 ( \32010 , \32008 , \32009 );
not \U$31668 ( \32011 , \8362 );
not \U$31669 ( \32012 , \31409 );
or \U$31670 ( \32013 , \32011 , \32012 );
nand \U$31671 ( \32014 , \24128 , \8353 );
nand \U$31672 ( \32015 , \32013 , \32014 );
xor \U$31673 ( \32016 , \32010 , \32015 );
not \U$31674 ( \32017 , \17563 );
not \U$31675 ( \32018 , \31354 );
or \U$31676 ( \32019 , \32017 , \32018 );
nand \U$31677 ( \32020 , \24196 , \14930 );
nand \U$31678 ( \32021 , \32019 , \32020 );
and \U$31679 ( \32022 , \32016 , \32021 );
and \U$31680 ( \32023 , \32010 , \32015 );
or \U$31681 ( \32024 , \32022 , \32023 );
xor \U$31682 ( \32025 , \32005 , \32024 );
xor \U$31683 ( \32026 , \31996 , \32025 );
not \U$31684 ( \32027 , \32026 );
or \U$31685 ( \32028 , \31932 , \32027 );
or \U$31686 ( \32029 , \32026 , \31931 );
nand \U$31687 ( \32030 , \31608 , \31649 );
and \U$31688 ( \32031 , \32030 , \31576 );
nor \U$31689 ( \32032 , \31649 , \31608 );
nor \U$31690 ( \32033 , \32031 , \32032 );
not \U$31691 ( \32034 , \32033 );
not \U$31692 ( \32035 , \32034 );
xor \U$31693 ( \32036 , \31935 , \31942 );
xor \U$31694 ( \32037 , \32036 , \31959 );
not \U$31695 ( \32038 , \32037 );
not \U$31696 ( \32039 , \32038 );
or \U$31697 ( \32040 , \32035 , \32039 );
not \U$31698 ( \32041 , \32033 );
not \U$31699 ( \32042 , \32037 );
or \U$31700 ( \32043 , \32041 , \32042 );
not \U$31701 ( \32044 , \31340 );
not \U$31702 ( \32045 , \31365 );
or \U$31703 ( \32046 , \32044 , \32045 );
or \U$31704 ( \32047 , \31365 , \31340 );
nand \U$31705 ( \32048 , \32047 , \31334 );
nand \U$31706 ( \32049 , \32046 , \32048 );
nand \U$31707 ( \32050 , \32043 , \32049 );
nand \U$31708 ( \32051 , \32040 , \32050 );
nand \U$31709 ( \32052 , \32029 , \32051 );
nand \U$31710 ( \32053 , \32028 , \32052 );
xor \U$31711 ( \32054 , \31928 , \32053 );
xor \U$31712 ( \32055 , \24283 , \24318 );
xor \U$31713 ( \32056 , \32055 , \24328 );
xor \U$31714 ( \32057 , \31807 , \31809 );
and \U$31715 ( \32058 , \32057 , \31831 );
and \U$31716 ( \32059 , \31807 , \31809 );
or \U$31717 ( \32060 , \32058 , \32059 );
xor \U$31718 ( \32061 , \32056 , \32060 );
or \U$31719 ( \32062 , \32004 , \32024 );
nand \U$31720 ( \32063 , \32062 , \32000 );
nand \U$31721 ( \32064 , \32004 , \32024 );
nand \U$31722 ( \32065 , \32063 , \32064 );
xor \U$31723 ( \32066 , \32061 , \32065 );
xor \U$31724 ( \32067 , \31962 , \31995 );
and \U$31725 ( \32068 , \32067 , \32025 );
and \U$31726 ( \32069 , \31962 , \31995 );
or \U$31727 ( \32070 , \32068 , \32069 );
xor \U$31728 ( \32071 , \32066 , \32070 );
xor \U$31729 ( \32072 , \23846 , \23848 );
xor \U$31730 ( \32073 , \32072 , \23880 );
xor \U$31731 ( \32074 , \31858 , \31863 );
and \U$31732 ( \32075 , \32074 , \31869 );
and \U$31733 ( \32076 , \31858 , \31863 );
or \U$31734 ( \32077 , \32075 , \32076 );
xor \U$31735 ( \32078 , \24382 , \24392 );
xor \U$31736 ( \32079 , \32078 , \24403 );
xor \U$31737 ( \32080 , \32077 , \32079 );
xor \U$31738 ( \32081 , \23877 , \23866 );
xor \U$31739 ( \32082 , \32081 , \23859 );
and \U$31740 ( \32083 , \32080 , \32082 );
and \U$31741 ( \32084 , \32077 , \32079 );
or \U$31742 ( \32085 , \32083 , \32084 );
xor \U$31743 ( \32086 , \32073 , \32085 );
xor \U$31744 ( \32087 , \24094 , \24104 );
xor \U$31745 ( \32088 , \32087 , \24115 );
not \U$31746 ( \32089 , \24198 );
not \U$31747 ( \32090 , \24185 );
or \U$31748 ( \32091 , \32089 , \32090 );
or \U$31749 ( \32092 , \24185 , \24198 );
nand \U$31750 ( \32093 , \32091 , \32092 );
not \U$31751 ( \32094 , \8450 );
not \U$31752 ( \32095 , \23584 );
or \U$31753 ( \32096 , \32094 , \32095 );
nand \U$31754 ( \32097 , \32096 , \24179 );
and \U$31755 ( \32098 , \32093 , \32097 );
not \U$31756 ( \32099 , \32093 );
not \U$31757 ( \32100 , \24182 );
and \U$31758 ( \32101 , \32099 , \32100 );
nor \U$31759 ( \32102 , \32098 , \32101 );
xor \U$31760 ( \32103 , \32088 , \32102 );
not \U$31761 ( \32104 , \24157 );
not \U$31762 ( \32105 , \24133 );
or \U$31763 ( \32106 , \32104 , \32105 );
or \U$31764 ( \32107 , \24157 , \24133 );
nand \U$31765 ( \32108 , \32106 , \32107 );
and \U$31766 ( \32109 , \32108 , \24144 );
not \U$31767 ( \32110 , \32108 );
and \U$31768 ( \32111 , \32110 , \24145 );
nor \U$31769 ( \32112 , \32109 , \32111 );
and \U$31770 ( \32113 , \32103 , \32112 );
and \U$31771 ( \32114 , \32088 , \32102 );
or \U$31772 ( \32115 , \32113 , \32114 );
xor \U$31773 ( \32116 , \32086 , \32115 );
xnor \U$31774 ( \32117 , \32071 , \32116 );
not \U$31775 ( \32118 , \32117 );
xor \U$31776 ( \32119 , \32054 , \32118 );
and \U$31777 ( \32120 , \31838 , \31851 );
not \U$31778 ( \32121 , \31838 );
not \U$31779 ( \32122 , \31851 );
and \U$31780 ( \32123 , \32121 , \32122 );
nor \U$31781 ( \32124 , \32120 , \32123 );
not \U$31782 ( \32125 , \31870 );
and \U$31783 ( \32126 , \32124 , \32125 );
not \U$31784 ( \32127 , \32124 );
and \U$31785 ( \32128 , \32127 , \31870 );
nor \U$31786 ( \32129 , \32126 , \32128 );
not \U$31787 ( \32130 , \32129 );
xor \U$31788 ( \32131 , \31739 , \31745 );
xor \U$31789 ( \32132 , \32131 , \31750 );
or \U$31790 ( \32133 , \32130 , \32132 );
xor \U$31791 ( \32134 , \31398 , \31402 );
and \U$31792 ( \32135 , \32134 , \31436 );
and \U$31793 ( \32136 , \31398 , \31402 );
or \U$31794 ( \32137 , \32135 , \32136 );
nand \U$31795 ( \32138 , \32133 , \32137 );
nand \U$31796 ( \32139 , \32130 , \32132 );
nand \U$31797 ( \32140 , \32138 , \32139 );
not \U$31798 ( \32141 , \31915 );
not \U$31799 ( \32142 , \31910 );
or \U$31800 ( \32143 , \32141 , \32142 );
or \U$31801 ( \32144 , \31910 , \31915 );
nand \U$31802 ( \32145 , \32143 , \32144 );
and \U$31803 ( \32146 , \32145 , \31907 );
not \U$31804 ( \32147 , \32145 );
not \U$31805 ( \32148 , \31907 );
and \U$31806 ( \32149 , \32147 , \32148 );
nor \U$31807 ( \32150 , \32146 , \32149 );
xor \U$31808 ( \32151 , \32010 , \32015 );
xor \U$31809 ( \32152 , \32151 , \32021 );
not \U$31810 ( \32153 , \32152 );
xor \U$31811 ( \32154 , \31778 , \31782 );
xor \U$31812 ( \32155 , \32154 , \31787 );
not \U$31813 ( \32156 , \32155 );
or \U$31814 ( \32157 , \32153 , \32156 );
or \U$31815 ( \32158 , \32155 , \32152 );
buf \U$31816 ( \32159 , \31474 );
or \U$31817 ( \32160 , \32159 , \31480 );
nand \U$31818 ( \32161 , \32160 , \31487 );
nand \U$31819 ( \32162 , \31480 , \32159 );
nand \U$31820 ( \32163 , \32161 , \32162 );
nand \U$31821 ( \32164 , \32158 , \32163 );
nand \U$31822 ( \32165 , \32157 , \32164 );
xor \U$31823 ( \32166 , \32150 , \32165 );
xor \U$31824 ( \32167 , \32088 , \32102 );
xor \U$31825 ( \32168 , \32167 , \32112 );
xor \U$31826 ( \32169 , \32166 , \32168 );
xor \U$31827 ( \32170 , \32140 , \32169 );
not \U$31828 ( \32171 , \31496 );
not \U$31829 ( \32172 , \31489 );
or \U$31830 ( \32173 , \32171 , \32172 );
not \U$31831 ( \32174 , \31497 );
not \U$31832 ( \32175 , \31488 );
or \U$31833 ( \32176 , \32174 , \32175 );
nand \U$31834 ( \32177 , \32176 , \31505 );
nand \U$31835 ( \32178 , \32173 , \32177 );
xor \U$31836 ( \32179 , \32163 , \32152 );
xor \U$31837 ( \32180 , \32179 , \32155 );
or \U$31838 ( \32181 , \32178 , \32180 );
xor \U$31839 ( \32182 , \31993 , \31986 );
xnor \U$31840 ( \32183 , \32182 , \31968 );
not \U$31841 ( \32184 , \32183 );
nand \U$31842 ( \32185 , \32181 , \32184 );
nand \U$31843 ( \32186 , \32178 , \32180 );
nand \U$31844 ( \32187 , \32185 , \32186 );
and \U$31845 ( \32188 , \32170 , \32187 );
and \U$31846 ( \32189 , \32140 , \32169 );
or \U$31847 ( \32190 , \32188 , \32189 );
xor \U$31848 ( \32191 , \32150 , \32165 );
and \U$31849 ( \32192 , \32191 , \32168 );
and \U$31850 ( \32193 , \32150 , \32165 );
or \U$31851 ( \32194 , \32192 , \32193 );
not \U$31852 ( \32195 , \24160 );
not \U$31853 ( \32196 , \24200 );
not \U$31854 ( \32197 , \24205 );
and \U$31855 ( \32198 , \32196 , \32197 );
and \U$31856 ( \32199 , \24205 , \24200 );
nor \U$31857 ( \32200 , \32198 , \32199 );
not \U$31858 ( \32201 , \32200 );
or \U$31859 ( \32202 , \32195 , \32201 );
or \U$31860 ( \32203 , \24160 , \32200 );
nand \U$31861 ( \32204 , \32202 , \32203 );
xor \U$31862 ( \32205 , \24356 , \24406 );
xor \U$31863 ( \32206 , \32205 , \24409 );
xor \U$31864 ( \32207 , \32204 , \32206 );
xor \U$31865 ( \32208 , \24420 , \24422 );
xor \U$31866 ( \32209 , \32208 , \24502 );
xor \U$31867 ( \32210 , \32207 , \32209 );
xor \U$31868 ( \32211 , \32194 , \32210 );
xor \U$31869 ( \32212 , \32077 , \32079 );
xor \U$31870 ( \32213 , \32212 , \32082 );
not \U$31871 ( \32214 , \31753 );
not \U$31872 ( \32215 , \32214 );
not \U$31873 ( \32216 , \31791 );
not \U$31874 ( \32217 , \31773 );
or \U$31875 ( \32218 , \32216 , \32217 );
or \U$31876 ( \32219 , \31773 , \31791 );
nand \U$31877 ( \32220 , \32218 , \32219 );
not \U$31878 ( \32221 , \32220 );
or \U$31879 ( \32222 , \32215 , \32221 );
or \U$31880 ( \32223 , \32214 , \32220 );
nand \U$31881 ( \32224 , \32222 , \32223 );
xor \U$31882 ( \32225 , \32213 , \32224 );
xor \U$31883 ( \32226 , \31529 , \31533 );
and \U$31884 ( \32227 , \32226 , \31538 );
and \U$31885 ( \32228 , \31529 , \31533 );
or \U$31886 ( \32229 , \32227 , \32228 );
xor \U$31887 ( \32230 , \31764 , \31756 );
xnor \U$31888 ( \32231 , \32230 , \31771 );
nor \U$31889 ( \32232 , \32229 , \32231 );
not \U$31890 ( \32233 , \31694 );
not \U$31891 ( \32234 , \31659 );
or \U$31892 ( \32235 , \32233 , \32234 );
or \U$31893 ( \32236 , \31659 , \31694 );
nand \U$31894 ( \32237 , \32236 , \31655 );
nand \U$31895 ( \32238 , \32235 , \32237 );
not \U$31896 ( \32239 , \32238 );
or \U$31897 ( \32240 , \32232 , \32239 );
nand \U$31898 ( \32241 , \32229 , \32231 );
nand \U$31899 ( \32242 , \32240 , \32241 );
and \U$31900 ( \32243 , \32225 , \32242 );
and \U$31901 ( \32244 , \32213 , \32224 );
or \U$31902 ( \32245 , \32243 , \32244 );
xnor \U$31903 ( \32246 , \32211 , \32245 );
xnor \U$31904 ( \32247 , \32190 , \32246 );
not \U$31905 ( \32248 , \32247 );
xor \U$31906 ( \32249 , \31930 , \32051 );
xnor \U$31907 ( \32250 , \32249 , \32026 );
not \U$31908 ( \32251 , \32250 );
not \U$31909 ( \32252 , \32251 );
xor \U$31910 ( \32253 , \32213 , \32224 );
xor \U$31911 ( \32254 , \32253 , \32242 );
not \U$31912 ( \32255 , \32254 );
not \U$31913 ( \32256 , \32255 );
not \U$31914 ( \32257 , \32256 );
or \U$31915 ( \32258 , \32252 , \32257 );
not \U$31916 ( \32259 , \32255 );
not \U$31917 ( \32260 , \32250 );
or \U$31918 ( \32261 , \32259 , \32260 );
or \U$31919 ( \32262 , \31559 , \31650 );
nand \U$31920 ( \32263 , \32262 , \31695 );
nand \U$31921 ( \32264 , \31650 , \31559 );
nand \U$31922 ( \32265 , \32263 , \32264 );
and \U$31923 ( \32266 , \32231 , \32238 );
not \U$31924 ( \32267 , \32231 );
and \U$31925 ( \32268 , \32267 , \32239 );
nor \U$31926 ( \32269 , \32266 , \32268 );
and \U$31927 ( \32270 , \32269 , \32229 );
not \U$31928 ( \32271 , \32269 );
not \U$31929 ( \32272 , \32229 );
and \U$31930 ( \32273 , \32271 , \32272 );
nor \U$31931 ( \32274 , \32270 , \32273 );
xor \U$31932 ( \32275 , \32265 , \32274 );
and \U$31933 ( \32276 , \32049 , \32033 );
not \U$31934 ( \32277 , \32049 );
and \U$31935 ( \32278 , \32277 , \32034 );
or \U$31936 ( \32279 , \32276 , \32278 );
buf \U$31937 ( \32280 , \32037 );
not \U$31938 ( \32281 , \32280 );
and \U$31939 ( \32282 , \32279 , \32281 );
not \U$31940 ( \32283 , \32279 );
and \U$31941 ( \32284 , \32283 , \32280 );
nor \U$31942 ( \32285 , \32282 , \32284 );
and \U$31943 ( \32286 , \32275 , \32285 );
and \U$31944 ( \32287 , \32265 , \32274 );
or \U$31945 ( \32288 , \32286 , \32287 );
nand \U$31946 ( \32289 , \32261 , \32288 );
nand \U$31947 ( \32290 , \32258 , \32289 );
not \U$31948 ( \32291 , \32290 );
not \U$31949 ( \32292 , \32291 );
and \U$31950 ( \32293 , \32248 , \32292 );
and \U$31951 ( \32294 , \32291 , \32247 );
nor \U$31952 ( \32295 , \32293 , \32294 );
xor \U$31953 ( \32296 , \32119 , \32295 );
xor \U$31954 ( \32297 , \32140 , \32169 );
xor \U$31955 ( \32298 , \32297 , \32187 );
buf \U$31956 ( \32299 , \32298 );
not \U$31957 ( \32300 , \32299 );
not \U$31958 ( \32301 , \32132 );
not \U$31959 ( \32302 , \32301 );
not \U$31960 ( \32303 , \32129 );
not \U$31961 ( \32304 , \32303 );
or \U$31962 ( \32305 , \32302 , \32304 );
nand \U$31963 ( \32306 , \32129 , \32132 );
nand \U$31964 ( \32307 , \32305 , \32306 );
not \U$31965 ( \32308 , \32137 );
and \U$31966 ( \32309 , \32307 , \32308 );
not \U$31967 ( \32310 , \32307 );
and \U$31968 ( \32311 , \32310 , \32137 );
nor \U$31969 ( \32312 , \32309 , \32311 );
not \U$31970 ( \32313 , \32312 );
xor \U$31971 ( \32314 , \31525 , \31539 );
and \U$31972 ( \32315 , \32314 , \31545 );
and \U$31973 ( \32316 , \31525 , \31539 );
or \U$31974 ( \32317 , \32315 , \32316 );
or \U$31975 ( \32318 , \32313 , \32317 );
not \U$31976 ( \32319 , \31442 );
not \U$31977 ( \32320 , \31366 );
or \U$31978 ( \32321 , \32319 , \32320 );
or \U$31979 ( \32322 , \31442 , \31366 );
nand \U$31980 ( \32323 , \32322 , \31437 );
nand \U$31981 ( \32324 , \32321 , \32323 );
nand \U$31982 ( \32325 , \32318 , \32324 );
not \U$31983 ( \32326 , \32317 );
not \U$31984 ( \32327 , \32326 );
nand \U$31985 ( \32328 , \32327 , \32313 );
nand \U$31986 ( \32329 , \32325 , \32328 );
not \U$31987 ( \32330 , \32329 );
nand \U$31988 ( \32331 , \32300 , \32330 );
not \U$31989 ( \32332 , \32331 );
not \U$31990 ( \32333 , \32178 );
not \U$31991 ( \32334 , \32183 );
or \U$31992 ( \32335 , \32333 , \32334 );
or \U$31993 ( \32336 , \32178 , \32183 );
nand \U$31994 ( \32337 , \32335 , \32336 );
xor \U$31995 ( \32338 , \32180 , \32337 );
not \U$31996 ( \32339 , \31506 );
not \U$31997 ( \32340 , \31457 );
or \U$31998 ( \32341 , \32339 , \32340 );
or \U$31999 ( \32342 , \31457 , \31506 );
nand \U$32000 ( \32343 , \32342 , \31452 );
nand \U$32001 ( \32344 , \32341 , \32343 );
xor \U$32002 ( \32345 , \32338 , \32344 );
xor \U$32003 ( \32346 , \32265 , \32274 );
xor \U$32004 ( \32347 , \32346 , \32285 );
and \U$32005 ( \32348 , \32345 , \32347 );
and \U$32006 ( \32349 , \32338 , \32344 );
or \U$32007 ( \32350 , \32348 , \32349 );
not \U$32008 ( \32351 , \32350 );
or \U$32009 ( \32352 , \32332 , \32351 );
not \U$32010 ( \32353 , \32330 );
nand \U$32011 ( \32354 , \32353 , \32299 );
nand \U$32012 ( \32355 , \32352 , \32354 );
xor \U$32013 ( \32356 , \32296 , \32355 );
xor \U$32014 ( \32357 , \32254 , \32288 );
xor \U$32015 ( \32358 , \31930 , \32051 );
xor \U$32016 ( \32359 , \32358 , \32026 );
xnor \U$32017 ( \32360 , \32357 , \32359 );
buf \U$32018 ( \32361 , \32360 );
not \U$32019 ( \32362 , \32361 );
and \U$32020 ( \32363 , \32298 , \32330 );
not \U$32021 ( \32364 , \32298 );
and \U$32022 ( \32365 , \32364 , \32329 );
nor \U$32023 ( \32366 , \32363 , \32365 );
not \U$32024 ( \32367 , \32366 );
not \U$32025 ( \32368 , \32367 );
not \U$32026 ( \32369 , \32350 );
not \U$32027 ( \32370 , \32369 );
or \U$32028 ( \32371 , \32368 , \32370 );
nand \U$32029 ( \32372 , \32366 , \32350 );
nand \U$32030 ( \32373 , \32371 , \32372 );
buf \U$32031 ( \32374 , \32373 );
not \U$32032 ( \32375 , \32374 );
not \U$32033 ( \32376 , \32375 );
or \U$32034 ( \32377 , \32362 , \32376 );
xor \U$32035 ( \32378 , \32338 , \32344 );
xor \U$32036 ( \32379 , \32378 , \32347 );
not \U$32037 ( \32380 , \32379 );
xnor \U$32038 ( \32381 , \32317 , \32312 );
xnor \U$32039 ( \32382 , \32381 , \32324 );
buf \U$32040 ( \32383 , \32382 );
xor \U$32041 ( \32384 , \31546 , \31552 );
and \U$32042 ( \32385 , \32384 , \31696 );
and \U$32043 ( \32386 , \31546 , \31552 );
or \U$32044 ( \32387 , \32385 , \32386 );
not \U$32045 ( \32388 , \32387 );
nand \U$32046 ( \32389 , \32383 , \32388 );
not \U$32047 ( \32390 , \32389 );
or \U$32048 ( \32391 , \32380 , \32390 );
or \U$32049 ( \32392 , \32383 , \32388 );
nand \U$32050 ( \32393 , \32391 , \32392 );
not \U$32051 ( \32394 , \32393 );
not \U$32052 ( \32395 , \32394 );
nand \U$32053 ( \32396 , \32377 , \32395 );
not \U$32054 ( \32397 , \32361 );
nand \U$32055 ( \32398 , \32397 , \32374 );
nand \U$32056 ( \32399 , \32396 , \32398 );
not \U$32057 ( \32400 , \32399 );
nand \U$32058 ( \32401 , \32356 , \32400 );
xor \U$32059 ( \32402 , \24044 , \24047 );
xor \U$32060 ( \32403 , \32402 , \23883 );
xor \U$32061 ( \32404 , \24122 , \24208 );
xor \U$32062 ( \32405 , \32404 , \24211 );
xor \U$32063 ( \32406 , \32403 , \32405 );
xor \U$32064 ( \32407 , \24351 , \24353 );
xor \U$32065 ( \32408 , \32407 , \24412 );
xor \U$32066 ( \32409 , \32406 , \32408 );
not \U$32067 ( \32410 , \32409 );
buf \U$32068 ( \32411 , \32410 );
not \U$32069 ( \32412 , \32411 );
buf \U$32070 ( \32413 , \32066 );
not \U$32071 ( \32414 , \32413 );
not \U$32072 ( \32415 , \32116 );
or \U$32073 ( \32416 , \32414 , \32415 );
or \U$32074 ( \32417 , \32116 , \32413 );
nand \U$32075 ( \32418 , \32417 , \32070 );
nand \U$32076 ( \32419 , \32416 , \32418 );
not \U$32077 ( \32420 , \31926 );
not \U$32078 ( \32421 , \31918 );
or \U$32079 ( \32422 , \32420 , \32421 );
or \U$32080 ( \32423 , \31926 , \31918 );
buf \U$32081 ( \32424 , \31886 );
nand \U$32082 ( \32425 , \32423 , \32424 );
nand \U$32083 ( \32426 , \32422 , \32425 );
xor \U$32084 ( \32427 , \32056 , \32060 );
and \U$32085 ( \32428 , \32427 , \32065 );
and \U$32086 ( \32429 , \32056 , \32060 );
or \U$32087 ( \32430 , \32428 , \32429 );
xor \U$32088 ( \32431 , \32426 , \32430 );
not \U$32089 ( \32432 , \32073 );
not \U$32090 ( \32433 , \32115 );
or \U$32091 ( \32434 , \32432 , \32433 );
or \U$32092 ( \32435 , \32115 , \32073 );
nand \U$32093 ( \32436 , \32435 , \32085 );
nand \U$32094 ( \32437 , \32434 , \32436 );
xnor \U$32095 ( \32438 , \32431 , \32437 );
not \U$32096 ( \32439 , \32438 );
xnor \U$32097 ( \32440 , \32419 , \32439 );
not \U$32098 ( \32441 , \32440 );
or \U$32099 ( \32442 , \32412 , \32441 );
not \U$32100 ( \32443 , \32440 );
not \U$32101 ( \32444 , \32411 );
nand \U$32102 ( \32445 , \32443 , \32444 );
nand \U$32103 ( \32446 , \32442 , \32445 );
not \U$32104 ( \32447 , \32118 );
not \U$32105 ( \32448 , \31928 );
or \U$32106 ( \32449 , \32447 , \32448 );
not \U$32107 ( \32450 , \31928 );
not \U$32108 ( \32451 , \32450 );
not \U$32109 ( \32452 , \32117 );
or \U$32110 ( \32453 , \32451 , \32452 );
nand \U$32111 ( \32454 , \32453 , \32053 );
nand \U$32112 ( \32455 , \32449 , \32454 );
not \U$32113 ( \32456 , \32455 );
xor \U$32114 ( \32457 , \32204 , \32206 );
and \U$32115 ( \32458 , \32457 , \32209 );
and \U$32116 ( \32459 , \32204 , \32206 );
or \U$32117 ( \32460 , \32458 , \32459 );
or \U$32118 ( \32461 , \31796 , \31878 );
nand \U$32119 ( \32462 , \32461 , \31927 );
nand \U$32120 ( \32463 , \31878 , \31796 );
nand \U$32121 ( \32464 , \32462 , \32463 );
xor \U$32122 ( \32465 , \32460 , \32464 );
xor \U$32123 ( \32466 , \24505 , \24507 );
xor \U$32124 ( \32467 , \32466 , \24510 );
xor \U$32125 ( \32468 , \32465 , \32467 );
not \U$32126 ( \32469 , \32468 );
or \U$32127 ( \32470 , \32210 , \32194 );
nand \U$32128 ( \32471 , \32470 , \32245 );
nand \U$32129 ( \32472 , \32210 , \32194 );
nand \U$32130 ( \32473 , \32471 , \32472 );
not \U$32131 ( \32474 , \32473 );
not \U$32132 ( \32475 , \32474 );
and \U$32133 ( \32476 , \32469 , \32475 );
and \U$32134 ( \32477 , \32468 , \32474 );
nor \U$32135 ( \32478 , \32476 , \32477 );
not \U$32136 ( \32479 , \32478 );
or \U$32137 ( \32480 , \32456 , \32479 );
not \U$32138 ( \32481 , \32455 );
not \U$32139 ( \32482 , \32478 );
nand \U$32140 ( \32483 , \32481 , \32482 );
nand \U$32141 ( \32484 , \32480 , \32483 );
xor \U$32142 ( \32485 , \32446 , \32484 );
not \U$32143 ( \32486 , \32290 );
buf \U$32144 ( \32487 , \32246 );
not \U$32145 ( \32488 , \32487 );
not \U$32146 ( \32489 , \32488 );
or \U$32147 ( \32490 , \32486 , \32489 );
not \U$32148 ( \32491 , \32487 );
not \U$32149 ( \32492 , \32291 );
or \U$32150 ( \32493 , \32491 , \32492 );
nand \U$32151 ( \32494 , \32493 , \32190 );
nand \U$32152 ( \32495 , \32490 , \32494 );
xnor \U$32153 ( \32496 , \32485 , \32495 );
nand \U$32154 ( \32497 , \32355 , \32119 );
not \U$32155 ( \32498 , \32497 );
not \U$32156 ( \32499 , \32355 );
not \U$32157 ( \32500 , \32119 );
and \U$32158 ( \32501 , \32499 , \32500 );
buf \U$32159 ( \32502 , \32295 );
nor \U$32160 ( \32503 , \32501 , \32502 );
nor \U$32161 ( \32504 , \32498 , \32503 );
nand \U$32162 ( \32505 , \32496 , \32504 );
xor \U$32163 ( \32506 , \32360 , \32373 );
xnor \U$32164 ( \32507 , \32506 , \32394 );
not \U$32165 ( \32508 , \31447 );
buf \U$32166 ( \32509 , \31443 );
not \U$32167 ( \32510 , \32509 );
nand \U$32168 ( \32511 , \32508 , \32510 );
and \U$32169 ( \32512 , \32511 , \31515 );
and \U$32170 ( \32513 , \31447 , \32509 );
nor \U$32171 ( \32514 , \32512 , \32513 );
not \U$32172 ( \32515 , \31702 );
not \U$32173 ( \32516 , \31697 );
or \U$32174 ( \32517 , \32515 , \32516 );
not \U$32175 ( \32518 , \31703 );
not \U$32176 ( \32519 , \31697 );
not \U$32177 ( \32520 , \32519 );
or \U$32178 ( \32521 , \32518 , \32520 );
nand \U$32179 ( \32522 , \32521 , \31714 );
nand \U$32180 ( \32523 , \32517 , \32522 );
not \U$32181 ( \32524 , \32523 );
xor \U$32182 ( \32525 , \32514 , \32524 );
not \U$32183 ( \32526 , \32382 );
not \U$32184 ( \32527 , \32387 );
and \U$32185 ( \32528 , \32526 , \32527 );
and \U$32186 ( \32529 , \32382 , \32387 );
nor \U$32187 ( \32530 , \32528 , \32529 );
not \U$32188 ( \32531 , \32530 );
not \U$32189 ( \32532 , \32379 );
and \U$32190 ( \32533 , \32531 , \32532 );
and \U$32191 ( \32534 , \32379 , \32530 );
nor \U$32192 ( \32535 , \32533 , \32534 );
and \U$32193 ( \32536 , \32525 , \32535 );
and \U$32194 ( \32537 , \32514 , \32524 );
or \U$32195 ( \32538 , \32536 , \32537 );
nand \U$32196 ( \32539 , \32507 , \32538 );
xor \U$32197 ( \32540 , \32514 , \32524 );
xor \U$32198 ( \32541 , \32540 , \32535 );
buf \U$32199 ( \32542 , \32541 );
not \U$32200 ( \32543 , \31516 );
nand \U$32201 ( \32544 , \31719 , \32543 );
and \U$32202 ( \32545 , \32544 , \31520 );
nor \U$32203 ( \32546 , \31719 , \32543 );
nor \U$32204 ( \32547 , \32545 , \32546 );
buf \U$32205 ( \32548 , \32547 );
nand \U$32206 ( \32549 , \32542 , \32548 );
and \U$32207 ( \32550 , \32401 , \32505 , \32539 , \32549 );
nand \U$32208 ( \32551 , \31737 , \32550 );
not \U$32209 ( \32552 , \32551 );
not \U$32210 ( \32553 , \32401 );
nor \U$32211 ( \32554 , \32541 , \32547 );
nand \U$32212 ( \32555 , \32539 , \32554 );
not \U$32213 ( \32556 , \32507 );
not \U$32214 ( \32557 , \32538 );
nand \U$32215 ( \32558 , \32556 , \32557 );
nand \U$32216 ( \32559 , \32555 , \32558 );
not \U$32217 ( \32560 , \32559 );
or \U$32218 ( \32561 , \32553 , \32560 );
not \U$32219 ( \32562 , \32356 );
not \U$32220 ( \32563 , \32400 );
nand \U$32221 ( \32564 , \32562 , \32563 );
nand \U$32222 ( \32565 , \32561 , \32564 );
buf \U$32223 ( \32566 , \32505 );
nand \U$32224 ( \32567 , \32565 , \32566 );
not \U$32225 ( \32568 , \32496 );
not \U$32226 ( \32569 , \32504 );
nand \U$32227 ( \32570 , \32568 , \32569 );
nand \U$32228 ( \32571 , \32567 , \32570 );
not \U$32229 ( \32572 , \32571 );
not \U$32230 ( \32573 , \32572 );
or \U$32231 ( \32574 , \32552 , \32573 );
xor \U$32232 ( \32575 , \24216 , \24219 );
not \U$32233 ( \32576 , \24214 );
xnor \U$32234 ( \32577 , \32575 , \32576 );
buf \U$32235 ( \32578 , \32405 );
not \U$32236 ( \32579 , \32403 );
or \U$32237 ( \32580 , \32578 , \32579 );
nand \U$32238 ( \32581 , \32580 , \32408 );
nand \U$32239 ( \32582 , \32578 , \32579 );
nand \U$32240 ( \32583 , \32581 , \32582 );
xnor \U$32241 ( \32584 , \32577 , \32583 );
xor \U$32242 ( \32585 , \24415 , \24417 );
xor \U$32243 ( \32586 , \32585 , \24513 );
and \U$32244 ( \32587 , \32584 , \32586 );
not \U$32245 ( \32588 , \32584 );
not \U$32246 ( \32589 , \32586 );
and \U$32247 ( \32590 , \32588 , \32589 );
nor \U$32248 ( \32591 , \32587 , \32590 );
xor \U$32249 ( \32592 , \32460 , \32464 );
and \U$32250 ( \32593 , \32592 , \32467 );
and \U$32251 ( \32594 , \32460 , \32464 );
or \U$32252 ( \32595 , \32593 , \32594 );
not \U$32253 ( \32596 , \32595 );
or \U$32254 ( \32597 , \32430 , \32437 );
buf \U$32255 ( \32598 , \32426 );
nand \U$32256 ( \32599 , \32597 , \32598 );
nand \U$32257 ( \32600 , \32437 , \32430 );
nand \U$32258 ( \32601 , \32599 , \32600 );
xor \U$32259 ( \32602 , \24244 , \24339 );
xor \U$32260 ( \32603 , \32602 , \24342 );
not \U$32261 ( \32604 , \32603 );
and \U$32262 ( \32605 , \24056 , \24070 );
not \U$32263 ( \32606 , \24056 );
and \U$32264 ( \32607 , \32606 , \24071 );
nor \U$32265 ( \32608 , \32605 , \32607 );
not \U$32266 ( \32609 , \24053 );
and \U$32267 ( \32610 , \32608 , \32609 );
not \U$32268 ( \32611 , \32608 );
and \U$32269 ( \32612 , \32611 , \24053 );
nor \U$32270 ( \32613 , \32610 , \32612 );
not \U$32271 ( \32614 , \32613 );
or \U$32272 ( \32615 , \32604 , \32614 );
or \U$32273 ( \32616 , \32613 , \32603 );
nand \U$32274 ( \32617 , \32615 , \32616 );
xnor \U$32275 ( \32618 , \32601 , \32617 );
xor \U$32276 ( \32619 , \32596 , \32618 );
not \U$32277 ( \32620 , \32438 );
not \U$32278 ( \32621 , \32409 );
or \U$32279 ( \32622 , \32620 , \32621 );
nand \U$32280 ( \32623 , \32622 , \32419 );
nand \U$32281 ( \32624 , \32410 , \32439 );
nand \U$32282 ( \32625 , \32623 , \32624 );
not \U$32283 ( \32626 , \32625 );
xor \U$32284 ( \32627 , \32619 , \32626 );
xor \U$32285 ( \32628 , \32591 , \32627 );
not \U$32286 ( \32629 , \32455 );
nand \U$32287 ( \32630 , \32629 , \32474 );
buf \U$32288 ( \32631 , \32468 );
and \U$32289 ( \32632 , \32630 , \32631 );
and \U$32290 ( \32633 , \32455 , \32473 );
nor \U$32291 ( \32634 , \32632 , \32633 );
xnor \U$32292 ( \32635 , \32628 , \32634 );
or \U$32293 ( \32636 , \32446 , \32495 );
nand \U$32294 ( \32637 , \32636 , \32484 );
not \U$32295 ( \32638 , \32446 );
not \U$32296 ( \32639 , \32638 );
nand \U$32297 ( \32640 , \32639 , \32495 );
nand \U$32298 ( \32641 , \32637 , \32640 );
not \U$32299 ( \32642 , \32641 );
nand \U$32300 ( \32643 , \32635 , \32642 );
xor \U$32301 ( \32644 , \24348 , \24516 );
buf \U$32302 ( \32645 , \24346 );
not \U$32303 ( \32646 , \32645 );
and \U$32304 ( \32647 , \32644 , \32646 );
not \U$32305 ( \32648 , \32644 );
and \U$32306 ( \32649 , \32648 , \32645 );
nor \U$32307 ( \32650 , \32647 , \32649 );
xor \U$32308 ( \32651 , \24076 , \24083 );
xor \U$32309 ( \32652 , \32651 , \24222 );
not \U$32310 ( \32653 , \32603 );
nand \U$32311 ( \32654 , \32613 , \32653 );
not \U$32312 ( \32655 , \32654 );
not \U$32313 ( \32656 , \32601 );
or \U$32314 ( \32657 , \32655 , \32656 );
or \U$32315 ( \32658 , \32613 , \32653 );
nand \U$32316 ( \32659 , \32657 , \32658 );
xor \U$32317 ( \32660 , \32652 , \32659 );
not \U$32318 ( \32661 , \32577 );
nand \U$32319 ( \32662 , \32661 , \32583 );
not \U$32320 ( \32663 , \32577 );
not \U$32321 ( \32664 , \32583 );
not \U$32322 ( \32665 , \32664 );
or \U$32323 ( \32666 , \32663 , \32665 );
nand \U$32324 ( \32667 , \32666 , \32586 );
nand \U$32325 ( \32668 , \32662 , \32667 );
xor \U$32326 ( \32669 , \32660 , \32668 );
xor \U$32327 ( \32670 , \32650 , \32669 );
xor \U$32328 ( \32671 , \32596 , \32618 );
and \U$32329 ( \32672 , \32671 , \32626 );
and \U$32330 ( \32673 , \32596 , \32618 );
or \U$32331 ( \32674 , \32672 , \32673 );
xor \U$32332 ( \32675 , \32670 , \32674 );
not \U$32333 ( \32676 , \32627 );
not \U$32334 ( \32677 , \32591 );
not \U$32335 ( \32678 , \32677 );
nand \U$32336 ( \32679 , \32676 , \32678 );
not \U$32337 ( \32680 , \32677 );
not \U$32338 ( \32681 , \32627 );
or \U$32339 ( \32682 , \32680 , \32681 );
not \U$32340 ( \32683 , \32634 );
nand \U$32341 ( \32684 , \32682 , \32683 );
nand \U$32342 ( \32685 , \32679 , \32684 );
not \U$32343 ( \32686 , \32685 );
nand \U$32344 ( \32687 , \32675 , \32686 );
xor \U$32345 ( \32688 , \32650 , \32669 );
and \U$32346 ( \32689 , \32688 , \32674 );
and \U$32347 ( \32690 , \32650 , \32669 );
or \U$32348 ( \32691 , \32689 , \32690 );
xor \U$32349 ( \32692 , \24533 , \24526 );
xnor \U$32350 ( \32693 , \32692 , \24537 );
xor \U$32351 ( \32694 , \24225 , \24227 );
xor \U$32352 ( \32695 , \32694 , \24519 );
xor \U$32353 ( \32696 , \32693 , \32695 );
not \U$32354 ( \32697 , \32652 );
not \U$32355 ( \32698 , \32697 );
not \U$32356 ( \32699 , \32659 );
or \U$32357 ( \32700 , \32698 , \32699 );
not \U$32358 ( \32701 , \32652 );
not \U$32359 ( \32702 , \32659 );
not \U$32360 ( \32703 , \32702 );
or \U$32361 ( \32704 , \32701 , \32703 );
nand \U$32362 ( \32705 , \32704 , \32668 );
nand \U$32363 ( \32706 , \32700 , \32705 );
xor \U$32364 ( \32707 , \32696 , \32706 );
nand \U$32365 ( \32708 , \32691 , \32707 );
xor \U$32366 ( \32709 , \24540 , \24522 );
xnor \U$32367 ( \32710 , \32709 , \23843 );
not \U$32368 ( \32711 , \32693 );
not \U$32369 ( \32712 , \32711 );
not \U$32370 ( \32713 , \32706 );
or \U$32371 ( \32714 , \32712 , \32713 );
or \U$32372 ( \32715 , \32706 , \32711 );
buf \U$32373 ( \32716 , \32695 );
nand \U$32374 ( \32717 , \32715 , \32716 );
nand \U$32375 ( \32718 , \32714 , \32717 );
not \U$32376 ( \32719 , \32718 );
nand \U$32377 ( \32720 , \32710 , \32719 );
and \U$32378 ( \32721 , \32643 , \32687 , \32708 , \32720 );
buf \U$32379 ( \32722 , \32721 );
nand \U$32380 ( \32723 , \32574 , \32722 );
buf \U$32381 ( \32724 , \32720 );
not \U$32382 ( \32725 , \32724 );
nand \U$32383 ( \32726 , \32707 , \32691 );
not \U$32384 ( \32727 , \32726 );
not \U$32385 ( \32728 , \32687 );
nor \U$32386 ( \32729 , \32635 , \32642 );
not \U$32387 ( \32730 , \32729 );
or \U$32388 ( \32731 , \32728 , \32730 );
not \U$32389 ( \32732 , \32675 );
not \U$32390 ( \32733 , \32686 );
nand \U$32391 ( \32734 , \32732 , \32733 );
nand \U$32392 ( \32735 , \32731 , \32734 );
not \U$32393 ( \32736 , \32735 );
or \U$32394 ( \32737 , \32727 , \32736 );
or \U$32395 ( \32738 , \32707 , \32691 );
nand \U$32396 ( \32739 , \32737 , \32738 );
not \U$32397 ( \32740 , \32739 );
or \U$32398 ( \32741 , \32725 , \32740 );
or \U$32399 ( \32742 , \32710 , \32719 );
nand \U$32400 ( \32743 , \32741 , \32742 );
not \U$32401 ( \32744 , \32743 );
xor \U$32402 ( \32745 , \28639 , \28651 );
xor \U$32403 ( \32746 , \32745 , \28662 );
xor \U$32404 ( \32747 , \28748 , \28758 );
xor \U$32405 ( \32748 , \32747 , \28769 );
xor \U$32406 ( \32749 , \32746 , \32748 );
xor \U$32407 ( \32750 , \28615 , \28625 );
xor \U$32408 ( \32751 , \32750 , \28636 );
not \U$32409 ( \32752 , \4075 );
not \U$32410 ( \32753 , \28754 );
or \U$32411 ( \32754 , \32752 , \32753 );
not \U$32412 ( \32755 , RIbb2e710_33);
not \U$32413 ( \32756 , \15031 );
or \U$32414 ( \32757 , \32755 , \32756 );
nand \U$32415 ( \32758 , \17682 , \2935 );
nand \U$32416 ( \32759 , \32757 , \32758 );
nand \U$32417 ( \32760 , \32759 , \3887 );
nand \U$32418 ( \32761 , \32754 , \32760 );
xor \U$32419 ( \32762 , \32751 , \32761 );
not \U$32420 ( \32763 , \7104 );
not \U$32421 ( \32764 , \28878 );
or \U$32422 ( \32765 , \32763 , \32764 );
and \U$32423 ( \32766 , RIbb2e440_39, \12323 );
not \U$32424 ( \32767 , RIbb2e440_39);
and \U$32425 ( \32768 , \32767 , \12324 );
or \U$32426 ( \32769 , \32766 , \32768 );
nand \U$32427 ( \32770 , \32769 , \7103 );
nand \U$32428 ( \32771 , \32765 , \32770 );
and \U$32429 ( \32772 , \32762 , \32771 );
and \U$32430 ( \32773 , \32751 , \32761 );
or \U$32431 ( \32774 , \32772 , \32773 );
xor \U$32432 ( \32775 , \32749 , \32774 );
not \U$32433 ( \32776 , \4712 );
not \U$32434 ( \32777 , RIbb2e620_35);
not \U$32435 ( \32778 , \15456 );
or \U$32436 ( \32779 , \32777 , \32778 );
nand \U$32437 ( \32780 , \16320 , \3866 );
nand \U$32438 ( \32781 , \32779 , \32780 );
not \U$32439 ( \32782 , \32781 );
or \U$32440 ( \32783 , \32776 , \32782 );
nand \U$32441 ( \32784 , \28765 , \4714 );
nand \U$32442 ( \32785 , \32783 , \32784 );
not \U$32443 ( \32786 , \6251 );
not \U$32444 ( \32787 , RIbb2e530_37);
not \U$32445 ( \32788 , \13475 );
or \U$32446 ( \32789 , \32787 , \32788 );
nand \U$32447 ( \32790 , \26964 , \7473 );
nand \U$32448 ( \32791 , \32789 , \32790 );
not \U$32449 ( \32792 , \32791 );
or \U$32450 ( \32793 , \32786 , \32792 );
nand \U$32451 ( \32794 , \28658 , \6242 );
nand \U$32452 ( \32795 , \32793 , \32794 );
xor \U$32453 ( \32796 , \32785 , \32795 );
not \U$32454 ( \32797 , \12167 );
not \U$32455 ( \32798 , RIbb2df90_49);
not \U$32456 ( \32799 , \9071 );
or \U$32457 ( \32800 , \32798 , \32799 );
nand \U$32458 ( \32801 , \7299 , \12278 );
nand \U$32459 ( \32802 , \32800 , \32801 );
not \U$32460 ( \32803 , \32802 );
or \U$32461 ( \32804 , \32797 , \32803 );
nand \U$32462 ( \32805 , \28730 , \16427 );
nand \U$32463 ( \32806 , \32804 , \32805 );
and \U$32464 ( \32807 , \32796 , \32806 );
and \U$32465 ( \32808 , \32785 , \32795 );
or \U$32466 ( \32809 , \32807 , \32808 );
xor \U$32467 ( \32810 , \28837 , \28846 );
not \U$32468 ( \32811 , \3465 );
not \U$32469 ( \32812 , \28632 );
or \U$32470 ( \32813 , \32811 , \32812 );
not \U$32471 ( \32814 , RIbb2e9e0_27);
not \U$32472 ( \32815 , \16820 );
or \U$32473 ( \32816 , \32814 , \32815 );
buf \U$32474 ( \32817 , \16818 );
nand \U$32475 ( \32818 , \32817 , \4598 );
nand \U$32476 ( \32819 , \32816 , \32818 );
nand \U$32477 ( \32820 , \32819 , \3445 );
nand \U$32478 ( \32821 , \32813 , \32820 );
xor \U$32479 ( \32822 , \32810 , \32821 );
not \U$32480 ( \32823 , \2925 );
not \U$32481 ( \32824 , \28855 );
or \U$32482 ( \32825 , \32823 , \32824 );
not \U$32483 ( \32826 , RIbb2e8f0_29);
not \U$32484 ( \32827 , \16555 );
or \U$32485 ( \32828 , \32826 , \32827 );
nand \U$32486 ( \32829 , \16706 , \3800 );
nand \U$32487 ( \32830 , \32828 , \32829 );
nand \U$32488 ( \32831 , \32830 , \2922 );
nand \U$32489 ( \32832 , \32825 , \32831 );
and \U$32490 ( \32833 , \32822 , \32832 );
and \U$32491 ( \32834 , \32810 , \32821 );
or \U$32492 ( \32835 , \32833 , \32834 );
not \U$32493 ( \32836 , \8361 );
not \U$32494 ( \32837 , RIbb2e350_41);
not \U$32495 ( \32838 , \11580 );
or \U$32496 ( \32839 , \32837 , \32838 );
not \U$32497 ( \32840 , RIbb2e350_41);
nand \U$32498 ( \32841 , \32840 , \14885 );
nand \U$32499 ( \32842 , \32839 , \32841 );
not \U$32500 ( \32843 , \32842 );
or \U$32501 ( \32844 , \32836 , \32843 );
nand \U$32502 ( \32845 , \28808 , \8354 );
nand \U$32503 ( \32846 , \32844 , \32845 );
xor \U$32504 ( \32847 , \32835 , \32846 );
not \U$32505 ( \32848 , \17563 );
not \U$32506 ( \32849 , RIbb2ddb0_53);
not \U$32507 ( \32850 , \10126 );
or \U$32508 ( \32851 , \32849 , \32850 );
not \U$32509 ( \32852 , \8388 );
nand \U$32510 ( \32853 , \32852 , \12681 );
nand \U$32511 ( \32854 , \32851 , \32853 );
not \U$32512 ( \32855 , \32854 );
or \U$32513 ( \32856 , \32848 , \32855 );
nand \U$32514 ( \32857 , \28887 , \14930 );
nand \U$32515 ( \32858 , \32856 , \32857 );
and \U$32516 ( \32859 , \32847 , \32858 );
and \U$32517 ( \32860 , \32835 , \32846 );
or \U$32518 ( \32861 , \32859 , \32860 );
xor \U$32519 ( \32862 , \32809 , \32861 );
not \U$32520 ( \32863 , \10599 );
not \U$32521 ( \32864 , RIbb2e170_45);
not \U$32522 ( \32865 , \10306 );
or \U$32523 ( \32866 , \32864 , \32865 );
nand \U$32524 ( \32867 , \9841 , \12003 );
nand \U$32525 ( \32868 , \32866 , \32867 );
not \U$32526 ( \32869 , \32868 );
or \U$32527 ( \32870 , \32863 , \32869 );
nand \U$32528 ( \32871 , \28821 , \10119 );
nand \U$32529 ( \32872 , \32870 , \32871 );
not \U$32530 ( \32873 , \12965 );
not \U$32531 ( \32874 , \28718 );
or \U$32532 ( \32875 , \32873 , \32874 );
not \U$32533 ( \32876 , RIbb2e080_47);
not \U$32534 ( \32877 , \12194 );
or \U$32535 ( \32878 , \32876 , \32877 );
nand \U$32536 ( \32879 , \8631 , \10113 );
nand \U$32537 ( \32880 , \32878 , \32879 );
nand \U$32538 ( \32881 , \32880 , \11176 );
nand \U$32539 ( \32882 , \32875 , \32881 );
xor \U$32540 ( \32883 , \32872 , \32882 );
not \U$32541 ( \32884 , \10449 );
not \U$32542 ( \32885 , RIbb2e260_43);
not \U$32543 ( \32886 , \12764 );
or \U$32544 ( \32887 , \32885 , \32886 );
not \U$32545 ( \32888 , \12764 );
nand \U$32546 ( \32889 , \32888 , \9847 );
nand \U$32547 ( \32890 , \32887 , \32889 );
not \U$32548 ( \32891 , \32890 );
or \U$32549 ( \32892 , \32884 , \32891 );
nand \U$32550 ( \32893 , \28797 , \9099 );
nand \U$32551 ( \32894 , \32892 , \32893 );
and \U$32552 ( \32895 , \32883 , \32894 );
and \U$32553 ( \32896 , \32872 , \32882 );
or \U$32554 ( \32897 , \32895 , \32896 );
xor \U$32555 ( \32898 , \32862 , \32897 );
xor \U$32556 ( \32899 , \32775 , \32898 );
xor \U$32557 ( \32900 , \32835 , \32846 );
xor \U$32558 ( \32901 , \32900 , \32858 );
xor \U$32559 ( \32902 , \32872 , \32882 );
xor \U$32560 ( \32903 , \32902 , \32894 );
xor \U$32561 ( \32904 , \32901 , \32903 );
not \U$32562 ( \32905 , \17275 );
not \U$32563 ( \32906 , RIbb2d900_63);
not \U$32564 ( \32907 , \6173 );
or \U$32565 ( \32908 , \32906 , \32907 );
nand \U$32566 ( \32909 , \3228 , \20254 );
nand \U$32567 ( \32910 , \32908 , \32909 );
not \U$32568 ( \32911 , \32910 );
or \U$32569 ( \32912 , \32905 , \32911 );
not \U$32570 ( \32913 , RIbb2d900_63);
not \U$32571 ( \32914 , \3203 );
or \U$32572 ( \32915 , \32913 , \32914 );
nand \U$32573 ( \32916 , \4640 , \17262 );
nand \U$32574 ( \32917 , \32915 , \32916 );
nand \U$32575 ( \32918 , \32917 , RIbb2d888_64);
nand \U$32576 ( \32919 , \32912 , \32918 );
not \U$32577 ( \32920 , \17100 );
not \U$32578 ( \32921 , RIbb2dbd0_57);
not \U$32579 ( \32922 , \4752 );
or \U$32580 ( \32923 , \32921 , \32922 );
nand \U$32581 ( \32924 , \6013 , \17411 );
nand \U$32582 ( \32925 , \32923 , \32924 );
not \U$32583 ( \32926 , \32925 );
or \U$32584 ( \32927 , \32920 , \32926 );
not \U$32585 ( \32928 , RIbb2dbd0_57);
not \U$32586 ( \32929 , \13756 );
or \U$32587 ( \32930 , \32928 , \32929 );
not \U$32588 ( \32931 , RIbb2dbd0_57);
nand \U$32589 ( \32932 , \32931 , \16153 );
nand \U$32590 ( \32933 , \32930 , \32932 );
nand \U$32591 ( \32934 , \32933 , \16675 );
nand \U$32592 ( \32935 , \32927 , \32934 );
nor \U$32593 ( \32936 , \32919 , \32935 );
not \U$32594 ( \32937 , \15181 );
and \U$32595 ( \32938 , RIbb2dcc0_55, \6268 );
not \U$32596 ( \32939 , RIbb2dcc0_55);
and \U$32597 ( \32940 , \32939 , \8375 );
or \U$32598 ( \32941 , \32938 , \32940 );
not \U$32599 ( \32942 , \32941 );
or \U$32600 ( \32943 , \32937 , \32942 );
not \U$32601 ( \32944 , \9023 );
xor \U$32602 ( \32945 , RIbb2dcc0_55, \32944 );
nand \U$32603 ( \32946 , \32945 , \14613 );
nand \U$32604 ( \32947 , \32943 , \32946 );
not \U$32605 ( \32948 , \32947 );
or \U$32606 ( \32949 , \32936 , \32948 );
nand \U$32607 ( \32950 , \32935 , \32919 );
nand \U$32608 ( \32951 , \32949 , \32950 );
and \U$32609 ( \32952 , \32904 , \32951 );
and \U$32610 ( \32953 , \32901 , \32903 );
or \U$32611 ( \32954 , \32952 , \32953 );
xnor \U$32612 ( \32955 , \32899 , \32954 );
not \U$32613 ( \32956 , \32955 );
not \U$32614 ( \32957 , \32956 );
xor \U$32615 ( \32958 , \32751 , \32761 );
xor \U$32616 ( \32959 , \32958 , \32771 );
xor \U$32617 ( \32960 , \32785 , \32795 );
xor \U$32618 ( \32961 , \32960 , \32806 );
xor \U$32619 ( \32962 , \32959 , \32961 );
or \U$32620 ( \32963 , RIbb2e968_28, RIbb2e8f0_29);
nand \U$32621 ( \32964 , \32963 , \17506 );
and \U$32622 ( \32965 , RIbb2e968_28, RIbb2e8f0_29);
nor \U$32623 ( \32966 , \32965 , \3462 );
and \U$32624 ( \32967 , \32964 , \32966 );
not \U$32625 ( \32968 , \3465 );
not \U$32626 ( \32969 , RIbb2e9e0_27);
not \U$32627 ( \32970 , \17745 );
or \U$32628 ( \32971 , \32969 , \32970 );
nand \U$32629 ( \32972 , \17518 , \6065 );
nand \U$32630 ( \32973 , \32971 , \32972 );
not \U$32631 ( \32974 , \32973 );
or \U$32632 ( \32975 , \32968 , \32974 );
or \U$32633 ( \32976 , \19064 , \3462 );
or \U$32634 ( \32977 , \20747 , RIbb2e9e0_27);
nand \U$32635 ( \32978 , \32976 , \32977 );
nand \U$32636 ( \32979 , \32978 , \3444 );
nand \U$32637 ( \32980 , \32975 , \32979 );
and \U$32638 ( \32981 , \32967 , \32980 );
not \U$32639 ( \32982 , \2941 );
not \U$32640 ( \32983 , RIbb2e800_31);
not \U$32641 ( \32984 , \16856 );
not \U$32642 ( \32985 , \32984 );
or \U$32643 ( \32986 , \32983 , \32985 );
not \U$32644 ( \32987 , \32984 );
nand \U$32645 ( \32988 , \32987 , \9169 );
nand \U$32646 ( \32989 , \32986 , \32988 );
not \U$32647 ( \32990 , \32989 );
or \U$32648 ( \32991 , \32982 , \32990 );
not \U$32649 ( \32992 , RIbb2e800_31);
buf \U$32650 ( \32993 , \27577 );
not \U$32651 ( \32994 , \32993 );
or \U$32652 ( \32995 , \32992 , \32994 );
buf \U$32653 ( \32996 , \16829 );
nand \U$32654 ( \32997 , \32996 , \4096 );
nand \U$32655 ( \32998 , \32995 , \32997 );
nand \U$32656 ( \32999 , \32998 , \2939 );
nand \U$32657 ( \33000 , \32991 , \32999 );
xor \U$32658 ( \33001 , \32981 , \33000 );
not \U$32659 ( \33002 , \4790 );
not \U$32660 ( \33003 , RIbb2e710_33);
not \U$32661 ( \33004 , \21665 );
or \U$32662 ( \33005 , \33003 , \33004 );
nand \U$32663 ( \33006 , \23098 , \2935 );
nand \U$32664 ( \33007 , \33005 , \33006 );
not \U$32665 ( \33008 , \33007 );
or \U$32666 ( \33009 , \33002 , \33008 );
not \U$32667 ( \33010 , RIbb2e710_33);
not \U$32668 ( \33011 , \20716 );
or \U$32669 ( \33012 , \33010 , \33011 );
nand \U$32670 ( \33013 , \15825 , \3882 );
nand \U$32671 ( \33014 , \33012 , \33013 );
nand \U$32672 ( \33015 , \33014 , \3886 );
nand \U$32673 ( \33016 , \33009 , \33015 );
and \U$32674 ( \33017 , \33001 , \33016 );
and \U$32675 ( \33018 , \32981 , \33000 );
or \U$32676 ( \33019 , \33017 , \33018 );
not \U$32677 ( \33020 , \10451 );
not \U$32678 ( \33021 , \32890 );
or \U$32679 ( \33022 , \33020 , \33021 );
not \U$32680 ( \33023 , RIbb2e260_43);
not \U$32681 ( \33024 , \16601 );
or \U$32682 ( \33025 , \33023 , \33024 );
not \U$32683 ( \33026 , \17294 );
nand \U$32684 ( \33027 , \33026 , \10444 );
nand \U$32685 ( \33028 , \33025 , \33027 );
nand \U$32686 ( \33029 , \33028 , \9098 );
nand \U$32687 ( \33030 , \33022 , \33029 );
xor \U$32688 ( \33031 , \33019 , \33030 );
not \U$32689 ( \33032 , \10599 );
not \U$32690 ( \33033 , RIbb2e170_45);
not \U$32691 ( \33034 , \12234 );
or \U$32692 ( \33035 , \33033 , \33034 );
nand \U$32693 ( \33036 , \10301 , \12451 );
nand \U$32694 ( \33037 , \33035 , \33036 );
not \U$32695 ( \33038 , \33037 );
or \U$32696 ( \33039 , \33032 , \33038 );
nand \U$32697 ( \33040 , \32868 , \10119 );
nand \U$32698 ( \33041 , \33039 , \33040 );
and \U$32699 ( \33042 , \33031 , \33041 );
and \U$32700 ( \33043 , \33019 , \33030 );
or \U$32701 ( \33044 , \33042 , \33043 );
xor \U$32702 ( \33045 , \32962 , \33044 );
not \U$32703 ( \33046 , \8354 );
not \U$32704 ( \33047 , \32842 );
or \U$32705 ( \33048 , \33046 , \33047 );
not \U$32706 ( \33049 , \22070 );
xor \U$32707 ( \33050 , RIbb2e350_41, \33049 );
nand \U$32708 ( \33051 , \33050 , \8362 );
nand \U$32709 ( \33052 , \33048 , \33051 );
not \U$32710 ( \33053 , \12692 );
and \U$32711 ( \33054 , RIbb2dea0_51, \13876 );
not \U$32712 ( \33055 , RIbb2dea0_51);
and \U$32713 ( \33056 , \33055 , \6604 );
or \U$32714 ( \33057 , \33054 , \33056 );
not \U$32715 ( \33058 , \33057 );
or \U$32716 ( \33059 , \33053 , \33058 );
not \U$32717 ( \33060 , RIbb2dea0_51);
not \U$32718 ( \33061 , \11535 );
or \U$32719 ( \33062 , \33060 , \33061 );
nand \U$32720 ( \33063 , \28728 , \21882 );
nand \U$32721 ( \33064 , \33062 , \33063 );
nand \U$32722 ( \33065 , \33064 , \12774 );
nand \U$32723 ( \33066 , \33059 , \33065 );
xor \U$32724 ( \33067 , \33052 , \33066 );
not \U$32725 ( \33068 , \14930 );
not \U$32726 ( \33069 , \32854 );
or \U$32727 ( \33070 , \33068 , \33069 );
not \U$32728 ( \33071 , RIbb2ddb0_53);
not \U$32729 ( \33072 , \9010 );
or \U$32730 ( \33073 , \33071 , \33072 );
nand \U$32731 ( \33074 , \16952 , \13463 );
nand \U$32732 ( \33075 , \33073 , \33074 );
nand \U$32733 ( \33076 , \33075 , \13467 );
nand \U$32734 ( \33077 , \33070 , \33076 );
and \U$32735 ( \33078 , \33067 , \33077 );
and \U$32736 ( \33079 , \33052 , \33066 );
or \U$32737 ( \33080 , \33078 , \33079 );
xor \U$32738 ( \33081 , \32810 , \32821 );
xor \U$32739 ( \33082 , \33081 , \32832 );
not \U$32740 ( \33083 , \11176 );
not \U$32741 ( \33084 , RIbb2e080_47);
not \U$32742 ( \33085 , \9857 );
or \U$32743 ( \33086 , \33084 , \33085 );
nand \U$32744 ( \33087 , \15128 , \10113 );
nand \U$32745 ( \33088 , \33086 , \33087 );
not \U$32746 ( \33089 , \33088 );
or \U$32747 ( \33090 , \33083 , \33089 );
nand \U$32748 ( \33091 , \32880 , \12965 );
nand \U$32749 ( \33092 , \33090 , \33091 );
xor \U$32750 ( \33093 , \33082 , \33092 );
not \U$32751 ( \33094 , \12285 );
not \U$32752 ( \33095 , \32802 );
or \U$32753 ( \33096 , \33094 , \33095 );
not \U$32754 ( \33097 , RIbb2df90_49);
not \U$32755 ( \33098 , \12801 );
or \U$32756 ( \33099 , \33097 , \33098 );
nand \U$32757 ( \33100 , \9819 , \12278 );
nand \U$32758 ( \33101 , \33099 , \33100 );
nand \U$32759 ( \33102 , \33101 , \12167 );
nand \U$32760 ( \33103 , \33096 , \33102 );
and \U$32761 ( \33104 , \33093 , \33103 );
and \U$32762 ( \33105 , \33082 , \33092 );
or \U$32763 ( \33106 , \33104 , \33105 );
xor \U$32764 ( \33107 , \33080 , \33106 );
not \U$32765 ( \33108 , \15181 );
not \U$32766 ( \33109 , RIbb2dcc0_55);
not \U$32767 ( \33110 , \13756 );
or \U$32768 ( \33111 , \33109 , \33110 );
not \U$32769 ( \33112 , RIbb2dcc0_55);
nand \U$32770 ( \33113 , \33112 , \16153 );
nand \U$32771 ( \33114 , \33111 , \33113 );
not \U$32772 ( \33115 , \33114 );
or \U$32773 ( \33116 , \33108 , \33115 );
nand \U$32774 ( \33117 , \32941 , \14613 );
nand \U$32775 ( \33118 , \33116 , \33117 );
not \U$32776 ( \33119 , \14067 );
not \U$32777 ( \33120 , \33057 );
or \U$32778 ( \33121 , \33119 , \33120 );
and \U$32779 ( \33122 , RIbb2dea0_51, \21570 );
not \U$32780 ( \33123 , RIbb2dea0_51);
and \U$32781 ( \33124 , \33123 , \7308 );
or \U$32782 ( \33125 , \33122 , \33124 );
nand \U$32783 ( \33126 , \33125 , \12692 );
nand \U$32784 ( \33127 , \33121 , \33126 );
xor \U$32785 ( \33128 , \33118 , \33127 );
not \U$32786 ( \33129 , \16675 );
not \U$32787 ( \33130 , \32925 );
or \U$32788 ( \33131 , \33129 , \33130 );
not \U$32789 ( \33132 , RIbb2dbd0_57);
not \U$32790 ( \33133 , \13728 );
or \U$32791 ( \33134 , \33132 , \33133 );
nand \U$32792 ( \33135 , \3002 , \14602 );
nand \U$32793 ( \33136 , \33134 , \33135 );
nand \U$32794 ( \33137 , \33136 , \15738 );
nand \U$32795 ( \33138 , \33131 , \33137 );
xor \U$32796 ( \33139 , \33128 , \33138 );
xor \U$32797 ( \33140 , \33107 , \33139 );
xor \U$32798 ( \33141 , \33045 , \33140 );
xor \U$32799 ( \33142 , \33019 , \33030 );
xor \U$32800 ( \33143 , \33142 , \33041 );
not \U$32801 ( \33144 , \33143 );
not \U$32802 ( \33145 , \33144 );
xor \U$32803 ( \33146 , \32947 , \32935 );
xnor \U$32804 ( \33147 , \33146 , \32919 );
not \U$32805 ( \33148 , \33147 );
or \U$32806 ( \33149 , \33145 , \33148 );
not \U$32807 ( \33150 , \2939 );
not \U$32808 ( \33151 , \32989 );
or \U$32809 ( \33152 , \33150 , \33151 );
nand \U$32810 ( \33153 , \28866 , \3613 );
nand \U$32811 ( \33154 , \33152 , \33153 );
and \U$32812 ( \33155 , \19064 , \2962 );
not \U$32813 ( \33156 , \3465 );
not \U$32814 ( \33157 , \32819 );
or \U$32815 ( \33158 , \33156 , \33157 );
nand \U$32816 ( \33159 , \32973 , \3444 );
nand \U$32817 ( \33160 , \33158 , \33159 );
xor \U$32818 ( \33161 , \33155 , \33160 );
not \U$32819 ( \33162 , \2921 );
not \U$32820 ( \33163 , RIbb2e8f0_29);
not \U$32821 ( \33164 , \27234 );
or \U$32822 ( \33165 , \33163 , \33164 );
nand \U$32823 ( \33166 , \16704 , \3265 );
nand \U$32824 ( \33167 , \33165 , \33166 );
not \U$32825 ( \33168 , \33167 );
or \U$32826 ( \33169 , \33162 , \33168 );
nand \U$32827 ( \33170 , \32830 , \2924 );
nand \U$32828 ( \33171 , \33169 , \33170 );
and \U$32829 ( \33172 , \33161 , \33171 );
and \U$32830 ( \33173 , \33155 , \33160 );
or \U$32831 ( \33174 , \33172 , \33173 );
xor \U$32832 ( \33175 , \33154 , \33174 );
not \U$32833 ( \33176 , \7104 );
not \U$32834 ( \33177 , \32769 );
or \U$32835 ( \33178 , \33176 , \33177 );
and \U$32836 ( \33179 , RIbb2e440_39, \21756 );
not \U$32837 ( \33180 , RIbb2e440_39);
and \U$32838 ( \33181 , \33180 , \27199 );
or \U$32839 ( \33182 , \33179 , \33181 );
nand \U$32840 ( \33183 , \33182 , \7103 );
nand \U$32841 ( \33184 , \33178 , \33183 );
xor \U$32842 ( \33185 , \33175 , \33184 );
not \U$32843 ( \33186 , \16541 );
not \U$32844 ( \33187 , RIbb2d9f0_61);
not \U$32845 ( \33188 , \3023 );
or \U$32846 ( \33189 , \33187 , \33188 );
nand \U$32847 ( \33190 , \8874 , \19746 );
nand \U$32848 ( \33191 , \33189 , \33190 );
not \U$32849 ( \33192 , \33191 );
or \U$32850 ( \33193 , \33186 , \33192 );
not \U$32851 ( \33194 , RIbb2d9f0_61);
not \U$32852 ( \33195 , \7018 );
or \U$32853 ( \33196 , \33194 , \33195 );
nand \U$32854 ( \33197 , \3762 , \19746 );
nand \U$32855 ( \33198 , \33196 , \33197 );
nand \U$32856 ( \33199 , \33198 , \26834 );
nand \U$32857 ( \33200 , \33193 , \33199 );
xor \U$32858 ( \33201 , \33185 , \33200 );
not \U$32859 ( \33202 , \17470 );
and \U$32860 ( \33203 , RIbb2dae0_59, \4029 );
not \U$32861 ( \33204 , RIbb2dae0_59);
and \U$32862 ( \33205 , \33204 , \16180 );
or \U$32863 ( \33206 , \33203 , \33205 );
not \U$32864 ( \33207 , \33206 );
or \U$32865 ( \33208 , \33202 , \33207 );
and \U$32866 ( \33209 , RIbb2dae0_59, \3276 );
not \U$32867 ( \33210 , RIbb2dae0_59);
and \U$32868 ( \33211 , \33210 , \3275 );
or \U$32869 ( \33212 , \33209 , \33211 );
nand \U$32870 ( \33213 , \33212 , \16271 );
nand \U$32871 ( \33214 , \33208 , \33213 );
xor \U$32872 ( \33215 , \33201 , \33214 );
nand \U$32873 ( \33216 , \33149 , \33215 );
not \U$32874 ( \33217 , \33147 );
nand \U$32875 ( \33218 , \33217 , \33143 );
nand \U$32876 ( \33219 , \33216 , \33218 );
and \U$32877 ( \33220 , \33141 , \33219 );
and \U$32878 ( \33221 , \33045 , \33140 );
or \U$32879 ( \33222 , \33220 , \33221 );
not \U$32880 ( \33223 , \33222 );
not \U$32881 ( \33224 , \33223 );
or \U$32882 ( \33225 , \32957 , \33224 );
nand \U$32883 ( \33226 , \33222 , \32955 );
nand \U$32884 ( \33227 , \33225 , \33226 );
and \U$32885 ( \33228 , \28825 , \28801 );
not \U$32886 ( \33229 , \28825 );
not \U$32887 ( \33230 , \28801 );
and \U$32888 ( \33231 , \33229 , \33230 );
nor \U$32889 ( \33232 , \33228 , \33231 );
not \U$32890 ( \33233 , \28812 );
and \U$32891 ( \33234 , \33232 , \33233 );
not \U$32892 ( \33235 , \33232 );
and \U$32893 ( \33236 , \33235 , \28812 );
nor \U$32894 ( \33237 , \33234 , \33236 );
not \U$32895 ( \33238 , \16271 );
not \U$32896 ( \33239 , \33206 );
or \U$32897 ( \33240 , \33238 , \33239 );
and \U$32898 ( \33241 , RIbb2dae0_59, \3023 );
not \U$32899 ( \33242 , RIbb2dae0_59);
and \U$32900 ( \33243 , \33242 , \15444 );
or \U$32901 ( \33244 , \33241 , \33243 );
nand \U$32902 ( \33245 , \33244 , \17470 );
nand \U$32903 ( \33246 , \33240 , \33245 );
not \U$32904 ( \33247 , \33246 );
not \U$32905 ( \33248 , \4075 );
not \U$32906 ( \33249 , \32759 );
or \U$32907 ( \33250 , \33248 , \33249 );
nand \U$32908 ( \33251 , \33007 , \3886 );
nand \U$32909 ( \33252 , \33250 , \33251 );
not \U$32910 ( \33253 , \6241 );
not \U$32911 ( \33254 , \32791 );
or \U$32912 ( \33255 , \33253 , \33254 );
not \U$32913 ( \33256 , RIbb2e530_37);
not \U$32914 ( \33257 , \17315 );
or \U$32915 ( \33258 , \33256 , \33257 );
nand \U$32916 ( \33259 , \13989 , \8701 );
nand \U$32917 ( \33260 , \33258 , \33259 );
nand \U$32918 ( \33261 , \33260 , \6251 );
nand \U$32919 ( \33262 , \33255 , \33261 );
xor \U$32920 ( \33263 , \33252 , \33262 );
not \U$32921 ( \33264 , \4712 );
and \U$32922 ( \33265 , \3866 , \16309 );
not \U$32923 ( \33266 , \3866 );
and \U$32924 ( \33267 , \33266 , \15036 );
nor \U$32925 ( \33268 , \33265 , \33267 );
not \U$32926 ( \33269 , \33268 );
or \U$32927 ( \33270 , \33264 , \33269 );
nand \U$32928 ( \33271 , \32781 , \5845 );
nand \U$32929 ( \33272 , \33270 , \33271 );
and \U$32930 ( \33273 , \33263 , \33272 );
and \U$32931 ( \33274 , \33252 , \33262 );
or \U$32932 ( \33275 , \33273 , \33274 );
not \U$32933 ( \33276 , \33275 );
nand \U$32934 ( \33277 , \33247 , \33276 );
xor \U$32935 ( \33278 , \33154 , \33174 );
and \U$32936 ( \33279 , \33278 , \33184 );
and \U$32937 ( \33280 , \33154 , \33174 );
or \U$32938 ( \33281 , \33279 , \33280 );
and \U$32939 ( \33282 , \33277 , \33281 );
not \U$32940 ( \33283 , \33246 );
nor \U$32941 ( \33284 , \33283 , \33276 );
nor \U$32942 ( \33285 , \33282 , \33284 );
not \U$32943 ( \33286 , \33285 );
xor \U$32944 ( \33287 , \33237 , \33286 );
xor \U$32945 ( \33288 , \28847 , \28857 );
xor \U$32946 ( \33289 , \33288 , \28868 );
not \U$32947 ( \33290 , \17275 );
not \U$32948 ( \33291 , \32917 );
or \U$32949 ( \33292 , \33290 , \33291 );
not \U$32950 ( \33293 , RIbb2d900_63);
not \U$32951 ( \33294 , \15398 );
or \U$32952 ( \33295 , \33293 , \33294 );
not \U$32953 ( \33296 , RIbb2d900_63);
nand \U$32954 ( \33297 , \3146 , \33296 );
nand \U$32955 ( \33298 , \33295 , \33297 );
nand \U$32956 ( \33299 , \33298 , RIbb2d888_64);
nand \U$32957 ( \33300 , \33292 , \33299 );
xor \U$32958 ( \33301 , \33289 , \33300 );
not \U$32959 ( \33302 , \16541 );
not \U$32960 ( \33303 , \33198 );
or \U$32961 ( \33304 , \33302 , \33303 );
not \U$32962 ( \33305 , RIbb2d9f0_61);
not \U$32963 ( \33306 , \6173 );
or \U$32964 ( \33307 , \33305 , \33306 );
nand \U$32965 ( \33308 , \27437 , \21449 );
nand \U$32966 ( \33309 , \33307 , \33308 );
nand \U$32967 ( \33310 , \33309 , \26834 );
nand \U$32968 ( \33311 , \33304 , \33310 );
and \U$32969 ( \33312 , \33301 , \33311 );
and \U$32970 ( \33313 , \33289 , \33300 );
or \U$32971 ( \33314 , \33312 , \33313 );
xnor \U$32972 ( \33315 , \33287 , \33314 );
buf \U$32973 ( \33316 , \33315 );
not \U$32974 ( \33317 , \33316 );
not \U$32975 ( \33318 , \33317 );
xor \U$32976 ( \33319 , \28871 , \28880 );
xor \U$32977 ( \33320 , \33319 , \28891 );
xor \U$32978 ( \33321 , \28712 , \28722 );
xor \U$32979 ( \33322 , \33321 , \28734 );
xor \U$32980 ( \33323 , \33320 , \33322 );
xor \U$32981 ( \33324 , \33118 , \33127 );
and \U$32982 ( \33325 , \33324 , \33138 );
and \U$32983 ( \33326 , \33118 , \33127 );
or \U$32984 ( \33327 , \33325 , \33326 );
not \U$32985 ( \33328 , \33327 );
xor \U$32986 ( \33329 , \33323 , \33328 );
not \U$32987 ( \33330 , \33329 );
not \U$32988 ( \33331 , \33330 );
xor \U$32989 ( \33332 , \33080 , \33106 );
and \U$32990 ( \33333 , \33332 , \33139 );
and \U$32991 ( \33334 , \33080 , \33106 );
or \U$32992 ( \33335 , \33333 , \33334 );
not \U$32993 ( \33336 , \33335 );
not \U$32994 ( \33337 , \33336 );
or \U$32995 ( \33338 , \33331 , \33337 );
nand \U$32996 ( \33339 , \33329 , \33335 );
nand \U$32997 ( \33340 , \33338 , \33339 );
not \U$32998 ( \33341 , \33340 );
or \U$32999 ( \33342 , \33318 , \33341 );
or \U$33000 ( \33343 , \33340 , \33317 );
nand \U$33001 ( \33344 , \33342 , \33343 );
not \U$33002 ( \33345 , \33344 );
and \U$33003 ( \33346 , \33227 , \33345 );
not \U$33004 ( \33347 , \33227 );
and \U$33005 ( \33348 , \33347 , \33344 );
nor \U$33006 ( \33349 , \33346 , \33348 );
xor \U$33007 ( \33350 , \32967 , \32980 );
not \U$33008 ( \33351 , \2924 );
not \U$33009 ( \33352 , \33167 );
or \U$33010 ( \33353 , \33351 , \33352 );
not \U$33011 ( \33354 , RIbb2e8f0_29);
not \U$33012 ( \33355 , \16819 );
or \U$33013 ( \33356 , \33354 , \33355 );
nand \U$33014 ( \33357 , \16818 , \3800 );
nand \U$33015 ( \33358 , \33356 , \33357 );
nand \U$33016 ( \33359 , \33358 , \2921 );
nand \U$33017 ( \33360 , \33353 , \33359 );
xor \U$33018 ( \33361 , \33350 , \33360 );
not \U$33019 ( \33362 , \4790 );
not \U$33020 ( \33363 , \33014 );
or \U$33021 ( \33364 , \33362 , \33363 );
and \U$33022 ( \33365 , \16747 , RIbb2e710_33);
not \U$33023 ( \33366 , \16747 );
and \U$33024 ( \33367 , \33366 , \2935 );
or \U$33025 ( \33368 , \33365 , \33367 );
nand \U$33026 ( \33369 , \33368 , \3886 );
nand \U$33027 ( \33370 , \33364 , \33369 );
and \U$33028 ( \33371 , \33361 , \33370 );
and \U$33029 ( \33372 , \33350 , \33360 );
or \U$33030 ( \33373 , \33371 , \33372 );
not \U$33031 ( \33374 , \10449 );
not \U$33032 ( \33375 , RIbb2e260_43);
not \U$33033 ( \33376 , \11580 );
or \U$33034 ( \33377 , \33375 , \33376 );
nand \U$33035 ( \33378 , \22555 , \8347 );
nand \U$33036 ( \33379 , \33377 , \33378 );
not \U$33037 ( \33380 , \33379 );
or \U$33038 ( \33381 , \33374 , \33380 );
nand \U$33039 ( \33382 , \33028 , \9099 );
nand \U$33040 ( \33383 , \33381 , \33382 );
xor \U$33041 ( \33384 , \33373 , \33383 );
not \U$33042 ( \33385 , \15738 );
not \U$33043 ( \33386 , \32933 );
or \U$33044 ( \33387 , \33385 , \33386 );
not \U$33045 ( \33388 , RIbb2dbd0_57);
not \U$33046 ( \33389 , \6268 );
or \U$33047 ( \33390 , \33388 , \33389 );
nand \U$33048 ( \33391 , \8375 , \14602 );
nand \U$33049 ( \33392 , \33390 , \33391 );
nand \U$33050 ( \33393 , \33392 , \19101 );
nand \U$33051 ( \33394 , \33387 , \33393 );
xnor \U$33052 ( \33395 , \33384 , \33394 );
not \U$33053 ( \33396 , \33395 );
not \U$33054 ( \33397 , \33396 );
not \U$33055 ( \33398 , \12692 );
and \U$33056 ( \33399 , RIbb2dea0_51, \7298 );
not \U$33057 ( \33400 , RIbb2dea0_51);
and \U$33058 ( \33401 , \33400 , \26422 );
or \U$33059 ( \33402 , \33399 , \33401 );
not \U$33060 ( \33403 , \33402 );
or \U$33061 ( \33404 , \33398 , \33403 );
and \U$33062 ( \33405 , RIbb2dea0_51, \27507 );
not \U$33063 ( \33406 , RIbb2dea0_51);
and \U$33064 ( \33407 , \33406 , \14024 );
or \U$33065 ( \33408 , \33405 , \33407 );
nand \U$33066 ( \33409 , \33408 , \12774 );
nand \U$33067 ( \33410 , \33404 , \33409 );
not \U$33068 ( \33411 , \33410 );
not \U$33069 ( \33412 , RIbb2d888_64);
not \U$33070 ( \33413 , RIbb2d900_63);
not \U$33071 ( \33414 , \7018 );
or \U$33072 ( \33415 , \33413 , \33414 );
nand \U$33073 ( \33416 , \3762 , \17262 );
nand \U$33074 ( \33417 , \33415 , \33416 );
not \U$33075 ( \33418 , \33417 );
or \U$33076 ( \33419 , \33412 , \33418 );
not \U$33077 ( \33420 , RIbb2d900_63);
not \U$33078 ( \33421 , \8492 );
or \U$33079 ( \33422 , \33420 , \33421 );
nand \U$33080 ( \33423 , \8491 , \17262 );
nand \U$33081 ( \33424 , \33422 , \33423 );
nand \U$33082 ( \33425 , \33424 , \17275 );
nand \U$33083 ( \33426 , \33419 , \33425 );
not \U$33084 ( \33427 , \33426 );
or \U$33085 ( \33428 , \33411 , \33427 );
or \U$33086 ( \33429 , \33426 , \33410 );
not \U$33087 ( \33430 , \16533 );
not \U$33088 ( \33431 , RIbb2d9f0_61);
not \U$33089 ( \33432 , \13738 );
or \U$33090 ( \33433 , \33431 , \33432 );
nand \U$33091 ( \33434 , \12596 , \16537 );
nand \U$33092 ( \33435 , \33433 , \33434 );
not \U$33093 ( \33436 , \33435 );
or \U$33094 ( \33437 , \33430 , \33436 );
not \U$33095 ( \33438 , RIbb2d9f0_61);
not \U$33096 ( \33439 , \25942 );
or \U$33097 ( \33440 , \33438 , \33439 );
nand \U$33098 ( \33441 , \3002 , \16254 );
nand \U$33099 ( \33442 , \33440 , \33441 );
nand \U$33100 ( \33443 , \33442 , \16541 );
nand \U$33101 ( \33444 , \33437 , \33443 );
nand \U$33102 ( \33445 , \33429 , \33444 );
nand \U$33103 ( \33446 , \33428 , \33445 );
not \U$33104 ( \33447 , \33446 );
or \U$33105 ( \33448 , \33397 , \33447 );
or \U$33106 ( \33449 , \33396 , \33446 );
not \U$33107 ( \33450 , \2941 );
not \U$33108 ( \33451 , \32998 );
or \U$33109 ( \33452 , \33450 , \33451 );
not \U$33110 ( \33453 , RIbb2e800_31);
not \U$33111 ( \33454 , \16555 );
or \U$33112 ( \33455 , \33453 , \33454 );
not \U$33113 ( \33456 , RIbb2e800_31);
nand \U$33114 ( \33457 , \33456 , \16706 );
nand \U$33115 ( \33458 , \33455 , \33457 );
nand \U$33116 ( \33459 , \33458 , \2940 );
nand \U$33117 ( \33460 , \33452 , \33459 );
and \U$33118 ( \33461 , \19064 , \3465 );
not \U$33119 ( \33462 , \2924 );
not \U$33120 ( \33463 , \33358 );
or \U$33121 ( \33464 , \33462 , \33463 );
not \U$33122 ( \33465 , RIbb2e8f0_29);
not \U$33123 ( \33466 , \17745 );
or \U$33124 ( \33467 , \33465 , \33466 );
nand \U$33125 ( \33468 , \26129 , \3800 );
nand \U$33126 ( \33469 , \33467 , \33468 );
nand \U$33127 ( \33470 , \33469 , \2921 );
nand \U$33128 ( \33471 , \33464 , \33470 );
xor \U$33129 ( \33472 , \33461 , \33471 );
not \U$33130 ( \33473 , \2939 );
not \U$33131 ( \33474 , RIbb2e800_31);
not \U$33132 ( \33475 , \17756 );
or \U$33133 ( \33476 , \33474 , \33475 );
not \U$33134 ( \33477 , \17756 );
nand \U$33135 ( \33478 , \33477 , \9169 );
nand \U$33136 ( \33479 , \33476 , \33478 );
not \U$33137 ( \33480 , \33479 );
or \U$33138 ( \33481 , \33473 , \33480 );
nand \U$33139 ( \33482 , \33458 , \2941 );
nand \U$33140 ( \33483 , \33481 , \33482 );
and \U$33141 ( \33484 , \33472 , \33483 );
and \U$33142 ( \33485 , \33461 , \33471 );
or \U$33143 ( \33486 , \33484 , \33485 );
xor \U$33144 ( \33487 , \33460 , \33486 );
not \U$33145 ( \33488 , \8354 );
not \U$33146 ( \33489 , RIbb2e350_41);
not \U$33147 ( \33490 , \12325 );
or \U$33148 ( \33491 , \33489 , \33490 );
nand \U$33149 ( \33492 , \12933 , \8357 );
nand \U$33150 ( \33493 , \33491 , \33492 );
not \U$33151 ( \33494 , \33493 );
or \U$33152 ( \33495 , \33488 , \33494 );
not \U$33153 ( \33496 , RIbb2e350_41);
not \U$33154 ( \33497 , \14844 );
not \U$33155 ( \33498 , \33497 );
or \U$33156 ( \33499 , \33496 , \33498 );
nand \U$33157 ( \33500 , \25984 , \9402 );
nand \U$33158 ( \33501 , \33499 , \33500 );
nand \U$33159 ( \33502 , \33501 , \8362 );
nand \U$33160 ( \33503 , \33495 , \33502 );
xor \U$33161 ( \33504 , \33487 , \33503 );
not \U$33162 ( \33505 , \33504 );
not \U$33163 ( \33506 , \16257 );
xor \U$33164 ( \33507 , RIbb2dae0_59, \10458 );
not \U$33165 ( \33508 , \33507 );
or \U$33166 ( \33509 , \33506 , \33508 );
not \U$33167 ( \33510 , RIbb2dae0_59);
not \U$33168 ( \33511 , \13756 );
or \U$33169 ( \33512 , \33510 , \33511 );
not \U$33170 ( \33513 , RIbb2dae0_59);
nand \U$33171 ( \33514 , \33513 , \4324 );
nand \U$33172 ( \33515 , \33512 , \33514 );
nand \U$33173 ( \33516 , \33515 , \16271 );
nand \U$33174 ( \33517 , \33509 , \33516 );
not \U$33175 ( \33518 , \33517 );
or \U$33176 ( \33519 , \33505 , \33518 );
or \U$33177 ( \33520 , \33517 , \33504 );
xor \U$33178 ( \33521 , \33461 , \33471 );
xor \U$33179 ( \33522 , \33521 , \33483 );
not \U$33180 ( \33523 , \7104 );
and \U$33181 ( \33524 , RIbb2e440_39, \15051 );
not \U$33182 ( \33525 , RIbb2e440_39);
and \U$33183 ( \33526 , \33525 , \15055 );
or \U$33184 ( \33527 , \33524 , \33526 );
not \U$33185 ( \33528 , \33527 );
or \U$33186 ( \33529 , \33523 , \33528 );
and \U$33187 ( \33530 , RIbb2e440_39, \16320 );
not \U$33188 ( \33531 , RIbb2e440_39);
and \U$33189 ( \33532 , \33531 , \14503 );
nor \U$33190 ( \33533 , \33530 , \33532 );
nand \U$33191 ( \33534 , \33533 , \7102 );
nand \U$33192 ( \33535 , \33529 , \33534 );
xor \U$33193 ( \33536 , \33522 , \33535 );
not \U$33194 ( \33537 , \9099 );
not \U$33195 ( \33538 , RIbb2e260_43);
not \U$33196 ( \33539 , \12839 );
or \U$33197 ( \33540 , \33538 , \33539 );
nand \U$33198 ( \33541 , \12175 , \8347 );
nand \U$33199 ( \33542 , \33540 , \33541 );
not \U$33200 ( \33543 , \33542 );
or \U$33201 ( \33544 , \33537 , \33543 );
not \U$33202 ( \33545 , RIbb2e260_43);
not \U$33203 ( \33546 , \12323 );
or \U$33204 ( \33547 , \33545 , \33546 );
nand \U$33205 ( \33548 , \12933 , \17231 );
nand \U$33206 ( \33549 , \33547 , \33548 );
nand \U$33207 ( \33550 , \33549 , \10449 );
nand \U$33208 ( \33551 , \33544 , \33550 );
and \U$33209 ( \33552 , \33536 , \33551 );
and \U$33210 ( \33553 , \33522 , \33535 );
or \U$33211 ( \33554 , \33552 , \33553 );
nand \U$33212 ( \33555 , \33520 , \33554 );
nand \U$33213 ( \33556 , \33519 , \33555 );
nand \U$33214 ( \33557 , \33449 , \33556 );
nand \U$33215 ( \33558 , \33448 , \33557 );
not \U$33216 ( \33559 , \33558 );
xor \U$33217 ( \33560 , \33143 , \33215 );
xnor \U$33218 ( \33561 , \33560 , \33217 );
nand \U$33219 ( \33562 , \33559 , \33561 );
not \U$33220 ( \33563 , \33562 );
xor \U$33221 ( \33564 , \32981 , \33000 );
xor \U$33222 ( \33565 , \33564 , \33016 );
not \U$33223 ( \33566 , RIbb2d888_64);
not \U$33224 ( \33567 , \32910 );
or \U$33225 ( \33568 , \33566 , \33567 );
nand \U$33226 ( \33569 , \33417 , \17275 );
nand \U$33227 ( \33570 , \33568 , \33569 );
xor \U$33228 ( \33571 , \33565 , \33570 );
not \U$33229 ( \33572 , \16271 );
not \U$33230 ( \33573 , \33507 );
or \U$33231 ( \33574 , \33572 , \33573 );
nand \U$33232 ( \33575 , \33212 , \16257 );
nand \U$33233 ( \33576 , \33574 , \33575 );
xnor \U$33234 ( \33577 , \33571 , \33576 );
not \U$33235 ( \33578 , \33577 );
not \U$33236 ( \33579 , \33578 );
xor \U$33237 ( \33580 , \33460 , \33486 );
and \U$33238 ( \33581 , \33580 , \33503 );
and \U$33239 ( \33582 , \33460 , \33486 );
or \U$33240 ( \33583 , \33581 , \33582 );
not \U$33241 ( \33584 , \4714 );
not \U$33242 ( \33585 , RIbb2e620_35);
not \U$33243 ( \33586 , \16783 );
or \U$33244 ( \33587 , \33585 , \33586 );
nand \U$33245 ( \33588 , \15474 , \6002 );
nand \U$33246 ( \33589 , \33587 , \33588 );
not \U$33247 ( \33590 , \33589 );
or \U$33248 ( \33591 , \33584 , \33590 );
not \U$33249 ( \33592 , RIbb2e620_35);
not \U$33250 ( \33593 , \16567 );
or \U$33251 ( \33594 , \33592 , \33593 );
nand \U$33252 ( \33595 , \16566 , \6002 );
nand \U$33253 ( \33596 , \33594 , \33595 );
nand \U$33254 ( \33597 , \33596 , \4712 );
nand \U$33255 ( \33598 , \33591 , \33597 );
not \U$33256 ( \33599 , \7103 );
not \U$33257 ( \33600 , \33527 );
or \U$33258 ( \33601 , \33599 , \33600 );
and \U$33259 ( \33602 , RIbb2e440_39, \13475 );
not \U$33260 ( \33603 , RIbb2e440_39);
and \U$33261 ( \33604 , \33603 , \13474 );
or \U$33262 ( \33605 , \33602 , \33604 );
nand \U$33263 ( \33606 , \33605 , \7104 );
nand \U$33264 ( \33607 , \33601 , \33606 );
xor \U$33265 ( \33608 , \33598 , \33607 );
not \U$33266 ( \33609 , \6251 );
not \U$33267 ( \33610 , RIbb2e530_37);
not \U$33268 ( \33611 , \14528 );
or \U$33269 ( \33612 , \33610 , \33611 );
nand \U$33270 ( \33613 , \14527 , \4708 );
nand \U$33271 ( \33614 , \33612 , \33613 );
not \U$33272 ( \33615 , \33614 );
or \U$33273 ( \33616 , \33609 , \33615 );
not \U$33274 ( \33617 , RIbb2e530_37);
not \U$33275 ( \33618 , \15456 );
or \U$33276 ( \33619 , \33617 , \33618 );
nand \U$33277 ( \33620 , \16320 , \4708 );
nand \U$33278 ( \33621 , \33619 , \33620 );
nand \U$33279 ( \33622 , \33621 , \6242 );
nand \U$33280 ( \33623 , \33616 , \33622 );
and \U$33281 ( \33624 , \33608 , \33623 );
and \U$33282 ( \33625 , \33598 , \33607 );
or \U$33283 ( \33626 , \33624 , \33625 );
xor \U$33284 ( \33627 , \33583 , \33626 );
xor \U$33285 ( \33628 , \33350 , \33360 );
xor \U$33286 ( \33629 , \33628 , \33370 );
not \U$33287 ( \33630 , \14613 );
and \U$33288 ( \33631 , RIbb2dcc0_55, \10577 );
not \U$33289 ( \33632 , RIbb2dcc0_55);
and \U$33290 ( \33633 , \33632 , \5955 );
or \U$33291 ( \33634 , \33631 , \33633 );
not \U$33292 ( \33635 , \33634 );
or \U$33293 ( \33636 , \33630 , \33635 );
and \U$33294 ( \33637 , RIbb2dcc0_55, \9109 );
not \U$33295 ( \33638 , RIbb2dcc0_55);
and \U$33296 ( \33639 , \33638 , \8387 );
or \U$33297 ( \33640 , \33637 , \33639 );
nand \U$33298 ( \33641 , \33640 , \15181 );
nand \U$33299 ( \33642 , \33636 , \33641 );
xor \U$33300 ( \33643 , \33629 , \33642 );
not \U$33301 ( \33644 , \12167 );
not \U$33302 ( \33645 , RIbb2df90_49);
not \U$33303 ( \33646 , \9857 );
or \U$33304 ( \33647 , \33645 , \33646 );
nand \U$33305 ( \33648 , \15128 , \12278 );
nand \U$33306 ( \33649 , \33647 , \33648 );
not \U$33307 ( \33650 , \33649 );
or \U$33308 ( \33651 , \33644 , \33650 );
not \U$33309 ( \33652 , RIbb2df90_49);
not \U$33310 ( \33653 , \12194 );
or \U$33311 ( \33654 , \33652 , \33653 );
nand \U$33312 ( \33655 , \8631 , \12278 );
nand \U$33313 ( \33656 , \33654 , \33655 );
nand \U$33314 ( \33657 , \33656 , \12169 );
nand \U$33315 ( \33658 , \33651 , \33657 );
and \U$33316 ( \33659 , \33643 , \33658 );
and \U$33317 ( \33660 , \33629 , \33642 );
or \U$33318 ( \33661 , \33659 , \33660 );
xor \U$33319 ( \33662 , \33627 , \33661 );
not \U$33320 ( \33663 , \33662 );
or \U$33321 ( \33664 , \33579 , \33663 );
or \U$33322 ( \33665 , \33578 , \33662 );
not \U$33323 ( \33666 , \8353 );
not \U$33324 ( \33667 , \33501 );
or \U$33325 ( \33668 , \33666 , \33667 );
not \U$33326 ( \33669 , RIbb2e350_41);
not \U$33327 ( \33670 , \18857 );
or \U$33328 ( \33671 , \33669 , \33670 );
nand \U$33329 ( \33672 , \28391 , \7097 );
nand \U$33330 ( \33673 , \33671 , \33672 );
nand \U$33331 ( \33674 , \33673 , \8362 );
nand \U$33332 ( \33675 , \33668 , \33674 );
not \U$33333 ( \33676 , \6242 );
not \U$33334 ( \33677 , \33614 );
or \U$33335 ( \33678 , \33676 , \33677 );
not \U$33336 ( \33679 , RIbb2e530_37);
not \U$33337 ( \33680 , \16783 );
or \U$33338 ( \33681 , \33679 , \33680 );
nand \U$33339 ( \33682 , \15470 , \6246 );
nand \U$33340 ( \33683 , \33681 , \33682 );
nand \U$33341 ( \33684 , \33683 , \6251 );
nand \U$33342 ( \33685 , \33678 , \33684 );
xor \U$33343 ( \33686 , \33675 , \33685 );
not \U$33344 ( \33687 , \12167 );
not \U$33345 ( \33688 , RIbb2df90_49);
not \U$33346 ( \33689 , \22580 );
or \U$33347 ( \33690 , \33688 , \33689 );
nand \U$33348 ( \33691 , \9841 , \12278 );
nand \U$33349 ( \33692 , \33690 , \33691 );
not \U$33350 ( \33693 , \33692 );
or \U$33351 ( \33694 , \33687 , \33693 );
nand \U$33352 ( \33695 , \33649 , \16427 );
nand \U$33353 ( \33696 , \33694 , \33695 );
and \U$33354 ( \33697 , \33686 , \33696 );
and \U$33355 ( \33698 , \33675 , \33685 );
or \U$33356 ( \33699 , \33697 , \33698 );
not \U$33357 ( \33700 , \33699 );
not \U$33358 ( \33701 , \16674 );
not \U$33359 ( \33702 , RIbb2dbd0_57);
not \U$33360 ( \33703 , \9108 );
or \U$33361 ( \33704 , \33702 , \33703 );
not \U$33362 ( \33705 , RIbb2dbd0_57);
nand \U$33363 ( \33706 , \33705 , \8387 );
nand \U$33364 ( \33707 , \33704 , \33706 );
not \U$33365 ( \33708 , \33707 );
or \U$33366 ( \33709 , \33701 , \33708 );
not \U$33367 ( \33710 , RIbb2dbd0_57);
not \U$33368 ( \33711 , \9021 );
or \U$33369 ( \33712 , \33710 , \33711 );
nand \U$33370 ( \33713 , \18623 , \15741 );
nand \U$33371 ( \33714 , \33712 , \33713 );
nand \U$33372 ( \33715 , \33714 , \15738 );
nand \U$33373 ( \33716 , \33709 , \33715 );
not \U$33374 ( \33717 , \16257 );
not \U$33375 ( \33718 , \33515 );
or \U$33376 ( \33719 , \33717 , \33718 );
not \U$33377 ( \33720 , RIbb2dae0_59);
not \U$33378 ( \33721 , \6268 );
or \U$33379 ( \33722 , \33720 , \33721 );
not \U$33380 ( \33723 , RIbb2dae0_59);
nand \U$33381 ( \33724 , \33723 , \4391 );
nand \U$33382 ( \33725 , \33722 , \33724 );
nand \U$33383 ( \33726 , \33725 , \16271 );
nand \U$33384 ( \33727 , \33719 , \33726 );
xor \U$33385 ( \33728 , \33716 , \33727 );
not \U$33386 ( \33729 , \11177 );
not \U$33387 ( \33730 , RIbb2e080_47);
not \U$33388 ( \33731 , \13929 );
or \U$33389 ( \33732 , \33730 , \33731 );
nand \U$33390 ( \33733 , \10300 , \12971 );
nand \U$33391 ( \33734 , \33732 , \33733 );
not \U$33392 ( \33735 , \33734 );
or \U$33393 ( \33736 , \33729 , \33735 );
not \U$33394 ( \33737 , RIbb2e080_47);
not \U$33395 ( \33738 , \12764 );
or \U$33396 ( \33739 , \33737 , \33738 );
nand \U$33397 ( \33740 , \13525 , \10113 );
nand \U$33398 ( \33741 , \33739 , \33740 );
nand \U$33399 ( \33742 , \33741 , \11176 );
nand \U$33400 ( \33743 , \33736 , \33742 );
and \U$33401 ( \33744 , \33728 , \33743 );
and \U$33402 ( \33745 , \33716 , \33727 );
or \U$33403 ( \33746 , \33744 , \33745 );
not \U$33404 ( \33747 , \33746 );
or \U$33405 ( \33748 , \33700 , \33747 );
or \U$33406 ( \33749 , \33699 , \33746 );
or \U$33407 ( \33750 , RIbb2e878_30, RIbb2e800_31);
nand \U$33408 ( \33751 , \33750 , \17506 );
and \U$33409 ( \33752 , RIbb2e878_30, RIbb2e800_31);
nor \U$33410 ( \33753 , \33752 , \3800 );
and \U$33411 ( \33754 , \33751 , \33753 );
not \U$33412 ( \33755 , \2924 );
not \U$33413 ( \33756 , \33469 );
or \U$33414 ( \33757 , \33755 , \33756 );
and \U$33415 ( \33758 , RIbb2e8f0_29, \17506 );
not \U$33416 ( \33759 , RIbb2e8f0_29);
and \U$33417 ( \33760 , \33759 , \19063 );
nor \U$33418 ( \33761 , \33758 , \33760 );
nand \U$33419 ( \33762 , \33761 , \2921 );
nand \U$33420 ( \33763 , \33757 , \33762 );
xor \U$33421 ( \33764 , \33754 , \33763 );
not \U$33422 ( \33765 , \2941 );
not \U$33423 ( \33766 , \33479 );
or \U$33424 ( \33767 , \33765 , \33766 );
not \U$33425 ( \33768 , RIbb2e800_31);
not \U$33426 ( \33769 , \16820 );
or \U$33427 ( \33770 , \33768 , \33769 );
nand \U$33428 ( \33771 , \17529 , \2917 );
nand \U$33429 ( \33772 , \33770 , \33771 );
nand \U$33430 ( \33773 , \33772 , \2939 );
nand \U$33431 ( \33774 , \33767 , \33773 );
xor \U$33432 ( \33775 , \33764 , \33774 );
not \U$33433 ( \33776 , \4714 );
not \U$33434 ( \33777 , RIbb2e620_35);
not \U$33435 ( \33778 , \16844 );
or \U$33436 ( \33779 , \33777 , \33778 );
nand \U$33437 ( \33780 , \16576 , \6002 );
nand \U$33438 ( \33781 , \33779 , \33780 );
not \U$33439 ( \33782 , \33781 );
or \U$33440 ( \33783 , \33776 , \33782 );
not \U$33441 ( \33784 , RIbb2e620_35);
not \U$33442 ( \33785 , \16747 );
or \U$33443 ( \33786 , \33784 , \33785 );
nand \U$33444 ( \33787 , \19077 , \3866 );
nand \U$33445 ( \33788 , \33786 , \33787 );
nand \U$33446 ( \33789 , \33788 , \4712 );
nand \U$33447 ( \33790 , \33783 , \33789 );
and \U$33448 ( \33791 , \33775 , \33790 );
and \U$33449 ( \33792 , \33764 , \33774 );
or \U$33450 ( \33793 , \33791 , \33792 );
not \U$33451 ( \33794 , \15182 );
not \U$33452 ( \33795 , \33634 );
or \U$33453 ( \33796 , \33794 , \33795 );
and \U$33454 ( \33797 , RIbb2dcc0_55, \9057 );
not \U$33455 ( \33798 , RIbb2dcc0_55);
and \U$33456 ( \33799 , \33798 , \26467 );
or \U$33457 ( \33800 , \33797 , \33799 );
nand \U$33458 ( \33801 , \33800 , \14613 );
nand \U$33459 ( \33802 , \33796 , \33801 );
xor \U$33460 ( \33803 , \33793 , \33802 );
not \U$33461 ( \33804 , \10119 );
not \U$33462 ( \33805 , RIbb2e170_45);
not \U$33463 ( \33806 , \16601 );
or \U$33464 ( \33807 , \33805 , \33806 );
nand \U$33465 ( \33808 , \16604 , \12451 );
nand \U$33466 ( \33809 , \33807 , \33808 );
not \U$33467 ( \33810 , \33809 );
or \U$33468 ( \33811 , \33804 , \33810 );
not \U$33469 ( \33812 , RIbb2e170_45);
not \U$33470 ( \33813 , \14886 );
or \U$33471 ( \33814 , \33812 , \33813 );
nand \U$33472 ( \33815 , \22555 , \12003 );
nand \U$33473 ( \33816 , \33814 , \33815 );
nand \U$33474 ( \33817 , \33816 , \10117 );
nand \U$33475 ( \33818 , \33811 , \33817 );
and \U$33476 ( \33819 , \33803 , \33818 );
and \U$33477 ( \33820 , \33793 , \33802 );
or \U$33478 ( \33821 , \33819 , \33820 );
nand \U$33479 ( \33822 , \33749 , \33821 );
nand \U$33480 ( \33823 , \33748 , \33822 );
nand \U$33481 ( \33824 , \33665 , \33823 );
nand \U$33482 ( \33825 , \33664 , \33824 );
not \U$33483 ( \33826 , \33825 );
or \U$33484 ( \33827 , \33563 , \33826 );
not \U$33485 ( \33828 , \33561 );
nand \U$33486 ( \33829 , \33828 , \33558 );
nand \U$33487 ( \33830 , \33827 , \33829 );
not \U$33488 ( \33831 , \33830 );
xor \U$33489 ( \33832 , \32901 , \32903 );
xor \U$33490 ( \33833 , \33832 , \32951 );
xor \U$33491 ( \33834 , \33252 , \33262 );
xor \U$33492 ( \33835 , \33834 , \33272 );
not \U$33493 ( \33836 , \33835 );
not \U$33494 ( \33837 , \6251 );
not \U$33495 ( \33838 , \33621 );
or \U$33496 ( \33839 , \33837 , \33838 );
nand \U$33497 ( \33840 , \33260 , \6242 );
nand \U$33498 ( \33841 , \33839 , \33840 );
not \U$33499 ( \33842 , \33841 );
not \U$33500 ( \33843 , \4712 );
not \U$33501 ( \33844 , \33589 );
or \U$33502 ( \33845 , \33843 , \33844 );
nand \U$33503 ( \33846 , \5845 , \33268 );
nand \U$33504 ( \33847 , \33845 , \33846 );
not \U$33505 ( \33848 , \33847 );
nand \U$33506 ( \33849 , \33842 , \33848 );
not \U$33507 ( \33850 , \33849 );
not \U$33508 ( \33851 , \15181 );
not \U$33509 ( \33852 , \32945 );
or \U$33510 ( \33853 , \33851 , \33852 );
nand \U$33511 ( \33854 , \33640 , \14613 );
nand \U$33512 ( \33855 , \33853 , \33854 );
not \U$33513 ( \33856 , \33855 );
or \U$33514 ( \33857 , \33850 , \33856 );
nand \U$33515 ( \33858 , \33847 , \33841 );
nand \U$33516 ( \33859 , \33857 , \33858 );
not \U$33517 ( \33860 , \33859 );
or \U$33518 ( \33861 , \33836 , \33860 );
or \U$33519 ( \33862 , \33859 , \33835 );
xor \U$33520 ( \33863 , \33155 , \33160 );
xor \U$33521 ( \33864 , \33863 , \33171 );
not \U$33522 ( \33865 , \7103 );
not \U$33523 ( \33866 , \33605 );
or \U$33524 ( \33867 , \33865 , \33866 );
nand \U$33525 ( \33868 , \33182 , \7104 );
nand \U$33526 ( \33869 , \33867 , \33868 );
xor \U$33527 ( \33870 , \33864 , \33869 );
not \U$33528 ( \33871 , \8354 );
not \U$33529 ( \33872 , \33050 );
or \U$33530 ( \33873 , \33871 , \33872 );
nand \U$33531 ( \33874 , \33493 , \8362 );
nand \U$33532 ( \33875 , \33873 , \33874 );
and \U$33533 ( \33876 , \33870 , \33875 );
and \U$33534 ( \33877 , \33864 , \33869 );
or \U$33535 ( \33878 , \33876 , \33877 );
nand \U$33536 ( \33879 , \33862 , \33878 );
nand \U$33537 ( \33880 , \33861 , \33879 );
xor \U$33538 ( \33881 , \33185 , \33200 );
and \U$33539 ( \33882 , \33881 , \33214 );
and \U$33540 ( \33883 , \33185 , \33200 );
or \U$33541 ( \33884 , \33882 , \33883 );
xor \U$33542 ( \33885 , \33880 , \33884 );
xor \U$33543 ( \33886 , \33289 , \33300 );
xor \U$33544 ( \33887 , \33886 , \33311 );
xor \U$33545 ( \33888 , \33885 , \33887 );
xor \U$33546 ( \33889 , \33833 , \33888 );
xor \U$33547 ( \33890 , \33841 , \33848 );
xnor \U$33548 ( \33891 , \33890 , \33855 );
not \U$33549 ( \33892 , \33891 );
not \U$33550 ( \33893 , \14920 );
not \U$33551 ( \33894 , RIbb2ddb0_53);
not \U$33552 ( \33895 , \8338 );
or \U$33553 ( \33896 , \33894 , \33895 );
nand \U$33554 ( \33897 , \15796 , \16210 );
nand \U$33555 ( \33898 , \33896 , \33897 );
not \U$33556 ( \33899 , \33898 );
or \U$33557 ( \33900 , \33893 , \33899 );
nand \U$33558 ( \33901 , \33075 , \15688 );
nand \U$33559 ( \33902 , \33900 , \33901 );
not \U$33560 ( \33903 , \12692 );
not \U$33561 ( \33904 , \33064 );
or \U$33562 ( \33905 , \33903 , \33904 );
nand \U$33563 ( \33906 , \33402 , \14067 );
nand \U$33564 ( \33907 , \33905 , \33906 );
xor \U$33565 ( \33908 , \33902 , \33907 );
not \U$33566 ( \33909 , \26834 );
not \U$33567 ( \33910 , \33191 );
or \U$33568 ( \33911 , \33909 , \33910 );
nand \U$33569 ( \33912 , \33435 , \16541 );
nand \U$33570 ( \33913 , \33911 , \33912 );
xor \U$33571 ( \33914 , \33908 , \33913 );
not \U$33572 ( \33915 , \33914 );
or \U$33573 ( \33916 , \33892 , \33915 );
or \U$33574 ( \33917 , \33914 , \33891 );
not \U$33575 ( \33918 , \12285 );
not \U$33576 ( \33919 , \33101 );
or \U$33577 ( \33920 , \33918 , \33919 );
nand \U$33578 ( \33921 , \33656 , \13295 );
nand \U$33579 ( \33922 , \33920 , \33921 );
not \U$33580 ( \33923 , \12965 );
not \U$33581 ( \33924 , \33088 );
or \U$33582 ( \33925 , \33923 , \33924 );
not \U$33583 ( \33926 , RIbb2e080_47);
not \U$33584 ( \33927 , \12222 );
or \U$33585 ( \33928 , \33926 , \33927 );
nand \U$33586 ( \33929 , \14553 , \15632 );
nand \U$33587 ( \33930 , \33928 , \33929 );
nand \U$33588 ( \33931 , \33930 , \11176 );
nand \U$33589 ( \33932 , \33925 , \33931 );
xor \U$33590 ( \33933 , \33922 , \33932 );
not \U$33591 ( \33934 , \10117 );
not \U$33592 ( \33935 , RIbb2e170_45);
not \U$33593 ( \33936 , \12764 );
or \U$33594 ( \33937 , \33935 , \33936 );
nand \U$33595 ( \33938 , \32888 , \12003 );
nand \U$33596 ( \33939 , \33937 , \33938 );
not \U$33597 ( \33940 , \33939 );
or \U$33598 ( \33941 , \33934 , \33940 );
nand \U$33599 ( \33942 , \33037 , \10119 );
nand \U$33600 ( \33943 , \33941 , \33942 );
and \U$33601 ( \33944 , \33933 , \33943 );
not \U$33602 ( \33945 , \33933 );
not \U$33603 ( \33946 , \33943 );
and \U$33604 ( \33947 , \33945 , \33946 );
nor \U$33605 ( \33948 , \33944 , \33947 );
nand \U$33606 ( \33949 , \33917 , \33948 );
nand \U$33607 ( \33950 , \33916 , \33949 );
xor \U$33608 ( \33951 , \33864 , \33869 );
xor \U$33609 ( \33952 , \33951 , \33875 );
not \U$33610 ( \33953 , \33952 );
not \U$33611 ( \33954 , \9099 );
not \U$33612 ( \33955 , \33379 );
or \U$33613 ( \33956 , \33954 , \33955 );
nand \U$33614 ( \33957 , \33542 , \10449 );
nand \U$33615 ( \33958 , \33956 , \33957 );
not \U$33616 ( \33959 , \11177 );
not \U$33617 ( \33960 , \33930 );
or \U$33618 ( \33961 , \33959 , \33960 );
nand \U$33619 ( \33962 , \33734 , \11176 );
nand \U$33620 ( \33963 , \33961 , \33962 );
xor \U$33621 ( \33964 , \33958 , \33963 );
not \U$33622 ( \33965 , \10119 );
not \U$33623 ( \33966 , \33939 );
or \U$33624 ( \33967 , \33965 , \33966 );
nand \U$33625 ( \33968 , \33809 , \10117 );
nand \U$33626 ( \33969 , \33967 , \33968 );
and \U$33627 ( \33970 , \33964 , \33969 );
and \U$33628 ( \33971 , \33958 , \33963 );
or \U$33629 ( \33972 , \33970 , \33971 );
not \U$33630 ( \33973 , \33972 );
or \U$33631 ( \33974 , \33953 , \33973 );
or \U$33632 ( \33975 , \33972 , \33952 );
not \U$33633 ( \33976 , \17397 );
not \U$33634 ( \33977 , \33392 );
or \U$33635 ( \33978 , \33976 , \33977 );
nand \U$33636 ( \33979 , \33714 , \19101 );
nand \U$33637 ( \33980 , \33978 , \33979 );
not \U$33638 ( \33981 , \33980 );
not \U$33639 ( \33982 , \14930 );
not \U$33640 ( \33983 , \33898 );
or \U$33641 ( \33984 , \33982 , \33983 );
not \U$33642 ( \33985 , RIbb2ddb0_53);
not \U$33643 ( \33986 , \12790 );
or \U$33644 ( \33987 , \33985 , \33986 );
nand \U$33645 ( \33988 , \6937 , \12681 );
nand \U$33646 ( \33989 , \33987 , \33988 );
nand \U$33647 ( \33990 , \33989 , \14920 );
nand \U$33648 ( \33991 , \33984 , \33990 );
not \U$33649 ( \33992 , \33991 );
nand \U$33650 ( \33993 , \33981 , \33992 );
and \U$33651 ( \33994 , \33754 , \33763 );
not \U$33652 ( \33995 , \3886 );
not \U$33653 ( \33996 , RIbb2e710_33);
not \U$33654 ( \33997 , \23185 );
or \U$33655 ( \33998 , \33996 , \33997 );
nand \U$33656 ( \33999 , \16829 , \2935 );
nand \U$33657 ( \34000 , \33998 , \33999 );
not \U$33658 ( \34001 , \34000 );
or \U$33659 ( \34002 , \33995 , \34001 );
nand \U$33660 ( \34003 , \33368 , \4075 );
nand \U$33661 ( \34004 , \34002 , \34003 );
xor \U$33662 ( \34005 , \33994 , \34004 );
not \U$33663 ( \34006 , \4714 );
not \U$33664 ( \34007 , \33596 );
or \U$33665 ( \34008 , \34006 , \34007 );
nand \U$33666 ( \34009 , \33781 , \4712 );
nand \U$33667 ( \34010 , \34008 , \34009 );
and \U$33668 ( \34011 , \34005 , \34010 );
and \U$33669 ( \34012 , \33994 , \34004 );
or \U$33670 ( \34013 , \34011 , \34012 );
and \U$33671 ( \34014 , \33993 , \34013 );
not \U$33672 ( \34015 , \33980 );
nor \U$33673 ( \34016 , \34015 , \33992 );
nor \U$33674 ( \34017 , \34014 , \34016 );
not \U$33675 ( \34018 , \34017 );
nand \U$33676 ( \34019 , \33975 , \34018 );
nand \U$33677 ( \34020 , \33974 , \34019 );
or \U$33678 ( \34021 , \33950 , \34020 );
xor \U$33679 ( \34022 , \33583 , \33626 );
and \U$33680 ( \34023 , \34022 , \33661 );
and \U$33681 ( \34024 , \33583 , \33626 );
or \U$33682 ( \34025 , \34023 , \34024 );
nand \U$33683 ( \34026 , \34021 , \34025 );
nand \U$33684 ( \34027 , \33950 , \34020 );
nand \U$33685 ( \34028 , \34026 , \34027 );
xor \U$33686 ( \34029 , \33889 , \34028 );
not \U$33687 ( \34030 , \34029 );
or \U$33688 ( \34031 , \33831 , \34030 );
or \U$33689 ( \34032 , \34029 , \33830 );
xor \U$33690 ( \34033 , \34025 , \34020 );
xnor \U$33691 ( \34034 , \34033 , \33950 );
not \U$33692 ( \34035 , \34034 );
not \U$33693 ( \34036 , \34035 );
xor \U$33694 ( \34037 , \33598 , \33607 );
xor \U$33695 ( \34038 , \34037 , \33623 );
not \U$33696 ( \34039 , \13467 );
not \U$33697 ( \34040 , RIbb2ddb0_53);
not \U$33698 ( \34041 , \7297 );
or \U$33699 ( \34042 , \34040 , \34041 );
nand \U$33700 ( \34043 , \7296 , \13463 );
nand \U$33701 ( \34044 , \34042 , \34043 );
not \U$33702 ( \34045 , \34044 );
or \U$33703 ( \34046 , \34039 , \34045 );
nand \U$33704 ( \34047 , \33989 , \14929 );
nand \U$33705 ( \34048 , \34046 , \34047 );
not \U$33706 ( \34049 , \34048 );
not \U$33707 ( \34050 , \12692 );
not \U$33708 ( \34051 , \33408 );
or \U$33709 ( \34052 , \34050 , \34051 );
and \U$33710 ( \34053 , RIbb2dea0_51, \13863 );
not \U$33711 ( \34054 , RIbb2dea0_51);
and \U$33712 ( \34055 , \34054 , \8630 );
or \U$33713 ( \34056 , \34053 , \34055 );
nand \U$33714 ( \34057 , \34056 , \12774 );
nand \U$33715 ( \34058 , \34052 , \34057 );
not \U$33716 ( \34059 , \34058 );
nand \U$33717 ( \34060 , \34049 , \34059 );
not \U$33718 ( \34061 , \34060 );
not \U$33719 ( \34062 , \16533 );
not \U$33720 ( \34063 , \33442 );
or \U$33721 ( \34064 , \34062 , \34063 );
and \U$33722 ( \34065 , RIbb2d9f0_61, \4748 );
not \U$33723 ( \34066 , RIbb2d9f0_61);
and \U$33724 ( \34067 , \34066 , \3089 );
or \U$33725 ( \34068 , \34065 , \34067 );
nand \U$33726 ( \34069 , \34068 , \16541 );
nand \U$33727 ( \34070 , \34064 , \34069 );
not \U$33728 ( \34071 , \34070 );
or \U$33729 ( \34072 , \34061 , \34071 );
not \U$33730 ( \34073 , \34059 );
nand \U$33731 ( \34074 , \34073 , \34048 );
nand \U$33732 ( \34075 , \34072 , \34074 );
xor \U$33733 ( \34076 , \34038 , \34075 );
xor \U$33734 ( \34077 , \33629 , \33642 );
xor \U$33735 ( \34078 , \34077 , \33658 );
and \U$33736 ( \34079 , \34076 , \34078 );
and \U$33737 ( \34080 , \34038 , \34075 );
or \U$33738 ( \34081 , \34079 , \34080 );
xor \U$33739 ( \34082 , \33952 , \34017 );
not \U$33740 ( \34083 , \33972 );
xor \U$33741 ( \34084 , \34082 , \34083 );
xor \U$33742 ( \34085 , \34081 , \34084 );
not \U$33743 ( \34086 , \33891 );
and \U$33744 ( \34087 , \33948 , \34086 );
not \U$33745 ( \34088 , \33948 );
and \U$33746 ( \34089 , \34088 , \33891 );
nor \U$33747 ( \34090 , \34087 , \34089 );
not \U$33748 ( \34091 , \34090 );
xor \U$33749 ( \34092 , \33914 , \34091 );
and \U$33750 ( \34093 , \34085 , \34092 );
and \U$33751 ( \34094 , \34081 , \34084 );
or \U$33752 ( \34095 , \34093 , \34094 );
not \U$33753 ( \34096 , \34095 );
or \U$33754 ( \34097 , \34036 , \34096 );
or \U$33755 ( \34098 , \34095 , \34035 );
xor \U$33756 ( \34099 , \33859 , \33835 );
xor \U$33757 ( \34100 , \34099 , \33878 );
not \U$33758 ( \34101 , \33932 );
not \U$33759 ( \34102 , \33943 );
or \U$33760 ( \34103 , \34101 , \34102 );
or \U$33761 ( \34104 , \33943 , \33932 );
nand \U$33762 ( \34105 , \34104 , \33922 );
nand \U$33763 ( \34106 , \34103 , \34105 );
or \U$33764 ( \34107 , \33383 , \33394 );
nand \U$33765 ( \34108 , \34107 , \33373 );
nand \U$33766 ( \34109 , \33394 , \33383 );
nand \U$33767 ( \34110 , \34108 , \34109 );
xor \U$33768 ( \34111 , \34106 , \34110 );
xor \U$33769 ( \34112 , \33052 , \33066 );
xor \U$33770 ( \34113 , \34112 , \33077 );
xnor \U$33771 ( \34114 , \34111 , \34113 );
xor \U$33772 ( \34115 , \34100 , \34114 );
xor \U$33773 ( \34116 , \33902 , \33907 );
and \U$33774 ( \34117 , \34116 , \33913 );
and \U$33775 ( \34118 , \33902 , \33907 );
or \U$33776 ( \34119 , \34117 , \34118 );
xor \U$33777 ( \34120 , \33082 , \33092 );
xor \U$33778 ( \34121 , \34120 , \33103 );
xor \U$33779 ( \34122 , \34119 , \34121 );
nor \U$33780 ( \34123 , \33576 , \33570 );
not \U$33781 ( \34124 , \33565 );
or \U$33782 ( \34125 , \34123 , \34124 );
nand \U$33783 ( \34126 , \33576 , \33570 );
nand \U$33784 ( \34127 , \34125 , \34126 );
xor \U$33785 ( \34128 , \34122 , \34127 );
xnor \U$33786 ( \34129 , \34115 , \34128 );
nand \U$33787 ( \34130 , \34098 , \34129 );
nand \U$33788 ( \34131 , \34097 , \34130 );
nand \U$33789 ( \34132 , \34032 , \34131 );
nand \U$33790 ( \34133 , \34031 , \34132 );
not \U$33791 ( \34134 , \34133 );
xor \U$33792 ( \34135 , \33349 , \34134 );
xor \U$33793 ( \34136 , \33833 , \33888 );
and \U$33794 ( \34137 , \34136 , \34028 );
and \U$33795 ( \34138 , \33833 , \33888 );
or \U$33796 ( \34139 , \34137 , \34138 );
not \U$33797 ( \34140 , \34139 );
not \U$33798 ( \34141 , \34140 );
xor \U$33799 ( \34142 , \33880 , \33884 );
and \U$33800 ( \34143 , \34142 , \33887 );
and \U$33801 ( \34144 , \33880 , \33884 );
or \U$33802 ( \34145 , \34143 , \34144 );
not \U$33803 ( \34146 , \34145 );
not \U$33804 ( \34147 , RIbb2d888_64);
not \U$33805 ( \34148 , \28672 );
or \U$33806 ( \34149 , \34147 , \34148 );
nand \U$33807 ( \34150 , \33298 , \17275 );
nand \U$33808 ( \34151 , \34149 , \34150 );
not \U$33809 ( \34152 , \15182 );
not \U$33810 ( \34153 , \28587 );
or \U$33811 ( \34154 , \34152 , \34153 );
nand \U$33812 ( \34155 , \33114 , \22952 );
nand \U$33813 ( \34156 , \34154 , \34155 );
xor \U$33814 ( \34157 , \34151 , \34156 );
not \U$33815 ( \34158 , \16271 );
not \U$33816 ( \34159 , \33244 );
or \U$33817 ( \34160 , \34158 , \34159 );
nand \U$33818 ( \34161 , \17470 , \28682 );
nand \U$33819 ( \34162 , \34160 , \34161 );
xor \U$33820 ( \34163 , \34157 , \34162 );
not \U$33821 ( \34164 , \34163 );
not \U$33822 ( \34165 , \12774 );
not \U$33823 ( \34166 , \33125 );
or \U$33824 ( \34167 , \34165 , \34166 );
nand \U$33825 ( \34168 , \28549 , \12692 );
nand \U$33826 ( \34169 , \34167 , \34168 );
not \U$33827 ( \34170 , \16674 );
not \U$33828 ( \34171 , \33136 );
or \U$33829 ( \34172 , \34170 , \34171 );
nand \U$33830 ( \34173 , \28558 , \15738 );
nand \U$33831 ( \34174 , \34172 , \34173 );
xor \U$33832 ( \34175 , \34169 , \34174 );
not \U$33833 ( \34176 , \16541 );
not \U$33834 ( \34177 , \33309 );
or \U$33835 ( \34178 , \34176 , \34177 );
nand \U$33836 ( \34179 , \28598 , \26834 );
nand \U$33837 ( \34180 , \34178 , \34179 );
xnor \U$33838 ( \34181 , \34175 , \34180 );
not \U$33839 ( \34182 , \34181 );
or \U$33840 ( \34183 , \34164 , \34182 );
or \U$33841 ( \34184 , \34163 , \34181 );
nand \U$33842 ( \34185 , \34183 , \34184 );
xor \U$33843 ( \34186 , \32959 , \32961 );
and \U$33844 ( \34187 , \34186 , \33044 );
and \U$33845 ( \34188 , \32959 , \32961 );
or \U$33846 ( \34189 , \34187 , \34188 );
not \U$33847 ( \34190 , \34189 );
and \U$33848 ( \34191 , \34185 , \34190 );
not \U$33849 ( \34192 , \34185 );
and \U$33850 ( \34193 , \34192 , \34189 );
nor \U$33851 ( \34194 , \34191 , \34193 );
not \U$33852 ( \34195 , \34194 );
or \U$33853 ( \34196 , \34146 , \34195 );
or \U$33854 ( \34197 , \34145 , \34194 );
nand \U$33855 ( \34198 , \34196 , \34197 );
xor \U$33856 ( \34199 , \33281 , \33275 );
xor \U$33857 ( \34200 , \34199 , \33246 );
buf \U$33858 ( \34201 , \34200 );
xor \U$33859 ( \34202 , \34119 , \34121 );
and \U$33860 ( \34203 , \34202 , \34127 );
and \U$33861 ( \34204 , \34119 , \34121 );
or \U$33862 ( \34205 , \34203 , \34204 );
or \U$33863 ( \34206 , \34201 , \34205 );
not \U$33864 ( \34207 , \34106 );
not \U$33865 ( \34208 , \34113 );
or \U$33866 ( \34209 , \34207 , \34208 );
or \U$33867 ( \34210 , \34106 , \34113 );
nand \U$33868 ( \34211 , \34210 , \34110 );
nand \U$33869 ( \34212 , \34209 , \34211 );
nand \U$33870 ( \34213 , \34206 , \34212 );
nand \U$33871 ( \34214 , \34205 , \34201 );
nand \U$33872 ( \34215 , \34213 , \34214 );
not \U$33873 ( \34216 , \34215 );
and \U$33874 ( \34217 , \34198 , \34216 );
not \U$33875 ( \34218 , \34198 );
and \U$33876 ( \34219 , \34218 , \34215 );
nor \U$33877 ( \34220 , \34217 , \34219 );
not \U$33878 ( \34221 , \34220 );
not \U$33879 ( \34222 , \34221 );
or \U$33880 ( \34223 , \34141 , \34222 );
nand \U$33881 ( \34224 , \34220 , \34139 );
nand \U$33882 ( \34225 , \34223 , \34224 );
xor \U$33883 ( \34226 , \34200 , \34212 );
xnor \U$33884 ( \34227 , \34226 , \34205 );
not \U$33885 ( \34228 , \34227 );
not \U$33886 ( \34229 , \34228 );
not \U$33887 ( \34230 , \34100 );
nand \U$33888 ( \34231 , \34230 , \34114 );
not \U$33889 ( \34232 , \34231 );
not \U$33890 ( \34233 , \34128 );
or \U$33891 ( \34234 , \34232 , \34233 );
not \U$33892 ( \34235 , \34114 );
nand \U$33893 ( \34236 , \34235 , \34100 );
nand \U$33894 ( \34237 , \34234 , \34236 );
not \U$33895 ( \34238 , \34237 );
or \U$33896 ( \34239 , \34229 , \34238 );
not \U$33897 ( \34240 , \34227 );
not \U$33898 ( \34241 , \34237 );
not \U$33899 ( \34242 , \34241 );
or \U$33900 ( \34243 , \34240 , \34242 );
xor \U$33901 ( \34244 , \33045 , \33140 );
xor \U$33902 ( \34245 , \34244 , \33219 );
nand \U$33903 ( \34246 , \34243 , \34245 );
nand \U$33904 ( \34247 , \34239 , \34246 );
not \U$33905 ( \34248 , \34247 );
and \U$33906 ( \34249 , \34225 , \34248 );
not \U$33907 ( \34250 , \34225 );
and \U$33908 ( \34251 , \34250 , \34247 );
nor \U$33909 ( \34252 , \34249 , \34251 );
xor \U$33910 ( \34253 , \34135 , \34252 );
not \U$33911 ( \34254 , \34228 );
not \U$33912 ( \34255 , \34241 );
or \U$33913 ( \34256 , \34254 , \34255 );
nand \U$33914 ( \34257 , \34227 , \34237 );
nand \U$33915 ( \34258 , \34256 , \34257 );
not \U$33916 ( \34259 , \34245 );
and \U$33917 ( \34260 , \34258 , \34259 );
not \U$33918 ( \34261 , \34258 );
and \U$33919 ( \34262 , \34261 , \34245 );
nor \U$33920 ( \34263 , \34260 , \34262 );
xor \U$33921 ( \34264 , \33558 , \33825 );
xnor \U$33922 ( \34265 , \34264 , \33828 );
not \U$33923 ( \34266 , \34265 );
not \U$33924 ( \34267 , \34266 );
xor \U$33925 ( \34268 , \34013 , \33991 );
xor \U$33926 ( \34269 , \34268 , \33980 );
xor \U$33927 ( \34270 , \33958 , \33963 );
xor \U$33928 ( \34271 , \34270 , \33969 );
xor \U$33929 ( \34272 , \34269 , \34271 );
xor \U$33930 ( \34273 , \33410 , \33444 );
xor \U$33931 ( \34274 , \34273 , \33426 );
and \U$33932 ( \34275 , \34272 , \34274 );
and \U$33933 ( \34276 , \34269 , \34271 );
or \U$33934 ( \34277 , \34275 , \34276 );
not \U$33935 ( \34278 , \34277 );
and \U$33936 ( \34279 , \33446 , \33395 );
not \U$33937 ( \34280 , \33446 );
and \U$33938 ( \34281 , \34280 , \33396 );
nor \U$33939 ( \34282 , \34279 , \34281 );
xor \U$33940 ( \34283 , \34282 , \33556 );
not \U$33941 ( \34284 , \34283 );
not \U$33942 ( \34285 , \34284 );
or \U$33943 ( \34286 , \34278 , \34285 );
xor \U$33944 ( \34287 , \33994 , \34004 );
xor \U$33945 ( \34288 , \34287 , \34010 );
not \U$33946 ( \34289 , \4075 );
not \U$33947 ( \34290 , \34000 );
or \U$33948 ( \34291 , \34289 , \34290 );
not \U$33949 ( \34292 , RIbb2e710_33);
not \U$33950 ( \34293 , \16706 );
not \U$33951 ( \34294 , \34293 );
or \U$33952 ( \34295 , \34292 , \34294 );
nand \U$33953 ( \34296 , \16706 , \3877 );
nand \U$33954 ( \34297 , \34295 , \34296 );
nand \U$33955 ( \34298 , \34297 , \3886 );
nand \U$33956 ( \34299 , \34291 , \34298 );
not \U$33957 ( \34300 , \34299 );
not \U$33958 ( \34301 , \9099 );
not \U$33959 ( \34302 , \33549 );
or \U$33960 ( \34303 , \34301 , \34302 );
not \U$33961 ( \34304 , RIbb2e260_43);
not \U$33962 ( \34305 , \21756 );
or \U$33963 ( \34306 , \34304 , \34305 );
nand \U$33964 ( \34307 , \14844 , \8347 );
nand \U$33965 ( \34308 , \34306 , \34307 );
nand \U$33966 ( \34309 , \34308 , \10449 );
nand \U$33967 ( \34310 , \34303 , \34309 );
not \U$33968 ( \34311 , \34310 );
or \U$33969 ( \34312 , \34300 , \34311 );
or \U$33970 ( \34313 , \34310 , \34299 );
and \U$33971 ( \34314 , \17506 , \2924 );
not \U$33972 ( \34315 , \2941 );
not \U$33973 ( \34316 , \33772 );
or \U$33974 ( \34317 , \34315 , \34316 );
and \U$33975 ( \34318 , RIbb2e800_31, \28621 );
not \U$33976 ( \34319 , RIbb2e800_31);
and \U$33977 ( \34320 , \34319 , \17519 );
nor \U$33978 ( \34321 , \34318 , \34320 );
nand \U$33979 ( \34322 , \34321 , \2938 );
nand \U$33980 ( \34323 , \34317 , \34322 );
xor \U$33981 ( \34324 , \34314 , \34323 );
not \U$33982 ( \34325 , \4075 );
not \U$33983 ( \34326 , \34297 );
or \U$33984 ( \34327 , \34325 , \34326 );
not \U$33985 ( \34328 , RIbb2e710_33);
not \U$33986 ( \34329 , \27234 );
or \U$33987 ( \34330 , \34328 , \34329 );
nand \U$33988 ( \34331 , \27237 , \3877 );
nand \U$33989 ( \34332 , \34330 , \34331 );
nand \U$33990 ( \34333 , \34332 , \3886 );
nand \U$33991 ( \34334 , \34327 , \34333 );
and \U$33992 ( \34335 , \34324 , \34334 );
and \U$33993 ( \34336 , \34314 , \34323 );
or \U$33994 ( \34337 , \34335 , \34336 );
nand \U$33995 ( \34338 , \34313 , \34337 );
nand \U$33996 ( \34339 , \34312 , \34338 );
xor \U$33997 ( \34340 , \34288 , \34339 );
not \U$33998 ( \34341 , \17275 );
not \U$33999 ( \34342 , RIbb2d900_63);
not \U$34000 ( \34343 , \4029 );
or \U$34001 ( \34344 , \34342 , \34343 );
nand \U$34002 ( \34345 , \16180 , \17262 );
nand \U$34003 ( \34346 , \34344 , \34345 );
not \U$34004 ( \34347 , \34346 );
or \U$34005 ( \34348 , \34341 , \34347 );
nand \U$34006 ( \34349 , \33424 , RIbb2d888_64);
nand \U$34007 ( \34350 , \34348 , \34349 );
and \U$34008 ( \34351 , \34340 , \34350 );
and \U$34009 ( \34352 , \34288 , \34339 );
or \U$34010 ( \34353 , \34351 , \34352 );
and \U$34011 ( \34354 , RIbb2e350_41, \13546 );
not \U$34012 ( \34355 , RIbb2e350_41);
and \U$34013 ( \34356 , \34355 , \13545 );
or \U$34014 ( \34357 , \34354 , \34356 );
not \U$34015 ( \34358 , \34357 );
not \U$34016 ( \34359 , \8361 );
or \U$34017 ( \34360 , \34358 , \34359 );
nand \U$34018 ( \34361 , \33673 , \8353 );
nand \U$34019 ( \34362 , \34360 , \34361 );
not \U$34020 ( \34363 , \7104 );
not \U$34021 ( \34364 , \33533 );
or \U$34022 ( \34365 , \34363 , \34364 );
and \U$34023 ( \34366 , RIbb2e440_39, \16309 );
not \U$34024 ( \34367 , RIbb2e440_39);
not \U$34025 ( \34368 , \20577 );
and \U$34026 ( \34369 , \34367 , \34368 );
or \U$34027 ( \34370 , \34366 , \34369 );
nand \U$34028 ( \34371 , \34370 , \8445 );
nand \U$34029 ( \34372 , \34365 , \34371 );
xor \U$34030 ( \34373 , \34362 , \34372 );
not \U$34031 ( \34374 , \6241 );
not \U$34032 ( \34375 , \33683 );
or \U$34033 ( \34376 , \34374 , \34375 );
not \U$34034 ( \34377 , RIbb2e530_37);
not \U$34035 ( \34378 , \15754 );
or \U$34036 ( \34379 , \34377 , \34378 );
nand \U$34037 ( \34380 , \16568 , \6246 );
nand \U$34038 ( \34381 , \34379 , \34380 );
nand \U$34039 ( \34382 , \34381 , \6251 );
nand \U$34040 ( \34383 , \34376 , \34382 );
and \U$34041 ( \34384 , \34373 , \34383 );
and \U$34042 ( \34385 , \34362 , \34372 );
or \U$34043 ( \34386 , \34384 , \34385 );
not \U$34044 ( \34387 , \11176 );
not \U$34045 ( \34388 , RIbb2e080_47);
not \U$34046 ( \34389 , \12260 );
or \U$34047 ( \34390 , \34388 , \34389 );
nand \U$34048 ( \34391 , \12261 , \10113 );
nand \U$34049 ( \34392 , \34390 , \34391 );
not \U$34050 ( \34393 , \34392 );
or \U$34051 ( \34394 , \34387 , \34393 );
nand \U$34052 ( \34395 , \33741 , \11177 );
nand \U$34053 ( \34396 , \34394 , \34395 );
not \U$34054 ( \34397 , \34396 );
not \U$34055 ( \34398 , \19101 );
and \U$34056 ( \34399 , RIbb2dbd0_57, \21570 );
not \U$34057 ( \34400 , RIbb2dbd0_57);
and \U$34058 ( \34401 , \34400 , \7308 );
or \U$34059 ( \34402 , \34399 , \34401 );
not \U$34060 ( \34403 , \34402 );
or \U$34061 ( \34404 , \34398 , \34403 );
nand \U$34062 ( \34405 , \33707 , \15738 );
nand \U$34063 ( \34406 , \34404 , \34405 );
not \U$34064 ( \34407 , \34406 );
or \U$34065 ( \34408 , \34397 , \34407 );
or \U$34066 ( \34409 , \34406 , \34396 );
not \U$34067 ( \34410 , \10119 );
not \U$34068 ( \34411 , \33816 );
or \U$34069 ( \34412 , \34410 , \34411 );
not \U$34070 ( \34413 , RIbb2e170_45);
not \U$34071 ( \34414 , \22070 );
or \U$34072 ( \34415 , \34413 , \34414 );
nand \U$34073 ( \34416 , \12838 , \13372 );
nand \U$34074 ( \34417 , \34415 , \34416 );
nand \U$34075 ( \34418 , \34417 , \10117 );
nand \U$34076 ( \34419 , \34412 , \34418 );
nand \U$34077 ( \34420 , \34409 , \34419 );
nand \U$34078 ( \34421 , \34408 , \34420 );
xor \U$34079 ( \34422 , \34386 , \34421 );
not \U$34080 ( \34423 , \16271 );
and \U$34081 ( \34424 , RIbb2dae0_59, \4698 );
not \U$34082 ( \34425 , RIbb2dae0_59);
and \U$34083 ( \34426 , \34425 , \4699 );
or \U$34084 ( \34427 , \34424 , \34426 );
not \U$34085 ( \34428 , \34427 );
or \U$34086 ( \34429 , \34423 , \34428 );
nand \U$34087 ( \34430 , \33725 , \17470 );
nand \U$34088 ( \34431 , \34429 , \34430 );
not \U$34089 ( \34432 , \12284 );
not \U$34090 ( \34433 , \33692 );
or \U$34091 ( \34434 , \34432 , \34433 );
not \U$34092 ( \34435 , RIbb2df90_49);
not \U$34093 ( \34436 , \13929 );
or \U$34094 ( \34437 , \34435 , \34436 );
nand \U$34095 ( \34438 , \10300 , \12278 );
nand \U$34096 ( \34439 , \34437 , \34438 );
nand \U$34097 ( \34440 , \34439 , \13295 );
nand \U$34098 ( \34441 , \34434 , \34440 );
or \U$34099 ( \34442 , \34431 , \34441 );
not \U$34100 ( \34443 , \34442 );
xor \U$34101 ( \34444 , \33764 , \33774 );
xor \U$34102 ( \34445 , \34444 , \33790 );
not \U$34103 ( \34446 , \34445 );
or \U$34104 ( \34447 , \34443 , \34446 );
nand \U$34105 ( \34448 , \34431 , \34441 );
nand \U$34106 ( \34449 , \34447 , \34448 );
and \U$34107 ( \34450 , \34422 , \34449 );
and \U$34108 ( \34451 , \34386 , \34421 );
or \U$34109 ( \34452 , \34450 , \34451 );
xor \U$34110 ( \34453 , \34353 , \34452 );
xor \U$34111 ( \34454 , \33522 , \33535 );
xor \U$34112 ( \34455 , \34454 , \33551 );
xor \U$34113 ( \34456 , \33675 , \33685 );
xor \U$34114 ( \34457 , \34456 , \33696 );
xor \U$34115 ( \34458 , \34455 , \34457 );
or \U$34116 ( \34459 , RIbb2e788_32, RIbb2e710_33);
nand \U$34117 ( \34460 , \34459 , \17506 );
and \U$34118 ( \34461 , RIbb2e788_32, RIbb2e710_33);
nor \U$34119 ( \34462 , \34461 , \8810 );
and \U$34120 ( \34463 , \34460 , \34462 );
not \U$34121 ( \34464 , \2941 );
not \U$34122 ( \34465 , \34321 );
or \U$34123 ( \34466 , \34464 , \34465 );
or \U$34124 ( \34467 , \17506 , \8810 );
or \U$34125 ( \34468 , \20747 , RIbb2e800_31);
nand \U$34126 ( \34469 , \34467 , \34468 );
nand \U$34127 ( \34470 , \34469 , \2938 );
nand \U$34128 ( \34471 , \34466 , \34470 );
and \U$34129 ( \34472 , \34463 , \34471 );
not \U$34130 ( \34473 , \4714 );
not \U$34131 ( \34474 , \33788 );
or \U$34132 ( \34475 , \34473 , \34474 );
not \U$34133 ( \34476 , RIbb2e620_35);
not \U$34134 ( \34477 , \16727 );
or \U$34135 ( \34478 , \34476 , \34477 );
nand \U$34136 ( \34479 , \19831 , \6002 );
nand \U$34137 ( \34480 , \34478 , \34479 );
nand \U$34138 ( \34481 , \34480 , \4712 );
nand \U$34139 ( \34482 , \34475 , \34481 );
xor \U$34140 ( \34483 , \34472 , \34482 );
not \U$34141 ( \34484 , \6241 );
not \U$34142 ( \34485 , \34381 );
or \U$34143 ( \34486 , \34484 , \34485 );
not \U$34144 ( \34487 , RIbb2e530_37);
not \U$34145 ( \34488 , \16844 );
or \U$34146 ( \34489 , \34487 , \34488 );
nand \U$34147 ( \34490 , \16576 , \8701 );
nand \U$34148 ( \34491 , \34489 , \34490 );
nand \U$34149 ( \34492 , \34491 , \6251 );
nand \U$34150 ( \34493 , \34486 , \34492 );
and \U$34151 ( \34494 , \34483 , \34493 );
and \U$34152 ( \34495 , \34472 , \34482 );
or \U$34153 ( \34496 , \34494 , \34495 );
not \U$34154 ( \34497 , \14920 );
not \U$34155 ( \34498 , RIbb2ddb0_53);
not \U$34156 ( \34499 , \12211 );
or \U$34157 ( \34500 , \34498 , \34499 );
not \U$34158 ( \34501 , \12210 );
nand \U$34159 ( \34502 , \34501 , \16210 );
nand \U$34160 ( \34503 , \34500 , \34502 );
not \U$34161 ( \34504 , \34503 );
or \U$34162 ( \34505 , \34497 , \34504 );
nand \U$34163 ( \34506 , \34044 , \15688 );
nand \U$34164 ( \34507 , \34505 , \34506 );
xor \U$34165 ( \34508 , \34496 , \34507 );
not \U$34166 ( \34509 , \22952 );
not \U$34167 ( \34510 , \8638 );
not \U$34168 ( \34511 , RIbb2dcc0_55);
not \U$34169 ( \34512 , \34511 );
and \U$34170 ( \34513 , \34510 , \34512 );
and \U$34171 ( \34514 , \19870 , \18174 );
nor \U$34172 ( \34515 , \34513 , \34514 );
not \U$34173 ( \34516 , \34515 );
not \U$34174 ( \34517 , \34516 );
or \U$34175 ( \34518 , \34509 , \34517 );
nand \U$34176 ( \34519 , \33800 , \15182 );
nand \U$34177 ( \34520 , \34518 , \34519 );
and \U$34178 ( \34521 , \34508 , \34520 );
and \U$34179 ( \34522 , \34496 , \34507 );
or \U$34180 ( \34523 , \34521 , \34522 );
and \U$34181 ( \34524 , \34458 , \34523 );
and \U$34182 ( \34525 , \34455 , \34457 );
or \U$34183 ( \34526 , \34524 , \34525 );
and \U$34184 ( \34527 , \34453 , \34526 );
and \U$34185 ( \34528 , \34353 , \34452 );
or \U$34186 ( \34529 , \34527 , \34528 );
not \U$34187 ( \34530 , \34277 );
nand \U$34188 ( \34531 , \34530 , \34283 );
nand \U$34189 ( \34532 , \34529 , \34531 );
nand \U$34190 ( \34533 , \34286 , \34532 );
not \U$34191 ( \34534 , \34533 );
or \U$34192 ( \34535 , \34267 , \34534 );
not \U$34193 ( \34536 , \34533 );
not \U$34194 ( \34537 , \34536 );
not \U$34195 ( \34538 , \34265 );
or \U$34196 ( \34539 , \34537 , \34538 );
xor \U$34197 ( \34540 , \33823 , \33577 );
xor \U$34198 ( \34541 , \34540 , \33662 );
not \U$34199 ( \34542 , \34541 );
xor \U$34200 ( \34543 , \33517 , \33554 );
xor \U$34201 ( \34544 , \34543 , \33504 );
xor \U$34202 ( \34545 , \33716 , \33727 );
xor \U$34203 ( \34546 , \34545 , \33743 );
not \U$34204 ( \34547 , \34546 );
and \U$34205 ( \34548 , \34048 , \34059 );
not \U$34206 ( \34549 , \34048 );
and \U$34207 ( \34550 , \34549 , \34058 );
nor \U$34208 ( \34551 , \34548 , \34550 );
and \U$34209 ( \34552 , \34551 , \34070 );
not \U$34210 ( \34553 , \34551 );
not \U$34211 ( \34554 , \34070 );
and \U$34212 ( \34555 , \34553 , \34554 );
nor \U$34213 ( \34556 , \34552 , \34555 );
not \U$34214 ( \34557 , \34556 );
not \U$34215 ( \34558 , \34557 );
or \U$34216 ( \34559 , \34547 , \34558 );
or \U$34217 ( \34560 , \34557 , \34546 );
not \U$34218 ( \34561 , \12774 );
and \U$34219 ( \34562 , RIbb2dea0_51, \12820 );
not \U$34220 ( \34563 , RIbb2dea0_51);
and \U$34221 ( \34564 , \34563 , \12821 );
or \U$34222 ( \34565 , \34562 , \34564 );
not \U$34223 ( \34566 , \34565 );
or \U$34224 ( \34567 , \34561 , \34566 );
nand \U$34225 ( \34568 , \34056 , \12692 );
nand \U$34226 ( \34569 , \34567 , \34568 );
not \U$34227 ( \34570 , \34569 );
not \U$34228 ( \34571 , \17275 );
not \U$34229 ( \34572 , RIbb2d900_63);
not \U$34230 ( \34573 , \3276 );
or \U$34231 ( \34574 , \34572 , \34573 );
nand \U$34232 ( \34575 , \3003 , \17262 );
nand \U$34233 ( \34576 , \34574 , \34575 );
not \U$34234 ( \34577 , \34576 );
or \U$34235 ( \34578 , \34571 , \34577 );
nand \U$34236 ( \34579 , \34346 , RIbb2d888_64);
nand \U$34237 ( \34580 , \34578 , \34579 );
not \U$34238 ( \34581 , \34580 );
or \U$34239 ( \34582 , \34570 , \34581 );
or \U$34240 ( \34583 , \34580 , \34569 );
not \U$34241 ( \34584 , \18717 );
not \U$34242 ( \34585 , RIbb2d9f0_61);
not \U$34243 ( \34586 , \4087 );
or \U$34244 ( \34587 , \34585 , \34586 );
nand \U$34245 ( \34588 , \16153 , \16254 );
nand \U$34246 ( \34589 , \34587 , \34588 );
not \U$34247 ( \34590 , \34589 );
or \U$34248 ( \34591 , \34584 , \34590 );
nand \U$34249 ( \34592 , \34068 , \26834 );
nand \U$34250 ( \34593 , \34591 , \34592 );
nand \U$34251 ( \34594 , \34583 , \34593 );
nand \U$34252 ( \34595 , \34582 , \34594 );
nand \U$34253 ( \34596 , \34560 , \34595 );
nand \U$34254 ( \34597 , \34559 , \34596 );
xor \U$34255 ( \34598 , \34544 , \34597 );
xor \U$34256 ( \34599 , \33699 , \33746 );
xor \U$34257 ( \34600 , \34599 , \33821 );
and \U$34258 ( \34601 , \34598 , \34600 );
and \U$34259 ( \34602 , \34544 , \34597 );
or \U$34260 ( \34603 , \34601 , \34602 );
not \U$34261 ( \34604 , \34603 );
not \U$34262 ( \34605 , \34604 );
or \U$34263 ( \34606 , \34542 , \34605 );
xor \U$34264 ( \34607 , \34081 , \34084 );
xor \U$34265 ( \34608 , \34607 , \34092 );
nand \U$34266 ( \34609 , \34606 , \34608 );
not \U$34267 ( \34610 , \34541 );
nand \U$34268 ( \34611 , \34603 , \34610 );
nand \U$34269 ( \34612 , \34609 , \34611 );
nand \U$34270 ( \34613 , \34539 , \34612 );
nand \U$34271 ( \34614 , \34535 , \34613 );
not \U$34272 ( \34615 , \34614 );
xor \U$34273 ( \34616 , \34263 , \34615 );
xor \U$34274 ( \34617 , \33830 , \34029 );
xnor \U$34275 ( \34618 , \34617 , \34131 );
and \U$34276 ( \34619 , \34616 , \34618 );
and \U$34277 ( \34620 , \34263 , \34615 );
or \U$34278 ( \34621 , \34619 , \34620 );
nand \U$34279 ( \34622 , \34253 , \34621 );
not \U$34280 ( \34623 , \33335 );
not \U$34281 ( \34624 , \33315 );
or \U$34282 ( \34625 , \34623 , \34624 );
or \U$34283 ( \34626 , \33335 , \33315 );
nand \U$34284 ( \34627 , \34626 , \33330 );
nand \U$34285 ( \34628 , \34625 , \34627 );
xor \U$34286 ( \34629 , \28830 , \28827 );
xnor \U$34287 ( \34630 , \34629 , \28894 );
not \U$34288 ( \34631 , \28782 );
xor \U$34289 ( \34632 , \28772 , \34631 );
xnor \U$34290 ( \34633 , \34632 , \28737 );
not \U$34291 ( \34634 , \34633 );
xor \U$34292 ( \34635 , \34630 , \34634 );
not \U$34293 ( \34636 , \33322 );
not \U$34294 ( \34637 , \33327 );
or \U$34295 ( \34638 , \34636 , \34637 );
not \U$34296 ( \34639 , \33322 );
nand \U$34297 ( \34640 , \34639 , \33328 );
nand \U$34298 ( \34641 , \34640 , \33320 );
nand \U$34299 ( \34642 , \34638 , \34641 );
xor \U$34300 ( \34643 , \34635 , \34642 );
xor \U$34301 ( \34644 , \34628 , \34643 );
not \U$34302 ( \34645 , \33285 );
not \U$34303 ( \34646 , \33237 );
or \U$34304 ( \34647 , \34645 , \34646 );
nand \U$34305 ( \34648 , \34647 , \33314 );
not \U$34306 ( \34649 , \33237 );
nand \U$34307 ( \34650 , \34649 , \33286 );
nand \U$34308 ( \34651 , \34648 , \34650 );
not \U$34309 ( \34652 , \34651 );
not \U$34310 ( \34653 , \34169 );
not \U$34311 ( \34654 , \34174 );
or \U$34312 ( \34655 , \34653 , \34654 );
or \U$34313 ( \34656 , \34174 , \34169 );
nand \U$34314 ( \34657 , \34656 , \34180 );
nand \U$34315 ( \34658 , \34655 , \34657 );
xor \U$34316 ( \34659 , \28504 , \28517 );
xor \U$34317 ( \34660 , \34659 , \28528 );
not \U$34318 ( \34661 , \34660 );
and \U$34319 ( \34662 , \34658 , \34661 );
not \U$34320 ( \34663 , \34658 );
and \U$34321 ( \34664 , \34663 , \34660 );
or \U$34322 ( \34665 , \34662 , \34664 );
and \U$34323 ( \34666 , \28575 , \28551 );
not \U$34324 ( \34667 , \28575 );
and \U$34325 ( \34668 , \34667 , \28552 );
nor \U$34326 ( \34669 , \34666 , \34668 );
and \U$34327 ( \34670 , \34669 , \28563 );
not \U$34328 ( \34671 , \34669 );
and \U$34329 ( \34672 , \34671 , \28562 );
nor \U$34330 ( \34673 , \34670 , \34672 );
not \U$34331 ( \34674 , \34673 );
buf \U$34332 ( \34675 , \34674 );
and \U$34333 ( \34676 , \34665 , \34675 );
not \U$34334 ( \34677 , \34665 );
not \U$34335 ( \34678 , \34675 );
and \U$34336 ( \34679 , \34677 , \34678 );
nor \U$34337 ( \34680 , \34676 , \34679 );
and \U$34338 ( \34681 , \34652 , \34680 );
not \U$34339 ( \34682 , \34652 );
not \U$34340 ( \34683 , \34680 );
and \U$34341 ( \34684 , \34682 , \34683 );
nor \U$34342 ( \34685 , \34681 , \34684 );
xor \U$34343 ( \34686 , \28440 , \28449 );
xor \U$34344 ( \34687 , \34686 , \28458 );
xor \U$34345 ( \34688 , \34151 , \34156 );
and \U$34346 ( \34689 , \34688 , \34162 );
and \U$34347 ( \34690 , \34151 , \34156 );
or \U$34348 ( \34691 , \34689 , \34690 );
xor \U$34349 ( \34692 , \34687 , \34691 );
xor \U$34350 ( \34693 , \28665 , \28676 );
xor \U$34351 ( \34694 , \34693 , \28686 );
xor \U$34352 ( \34695 , \34692 , \34694 );
and \U$34353 ( \34696 , \34685 , \34695 );
not \U$34354 ( \34697 , \34685 );
not \U$34355 ( \34698 , \34695 );
and \U$34356 ( \34699 , \34697 , \34698 );
nor \U$34357 ( \34700 , \34696 , \34699 );
xor \U$34358 ( \34701 , \34644 , \34700 );
not \U$34359 ( \34702 , \34139 );
not \U$34360 ( \34703 , \34221 );
or \U$34361 ( \34704 , \34702 , \34703 );
not \U$34362 ( \34705 , \34220 );
not \U$34363 ( \34706 , \34140 );
or \U$34364 ( \34707 , \34705 , \34706 );
nand \U$34365 ( \34708 , \34707 , \34247 );
nand \U$34366 ( \34709 , \34704 , \34708 );
xor \U$34367 ( \34710 , \34701 , \34709 );
not \U$34368 ( \34711 , \34145 );
not \U$34369 ( \34712 , \34711 );
not \U$34370 ( \34713 , \34194 );
or \U$34371 ( \34714 , \34712 , \34713 );
nand \U$34372 ( \34715 , \34714 , \34215 );
or \U$34373 ( \34716 , \34194 , \34711 );
nand \U$34374 ( \34717 , \34715 , \34716 );
not \U$34375 ( \34718 , \34181 );
not \U$34376 ( \34719 , \34718 );
not \U$34377 ( \34720 , \34163 );
or \U$34378 ( \34721 , \34719 , \34720 );
or \U$34379 ( \34722 , \34163 , \34718 );
nand \U$34380 ( \34723 , \34722 , \34189 );
nand \U$34381 ( \34724 , \34721 , \34723 );
xor \U$34382 ( \34725 , \32746 , \32748 );
and \U$34383 ( \34726 , \34725 , \32774 );
and \U$34384 ( \34727 , \32746 , \32748 );
or \U$34385 ( \34728 , \34726 , \34727 );
xor \U$34386 ( \34729 , \28582 , \28591 );
xor \U$34387 ( \34730 , \34729 , \28602 );
xnor \U$34388 ( \34731 , \34728 , \34730 );
xor \U$34389 ( \34732 , \32809 , \32861 );
and \U$34390 ( \34733 , \34732 , \32897 );
and \U$34391 ( \34734 , \32809 , \32861 );
or \U$34392 ( \34735 , \34733 , \34734 );
xor \U$34393 ( \34736 , \34731 , \34735 );
not \U$34394 ( \34737 , \34736 );
xor \U$34395 ( \34738 , \34724 , \34737 );
not \U$34396 ( \34739 , \32775 );
not \U$34397 ( \34740 , \32898 );
or \U$34398 ( \34741 , \34739 , \34740 );
or \U$34399 ( \34742 , \32775 , \32898 );
nand \U$34400 ( \34743 , \34742 , \32954 );
nand \U$34401 ( \34744 , \34741 , \34743 );
xnor \U$34402 ( \34745 , \34738 , \34744 );
not \U$34403 ( \34746 , \34745 );
xor \U$34404 ( \34747 , \34717 , \34746 );
not \U$34405 ( \34748 , \32955 );
not \U$34406 ( \34749 , \33223 );
or \U$34407 ( \34750 , \34748 , \34749 );
nand \U$34408 ( \34751 , \34750 , \33344 );
nand \U$34409 ( \34752 , \32956 , \33222 );
nand \U$34410 ( \34753 , \34751 , \34752 );
xnor \U$34411 ( \34754 , \34747 , \34753 );
xnor \U$34412 ( \34755 , \34710 , \34754 );
xor \U$34413 ( \34756 , \33349 , \34134 );
and \U$34414 ( \34757 , \34756 , \34252 );
and \U$34415 ( \34758 , \33349 , \34134 );
or \U$34416 ( \34759 , \34757 , \34758 );
nand \U$34417 ( \34760 , \34755 , \34759 );
xor \U$34418 ( \34761 , \34263 , \34615 );
xor \U$34419 ( \34762 , \34761 , \34618 );
xor \U$34420 ( \34763 , \34034 , \34095 );
xor \U$34421 ( \34764 , \34763 , \34129 );
xor \U$34422 ( \34765 , \34038 , \34075 );
xor \U$34423 ( \34766 , \34765 , \34078 );
not \U$34424 ( \34767 , \34766 );
xor \U$34425 ( \34768 , \34269 , \34271 );
xor \U$34426 ( \34769 , \34768 , \34274 );
not \U$34427 ( \34770 , \34769 );
or \U$34428 ( \34771 , \34767 , \34770 );
or \U$34429 ( \34772 , \34766 , \34769 );
xor \U$34430 ( \34773 , \34288 , \34339 );
xor \U$34431 ( \34774 , \34773 , \34350 );
not \U$34432 ( \34775 , \34774 );
xor \U$34433 ( \34776 , \33793 , \33802 );
xor \U$34434 ( \34777 , \34776 , \33818 );
not \U$34435 ( \34778 , \34777 );
nand \U$34436 ( \34779 , \34775 , \34778 );
not \U$34437 ( \34780 , \34779 );
xor \U$34438 ( \34781 , \34314 , \34323 );
xor \U$34439 ( \34782 , \34781 , \34334 );
not \U$34440 ( \34783 , \7103 );
and \U$34441 ( \34784 , RIbb2e440_39, \15469 );
not \U$34442 ( \34785 , RIbb2e440_39);
and \U$34443 ( \34786 , \34785 , \17682 );
or \U$34444 ( \34787 , \34784 , \34786 );
not \U$34445 ( \34788 , \34787 );
or \U$34446 ( \34789 , \34783 , \34788 );
nand \U$34447 ( \34790 , \34370 , \7104 );
nand \U$34448 ( \34791 , \34789 , \34790 );
xor \U$34449 ( \34792 , \34782 , \34791 );
not \U$34450 ( \34793 , RIbb2e260_43);
not \U$34451 ( \34794 , \13211 );
or \U$34452 ( \34795 , \34793 , \34794 );
nand \U$34453 ( \34796 , \13474 , \8347 );
nand \U$34454 ( \34797 , \34795 , \34796 );
not \U$34455 ( \34798 , \34797 );
not \U$34456 ( \34799 , \9098 );
or \U$34457 ( \34800 , \34798 , \34799 );
not \U$34458 ( \34801 , \34308 );
not \U$34459 ( \34802 , \10451 );
or \U$34460 ( \34803 , \34801 , \34802 );
nand \U$34461 ( \34804 , \34800 , \34803 );
and \U$34462 ( \34805 , \34792 , \34804 );
and \U$34463 ( \34806 , \34782 , \34791 );
or \U$34464 ( \34807 , \34805 , \34806 );
not \U$34465 ( \34808 , \34807 );
xor \U$34466 ( \34809 , \34299 , \34337 );
xnor \U$34467 ( \34810 , \34809 , \34310 );
nand \U$34468 ( \34811 , \34808 , \34810 );
not \U$34469 ( \34812 , \34811 );
not \U$34470 ( \34813 , \4075 );
not \U$34471 ( \34814 , \34332 );
or \U$34472 ( \34815 , \34813 , \34814 );
not \U$34473 ( \34816 , RIbb2e710_33);
not \U$34474 ( \34817 , \18908 );
or \U$34475 ( \34818 , \34816 , \34817 );
nand \U$34476 ( \34819 , \32817 , \2935 );
nand \U$34477 ( \34820 , \34818 , \34819 );
nand \U$34478 ( \34821 , \34820 , \3886 );
nand \U$34479 ( \34822 , \34815 , \34821 );
xor \U$34480 ( \34823 , \34463 , \34471 );
xor \U$34481 ( \34824 , \34822 , \34823 );
not \U$34482 ( \34825 , \6251 );
not \U$34483 ( \34826 , RIbb2e530_37);
not \U$34484 ( \34827 , \16747 );
or \U$34485 ( \34828 , \34826 , \34827 );
nand \U$34486 ( \34829 , \19077 , \6246 );
nand \U$34487 ( \34830 , \34828 , \34829 );
not \U$34488 ( \34831 , \34830 );
or \U$34489 ( \34832 , \34825 , \34831 );
nand \U$34490 ( \34833 , \34491 , \6241 );
nand \U$34491 ( \34834 , \34832 , \34833 );
and \U$34492 ( \34835 , \34824 , \34834 );
and \U$34493 ( \34836 , \34822 , \34823 );
or \U$34494 ( \34837 , \34835 , \34836 );
not \U$34495 ( \34838 , \16674 );
and \U$34496 ( \34839 , RIbb2dbd0_57, \13876 );
not \U$34497 ( \34840 , RIbb2dbd0_57);
and \U$34498 ( \34841 , \34840 , \26467 );
or \U$34499 ( \34842 , \34839 , \34841 );
not \U$34500 ( \34843 , \34842 );
or \U$34501 ( \34844 , \34838 , \34843 );
nand \U$34502 ( \34845 , \34402 , \17100 );
nand \U$34503 ( \34846 , \34844 , \34845 );
xor \U$34504 ( \34847 , \34837 , \34846 );
not \U$34505 ( \34848 , \17563 );
not \U$34506 ( \34849 , RIbb2ddb0_53);
not \U$34507 ( \34850 , \12194 );
or \U$34508 ( \34851 , \34849 , \34850 );
nand \U$34509 ( \34852 , \13866 , \13463 );
nand \U$34510 ( \34853 , \34851 , \34852 );
not \U$34511 ( \34854 , \34853 );
or \U$34512 ( \34855 , \34848 , \34854 );
nand \U$34513 ( \34856 , \34503 , \14930 );
nand \U$34514 ( \34857 , \34855 , \34856 );
and \U$34515 ( \34858 , \34847 , \34857 );
and \U$34516 ( \34859 , \34837 , \34846 );
or \U$34517 ( \34860 , \34858 , \34859 );
not \U$34518 ( \34861 , \34860 );
or \U$34519 ( \34862 , \34812 , \34861 );
not \U$34520 ( \34863 , \34810 );
nand \U$34521 ( \34864 , \34863 , \34807 );
nand \U$34522 ( \34865 , \34862 , \34864 );
not \U$34523 ( \34866 , \34865 );
or \U$34524 ( \34867 , \34780 , \34866 );
nand \U$34525 ( \34868 , \34774 , \34777 );
nand \U$34526 ( \34869 , \34867 , \34868 );
nand \U$34527 ( \34870 , \34772 , \34869 );
nand \U$34528 ( \34871 , \34771 , \34870 );
not \U$34529 ( \34872 , \34871 );
xor \U$34530 ( \34873 , \34277 , \34283 );
xor \U$34531 ( \34874 , \34873 , \34529 );
nand \U$34532 ( \34875 , \34872 , \34874 );
not \U$34533 ( \34876 , \34875 );
xor \U$34534 ( \34877 , \34386 , \34421 );
xor \U$34535 ( \34878 , \34877 , \34449 );
not \U$34536 ( \34879 , \34878 );
not \U$34537 ( \34880 , \34879 );
not \U$34538 ( \34881 , \34546 );
not \U$34539 ( \34882 , \34881 );
not \U$34540 ( \34883 , \34557 );
or \U$34541 ( \34884 , \34882 , \34883 );
nand \U$34542 ( \34885 , \34556 , \34546 );
nand \U$34543 ( \34886 , \34884 , \34885 );
not \U$34544 ( \34887 , \34595 );
and \U$34545 ( \34888 , \34886 , \34887 );
not \U$34546 ( \34889 , \34886 );
and \U$34547 ( \34890 , \34889 , \34595 );
nor \U$34548 ( \34891 , \34888 , \34890 );
not \U$34549 ( \34892 , \34891 );
or \U$34550 ( \34893 , \34880 , \34892 );
xor \U$34551 ( \34894 , \34472 , \34482 );
xor \U$34552 ( \34895 , \34894 , \34493 );
not \U$34553 ( \34896 , \34895 );
not \U$34554 ( \34897 , \7104 );
not \U$34555 ( \34898 , \34787 );
or \U$34556 ( \34899 , \34897 , \34898 );
not \U$34557 ( \34900 , RIbb2e440_39);
not \U$34558 ( \34901 , \15754 );
or \U$34559 ( \34902 , \34900 , \34901 );
not \U$34560 ( \34903 , RIbb2e440_39);
nand \U$34561 ( \34904 , \34903 , \16566 );
nand \U$34562 ( \34905 , \34902 , \34904 );
nand \U$34563 ( \34906 , \34905 , \7102 );
nand \U$34564 ( \34907 , \34899 , \34906 );
not \U$34565 ( \34908 , \10599 );
and \U$34566 ( \34909 , RIbb2e170_45, \12348 );
not \U$34567 ( \34910 , RIbb2e170_45);
and \U$34568 ( \34911 , \34910 , \16765 );
or \U$34569 ( \34912 , \34909 , \34911 );
not \U$34570 ( \34913 , \34912 );
or \U$34571 ( \34914 , \34908 , \34913 );
not \U$34572 ( \34915 , RIbb2e170_45);
not \U$34573 ( \34916 , \12323 );
or \U$34574 ( \34917 , \34915 , \34916 );
nand \U$34575 ( \34918 , \14635 , \9094 );
nand \U$34576 ( \34919 , \34917 , \34918 );
nand \U$34577 ( \34920 , \34919 , \10119 );
nand \U$34578 ( \34921 , \34914 , \34920 );
xor \U$34579 ( \34922 , \34907 , \34921 );
not \U$34580 ( \34923 , \8362 );
not \U$34581 ( \34924 , RIbb2e350_41);
not \U$34582 ( \34925 , \20577 );
or \U$34583 ( \34926 , \34924 , \34925 );
nand \U$34584 ( \34927 , \34368 , \7097 );
nand \U$34585 ( \34928 , \34926 , \34927 );
not \U$34586 ( \34929 , \34928 );
or \U$34587 ( \34930 , \34923 , \34929 );
not \U$34588 ( \34931 , RIbb2e350_41);
not \U$34589 ( \34932 , \27449 );
or \U$34590 ( \34933 , \34931 , \34932 );
nand \U$34591 ( \34934 , \13977 , \9402 );
nand \U$34592 ( \34935 , \34933 , \34934 );
nand \U$34593 ( \34936 , \34935 , \8354 );
nand \U$34594 ( \34937 , \34930 , \34936 );
and \U$34595 ( \34938 , \34922 , \34937 );
and \U$34596 ( \34939 , \34907 , \34921 );
or \U$34597 ( \34940 , \34938 , \34939 );
not \U$34598 ( \34941 , \34940 );
or \U$34599 ( \34942 , \34896 , \34941 );
or \U$34600 ( \34943 , \34940 , \34895 );
not \U$34601 ( \34944 , \4714 );
not \U$34602 ( \34945 , \34480 );
or \U$34603 ( \34946 , \34944 , \34945 );
not \U$34604 ( \34947 , RIbb2e620_35);
not \U$34605 ( \34948 , \17768 );
or \U$34606 ( \34949 , \34947 , \34948 );
nand \U$34607 ( \34950 , \26039 , \3866 );
nand \U$34608 ( \34951 , \34949 , \34950 );
nand \U$34609 ( \34952 , \34951 , \4712 );
nand \U$34610 ( \34953 , \34946 , \34952 );
and \U$34611 ( \34954 , \17506 , \2941 );
not \U$34612 ( \34955 , \4075 );
not \U$34613 ( \34956 , \34820 );
or \U$34614 ( \34957 , \34955 , \34956 );
not \U$34615 ( \34958 , \20552 );
and \U$34616 ( \34959 , RIbb2e710_33, \34958 );
not \U$34617 ( \34960 , RIbb2e710_33);
and \U$34618 ( \34961 , \34960 , \17745 );
nor \U$34619 ( \34962 , \34959 , \34961 );
nand \U$34620 ( \34963 , \34962 , \3886 );
nand \U$34621 ( \34964 , \34957 , \34963 );
xor \U$34622 ( \34965 , \34954 , \34964 );
not \U$34623 ( \34966 , \4712 );
not \U$34624 ( \34967 , RIbb2e620_35);
not \U$34625 ( \34968 , \17755 );
or \U$34626 ( \34969 , \34967 , \34968 );
nand \U$34627 ( \34970 , \18923 , \6002 );
nand \U$34628 ( \34971 , \34969 , \34970 );
not \U$34629 ( \34972 , \34971 );
or \U$34630 ( \34973 , \34966 , \34972 );
nand \U$34631 ( \34974 , \34951 , \4714 );
nand \U$34632 ( \34975 , \34973 , \34974 );
and \U$34633 ( \34976 , \34965 , \34975 );
and \U$34634 ( \34977 , \34954 , \34964 );
or \U$34635 ( \34978 , \34976 , \34977 );
xor \U$34636 ( \34979 , \34953 , \34978 );
not \U$34637 ( \34980 , \9098 );
not \U$34638 ( \34981 , RIbb2e260_43);
not \U$34639 ( \34982 , \13986 );
or \U$34640 ( \34983 , \34981 , \34982 );
nand \U$34641 ( \34984 , \13547 , \8347 );
nand \U$34642 ( \34985 , \34983 , \34984 );
not \U$34643 ( \34986 , \34985 );
or \U$34644 ( \34987 , \34980 , \34986 );
nand \U$34645 ( \34988 , \34797 , \10451 );
nand \U$34646 ( \34989 , \34987 , \34988 );
and \U$34647 ( \34990 , \34979 , \34989 );
and \U$34648 ( \34991 , \34953 , \34978 );
or \U$34649 ( \34992 , \34990 , \34991 );
nand \U$34650 ( \34993 , \34943 , \34992 );
nand \U$34651 ( \34994 , \34942 , \34993 );
not \U$34652 ( \34995 , \16271 );
and \U$34653 ( \34996 , RIbb2dae0_59, \8388 );
not \U$34654 ( \34997 , RIbb2dae0_59);
and \U$34655 ( \34998 , \34997 , \9110 );
or \U$34656 ( \34999 , \34996 , \34998 );
not \U$34657 ( \35000 , \34999 );
or \U$34658 ( \35001 , \34995 , \35000 );
nand \U$34659 ( \35002 , \34427 , \17470 );
nand \U$34660 ( \35003 , \35001 , \35002 );
not \U$34661 ( \35004 , \12774 );
and \U$34662 ( \35005 , RIbb2dea0_51, \12222 );
not \U$34663 ( \35006 , RIbb2dea0_51);
and \U$34664 ( \35007 , \35006 , \9841 );
or \U$34665 ( \35008 , \35005 , \35007 );
not \U$34666 ( \35009 , \35008 );
or \U$34667 ( \35010 , \35004 , \35009 );
nand \U$34668 ( \35011 , \34565 , \12692 );
nand \U$34669 ( \35012 , \35010 , \35011 );
xor \U$34670 ( \35013 , \35003 , \35012 );
not \U$34671 ( \35014 , \17275 );
not \U$34672 ( \35015 , RIbb2d900_63);
not \U$34673 ( \35016 , \3090 );
or \U$34674 ( \35017 , \35015 , \35016 );
nand \U$34675 ( \35018 , \3091 , \17262 );
nand \U$34676 ( \35019 , \35017 , \35018 );
not \U$34677 ( \35020 , \35019 );
or \U$34678 ( \35021 , \35014 , \35020 );
nand \U$34679 ( \35022 , \34576 , RIbb2d888_64);
nand \U$34680 ( \35023 , \35021 , \35022 );
and \U$34681 ( \35024 , \35013 , \35023 );
and \U$34682 ( \35025 , \35003 , \35012 );
or \U$34683 ( \35026 , \35024 , \35025 );
xor \U$34684 ( \35027 , \34994 , \35026 );
xor \U$34685 ( \35028 , \34593 , \34569 );
xor \U$34686 ( \35029 , \34580 , \35028 );
and \U$34687 ( \35030 , \35027 , \35029 );
and \U$34688 ( \35031 , \34994 , \35026 );
or \U$34689 ( \35032 , \35030 , \35031 );
nand \U$34690 ( \35033 , \34893 , \35032 );
not \U$34691 ( \35034 , \34891 );
nand \U$34692 ( \35035 , \35034 , \34878 );
nand \U$34693 ( \35036 , \35033 , \35035 );
xor \U$34694 ( \35037 , \34353 , \34452 );
xor \U$34695 ( \35038 , \35037 , \34526 );
or \U$34696 ( \35039 , \35036 , \35038 );
xor \U$34697 ( \35040 , \34362 , \34372 );
xor \U$34698 ( \35041 , \35040 , \34383 );
not \U$34699 ( \35042 , \8361 );
not \U$34700 ( \35043 , \34935 );
or \U$34701 ( \35044 , \35042 , \35043 );
nand \U$34702 ( \35045 , \34357 , \8354 );
nand \U$34703 ( \35046 , \35044 , \35045 );
not \U$34704 ( \35047 , \10119 );
not \U$34705 ( \35048 , \34417 );
or \U$34706 ( \35049 , \35047 , \35048 );
nand \U$34707 ( \35050 , \34919 , \10599 );
nand \U$34708 ( \35051 , \35049 , \35050 );
xor \U$34709 ( \35052 , \35046 , \35051 );
not \U$34710 ( \35053 , \12167 );
not \U$34711 ( \35054 , RIbb2df90_49);
not \U$34712 ( \35055 , \12764 );
or \U$34713 ( \35056 , \35054 , \35055 );
nand \U$34714 ( \35057 , \13525 , \12278 );
nand \U$34715 ( \35058 , \35056 , \35057 );
not \U$34716 ( \35059 , \35058 );
or \U$34717 ( \35060 , \35053 , \35059 );
nand \U$34718 ( \35061 , \34439 , \14752 );
nand \U$34719 ( \35062 , \35060 , \35061 );
and \U$34720 ( \35063 , \35052 , \35062 );
and \U$34721 ( \35064 , \35046 , \35051 );
or \U$34722 ( \35065 , \35063 , \35064 );
xor \U$34723 ( \35066 , \35041 , \35065 );
not \U$34724 ( \35067 , \11177 );
not \U$34725 ( \35068 , \34392 );
or \U$34726 ( \35069 , \35067 , \35068 );
not \U$34727 ( \35070 , RIbb2e080_47);
not \U$34728 ( \35071 , \11580 );
or \U$34729 ( \35072 , \35070 , \35071 );
nand \U$34730 ( \35073 , \14885 , \22357 );
nand \U$34731 ( \35074 , \35072 , \35073 );
nand \U$34732 ( \35075 , \35074 , \11176 );
nand \U$34733 ( \35076 , \35069 , \35075 );
not \U$34734 ( \35077 , \35076 );
not \U$34735 ( \35078 , \14613 );
not \U$34736 ( \35079 , \13854 );
not \U$34737 ( \35080 , \34511 );
and \U$34738 ( \35081 , \35079 , \35080 );
and \U$34739 ( \35082 , \13854 , \34511 );
nor \U$34740 ( \35083 , \35081 , \35082 );
nor \U$34741 ( \35084 , \35078 , \35083 );
not \U$34742 ( \35085 , \15181 );
nor \U$34743 ( \35086 , \35085 , \34515 );
nor \U$34744 ( \35087 , \35084 , \35086 );
nand \U$34745 ( \35088 , \35077 , \35087 );
not \U$34746 ( \35089 , \35088 );
not \U$34747 ( \35090 , \16533 );
not \U$34748 ( \35091 , \34589 );
or \U$34749 ( \35092 , \35090 , \35091 );
not \U$34750 ( \35093 , RIbb2d9f0_61);
not \U$34751 ( \35094 , \13560 );
or \U$34752 ( \35095 , \35093 , \35094 );
nand \U$34753 ( \35096 , \20390 , \19746 );
nand \U$34754 ( \35097 , \35095 , \35096 );
nand \U$34755 ( \35098 , \35097 , \18717 );
nand \U$34756 ( \35099 , \35092 , \35098 );
not \U$34757 ( \35100 , \35099 );
or \U$34758 ( \35101 , \35089 , \35100 );
not \U$34759 ( \35102 , \35087 );
nand \U$34760 ( \35103 , \35102 , \35076 );
nand \U$34761 ( \35104 , \35101 , \35103 );
and \U$34762 ( \35105 , \35066 , \35104 );
and \U$34763 ( \35106 , \35041 , \35065 );
or \U$34764 ( \35107 , \35105 , \35106 );
xor \U$34765 ( \35108 , \34496 , \34507 );
xor \U$34766 ( \35109 , \35108 , \34520 );
not \U$34767 ( \35110 , \35109 );
not \U$34768 ( \35111 , \34405 );
and \U$34769 ( \35112 , \34402 , \19101 );
nor \U$34770 ( \35113 , \35111 , \35112 );
and \U$34771 ( \35114 , \34419 , \35113 );
not \U$34772 ( \35115 , \34419 );
and \U$34773 ( \35116 , \35115 , \34406 );
nor \U$34774 ( \35117 , \35114 , \35116 );
xor \U$34775 ( \35118 , \35117 , \34396 );
not \U$34776 ( \35119 , \35118 );
not \U$34777 ( \35120 , \35119 );
or \U$34778 ( \35121 , \35110 , \35120 );
not \U$34779 ( \35122 , \35109 );
not \U$34780 ( \35123 , \35122 );
not \U$34781 ( \35124 , \35118 );
or \U$34782 ( \35125 , \35123 , \35124 );
xor \U$34783 ( \35126 , \34445 , \34441 );
xnor \U$34784 ( \35127 , \35126 , \34431 );
not \U$34785 ( \35128 , \35127 );
nand \U$34786 ( \35129 , \35125 , \35128 );
nand \U$34787 ( \35130 , \35121 , \35129 );
xor \U$34788 ( \35131 , \35107 , \35130 );
xor \U$34789 ( \35132 , \34455 , \34457 );
xor \U$34790 ( \35133 , \35132 , \34523 );
and \U$34791 ( \35134 , \35131 , \35133 );
and \U$34792 ( \35135 , \35107 , \35130 );
or \U$34793 ( \35136 , \35134 , \35135 );
nand \U$34794 ( \35137 , \35039 , \35136 );
nand \U$34795 ( \35138 , \35038 , \35036 );
nand \U$34796 ( \35139 , \35137 , \35138 );
not \U$34797 ( \35140 , \35139 );
or \U$34798 ( \35141 , \34876 , \35140 );
not \U$34799 ( \35142 , \34874 );
nand \U$34800 ( \35143 , \35142 , \34871 );
nand \U$34801 ( \35144 , \35141 , \35143 );
not \U$34802 ( \35145 , \35144 );
xor \U$34803 ( \35146 , \34764 , \35145 );
xor \U$34804 ( \35147 , \34533 , \34266 );
xnor \U$34805 ( \35148 , \35147 , \34612 );
and \U$34806 ( \35149 , \35146 , \35148 );
and \U$34807 ( \35150 , \34764 , \35145 );
or \U$34808 ( \35151 , \35149 , \35150 );
nand \U$34809 ( \35152 , \34762 , \35151 );
not \U$34810 ( \35153 , \34701 );
nor \U$34811 ( \35154 , \34709 , \35153 );
or \U$34812 ( \35155 , \34754 , \35154 );
nand \U$34813 ( \35156 , \34709 , \35153 );
nand \U$34814 ( \35157 , \35155 , \35156 );
not \U$34815 ( \35158 , \35157 );
not \U$34816 ( \35159 , \34651 );
not \U$34817 ( \35160 , \34683 );
or \U$34818 ( \35161 , \35159 , \35160 );
not \U$34819 ( \35162 , \34652 );
not \U$34820 ( \35163 , \34680 );
or \U$34821 ( \35164 , \35162 , \35163 );
nand \U$34822 ( \35165 , \35164 , \34695 );
nand \U$34823 ( \35166 , \35161 , \35165 );
not \U$34824 ( \35167 , \34661 );
not \U$34825 ( \35168 , \34674 );
or \U$34826 ( \35169 , \35167 , \35168 );
not \U$34827 ( \35170 , \34660 );
not \U$34828 ( \35171 , \34673 );
or \U$34829 ( \35172 , \35170 , \35171 );
nand \U$34830 ( \35173 , \35172 , \34658 );
nand \U$34831 ( \35174 , \35169 , \35173 );
xor \U$34832 ( \35175 , \28376 , \28415 );
xor \U$34833 ( \35176 , \35175 , \28461 );
xor \U$34834 ( \35177 , \35174 , \35176 );
xor \U$34835 ( \35178 , \28542 , \28579 );
xor \U$34836 ( \35179 , \35178 , \28605 );
not \U$34837 ( \35180 , \35179 );
and \U$34838 ( \35181 , \35177 , \35180 );
not \U$34839 ( \35182 , \35177 );
and \U$34840 ( \35183 , \35182 , \35179 );
nor \U$34841 ( \35184 , \35181 , \35183 );
not \U$34842 ( \35185 , \35184 );
and \U$34843 ( \35186 , \35166 , \35185 );
not \U$34844 ( \35187 , \35166 );
and \U$34845 ( \35188 , \35187 , \35184 );
nor \U$34846 ( \35189 , \35186 , \35188 );
xor \U$34847 ( \35190 , \28532 , \28534 );
xor \U$34848 ( \35191 , \35190 , \28537 );
xor \U$34849 ( \35192 , \34687 , \34691 );
and \U$34850 ( \35193 , \35192 , \34694 );
and \U$34851 ( \35194 , \34687 , \34691 );
or \U$34852 ( \35195 , \35193 , \35194 );
xor \U$34853 ( \35196 , \35191 , \35195 );
xor \U$34854 ( \35197 , \28611 , \28613 );
xor \U$34855 ( \35198 , \35197 , \28689 );
xor \U$34856 ( \35199 , \35196 , \35198 );
not \U$34857 ( \35200 , \35199 );
and \U$34858 ( \35201 , \35189 , \35200 );
not \U$34859 ( \35202 , \35189 );
and \U$34860 ( \35203 , \35202 , \35199 );
nor \U$34861 ( \35204 , \35201 , \35203 );
not \U$34862 ( \35205 , \34746 );
not \U$34863 ( \35206 , \34717 );
or \U$34864 ( \35207 , \35205 , \35206 );
not \U$34865 ( \35208 , \34717 );
not \U$34866 ( \35209 , \35208 );
not \U$34867 ( \35210 , \34745 );
or \U$34868 ( \35211 , \35209 , \35210 );
nand \U$34869 ( \35212 , \35211 , \34753 );
nand \U$34870 ( \35213 , \35207 , \35212 );
not \U$34871 ( \35214 , \35213 );
xor \U$34872 ( \35215 , \35204 , \35214 );
not \U$34873 ( \35216 , \34744 );
not \U$34874 ( \35217 , \34724 );
nand \U$34875 ( \35218 , \35217 , \34736 );
not \U$34876 ( \35219 , \35218 );
or \U$34877 ( \35220 , \35216 , \35219 );
nand \U$34878 ( \35221 , \34737 , \34724 );
nand \U$34879 ( \35222 , \35220 , \35221 );
not \U$34880 ( \35223 , \35222 );
not \U$34881 ( \35224 , \35223 );
not \U$34882 ( \35225 , \34730 );
not \U$34883 ( \35226 , \34728 );
nand \U$34884 ( \35227 , \35225 , \35226 );
not \U$34885 ( \35228 , \35227 );
not \U$34886 ( \35229 , \34735 );
or \U$34887 ( \35230 , \35228 , \35229 );
not \U$34888 ( \35231 , \35226 );
nand \U$34889 ( \35232 , \35231 , \34730 );
nand \U$34890 ( \35233 , \35230 , \35232 );
not \U$34891 ( \35234 , \35233 );
not \U$34892 ( \35235 , \35234 );
not \U$34893 ( \35236 , \28788 );
not \U$34894 ( \35237 , \28898 );
not \U$34895 ( \35238 , \35237 );
or \U$34896 ( \35239 , \35236 , \35238 );
not \U$34897 ( \35240 , \28788 );
nand \U$34898 ( \35241 , \35240 , \28898 );
nand \U$34899 ( \35242 , \35239 , \35241 );
not \U$34900 ( \35243 , \28790 );
and \U$34901 ( \35244 , \35242 , \35243 );
not \U$34902 ( \35245 , \35242 );
and \U$34903 ( \35246 , \35245 , \28790 );
nor \U$34904 ( \35247 , \35244 , \35246 );
not \U$34905 ( \35248 , \35247 );
not \U$34906 ( \35249 , \35248 );
or \U$34907 ( \35250 , \35235 , \35249 );
nand \U$34908 ( \35251 , \35247 , \35233 );
nand \U$34909 ( \35252 , \35250 , \35251 );
not \U$34910 ( \35253 , \34642 );
nand \U$34911 ( \35254 , \34630 , \34633 );
not \U$34912 ( \35255 , \35254 );
or \U$34913 ( \35256 , \35253 , \35255 );
not \U$34914 ( \35257 , \34630 );
nand \U$34915 ( \35258 , \35257 , \34634 );
nand \U$34916 ( \35259 , \35256 , \35258 );
not \U$34917 ( \35260 , \35259 );
and \U$34918 ( \35261 , \35252 , \35260 );
not \U$34919 ( \35262 , \35252 );
and \U$34920 ( \35263 , \35262 , \35259 );
nor \U$34921 ( \35264 , \35261 , \35263 );
not \U$34922 ( \35265 , \35264 );
not \U$34923 ( \35266 , \35265 );
or \U$34924 ( \35267 , \35224 , \35266 );
nand \U$34925 ( \35268 , \35264 , \35222 );
nand \U$34926 ( \35269 , \35267 , \35268 );
not \U$34927 ( \35270 , \34628 );
not \U$34928 ( \35271 , \34643 );
not \U$34929 ( \35272 , \35271 );
or \U$34930 ( \35273 , \35270 , \35272 );
or \U$34931 ( \35274 , \35271 , \34628 );
nand \U$34932 ( \35275 , \35274 , \34700 );
nand \U$34933 ( \35276 , \35273 , \35275 );
not \U$34934 ( \35277 , \35276 );
and \U$34935 ( \35278 , \35269 , \35277 );
not \U$34936 ( \35279 , \35269 );
and \U$34937 ( \35280 , \35279 , \35276 );
nor \U$34938 ( \35281 , \35278 , \35280 );
xor \U$34939 ( \35282 , \35215 , \35281 );
nand \U$34940 ( \35283 , \35158 , \35282 );
and \U$34941 ( \35284 , \34622 , \34760 , \35152 , \35283 );
not \U$34942 ( \35285 , \35284 );
not \U$34943 ( \35286 , \35285 );
and \U$34944 ( \35287 , \28363 , \28917 );
not \U$34945 ( \35288 , \28363 );
not \U$34946 ( \35289 , \28917 );
and \U$34947 ( \35290 , \35288 , \35289 );
nor \U$34948 ( \35291 , \35287 , \35290 );
and \U$34949 ( \35292 , \35291 , \28370 );
not \U$34950 ( \35293 , \35291 );
and \U$34951 ( \35294 , \35293 , \28920 );
nor \U$34952 ( \35295 , \35292 , \35294 );
xor \U$34953 ( \35296 , \28484 , \28912 );
xor \U$34954 ( \35297 , \35296 , \28915 );
not \U$34955 ( \35298 , \35297 );
not \U$34956 ( \35299 , \27428 );
not \U$34957 ( \35300 , \27420 );
or \U$34958 ( \35301 , \35299 , \35300 );
nand \U$34959 ( \35302 , \27419 , \27425 );
nand \U$34960 ( \35303 , \35301 , \35302 );
not \U$34961 ( \35304 , \27473 );
and \U$34962 ( \35305 , \35303 , \35304 );
not \U$34963 ( \35306 , \35303 );
and \U$34964 ( \35307 , \35306 , \27473 );
nor \U$34965 ( \35308 , \35305 , \35307 );
not \U$34966 ( \35309 , \35308 );
not \U$34967 ( \35310 , \28474 );
not \U$34968 ( \35311 , \28464 );
not \U$34969 ( \35312 , \35311 );
or \U$34970 ( \35313 , \35310 , \35312 );
nand \U$34971 ( \35314 , \28473 , \28464 );
nand \U$34972 ( \35315 , \35313 , \35314 );
not \U$34973 ( \35316 , \28467 );
and \U$34974 ( \35317 , \35315 , \35316 );
not \U$34975 ( \35318 , \35315 );
and \U$34976 ( \35319 , \35318 , \28467 );
nor \U$34977 ( \35320 , \35317 , \35319 );
not \U$34978 ( \35321 , \35320 );
or \U$34979 ( \35322 , \35309 , \35321 );
not \U$34980 ( \35323 , \35179 );
nor \U$34981 ( \35324 , \35174 , \35176 );
not \U$34982 ( \35325 , \35324 );
not \U$34983 ( \35326 , \35325 );
or \U$34984 ( \35327 , \35323 , \35326 );
nand \U$34985 ( \35328 , \35174 , \35176 );
nand \U$34986 ( \35329 , \35327 , \35328 );
nand \U$34987 ( \35330 , \35322 , \35329 );
not \U$34988 ( \35331 , \35308 );
not \U$34989 ( \35332 , \35320 );
nand \U$34990 ( \35333 , \35331 , \35332 );
nand \U$34991 ( \35334 , \35330 , \35333 );
buf \U$34992 ( \35335 , \35334 );
not \U$34993 ( \35336 , \35335 );
xor \U$34994 ( \35337 , \28476 , \28478 );
xor \U$34995 ( \35338 , \35337 , \28481 );
not \U$34996 ( \35339 , \35338 );
or \U$34997 ( \35340 , \35336 , \35339 );
or \U$34998 ( \35341 , \35338 , \35335 );
xor \U$34999 ( \35342 , \28540 , \28608 );
xor \U$35000 ( \35343 , \35342 , \28692 );
not \U$35001 ( \35344 , \35343 );
not \U$35002 ( \35345 , \35191 );
not \U$35003 ( \35346 , \35198 );
or \U$35004 ( \35347 , \35345 , \35346 );
or \U$35005 ( \35348 , \35198 , \35191 );
nand \U$35006 ( \35349 , \35348 , \35195 );
nand \U$35007 ( \35350 , \35347 , \35349 );
not \U$35008 ( \35351 , \35350 );
or \U$35009 ( \35352 , \35344 , \35351 );
or \U$35010 ( \35353 , \35343 , \35350 );
xor \U$35011 ( \35354 , \28698 , \28709 );
xor \U$35012 ( \35355 , \35354 , \28902 );
nand \U$35013 ( \35356 , \35353 , \35355 );
nand \U$35014 ( \35357 , \35352 , \35356 );
nand \U$35015 ( \35358 , \35341 , \35357 );
nand \U$35016 ( \35359 , \35340 , \35358 );
not \U$35017 ( \35360 , \35359 );
xor \U$35018 ( \35361 , \27127 , \27339 );
xnor \U$35019 ( \35362 , \35361 , \27327 );
nand \U$35020 ( \35363 , \35360 , \35362 );
not \U$35021 ( \35364 , \35363 );
or \U$35022 ( \35365 , \35298 , \35364 );
not \U$35023 ( \35366 , \35362 );
nand \U$35024 ( \35367 , \35366 , \35359 );
nand \U$35025 ( \35368 , \35365 , \35367 );
not \U$35026 ( \35369 , \35368 );
nand \U$35027 ( \35370 , \35295 , \35369 );
not \U$35028 ( \35371 , \35359 );
not \U$35029 ( \35372 , \35362 );
or \U$35030 ( \35373 , \35371 , \35372 );
or \U$35031 ( \35374 , \35359 , \35362 );
nand \U$35032 ( \35375 , \35373 , \35374 );
not \U$35033 ( \35376 , \35297 );
and \U$35034 ( \35377 , \35375 , \35376 );
not \U$35035 ( \35378 , \35375 );
and \U$35036 ( \35379 , \35378 , \35297 );
nor \U$35037 ( \35380 , \35377 , \35379 );
xor \U$35038 ( \35381 , \28905 , \28695 );
not \U$35039 ( \35382 , \28910 );
xor \U$35040 ( \35383 , \35381 , \35382 );
not \U$35041 ( \35384 , \35233 );
not \U$35042 ( \35385 , \35247 );
not \U$35043 ( \35386 , \35385 );
or \U$35044 ( \35387 , \35384 , \35386 );
or \U$35045 ( \35388 , \35385 , \35233 );
nand \U$35046 ( \35389 , \35388 , \35259 );
nand \U$35047 ( \35390 , \35387 , \35389 );
not \U$35048 ( \35391 , \35390 );
not \U$35049 ( \35392 , \35391 );
xor \U$35050 ( \35393 , \35308 , \35329 );
xor \U$35051 ( \35394 , \35393 , \35332 );
not \U$35052 ( \35395 , \35394 );
or \U$35053 ( \35396 , \35392 , \35395 );
not \U$35054 ( \35397 , \35199 );
not \U$35055 ( \35398 , \35166 );
nand \U$35056 ( \35399 , \35398 , \35184 );
not \U$35057 ( \35400 , \35399 );
or \U$35058 ( \35401 , \35397 , \35400 );
nand \U$35059 ( \35402 , \35185 , \35166 );
nand \U$35060 ( \35403 , \35401 , \35402 );
nand \U$35061 ( \35404 , \35396 , \35403 );
not \U$35062 ( \35405 , \35394 );
nand \U$35063 ( \35406 , \35405 , \35390 );
and \U$35064 ( \35407 , \35404 , \35406 );
xor \U$35065 ( \35408 , \35383 , \35407 );
xor \U$35066 ( \35409 , \35334 , \35357 );
xnor \U$35067 ( \35410 , \35409 , \35338 );
and \U$35068 ( \35411 , \35408 , \35410 );
and \U$35069 ( \35412 , \35383 , \35407 );
or \U$35070 ( \35413 , \35411 , \35412 );
nand \U$35071 ( \35414 , \35380 , \35413 );
nand \U$35072 ( \35415 , \35370 , \35414 );
xor \U$35073 ( \35416 , \35343 , \35350 );
not \U$35074 ( \35417 , \35355 );
xor \U$35075 ( \35418 , \35416 , \35417 );
not \U$35076 ( \35419 , \35222 );
not \U$35077 ( \35420 , \35265 );
or \U$35078 ( \35421 , \35419 , \35420 );
nand \U$35079 ( \35422 , \35264 , \35223 );
nand \U$35080 ( \35423 , \35276 , \35422 );
nand \U$35081 ( \35424 , \35421 , \35423 );
not \U$35082 ( \35425 , \35424 );
xor \U$35083 ( \35426 , \35418 , \35425 );
xor \U$35084 ( \35427 , \35390 , \35405 );
xnor \U$35085 ( \35428 , \35427 , \35403 );
and \U$35086 ( \35429 , \35426 , \35428 );
and \U$35087 ( \35430 , \35418 , \35425 );
or \U$35088 ( \35431 , \35429 , \35430 );
not \U$35089 ( \35432 , \35431 );
xor \U$35090 ( \35433 , \35383 , \35407 );
xor \U$35091 ( \35434 , \35433 , \35410 );
not \U$35092 ( \35435 , \35434 );
or \U$35093 ( \35436 , \35432 , \35435 );
xor \U$35094 ( \35437 , \35418 , \35425 );
xor \U$35095 ( \35438 , \35437 , \35428 );
xor \U$35096 ( \35439 , \35204 , \35214 );
and \U$35097 ( \35440 , \35439 , \35281 );
and \U$35098 ( \35441 , \35204 , \35214 );
or \U$35099 ( \35442 , \35440 , \35441 );
nand \U$35100 ( \35443 , \35438 , \35442 );
nand \U$35101 ( \35444 , \35436 , \35443 );
nor \U$35102 ( \35445 , \35415 , \35444 );
buf \U$35103 ( \35446 , \35445 );
or \U$35104 ( \35447 , RIbb2e698_34, RIbb2e620_35);
nand \U$35105 ( \35448 , \35447 , \17506 );
and \U$35106 ( \35449 , RIbb2e698_34, RIbb2e620_35);
nor \U$35107 ( \35450 , \35449 , \2935 );
and \U$35108 ( \35451 , \35448 , \35450 );
not \U$35109 ( \35452 , \4075 );
not \U$35110 ( \35453 , \34962 );
or \U$35111 ( \35454 , \35452 , \35453 );
and \U$35112 ( \35455 , RIbb2e710_33, \17506 );
not \U$35113 ( \35456 , RIbb2e710_33);
and \U$35114 ( \35457 , \35456 , \20747 );
nor \U$35115 ( \35458 , \35455 , \35457 );
nand \U$35116 ( \35459 , \35458 , \3885 );
nand \U$35117 ( \35460 , \35454 , \35459 );
xor \U$35118 ( \35461 , \35451 , \35460 );
not \U$35119 ( \35462 , \4714 );
not \U$35120 ( \35463 , \34971 );
or \U$35121 ( \35464 , \35462 , \35463 );
not \U$35122 ( \35465 , RIbb2e620_35);
not \U$35123 ( \35466 , \32817 );
not \U$35124 ( \35467 , \35466 );
or \U$35125 ( \35468 , \35465 , \35467 );
nand \U$35126 ( \35469 , \32817 , \6002 );
nand \U$35127 ( \35470 , \35468 , \35469 );
nand \U$35128 ( \35471 , \35470 , \4712 );
nand \U$35129 ( \35472 , \35464 , \35471 );
xor \U$35130 ( \35473 , \35461 , \35472 );
not \U$35131 ( \35474 , \7102 );
and \U$35132 ( \35475 , RIbb2e440_39, \16747 );
not \U$35133 ( \35476 , RIbb2e440_39);
and \U$35134 ( \35477 , \35476 , \18093 );
or \U$35135 ( \35478 , \35475 , \35477 );
not \U$35136 ( \35479 , \35478 );
or \U$35137 ( \35480 , \35474 , \35479 );
and \U$35138 ( \35481 , RIbb2e440_39, \15824 );
not \U$35139 ( \35482 , RIbb2e440_39);
and \U$35140 ( \35483 , \35482 , \16575 );
or \U$35141 ( \35484 , \35481 , \35483 );
nand \U$35142 ( \35485 , \35484 , \7104 );
nand \U$35143 ( \35486 , \35480 , \35485 );
xor \U$35144 ( \35487 , \35473 , \35486 );
not \U$35145 ( \35488 , \16427 );
not \U$35146 ( \35489 , RIbb2df90_49);
not \U$35147 ( \35490 , \11580 );
or \U$35148 ( \35491 , \35489 , \35490 );
nand \U$35149 ( \35492 , \14885 , \12278 );
nand \U$35150 ( \35493 , \35491 , \35492 );
not \U$35151 ( \35494 , \35493 );
or \U$35152 ( \35495 , \35488 , \35494 );
not \U$35153 ( \35496 , RIbb2df90_49);
not \U$35154 ( \35497 , \12839 );
or \U$35155 ( \35498 , \35496 , \35497 );
nand \U$35156 ( \35499 , \12175 , \12278 );
nand \U$35157 ( \35500 , \35498 , \35499 );
nand \U$35158 ( \35501 , \35500 , \13295 );
nand \U$35159 ( \35502 , \35495 , \35501 );
xor \U$35160 ( \35503 , \35487 , \35502 );
and \U$35161 ( \35504 , RIbb2d9f0_61, \8388 );
not \U$35162 ( \35505 , RIbb2d9f0_61);
and \U$35163 ( \35506 , \35505 , \9110 );
or \U$35164 ( \35507 , \35504 , \35506 );
not \U$35165 ( \35508 , \35507 );
not \U$35166 ( \35509 , \26834 );
or \U$35167 ( \35510 , \35508 , \35509 );
not \U$35168 ( \35511 , \5955 );
not \U$35169 ( \35512 , \16254 );
and \U$35170 ( \35513 , \35511 , \35512 );
and \U$35171 ( \35514 , \5955 , \16254 );
nor \U$35172 ( \35515 , \35513 , \35514 );
or \U$35173 ( \35516 , \35515 , \16542 );
nand \U$35174 ( \35517 , \35510 , \35516 );
xor \U$35175 ( \35518 , \35503 , \35517 );
not \U$35176 ( \35519 , \35518 );
not \U$35177 ( \35520 , \21882 );
not \U$35178 ( \35521 , \16601 );
not \U$35179 ( \35522 , \35521 );
or \U$35180 ( \35523 , \35520 , \35522 );
not \U$35181 ( \35524 , \16604 );
nand \U$35182 ( \35525 , \35524 , RIbb2dea0_51);
nand \U$35183 ( \35526 , \35523 , \35525 );
and \U$35184 ( \35527 , \12692 , \35526 );
and \U$35185 ( \35528 , RIbb2dea0_51, \11580 );
not \U$35186 ( \35529 , RIbb2dea0_51);
and \U$35187 ( \35530 , \35529 , \11581 );
or \U$35188 ( \35531 , \35528 , \35530 );
and \U$35189 ( \35532 , \35531 , \14067 );
nor \U$35190 ( \35533 , \35527 , \35532 );
or \U$35191 ( \35534 , RIbb2e5a8_36, RIbb2e530_37);
nand \U$35192 ( \35535 , \35534 , \17506 );
and \U$35193 ( \35536 , RIbb2e5a8_36, RIbb2e530_37);
nor \U$35194 ( \35537 , \35536 , \6002 );
and \U$35195 ( \35538 , \35535 , \35537 );
not \U$35196 ( \35539 , \4710 );
not \U$35197 ( \35540 , RIbb2e620_35);
not \U$35198 ( \35541 , \20552 );
or \U$35199 ( \35542 , \35540 , \35541 );
nand \U$35200 ( \35543 , \26129 , \6002 );
nand \U$35201 ( \35544 , \35542 , \35543 );
not \U$35202 ( \35545 , \35544 );
or \U$35203 ( \35546 , \35539 , \35545 );
or \U$35204 ( \35547 , \17506 , \3866 );
or \U$35205 ( \35548 , \18929 , RIbb2e620_35);
nand \U$35206 ( \35549 , \35547 , \35548 );
nand \U$35207 ( \35550 , \35549 , \4711 );
nand \U$35208 ( \35551 , \35546 , \35550 );
and \U$35209 ( \35552 , \35538 , \35551 );
not \U$35210 ( \35553 , \7104 );
not \U$35211 ( \35554 , \35478 );
or \U$35212 ( \35555 , \35553 , \35554 );
and \U$35213 ( \35556 , RIbb2e440_39, \32993 );
not \U$35214 ( \35557 , RIbb2e440_39);
and \U$35215 ( \35558 , \35557 , \32996 );
or \U$35216 ( \35559 , \35556 , \35558 );
nand \U$35217 ( \35560 , \35559 , \7102 );
nand \U$35218 ( \35561 , \35555 , \35560 );
xor \U$35219 ( \35562 , \35552 , \35561 );
not \U$35220 ( \35563 , \8354 );
not \U$35221 ( \35564 , RIbb2e350_41);
not \U$35222 ( \35565 , \16567 );
or \U$35223 ( \35566 , \35564 , \35565 );
nand \U$35224 ( \35567 , \23098 , \9402 );
nand \U$35225 ( \35568 , \35566 , \35567 );
not \U$35226 ( \35569 , \35568 );
or \U$35227 ( \35570 , \35563 , \35569 );
not \U$35228 ( \35571 , \16576 );
not \U$35229 ( \35572 , \8357 );
and \U$35230 ( \35573 , \35571 , \35572 );
and \U$35231 ( \35574 , \15825 , \7097 );
nor \U$35232 ( \35575 , \35573 , \35574 );
not \U$35233 ( \35576 , \35575 );
nand \U$35234 ( \35577 , \35576 , \8362 );
nand \U$35235 ( \35578 , \35570 , \35577 );
xor \U$35236 ( \35579 , \35562 , \35578 );
not \U$35237 ( \35580 , \35579 );
nand \U$35238 ( \35581 , \35533 , \35580 );
not \U$35239 ( \35582 , \7104 );
not \U$35240 ( \35583 , \35559 );
or \U$35241 ( \35584 , \35582 , \35583 );
xnor \U$35242 ( \35585 , RIbb2e440_39, \34293 );
nand \U$35243 ( \35586 , \35585 , \7102 );
nand \U$35244 ( \35587 , \35584 , \35586 );
and \U$35245 ( \35588 , \17506 , \4714 );
not \U$35246 ( \35589 , \6241 );
not \U$35247 ( \35590 , RIbb2e530_37);
not \U$35248 ( \35591 , \16820 );
or \U$35249 ( \35592 , \35590 , \35591 );
nand \U$35250 ( \35593 , \32817 , \8701 );
nand \U$35251 ( \35594 , \35592 , \35593 );
not \U$35252 ( \35595 , \35594 );
or \U$35253 ( \35596 , \35589 , \35595 );
not \U$35254 ( \35597 , \26129 );
not \U$35255 ( \35598 , \35597 );
and \U$35256 ( \35599 , RIbb2e530_37, \35598 );
not \U$35257 ( \35600 , RIbb2e530_37);
not \U$35258 ( \35601 , \26129 );
and \U$35259 ( \35602 , \35600 , \35601 );
nor \U$35260 ( \35603 , \35599 , \35602 );
nand \U$35261 ( \35604 , \35603 , \6250 );
nand \U$35262 ( \35605 , \35596 , \35604 );
xor \U$35263 ( \35606 , \35588 , \35605 );
not \U$35264 ( \35607 , \7102 );
not \U$35265 ( \35608 , RIbb2e440_39);
not \U$35266 ( \35609 , \27234 );
or \U$35267 ( \35610 , \35608 , \35609 );
not \U$35268 ( \35611 , RIbb2e440_39);
nand \U$35269 ( \35612 , \35611 , \18920 );
nand \U$35270 ( \35613 , \35610 , \35612 );
not \U$35271 ( \35614 , \35613 );
or \U$35272 ( \35615 , \35607 , \35614 );
nand \U$35273 ( \35616 , \35585 , \7104 );
nand \U$35274 ( \35617 , \35615 , \35616 );
and \U$35275 ( \35618 , \35606 , \35617 );
and \U$35276 ( \35619 , \35588 , \35605 );
or \U$35277 ( \35620 , \35618 , \35619 );
xor \U$35278 ( \35621 , \35587 , \35620 );
not \U$35279 ( \35622 , \11176 );
not \U$35280 ( \35623 , RIbb2e080_47);
not \U$35281 ( \35624 , \13546 );
or \U$35282 ( \35625 , \35623 , \35624 );
nand \U$35283 ( \35626 , \15055 , \12971 );
nand \U$35284 ( \35627 , \35625 , \35626 );
not \U$35285 ( \35628 , \35627 );
or \U$35286 ( \35629 , \35622 , \35628 );
not \U$35287 ( \35630 , RIbb2e080_47);
not \U$35288 ( \35631 , \15761 );
or \U$35289 ( \35632 , \35630 , \35631 );
buf \U$35290 ( \35633 , \26964 );
nand \U$35291 ( \35634 , \35633 , \11959 );
nand \U$35292 ( \35635 , \35632 , \35634 );
nand \U$35293 ( \35636 , \35635 , \12965 );
nand \U$35294 ( \35637 , \35629 , \35636 );
and \U$35295 ( \35638 , \35621 , \35637 );
and \U$35296 ( \35639 , \35587 , \35620 );
or \U$35297 ( \35640 , \35638 , \35639 );
and \U$35298 ( \35641 , \35581 , \35640 );
nor \U$35299 ( \35642 , \35533 , \35580 );
nor \U$35300 ( \35643 , \35641 , \35642 );
nand \U$35301 ( \35644 , \35519 , \35643 );
not \U$35302 ( \35645 , \35644 );
and \U$35303 ( \35646 , \17506 , \4075 );
not \U$35304 ( \35647 , \4710 );
not \U$35305 ( \35648 , \35470 );
or \U$35306 ( \35649 , \35647 , \35648 );
nand \U$35307 ( \35650 , \35544 , \4712 );
nand \U$35308 ( \35651 , \35649 , \35650 );
xor \U$35309 ( \35652 , \35646 , \35651 );
not \U$35310 ( \35653 , \6250 );
not \U$35311 ( \35654 , RIbb2e530_37);
not \U$35312 ( \35655 , \17756 );
or \U$35313 ( \35656 , \35654 , \35655 );
nand \U$35314 ( \35657 , \18923 , \4708 );
nand \U$35315 ( \35658 , \35656 , \35657 );
not \U$35316 ( \35659 , \35658 );
or \U$35317 ( \35660 , \35653 , \35659 );
not \U$35318 ( \35661 , RIbb2e530_37);
not \U$35319 ( \35662 , \34293 );
or \U$35320 ( \35663 , \35661 , \35662 );
nand \U$35321 ( \35664 , \16706 , \4708 );
nand \U$35322 ( \35665 , \35663 , \35664 );
nand \U$35323 ( \35666 , \35665 , \6240 );
nand \U$35324 ( \35667 , \35660 , \35666 );
xor \U$35325 ( \35668 , \35652 , \35667 );
not \U$35326 ( \35669 , \11177 );
not \U$35327 ( \35670 , RIbb2e080_47);
not \U$35328 ( \35671 , \21756 );
or \U$35329 ( \35672 , \35670 , \35671 );
nand \U$35330 ( \35673 , \14844 , \12971 );
nand \U$35331 ( \35674 , \35672 , \35673 );
not \U$35332 ( \35675 , \35674 );
or \U$35333 ( \35676 , \35669 , \35675 );
nand \U$35334 ( \35677 , \35635 , \11176 );
nand \U$35335 ( \35678 , \35676 , \35677 );
xor \U$35336 ( \35679 , \35668 , \35678 );
not \U$35337 ( \35680 , \10117 );
not \U$35338 ( \35681 , RIbb2e170_45);
not \U$35339 ( \35682 , \13980 );
not \U$35340 ( \35683 , \35682 );
or \U$35341 ( \35684 , \35681 , \35683 );
not \U$35342 ( \35685 , \15456 );
nand \U$35343 ( \35686 , \35685 , \9094 );
nand \U$35344 ( \35687 , \35684 , \35686 );
not \U$35345 ( \35688 , \35687 );
or \U$35346 ( \35689 , \35680 , \35688 );
not \U$35347 ( \35690 , RIbb2e170_45);
not \U$35348 ( \35691 , \17315 );
or \U$35349 ( \35692 , \35690 , \35691 );
nand \U$35350 ( \35693 , \13989 , \12003 );
nand \U$35351 ( \35694 , \35692 , \35693 );
nand \U$35352 ( \35695 , \35694 , \10119 );
nand \U$35353 ( \35696 , \35689 , \35695 );
xor \U$35354 ( \35697 , \35679 , \35696 );
not \U$35355 ( \35698 , \12692 );
not \U$35356 ( \35699 , \35531 );
or \U$35357 ( \35700 , \35698 , \35699 );
and \U$35358 ( \35701 , RIbb2dea0_51, \13680 );
not \U$35359 ( \35702 , RIbb2dea0_51);
and \U$35360 ( \35703 , \35702 , \22073 );
or \U$35361 ( \35704 , \35701 , \35703 );
nand \U$35362 ( \35705 , \35704 , \14067 );
nand \U$35363 ( \35706 , \35700 , \35705 );
not \U$35364 ( \35707 , \35706 );
and \U$35365 ( \35708 , RIbb2dae0_59, \12801 );
not \U$35366 ( \35709 , RIbb2dae0_59);
and \U$35367 ( \35710 , \35709 , \9819 );
nor \U$35368 ( \35711 , \35708 , \35710 );
not \U$35369 ( \35712 , \35711 );
not \U$35370 ( \35713 , \29399 );
and \U$35371 ( \35714 , \35712 , \35713 );
not \U$35372 ( \35715 , RIbb2dae0_59);
not \U$35373 ( \35716 , \11232 );
or \U$35374 ( \35717 , \35715 , \35716 );
nand \U$35375 ( \35718 , \9074 , \17024 );
nand \U$35376 ( \35719 , \35717 , \35718 );
and \U$35377 ( \35720 , \35719 , \17470 );
nor \U$35378 ( \35721 , \35714 , \35720 );
not \U$35379 ( \35722 , \35721 );
not \U$35380 ( \35723 , \35722 );
or \U$35381 ( \35724 , \35707 , \35723 );
not \U$35382 ( \35725 , \35721 );
not \U$35383 ( \35726 , \35706 );
not \U$35384 ( \35727 , \35726 );
or \U$35385 ( \35728 , \35725 , \35727 );
not \U$35386 ( \35729 , \13467 );
not \U$35387 ( \35730 , RIbb2ddb0_53);
not \U$35388 ( \35731 , \15188 );
or \U$35389 ( \35732 , \35730 , \35731 );
nand \U$35390 ( \35733 , \16604 , \26750 );
nand \U$35391 ( \35734 , \35732 , \35733 );
not \U$35392 ( \35735 , \35734 );
or \U$35393 ( \35736 , \35729 , \35735 );
not \U$35394 ( \35737 , RIbb2ddb0_53);
not \U$35395 ( \35738 , \12249 );
or \U$35396 ( \35739 , \35737 , \35738 );
nand \U$35397 ( \35740 , \10764 , \13941 );
nand \U$35398 ( \35741 , \35739 , \35740 );
nand \U$35399 ( \35742 , \35741 , \14930 );
nand \U$35400 ( \35743 , \35736 , \35742 );
nand \U$35401 ( \35744 , \35728 , \35743 );
nand \U$35402 ( \35745 , \35724 , \35744 );
xor \U$35403 ( \35746 , \35697 , \35745 );
or \U$35404 ( \35747 , RIbb2e4b8_38, RIbb2e440_39);
nand \U$35405 ( \35748 , \35747 , \17506 );
and \U$35406 ( \35749 , RIbb2e4b8_38, RIbb2e440_39);
nor \U$35407 ( \35750 , \35749 , \4708 );
and \U$35408 ( \35751 , \35748 , \35750 );
not \U$35409 ( \35752 , \6250 );
or \U$35410 ( \35753 , \17506 , \6246 );
or \U$35411 ( \35754 , \20747 , RIbb2e530_37);
nand \U$35412 ( \35755 , \35753 , \35754 );
not \U$35413 ( \35756 , \35755 );
or \U$35414 ( \35757 , \35752 , \35756 );
nand \U$35415 ( \35758 , \35603 , \6240 );
nand \U$35416 ( \35759 , \35757 , \35758 );
and \U$35417 ( \35760 , \35751 , \35759 );
not \U$35418 ( \35761 , \8361 );
not \U$35419 ( \35762 , RIbb2e350_41);
buf \U$35420 ( \35763 , \16727 );
not \U$35421 ( \35764 , \35763 );
or \U$35422 ( \35765 , \35762 , \35764 );
nand \U$35423 ( \35766 , \19831 , \8357 );
nand \U$35424 ( \35767 , \35765 , \35766 );
not \U$35425 ( \35768 , \35767 );
or \U$35426 ( \35769 , \35761 , \35768 );
not \U$35427 ( \35770 , \16751 );
not \U$35428 ( \35771 , \7097 );
and \U$35429 ( \35772 , \35770 , \35771 );
and \U$35430 ( \35773 , \18093 , \8357 );
nor \U$35431 ( \35774 , \35772 , \35773 );
not \U$35432 ( \35775 , \35774 );
nand \U$35433 ( \35776 , \35775 , \8354 );
nand \U$35434 ( \35777 , \35769 , \35776 );
xor \U$35435 ( \35778 , \35760 , \35777 );
not \U$35436 ( \35779 , \9099 );
not \U$35437 ( \35780 , RIbb2e260_43);
not \U$35438 ( \35781 , \15754 );
or \U$35439 ( \35782 , \35780 , \35781 );
nand \U$35440 ( \35783 , \15753 , \17231 );
nand \U$35441 ( \35784 , \35782 , \35783 );
not \U$35442 ( \35785 , \35784 );
or \U$35443 ( \35786 , \35779 , \35785 );
not \U$35444 ( \35787 , RIbb2e260_43);
not \U$35445 ( \35788 , \15824 );
or \U$35446 ( \35789 , \35787 , \35788 );
nand \U$35447 ( \35790 , \16576 , \26255 );
nand \U$35448 ( \35791 , \35789 , \35790 );
nand \U$35449 ( \35792 , \35791 , \9098 );
nand \U$35450 ( \35793 , \35786 , \35792 );
and \U$35451 ( \35794 , \35778 , \35793 );
and \U$35452 ( \35795 , \35760 , \35777 );
or \U$35453 ( \35796 , \35794 , \35795 );
not \U$35454 ( \35797 , \14613 );
not \U$35455 ( \35798 , RIbb2dcc0_55);
not \U$35456 ( \35799 , \12234 );
or \U$35457 ( \35800 , \35798 , \35799 );
or \U$35458 ( \35801 , \12744 , RIbb2dcc0_55);
nand \U$35459 ( \35802 , \35800 , \35801 );
not \U$35460 ( \35803 , \35802 );
or \U$35461 ( \35804 , \35797 , \35803 );
and \U$35462 ( \35805 , RIbb2dcc0_55, \22580 );
not \U$35463 ( \35806 , RIbb2dcc0_55);
and \U$35464 ( \35807 , \35806 , \9841 );
or \U$35465 ( \35808 , \35805 , \35807 );
nand \U$35466 ( \35809 , \35808 , \15181 );
nand \U$35467 ( \35810 , \35804 , \35809 );
xor \U$35468 ( \35811 , \35796 , \35810 );
not \U$35469 ( \35812 , \16541 );
not \U$35470 ( \35813 , RIbb2d9f0_61);
not \U$35471 ( \35814 , \6938 );
or \U$35472 ( \35815 , \35813 , \35814 );
nand \U$35473 ( \35816 , \11534 , \19746 );
nand \U$35474 ( \35817 , \35815 , \35816 );
not \U$35475 ( \35818 , \35817 );
or \U$35476 ( \35819 , \35812 , \35818 );
not \U$35477 ( \35820 , \13879 );
not \U$35478 ( \35821 , \16537 );
and \U$35479 ( \35822 , \35820 , \35821 );
not \U$35480 ( \35823 , \13876 );
and \U$35481 ( \35824 , \35823 , \19746 );
nor \U$35482 ( \35825 , \35822 , \35824 );
not \U$35483 ( \35826 , \35825 );
nand \U$35484 ( \35827 , \35826 , \26834 );
nand \U$35485 ( \35828 , \35819 , \35827 );
and \U$35486 ( \35829 , \35811 , \35828 );
and \U$35487 ( \35830 , \35796 , \35810 );
or \U$35488 ( \35831 , \35829 , \35830 );
and \U$35489 ( \35832 , \35746 , \35831 );
and \U$35490 ( \35833 , \35697 , \35745 );
or \U$35491 ( \35834 , \35832 , \35833 );
not \U$35492 ( \35835 , \35834 );
or \U$35493 ( \35836 , \35645 , \35835 );
not \U$35494 ( \35837 , \35643 );
nand \U$35495 ( \35838 , \35837 , \35518 );
nand \U$35496 ( \35839 , \35836 , \35838 );
not \U$35497 ( \35840 , \35839 );
not \U$35498 ( \35841 , \15181 );
and \U$35499 ( \35842 , RIbb2dcc0_55, \8319 );
not \U$35500 ( \35843 , RIbb2dcc0_55);
and \U$35501 ( \35844 , \35843 , \12214 );
or \U$35502 ( \35845 , \35842 , \35844 );
not \U$35503 ( \35846 , \35845 );
or \U$35504 ( \35847 , \35841 , \35846 );
not \U$35505 ( \35848 , RIbb2dcc0_55);
not \U$35506 ( \35849 , \23529 );
or \U$35507 ( \35850 , \35848 , \35849 );
or \U$35508 ( \35851 , \15786 , RIbb2dcc0_55);
nand \U$35509 ( \35852 , \35850 , \35851 );
nand \U$35510 ( \35853 , \35852 , \14613 );
nand \U$35511 ( \35854 , \35847 , \35853 );
not \U$35512 ( \35855 , \14920 );
not \U$35513 ( \35856 , RIbb2ddb0_53);
not \U$35514 ( \35857 , \12222 );
or \U$35515 ( \35858 , \35856 , \35857 );
nand \U$35516 ( \35859 , \20045 , \16210 );
nand \U$35517 ( \35860 , \35858 , \35859 );
not \U$35518 ( \35861 , \35860 );
or \U$35519 ( \35862 , \35855 , \35861 );
not \U$35520 ( \35863 , RIbb2ddb0_53);
not \U$35521 ( \35864 , \12820 );
or \U$35522 ( \35865 , \35863 , \35864 );
nand \U$35523 ( \35866 , \16475 , \16210 );
nand \U$35524 ( \35867 , \35865 , \35866 );
nand \U$35525 ( \35868 , \35867 , \15688 );
nand \U$35526 ( \35869 , \35862 , \35868 );
and \U$35527 ( \35870 , \35854 , \35869 );
not \U$35528 ( \35871 , \35854 );
and \U$35529 ( \35872 , \35860 , \17563 );
and \U$35530 ( \35873 , \35867 , \14930 );
nor \U$35531 ( \35874 , \35872 , \35873 );
and \U$35532 ( \35875 , \35871 , \35874 );
nor \U$35533 ( \35876 , \35870 , \35875 );
not \U$35534 ( \35877 , RIbb2d888_64);
not \U$35535 ( \35878 , RIbb2d900_63);
not \U$35536 ( \35879 , \13552 );
or \U$35537 ( \35880 , \35878 , \35879 );
nand \U$35538 ( \35881 , \4085 , \20254 );
nand \U$35539 ( \35882 , \35880 , \35881 );
not \U$35540 ( \35883 , \35882 );
or \U$35541 ( \35884 , \35877 , \35883 );
not \U$35542 ( \35885 , RIbb2d900_63);
not \U$35543 ( \35886 , \14536 );
or \U$35544 ( \35887 , \35885 , \35886 );
nand \U$35545 ( \35888 , \6269 , \17262 );
nand \U$35546 ( \35889 , \35887 , \35888 );
nand \U$35547 ( \35890 , \35889 , \17275 );
nand \U$35548 ( \35891 , \35884 , \35890 );
xor \U$35549 ( \35892 , \35876 , \35891 );
not \U$35550 ( \35893 , \6241 );
not \U$35551 ( \35894 , RIbb2e530_37);
not \U$35552 ( \35895 , \27577 );
or \U$35553 ( \35896 , \35894 , \35895 );
nand \U$35554 ( \35897 , \16829 , \4708 );
nand \U$35555 ( \35898 , \35896 , \35897 );
not \U$35556 ( \35899 , \35898 );
or \U$35557 ( \35900 , \35893 , \35899 );
nand \U$35558 ( \35901 , \35665 , \6251 );
nand \U$35559 ( \35902 , \35900 , \35901 );
xor \U$35560 ( \35903 , \35646 , \35651 );
and \U$35561 ( \35904 , \35903 , \35667 );
and \U$35562 ( \35905 , \35646 , \35651 );
or \U$35563 ( \35906 , \35904 , \35905 );
xor \U$35564 ( \35907 , \35902 , \35906 );
not \U$35565 ( \35908 , \10119 );
not \U$35566 ( \35909 , RIbb2e170_45);
not \U$35567 ( \35910 , \14624 );
or \U$35568 ( \35911 , \35909 , \35910 );
nand \U$35569 ( \35912 , \13474 , \13372 );
nand \U$35570 ( \35913 , \35911 , \35912 );
not \U$35571 ( \35914 , \35913 );
or \U$35572 ( \35915 , \35908 , \35914 );
nand \U$35573 ( \35916 , \35694 , \10599 );
nand \U$35574 ( \35917 , \35915 , \35916 );
xor \U$35575 ( \35918 , \35907 , \35917 );
not \U$35576 ( \35919 , \14067 );
not \U$35577 ( \35920 , \35526 );
or \U$35578 ( \35921 , \35919 , \35920 );
and \U$35579 ( \35922 , RIbb2dea0_51, \14563 );
not \U$35580 ( \35923 , RIbb2dea0_51);
and \U$35581 ( \35924 , \35923 , \13525 );
or \U$35582 ( \35925 , \35922 , \35924 );
nand \U$35583 ( \35926 , \35925 , \12692 );
nand \U$35584 ( \35927 , \35921 , \35926 );
xor \U$35585 ( \35928 , \35918 , \35927 );
xor \U$35586 ( \35929 , \35668 , \35678 );
and \U$35587 ( \35930 , \35929 , \35696 );
and \U$35588 ( \35931 , \35668 , \35678 );
or \U$35589 ( \35932 , \35930 , \35931 );
and \U$35590 ( \35933 , \35928 , \35932 );
and \U$35591 ( \35934 , \35918 , \35927 );
or \U$35592 ( \35935 , \35933 , \35934 );
xor \U$35593 ( \35936 , \35892 , \35935 );
xor \U$35594 ( \35937 , \35902 , \35906 );
and \U$35595 ( \35938 , \35937 , \35917 );
and \U$35596 ( \35939 , \35902 , \35906 );
or \U$35597 ( \35940 , \35938 , \35939 );
not \U$35598 ( \35941 , \8353 );
not \U$35599 ( \35942 , RIbb2e350_41);
not \U$35600 ( \35943 , \15031 );
or \U$35601 ( \35944 , \35942 , \35943 );
nand \U$35602 ( \35945 , \17682 , \7097 );
nand \U$35603 ( \35946 , \35944 , \35945 );
not \U$35604 ( \35947 , \35946 );
or \U$35605 ( \35948 , \35941 , \35947 );
nand \U$35606 ( \35949 , \35568 , \8362 );
nand \U$35607 ( \35950 , \35948 , \35949 );
not \U$35608 ( \35951 , \35950 );
not \U$35609 ( \35952 , \11176 );
not \U$35610 ( \35953 , \35674 );
or \U$35611 ( \35954 , \35952 , \35953 );
not \U$35612 ( \35955 , RIbb2e080_47);
not \U$35613 ( \35956 , \16865 );
or \U$35614 ( \35957 , \35955 , \35956 );
nand \U$35615 ( \35958 , \12932 , \10113 );
nand \U$35616 ( \35959 , \35957 , \35958 );
nand \U$35617 ( \35960 , \35959 , \11177 );
nand \U$35618 ( \35961 , \35954 , \35960 );
not \U$35619 ( \35962 , \35961 );
or \U$35620 ( \35963 , \35951 , \35962 );
or \U$35621 ( \35964 , \35961 , \35950 );
not \U$35622 ( \35965 , \9099 );
not \U$35623 ( \35966 , RIbb2e260_43);
not \U$35624 ( \35967 , \13978 );
or \U$35625 ( \35968 , \35966 , \35967 );
nand \U$35626 ( \35969 , \13979 , \17231 );
nand \U$35627 ( \35970 , \35968 , \35969 );
not \U$35628 ( \35971 , \35970 );
or \U$35629 ( \35972 , \35965 , \35971 );
not \U$35630 ( \35973 , RIbb2e260_43);
not \U$35631 ( \35974 , \14528 );
or \U$35632 ( \35975 , \35973 , \35974 );
nand \U$35633 ( \35976 , \15036 , \8347 );
nand \U$35634 ( \35977 , \35975 , \35976 );
nand \U$35635 ( \35978 , \35977 , \9098 );
nand \U$35636 ( \35979 , \35972 , \35978 );
nand \U$35637 ( \35980 , \35964 , \35979 );
nand \U$35638 ( \35981 , \35963 , \35980 );
not \U$35639 ( \35982 , \35981 );
xor \U$35640 ( \35983 , \35940 , \35982 );
not \U$35641 ( \35984 , \13295 );
not \U$35642 ( \35985 , \35493 );
or \U$35643 ( \35986 , \35984 , \35985 );
not \U$35644 ( \35987 , RIbb2df90_49);
not \U$35645 ( \35988 , \12257 );
or \U$35646 ( \35989 , \35987 , \35988 );
nand \U$35647 ( \35990 , \12755 , \12278 );
nand \U$35648 ( \35991 , \35989 , \35990 );
nand \U$35649 ( \35992 , \35991 , \14752 );
nand \U$35650 ( \35993 , \35986 , \35992 );
not \U$35651 ( \35994 , \8354 );
not \U$35652 ( \35995 , \34928 );
or \U$35653 ( \35996 , \35994 , \35995 );
nand \U$35654 ( \35997 , \35946 , \8361 );
nand \U$35655 ( \35998 , \35996 , \35997 );
not \U$35656 ( \35999 , \35998 );
not \U$35657 ( \36000 , \35999 );
not \U$35658 ( \36001 , \11177 );
not \U$35659 ( \36002 , RIbb2e080_47);
not \U$35660 ( \36003 , \19894 );
or \U$35661 ( \36004 , \36002 , \36003 );
nand \U$35662 ( \36005 , \12174 , \12971 );
nand \U$35663 ( \36006 , \36004 , \36005 );
not \U$35664 ( \36007 , \36006 );
or \U$35665 ( \36008 , \36001 , \36007 );
nand \U$35666 ( \36009 , \35959 , \11176 );
nand \U$35667 ( \36010 , \36008 , \36009 );
not \U$35668 ( \36011 , \36010 );
and \U$35669 ( \36012 , \36000 , \36011 );
and \U$35670 ( \36013 , \36010 , \35999 );
nor \U$35671 ( \36014 , \36012 , \36013 );
xor \U$35672 ( \36015 , \35993 , \36014 );
xor \U$35673 ( \36016 , \35983 , \36015 );
xor \U$35674 ( \36017 , \35936 , \36016 );
not \U$35675 ( \36018 , \36017 );
xor \U$35676 ( \36019 , \35487 , \35502 );
and \U$35677 ( \36020 , \36019 , \35517 );
and \U$35678 ( \36021 , \35487 , \35502 );
or \U$35679 ( \36022 , \36020 , \36021 );
and \U$35680 ( \36023 , \35451 , \35460 );
not \U$35681 ( \36024 , \6250 );
not \U$35682 ( \36025 , \35898 );
or \U$35683 ( \36026 , \36024 , \36025 );
not \U$35684 ( \36027 , \6245 );
nand \U$35685 ( \36028 , \36027 , \34830 );
nand \U$35686 ( \36029 , \36026 , \36028 );
xor \U$35687 ( \36030 , \36023 , \36029 );
not \U$35688 ( \36031 , \7104 );
not \U$35689 ( \36032 , \34905 );
or \U$35690 ( \36033 , \36031 , \36032 );
nand \U$35691 ( \36034 , \35484 , \7102 );
nand \U$35692 ( \36035 , \36033 , \36034 );
xor \U$35693 ( \36036 , \36030 , \36035 );
not \U$35694 ( \36037 , \12690 );
not \U$35695 ( \36038 , \35925 );
or \U$35696 ( \36039 , \36037 , \36038 );
not \U$35697 ( \36040 , \25687 );
and \U$35698 ( \36041 , RIbb2dea0_51, \12233 );
not \U$35699 ( \36042 , RIbb2dea0_51);
and \U$35700 ( \36043 , \36042 , \10300 );
or \U$35701 ( \36044 , \36041 , \36043 );
nand \U$35702 ( \36045 , \36040 , \36044 );
nand \U$35703 ( \36046 , \36039 , \36045 );
xor \U$35704 ( \36047 , \36036 , \36046 );
not \U$35705 ( \36048 , \17470 );
and \U$35706 ( \36049 , RIbb2dae0_59, \9010 );
not \U$35707 ( \36050 , RIbb2dae0_59);
and \U$35708 ( \36051 , \36050 , \5955 );
or \U$35709 ( \36052 , \36049 , \36051 );
not \U$35710 ( \36053 , \36052 );
or \U$35711 ( \36054 , \36048 , \36053 );
and \U$35712 ( \36055 , RIbb2dae0_59, \6943 );
not \U$35713 ( \36056 , RIbb2dae0_59);
and \U$35714 ( \36057 , \36056 , \9056 );
or \U$35715 ( \36058 , \36055 , \36057 );
nand \U$35716 ( \36059 , \36058 , \16271 );
nand \U$35717 ( \36060 , \36054 , \36059 );
xnor \U$35718 ( \36061 , \36047 , \36060 );
and \U$35719 ( \36062 , \36022 , \36061 );
not \U$35720 ( \36063 , \36022 );
not \U$35721 ( \36064 , \36061 );
and \U$35722 ( \36065 , \36063 , \36064 );
or \U$35723 ( \36066 , \36062 , \36065 );
xor \U$35724 ( \36067 , \35461 , \35472 );
and \U$35725 ( \36068 , \36067 , \35486 );
and \U$35726 ( \36069 , \35461 , \35472 );
or \U$35727 ( \36070 , \36068 , \36069 );
not \U$35728 ( \36071 , \16674 );
and \U$35729 ( \36072 , RIbb2dbd0_57, \13853 );
not \U$35730 ( \36073 , RIbb2dbd0_57);
and \U$35731 ( \36074 , \36073 , \14673 );
or \U$35732 ( \36075 , \36072 , \36074 );
not \U$35733 ( \36076 , \36075 );
or \U$35734 ( \36077 , \36071 , \36076 );
not \U$35735 ( \36078 , RIbb2dbd0_57);
not \U$35736 ( \36079 , \20772 );
or \U$35737 ( \36080 , \36078 , \36079 );
nand \U$35738 ( \36081 , \25844 , \16671 );
nand \U$35739 ( \36082 , \36080 , \36081 );
nand \U$35740 ( \36083 , \36082 , \15738 );
nand \U$35741 ( \36084 , \36077 , \36083 );
xor \U$35742 ( \36085 , \36070 , \36084 );
not \U$35743 ( \36086 , \18717 );
not \U$35744 ( \36087 , \35507 );
or \U$35745 ( \36088 , \36086 , \36087 );
not \U$35746 ( \36089 , RIbb2d9f0_61);
not \U$35747 ( \36090 , \14000 );
or \U$35748 ( \36091 , \36089 , \36090 );
nand \U$35749 ( \36092 , \6198 , \19746 );
nand \U$35750 ( \36093 , \36091 , \36092 );
nand \U$35751 ( \36094 , \36093 , \16533 );
nand \U$35752 ( \36095 , \36088 , \36094 );
xnor \U$35753 ( \36096 , \36085 , \36095 );
buf \U$35754 ( \36097 , \36096 );
and \U$35755 ( \36098 , \36066 , \36097 );
not \U$35756 ( \36099 , \36066 );
not \U$35757 ( \36100 , \36097 );
and \U$35758 ( \36101 , \36099 , \36100 );
nor \U$35759 ( \36102 , \36098 , \36101 );
not \U$35760 ( \36103 , \36102 );
and \U$35761 ( \36104 , \36018 , \36103 );
and \U$35762 ( \36105 , \36017 , \36102 );
nor \U$35763 ( \36106 , \36104 , \36105 );
not \U$35764 ( \36107 , \36106 );
or \U$35765 ( \36108 , \35840 , \36107 );
or \U$35766 ( \36109 , \36106 , \35839 );
nand \U$35767 ( \36110 , \36108 , \36109 );
xor \U$35768 ( \36111 , \35587 , \35620 );
xor \U$35769 ( \36112 , \36111 , \35637 );
xor \U$35770 ( \36113 , \35588 , \35605 );
xor \U$35771 ( \36114 , \36113 , \35617 );
not \U$35772 ( \36115 , \11176 );
not \U$35773 ( \36116 , RIbb2e080_47);
not \U$35774 ( \36117 , \14503 );
or \U$35775 ( \36118 , \36116 , \36117 );
nand \U$35776 ( \36119 , \35685 , \16171 );
nand \U$35777 ( \36120 , \36118 , \36119 );
not \U$35778 ( \36121 , \36120 );
or \U$35779 ( \36122 , \36115 , \36121 );
nand \U$35780 ( \36123 , \35627 , \12965 );
nand \U$35781 ( \36124 , \36122 , \36123 );
xor \U$35782 ( \36125 , \36114 , \36124 );
not \U$35783 ( \36126 , \12692 );
not \U$35784 ( \36127 , \35704 );
or \U$35785 ( \36128 , \36126 , \36127 );
and \U$35786 ( \36129 , RIbb2dea0_51, \15484 );
not \U$35787 ( \36130 , RIbb2dea0_51);
and \U$35788 ( \36131 , \36130 , \12933 );
or \U$35789 ( \36132 , \36129 , \36131 );
nand \U$35790 ( \36133 , \36132 , \14067 );
nand \U$35791 ( \36134 , \36128 , \36133 );
and \U$35792 ( \36135 , \36125 , \36134 );
and \U$35793 ( \36136 , \36114 , \36124 );
or \U$35794 ( \36137 , \36135 , \36136 );
xor \U$35795 ( \36138 , \36112 , \36137 );
not \U$35796 ( \36139 , \26834 );
not \U$35797 ( \36140 , \35817 );
or \U$35798 ( \36141 , \36139 , \36140 );
not \U$35799 ( \36142 , RIbb2d9f0_61);
not \U$35800 ( \36143 , \9071 );
or \U$35801 ( \36144 , \36142 , \36143 );
nand \U$35802 ( \36145 , \9074 , \16254 );
nand \U$35803 ( \36146 , \36144 , \36145 );
nand \U$35804 ( \36147 , \36146 , \18717 );
nand \U$35805 ( \36148 , \36141 , \36147 );
not \U$35806 ( \36149 , \36148 );
not \U$35807 ( \36150 , \14613 );
and \U$35808 ( \36151 , RIbb2dcc0_55, \14563 );
not \U$35809 ( \36152 , RIbb2dcc0_55);
and \U$35810 ( \36153 , \36152 , \10764 );
or \U$35811 ( \36154 , \36151 , \36153 );
not \U$35812 ( \36155 , \36154 );
or \U$35813 ( \36156 , \36150 , \36155 );
nand \U$35814 ( \36157 , \35802 , \15182 );
nand \U$35815 ( \36158 , \36156 , \36157 );
not \U$35816 ( \36159 , \36158 );
or \U$35817 ( \36160 , \36149 , \36159 );
or \U$35818 ( \36161 , \36158 , \36148 );
xor \U$35819 ( \36162 , \35751 , \35759 );
not \U$35820 ( \36163 , \7104 );
not \U$35821 ( \36164 , \35613 );
or \U$35822 ( \36165 , \36163 , \36164 );
and \U$35823 ( \36166 , RIbb2e440_39, \26050 );
not \U$35824 ( \36167 , RIbb2e440_39);
and \U$35825 ( \36168 , \36167 , \17529 );
or \U$35826 ( \36169 , \36166 , \36168 );
nand \U$35827 ( \36170 , \36169 , \7102 );
nand \U$35828 ( \36171 , \36165 , \36170 );
xor \U$35829 ( \36172 , \36162 , \36171 );
not \U$35830 ( \36173 , \8362 );
not \U$35831 ( \36174 , RIbb2e350_41);
not \U$35832 ( \36175 , \34293 );
or \U$35833 ( \36176 , \36174 , \36175 );
nand \U$35834 ( \36177 , \16556 , \9402 );
nand \U$35835 ( \36178 , \36176 , \36177 );
not \U$35836 ( \36179 , \36178 );
or \U$35837 ( \36180 , \36173 , \36179 );
nand \U$35838 ( \36181 , \35767 , \8354 );
nand \U$35839 ( \36182 , \36180 , \36181 );
and \U$35840 ( \36183 , \36172 , \36182 );
and \U$35841 ( \36184 , \36162 , \36171 );
or \U$35842 ( \36185 , \36183 , \36184 );
nand \U$35843 ( \36186 , \36161 , \36185 );
nand \U$35844 ( \36187 , \36160 , \36186 );
and \U$35845 ( \36188 , \36138 , \36187 );
and \U$35846 ( \36189 , \36112 , \36137 );
or \U$35847 ( \36190 , \36188 , \36189 );
not \U$35848 ( \36191 , RIbb2e260_43);
not \U$35849 ( \36192 , \17681 );
or \U$35850 ( \36193 , \36191 , \36192 );
nand \U$35851 ( \36194 , \15474 , \26255 );
nand \U$35852 ( \36195 , \36193 , \36194 );
not \U$35853 ( \36196 , \36195 );
not \U$35854 ( \36197 , \9099 );
or \U$35855 ( \36198 , \36196 , \36197 );
nand \U$35856 ( \36199 , \35784 , \9098 );
nand \U$35857 ( \36200 , \36198 , \36199 );
not \U$35858 ( \36201 , \13295 );
not \U$35859 ( \36202 , RIbb2df90_49);
not \U$35860 ( \36203 , \33497 );
or \U$35861 ( \36204 , \36202 , \36203 );
nand \U$35862 ( \36205 , \12349 , \12278 );
nand \U$35863 ( \36206 , \36204 , \36205 );
not \U$35864 ( \36207 , \36206 );
or \U$35865 ( \36208 , \36201 , \36207 );
not \U$35866 ( \36209 , RIbb2df90_49);
not \U$35867 ( \36210 , \12934 );
or \U$35868 ( \36211 , \36209 , \36210 );
nand \U$35869 ( \36212 , \12324 , \12278 );
nand \U$35870 ( \36213 , \36211 , \36212 );
nand \U$35871 ( \36214 , \36213 , \14752 );
nand \U$35872 ( \36215 , \36208 , \36214 );
xor \U$35873 ( \36216 , \36200 , \36215 );
not \U$35874 ( \36217 , \10119 );
not \U$35875 ( \36218 , \35687 );
or \U$35876 ( \36219 , \36217 , \36218 );
not \U$35877 ( \36220 , RIbb2e170_45);
not \U$35878 ( \36221 , \21770 );
or \U$35879 ( \36222 , \36220 , \36221 );
nand \U$35880 ( \36223 , \14527 , \11065 );
nand \U$35881 ( \36224 , \36222 , \36223 );
nand \U$35882 ( \36225 , \36224 , \10117 );
nand \U$35883 ( \36226 , \36219 , \36225 );
xor \U$35884 ( \36227 , \36216 , \36226 );
not \U$35885 ( \36228 , \10117 );
not \U$35886 ( \36229 , RIbb2e170_45);
not \U$35887 ( \36230 , \15031 );
or \U$35888 ( \36231 , \36229 , \36230 );
nand \U$35889 ( \36232 , \15474 , \9094 );
nand \U$35890 ( \36233 , \36231 , \36232 );
not \U$35891 ( \36234 , \36233 );
or \U$35892 ( \36235 , \36228 , \36234 );
nand \U$35893 ( \36236 , \36224 , \10119 );
nand \U$35894 ( \36237 , \36235 , \36236 );
not \U$35895 ( \36238 , \12169 );
not \U$35896 ( \36239 , \36206 );
or \U$35897 ( \36240 , \36238 , \36239 );
not \U$35898 ( \36241 , RIbb2df90_49);
not \U$35899 ( \36242 , \13211 );
or \U$35900 ( \36243 , \36241 , \36242 );
nand \U$35901 ( \36244 , \35633 , \12278 );
nand \U$35902 ( \36245 , \36243 , \36244 );
nand \U$35903 ( \36246 , \36245 , \12167 );
nand \U$35904 ( \36247 , \36240 , \36246 );
xor \U$35905 ( \36248 , \36237 , \36247 );
not \U$35906 ( \36249 , \17397 );
not \U$35907 ( \36250 , RIbb2dbd0_57);
not \U$35908 ( \36251 , \12820 );
or \U$35909 ( \36252 , \36250 , \36251 );
nand \U$35910 ( \36253 , \9280 , \15741 );
nand \U$35911 ( \36254 , \36252 , \36253 );
not \U$35912 ( \36255 , \36254 );
or \U$35913 ( \36256 , \36249 , \36255 );
not \U$35914 ( \36257 , RIbb2dbd0_57);
not \U$35915 ( \36258 , \22580 );
or \U$35916 ( \36259 , \36257 , \36258 );
nand \U$35917 ( \36260 , \9841 , \15741 );
nand \U$35918 ( \36261 , \36259 , \36260 );
nand \U$35919 ( \36262 , \36261 , \16675 );
nand \U$35920 ( \36263 , \36256 , \36262 );
and \U$35921 ( \36264 , \36248 , \36263 );
and \U$35922 ( \36265 , \36237 , \36247 );
or \U$35923 ( \36266 , \36264 , \36265 );
xor \U$35924 ( \36267 , \36227 , \36266 );
not \U$35925 ( \36268 , \16271 );
and \U$35926 ( \36269 , RIbb2dae0_59, \12194 );
not \U$35927 ( \36270 , RIbb2dae0_59);
and \U$35928 ( \36271 , \36270 , \8631 );
or \U$35929 ( \36272 , \36269 , \36271 );
not \U$35930 ( \36273 , \36272 );
or \U$35931 ( \36274 , \36268 , \36273 );
not \U$35932 ( \36275 , \35711 );
nand \U$35933 ( \36276 , \36275 , \17470 );
nand \U$35934 ( \36277 , \36274 , \36276 );
not \U$35935 ( \36278 , RIbb2d888_64);
not \U$35936 ( \36279 , RIbb2d900_63);
not \U$35937 ( \36280 , \5956 );
or \U$35938 ( \36281 , \36279 , \36280 );
nand \U$35939 ( \36282 , \5955 , \17262 );
nand \U$35940 ( \36283 , \36281 , \36282 );
not \U$35941 ( \36284 , \36283 );
or \U$35942 ( \36285 , \36278 , \36284 );
not \U$35943 ( \36286 , RIbb2d900_63);
not \U$35944 ( \36287 , \8338 );
or \U$35945 ( \36288 , \36286 , \36287 );
nand \U$35946 ( \36289 , \10156 , \20254 );
nand \U$35947 ( \36290 , \36288 , \36289 );
nand \U$35948 ( \36291 , \36290 , \17275 );
nand \U$35949 ( \36292 , \36285 , \36291 );
nor \U$35950 ( \36293 , \36277 , \36292 );
not \U$35951 ( \36294 , \17563 );
not \U$35952 ( \36295 , RIbb2ddb0_53);
not \U$35953 ( \36296 , \22555 );
not \U$35954 ( \36297 , \36296 );
or \U$35955 ( \36298 , \36295 , \36297 );
nand \U$35956 ( \36299 , \11581 , \13463 );
nand \U$35957 ( \36300 , \36298 , \36299 );
not \U$35958 ( \36301 , \36300 );
or \U$35959 ( \36302 , \36294 , \36301 );
nand \U$35960 ( \36303 , \35734 , \14930 );
nand \U$35961 ( \36304 , \36302 , \36303 );
not \U$35962 ( \36305 , \36304 );
or \U$35963 ( \36306 , \36293 , \36305 );
nand \U$35964 ( \36307 , \36277 , \36292 );
nand \U$35965 ( \36308 , \36306 , \36307 );
and \U$35966 ( \36309 , \36267 , \36308 );
and \U$35967 ( \36310 , \36227 , \36266 );
or \U$35968 ( \36311 , \36309 , \36310 );
xor \U$35969 ( \36312 , \36190 , \36311 );
xor \U$35970 ( \36313 , \35697 , \35745 );
xor \U$35971 ( \36314 , \36313 , \35831 );
and \U$35972 ( \36315 , \36312 , \36314 );
and \U$35973 ( \36316 , \36190 , \36311 );
or \U$35974 ( \36317 , \36315 , \36316 );
not \U$35975 ( \36318 , \36317 );
xor \U$35976 ( \36319 , \35918 , \35927 );
xor \U$35977 ( \36320 , \36319 , \35932 );
xor \U$35978 ( \36321 , \36200 , \36215 );
and \U$35979 ( \36322 , \36321 , \36226 );
and \U$35980 ( \36323 , \36200 , \36215 );
or \U$35981 ( \36324 , \36322 , \36323 );
not \U$35982 ( \36325 , \16675 );
not \U$35983 ( \36326 , \36254 );
or \U$35984 ( \36327 , \36325 , \36326 );
not \U$35985 ( \36328 , RIbb2dbd0_57);
not \U$35986 ( \36329 , \12194 );
or \U$35987 ( \36330 , \36328 , \36329 );
nand \U$35988 ( \36331 , \13866 , \14602 );
nand \U$35989 ( \36332 , \36330 , \36331 );
nand \U$35990 ( \36333 , \36332 , \17397 );
nand \U$35991 ( \36334 , \36327 , \36333 );
not \U$35992 ( \36335 , \17275 );
not \U$35993 ( \36336 , \36283 );
or \U$35994 ( \36337 , \36335 , \36336 );
not \U$35995 ( \36338 , \8387 );
not \U$35996 ( \36339 , \19721 );
and \U$35997 ( \36340 , \36338 , \36339 );
and \U$35998 ( \36341 , \7111 , \19721 );
nor \U$35999 ( \36342 , \36340 , \36341 );
not \U$36000 ( \36343 , \36342 );
nand \U$36001 ( \36344 , \36343 , RIbb2d888_64);
nand \U$36002 ( \36345 , \36337 , \36344 );
nor \U$36003 ( \36346 , \36334 , \36345 );
xor \U$36004 ( \36347 , \35538 , \35551 );
not \U$36005 ( \36348 , \6241 );
not \U$36006 ( \36349 , \35658 );
or \U$36007 ( \36350 , \36348 , \36349 );
nand \U$36008 ( \36351 , \35594 , \6250 );
nand \U$36009 ( \36352 , \36350 , \36351 );
xor \U$36010 ( \36353 , \36347 , \36352 );
or \U$36011 ( \36354 , \35774 , \8363 );
or \U$36012 ( \36355 , \35575 , \8352 );
nand \U$36013 ( \36356 , \36354 , \36355 );
xor \U$36014 ( \36357 , \36353 , \36356 );
not \U$36015 ( \36358 , \36357 );
or \U$36016 ( \36359 , \36346 , \36358 );
nand \U$36017 ( \36360 , \36334 , \36345 );
nand \U$36018 ( \36361 , \36359 , \36360 );
xor \U$36019 ( \36362 , \36324 , \36361 );
not \U$36020 ( \36363 , \9099 );
not \U$36021 ( \36364 , \35977 );
or \U$36022 ( \36365 , \36363 , \36364 );
nand \U$36023 ( \36366 , \36195 , \9098 );
nand \U$36024 ( \36367 , \36365 , \36366 );
not \U$36025 ( \36368 , \14752 );
not \U$36026 ( \36369 , \35500 );
or \U$36027 ( \36370 , \36368 , \36369 );
nand \U$36028 ( \36371 , \36213 , \13295 );
nand \U$36029 ( \36372 , \36370 , \36371 );
xor \U$36030 ( \36373 , \36367 , \36372 );
not \U$36031 ( \36374 , \16675 );
not \U$36032 ( \36375 , \36332 );
or \U$36033 ( \36376 , \36374 , \36375 );
not \U$36034 ( \36377 , RIbb2dbd0_57);
not \U$36035 ( \36378 , \12211 );
or \U$36036 ( \36379 , \36377 , \36378 );
nand \U$36037 ( \36380 , \34501 , \14602 );
nand \U$36038 ( \36381 , \36379 , \36380 );
nand \U$36039 ( \36382 , \36381 , \15738 );
nand \U$36040 ( \36383 , \36376 , \36382 );
xor \U$36041 ( \36384 , \36373 , \36383 );
and \U$36042 ( \36385 , \36362 , \36384 );
and \U$36043 ( \36386 , \36324 , \36361 );
or \U$36044 ( \36387 , \36385 , \36386 );
xor \U$36045 ( \36388 , \36320 , \36387 );
xor \U$36046 ( \36389 , \36367 , \36372 );
and \U$36047 ( \36390 , \36389 , \36383 );
and \U$36048 ( \36391 , \36367 , \36372 );
or \U$36049 ( \36392 , \36390 , \36391 );
xor \U$36050 ( \36393 , \36347 , \36352 );
and \U$36051 ( \36394 , \36393 , \36356 );
and \U$36052 ( \36395 , \36347 , \36352 );
or \U$36053 ( \36396 , \36394 , \36395 );
not \U$36054 ( \36397 , RIbb2d888_64);
and \U$36055 ( \36398 , \6198 , \20254 );
not \U$36056 ( \36399 , \6198 );
and \U$36057 ( \36400 , \36399 , RIbb2d900_63);
or \U$36058 ( \36401 , \36398 , \36400 );
not \U$36059 ( \36402 , \36401 );
or \U$36060 ( \36403 , \36397 , \36402 );
not \U$36061 ( \36404 , \17275 );
or \U$36062 ( \36405 , \36342 , \36404 );
nand \U$36063 ( \36406 , \36403 , \36405 );
xor \U$36064 ( \36407 , \36396 , \36406 );
or \U$36065 ( \36408 , \35825 , \16542 );
or \U$36066 ( \36409 , \35515 , \16534 );
nand \U$36067 ( \36410 , \36408 , \36409 );
and \U$36068 ( \36411 , \36407 , \36410 );
and \U$36069 ( \36412 , \36396 , \36406 );
or \U$36070 ( \36413 , \36411 , \36412 );
xor \U$36071 ( \36414 , \36392 , \36413 );
not \U$36072 ( \36415 , \14613 );
not \U$36073 ( \36416 , \35808 );
or \U$36074 ( \36417 , \36415 , \36416 );
and \U$36075 ( \36418 , RIbb2dcc0_55, \13916 );
not \U$36076 ( \36419 , RIbb2dcc0_55);
and \U$36077 ( \36420 , \36419 , \16475 );
or \U$36078 ( \36421 , \36418 , \36420 );
nand \U$36079 ( \36422 , \36421 , \15181 );
nand \U$36080 ( \36423 , \36417 , \36422 );
not \U$36081 ( \36424 , \36423 );
not \U$36082 ( \36425 , \36424 );
not \U$36083 ( \36426 , \16271 );
not \U$36084 ( \36427 , \35719 );
or \U$36085 ( \36428 , \36426 , \36427 );
not \U$36086 ( \36429 , RIbb2dae0_59);
not \U$36087 ( \36430 , \9791 );
or \U$36088 ( \36431 , \36429 , \36430 );
not \U$36089 ( \36432 , \8639 );
nand \U$36090 ( \36433 , \36432 , \25675 );
nand \U$36091 ( \36434 , \36431 , \36433 );
nand \U$36092 ( \36435 , \36434 , \17470 );
nand \U$36093 ( \36436 , \36428 , \36435 );
not \U$36094 ( \36437 , \36436 );
not \U$36095 ( \36438 , \36437 );
or \U$36096 ( \36439 , \36425 , \36438 );
not \U$36097 ( \36440 , \13467 );
not \U$36098 ( \36441 , \35741 );
or \U$36099 ( \36442 , \36440 , \36441 );
and \U$36100 ( \36443 , \12234 , RIbb2ddb0_53);
not \U$36101 ( \36444 , \12234 );
and \U$36102 ( \36445 , \36444 , \16210 );
or \U$36103 ( \36446 , \36443 , \36445 );
nand \U$36104 ( \36447 , \36446 , \14930 );
nand \U$36105 ( \36448 , \36442 , \36447 );
nand \U$36106 ( \36449 , \36439 , \36448 );
nand \U$36107 ( \36450 , \36436 , \36423 );
nand \U$36108 ( \36451 , \36449 , \36450 );
xor \U$36109 ( \36452 , \36414 , \36451 );
xor \U$36110 ( \36453 , \36388 , \36452 );
not \U$36111 ( \36454 , \36453 );
or \U$36112 ( \36455 , \36318 , \36454 );
or \U$36113 ( \36456 , \36453 , \36317 );
xor \U$36114 ( \36457 , \36324 , \36361 );
xor \U$36115 ( \36458 , \36457 , \36384 );
xor \U$36116 ( \36459 , \35796 , \35810 );
xor \U$36117 ( \36460 , \36459 , \35828 );
and \U$36118 ( \36461 , \36334 , \36358 );
not \U$36119 ( \36462 , \36334 );
and \U$36120 ( \36463 , \36462 , \36357 );
nor \U$36121 ( \36464 , \36461 , \36463 );
xnor \U$36122 ( \36465 , \36464 , \36345 );
xor \U$36123 ( \36466 , \36460 , \36465 );
and \U$36124 ( \36467 , \35743 , \35726 );
not \U$36125 ( \36468 , \35743 );
and \U$36126 ( \36469 , \36468 , \35706 );
or \U$36127 ( \36470 , \36467 , \36469 );
xor \U$36128 ( \36471 , \36470 , \35722 );
and \U$36129 ( \36472 , \36466 , \36471 );
and \U$36130 ( \36473 , \36460 , \36465 );
or \U$36131 ( \36474 , \36472 , \36473 );
xor \U$36132 ( \36475 , \36458 , \36474 );
xor \U$36133 ( \36476 , \35579 , \35640 );
xnor \U$36134 ( \36477 , \36476 , \35533 );
xor \U$36135 ( \36478 , \36396 , \36406 );
xor \U$36136 ( \36479 , \36478 , \36410 );
not \U$36137 ( \36480 , \36479 );
and \U$36138 ( \36481 , \36437 , \36424 );
not \U$36139 ( \36482 , \36437 );
and \U$36140 ( \36483 , \36482 , \36423 );
nor \U$36141 ( \36484 , \36481 , \36483 );
and \U$36142 ( \36485 , \36484 , \36448 );
not \U$36143 ( \36486 , \36484 );
not \U$36144 ( \36487 , \36448 );
and \U$36145 ( \36488 , \36486 , \36487 );
nor \U$36146 ( \36489 , \36485 , \36488 );
not \U$36147 ( \36490 , \36489 );
xor \U$36148 ( \36491 , \36480 , \36490 );
xor \U$36149 ( \36492 , \36477 , \36491 );
and \U$36150 ( \36493 , \36475 , \36492 );
and \U$36151 ( \36494 , \36458 , \36474 );
or \U$36152 ( \36495 , \36493 , \36494 );
nand \U$36153 ( \36496 , \36456 , \36495 );
nand \U$36154 ( \36497 , \36455 , \36496 );
xor \U$36155 ( \36498 , \36110 , \36497 );
xor \U$36156 ( \36499 , \36320 , \36387 );
and \U$36157 ( \36500 , \36499 , \36452 );
and \U$36158 ( \36501 , \36320 , \36387 );
or \U$36159 ( \36502 , \36500 , \36501 );
not \U$36160 ( \36503 , \36502 );
not \U$36161 ( \36504 , \36503 );
xor \U$36162 ( \36505 , \34954 , \34964 );
xor \U$36163 ( \36506 , \36505 , \34975 );
not \U$36164 ( \36507 , \10117 );
not \U$36165 ( \36508 , \35913 );
or \U$36166 ( \36509 , \36507 , \36508 );
nand \U$36167 ( \36510 , \34912 , \10119 );
nand \U$36168 ( \36511 , \36509 , \36510 );
xor \U$36169 ( \36512 , \36506 , \36511 );
not \U$36170 ( \36513 , \9098 );
not \U$36171 ( \36514 , \35970 );
or \U$36172 ( \36515 , \36513 , \36514 );
nand \U$36173 ( \36516 , \34985 , \9099 );
nand \U$36174 ( \36517 , \36515 , \36516 );
xor \U$36175 ( \36518 , \36512 , \36517 );
not \U$36176 ( \36519 , \14613 );
not \U$36177 ( \36520 , \36421 );
or \U$36178 ( \36521 , \36519 , \36520 );
nand \U$36179 ( \36522 , \35852 , \15181 );
nand \U$36180 ( \36523 , \36521 , \36522 );
not \U$36181 ( \36524 , \36523 );
not \U$36182 ( \36525 , \16674 );
not \U$36183 ( \36526 , \36381 );
or \U$36184 ( \36527 , \36525 , \36526 );
nand \U$36185 ( \36528 , \36075 , \15738 );
nand \U$36186 ( \36529 , \36527 , \36528 );
not \U$36187 ( \36530 , \36529 );
or \U$36188 ( \36531 , \36524 , \36530 );
or \U$36189 ( \36532 , \36529 , \36523 );
xor \U$36190 ( \36533 , \35552 , \35561 );
and \U$36191 ( \36534 , \36533 , \35578 );
and \U$36192 ( \36535 , \35552 , \35561 );
or \U$36193 ( \36536 , \36534 , \36535 );
nand \U$36194 ( \36537 , \36532 , \36536 );
nand \U$36195 ( \36538 , \36531 , \36537 );
xor \U$36196 ( \36539 , \36518 , \36538 );
not \U$36197 ( \36540 , \17275 );
not \U$36198 ( \36541 , \36401 );
or \U$36199 ( \36542 , \36540 , \36541 );
nand \U$36200 ( \36543 , \35889 , RIbb2d888_64);
nand \U$36201 ( \36544 , \36542 , \36543 );
not \U$36202 ( \36545 , \36544 );
not \U$36203 ( \36546 , \16271 );
not \U$36204 ( \36547 , \36434 );
or \U$36205 ( \36548 , \36546 , \36547 );
nand \U$36206 ( \36549 , \36058 , \17470 );
nand \U$36207 ( \36550 , \36548 , \36549 );
not \U$36208 ( \36551 , \36550 );
or \U$36209 ( \36552 , \36545 , \36551 );
or \U$36210 ( \36553 , \36550 , \36544 );
not \U$36211 ( \36554 , \13467 );
not \U$36212 ( \36555 , \36446 );
or \U$36213 ( \36556 , \36554 , \36555 );
nand \U$36214 ( \36557 , \35860 , \14930 );
nand \U$36215 ( \36558 , \36556 , \36557 );
nand \U$36216 ( \36559 , \36553 , \36558 );
nand \U$36217 ( \36560 , \36552 , \36559 );
xnor \U$36218 ( \36561 , \36539 , \36560 );
xor \U$36219 ( \36562 , \36392 , \36413 );
and \U$36220 ( \36563 , \36562 , \36451 );
and \U$36221 ( \36564 , \36392 , \36413 );
or \U$36222 ( \36565 , \36563 , \36564 );
xor \U$36223 ( \36566 , \36561 , \36565 );
xor \U$36224 ( \36567 , \35979 , \35950 );
xor \U$36225 ( \36568 , \36567 , \35961 );
xor \U$36226 ( \36569 , \36529 , \36523 );
xor \U$36227 ( \36570 , \36536 , \36569 );
xor \U$36228 ( \36571 , \36568 , \36570 );
xor \U$36229 ( \36572 , \36558 , \36550 );
xor \U$36230 ( \36573 , \36544 , \36572 );
and \U$36231 ( \36574 , \36571 , \36573 );
and \U$36232 ( \36575 , \36568 , \36570 );
or \U$36233 ( \36576 , \36574 , \36575 );
xor \U$36234 ( \36577 , \36566 , \36576 );
not \U$36235 ( \36578 , \36577 );
not \U$36236 ( \36579 , \36578 );
or \U$36237 ( \36580 , \36504 , \36579 );
nand \U$36238 ( \36581 , \36577 , \36502 );
nand \U$36239 ( \36582 , \36580 , \36581 );
xor \U$36240 ( \36583 , \36568 , \36570 );
xor \U$36241 ( \36584 , \36583 , \36573 );
not \U$36242 ( \36585 , \36584 );
not \U$36243 ( \36586 , \36479 );
not \U$36244 ( \36587 , \36489 );
or \U$36245 ( \36588 , \36586 , \36587 );
not \U$36246 ( \36589 , \36489 );
and \U$36247 ( \36590 , \36480 , \36589 );
not \U$36248 ( \36591 , \36590 );
nand \U$36249 ( \36592 , \36591 , \36477 );
nand \U$36250 ( \36593 , \36588 , \36592 );
not \U$36251 ( \36594 , \36593 );
or \U$36252 ( \36595 , \36585 , \36594 );
or \U$36253 ( \36596 , \36593 , \36584 );
not \U$36254 ( \36597 , \35643 );
not \U$36255 ( \36598 , \35518 );
and \U$36256 ( \36599 , \36597 , \36598 );
and \U$36257 ( \36600 , \35518 , \35643 );
nor \U$36258 ( \36601 , \36599 , \36600 );
not \U$36259 ( \36602 , \36601 );
not \U$36260 ( \36603 , \35834 );
or \U$36261 ( \36604 , \36602 , \36603 );
or \U$36262 ( \36605 , \35834 , \36601 );
nand \U$36263 ( \36606 , \36604 , \36605 );
nand \U$36264 ( \36607 , \36596 , \36606 );
nand \U$36265 ( \36608 , \36595 , \36607 );
and \U$36266 ( \36609 , \36582 , \36608 );
not \U$36267 ( \36610 , \36582 );
not \U$36268 ( \36611 , \36608 );
and \U$36269 ( \36612 , \36610 , \36611 );
nor \U$36270 ( \36613 , \36609 , \36612 );
xor \U$36271 ( \36614 , \36498 , \36613 );
not \U$36272 ( \36615 , \36614 );
xor \U$36273 ( \36616 , \36317 , \36453 );
xor \U$36274 ( \36617 , \36616 , \36495 );
not \U$36275 ( \36618 , \36617 );
xor \U$36276 ( \36619 , \36227 , \36266 );
xor \U$36277 ( \36620 , \36619 , \36308 );
xor \U$36278 ( \36621 , \36277 , \36305 );
xnor \U$36279 ( \36622 , \36621 , \36292 );
xor \U$36280 ( \36623 , \36114 , \36124 );
xor \U$36281 ( \36624 , \36623 , \36134 );
or \U$36282 ( \36625 , \36622 , \36624 );
xor \U$36283 ( \36626 , \36158 , \36148 );
xor \U$36284 ( \36627 , \36626 , \36185 );
nand \U$36285 ( \36628 , \36625 , \36627 );
nand \U$36286 ( \36629 , \36622 , \36624 );
nand \U$36287 ( \36630 , \36628 , \36629 );
xor \U$36288 ( \36631 , \36620 , \36630 );
xor \U$36289 ( \36632 , \36460 , \36465 );
xor \U$36290 ( \36633 , \36632 , \36471 );
and \U$36291 ( \36634 , \36631 , \36633 );
and \U$36292 ( \36635 , \36620 , \36630 );
or \U$36293 ( \36636 , \36634 , \36635 );
xor \U$36294 ( \36637 , \36190 , \36311 );
xor \U$36295 ( \36638 , \36637 , \36314 );
not \U$36296 ( \36639 , \36638 );
xor \U$36297 ( \36640 , \35760 , \35777 );
xor \U$36298 ( \36641 , \36640 , \35793 );
and \U$36299 ( \36642 , \19064 , \6240 );
not \U$36300 ( \36643 , \7104 );
not \U$36301 ( \36644 , \36169 );
or \U$36302 ( \36645 , \36643 , \36644 );
and \U$36303 ( \36646 , RIbb2e440_39, \35597 );
not \U$36304 ( \36647 , RIbb2e440_39);
and \U$36305 ( \36648 , \36647 , \28621 );
or \U$36306 ( \36649 , \36646 , \36648 );
nand \U$36307 ( \36650 , \36649 , \7102 );
nand \U$36308 ( \36651 , \36645 , \36650 );
xor \U$36309 ( \36652 , \36642 , \36651 );
not \U$36310 ( \36653 , \8353 );
not \U$36311 ( \36654 , \36178 );
or \U$36312 ( \36655 , \36653 , \36654 );
not \U$36313 ( \36656 , RIbb2e350_41);
not \U$36314 ( \36657 , \27234 );
or \U$36315 ( \36658 , \36656 , \36657 );
nand \U$36316 ( \36659 , \16704 , \9402 );
nand \U$36317 ( \36660 , \36658 , \36659 );
nand \U$36318 ( \36661 , \36660 , \8361 );
nand \U$36319 ( \36662 , \36655 , \36661 );
and \U$36320 ( \36663 , \36652 , \36662 );
and \U$36321 ( \36664 , \36642 , \36651 );
or \U$36322 ( \36665 , \36663 , \36664 );
not \U$36323 ( \36666 , \9098 );
and \U$36324 ( \36667 , \16747 , RIbb2e260_43);
not \U$36325 ( \36668 , \16747 );
and \U$36326 ( \36669 , \36668 , \8347 );
or \U$36327 ( \36670 , \36667 , \36669 );
not \U$36328 ( \36671 , \36670 );
or \U$36329 ( \36672 , \36666 , \36671 );
nand \U$36330 ( \36673 , \35791 , \10451 );
nand \U$36331 ( \36674 , \36672 , \36673 );
xor \U$36332 ( \36675 , \36665 , \36674 );
not \U$36333 ( \36676 , \12774 );
not \U$36334 ( \36677 , \33497 );
xor \U$36335 ( \36678 , RIbb2dea0_51, \36677 );
not \U$36336 ( \36679 , \36678 );
or \U$36337 ( \36680 , \36676 , \36679 );
nand \U$36338 ( \36681 , \36132 , \12692 );
nand \U$36339 ( \36682 , \36680 , \36681 );
and \U$36340 ( \36683 , \36675 , \36682 );
and \U$36341 ( \36684 , \36665 , \36674 );
or \U$36342 ( \36685 , \36683 , \36684 );
xor \U$36343 ( \36686 , \36641 , \36685 );
not \U$36344 ( \36687 , \10119 );
not \U$36345 ( \36688 , \36233 );
or \U$36346 ( \36689 , \36687 , \36688 );
not \U$36347 ( \36690 , RIbb2e170_45);
not \U$36348 ( \36691 , \21665 );
or \U$36349 ( \36692 , \36690 , \36691 );
nand \U$36350 ( \36693 , \15753 , \9094 );
nand \U$36351 ( \36694 , \36692 , \36693 );
nand \U$36352 ( \36695 , \36694 , \10117 );
nand \U$36353 ( \36696 , \36689 , \36695 );
not \U$36354 ( \36697 , \11176 );
not \U$36355 ( \36698 , RIbb2e080_47);
not \U$36356 ( \36699 , \21770 );
or \U$36357 ( \36700 , \36698 , \36699 );
nand \U$36358 ( \36701 , \14527 , \15632 );
nand \U$36359 ( \36702 , \36700 , \36701 );
not \U$36360 ( \36703 , \36702 );
or \U$36361 ( \36704 , \36697 , \36703 );
nand \U$36362 ( \36705 , \36120 , \12965 );
nand \U$36363 ( \36706 , \36704 , \36705 );
xor \U$36364 ( \36707 , \36696 , \36706 );
not \U$36365 ( \36708 , \12167 );
not \U$36366 ( \36709 , RIbb2df90_49);
not \U$36367 ( \36710 , \15054 );
or \U$36368 ( \36711 , \36709 , \36710 );
nand \U$36369 ( \36712 , \13547 , \12278 );
nand \U$36370 ( \36713 , \36711 , \36712 );
not \U$36371 ( \36714 , \36713 );
or \U$36372 ( \36715 , \36708 , \36714 );
nand \U$36373 ( \36716 , \36245 , \14752 );
nand \U$36374 ( \36717 , \36715 , \36716 );
and \U$36375 ( \36718 , \36707 , \36717 );
and \U$36376 ( \36719 , \36696 , \36706 );
or \U$36377 ( \36720 , \36718 , \36719 );
and \U$36378 ( \36721 , \36686 , \36720 );
and \U$36379 ( \36722 , \36641 , \36685 );
or \U$36380 ( \36723 , \36721 , \36722 );
xor \U$36381 ( \36724 , \36112 , \36137 );
xor \U$36382 ( \36725 , \36724 , \36187 );
xor \U$36383 ( \36726 , \36723 , \36725 );
xor \U$36384 ( \36727 , \36237 , \36247 );
xor \U$36385 ( \36728 , \36727 , \36263 );
not \U$36386 ( \36729 , \36728 );
not \U$36387 ( \36730 , \14930 );
not \U$36388 ( \36731 , \36300 );
or \U$36389 ( \36732 , \36730 , \36731 );
not \U$36390 ( \36733 , RIbb2ddb0_53);
not \U$36391 ( \36734 , \13680 );
or \U$36392 ( \36735 , \36733 , \36734 );
not \U$36393 ( \36736 , \13680 );
nand \U$36394 ( \36737 , \36736 , \12681 );
nand \U$36395 ( \36738 , \36735 , \36737 );
nand \U$36396 ( \36739 , \36738 , \17563 );
nand \U$36397 ( \36740 , \36732 , \36739 );
not \U$36398 ( \36741 , \36740 );
not \U$36399 ( \36742 , \17275 );
not \U$36400 ( \36743 , RIbb2d900_63);
not \U$36401 ( \36744 , \8639 );
or \U$36402 ( \36745 , \36743 , \36744 );
nand \U$36403 ( \36746 , \8638 , \19721 );
nand \U$36404 ( \36747 , \36745 , \36746 );
not \U$36405 ( \36748 , \36747 );
or \U$36406 ( \36749 , \36742 , \36748 );
nand \U$36407 ( \36750 , \36290 , RIbb2d888_64);
nand \U$36408 ( \36751 , \36749 , \36750 );
not \U$36409 ( \36752 , \36751 );
or \U$36410 ( \36753 , \36741 , \36752 );
or \U$36411 ( \36754 , \36751 , \36740 );
not \U$36412 ( \36755 , \14613 );
and \U$36413 ( \36756 , RIbb2dcc0_55, \16601 );
not \U$36414 ( \36757 , RIbb2dcc0_55);
and \U$36415 ( \36758 , \36757 , \16604 );
or \U$36416 ( \36759 , \36756 , \36758 );
not \U$36417 ( \36760 , \36759 );
or \U$36418 ( \36761 , \36755 , \36760 );
not \U$36419 ( \36762 , \27954 );
nand \U$36420 ( \36763 , \36762 , \36154 );
nand \U$36421 ( \36764 , \36761 , \36763 );
nand \U$36422 ( \36765 , \36754 , \36764 );
nand \U$36423 ( \36766 , \36753 , \36765 );
not \U$36424 ( \36767 , \36766 );
or \U$36425 ( \36768 , \36729 , \36767 );
or \U$36426 ( \36769 , \36766 , \36728 );
not \U$36427 ( \36770 , \16675 );
not \U$36428 ( \36771 , RIbb2dbd0_57);
not \U$36429 ( \36772 , \12744 );
or \U$36430 ( \36773 , \36771 , \36772 );
nand \U$36431 ( \36774 , \10301 , \15741 );
nand \U$36432 ( \36775 , \36773 , \36774 );
not \U$36433 ( \36776 , \36775 );
or \U$36434 ( \36777 , \36770 , \36776 );
nand \U$36435 ( \36778 , \36261 , \17100 );
nand \U$36436 ( \36779 , \36777 , \36778 );
not \U$36437 ( \36780 , \36779 );
not \U$36438 ( \36781 , \16541 );
not \U$36439 ( \36782 , RIbb2d9f0_61);
not \U$36440 ( \36783 , \12211 );
or \U$36441 ( \36784 , \36782 , \36783 );
nand \U$36442 ( \36785 , \8321 , \21449 );
nand \U$36443 ( \36786 , \36784 , \36785 );
not \U$36444 ( \36787 , \36786 );
or \U$36445 ( \36788 , \36781 , \36787 );
nand \U$36446 ( \36789 , \36146 , \26834 );
nand \U$36447 ( \36790 , \36788 , \36789 );
not \U$36448 ( \36791 , \36790 );
or \U$36449 ( \36792 , \36780 , \36791 );
or \U$36450 ( \36793 , \36790 , \36779 );
not \U$36451 ( \36794 , \10119 );
not \U$36452 ( \36795 , \36694 );
or \U$36453 ( \36796 , \36794 , \36795 );
not \U$36454 ( \36797 , RIbb2e170_45);
not \U$36455 ( \36798 , \16844 );
or \U$36456 ( \36799 , \36797 , \36798 );
nand \U$36457 ( \36800 , \15825 , \17970 );
nand \U$36458 ( \36801 , \36799 , \36800 );
nand \U$36459 ( \36802 , \36801 , \10599 );
nand \U$36460 ( \36803 , \36796 , \36802 );
not \U$36461 ( \36804 , \36803 );
not \U$36462 ( \36805 , \9099 );
not \U$36463 ( \36806 , \36670 );
or \U$36464 ( \36807 , \36805 , \36806 );
not \U$36465 ( \36808 , RIbb2e260_43);
not \U$36466 ( \36809 , \27577 );
or \U$36467 ( \36810 , \36808 , \36809 );
not \U$36468 ( \36811 , \35763 );
nand \U$36469 ( \36812 , \36811 , \13772 );
nand \U$36470 ( \36813 , \36810 , \36812 );
nand \U$36471 ( \36814 , \36813 , \9098 );
nand \U$36472 ( \36815 , \36807 , \36814 );
not \U$36473 ( \36816 , \36815 );
and \U$36474 ( \36817 , \36804 , \36816 );
or \U$36475 ( \36818 , RIbb2e3c8_40, RIbb2e350_41);
nand \U$36476 ( \36819 , \36818 , \17506 );
and \U$36477 ( \36820 , RIbb2e3c8_40, RIbb2e350_41);
nor \U$36478 ( \36821 , \36820 , \10908 );
nand \U$36479 ( \36822 , \36819 , \36821 );
not \U$36480 ( \36823 , \36822 );
not \U$36481 ( \36824 , \7104 );
not \U$36482 ( \36825 , \36649 );
or \U$36483 ( \36826 , \36824 , \36825 );
and \U$36484 ( \36827 , RIbb2e440_39, \17506 );
not \U$36485 ( \36828 , RIbb2e440_39);
and \U$36486 ( \36829 , \36828 , \20747 );
nor \U$36487 ( \36830 , \36827 , \36829 );
nand \U$36488 ( \36831 , \36830 , \7102 );
nand \U$36489 ( \36832 , \36826 , \36831 );
nand \U$36490 ( \36833 , \36823 , \36832 );
nor \U$36491 ( \36834 , \36817 , \36833 );
and \U$36492 ( \36835 , \36803 , \36815 );
nor \U$36493 ( \36836 , \36834 , \36835 );
not \U$36494 ( \36837 , \36836 );
nand \U$36495 ( \36838 , \36793 , \36837 );
nand \U$36496 ( \36839 , \36792 , \36838 );
nand \U$36497 ( \36840 , \36769 , \36839 );
nand \U$36498 ( \36841 , \36768 , \36840 );
and \U$36499 ( \36842 , \36726 , \36841 );
and \U$36500 ( \36843 , \36723 , \36725 );
or \U$36501 ( \36844 , \36842 , \36843 );
not \U$36502 ( \36845 , \36844 );
nand \U$36503 ( \36846 , \36639 , \36845 );
and \U$36504 ( \36847 , \36636 , \36846 );
nor \U$36505 ( \36848 , \36639 , \36845 );
nor \U$36506 ( \36849 , \36847 , \36848 );
xor \U$36507 ( \36850 , \36584 , \36593 );
xnor \U$36508 ( \36851 , \36850 , \36606 );
nand \U$36509 ( \36852 , \36849 , \36851 );
not \U$36510 ( \36853 , \36852 );
or \U$36511 ( \36854 , \36618 , \36853 );
not \U$36512 ( \36855 , \36849 );
not \U$36513 ( \36856 , \36851 );
nand \U$36514 ( \36857 , \36855 , \36856 );
nand \U$36515 ( \36858 , \36854 , \36857 );
not \U$36516 ( \36859 , \36858 );
nand \U$36517 ( \36860 , \36615 , \36859 );
xor \U$36518 ( \36861 , \36110 , \36497 );
and \U$36519 ( \36862 , \36861 , \36613 );
and \U$36520 ( \36863 , \36110 , \36497 );
or \U$36521 ( \36864 , \36862 , \36863 );
not \U$36522 ( \36865 , \36864 );
or \U$36523 ( \36866 , \36565 , \36576 );
not \U$36524 ( \36867 , \36561 );
nand \U$36525 ( \36868 , \36866 , \36867 );
nand \U$36526 ( \36869 , \36565 , \36576 );
nand \U$36527 ( \36870 , \36868 , \36869 );
not \U$36528 ( \36871 , \36870 );
not \U$36529 ( \36872 , \36046 );
not \U$36530 ( \36873 , \36060 );
or \U$36531 ( \36874 , \36872 , \36873 );
or \U$36532 ( \36875 , \36060 , \36046 );
nand \U$36533 ( \36876 , \36875 , \36036 );
nand \U$36534 ( \36877 , \36874 , \36876 );
xor \U$36535 ( \36878 , \36023 , \36029 );
and \U$36536 ( \36879 , \36878 , \36035 );
and \U$36537 ( \36880 , \36023 , \36029 );
or \U$36538 ( \36881 , \36879 , \36880 );
not \U$36539 ( \36882 , \16533 );
not \U$36540 ( \36883 , \35097 );
or \U$36541 ( \36884 , \36882 , \36883 );
nand \U$36542 ( \36885 , \36093 , \18717 );
nand \U$36543 ( \36886 , \36884 , \36885 );
xor \U$36544 ( \36887 , \36881 , \36886 );
or \U$36545 ( \36888 , \35083 , \27954 );
nand \U$36546 ( \36889 , \35845 , \14613 );
nand \U$36547 ( \36890 , \36888 , \36889 );
xor \U$36548 ( \36891 , \36887 , \36890 );
xor \U$36549 ( \36892 , \36877 , \36891 );
not \U$36550 ( \36893 , \14930 );
not \U$36551 ( \36894 , \34853 );
or \U$36552 ( \36895 , \36893 , \36894 );
nand \U$36553 ( \36896 , \35867 , \17562 );
nand \U$36554 ( \36897 , \36895 , \36896 );
not \U$36555 ( \36898 , \17100 );
not \U$36556 ( \36899 , \34842 );
or \U$36557 ( \36900 , \36898 , \36899 );
nand \U$36558 ( \36901 , \36082 , \19101 );
nand \U$36559 ( \36902 , \36900 , \36901 );
and \U$36560 ( \36903 , \36897 , \36902 );
not \U$36561 ( \36904 , \36897 );
not \U$36562 ( \36905 , \36902 );
and \U$36563 ( \36906 , \36904 , \36905 );
nor \U$36564 ( \36907 , \36903 , \36906 );
not \U$36565 ( \36908 , \17470 );
not \U$36566 ( \36909 , \34999 );
or \U$36567 ( \36910 , \36908 , \36909 );
nand \U$36568 ( \36911 , \36052 , \16271 );
nand \U$36569 ( \36912 , \36910 , \36911 );
and \U$36570 ( \36913 , \36907 , \36912 );
not \U$36571 ( \36914 , \36907 );
not \U$36572 ( \36915 , \36912 );
and \U$36573 ( \36916 , \36914 , \36915 );
nor \U$36574 ( \36917 , \36913 , \36916 );
xnor \U$36575 ( \36918 , \36892 , \36917 );
not \U$36576 ( \36919 , \36918 );
xor \U$36577 ( \36920 , \35892 , \35935 );
and \U$36578 ( \36921 , \36920 , \36016 );
and \U$36579 ( \36922 , \35892 , \35935 );
or \U$36580 ( \36923 , \36921 , \36922 );
not \U$36581 ( \36924 , \36923 );
and \U$36582 ( \36925 , \36919 , \36924 );
and \U$36583 ( \36926 , \36918 , \36923 );
nor \U$36584 ( \36927 , \36925 , \36926 );
not \U$36585 ( \36928 , \36927 );
or \U$36586 ( \36929 , \36871 , \36928 );
or \U$36587 ( \36930 , \36870 , \36927 );
nand \U$36588 ( \36931 , \36929 , \36930 );
not \U$36589 ( \36932 , \36502 );
not \U$36590 ( \36933 , \36577 );
not \U$36591 ( \36934 , \36933 );
or \U$36592 ( \36935 , \36932 , \36934 );
or \U$36593 ( \36936 , \36933 , \36502 );
nand \U$36594 ( \36937 , \36936 , \36608 );
nand \U$36595 ( \36938 , \36935 , \36937 );
xor \U$36596 ( \36939 , \36931 , \36938 );
not \U$36597 ( \36940 , \35981 );
nand \U$36598 ( \36941 , \36940 , \36015 );
and \U$36599 ( \36942 , \36941 , \35940 );
nor \U$36600 ( \36943 , \36015 , \35982 );
nor \U$36601 ( \36944 , \36942 , \36943 );
not \U$36602 ( \36945 , \36944 );
not \U$36603 ( \36946 , \12692 );
not \U$36604 ( \36947 , \35008 );
or \U$36605 ( \36948 , \36946 , \36947 );
nand \U$36606 ( \36949 , \36044 , \14067 );
nand \U$36607 ( \36950 , \36948 , \36949 );
not \U$36608 ( \36951 , RIbb2d888_64);
not \U$36609 ( \36952 , \35019 );
or \U$36610 ( \36953 , \36951 , \36952 );
nand \U$36611 ( \36954 , \35882 , \17275 );
nand \U$36612 ( \36955 , \36953 , \36954 );
xor \U$36613 ( \36956 , \36950 , \36955 );
xor \U$36614 ( \36957 , \36506 , \36511 );
and \U$36615 ( \36958 , \36957 , \36517 );
and \U$36616 ( \36959 , \36506 , \36511 );
or \U$36617 ( \36960 , \36958 , \36959 );
xnor \U$36618 ( \36961 , \36956 , \36960 );
and \U$36619 ( \36962 , \36945 , \36961 );
not \U$36620 ( \36963 , \36945 );
not \U$36621 ( \36964 , \36961 );
and \U$36622 ( \36965 , \36963 , \36964 );
or \U$36623 ( \36966 , \36962 , \36965 );
nor \U$36624 ( \36967 , \36560 , \36518 );
not \U$36625 ( \36968 , \36538 );
or \U$36626 ( \36969 , \36967 , \36968 );
nand \U$36627 ( \36970 , \36560 , \36518 );
nand \U$36628 ( \36971 , \36969 , \36970 );
buf \U$36629 ( \36972 , \36971 );
xor \U$36630 ( \36973 , \36966 , \36972 );
not \U$36631 ( \36974 , \36064 );
not \U$36632 ( \36975 , \36096 );
not \U$36633 ( \36976 , \36975 );
or \U$36634 ( \36977 , \36974 , \36976 );
not \U$36635 ( \36978 , \36061 );
not \U$36636 ( \36979 , \36096 );
or \U$36637 ( \36980 , \36978 , \36979 );
nand \U$36638 ( \36981 , \36980 , \36022 );
nand \U$36639 ( \36982 , \36977 , \36981 );
xor \U$36640 ( \36983 , \34907 , \34921 );
xor \U$36641 ( \36984 , \36983 , \34937 );
or \U$36642 ( \36985 , \35891 , \35869 );
nand \U$36643 ( \36986 , \36985 , \35854 );
nand \U$36644 ( \36987 , \35891 , \35869 );
nand \U$36645 ( \36988 , \36986 , \36987 );
xor \U$36646 ( \36989 , \36984 , \36988 );
xor \U$36647 ( \36990 , \34822 , \34823 );
xor \U$36648 ( \36991 , \36990 , \34834 );
not \U$36649 ( \36992 , \12965 );
not \U$36650 ( \36993 , \35074 );
or \U$36651 ( \36994 , \36992 , \36993 );
nand \U$36652 ( \36995 , \36006 , \11176 );
nand \U$36653 ( \36996 , \36994 , \36995 );
xor \U$36654 ( \36997 , \36991 , \36996 );
not \U$36655 ( \36998 , \12167 );
not \U$36656 ( \36999 , \35991 );
or \U$36657 ( \37000 , \36998 , \36999 );
nand \U$36658 ( \37001 , \35058 , \16427 );
nand \U$36659 ( \37002 , \37000 , \37001 );
xor \U$36660 ( \37003 , \36997 , \37002 );
xor \U$36661 ( \37004 , \36989 , \37003 );
xor \U$36662 ( \37005 , \36982 , \37004 );
xor \U$36663 ( \37006 , \34953 , \34978 );
xor \U$36664 ( \37007 , \37006 , \34989 );
not \U$36665 ( \37008 , \36010 );
nand \U$36666 ( \37009 , \37008 , \35999 );
not \U$36667 ( \37010 , \37009 );
not \U$36668 ( \37011 , \35993 );
or \U$36669 ( \37012 , \37010 , \37011 );
nand \U$36670 ( \37013 , \36010 , \35998 );
nand \U$36671 ( \37014 , \37012 , \37013 );
xor \U$36672 ( \37015 , \37007 , \37014 );
not \U$36673 ( \37016 , \36095 );
not \U$36674 ( \37017 , \36084 );
or \U$36675 ( \37018 , \37016 , \37017 );
or \U$36676 ( \37019 , \36084 , \36095 );
nand \U$36677 ( \37020 , \37019 , \36070 );
nand \U$36678 ( \37021 , \37018 , \37020 );
xor \U$36679 ( \37022 , \37015 , \37021 );
xor \U$36680 ( \37023 , \37005 , \37022 );
xor \U$36681 ( \37024 , \36973 , \37023 );
not \U$36682 ( \37025 , \36102 );
or \U$36683 ( \37026 , \35839 , \37025 );
nand \U$36684 ( \37027 , \37026 , \36017 );
nand \U$36685 ( \37028 , \35839 , \37025 );
nand \U$36686 ( \37029 , \37027 , \37028 );
xor \U$36687 ( \37030 , \37024 , \37029 );
xor \U$36688 ( \37031 , \36939 , \37030 );
not \U$36689 ( \37032 , \37031 );
nand \U$36690 ( \37033 , \36865 , \37032 );
and \U$36691 ( \37034 , \36860 , \37033 );
xor \U$36692 ( \37035 , \35041 , \35065 );
xor \U$36693 ( \37036 , \37035 , \35104 );
xor \U$36694 ( \37037 , \35046 , \35051 );
xor \U$36695 ( \37038 , \37037 , \35062 );
not \U$36696 ( \37039 , \37038 );
xor \U$36697 ( \37040 , \36991 , \36996 );
and \U$36698 ( \37041 , \37040 , \37002 );
and \U$36699 ( \37042 , \36991 , \36996 );
or \U$36700 ( \37043 , \37041 , \37042 );
not \U$36701 ( \37044 , \37043 );
or \U$36702 ( \37045 , \37039 , \37044 );
or \U$36703 ( \37046 , \37043 , \37038 );
xor \U$36704 ( \37047 , \36881 , \36886 );
and \U$36705 ( \37048 , \37047 , \36890 );
and \U$36706 ( \37049 , \36881 , \36886 );
or \U$36707 ( \37050 , \37048 , \37049 );
nand \U$36708 ( \37051 , \37046 , \37050 );
nand \U$36709 ( \37052 , \37045 , \37051 );
xor \U$36710 ( \37053 , \37036 , \37052 );
not \U$36711 ( \37054 , \34807 );
not \U$36712 ( \37055 , \34810 );
and \U$36713 ( \37056 , \37054 , \37055 );
and \U$36714 ( \37057 , \34807 , \34810 );
nor \U$36715 ( \37058 , \37056 , \37057 );
xor \U$36716 ( \37059 , \37058 , \34860 );
not \U$36717 ( \37060 , \37059 );
and \U$36718 ( \37061 , \37053 , \37060 );
not \U$36719 ( \37062 , \37053 );
and \U$36720 ( \37063 , \37062 , \37059 );
nor \U$36721 ( \37064 , \37061 , \37063 );
xor \U$36722 ( \37065 , \34994 , \35026 );
xor \U$36723 ( \37066 , \37065 , \35029 );
and \U$36724 ( \37067 , \37064 , \37066 );
not \U$36725 ( \37068 , \37064 );
not \U$36726 ( \37069 , \37066 );
and \U$36727 ( \37070 , \37068 , \37069 );
nor \U$36728 ( \37071 , \37067 , \37070 );
xor \U$36729 ( \37072 , \36984 , \36988 );
and \U$36730 ( \37073 , \37072 , \37003 );
and \U$36731 ( \37074 , \36984 , \36988 );
or \U$36732 ( \37075 , \37073 , \37074 );
not \U$36733 ( \37076 , \37075 );
or \U$36734 ( \37077 , \36917 , \36891 );
nand \U$36735 ( \37078 , \37077 , \36877 );
nand \U$36736 ( \37079 , \36917 , \36891 );
nand \U$36737 ( \37080 , \37078 , \37079 );
not \U$36738 ( \37081 , \37080 );
or \U$36739 ( \37082 , \37076 , \37081 );
or \U$36740 ( \37083 , \37080 , \37075 );
xor \U$36741 ( \37084 , \34782 , \34791 );
xor \U$36742 ( \37085 , \37084 , \34804 );
not \U$36743 ( \37086 , \36905 );
not \U$36744 ( \37087 , \36915 );
or \U$36745 ( \37088 , \37086 , \37087 );
nand \U$36746 ( \37089 , \37088 , \36897 );
nand \U$36747 ( \37090 , \36912 , \36902 );
nand \U$36748 ( \37091 , \37089 , \37090 );
xor \U$36749 ( \37092 , \37085 , \37091 );
xor \U$36750 ( \37093 , \35076 , \35099 );
xor \U$36751 ( \37094 , \37093 , \35102 );
xor \U$36752 ( \37095 , \37092 , \37094 );
nand \U$36753 ( \37096 , \37083 , \37095 );
nand \U$36754 ( \37097 , \37082 , \37096 );
and \U$36755 ( \37098 , \37071 , \37097 );
not \U$36756 ( \37099 , \37071 );
not \U$36757 ( \37100 , \37097 );
and \U$36758 ( \37101 , \37099 , \37100 );
nor \U$36759 ( \37102 , \37098 , \37101 );
xor \U$36760 ( \37103 , \37075 , \37095 );
xnor \U$36761 ( \37104 , \37103 , \37080 );
xor \U$36762 ( \37105 , \34940 , \34992 );
xnor \U$36763 ( \37106 , \37105 , \34895 );
xor \U$36764 ( \37107 , \37007 , \37014 );
and \U$36765 ( \37108 , \37107 , \37021 );
and \U$36766 ( \37109 , \37007 , \37014 );
or \U$36767 ( \37110 , \37108 , \37109 );
xor \U$36768 ( \37111 , \37106 , \37110 );
xor \U$36769 ( \37112 , \37050 , \37038 );
xnor \U$36770 ( \37113 , \37112 , \37043 );
not \U$36771 ( \37114 , \37113 );
and \U$36772 ( \37115 , \37111 , \37114 );
not \U$36773 ( \37116 , \37111 );
and \U$36774 ( \37117 , \37116 , \37113 );
nor \U$36775 ( \37118 , \37115 , \37117 );
nand \U$36776 ( \37119 , \37104 , \37118 );
not \U$36777 ( \37120 , \37119 );
xor \U$36778 ( \37121 , \34837 , \34846 );
xor \U$36779 ( \37122 , \37121 , \34857 );
not \U$36780 ( \37123 , \36950 );
not \U$36781 ( \37124 , \36955 );
or \U$36782 ( \37125 , \37123 , \37124 );
or \U$36783 ( \37126 , \36955 , \36950 );
nand \U$36784 ( \37127 , \37126 , \36960 );
nand \U$36785 ( \37128 , \37125 , \37127 );
xnor \U$36786 ( \37129 , \37122 , \37128 );
xor \U$36787 ( \37130 , \35003 , \35012 );
xor \U$36788 ( \37131 , \37130 , \35023 );
xor \U$36789 ( \37132 , \37129 , \37131 );
not \U$36790 ( \37133 , \37132 );
not \U$36791 ( \37134 , \37133 );
not \U$36792 ( \37135 , \36945 );
not \U$36793 ( \37136 , \36964 );
or \U$36794 ( \37137 , \37135 , \37136 );
not \U$36795 ( \37138 , \36944 );
not \U$36796 ( \37139 , \36961 );
or \U$36797 ( \37140 , \37138 , \37139 );
nand \U$36798 ( \37141 , \37140 , \36971 );
nand \U$36799 ( \37142 , \37137 , \37141 );
not \U$36800 ( \37143 , \37142 );
not \U$36801 ( \37144 , \37143 );
or \U$36802 ( \37145 , \37134 , \37144 );
nand \U$36803 ( \37146 , \37142 , \37132 );
nand \U$36804 ( \37147 , \37145 , \37146 );
or \U$36805 ( \37148 , \37022 , \37004 );
nand \U$36806 ( \37149 , \37148 , \36982 );
nand \U$36807 ( \37150 , \37004 , \37022 );
nand \U$36808 ( \37151 , \37149 , \37150 );
and \U$36809 ( \37152 , \37147 , \37151 );
not \U$36810 ( \37153 , \37147 );
not \U$36811 ( \37154 , \37151 );
and \U$36812 ( \37155 , \37153 , \37154 );
nor \U$36813 ( \37156 , \37152 , \37155 );
not \U$36814 ( \37157 , \37156 );
or \U$36815 ( \37158 , \37120 , \37157 );
not \U$36816 ( \37159 , \37104 );
not \U$36817 ( \37160 , \37118 );
nand \U$36818 ( \37161 , \37159 , \37160 );
nand \U$36819 ( \37162 , \37158 , \37161 );
not \U$36820 ( \37163 , \37162 );
not \U$36821 ( \37164 , \37163 );
xor \U$36822 ( \37165 , \37102 , \37164 );
not \U$36823 ( \37166 , \37106 );
not \U$36824 ( \37167 , \37113 );
or \U$36825 ( \37168 , \37166 , \37167 );
nand \U$36826 ( \37169 , \37168 , \37110 );
not \U$36827 ( \37170 , \37106 );
nand \U$36828 ( \37171 , \37170 , \37114 );
nand \U$36829 ( \37172 , \37169 , \37171 );
not \U$36830 ( \37173 , \37133 );
not \U$36831 ( \37174 , \37142 );
or \U$36832 ( \37175 , \37173 , \37174 );
not \U$36833 ( \37176 , \37132 );
not \U$36834 ( \37177 , \37143 );
or \U$36835 ( \37178 , \37176 , \37177 );
nand \U$36836 ( \37179 , \37178 , \37151 );
nand \U$36837 ( \37180 , \37175 , \37179 );
xor \U$36838 ( \37181 , \37172 , \37180 );
xor \U$36839 ( \37182 , \37085 , \37091 );
and \U$36840 ( \37183 , \37182 , \37094 );
and \U$36841 ( \37184 , \37085 , \37091 );
or \U$36842 ( \37185 , \37183 , \37184 );
not \U$36843 ( \37186 , \35122 );
not \U$36844 ( \37187 , \35128 );
or \U$36845 ( \37188 , \37186 , \37187 );
nand \U$36846 ( \37189 , \35127 , \35109 );
nand \U$36847 ( \37190 , \37188 , \37189 );
xor \U$36848 ( \37191 , \37190 , \35119 );
xor \U$36849 ( \37192 , \37185 , \37191 );
or \U$36850 ( \37193 , \37131 , \37122 );
not \U$36851 ( \37194 , \37193 );
not \U$36852 ( \37195 , \37128 );
or \U$36853 ( \37196 , \37194 , \37195 );
nand \U$36854 ( \37197 , \37131 , \37122 );
nand \U$36855 ( \37198 , \37196 , \37197 );
xor \U$36856 ( \37199 , \37192 , \37198 );
xor \U$36857 ( \37200 , \37181 , \37199 );
xnor \U$36858 ( \37201 , \37165 , \37200 );
not \U$36859 ( \37202 , \37160 );
not \U$36860 ( \37203 , \37104 );
or \U$36861 ( \37204 , \37202 , \37203 );
nand \U$36862 ( \37205 , \37159 , \37118 );
nand \U$36863 ( \37206 , \37204 , \37205 );
buf \U$36864 ( \37207 , \37156 );
not \U$36865 ( \37208 , \37207 );
and \U$36866 ( \37209 , \37206 , \37208 );
not \U$36867 ( \37210 , \37206 );
and \U$36868 ( \37211 , \37210 , \37207 );
nor \U$36869 ( \37212 , \37209 , \37211 );
not \U$36870 ( \37213 , \36923 );
nand \U$36871 ( \37214 , \37213 , \36918 );
not \U$36872 ( \37215 , \37214 );
not \U$36873 ( \37216 , \36870 );
or \U$36874 ( \37217 , \37215 , \37216 );
not \U$36875 ( \37218 , \36918 );
nand \U$36876 ( \37219 , \37218 , \36923 );
nand \U$36877 ( \37220 , \37217 , \37219 );
not \U$36878 ( \37221 , \37220 );
nand \U$36879 ( \37222 , \37212 , \37221 );
xor \U$36880 ( \37223 , \36973 , \37023 );
and \U$36881 ( \37224 , \37223 , \37029 );
and \U$36882 ( \37225 , \36973 , \37023 );
or \U$36883 ( \37226 , \37224 , \37225 );
and \U$36884 ( \37227 , \37222 , \37226 );
nor \U$36885 ( \37228 , \37212 , \37221 );
nor \U$36886 ( \37229 , \37227 , \37228 );
nand \U$36887 ( \37230 , \37201 , \37229 );
xor \U$36888 ( \37231 , \36931 , \36938 );
and \U$36889 ( \37232 , \37231 , \37030 );
and \U$36890 ( \37233 , \36931 , \36938 );
or \U$36891 ( \37234 , \37232 , \37233 );
not \U$36892 ( \37235 , \37234 );
not \U$36893 ( \37236 , \37220 );
not \U$36894 ( \37237 , \37226 );
not \U$36895 ( \37238 , \37237 );
or \U$36896 ( \37239 , \37236 , \37238 );
nand \U$36897 ( \37240 , \37226 , \37221 );
nand \U$36898 ( \37241 , \37239 , \37240 );
not \U$36899 ( \37242 , \37212 );
and \U$36900 ( \37243 , \37241 , \37242 );
not \U$36901 ( \37244 , \37241 );
and \U$36902 ( \37245 , \37244 , \37212 );
or \U$36903 ( \37246 , \37243 , \37245 );
nand \U$36904 ( \37247 , \37235 , \37246 );
and \U$36905 ( \37248 , \37034 , \37230 , \37247 );
xor \U$36906 ( \37249 , \35038 , \35136 );
xnor \U$36907 ( \37250 , \37249 , \35036 );
not \U$36908 ( \37251 , \37066 );
not \U$36909 ( \37252 , \37064 );
or \U$36910 ( \37253 , \37251 , \37252 );
or \U$36911 ( \37254 , \37066 , \37064 );
nand \U$36912 ( \37255 , \37254 , \37097 );
nand \U$36913 ( \37256 , \37253 , \37255 );
not \U$36914 ( \37257 , \37256 );
xor \U$36915 ( \37258 , \34878 , \34891 );
xor \U$36916 ( \37259 , \37258 , \35032 );
xor \U$36917 ( \37260 , \35107 , \35130 );
xor \U$36918 ( \37261 , \37260 , \35133 );
not \U$36919 ( \37262 , \37261 );
nand \U$36920 ( \37263 , \37259 , \37262 );
not \U$36921 ( \37264 , \37263 );
or \U$36922 ( \37265 , \37257 , \37264 );
not \U$36923 ( \37266 , \37259 );
nand \U$36924 ( \37267 , \37266 , \37261 );
nand \U$36925 ( \37268 , \37265 , \37267 );
not \U$36926 ( \37269 , \37268 );
xor \U$36927 ( \37270 , \37250 , \37269 );
xor \U$36928 ( \37271 , \34544 , \34597 );
xor \U$36929 ( \37272 , \37271 , \34600 );
not \U$36930 ( \37273 , \37272 );
not \U$36931 ( \37274 , \37273 );
xor \U$36932 ( \37275 , \34766 , \34769 );
xnor \U$36933 ( \37276 , \37275 , \34869 );
not \U$36934 ( \37277 , \37276 );
not \U$36935 ( \37278 , \37277 );
or \U$36936 ( \37279 , \37274 , \37278 );
nand \U$36937 ( \37280 , \37276 , \37272 );
nand \U$36938 ( \37281 , \37279 , \37280 );
not \U$36939 ( \37282 , \34777 );
not \U$36940 ( \37283 , \34775 );
or \U$36941 ( \37284 , \37282 , \37283 );
nand \U$36942 ( \37285 , \34774 , \34778 );
nand \U$36943 ( \37286 , \37284 , \37285 );
xnor \U$36944 ( \37287 , \37286 , \34865 );
not \U$36945 ( \37288 , \37287 );
not \U$36946 ( \37289 , \37288 );
not \U$36947 ( \37290 , \37060 );
not \U$36948 ( \37291 , \37036 );
or \U$36949 ( \37292 , \37290 , \37291 );
not \U$36950 ( \37293 , \37059 );
not \U$36951 ( \37294 , \37036 );
not \U$36952 ( \37295 , \37294 );
or \U$36953 ( \37296 , \37293 , \37295 );
nand \U$36954 ( \37297 , \37296 , \37052 );
nand \U$36955 ( \37298 , \37292 , \37297 );
not \U$36956 ( \37299 , \37298 );
or \U$36957 ( \37300 , \37289 , \37299 );
not \U$36958 ( \37301 , \37298 );
not \U$36959 ( \37302 , \37301 );
not \U$36960 ( \37303 , \37287 );
or \U$36961 ( \37304 , \37302 , \37303 );
xor \U$36962 ( \37305 , \37185 , \37191 );
and \U$36963 ( \37306 , \37305 , \37198 );
and \U$36964 ( \37307 , \37185 , \37191 );
or \U$36965 ( \37308 , \37306 , \37307 );
nand \U$36966 ( \37309 , \37304 , \37308 );
nand \U$36967 ( \37310 , \37300 , \37309 );
not \U$36968 ( \37311 , \37310 );
and \U$36969 ( \37312 , \37281 , \37311 );
not \U$36970 ( \37313 , \37281 );
and \U$36971 ( \37314 , \37313 , \37310 );
nor \U$36972 ( \37315 , \37312 , \37314 );
xor \U$36973 ( \37316 , \37270 , \37315 );
xor \U$36974 ( \37317 , \37287 , \37298 );
xor \U$36975 ( \37318 , \37317 , \37308 );
xor \U$36976 ( \37319 , \37172 , \37180 );
and \U$36977 ( \37320 , \37319 , \37199 );
and \U$36978 ( \37321 , \37172 , \37180 );
or \U$36979 ( \37322 , \37320 , \37321 );
not \U$36980 ( \37323 , \37322 );
xor \U$36981 ( \37324 , \37318 , \37323 );
xor \U$36982 ( \37325 , \37261 , \37259 );
xor \U$36983 ( \37326 , \37325 , \37256 );
and \U$36984 ( \37327 , \37324 , \37326 );
and \U$36985 ( \37328 , \37318 , \37323 );
or \U$36986 ( \37329 , \37327 , \37328 );
nand \U$36987 ( \37330 , \37316 , \37329 );
buf \U$36988 ( \37331 , \37330 );
xor \U$36989 ( \37332 , \37318 , \37323 );
xor \U$36990 ( \37333 , \37332 , \37326 );
buf \U$36991 ( \37334 , \37333 );
not \U$36992 ( \37335 , \37102 );
not \U$36993 ( \37336 , \37162 );
or \U$36994 ( \37337 , \37335 , \37336 );
not \U$36995 ( \37338 , \37162 );
not \U$36996 ( \37339 , \37102 );
nand \U$36997 ( \37340 , \37338 , \37339 );
nand \U$36998 ( \37341 , \37200 , \37340 );
nand \U$36999 ( \37342 , \37337 , \37341 );
not \U$37000 ( \37343 , \37342 );
nand \U$37001 ( \37344 , \37334 , \37343 );
and \U$37002 ( \37345 , \37331 , \37344 );
and \U$37003 ( \37346 , \34604 , \34541 );
not \U$37004 ( \37347 , \34604 );
and \U$37005 ( \37348 , \37347 , \34610 );
nor \U$37006 ( \37349 , \37346 , \37348 );
not \U$37007 ( \37350 , \34608 );
and \U$37008 ( \37351 , \37349 , \37350 );
not \U$37009 ( \37352 , \37349 );
and \U$37010 ( \37353 , \37352 , \34608 );
nor \U$37011 ( \37354 , \37351 , \37353 );
not \U$37012 ( \37355 , \37272 );
not \U$37013 ( \37356 , \37277 );
not \U$37014 ( \37357 , \37356 );
not \U$37015 ( \37358 , \37357 );
or \U$37016 ( \37359 , \37355 , \37358 );
not \U$37017 ( \37360 , \37273 );
not \U$37018 ( \37361 , \37356 );
or \U$37019 ( \37362 , \37360 , \37361 );
nand \U$37020 ( \37363 , \37362 , \37310 );
nand \U$37021 ( \37364 , \37359 , \37363 );
not \U$37022 ( \37365 , \37364 );
xor \U$37023 ( \37366 , \37354 , \37365 );
xor \U$37024 ( \37367 , \34871 , \34874 );
xor \U$37025 ( \37368 , \37367 , \35139 );
xor \U$37026 ( \37369 , \37366 , \37368 );
xor \U$37027 ( \37370 , \37250 , \37269 );
and \U$37028 ( \37371 , \37370 , \37315 );
and \U$37029 ( \37372 , \37250 , \37269 );
or \U$37030 ( \37373 , \37371 , \37372 );
nand \U$37031 ( \37374 , \37369 , \37373 );
buf \U$37032 ( \37375 , \37374 );
xor \U$37033 ( \37376 , \34764 , \35145 );
xor \U$37034 ( \37377 , \37376 , \35148 );
xor \U$37035 ( \37378 , \37354 , \37365 );
and \U$37036 ( \37379 , \37378 , \37368 );
and \U$37037 ( \37380 , \37354 , \37365 );
or \U$37038 ( \37381 , \37379 , \37380 );
nand \U$37039 ( \37382 , \37377 , \37381 );
buf \U$37040 ( \37383 , \37382 );
nand \U$37041 ( \37384 , \37248 , \37345 , \37375 , \37383 );
not \U$37042 ( \37385 , \37384 );
or \U$37043 ( \37386 , RIbb2e2d8_42, RIbb2e260_43);
nand \U$37044 ( \37387 , \37386 , \17506 );
and \U$37045 ( \37388 , RIbb2e2d8_42, RIbb2e260_43);
nor \U$37046 ( \37389 , \37388 , \8357 );
and \U$37047 ( \37390 , \37387 , \37389 );
not \U$37048 ( \37391 , \8353 );
not \U$37049 ( \37392 , RIbb2e350_41);
not \U$37050 ( \37393 , \35601 );
or \U$37051 ( \37394 , \37392 , \37393 );
nand \U$37052 ( \37395 , \34958 , \8357 );
nand \U$37053 ( \37396 , \37394 , \37395 );
not \U$37054 ( \37397 , \37396 );
or \U$37055 ( \37398 , \37391 , \37397 );
or \U$37056 ( \37399 , \19064 , \8357 );
or \U$37057 ( \37400 , \18929 , RIbb2e350_41);
nand \U$37058 ( \37401 , \37399 , \37400 );
nand \U$37059 ( \37402 , \37401 , \8361 );
nand \U$37060 ( \37403 , \37398 , \37402 );
xor \U$37061 ( \37404 , \37390 , \37403 );
not \U$37062 ( \37405 , \9099 );
not \U$37063 ( \37406 , RIbb2e260_43);
not \U$37064 ( \37407 , \27234 );
or \U$37065 ( \37408 , \37406 , \37407 );
nand \U$37066 ( \37409 , \16704 , \10444 );
nand \U$37067 ( \37410 , \37408 , \37409 );
not \U$37068 ( \37411 , \37410 );
or \U$37069 ( \37412 , \37405 , \37411 );
and \U$37070 ( \37413 , \8347 , \16820 );
not \U$37071 ( \37414 , \8347 );
and \U$37072 ( \37415 , \37414 , \16821 );
nor \U$37073 ( \37416 , \37413 , \37415 );
nand \U$37074 ( \37417 , \37416 , \10449 );
nand \U$37075 ( \37418 , \37412 , \37417 );
xor \U$37076 ( \37419 , \37404 , \37418 );
not \U$37077 ( \37420 , \11177 );
not \U$37078 ( \37421 , RIbb2e080_47);
not \U$37079 ( \37422 , \16844 );
or \U$37080 ( \37423 , \37421 , \37422 );
nand \U$37081 ( \37424 , \15825 , \10113 );
nand \U$37082 ( \37425 , \37423 , \37424 );
not \U$37083 ( \37426 , \37425 );
or \U$37084 ( \37427 , \37420 , \37426 );
not \U$37085 ( \37428 , RIbb2e080_47);
not \U$37086 ( \37429 , \32984 );
or \U$37087 ( \37430 , \37428 , \37429 );
nand \U$37088 ( \37431 , \32987 , \22357 );
nand \U$37089 ( \37432 , \37430 , \37431 );
nand \U$37090 ( \37433 , \37432 , \11176 );
nand \U$37091 ( \37434 , \37427 , \37433 );
and \U$37092 ( \37435 , \37419 , \37434 );
and \U$37093 ( \37436 , \37404 , \37418 );
or \U$37094 ( \37437 , \37435 , \37436 );
and \U$37095 ( \37438 , \37390 , \37403 );
not \U$37096 ( \37439 , \10119 );
not \U$37097 ( \37440 , RIbb2e170_45);
not \U$37098 ( \37441 , \16747 );
or \U$37099 ( \37442 , \37440 , \37441 );
nand \U$37100 ( \37443 , \16751 , \12003 );
nand \U$37101 ( \37444 , \37442 , \37443 );
not \U$37102 ( \37445 , \37444 );
or \U$37103 ( \37446 , \37439 , \37445 );
not \U$37104 ( \37447 , RIbb2e170_45);
not \U$37105 ( \37448 , \32993 );
or \U$37106 ( \37449 , \37447 , \37448 );
nand \U$37107 ( \37450 , \36811 , \12003 );
nand \U$37108 ( \37451 , \37449 , \37450 );
nand \U$37109 ( \37452 , \37451 , \10117 );
nand \U$37110 ( \37453 , \37446 , \37452 );
xor \U$37111 ( \37454 , \37438 , \37453 );
not \U$37112 ( \37455 , \11177 );
not \U$37113 ( \37456 , RIbb2e080_47);
not \U$37114 ( \37457 , \15754 );
or \U$37115 ( \37458 , \37456 , \37457 );
nand \U$37116 ( \37459 , \16566 , \10113 );
nand \U$37117 ( \37460 , \37458 , \37459 );
not \U$37118 ( \37461 , \37460 );
or \U$37119 ( \37462 , \37455 , \37461 );
nand \U$37120 ( \37463 , \37425 , \11176 );
nand \U$37121 ( \37464 , \37462 , \37463 );
xor \U$37122 ( \37465 , \37454 , \37464 );
xor \U$37123 ( \37466 , \37437 , \37465 );
not \U$37124 ( \37467 , \14930 );
not \U$37125 ( \37468 , RIbb2ddb0_53);
not \U$37126 ( \37469 , \35633 );
not \U$37127 ( \37470 , \37469 );
or \U$37128 ( \37471 , \37468 , \37470 );
not \U$37129 ( \37472 , \15761 );
nand \U$37130 ( \37473 , \37472 , \13463 );
nand \U$37131 ( \37474 , \37471 , \37473 );
not \U$37132 ( \37475 , \37474 );
or \U$37133 ( \37476 , \37467 , \37475 );
not \U$37134 ( \37477 , RIbb2ddb0_53);
not \U$37135 ( \37478 , \15051 );
or \U$37136 ( \37479 , \37477 , \37478 );
nand \U$37137 ( \37480 , \13547 , \16210 );
nand \U$37138 ( \37481 , \37479 , \37480 );
nand \U$37139 ( \37482 , \37481 , \17562 );
nand \U$37140 ( \37483 , \37476 , \37482 );
not \U$37141 ( \37484 , \12692 );
not \U$37142 ( \37485 , RIbb2dea0_51);
not \U$37143 ( \37486 , \35682 );
or \U$37144 ( \37487 , \37485 , \37486 );
not \U$37145 ( \37488 , RIbb2dea0_51);
not \U$37146 ( \37489 , \14503 );
nand \U$37147 ( \37490 , \37488 , \37489 );
nand \U$37148 ( \37491 , \37487 , \37490 );
not \U$37149 ( \37492 , \37491 );
or \U$37150 ( \37493 , \37484 , \37492 );
and \U$37151 ( \37494 , RIbb2dea0_51, \15037 );
not \U$37152 ( \37495 , RIbb2dea0_51);
and \U$37153 ( \37496 , \37495 , \15036 );
or \U$37154 ( \37497 , \37494 , \37496 );
nand \U$37155 ( \37498 , \37497 , \14067 );
nand \U$37156 ( \37499 , \37493 , \37498 );
xor \U$37157 ( \37500 , \37483 , \37499 );
not \U$37158 ( \37501 , \14613 );
and \U$37159 ( \37502 , RIbb2dcc0_55, \12348 );
not \U$37160 ( \37503 , RIbb2dcc0_55);
and \U$37161 ( \37504 , \37503 , \25984 );
or \U$37162 ( \37505 , \37502 , \37504 );
not \U$37163 ( \37506 , \37505 );
or \U$37164 ( \37507 , \37501 , \37506 );
and \U$37165 ( \37508 , RIbb2dcc0_55, \12934 );
not \U$37166 ( \37509 , RIbb2dcc0_55);
not \U$37167 ( \37510 , \15484 );
and \U$37168 ( \37511 , \37509 , \37510 );
or \U$37169 ( \37512 , \37508 , \37511 );
nand \U$37170 ( \37513 , \37512 , \15181 );
nand \U$37171 ( \37514 , \37507 , \37513 );
and \U$37172 ( \37515 , \37500 , \37514 );
and \U$37173 ( \37516 , \37483 , \37499 );
or \U$37174 ( \37517 , \37515 , \37516 );
xor \U$37175 ( \37518 , \37466 , \37517 );
not \U$37176 ( \37519 , \10119 );
not \U$37177 ( \37520 , \37451 );
or \U$37178 ( \37521 , \37519 , \37520 );
not \U$37179 ( \37522 , RIbb2e170_45);
not \U$37180 ( \37523 , \16706 );
not \U$37181 ( \37524 , \37523 );
or \U$37182 ( \37525 , \37522 , \37524 );
not \U$37183 ( \37526 , \16710 );
nand \U$37184 ( \37527 , \37526 , \13372 );
nand \U$37185 ( \37528 , \37525 , \37527 );
nand \U$37186 ( \37529 , \37528 , \10599 );
nand \U$37187 ( \37530 , \37521 , \37529 );
and \U$37188 ( \37531 , \17506 , \8353 );
not \U$37189 ( \37532 , \37416 );
not \U$37190 ( \37533 , \9099 );
or \U$37191 ( \37534 , \37532 , \37533 );
not \U$37192 ( \37535 , RIbb2e260_43);
not \U$37193 ( \37536 , \35601 );
or \U$37194 ( \37537 , \37535 , \37536 );
nand \U$37195 ( \37538 , \17518 , \17231 );
nand \U$37196 ( \37539 , \37537 , \37538 );
nand \U$37197 ( \37540 , \37539 , \9097 );
nand \U$37198 ( \37541 , \37534 , \37540 );
xor \U$37199 ( \37542 , \37531 , \37541 );
not \U$37200 ( \37543 , \10118 );
not \U$37201 ( \37544 , \37528 );
or \U$37202 ( \37545 , \37543 , \37544 );
not \U$37203 ( \37546 , RIbb2e170_45);
not \U$37204 ( \37547 , \27234 );
or \U$37205 ( \37548 , \37546 , \37547 );
nand \U$37206 ( \37549 , \16704 , \12003 );
nand \U$37207 ( \37550 , \37548 , \37549 );
nand \U$37208 ( \37551 , \37550 , \10117 );
nand \U$37209 ( \37552 , \37545 , \37551 );
and \U$37210 ( \37553 , \37542 , \37552 );
and \U$37211 ( \37554 , \37531 , \37541 );
or \U$37212 ( \37555 , \37553 , \37554 );
xor \U$37213 ( \37556 , \37530 , \37555 );
not \U$37214 ( \37557 , \12285 );
not \U$37215 ( \37558 , RIbb2df90_49);
not \U$37216 ( \37559 , \15471 );
not \U$37217 ( \37560 , \37559 );
not \U$37218 ( \37561 , \37560 );
or \U$37219 ( \37562 , \37558 , \37561 );
nand \U$37220 ( \37563 , \15032 , \12278 );
nand \U$37221 ( \37564 , \37562 , \37563 );
not \U$37222 ( \37565 , \37564 );
or \U$37223 ( \37566 , \37557 , \37565 );
and \U$37224 ( \37567 , RIbb2df90_49, \16568 );
not \U$37225 ( \37568 , RIbb2df90_49);
and \U$37226 ( \37569 , \37568 , \15755 );
nor \U$37227 ( \37570 , \37567 , \37569 );
nand \U$37228 ( \37571 , \37570 , \12167 );
nand \U$37229 ( \37572 , \37566 , \37571 );
xor \U$37230 ( \37573 , \37556 , \37572 );
xor \U$37231 ( \37574 , \37531 , \37541 );
xor \U$37232 ( \37575 , \37574 , \37552 );
not \U$37233 ( \37576 , \15181 );
not \U$37234 ( \37577 , \37505 );
or \U$37235 ( \37578 , \37576 , \37577 );
and \U$37236 ( \37579 , RIbb2dcc0_55, \15761 );
not \U$37237 ( \37580 , RIbb2dcc0_55);
and \U$37238 ( \37581 , \37580 , \13474 );
or \U$37239 ( \37582 , \37579 , \37581 );
nand \U$37240 ( \37583 , \37582 , \14613 );
nand \U$37241 ( \37584 , \37578 , \37583 );
xor \U$37242 ( \37585 , \37575 , \37584 );
not \U$37243 ( \37586 , \17397 );
not \U$37244 ( \37587 , RIbb2dbd0_57);
not \U$37245 ( \37588 , \22070 );
or \U$37246 ( \37589 , \37587 , \37588 );
nand \U$37247 ( \37590 , \22073 , \16671 );
nand \U$37248 ( \37591 , \37589 , \37590 );
not \U$37249 ( \37592 , \37591 );
or \U$37250 ( \37593 , \37586 , \37592 );
not \U$37251 ( \37594 , RIbb2dbd0_57);
not \U$37252 ( \37595 , \12934 );
or \U$37253 ( \37596 , \37594 , \37595 );
nand \U$37254 ( \37597 , \12933 , \15741 );
nand \U$37255 ( \37598 , \37596 , \37597 );
nand \U$37256 ( \37599 , \37598 , \19101 );
nand \U$37257 ( \37600 , \37593 , \37599 );
and \U$37258 ( \37601 , \37585 , \37600 );
and \U$37259 ( \37602 , \37575 , \37584 );
or \U$37260 ( \37603 , \37601 , \37602 );
xor \U$37261 ( \37604 , \37573 , \37603 );
xor \U$37262 ( \37605 , \37483 , \37499 );
xor \U$37263 ( \37606 , \37605 , \37514 );
and \U$37264 ( \37607 , \37604 , \37606 );
and \U$37265 ( \37608 , \37573 , \37603 );
or \U$37266 ( \37609 , \37607 , \37608 );
xor \U$37267 ( \37610 , \37518 , \37609 );
and \U$37268 ( \37611 , \17506 , \7104 );
not \U$37269 ( \37612 , \8353 );
and \U$37270 ( \37613 , RIbb2e350_41, \32817 );
not \U$37271 ( \37614 , RIbb2e350_41);
and \U$37272 ( \37615 , \37614 , \16820 );
nor \U$37273 ( \37616 , \37613 , \37615 );
not \U$37274 ( \37617 , \37616 );
or \U$37275 ( \37618 , \37612 , \37617 );
nand \U$37276 ( \37619 , \37396 , \8361 );
nand \U$37277 ( \37620 , \37618 , \37619 );
xor \U$37278 ( \37621 , \37611 , \37620 );
not \U$37279 ( \37622 , \9099 );
not \U$37280 ( \37623 , RIbb2e260_43);
not \U$37281 ( \37624 , \34293 );
or \U$37282 ( \37625 , \37623 , \37624 );
not \U$37283 ( \37626 , \37523 );
nand \U$37284 ( \37627 , \37626 , \8347 );
nand \U$37285 ( \37628 , \37625 , \37627 );
not \U$37286 ( \37629 , \37628 );
or \U$37287 ( \37630 , \37622 , \37629 );
nand \U$37288 ( \37631 , \37410 , \9098 );
nand \U$37289 ( \37632 , \37630 , \37631 );
xor \U$37290 ( \37633 , \37621 , \37632 );
not \U$37291 ( \37634 , \16427 );
not \U$37292 ( \37635 , RIbb2df90_49);
not \U$37293 ( \37636 , \14528 );
or \U$37294 ( \37637 , \37635 , \37636 );
nand \U$37295 ( \37638 , \14527 , \12278 );
nand \U$37296 ( \37639 , \37637 , \37638 );
not \U$37297 ( \37640 , \37639 );
or \U$37298 ( \37641 , \37634 , \37640 );
nand \U$37299 ( \37642 , \37564 , \12167 );
nand \U$37300 ( \37643 , \37641 , \37642 );
xor \U$37301 ( \37644 , \37633 , \37643 );
not \U$37302 ( \37645 , \15182 );
not \U$37303 ( \37646 , \22073 );
and \U$37304 ( \37647 , RIbb2dcc0_55, \37646 );
not \U$37305 ( \37648 , RIbb2dcc0_55);
and \U$37306 ( \37649 , \37648 , \36736 );
or \U$37307 ( \37650 , \37647 , \37649 );
not \U$37308 ( \37651 , \37650 );
or \U$37309 ( \37652 , \37645 , \37651 );
nand \U$37310 ( \37653 , \37512 , \14613 );
nand \U$37311 ( \37654 , \37652 , \37653 );
xor \U$37312 ( \37655 , \37644 , \37654 );
not \U$37313 ( \37656 , RIbb2d888_64);
not \U$37314 ( \37657 , RIbb2d900_63);
not \U$37315 ( \37658 , \10175 );
or \U$37316 ( \37659 , \37657 , \37658 );
nand \U$37317 ( \37660 , \8631 , \19721 );
nand \U$37318 ( \37661 , \37659 , \37660 );
not \U$37319 ( \37662 , \37661 );
or \U$37320 ( \37663 , \37656 , \37662 );
not \U$37321 ( \37664 , RIbb2d900_63);
not \U$37322 ( \37665 , \9279 );
or \U$37323 ( \37666 , \37664 , \37665 );
nand \U$37324 ( \37667 , \9860 , \17262 );
nand \U$37325 ( \37668 , \37666 , \37667 );
nand \U$37326 ( \37669 , \37668 , \17275 );
nand \U$37327 ( \37670 , \37663 , \37669 );
not \U$37328 ( \37671 , \37670 );
not \U$37329 ( \37672 , \37671 );
not \U$37330 ( \37673 , \15738 );
not \U$37331 ( \37674 , RIbb2dbd0_57);
not \U$37332 ( \37675 , \11580 );
or \U$37333 ( \37676 , \37674 , \37675 );
nand \U$37334 ( \37677 , \11581 , \15741 );
nand \U$37335 ( \37678 , \37676 , \37677 );
not \U$37336 ( \37679 , \37678 );
or \U$37337 ( \37680 , \37673 , \37679 );
nand \U$37338 ( \37681 , \37591 , \16675 );
nand \U$37339 ( \37682 , \37680 , \37681 );
not \U$37340 ( \37683 , \37682 );
not \U$37341 ( \37684 , \37683 );
or \U$37342 ( \37685 , \37672 , \37684 );
not \U$37343 ( \37686 , \26834 );
not \U$37344 ( \37687 , RIbb2d9f0_61);
not \U$37345 ( \37688 , \12222 );
or \U$37346 ( \37689 , \37687 , \37688 );
nand \U$37347 ( \37690 , \9841 , \16537 );
nand \U$37348 ( \37691 , \37689 , \37690 );
not \U$37349 ( \37692 , \37691 );
or \U$37350 ( \37693 , \37686 , \37692 );
not \U$37351 ( \37694 , RIbb2d9f0_61);
not \U$37352 ( \37695 , \12744 );
or \U$37353 ( \37696 , \37694 , \37695 );
nand \U$37354 ( \37697 , \10301 , \19746 );
nand \U$37355 ( \37698 , \37696 , \37697 );
nand \U$37356 ( \37699 , \37698 , \16541 );
nand \U$37357 ( \37700 , \37693 , \37699 );
nand \U$37358 ( \37701 , \37685 , \37700 );
nand \U$37359 ( \37702 , \37682 , \37670 );
nand \U$37360 ( \37703 , \37701 , \37702 );
xor \U$37361 ( \37704 , \37655 , \37703 );
not \U$37362 ( \37705 , \16541 );
not \U$37363 ( \37706 , \37691 );
or \U$37364 ( \37707 , \37705 , \37706 );
not \U$37365 ( \37708 , RIbb2d9f0_61);
not \U$37366 ( \37709 , \9857 );
or \U$37367 ( \37710 , \37708 , \37709 );
nand \U$37368 ( \37711 , \15128 , \19746 );
nand \U$37369 ( \37712 , \37710 , \37711 );
nand \U$37370 ( \37713 , \37712 , \26834 );
nand \U$37371 ( \37714 , \37707 , \37713 );
not \U$37372 ( \37715 , \16271 );
and \U$37373 ( \37716 , RIbb2dae0_59, \14563 );
not \U$37374 ( \37717 , RIbb2dae0_59);
and \U$37375 ( \37718 , \37717 , \10764 );
or \U$37376 ( \37719 , \37716 , \37718 );
not \U$37377 ( \37720 , \37719 );
or \U$37378 ( \37721 , \37715 , \37720 );
not \U$37379 ( \37722 , RIbb2dae0_59);
not \U$37380 ( \37723 , \12744 );
or \U$37381 ( \37724 , \37722 , \37723 );
not \U$37382 ( \37725 , RIbb2dae0_59);
nand \U$37383 ( \37726 , \37725 , \10301 );
nand \U$37384 ( \37727 , \37724 , \37726 );
nand \U$37385 ( \37728 , \37727 , \17470 );
nand \U$37386 ( \37729 , \37721 , \37728 );
xor \U$37387 ( \37730 , \37714 , \37729 );
not \U$37388 ( \37731 , RIbb2d888_64);
not \U$37389 ( \37732 , RIbb2d900_63);
not \U$37390 ( \37733 , \8320 );
or \U$37391 ( \37734 , \37732 , \37733 );
nand \U$37392 ( \37735 , \8321 , \33296 );
nand \U$37393 ( \37736 , \37734 , \37735 );
not \U$37394 ( \37737 , \37736 );
or \U$37395 ( \37738 , \37731 , \37737 );
nand \U$37396 ( \37739 , \37661 , \17275 );
nand \U$37397 ( \37740 , \37738 , \37739 );
xor \U$37398 ( \37741 , \37730 , \37740 );
xor \U$37399 ( \37742 , \37704 , \37741 );
and \U$37400 ( \37743 , \37610 , \37742 );
and \U$37401 ( \37744 , \37518 , \37609 );
or \U$37402 ( \37745 , \37743 , \37744 );
xor \U$37403 ( \37746 , \37714 , \37729 );
and \U$37404 ( \37747 , \37746 , \37740 );
and \U$37405 ( \37748 , \37714 , \37729 );
or \U$37406 ( \37749 , \37747 , \37748 );
not \U$37407 ( \37750 , \37749 );
not \U$37408 ( \37751 , \12692 );
and \U$37409 ( \37752 , RIbb2dea0_51, \37469 );
not \U$37410 ( \37753 , RIbb2dea0_51);
and \U$37411 ( \37754 , \37753 , \37472 );
or \U$37412 ( \37755 , \37752 , \37754 );
not \U$37413 ( \37756 , \37755 );
or \U$37414 ( \37757 , \37751 , \37756 );
and \U$37415 ( \37758 , RIbb2dea0_51, \13546 );
not \U$37416 ( \37759 , RIbb2dea0_51);
and \U$37417 ( \37760 , \37759 , \15055 );
or \U$37418 ( \37761 , \37758 , \37760 );
nand \U$37419 ( \37762 , \37761 , \12774 );
nand \U$37420 ( \37763 , \37757 , \37762 );
not \U$37421 ( \37764 , \12169 );
not \U$37422 ( \37765 , RIbb2df90_49);
not \U$37423 ( \37766 , \35682 );
or \U$37424 ( \37767 , \37765 , \37766 );
nand \U$37425 ( \37768 , \13980 , \12278 );
nand \U$37426 ( \37769 , \37767 , \37768 );
not \U$37427 ( \37770 , \37769 );
or \U$37428 ( \37771 , \37764 , \37770 );
nand \U$37429 ( \37772 , \37639 , \12167 );
nand \U$37430 ( \37773 , \37771 , \37772 );
xor \U$37431 ( \37774 , \37763 , \37773 );
not \U$37432 ( \37775 , \14930 );
not \U$37433 ( \37776 , RIbb2ddb0_53);
not \U$37434 ( \37777 , \15484 );
or \U$37435 ( \37778 , \37776 , \37777 );
nand \U$37436 ( \37779 , \12933 , \13463 );
nand \U$37437 ( \37780 , \37778 , \37779 );
not \U$37438 ( \37781 , \37780 );
or \U$37439 ( \37782 , \37775 , \37781 );
not \U$37440 ( \37783 , RIbb2ddb0_53);
not \U$37441 ( \37784 , \33497 );
or \U$37442 ( \37785 , \37783 , \37784 );
nand \U$37443 ( \37786 , \25984 , \12681 );
nand \U$37444 ( \37787 , \37785 , \37786 );
nand \U$37445 ( \37788 , \37787 , \17563 );
nand \U$37446 ( \37789 , \37782 , \37788 );
xor \U$37447 ( \37790 , \37774 , \37789 );
not \U$37448 ( \37791 , \15688 );
not \U$37449 ( \37792 , \37787 );
or \U$37450 ( \37793 , \37791 , \37792 );
nand \U$37451 ( \37794 , \37474 , \14920 );
nand \U$37452 ( \37795 , \37793 , \37794 );
not \U$37453 ( \37796 , \12774 );
not \U$37454 ( \37797 , \37491 );
or \U$37455 ( \37798 , \37796 , \37797 );
nand \U$37456 ( \37799 , \37761 , \12692 );
nand \U$37457 ( \37800 , \37798 , \37799 );
xor \U$37458 ( \37801 , \37795 , \37800 );
not \U$37459 ( \37802 , \15738 );
not \U$37460 ( \37803 , RIbb2dbd0_57);
not \U$37461 ( \37804 , \16601 );
or \U$37462 ( \37805 , \37803 , \37804 );
nand \U$37463 ( \37806 , \16604 , \17097 );
nand \U$37464 ( \37807 , \37805 , \37806 );
not \U$37465 ( \37808 , \37807 );
or \U$37466 ( \37809 , \37802 , \37808 );
nand \U$37467 ( \37810 , \37678 , \19101 );
nand \U$37468 ( \37811 , \37809 , \37810 );
and \U$37469 ( \37812 , \37801 , \37811 );
and \U$37470 ( \37813 , \37795 , \37800 );
or \U$37471 ( \37814 , \37812 , \37813 );
xnor \U$37472 ( \37815 , \37790 , \37814 );
not \U$37473 ( \37816 , \37815 );
or \U$37474 ( \37817 , \37750 , \37816 );
or \U$37475 ( \37818 , \37815 , \37749 );
nand \U$37476 ( \37819 , \37817 , \37818 );
not \U$37477 ( \37820 , \36822 );
not \U$37478 ( \37821 , \36832 );
or \U$37479 ( \37822 , \37820 , \37821 );
or \U$37480 ( \37823 , \36832 , \36822 );
nand \U$37481 ( \37824 , \37822 , \37823 );
not \U$37482 ( \37825 , \8353 );
not \U$37483 ( \37826 , \36660 );
or \U$37484 ( \37827 , \37825 , \37826 );
nand \U$37485 ( \37828 , \37616 , \8361 );
nand \U$37486 ( \37829 , \37827 , \37828 );
xor \U$37487 ( \37830 , \37824 , \37829 );
not \U$37488 ( \37831 , \9099 );
not \U$37489 ( \37832 , \36813 );
or \U$37490 ( \37833 , \37831 , \37832 );
nand \U$37491 ( \37834 , \37628 , \10449 );
nand \U$37492 ( \37835 , \37833 , \37834 );
xor \U$37493 ( \37836 , \37830 , \37835 );
not \U$37494 ( \37837 , \15182 );
and \U$37495 ( \37838 , RIbb2dcc0_55, \36296 );
not \U$37496 ( \37839 , RIbb2dcc0_55);
and \U$37497 ( \37840 , \37839 , \22555 );
or \U$37498 ( \37841 , \37838 , \37840 );
not \U$37499 ( \37842 , \37841 );
or \U$37500 ( \37843 , \37837 , \37842 );
nand \U$37501 ( \37844 , \37650 , \14613 );
nand \U$37502 ( \37845 , \37843 , \37844 );
xor \U$37503 ( \37846 , \37836 , \37845 );
not \U$37504 ( \37847 , \17470 );
and \U$37505 ( \37848 , RIbb2dae0_59, \12222 );
not \U$37506 ( \37849 , RIbb2dae0_59);
and \U$37507 ( \37850 , \37849 , \9841 );
or \U$37508 ( \37851 , \37848 , \37850 );
not \U$37509 ( \37852 , \37851 );
or \U$37510 ( \37853 , \37847 , \37852 );
nand \U$37511 ( \37854 , \37727 , \16271 );
nand \U$37512 ( \37855 , \37853 , \37854 );
xor \U$37513 ( \37856 , \37846 , \37855 );
not \U$37514 ( \37857 , \37856 );
not \U$37515 ( \37858 , \37857 );
xor \U$37516 ( \37859 , \37438 , \37453 );
and \U$37517 ( \37860 , \37859 , \37464 );
and \U$37518 ( \37861 , \37438 , \37453 );
or \U$37519 ( \37862 , \37860 , \37861 );
not \U$37520 ( \37863 , \26834 );
not \U$37521 ( \37864 , RIbb2d9f0_61);
not \U$37522 ( \37865 , \12194 );
or \U$37523 ( \37866 , \37864 , \37865 );
nand \U$37524 ( \37867 , \10178 , \16254 );
nand \U$37525 ( \37868 , \37866 , \37867 );
not \U$37526 ( \37869 , \37868 );
or \U$37527 ( \37870 , \37863 , \37869 );
nand \U$37528 ( \37871 , \37712 , \16541 );
nand \U$37529 ( \37872 , \37870 , \37871 );
xor \U$37530 ( \37873 , \37862 , \37872 );
not \U$37531 ( \37874 , \16675 );
not \U$37532 ( \37875 , \37807 );
or \U$37533 ( \37876 , \37874 , \37875 );
and \U$37534 ( \37877 , RIbb2dbd0_57, \12249 );
not \U$37535 ( \37878 , RIbb2dbd0_57);
and \U$37536 ( \37879 , \37878 , \26937 );
or \U$37537 ( \37880 , \37877 , \37879 );
nand \U$37538 ( \37881 , \37880 , \15738 );
nand \U$37539 ( \37882 , \37876 , \37881 );
xnor \U$37540 ( \37883 , \37873 , \37882 );
not \U$37541 ( \37884 , \37883 );
not \U$37542 ( \37885 , \37884 );
or \U$37543 ( \37886 , \37858 , \37885 );
nand \U$37544 ( \37887 , \37883 , \37856 );
nand \U$37545 ( \37888 , \37886 , \37887 );
xor \U$37546 ( \37889 , \37437 , \37465 );
and \U$37547 ( \37890 , \37889 , \37517 );
and \U$37548 ( \37891 , \37437 , \37465 );
or \U$37549 ( \37892 , \37890 , \37891 );
not \U$37550 ( \37893 , \37892 );
and \U$37551 ( \37894 , \37888 , \37893 );
not \U$37552 ( \37895 , \37888 );
and \U$37553 ( \37896 , \37895 , \37892 );
nor \U$37554 ( \37897 , \37894 , \37896 );
xor \U$37555 ( \37898 , \37819 , \37897 );
not \U$37556 ( \37899 , \10117 );
not \U$37557 ( \37900 , \37444 );
or \U$37558 ( \37901 , \37899 , \37900 );
nand \U$37559 ( \37902 , \36801 , \10119 );
nand \U$37560 ( \37903 , \37901 , \37902 );
xor \U$37561 ( \37904 , \37611 , \37620 );
and \U$37562 ( \37905 , \37904 , \37632 );
and \U$37563 ( \37906 , \37611 , \37620 );
or \U$37564 ( \37907 , \37905 , \37906 );
xor \U$37565 ( \37908 , \37903 , \37907 );
not \U$37566 ( \37909 , \11177 );
not \U$37567 ( \37910 , RIbb2e080_47);
not \U$37568 ( \37911 , \37559 );
not \U$37569 ( \37912 , \37911 );
or \U$37570 ( \37913 , \37910 , \37912 );
nand \U$37571 ( \37914 , \15032 , \16163 );
nand \U$37572 ( \37915 , \37913 , \37914 );
not \U$37573 ( \37916 , \37915 );
or \U$37574 ( \37917 , \37909 , \37916 );
nand \U$37575 ( \37918 , \37460 , \11176 );
nand \U$37576 ( \37919 , \37917 , \37918 );
xor \U$37577 ( \37920 , \37908 , \37919 );
not \U$37578 ( \37921 , \17275 );
not \U$37579 ( \37922 , \37736 );
or \U$37580 ( \37923 , \37921 , \37922 );
not \U$37581 ( \37924 , RIbb2d900_63);
not \U$37582 ( \37925 , \10165 );
or \U$37583 ( \37926 , \37924 , \37925 );
nand \U$37584 ( \37927 , \7300 , \17262 );
nand \U$37585 ( \37928 , \37926 , \37927 );
nand \U$37586 ( \37929 , \37928 , RIbb2d888_64);
nand \U$37587 ( \37930 , \37923 , \37929 );
xor \U$37588 ( \37931 , \37920 , \37930 );
xor \U$37589 ( \37932 , \37633 , \37643 );
and \U$37590 ( \37933 , \37932 , \37654 );
and \U$37591 ( \37934 , \37633 , \37643 );
or \U$37592 ( \37935 , \37933 , \37934 );
xor \U$37593 ( \37936 , \37931 , \37935 );
xor \U$37594 ( \37937 , \37530 , \37555 );
and \U$37595 ( \37938 , \37937 , \37572 );
and \U$37596 ( \37939 , \37530 , \37555 );
or \U$37597 ( \37940 , \37938 , \37939 );
xor \U$37598 ( \37941 , \37795 , \37800 );
xor \U$37599 ( \37942 , \37941 , \37811 );
xor \U$37600 ( \37943 , \37940 , \37942 );
xor \U$37601 ( \37944 , \37404 , \37418 );
xor \U$37602 ( \37945 , \37944 , \37434 );
or \U$37603 ( \37946 , RIbb2e1e8_44, RIbb2e170_45);
nand \U$37604 ( \37947 , \37946 , \17506 );
and \U$37605 ( \37948 , RIbb2e1e8_44, RIbb2e170_45);
nor \U$37606 ( \37949 , \37948 , \17231 );
and \U$37607 ( \37950 , \37947 , \37949 );
not \U$37608 ( \37951 , \37539 );
not \U$37609 ( \37952 , \9099 );
or \U$37610 ( \37953 , \37951 , \37952 );
or \U$37611 ( \37954 , \17506 , \17231 );
or \U$37612 ( \37955 , \18929 , RIbb2e260_43);
nand \U$37613 ( \37956 , \37954 , \37955 );
nand \U$37614 ( \37957 , \37956 , \9097 );
nand \U$37615 ( \37958 , \37953 , \37957 );
and \U$37616 ( \37959 , \37950 , \37958 );
not \U$37617 ( \37960 , \11177 );
not \U$37618 ( \37961 , \37432 );
or \U$37619 ( \37962 , \37960 , \37961 );
not \U$37620 ( \37963 , RIbb2e080_47);
not \U$37621 ( \37964 , \32996 );
not \U$37622 ( \37965 , \37964 );
or \U$37623 ( \37966 , \37963 , \37965 );
nand \U$37624 ( \37967 , \32996 , \22357 );
nand \U$37625 ( \37968 , \37966 , \37967 );
nand \U$37626 ( \37969 , \37968 , \11176 );
nand \U$37627 ( \37970 , \37962 , \37969 );
xor \U$37628 ( \37971 , \37959 , \37970 );
not \U$37629 ( \37972 , \12169 );
not \U$37630 ( \37973 , \37570 );
or \U$37631 ( \37974 , \37972 , \37973 );
not \U$37632 ( \37975 , RIbb2df90_49);
not \U$37633 ( \37976 , \16844 );
or \U$37634 ( \37977 , \37975 , \37976 );
nand \U$37635 ( \37978 , \15825 , \12278 );
nand \U$37636 ( \37979 , \37977 , \37978 );
nand \U$37637 ( \37980 , \37979 , \12167 );
nand \U$37638 ( \37981 , \37974 , \37980 );
and \U$37639 ( \37982 , \37971 , \37981 );
and \U$37640 ( \37983 , \37959 , \37970 );
or \U$37641 ( \37984 , \37982 , \37983 );
xor \U$37642 ( \37985 , \37945 , \37984 );
not \U$37643 ( \37986 , \16271 );
and \U$37644 ( \37987 , RIbb2dae0_59, \15188 );
not \U$37645 ( \37988 , RIbb2dae0_59);
and \U$37646 ( \37989 , \37988 , \11145 );
or \U$37647 ( \37990 , \37987 , \37989 );
not \U$37648 ( \37991 , \37990 );
or \U$37649 ( \37992 , \37986 , \37991 );
nand \U$37650 ( \37993 , \37719 , \17470 );
nand \U$37651 ( \37994 , \37992 , \37993 );
and \U$37652 ( \37995 , \37985 , \37994 );
and \U$37653 ( \37996 , \37945 , \37984 );
or \U$37654 ( \37997 , \37995 , \37996 );
and \U$37655 ( \37998 , \37943 , \37997 );
and \U$37656 ( \37999 , \37940 , \37942 );
or \U$37657 ( \38000 , \37998 , \37999 );
xor \U$37658 ( \38001 , \37936 , \38000 );
xor \U$37659 ( \38002 , \37655 , \37703 );
and \U$37660 ( \38003 , \38002 , \37741 );
and \U$37661 ( \38004 , \37655 , \37703 );
or \U$37662 ( \38005 , \38003 , \38004 );
xor \U$37663 ( \38006 , \38001 , \38005 );
xnor \U$37664 ( \38007 , \37898 , \38006 );
or \U$37665 ( \38008 , \37745 , \38007 );
xor \U$37666 ( \38009 , \37940 , \37942 );
xor \U$37667 ( \38010 , \38009 , \37997 );
xor \U$37668 ( \38011 , \37959 , \37970 );
xor \U$37669 ( \38012 , \38011 , \37981 );
not \U$37670 ( \38013 , \15181 );
not \U$37671 ( \38014 , \37582 );
or \U$37672 ( \38015 , \38013 , \38014 );
and \U$37673 ( \38016 , RIbb2dcc0_55, \15051 );
not \U$37674 ( \38017 , RIbb2dcc0_55);
and \U$37675 ( \38018 , \38017 , \13547 );
or \U$37676 ( \38019 , \38016 , \38018 );
nand \U$37677 ( \38020 , \38019 , \14613 );
nand \U$37678 ( \38021 , \38015 , \38020 );
not \U$37679 ( \38022 , \38021 );
not \U$37680 ( \38023 , \38022 );
not \U$37681 ( \38024 , \14929 );
not \U$37682 ( \38025 , RIbb2ddb0_53);
not \U$37683 ( \38026 , \14503 );
or \U$37684 ( \38027 , \38025 , \38026 );
nand \U$37685 ( \38028 , \16320 , \16210 );
nand \U$37686 ( \38029 , \38027 , \38028 );
not \U$37687 ( \38030 , \38029 );
or \U$37688 ( \38031 , \38024 , \38030 );
not \U$37689 ( \38032 , RIbb2ddb0_53);
not \U$37690 ( \38033 , \21770 );
or \U$37691 ( \38034 , \38032 , \38033 );
nand \U$37692 ( \38035 , \14527 , \16210 );
nand \U$37693 ( \38036 , \38034 , \38035 );
nand \U$37694 ( \38037 , \38036 , \17562 );
nand \U$37695 ( \38038 , \38031 , \38037 );
not \U$37696 ( \38039 , \38038 );
not \U$37697 ( \38040 , \38039 );
or \U$37698 ( \38041 , \38023 , \38040 );
not \U$37699 ( \38042 , \12692 );
and \U$37700 ( \38043 , RIbb2dea0_51, \15031 );
not \U$37701 ( \38044 , RIbb2dea0_51);
and \U$37702 ( \38045 , \38044 , \15474 );
or \U$37703 ( \38046 , \38043 , \38045 );
not \U$37704 ( \38047 , \38046 );
or \U$37705 ( \38048 , \38042 , \38047 );
not \U$37706 ( \38049 , RIbb2dea0_51);
not \U$37707 ( \38050 , \16567 );
or \U$37708 ( \38051 , \38049 , \38050 );
or \U$37709 ( \38052 , \21665 , RIbb2dea0_51);
nand \U$37710 ( \38053 , \38051 , \38052 );
nand \U$37711 ( \38054 , \38053 , \14067 );
nand \U$37712 ( \38055 , \38048 , \38054 );
nand \U$37713 ( \38056 , \38041 , \38055 );
nand \U$37714 ( \38057 , \38038 , \38021 );
nand \U$37715 ( \38058 , \38056 , \38057 );
xor \U$37716 ( \38059 , \38012 , \38058 );
not \U$37717 ( \38060 , \11177 );
not \U$37718 ( \38061 , \37968 );
or \U$37719 ( \38062 , \38060 , \38061 );
not \U$37720 ( \38063 , RIbb2e080_47);
not \U$37721 ( \38064 , \16555 );
or \U$37722 ( \38065 , \38063 , \38064 );
nand \U$37723 ( \38066 , \37626 , \10113 );
nand \U$37724 ( \38067 , \38065 , \38066 );
nand \U$37725 ( \38068 , \38067 , \11176 );
nand \U$37726 ( \38069 , \38062 , \38068 );
and \U$37727 ( \38070 , \17506 , \9099 );
not \U$37728 ( \38071 , \10118 );
not \U$37729 ( \38072 , RIbb2e170_45);
not \U$37730 ( \38073 , \16820 );
or \U$37731 ( \38074 , \38072 , \38073 );
nand \U$37732 ( \38075 , \32817 , \12003 );
nand \U$37733 ( \38076 , \38074 , \38075 );
not \U$37734 ( \38077 , \38076 );
or \U$37735 ( \38078 , \38071 , \38077 );
not \U$37736 ( \38079 , \35601 );
and \U$37737 ( \38080 , RIbb2e170_45, \38079 );
not \U$37738 ( \38081 , RIbb2e170_45);
and \U$37739 ( \38082 , \38081 , \17520 );
nor \U$37740 ( \38083 , \38080 , \38082 );
nand \U$37741 ( \38084 , \38083 , \10116 );
nand \U$37742 ( \38085 , \38078 , \38084 );
xor \U$37743 ( \38086 , \38070 , \38085 );
not \U$37744 ( \38087 , \11175 );
not \U$37745 ( \38088 , RIbb2e080_47);
not \U$37746 ( \38089 , \27234 );
or \U$37747 ( \38090 , \38088 , \38089 );
nand \U$37748 ( \38091 , \16704 , \12971 );
nand \U$37749 ( \38092 , \38090 , \38091 );
not \U$37750 ( \38093 , \38092 );
or \U$37751 ( \38094 , \38087 , \38093 );
nand \U$37752 ( \38095 , \38067 , \11174 );
nand \U$37753 ( \38096 , \38094 , \38095 );
and \U$37754 ( \38097 , \38086 , \38096 );
and \U$37755 ( \38098 , \38070 , \38085 );
or \U$37756 ( \38099 , \38097 , \38098 );
xor \U$37757 ( \38100 , \38069 , \38099 );
not \U$37758 ( \38101 , \15738 );
not \U$37759 ( \38102 , \37598 );
or \U$37760 ( \38103 , \38101 , \38102 );
not \U$37761 ( \38104 , RIbb2dbd0_57);
not \U$37762 ( \38105 , \33497 );
or \U$37763 ( \38106 , \38104 , \38105 );
nand \U$37764 ( \38107 , \12349 , \15741 );
nand \U$37765 ( \38108 , \38106 , \38107 );
nand \U$37766 ( \38109 , \38108 , \16674 );
nand \U$37767 ( \38110 , \38103 , \38109 );
and \U$37768 ( \38111 , \38100 , \38110 );
and \U$37769 ( \38112 , \38069 , \38099 );
or \U$37770 ( \38113 , \38111 , \38112 );
and \U$37771 ( \38114 , \38059 , \38113 );
and \U$37772 ( \38115 , \38012 , \38058 );
or \U$37773 ( \38116 , \38114 , \38115 );
not \U$37774 ( \38117 , \38116 );
xnor \U$37775 ( \38118 , \37700 , \37683 );
and \U$37776 ( \38119 , \38118 , \37671 );
not \U$37777 ( \38120 , \38118 );
and \U$37778 ( \38121 , \38120 , \37670 );
nor \U$37779 ( \38122 , \38119 , \38121 );
not \U$37780 ( \38123 , \38122 );
not \U$37781 ( \38124 , \38123 );
or \U$37782 ( \38125 , \38117 , \38124 );
xor \U$37783 ( \38126 , \37575 , \37584 );
xor \U$37784 ( \38127 , \38126 , \37600 );
xor \U$37785 ( \38128 , \37950 , \37958 );
not \U$37786 ( \38129 , \10119 );
not \U$37787 ( \38130 , \37550 );
or \U$37788 ( \38131 , \38129 , \38130 );
nand \U$37789 ( \38132 , \38076 , \10117 );
nand \U$37790 ( \38133 , \38131 , \38132 );
xor \U$37791 ( \38134 , \38128 , \38133 );
not \U$37792 ( \38135 , \12168 );
not \U$37793 ( \38136 , \37979 );
or \U$37794 ( \38137 , \38135 , \38136 );
not \U$37795 ( \38138 , RIbb2df90_49);
not \U$37796 ( \38139 , \32984 );
or \U$37797 ( \38140 , \38138 , \38139 );
nand \U$37798 ( \38141 , \32987 , \12278 );
nand \U$37799 ( \38142 , \38140 , \38141 );
nand \U$37800 ( \38143 , \38142 , \12167 );
nand \U$37801 ( \38144 , \38137 , \38143 );
xor \U$37802 ( \38145 , \38134 , \38144 );
not \U$37803 ( \38146 , \26834 );
not \U$37804 ( \38147 , RIbb2d9f0_61);
not \U$37805 ( \38148 , \12764 );
or \U$37806 ( \38149 , \38147 , \38148 );
nand \U$37807 ( \38150 , \10764 , \19746 );
nand \U$37808 ( \38151 , \38149 , \38150 );
not \U$37809 ( \38152 , \38151 );
or \U$37810 ( \38153 , \38146 , \38152 );
not \U$37811 ( \38154 , RIbb2d9f0_61);
not \U$37812 ( \38155 , \16601 );
or \U$37813 ( \38156 , \38154 , \38155 );
nand \U$37814 ( \38157 , \16604 , \16254 );
nand \U$37815 ( \38158 , \38156 , \38157 );
nand \U$37816 ( \38159 , \38158 , \16541 );
nand \U$37817 ( \38160 , \38153 , \38159 );
xor \U$37818 ( \38161 , \38145 , \38160 );
not \U$37819 ( \38162 , RIbb2d888_64);
not \U$37820 ( \38163 , RIbb2d900_63);
not \U$37821 ( \38164 , \12222 );
or \U$37822 ( \38165 , \38163 , \38164 );
nand \U$37823 ( \38166 , \9841 , \22946 );
nand \U$37824 ( \38167 , \38165 , \38166 );
not \U$37825 ( \38168 , \38167 );
or \U$37826 ( \38169 , \38162 , \38168 );
not \U$37827 ( \38170 , RIbb2d900_63);
not \U$37828 ( \38171 , \12744 );
or \U$37829 ( \38172 , \38170 , \38171 );
nand \U$37830 ( \38173 , \12235 , \17262 );
nand \U$37831 ( \38174 , \38172 , \38173 );
nand \U$37832 ( \38175 , \38174 , \17275 );
nand \U$37833 ( \38176 , \38169 , \38175 );
and \U$37834 ( \38177 , \38161 , \38176 );
and \U$37835 ( \38178 , \38145 , \38160 );
or \U$37836 ( \38179 , \38177 , \38178 );
xor \U$37837 ( \38180 , \38127 , \38179 );
not \U$37838 ( \38181 , \14929 );
not \U$37839 ( \38182 , \37481 );
or \U$37840 ( \38183 , \38181 , \38182 );
nand \U$37841 ( \38184 , \38029 , \17562 );
nand \U$37842 ( \38185 , \38183 , \38184 );
not \U$37843 ( \38186 , \38185 );
not \U$37844 ( \38187 , \12692 );
not \U$37845 ( \38188 , \37497 );
or \U$37846 ( \38189 , \38187 , \38188 );
nand \U$37847 ( \38190 , \38046 , \12774 );
nand \U$37848 ( \38191 , \38189 , \38190 );
xor \U$37849 ( \38192 , \38186 , \38191 );
not \U$37850 ( \38193 , \26834 );
not \U$37851 ( \38194 , \37698 );
or \U$37852 ( \38195 , \38193 , \38194 );
nand \U$37853 ( \38196 , \38151 , \16541 );
nand \U$37854 ( \38197 , \38195 , \38196 );
xnor \U$37855 ( \38198 , \38192 , \38197 );
and \U$37856 ( \38199 , \38180 , \38198 );
and \U$37857 ( \38200 , \38127 , \38179 );
or \U$37858 ( \38201 , \38199 , \38200 );
not \U$37859 ( \38202 , \38116 );
nand \U$37860 ( \38203 , \38122 , \38202 );
nand \U$37861 ( \38204 , \38201 , \38203 );
nand \U$37862 ( \38205 , \38125 , \38204 );
nor \U$37863 ( \38206 , \38010 , \38205 );
not \U$37864 ( \38207 , \38191 );
nand \U$37865 ( \38208 , \38207 , \38186 );
not \U$37866 ( \38209 , \38208 );
not \U$37867 ( \38210 , \38197 );
or \U$37868 ( \38211 , \38209 , \38210 );
nand \U$37869 ( \38212 , \38191 , \38185 );
nand \U$37870 ( \38213 , \38211 , \38212 );
xor \U$37871 ( \38214 , \37945 , \37984 );
xor \U$37872 ( \38215 , \38214 , \37994 );
xor \U$37873 ( \38216 , \38213 , \38215 );
not \U$37874 ( \38217 , \17470 );
not \U$37875 ( \38218 , \37990 );
or \U$37876 ( \38219 , \38217 , \38218 );
not \U$37877 ( \38220 , \29399 );
and \U$37878 ( \38221 , RIbb2dae0_59, \36296 );
not \U$37879 ( \38222 , RIbb2dae0_59);
and \U$37880 ( \38223 , \38222 , \22555 );
or \U$37881 ( \38224 , \38221 , \38223 );
nand \U$37882 ( \38225 , \38220 , \38224 );
nand \U$37883 ( \38226 , \38219 , \38225 );
not \U$37884 ( \38227 , \38226 );
not \U$37885 ( \38228 , \17275 );
not \U$37886 ( \38229 , \38167 );
or \U$37887 ( \38230 , \38228 , \38229 );
nand \U$37888 ( \38231 , \37668 , RIbb2d888_64);
nand \U$37889 ( \38232 , \38230 , \38231 );
not \U$37890 ( \38233 , \38232 );
or \U$37891 ( \38234 , \38227 , \38233 );
or \U$37892 ( \38235 , \38232 , \38226 );
xor \U$37893 ( \38236 , \38128 , \38133 );
and \U$37894 ( \38237 , \38236 , \38144 );
and \U$37895 ( \38238 , \38128 , \38133 );
or \U$37896 ( \38239 , \38237 , \38238 );
nand \U$37897 ( \38240 , \38235 , \38239 );
nand \U$37898 ( \38241 , \38234 , \38240 );
and \U$37899 ( \38242 , \38216 , \38241 );
and \U$37900 ( \38243 , \38213 , \38215 );
or \U$37901 ( \38244 , \38242 , \38243 );
not \U$37902 ( \38245 , \38244 );
or \U$37903 ( \38246 , \38206 , \38245 );
nand \U$37904 ( \38247 , \38205 , \38010 );
nand \U$37905 ( \38248 , \38246 , \38247 );
buf \U$37906 ( \38249 , \38248 );
nand \U$37907 ( \38250 , \38008 , \38249 );
nand \U$37908 ( \38251 , \38007 , \37745 );
nand \U$37909 ( \38252 , \38250 , \38251 );
not \U$37910 ( \38253 , \38252 );
xor \U$37911 ( \38254 , \37903 , \37907 );
and \U$37912 ( \38255 , \38254 , \37919 );
and \U$37913 ( \38256 , \37903 , \37907 );
or \U$37914 ( \38257 , \38255 , \38256 );
xor \U$37915 ( \38258 , \37763 , \37773 );
and \U$37916 ( \38259 , \38258 , \37789 );
and \U$37917 ( \38260 , \37763 , \37773 );
or \U$37918 ( \38261 , \38259 , \38260 );
xor \U$37919 ( \38262 , \38257 , \38261 );
not \U$37920 ( \38263 , \12167 );
not \U$37921 ( \38264 , \37769 );
or \U$37922 ( \38265 , \38263 , \38264 );
nand \U$37923 ( \38266 , \36713 , \12285 );
nand \U$37924 ( \38267 , \38265 , \38266 );
not \U$37925 ( \38268 , \12774 );
not \U$37926 ( \38269 , \37755 );
or \U$37927 ( \38270 , \38268 , \38269 );
nand \U$37928 ( \38271 , \36678 , \12692 );
nand \U$37929 ( \38272 , \38270 , \38271 );
xor \U$37930 ( \38273 , \38267 , \38272 );
not \U$37931 ( \38274 , \17470 );
and \U$37932 ( \38275 , RIbb2dae0_59, \11700 );
not \U$37933 ( \38276 , RIbb2dae0_59);
and \U$37934 ( \38277 , \38276 , \9280 );
or \U$37935 ( \38278 , \38275 , \38277 );
not \U$37936 ( \38279 , \38278 );
or \U$37937 ( \38280 , \38274 , \38279 );
nand \U$37938 ( \38281 , \37851 , \16271 );
nand \U$37939 ( \38282 , \38280 , \38281 );
xor \U$37940 ( \38283 , \38273 , \38282 );
xor \U$37941 ( \38284 , \38262 , \38283 );
or \U$37942 ( \38285 , \37749 , \37814 );
and \U$37943 ( \38286 , \38285 , \37790 );
and \U$37944 ( \38287 , \37749 , \37814 );
nor \U$37945 ( \38288 , \38286 , \38287 );
not \U$37946 ( \38289 , \38288 );
xor \U$37947 ( \38290 , \38284 , \38289 );
xor \U$37948 ( \38291 , \36642 , \36651 );
xor \U$37949 ( \38292 , \38291 , \36662 );
not \U$37950 ( \38293 , \12965 );
not \U$37951 ( \38294 , \36702 );
or \U$37952 ( \38295 , \38293 , \38294 );
nand \U$37953 ( \38296 , \37915 , \11176 );
nand \U$37954 ( \38297 , \38295 , \38296 );
xor \U$37955 ( \38298 , \38292 , \38297 );
not \U$37956 ( \38299 , \14930 );
not \U$37957 ( \38300 , \36738 );
or \U$37958 ( \38301 , \38299 , \38300 );
nand \U$37959 ( \38302 , \37780 , \17563 );
nand \U$37960 ( \38303 , \38301 , \38302 );
xor \U$37961 ( \38304 , \38298 , \38303 );
xor \U$37962 ( \38305 , \37836 , \37845 );
and \U$37963 ( \38306 , \38305 , \37855 );
and \U$37964 ( \38307 , \37836 , \37845 );
or \U$37965 ( \38308 , \38306 , \38307 );
xor \U$37966 ( \38309 , \38304 , \38308 );
or \U$37967 ( \38310 , \37882 , \37872 );
nand \U$37968 ( \38311 , \38310 , \37862 );
nand \U$37969 ( \38312 , \37882 , \37872 );
nand \U$37970 ( \38313 , \38311 , \38312 );
xor \U$37971 ( \38314 , \38309 , \38313 );
xnor \U$37972 ( \38315 , \38290 , \38314 );
xor \U$37973 ( \38316 , \37936 , \38000 );
and \U$37974 ( \38317 , \38316 , \38005 );
and \U$37975 ( \38318 , \37936 , \38000 );
or \U$37976 ( \38319 , \38317 , \38318 );
not \U$37977 ( \38320 , \38319 );
not \U$37978 ( \38321 , \37884 );
or \U$37979 ( \38322 , \37857 , \38321 );
not \U$37980 ( \38323 , \37857 );
not \U$37981 ( \38324 , \38321 );
or \U$37982 ( \38325 , \38323 , \38324 );
nand \U$37983 ( \38326 , \38325 , \37892 );
nand \U$37984 ( \38327 , \38322 , \38326 );
xor \U$37985 ( \38328 , \36833 , \36815 );
xnor \U$37986 ( \38329 , \38328 , \36803 );
not \U$37987 ( \38330 , \15181 );
not \U$37988 ( \38331 , \36759 );
or \U$37989 ( \38332 , \38330 , \38331 );
nand \U$37990 ( \38333 , \37841 , \14613 );
nand \U$37991 ( \38334 , \38332 , \38333 );
xor \U$37992 ( \38335 , \38329 , \38334 );
not \U$37993 ( \38336 , RIbb2d888_64);
not \U$37994 ( \38337 , \36747 );
or \U$37995 ( \38338 , \38336 , \38337 );
nand \U$37996 ( \38339 , \37928 , \17275 );
nand \U$37997 ( \38340 , \38338 , \38339 );
xnor \U$37998 ( \38341 , \38335 , \38340 );
not \U$37999 ( \38342 , \38341 );
xor \U$38000 ( \38343 , \37824 , \37829 );
and \U$38001 ( \38344 , \38343 , \37835 );
and \U$38002 ( \38345 , \37824 , \37829 );
or \U$38003 ( \38346 , \38344 , \38345 );
not \U$38004 ( \38347 , \16533 );
not \U$38005 ( \38348 , \36786 );
or \U$38006 ( \38349 , \38347 , \38348 );
nand \U$38007 ( \38350 , \18717 , \37868 );
nand \U$38008 ( \38351 , \38349 , \38350 );
xor \U$38009 ( \38352 , \38346 , \38351 );
not \U$38010 ( \38353 , \16675 );
not \U$38011 ( \38354 , \37880 );
or \U$38012 ( \38355 , \38353 , \38354 );
nand \U$38013 ( \38356 , \36775 , \15738 );
nand \U$38014 ( \38357 , \38355 , \38356 );
xnor \U$38015 ( \38358 , \38352 , \38357 );
not \U$38016 ( \38359 , \38358 );
not \U$38017 ( \38360 , \38359 );
or \U$38018 ( \38361 , \38342 , \38360 );
not \U$38019 ( \38362 , \38341 );
nand \U$38020 ( \38363 , \38362 , \38358 );
nand \U$38021 ( \38364 , \38361 , \38363 );
xor \U$38022 ( \38365 , \37920 , \37930 );
and \U$38023 ( \38366 , \38365 , \37935 );
and \U$38024 ( \38367 , \37920 , \37930 );
or \U$38025 ( \38368 , \38366 , \38367 );
and \U$38026 ( \38369 , \38364 , \38368 );
not \U$38027 ( \38370 , \38364 );
not \U$38028 ( \38371 , \38368 );
and \U$38029 ( \38372 , \38370 , \38371 );
nor \U$38030 ( \38373 , \38369 , \38372 );
not \U$38031 ( \38374 , \38373 );
and \U$38032 ( \38375 , \38327 , \38374 );
not \U$38033 ( \38376 , \38327 );
and \U$38034 ( \38377 , \38376 , \38373 );
nor \U$38035 ( \38378 , \38375 , \38377 );
not \U$38036 ( \38379 , \38378 );
and \U$38037 ( \38380 , \38320 , \38379 );
and \U$38038 ( \38381 , \38319 , \38378 );
nor \U$38039 ( \38382 , \38380 , \38381 );
xor \U$38040 ( \38383 , \38315 , \38382 );
not \U$38041 ( \38384 , \37819 );
nand \U$38042 ( \38385 , \38384 , \37897 );
not \U$38043 ( \38386 , \38385 );
not \U$38044 ( \38387 , \38006 );
or \U$38045 ( \38388 , \38386 , \38387 );
not \U$38046 ( \38389 , \37897 );
nand \U$38047 ( \38390 , \38389 , \37819 );
nand \U$38048 ( \38391 , \38388 , \38390 );
not \U$38049 ( \38392 , \38391 );
xor \U$38050 ( \38393 , \38383 , \38392 );
nand \U$38051 ( \38394 , \38253 , \38393 );
not \U$38052 ( \38395 , \38394 );
xor \U$38053 ( \38396 , \37518 , \37609 );
xor \U$38054 ( \38397 , \38396 , \37742 );
not \U$38055 ( \38398 , \38397 );
not \U$38056 ( \38399 , \38205 );
not \U$38057 ( \38400 , \38399 );
not \U$38058 ( \38401 , \38010 );
not \U$38059 ( \38402 , \38245 );
or \U$38060 ( \38403 , \38401 , \38402 );
or \U$38061 ( \38404 , \38245 , \38010 );
nand \U$38062 ( \38405 , \38403 , \38404 );
not \U$38063 ( \38406 , \38405 );
and \U$38064 ( \38407 , \38400 , \38406 );
and \U$38065 ( \38408 , \38399 , \38405 );
nor \U$38066 ( \38409 , \38407 , \38408 );
not \U$38067 ( \38410 , \38409 );
or \U$38068 ( \38411 , \38398 , \38410 );
or \U$38069 ( \38412 , \38409 , \38397 );
nand \U$38070 ( \38413 , \38411 , \38412 );
xor \U$38071 ( \38414 , \37573 , \37603 );
xor \U$38072 ( \38415 , \38414 , \37606 );
xor \U$38073 ( \38416 , \38213 , \38215 );
xor \U$38074 ( \38417 , \38416 , \38241 );
xor \U$38075 ( \38418 , \38415 , \38417 );
xor \U$38076 ( \38419 , \38239 , \38226 );
xnor \U$38077 ( \38420 , \38419 , \38232 );
not \U$38078 ( \38421 , \38420 );
not \U$38079 ( \38422 , \17100 );
not \U$38080 ( \38423 , \38108 );
or \U$38081 ( \38424 , \38422 , \38423 );
not \U$38082 ( \38425 , RIbb2dbd0_57);
not \U$38083 ( \38426 , \13475 );
or \U$38084 ( \38427 , \38425 , \38426 );
nand \U$38085 ( \38428 , \13212 , \15741 );
nand \U$38086 ( \38429 , \38427 , \38428 );
nand \U$38087 ( \38430 , \38429 , \19101 );
nand \U$38088 ( \38431 , \38424 , \38430 );
not \U$38089 ( \38432 , \14613 );
not \U$38090 ( \38433 , RIbb2dcc0_55);
not \U$38091 ( \38434 , \13978 );
or \U$38092 ( \38435 , \38433 , \38434 );
not \U$38093 ( \38436 , RIbb2dcc0_55);
nand \U$38094 ( \38437 , \38436 , \37489 );
nand \U$38095 ( \38438 , \38435 , \38437 );
not \U$38096 ( \38439 , \38438 );
or \U$38097 ( \38440 , \38432 , \38439 );
nand \U$38098 ( \38441 , \38019 , \15182 );
nand \U$38099 ( \38442 , \38440 , \38441 );
or \U$38100 ( \38443 , \38431 , \38442 );
xor \U$38101 ( \38444 , \38070 , \38085 );
xor \U$38102 ( \38445 , \38444 , \38096 );
nand \U$38103 ( \38446 , \38443 , \38445 );
nand \U$38104 ( \38447 , \38431 , \38442 );
nand \U$38105 ( \38448 , \38446 , \38447 );
and \U$38106 ( \38449 , \38039 , \38022 );
not \U$38107 ( \38450 , \38039 );
and \U$38108 ( \38451 , \38450 , \38021 );
nor \U$38109 ( \38452 , \38449 , \38451 );
xor \U$38110 ( \38453 , \38452 , \38055 );
xor \U$38111 ( \38454 , \38448 , \38453 );
not \U$38112 ( \38455 , \16541 );
not \U$38113 ( \38456 , RIbb2d9f0_61);
not \U$38114 ( \38457 , \36296 );
or \U$38115 ( \38458 , \38456 , \38457 );
nand \U$38116 ( \38459 , \11581 , \21449 );
nand \U$38117 ( \38460 , \38458 , \38459 );
not \U$38118 ( \38461 , \38460 );
or \U$38119 ( \38462 , \38455 , \38461 );
nand \U$38120 ( \38463 , \38158 , \26834 );
nand \U$38121 ( \38464 , \38462 , \38463 );
not \U$38122 ( \38465 , \38464 );
not \U$38123 ( \38466 , \16257 );
and \U$38124 ( \38467 , RIbb2dae0_59, \12839 );
not \U$38125 ( \38468 , RIbb2dae0_59);
and \U$38126 ( \38469 , \38468 , \12838 );
or \U$38127 ( \38470 , \38467 , \38469 );
not \U$38128 ( \38471 , \38470 );
or \U$38129 ( \38472 , \38466 , \38471 );
and \U$38130 ( \38473 , RIbb2dae0_59, \12323 );
not \U$38131 ( \38474 , RIbb2dae0_59);
and \U$38132 ( \38475 , \38474 , \12324 );
or \U$38133 ( \38476 , \38473 , \38475 );
nand \U$38134 ( \38477 , \38476 , \16271 );
nand \U$38135 ( \38478 , \38472 , \38477 );
not \U$38136 ( \38479 , \38478 );
not \U$38137 ( \38480 , \38036 );
not \U$38138 ( \38481 , \38480 );
not \U$38139 ( \38482 , \13937 );
and \U$38140 ( \38483 , \38481 , \38482 );
not \U$38141 ( \38484 , RIbb2ddb0_53);
not \U$38142 ( \38485 , \15471 );
or \U$38143 ( \38486 , \38484 , \38485 );
nand \U$38144 ( \38487 , \37559 , \26750 );
nand \U$38145 ( \38488 , \38486 , \38487 );
and \U$38146 ( \38489 , \38488 , \14920 );
nor \U$38147 ( \38490 , \38483 , \38489 );
nand \U$38148 ( \38491 , \38479 , \38490 );
not \U$38149 ( \38492 , \38491 );
or \U$38150 ( \38493 , \38465 , \38492 );
not \U$38151 ( \38494 , \38490 );
nand \U$38152 ( \38495 , \38494 , \38478 );
nand \U$38153 ( \38496 , \38493 , \38495 );
and \U$38154 ( \38497 , \38454 , \38496 );
and \U$38155 ( \38498 , \38448 , \38453 );
or \U$38156 ( \38499 , \38497 , \38498 );
not \U$38157 ( \38500 , \38499 );
not \U$38158 ( \38501 , \38500 );
or \U$38159 ( \38502 , \38421 , \38501 );
or \U$38160 ( \38503 , RIbb2e0f8_46, RIbb2e080_47);
nand \U$38161 ( \38504 , \38503 , \17506 );
and \U$38162 ( \38505 , RIbb2e0f8_46, RIbb2e080_47);
nor \U$38163 ( \38506 , \38505 , \11065 );
and \U$38164 ( \38507 , \38504 , \38506 );
not \U$38165 ( \38508 , \10118 );
not \U$38166 ( \38509 , \38083 );
or \U$38167 ( \38510 , \38508 , \38509 );
or \U$38168 ( \38511 , \17506 , \9094 );
or \U$38169 ( \38512 , \18929 , RIbb2e170_45);
nand \U$38170 ( \38513 , \38511 , \38512 );
nand \U$38171 ( \38514 , \38513 , \10116 );
nand \U$38172 ( \38515 , \38510 , \38514 );
and \U$38173 ( \38516 , \38507 , \38515 );
not \U$38174 ( \38517 , \12168 );
not \U$38175 ( \38518 , \38142 );
or \U$38176 ( \38519 , \38517 , \38518 );
not \U$38177 ( \38520 , RIbb2df90_49);
not \U$38178 ( \38521 , \27577 );
or \U$38179 ( \38522 , \38520 , \38521 );
nand \U$38180 ( \38523 , \19831 , \12278 );
nand \U$38181 ( \38524 , \38522 , \38523 );
nand \U$38182 ( \38525 , \38524 , \12167 );
nand \U$38183 ( \38526 , \38519 , \38525 );
xor \U$38184 ( \38527 , \38516 , \38526 );
not \U$38185 ( \38528 , \12692 );
not \U$38186 ( \38529 , \38053 );
or \U$38187 ( \38530 , \38528 , \38529 );
and \U$38188 ( \38531 , RIbb2dea0_51, \16577 );
not \U$38189 ( \38532 , RIbb2dea0_51);
and \U$38190 ( \38533 , \38532 , \15825 );
or \U$38191 ( \38534 , \38531 , \38533 );
nand \U$38192 ( \38535 , \38534 , \12690 );
nand \U$38193 ( \38536 , \38530 , \38535 );
and \U$38194 ( \38537 , \38527 , \38536 );
and \U$38195 ( \38538 , \38516 , \38526 );
or \U$38196 ( \38539 , \38537 , \38538 );
not \U$38197 ( \38540 , \17470 );
not \U$38198 ( \38541 , \38224 );
or \U$38199 ( \38542 , \38540 , \38541 );
nand \U$38200 ( \38543 , \38470 , \16271 );
nand \U$38201 ( \38544 , \38542 , \38543 );
xor \U$38202 ( \38545 , \38539 , \38544 );
xor \U$38203 ( \38546 , \38069 , \38099 );
xor \U$38204 ( \38547 , \38546 , \38110 );
and \U$38205 ( \38548 , \38545 , \38547 );
and \U$38206 ( \38549 , \38539 , \38544 );
or \U$38207 ( \38550 , \38548 , \38549 );
nand \U$38208 ( \38551 , \38502 , \38550 );
not \U$38209 ( \38552 , \38420 );
nand \U$38210 ( \38553 , \38552 , \38499 );
nand \U$38211 ( \38554 , \38551 , \38553 );
and \U$38212 ( \38555 , \38418 , \38554 );
and \U$38213 ( \38556 , \38415 , \38417 );
or \U$38214 ( \38557 , \38555 , \38556 );
not \U$38215 ( \38558 , \38557 );
and \U$38216 ( \38559 , \38413 , \38558 );
not \U$38217 ( \38560 , \38413 );
and \U$38218 ( \38561 , \38560 , \38557 );
nor \U$38219 ( \38562 , \38559 , \38561 );
xor \U$38220 ( \38563 , \38415 , \38417 );
xor \U$38221 ( \38564 , \38563 , \38554 );
not \U$38222 ( \38565 , \38564 );
xor \U$38223 ( \38566 , \38202 , \38123 );
xor \U$38224 ( \38567 , \38566 , \38201 );
nand \U$38225 ( \38568 , \38565 , \38567 );
xor \U$38226 ( \38569 , \38012 , \38058 );
xor \U$38227 ( \38570 , \38569 , \38113 );
not \U$38228 ( \38571 , \38570 );
xor \U$38229 ( \38572 , \38127 , \38179 );
xor \U$38230 ( \38573 , \38572 , \38198 );
not \U$38231 ( \38574 , \38573 );
or \U$38232 ( \38575 , \38571 , \38574 );
or \U$38233 ( \38576 , \38573 , \38570 );
xor \U$38234 ( \38577 , \38539 , \38544 );
xor \U$38235 ( \38578 , \38577 , \38547 );
not \U$38236 ( \38579 , \38578 );
xor \U$38237 ( \38580 , \38145 , \38160 );
xor \U$38238 ( \38581 , \38580 , \38176 );
not \U$38239 ( \38582 , \38581 );
or \U$38240 ( \38583 , \38579 , \38582 );
or \U$38241 ( \38584 , \38581 , \38578 );
xor \U$38242 ( \38585 , \38507 , \38515 );
not \U$38243 ( \38586 , \11174 );
not \U$38244 ( \38587 , \38092 );
or \U$38245 ( \38588 , \38586 , \38587 );
not \U$38246 ( \38589 , RIbb2e080_47);
not \U$38247 ( \38590 , \16820 );
or \U$38248 ( \38591 , \38589 , \38590 );
nand \U$38249 ( \38592 , \18909 , \10113 );
nand \U$38250 ( \38593 , \38591 , \38592 );
nand \U$38251 ( \38594 , \38593 , \11175 );
nand \U$38252 ( \38595 , \38588 , \38594 );
xor \U$38253 ( \38596 , \38585 , \38595 );
not \U$38254 ( \38597 , \12168 );
not \U$38255 ( \38598 , \38524 );
or \U$38256 ( \38599 , \38597 , \38598 );
not \U$38257 ( \38600 , RIbb2df90_49);
not \U$38258 ( \38601 , \34293 );
or \U$38259 ( \38602 , \38600 , \38601 );
nand \U$38260 ( \38603 , \26039 , \12278 );
nand \U$38261 ( \38604 , \38602 , \38603 );
nand \U$38262 ( \38605 , \38604 , \12167 );
nand \U$38263 ( \38606 , \38599 , \38605 );
and \U$38264 ( \38607 , \38596 , \38606 );
and \U$38265 ( \38608 , \38585 , \38595 );
or \U$38266 ( \38609 , \38607 , \38608 );
xor \U$38267 ( \38610 , \38516 , \38526 );
xor \U$38268 ( \38611 , \38610 , \38536 );
xor \U$38269 ( \38612 , \38609 , \38611 );
not \U$38270 ( \38613 , \17275 );
not \U$38271 ( \38614 , RIbb2d900_63);
not \U$38272 ( \38615 , \12249 );
or \U$38273 ( \38616 , \38614 , \38615 );
nand \U$38274 ( \38617 , \10764 , \33296 );
nand \U$38275 ( \38618 , \38616 , \38617 );
not \U$38276 ( \38619 , \38618 );
or \U$38277 ( \38620 , \38613 , \38619 );
nand \U$38278 ( \38621 , \38174 , RIbb2d888_64);
nand \U$38279 ( \38622 , \38620 , \38621 );
and \U$38280 ( \38623 , \38612 , \38622 );
and \U$38281 ( \38624 , \38609 , \38611 );
or \U$38282 ( \38625 , \38623 , \38624 );
nand \U$38283 ( \38626 , \38584 , \38625 );
nand \U$38284 ( \38627 , \38583 , \38626 );
nand \U$38285 ( \38628 , \38576 , \38627 );
nand \U$38286 ( \38629 , \38575 , \38628 );
and \U$38287 ( \38630 , \38568 , \38629 );
nor \U$38288 ( \38631 , \38565 , \38567 );
nor \U$38289 ( \38632 , \38630 , \38631 );
nor \U$38290 ( \38633 , \38562 , \38632 );
not \U$38291 ( \38634 , \38633 );
not \U$38292 ( \38635 , \38397 );
not \U$38293 ( \38636 , \38557 );
or \U$38294 ( \38637 , \38635 , \38636 );
not \U$38295 ( \38638 , \38397 );
not \U$38296 ( \38639 , \38638 );
not \U$38297 ( \38640 , \38558 );
or \U$38298 ( \38641 , \38639 , \38640 );
not \U$38299 ( \38642 , \38409 );
nand \U$38300 ( \38643 , \38641 , \38642 );
nand \U$38301 ( \38644 , \38637 , \38643 );
not \U$38302 ( \38645 , \38644 );
not \U$38303 ( \38646 , \37745 );
and \U$38304 ( \38647 , \38248 , \38646 );
not \U$38305 ( \38648 , \38248 );
and \U$38306 ( \38649 , \38648 , \37745 );
nor \U$38307 ( \38650 , \38647 , \38649 );
xor \U$38308 ( \38651 , \38650 , \38007 );
nand \U$38309 ( \38652 , \38645 , \38651 );
not \U$38310 ( \38653 , \38652 );
or \U$38311 ( \38654 , \38634 , \38653 );
not \U$38312 ( \38655 , \38651 );
nand \U$38313 ( \38656 , \38655 , \38644 );
nand \U$38314 ( \38657 , \38654 , \38656 );
not \U$38315 ( \38658 , \38657 );
or \U$38316 ( \38659 , \38395 , \38658 );
not \U$38317 ( \38660 , \38393 );
buf \U$38318 ( \38661 , \38252 );
nand \U$38319 ( \38662 , \38660 , \38661 );
nand \U$38320 ( \38663 , \38659 , \38662 );
xor \U$38321 ( \38664 , \38315 , \38382 );
and \U$38322 ( \38665 , \38664 , \38392 );
and \U$38323 ( \38666 , \38315 , \38382 );
or \U$38324 ( \38667 , \38665 , \38666 );
or \U$38325 ( \38668 , \38357 , \38351 );
nand \U$38326 ( \38669 , \38668 , \38346 );
nand \U$38327 ( \38670 , \38357 , \38351 );
nand \U$38328 ( \38671 , \38669 , \38670 );
xor \U$38329 ( \38672 , \36696 , \36706 );
xor \U$38330 ( \38673 , \38672 , \36717 );
xor \U$38331 ( \38674 , \36665 , \36674 );
xor \U$38332 ( \38675 , \38674 , \36682 );
and \U$38333 ( \38676 , \38673 , \38675 );
not \U$38334 ( \38677 , \38673 );
not \U$38335 ( \38678 , \38675 );
and \U$38336 ( \38679 , \38677 , \38678 );
nor \U$38337 ( \38680 , \38676 , \38679 );
xor \U$38338 ( \38681 , \38671 , \38680 );
not \U$38339 ( \38682 , \38362 );
not \U$38340 ( \38683 , \38359 );
or \U$38341 ( \38684 , \38682 , \38683 );
not \U$38342 ( \38685 , \38341 );
not \U$38343 ( \38686 , \38358 );
or \U$38344 ( \38687 , \38685 , \38686 );
nand \U$38345 ( \38688 , \38687 , \38368 );
nand \U$38346 ( \38689 , \38684 , \38688 );
xor \U$38347 ( \38690 , \38681 , \38689 );
xor \U$38348 ( \38691 , \38304 , \38308 );
and \U$38349 ( \38692 , \38691 , \38313 );
and \U$38350 ( \38693 , \38304 , \38308 );
or \U$38351 ( \38694 , \38692 , \38693 );
not \U$38352 ( \38695 , \38694 );
xnor \U$38353 ( \38696 , \38690 , \38695 );
not \U$38354 ( \38697 , \38327 );
nand \U$38355 ( \38698 , \38697 , \38374 );
not \U$38356 ( \38699 , \38698 );
not \U$38357 ( \38700 , \38319 );
or \U$38358 ( \38701 , \38699 , \38700 );
nand \U$38359 ( \38702 , \38373 , \38327 );
nand \U$38360 ( \38703 , \38701 , \38702 );
xor \U$38361 ( \38704 , \38696 , \38703 );
xor \U$38362 ( \38705 , \38267 , \38272 );
and \U$38363 ( \38706 , \38705 , \38282 );
and \U$38364 ( \38707 , \38267 , \38272 );
or \U$38365 ( \38708 , \38706 , \38707 );
not \U$38366 ( \38709 , \38334 );
not \U$38367 ( \38710 , \38340 );
or \U$38368 ( \38711 , \38709 , \38710 );
or \U$38369 ( \38712 , \38340 , \38334 );
nand \U$38370 ( \38713 , \38712 , \38329 );
nand \U$38371 ( \38714 , \38711 , \38713 );
xor \U$38372 ( \38715 , \38708 , \38714 );
xor \U$38373 ( \38716 , \36779 , \36836 );
xnor \U$38374 ( \38717 , \38716 , \36790 );
xnor \U$38375 ( \38718 , \38715 , \38717 );
not \U$38376 ( \38719 , \38718 );
xor \U$38377 ( \38720 , \36751 , \36740 );
xnor \U$38378 ( \38721 , \38720 , \36764 );
xor \U$38379 ( \38722 , \36162 , \36171 );
xor \U$38380 ( \38723 , \38722 , \36182 );
not \U$38381 ( \38724 , \16271 );
not \U$38382 ( \38725 , \38278 );
or \U$38383 ( \38726 , \38724 , \38725 );
nand \U$38384 ( \38727 , \36272 , \17470 );
nand \U$38385 ( \38728 , \38726 , \38727 );
xor \U$38386 ( \38729 , \38723 , \38728 );
xor \U$38387 ( \38730 , \38292 , \38297 );
and \U$38388 ( \38731 , \38730 , \38303 );
and \U$38389 ( \38732 , \38292 , \38297 );
or \U$38390 ( \38733 , \38731 , \38732 );
xor \U$38391 ( \38734 , \38729 , \38733 );
xor \U$38392 ( \38735 , \38721 , \38734 );
xor \U$38393 ( \38736 , \38257 , \38261 );
and \U$38394 ( \38737 , \38736 , \38283 );
and \U$38395 ( \38738 , \38257 , \38261 );
or \U$38396 ( \38739 , \38737 , \38738 );
xor \U$38397 ( \38740 , \38735 , \38739 );
xor \U$38398 ( \38741 , \38719 , \38740 );
not \U$38399 ( \38742 , \38284 );
not \U$38400 ( \38743 , \38289 );
or \U$38401 ( \38744 , \38742 , \38743 );
not \U$38402 ( \38745 , \38284 );
not \U$38403 ( \38746 , \38745 );
not \U$38404 ( \38747 , \38288 );
or \U$38405 ( \38748 , \38746 , \38747 );
nand \U$38406 ( \38749 , \38748 , \38314 );
nand \U$38407 ( \38750 , \38744 , \38749 );
xnor \U$38408 ( \38751 , \38741 , \38750 );
xnor \U$38409 ( \38752 , \38704 , \38751 );
nand \U$38410 ( \38753 , \38667 , \38752 );
and \U$38411 ( \38754 , \38663 , \38753 );
nor \U$38412 ( \38755 , \38667 , \38752 );
nor \U$38413 ( \38756 , \38754 , \38755 );
xor \U$38414 ( \38757 , \38625 , \38581 );
xnor \U$38415 ( \38758 , \38757 , \38578 );
and \U$38416 ( \38759 , \17506 , \10118 );
not \U$38417 ( \38760 , \11174 );
not \U$38418 ( \38761 , \38593 );
or \U$38419 ( \38762 , \38760 , \38761 );
and \U$38420 ( \38763 , RIbb2e080_47, \26129 );
not \U$38421 ( \38764 , RIbb2e080_47);
and \U$38422 ( \38765 , \38764 , \20552 );
nor \U$38423 ( \38766 , \38763 , \38765 );
nand \U$38424 ( \38767 , \38766 , \11175 );
nand \U$38425 ( \38768 , \38762 , \38767 );
xor \U$38426 ( \38769 , \38759 , \38768 );
not \U$38427 ( \38770 , \12168 );
not \U$38428 ( \38771 , \38604 );
or \U$38429 ( \38772 , \38770 , \38771 );
not \U$38430 ( \38773 , RIbb2df90_49);
not \U$38431 ( \38774 , \27234 );
or \U$38432 ( \38775 , \38773 , \38774 );
nand \U$38433 ( \38776 , \33477 , \12278 );
nand \U$38434 ( \38777 , \38775 , \38776 );
nand \U$38435 ( \38778 , \38777 , \12167 );
nand \U$38436 ( \38779 , \38772 , \38778 );
and \U$38437 ( \38780 , \38769 , \38779 );
and \U$38438 ( \38781 , \38759 , \38768 );
or \U$38439 ( \38782 , \38780 , \38781 );
not \U$38440 ( \38783 , \12690 );
not \U$38441 ( \38784 , RIbb2dea0_51);
not \U$38442 ( \38785 , \16747 );
or \U$38443 ( \38786 , \38784 , \38785 );
or \U$38444 ( \38787 , \16747 , RIbb2dea0_51);
nand \U$38445 ( \38788 , \38786 , \38787 );
not \U$38446 ( \38789 , \38788 );
or \U$38447 ( \38790 , \38783 , \38789 );
nand \U$38448 ( \38791 , \38534 , \12692 );
nand \U$38449 ( \38792 , \38790 , \38791 );
xor \U$38450 ( \38793 , \38782 , \38792 );
not \U$38451 ( \38794 , \19101 );
not \U$38452 ( \38795 , RIbb2dbd0_57);
not \U$38453 ( \38796 , \13986 );
or \U$38454 ( \38797 , \38795 , \38796 );
nand \U$38455 ( \38798 , \15055 , \15741 );
nand \U$38456 ( \38799 , \38797 , \38798 );
not \U$38457 ( \38800 , \38799 );
or \U$38458 ( \38801 , \38794 , \38800 );
nand \U$38459 ( \38802 , \38429 , \15738 );
nand \U$38460 ( \38803 , \38801 , \38802 );
and \U$38461 ( \38804 , \38793 , \38803 );
and \U$38462 ( \38805 , \38782 , \38792 );
or \U$38463 ( \38806 , \38804 , \38805 );
not \U$38464 ( \38807 , \38806 );
not \U$38465 ( \38808 , \16271 );
and \U$38466 ( \38809 , RIbb2dae0_59, \13809 );
not \U$38467 ( \38810 , RIbb2dae0_59);
and \U$38468 ( \38811 , \38810 , \14839 );
or \U$38469 ( \38812 , \38809 , \38811 );
not \U$38470 ( \38813 , \38812 );
or \U$38471 ( \38814 , \38808 , \38813 );
nand \U$38472 ( \38815 , \38476 , \16257 );
nand \U$38473 ( \38816 , \38814 , \38815 );
not \U$38474 ( \38817 , \15181 );
not \U$38475 ( \38818 , \38438 );
or \U$38476 ( \38819 , \38817 , \38818 );
not \U$38477 ( \38820 , RIbb2dcc0_55);
not \U$38478 ( \38821 , \14528 );
or \U$38479 ( \38822 , \38820 , \38821 );
not \U$38480 ( \38823 , RIbb2dcc0_55);
nand \U$38481 ( \38824 , \38823 , \15036 );
nand \U$38482 ( \38825 , \38822 , \38824 );
nand \U$38483 ( \38826 , \38825 , \14613 );
nand \U$38484 ( \38827 , \38819 , \38826 );
nor \U$38485 ( \38828 , \38816 , \38827 );
not \U$38486 ( \38829 , \14929 );
not \U$38487 ( \38830 , \38488 );
or \U$38488 ( \38831 , \38829 , \38830 );
and \U$38489 ( \38832 , RIbb2ddb0_53, \21665 );
not \U$38490 ( \38833 , RIbb2ddb0_53);
and \U$38491 ( \38834 , \38833 , \15756 );
nor \U$38492 ( \38835 , \38832 , \38834 );
not \U$38493 ( \38836 , \38835 );
nand \U$38494 ( \38837 , \38836 , \13467 );
nand \U$38495 ( \38838 , \38831 , \38837 );
not \U$38496 ( \38839 , \38838 );
or \U$38497 ( \38840 , \38828 , \38839 );
nand \U$38498 ( \38841 , \38827 , \38816 );
nand \U$38499 ( \38842 , \38840 , \38841 );
not \U$38500 ( \38843 , \38842 );
not \U$38501 ( \38844 , \38843 );
or \U$38502 ( \38845 , \38807 , \38844 );
not \U$38503 ( \38846 , \38806 );
nand \U$38504 ( \38847 , \38846 , \38842 );
nand \U$38505 ( \38848 , \38845 , \38847 );
xor \U$38506 ( \38849 , \38445 , \38442 );
xnor \U$38507 ( \38850 , \38849 , \38431 );
and \U$38508 ( \38851 , \38848 , \38850 );
not \U$38509 ( \38852 , \38848 );
not \U$38510 ( \38853 , \38850 );
and \U$38511 ( \38854 , \38852 , \38853 );
nor \U$38512 ( \38855 , \38851 , \38854 );
xor \U$38513 ( \38856 , \38782 , \38792 );
xor \U$38514 ( \38857 , \38856 , \38803 );
not \U$38515 ( \38858 , \16674 );
not \U$38516 ( \38859 , RIbb2dbd0_57);
not \U$38517 ( \38860 , \15456 );
or \U$38518 ( \38861 , \38859 , \38860 );
nand \U$38519 ( \38862 , \13980 , \17097 );
nand \U$38520 ( \38863 , \38861 , \38862 );
not \U$38521 ( \38864 , \38863 );
or \U$38522 ( \38865 , \38858 , \38864 );
nand \U$38523 ( \38866 , \38799 , \17397 );
nand \U$38524 ( \38867 , \38865 , \38866 );
not \U$38525 ( \38868 , \14613 );
and \U$38526 ( \38869 , RIbb2dcc0_55, \37911 );
not \U$38527 ( \38870 , RIbb2dcc0_55);
and \U$38528 ( \38871 , \38870 , \37559 );
or \U$38529 ( \38872 , \38869 , \38871 );
not \U$38530 ( \38873 , \38872 );
or \U$38531 ( \38874 , \38868 , \38873 );
nand \U$38532 ( \38875 , \38825 , \15181 );
nand \U$38533 ( \38876 , \38874 , \38875 );
nor \U$38534 ( \38877 , \38867 , \38876 );
xor \U$38535 ( \38878 , \38759 , \38768 );
xor \U$38536 ( \38879 , \38878 , \38779 );
not \U$38537 ( \38880 , \38879 );
or \U$38538 ( \38881 , \38877 , \38880 );
nand \U$38539 ( \38882 , \38876 , \38867 );
nand \U$38540 ( \38883 , \38881 , \38882 );
xor \U$38541 ( \38884 , \38857 , \38883 );
not \U$38542 ( \38885 , RIbb2d888_64);
not \U$38543 ( \38886 , \38618 );
or \U$38544 ( \38887 , \38885 , \38886 );
not \U$38545 ( \38888 , RIbb2d900_63);
not \U$38546 ( \38889 , \11145 );
not \U$38547 ( \38890 , \38889 );
or \U$38548 ( \38891 , \38888 , \38890 );
nand \U$38549 ( \38892 , \35521 , \17270 );
nand \U$38550 ( \38893 , \38891 , \38892 );
nand \U$38551 ( \38894 , \38893 , \17275 );
nand \U$38552 ( \38895 , \38887 , \38894 );
and \U$38553 ( \38896 , \38884 , \38895 );
and \U$38554 ( \38897 , \38857 , \38883 );
or \U$38555 ( \38898 , \38896 , \38897 );
not \U$38556 ( \38899 , \38898 );
nand \U$38557 ( \38900 , \38855 , \38899 );
not \U$38558 ( \38901 , \38900 );
xor \U$38559 ( \38902 , \38827 , \38816 );
and \U$38560 ( \38903 , \38902 , \38838 );
not \U$38561 ( \38904 , \38902 );
and \U$38562 ( \38905 , \38904 , \38839 );
nor \U$38563 ( \38906 , \38903 , \38905 );
buf \U$38564 ( \38907 , \38906 );
not \U$38565 ( \38908 , \38907 );
not \U$38566 ( \38909 , \17470 );
not \U$38567 ( \38910 , \38812 );
or \U$38568 ( \38911 , \38909 , \38910 );
and \U$38569 ( \38912 , RIbb2dae0_59, \13211 );
not \U$38570 ( \38913 , RIbb2dae0_59);
and \U$38571 ( \38914 , \38913 , \35633 );
or \U$38572 ( \38915 , \38912 , \38914 );
nand \U$38573 ( \38916 , \38915 , \16271 );
nand \U$38574 ( \38917 , \38911 , \38916 );
not \U$38575 ( \38918 , \26834 );
not \U$38576 ( \38919 , RIbb2d9f0_61);
not \U$38577 ( \38920 , \13680 );
or \U$38578 ( \38921 , \38919 , \38920 );
nand \U$38579 ( \38922 , \36736 , \19746 );
nand \U$38580 ( \38923 , \38921 , \38922 );
not \U$38581 ( \38924 , \38923 );
or \U$38582 ( \38925 , \38918 , \38924 );
not \U$38583 ( \38926 , RIbb2d9f0_61);
not \U$38584 ( \38927 , \12934 );
or \U$38585 ( \38928 , \38926 , \38927 );
nand \U$38586 ( \38929 , \12933 , \16254 );
nand \U$38587 ( \38930 , \38928 , \38929 );
nand \U$38588 ( \38931 , \38930 , \16541 );
nand \U$38589 ( \38932 , \38925 , \38931 );
xor \U$38590 ( \38933 , \38917 , \38932 );
not \U$38591 ( \38934 , RIbb2d888_64);
not \U$38592 ( \38935 , \38893 );
or \U$38593 ( \38936 , \38934 , \38935 );
not \U$38594 ( \38937 , RIbb2d900_63);
not \U$38595 ( \38938 , \11580 );
or \U$38596 ( \38939 , \38937 , \38938 );
nand \U$38597 ( \38940 , \22555 , \17262 );
nand \U$38598 ( \38941 , \38939 , \38940 );
nand \U$38599 ( \38942 , \38941 , \17275 );
nand \U$38600 ( \38943 , \38936 , \38942 );
and \U$38601 ( \38944 , \38933 , \38943 );
and \U$38602 ( \38945 , \38917 , \38932 );
or \U$38603 ( \38946 , \38944 , \38945 );
not \U$38604 ( \38947 , \38946 );
or \U$38605 ( \38948 , \38908 , \38947 );
or \U$38606 ( \38949 , \38946 , \38907 );
xor \U$38607 ( \38950 , \38585 , \38595 );
xor \U$38608 ( \38951 , \38950 , \38606 );
or \U$38609 ( \38952 , RIbb2e008_48, RIbb2df90_49);
nand \U$38610 ( \38953 , \38952 , \17506 );
and \U$38611 ( \38954 , RIbb2e008_48, RIbb2df90_49);
nor \U$38612 ( \38955 , \38954 , \10113 );
and \U$38613 ( \38956 , \38953 , \38955 );
not \U$38614 ( \38957 , \11175 );
or \U$38615 ( \38958 , \17506 , \10113 );
or \U$38616 ( \38959 , \18929 , RIbb2e080_47);
nand \U$38617 ( \38960 , \38958 , \38959 );
not \U$38618 ( \38961 , \38960 );
or \U$38619 ( \38962 , \38957 , \38961 );
not \U$38620 ( \38963 , \38766 );
not \U$38621 ( \38964 , \11174 );
or \U$38622 ( \38965 , \38963 , \38964 );
nand \U$38623 ( \38966 , \38962 , \38965 );
and \U$38624 ( \38967 , \38956 , \38966 );
not \U$38625 ( \38968 , \12692 );
not \U$38626 ( \38969 , \38788 );
or \U$38627 ( \38970 , \38968 , \38969 );
and \U$38628 ( \38971 , RIbb2dea0_51, \35763 );
not \U$38629 ( \38972 , RIbb2dea0_51);
and \U$38630 ( \38973 , \38972 , \32996 );
or \U$38631 ( \38974 , \38971 , \38973 );
nand \U$38632 ( \38975 , \38974 , \12690 );
nand \U$38633 ( \38976 , \38970 , \38975 );
xor \U$38634 ( \38977 , \38967 , \38976 );
not \U$38635 ( \38978 , RIbb2ddb0_53);
not \U$38636 ( \38979 , \16577 );
or \U$38637 ( \38980 , \38978 , \38979 );
nand \U$38638 ( \38981 , \15825 , \12681 );
nand \U$38639 ( \38982 , \38980 , \38981 );
not \U$38640 ( \38983 , \38982 );
not \U$38641 ( \38984 , \13467 );
or \U$38642 ( \38985 , \38983 , \38984 );
not \U$38643 ( \38986 , \14929 );
or \U$38644 ( \38987 , \38835 , \38986 );
nand \U$38645 ( \38988 , \38985 , \38987 );
and \U$38646 ( \38989 , \38977 , \38988 );
and \U$38647 ( \38990 , \38967 , \38976 );
or \U$38648 ( \38991 , \38989 , \38990 );
xor \U$38649 ( \38992 , \38951 , \38991 );
not \U$38650 ( \38993 , \26834 );
not \U$38651 ( \38994 , \38460 );
or \U$38652 ( \38995 , \38993 , \38994 );
nand \U$38653 ( \38996 , \38923 , \18717 );
nand \U$38654 ( \38997 , \38995 , \38996 );
xor \U$38655 ( \38998 , \38992 , \38997 );
nand \U$38656 ( \38999 , \38949 , \38998 );
nand \U$38657 ( \39000 , \38948 , \38999 );
not \U$38658 ( \39001 , \39000 );
or \U$38659 ( \39002 , \38901 , \39001 );
not \U$38660 ( \39003 , \38855 );
nand \U$38661 ( \39004 , \39003 , \38898 );
nand \U$38662 ( \39005 , \39002 , \39004 );
not \U$38663 ( \39006 , \39005 );
xor \U$38664 ( \39007 , \38758 , \39006 );
not \U$38665 ( \39008 , \38843 );
not \U$38666 ( \39009 , \38846 );
or \U$38667 ( \39010 , \39008 , \39009 );
nand \U$38668 ( \39011 , \39010 , \38853 );
not \U$38669 ( \39012 , \38843 );
nand \U$38670 ( \39013 , \39012 , \38806 );
nand \U$38671 ( \39014 , \39011 , \39013 );
xor \U$38672 ( \39015 , \38448 , \38453 );
xor \U$38673 ( \39016 , \39015 , \38496 );
xor \U$38674 ( \39017 , \39014 , \39016 );
not \U$38675 ( \39018 , \38464 );
not \U$38676 ( \39019 , \38478 );
not \U$38677 ( \39020 , \38490 );
and \U$38678 ( \39021 , \39019 , \39020 );
and \U$38679 ( \39022 , \38478 , \38490 );
nor \U$38680 ( \39023 , \39021 , \39022 );
not \U$38681 ( \39024 , \39023 );
or \U$38682 ( \39025 , \39018 , \39024 );
or \U$38683 ( \39026 , \38464 , \39023 );
nand \U$38684 ( \39027 , \39025 , \39026 );
not \U$38685 ( \39028 , \39027 );
not \U$38686 ( \39029 , \39028 );
xor \U$38687 ( \39030 , \38951 , \38991 );
and \U$38688 ( \39031 , \39030 , \38997 );
and \U$38689 ( \39032 , \38951 , \38991 );
or \U$38690 ( \39033 , \39031 , \39032 );
not \U$38691 ( \39034 , \39033 );
not \U$38692 ( \39035 , \39034 );
or \U$38693 ( \39036 , \39029 , \39035 );
xor \U$38694 ( \39037 , \38609 , \38611 );
xor \U$38695 ( \39038 , \39037 , \38622 );
nand \U$38696 ( \39039 , \39036 , \39038 );
nand \U$38697 ( \39040 , \39033 , \39027 );
nand \U$38698 ( \39041 , \39039 , \39040 );
xor \U$38699 ( \39042 , \39017 , \39041 );
xnor \U$38700 ( \39043 , \39007 , \39042 );
xor \U$38701 ( \39044 , \39027 , \39034 );
xor \U$38702 ( \39045 , \39044 , \39038 );
not \U$38703 ( \39046 , \39045 );
and \U$38704 ( \39047 , \38899 , \39003 );
not \U$38705 ( \39048 , \38899 );
and \U$38706 ( \39049 , \39048 , \38855 );
nor \U$38707 ( \39050 , \39047 , \39049 );
not \U$38708 ( \39051 , \39050 );
not \U$38709 ( \39052 , \39000 );
and \U$38710 ( \39053 , \39051 , \39052 );
and \U$38711 ( \39054 , \39000 , \39050 );
nor \U$38712 ( \39055 , \39053 , \39054 );
not \U$38713 ( \39056 , \39055 );
or \U$38714 ( \39057 , \39046 , \39056 );
xor \U$38715 ( \39058 , \38956 , \38966 );
not \U$38716 ( \39059 , \12168 );
not \U$38717 ( \39060 , \38777 );
or \U$38718 ( \39061 , \39059 , \39060 );
and \U$38719 ( \39062 , \12278 , \16820 );
not \U$38720 ( \39063 , \12278 );
and \U$38721 ( \39064 , \39063 , \32817 );
or \U$38722 ( \39065 , \39062 , \39064 );
not \U$38723 ( \39066 , \39065 );
nand \U$38724 ( \39067 , \39066 , \12167 );
nand \U$38725 ( \39068 , \39061 , \39067 );
xor \U$38726 ( \39069 , \39058 , \39068 );
not \U$38727 ( \39070 , \14929 );
not \U$38728 ( \39071 , \38982 );
or \U$38729 ( \39072 , \39070 , \39071 );
not \U$38730 ( \39073 , RIbb2ddb0_53);
not \U$38731 ( \39074 , \32984 );
or \U$38732 ( \39075 , \39073 , \39074 );
nand \U$38733 ( \39076 , \13463 , \16856 );
nand \U$38734 ( \39077 , \39075 , \39076 );
nand \U$38735 ( \39078 , \39077 , \13467 );
nand \U$38736 ( \39079 , \39072 , \39078 );
and \U$38737 ( \39080 , \39069 , \39079 );
and \U$38738 ( \39081 , \39058 , \39068 );
or \U$38739 ( \39082 , \39080 , \39081 );
xor \U$38740 ( \39083 , \38967 , \38976 );
xor \U$38741 ( \39084 , \39083 , \38988 );
xor \U$38742 ( \39085 , \39082 , \39084 );
not \U$38743 ( \39086 , \12692 );
not \U$38744 ( \39087 , \38974 );
or \U$38745 ( \39088 , \39086 , \39087 );
not \U$38746 ( \39089 , RIbb2dea0_51);
not \U$38747 ( \39090 , \17768 );
or \U$38748 ( \39091 , \39089 , \39090 );
not \U$38749 ( \39092 , RIbb2dea0_51);
nand \U$38750 ( \39093 , \39092 , \16706 );
nand \U$38751 ( \39094 , \39091 , \39093 );
nand \U$38752 ( \39095 , \39094 , \12774 );
nand \U$38753 ( \39096 , \39088 , \39095 );
nor \U$38754 ( \39097 , \18929 , \38964 );
not \U$38755 ( \39098 , RIbb2df90_49);
not \U$38756 ( \39099 , \17745 );
or \U$38757 ( \39100 , \39098 , \39099 );
nand \U$38758 ( \39101 , \26129 , \12278 );
nand \U$38759 ( \39102 , \39100 , \39101 );
not \U$38760 ( \39103 , \39102 );
not \U$38761 ( \39104 , \12167 );
or \U$38762 ( \39105 , \39103 , \39104 );
or \U$38763 ( \39106 , \39065 , \12283 );
nand \U$38764 ( \39107 , \39105 , \39106 );
xor \U$38765 ( \39108 , \39097 , \39107 );
not \U$38766 ( \39109 , \12690 );
not \U$38767 ( \39110 , RIbb2dea0_51);
not \U$38768 ( \39111 , \17750 );
or \U$38769 ( \39112 , \39110 , \39111 );
not \U$38770 ( \39113 , RIbb2dea0_51);
nand \U$38771 ( \39114 , \39113 , \18920 );
nand \U$38772 ( \39115 , \39112 , \39114 );
not \U$38773 ( \39116 , \39115 );
or \U$38774 ( \39117 , \39109 , \39116 );
nand \U$38775 ( \39118 , \39094 , \12692 );
nand \U$38776 ( \39119 , \39117 , \39118 );
and \U$38777 ( \39120 , \39108 , \39119 );
and \U$38778 ( \39121 , \39097 , \39107 );
or \U$38779 ( \39122 , \39120 , \39121 );
xor \U$38780 ( \39123 , \39096 , \39122 );
not \U$38781 ( \39124 , \17397 );
not \U$38782 ( \39125 , \38863 );
or \U$38783 ( \39126 , \39124 , \39125 );
not \U$38784 ( \39127 , RIbb2dbd0_57);
not \U$38785 ( \39128 , \14528 );
or \U$38786 ( \39129 , \39127 , \39128 );
not \U$38787 ( \39130 , RIbb2dbd0_57);
nand \U$38788 ( \39131 , \39130 , \14527 );
nand \U$38789 ( \39132 , \39129 , \39131 );
nand \U$38790 ( \39133 , \39132 , \15746 );
nand \U$38791 ( \39134 , \39126 , \39133 );
and \U$38792 ( \39135 , \39123 , \39134 );
and \U$38793 ( \39136 , \39096 , \39122 );
or \U$38794 ( \39137 , \39135 , \39136 );
and \U$38795 ( \39138 , \39085 , \39137 );
and \U$38796 ( \39139 , \39082 , \39084 );
or \U$38797 ( \39140 , \39138 , \39139 );
not \U$38798 ( \39141 , \39140 );
not \U$38799 ( \39142 , \15182 );
not \U$38800 ( \39143 , \38872 );
or \U$38801 ( \39144 , \39142 , \39143 );
not \U$38802 ( \39145 , RIbb2dcc0_55);
not \U$38803 ( \39146 , \21665 );
or \U$38804 ( \39147 , \39145 , \39146 );
not \U$38805 ( \39148 , RIbb2dcc0_55);
nand \U$38806 ( \39149 , \39148 , \15756 );
nand \U$38807 ( \39150 , \39147 , \39149 );
nand \U$38808 ( \39151 , \39150 , \14613 );
nand \U$38809 ( \39152 , \39144 , \39151 );
not \U$38810 ( \39153 , \39152 );
not \U$38811 ( \39154 , \39153 );
not \U$38812 ( \39155 , \16271 );
and \U$38813 ( \39156 , RIbb2dae0_59, \15054 );
not \U$38814 ( \39157 , RIbb2dae0_59);
and \U$38815 ( \39158 , \39157 , \15055 );
or \U$38816 ( \39159 , \39156 , \39158 );
not \U$38817 ( \39160 , \39159 );
or \U$38818 ( \39161 , \39155 , \39160 );
nand \U$38819 ( \39162 , \38915 , \17470 );
nand \U$38820 ( \39163 , \39161 , \39162 );
not \U$38821 ( \39164 , \39163 );
not \U$38822 ( \39165 , \39164 );
or \U$38823 ( \39166 , \39154 , \39165 );
not \U$38824 ( \39167 , \18717 );
not \U$38825 ( \39168 , \25984 );
and \U$38826 ( \39169 , \39168 , RIbb2d9f0_61);
not \U$38827 ( \39170 , \39168 );
and \U$38828 ( \39171 , \39170 , \21449 );
or \U$38829 ( \39172 , \39169 , \39171 );
not \U$38830 ( \39173 , \39172 );
or \U$38831 ( \39174 , \39167 , \39173 );
nand \U$38832 ( \39175 , \38930 , \16533 );
nand \U$38833 ( \39176 , \39174 , \39175 );
nand \U$38834 ( \39177 , \39166 , \39176 );
nand \U$38835 ( \39178 , \39163 , \39152 );
nand \U$38836 ( \39179 , \39177 , \39178 );
not \U$38837 ( \39180 , \39179 );
xor \U$38838 ( \39181 , \38917 , \38932 );
xor \U$38839 ( \39182 , \39181 , \38943 );
not \U$38840 ( \39183 , \39182 );
or \U$38841 ( \39184 , \39180 , \39183 );
or \U$38842 ( \39185 , \39182 , \39179 );
xor \U$38843 ( \39186 , \39058 , \39068 );
xor \U$38844 ( \39187 , \39186 , \39079 );
or \U$38845 ( \39188 , RIbb2df18_50, RIbb2dea0_51);
nand \U$38846 ( \39189 , \39188 , \19064 );
and \U$38847 ( \39190 , RIbb2df18_50, RIbb2dea0_51);
nor \U$38848 ( \39191 , \39190 , \12278 );
and \U$38849 ( \39192 , \39189 , \39191 );
not \U$38850 ( \39193 , \12168 );
not \U$38851 ( \39194 , \39102 );
or \U$38852 ( \39195 , \39193 , \39194 );
or \U$38853 ( \39196 , \17506 , \12278 );
or \U$38854 ( \39197 , \18929 , RIbb2df90_49);
nand \U$38855 ( \39198 , \39196 , \39197 );
nand \U$38856 ( \39199 , \39198 , \12166 );
nand \U$38857 ( \39200 , \39195 , \39199 );
and \U$38858 ( \39201 , \39192 , \39200 );
not \U$38859 ( \39202 , \17562 );
not \U$38860 ( \39203 , RIbb2ddb0_53);
not \U$38861 ( \39204 , \35763 );
or \U$38862 ( \39205 , \39203 , \39204 );
nand \U$38863 ( \39206 , \19831 , \13463 );
nand \U$38864 ( \39207 , \39205 , \39206 );
not \U$38865 ( \39208 , \39207 );
or \U$38866 ( \39209 , \39202 , \39208 );
nand \U$38867 ( \39210 , \39077 , \14929 );
nand \U$38868 ( \39211 , \39209 , \39210 );
xor \U$38869 ( \39212 , \39201 , \39211 );
not \U$38870 ( \39213 , \15181 );
not \U$38871 ( \39214 , \39150 );
or \U$38872 ( \39215 , \39213 , \39214 );
and \U$38873 ( \39216 , RIbb2dcc0_55, \16577 );
not \U$38874 ( \39217 , RIbb2dcc0_55);
and \U$38875 ( \39218 , \39217 , \15825 );
or \U$38876 ( \39219 , \39216 , \39218 );
nand \U$38877 ( \39220 , \39219 , \14613 );
nand \U$38878 ( \39221 , \39215 , \39220 );
and \U$38879 ( \39222 , \39212 , \39221 );
and \U$38880 ( \39223 , \39201 , \39211 );
or \U$38881 ( \39224 , \39222 , \39223 );
xor \U$38882 ( \39225 , \39187 , \39224 );
not \U$38883 ( \39226 , RIbb2d888_64);
not \U$38884 ( \39227 , \38941 );
or \U$38885 ( \39228 , \39226 , \39227 );
and \U$38886 ( \39229 , \37646 , RIbb2d900_63);
not \U$38887 ( \39230 , \37646 );
and \U$38888 ( \39231 , \39230 , \17262 );
or \U$38889 ( \39232 , \39229 , \39231 );
nand \U$38890 ( \39233 , \39232 , \17275 );
nand \U$38891 ( \39234 , \39228 , \39233 );
and \U$38892 ( \39235 , \39225 , \39234 );
and \U$38893 ( \39236 , \39187 , \39224 );
or \U$38894 ( \39237 , \39235 , \39236 );
nand \U$38895 ( \39238 , \39185 , \39237 );
nand \U$38896 ( \39239 , \39184 , \39238 );
not \U$38897 ( \39240 , \39239 );
or \U$38898 ( \39241 , \39141 , \39240 );
or \U$38899 ( \39242 , \39239 , \39140 );
xor \U$38900 ( \39243 , \38857 , \38883 );
xor \U$38901 ( \39244 , \39243 , \38895 );
nand \U$38902 ( \39245 , \39242 , \39244 );
nand \U$38903 ( \39246 , \39241 , \39245 );
nand \U$38904 ( \39247 , \39057 , \39246 );
not \U$38905 ( \39248 , \39055 );
not \U$38906 ( \39249 , \39045 );
nand \U$38907 ( \39250 , \39248 , \39249 );
and \U$38908 ( \39251 , \39247 , \39250 );
nand \U$38909 ( \39252 , \39043 , \39251 );
xor \U$38910 ( \39253 , \39045 , \39246 );
xnor \U$38911 ( \39254 , \39253 , \39055 );
xor \U$38912 ( \39255 , \38906 , \38998 );
xnor \U$38913 ( \39256 , \39255 , \38946 );
xor \U$38914 ( \39257 , \38876 , \38867 );
and \U$38915 ( \39258 , \39257 , \38879 );
not \U$38916 ( \39259 , \39257 );
and \U$38917 ( \39260 , \39259 , \38880 );
nor \U$38918 ( \39261 , \39258 , \39260 );
xor \U$38919 ( \39262 , \39082 , \39084 );
xor \U$38920 ( \39263 , \39262 , \39137 );
and \U$38921 ( \39264 , \39261 , \39263 );
xor \U$38922 ( \39265 , \39096 , \39122 );
xor \U$38923 ( \39266 , \39265 , \39134 );
xor \U$38924 ( \39267 , \39192 , \39200 );
not \U$38925 ( \39268 , \12692 );
not \U$38926 ( \39269 , \39115 );
or \U$38927 ( \39270 , \39268 , \39269 );
and \U$38928 ( \39271 , RIbb2dea0_51, \16820 );
not \U$38929 ( \39272 , RIbb2dea0_51);
and \U$38930 ( \39273 , \39272 , \32817 );
or \U$38931 ( \39274 , \39271 , \39273 );
nand \U$38932 ( \39275 , \39274 , \12690 );
nand \U$38933 ( \39276 , \39270 , \39275 );
xor \U$38934 ( \39277 , \39267 , \39276 );
not \U$38935 ( \39278 , \14929 );
not \U$38936 ( \39279 , \39207 );
or \U$38937 ( \39280 , \39278 , \39279 );
not \U$38938 ( \39281 , RIbb2ddb0_53);
not \U$38939 ( \39282 , \34293 );
or \U$38940 ( \39283 , \39281 , \39282 );
nand \U$38941 ( \39284 , \16556 , \13463 );
nand \U$38942 ( \39285 , \39283 , \39284 );
nand \U$38943 ( \39286 , \39285 , \13467 );
nand \U$38944 ( \39287 , \39280 , \39286 );
and \U$38945 ( \39288 , \39277 , \39287 );
and \U$38946 ( \39289 , \39267 , \39276 );
or \U$38947 ( \39290 , \39288 , \39289 );
not \U$38948 ( \39291 , \16271 );
not \U$38949 ( \39292 , RIbb2dae0_59);
not \U$38950 ( \39293 , \35682 );
or \U$38951 ( \39294 , \39292 , \39293 );
not \U$38952 ( \39295 , RIbb2dae0_59);
nand \U$38953 ( \39296 , \39295 , \37489 );
nand \U$38954 ( \39297 , \39294 , \39296 );
not \U$38955 ( \39298 , \39297 );
or \U$38956 ( \39299 , \39291 , \39298 );
nand \U$38957 ( \39300 , \39159 , \16257 );
nand \U$38958 ( \39301 , \39299 , \39300 );
xor \U$38959 ( \39302 , \39290 , \39301 );
not \U$38960 ( \39303 , \26834 );
not \U$38961 ( \39304 , \39172 );
or \U$38962 ( \39305 , \39303 , \39304 );
not \U$38963 ( \39306 , RIbb2d9f0_61);
not \U$38964 ( \39307 , \13211 );
or \U$38965 ( \39308 , \39306 , \39307 );
nand \U$38966 ( \39309 , \13212 , \16254 );
nand \U$38967 ( \39310 , \39308 , \39309 );
nand \U$38968 ( \39311 , \39310 , \16541 );
nand \U$38969 ( \39312 , \39305 , \39311 );
and \U$38970 ( \39313 , \39302 , \39312 );
and \U$38971 ( \39314 , \39290 , \39301 );
or \U$38972 ( \39315 , \39313 , \39314 );
xor \U$38973 ( \39316 , \39266 , \39315 );
xor \U$38974 ( \39317 , \39097 , \39107 );
xor \U$38975 ( \39318 , \39317 , \39119 );
not \U$38976 ( \39319 , \15746 );
not \U$38977 ( \39320 , RIbb2dbd0_57);
not \U$38978 ( \39321 , \37560 );
or \U$38979 ( \39322 , \39320 , \39321 );
nand \U$38980 ( \39323 , \15032 , \15741 );
nand \U$38981 ( \39324 , \39322 , \39323 );
not \U$38982 ( \39325 , \39324 );
or \U$38983 ( \39326 , \39319 , \39325 );
nand \U$38984 ( \39327 , \39132 , \17100 );
nand \U$38985 ( \39328 , \39326 , \39327 );
xor \U$38986 ( \39329 , \39318 , \39328 );
not \U$38987 ( \39330 , RIbb2d888_64);
not \U$38988 ( \39331 , \39232 );
or \U$38989 ( \39332 , \39330 , \39331 );
not \U$38990 ( \39333 , RIbb2d900_63);
not \U$38991 ( \39334 , \12934 );
or \U$38992 ( \39335 , \39333 , \39334 );
nand \U$38993 ( \39336 , \37510 , \17262 );
nand \U$38994 ( \39337 , \39335 , \39336 );
nand \U$38995 ( \39338 , \39337 , \17275 );
nand \U$38996 ( \39339 , \39332 , \39338 );
and \U$38997 ( \39340 , \39329 , \39339 );
and \U$38998 ( \39341 , \39318 , \39328 );
or \U$38999 ( \39342 , \39340 , \39341 );
and \U$39000 ( \39343 , \39316 , \39342 );
and \U$39001 ( \39344 , \39266 , \39315 );
or \U$39002 ( \39345 , \39343 , \39344 );
not \U$39003 ( \39346 , \39261 );
not \U$39004 ( \39347 , \39263 );
nand \U$39005 ( \39348 , \39346 , \39347 );
and \U$39006 ( \39349 , \39345 , \39348 );
nor \U$39007 ( \39350 , \39264 , \39349 );
xor \U$39008 ( \39351 , \39256 , \39350 );
xor \U$39009 ( \39352 , \39140 , \39244 );
xnor \U$39010 ( \39353 , \39352 , \39239 );
and \U$39011 ( \39354 , \39351 , \39353 );
and \U$39012 ( \39355 , \39256 , \39350 );
or \U$39013 ( \39356 , \39354 , \39355 );
nand \U$39014 ( \39357 , \39254 , \39356 );
nand \U$39015 ( \39358 , \39252 , \39357 );
not \U$39016 ( \39359 , \39358 );
xor \U$39017 ( \39360 , \38550 , \38420 );
xnor \U$39018 ( \39361 , \39360 , \38500 );
not \U$39019 ( \39362 , \39361 );
xor \U$39020 ( \39363 , \38570 , \38573 );
xnor \U$39021 ( \39364 , \39363 , \38627 );
not \U$39022 ( \39365 , \39364 );
or \U$39023 ( \39366 , \39362 , \39365 );
xor \U$39024 ( \39367 , \39014 , \39016 );
and \U$39025 ( \39368 , \39367 , \39041 );
and \U$39026 ( \39369 , \39014 , \39016 );
or \U$39027 ( \39370 , \39368 , \39369 );
nand \U$39028 ( \39371 , \39366 , \39370 );
or \U$39029 ( \39372 , \39364 , \39361 );
nand \U$39030 ( \39373 , \39371 , \39372 );
not \U$39031 ( \39374 , \39373 );
not \U$39032 ( \39375 , \38567 );
not \U$39033 ( \39376 , \38629 );
or \U$39034 ( \39377 , \39375 , \39376 );
or \U$39035 ( \39378 , \38629 , \38567 );
nand \U$39036 ( \39379 , \39377 , \39378 );
and \U$39037 ( \39380 , \39379 , \38565 );
not \U$39038 ( \39381 , \39379 );
and \U$39039 ( \39382 , \39381 , \38564 );
nor \U$39040 ( \39383 , \39380 , \39382 );
nand \U$39041 ( \39384 , \39374 , \39383 );
not \U$39042 ( \39385 , \38758 );
not \U$39043 ( \39386 , \39385 );
not \U$39044 ( \39387 , \39005 );
or \U$39045 ( \39388 , \39386 , \39387 );
not \U$39046 ( \39389 , \38758 );
not \U$39047 ( \39390 , \39006 );
or \U$39048 ( \39391 , \39389 , \39390 );
nand \U$39049 ( \39392 , \39391 , \39042 );
nand \U$39050 ( \39393 , \39388 , \39392 );
not \U$39051 ( \39394 , \39393 );
xor \U$39052 ( \39395 , \39361 , \39370 );
xnor \U$39053 ( \39396 , \39395 , \39364 );
nand \U$39054 ( \39397 , \39394 , \39396 );
and \U$39055 ( \39398 , \39359 , \39384 , \39397 );
xor \U$39056 ( \39399 , \39256 , \39350 );
xor \U$39057 ( \39400 , \39399 , \39353 );
xor \U$39058 ( \39401 , \39179 , \39237 );
xnor \U$39059 ( \39402 , \39401 , \39182 );
xnor \U$39060 ( \39403 , \39176 , \39164 );
and \U$39061 ( \39404 , \39403 , \39152 );
not \U$39062 ( \39405 , \39403 );
and \U$39063 ( \39406 , \39405 , \39153 );
nor \U$39064 ( \39407 , \39404 , \39406 );
xor \U$39065 ( \39408 , \39187 , \39224 );
xor \U$39066 ( \39409 , \39408 , \39234 );
xor \U$39067 ( \39410 , \39407 , \39409 );
xor \U$39068 ( \39411 , \39201 , \39211 );
xor \U$39069 ( \39412 , \39411 , \39221 );
not \U$39070 ( \39413 , \16271 );
and \U$39071 ( \39414 , RIbb2dae0_59, \14528 );
not \U$39072 ( \39415 , RIbb2dae0_59);
and \U$39073 ( \39416 , \39415 , \14527 );
or \U$39074 ( \39417 , \39414 , \39416 );
not \U$39075 ( \39418 , \39417 );
or \U$39076 ( \39419 , \39413 , \39418 );
nand \U$39077 ( \39420 , \39297 , \16257 );
nand \U$39078 ( \39421 , \39419 , \39420 );
not \U$39079 ( \39422 , \39421 );
not \U$39080 ( \39423 , \39422 );
not \U$39081 ( \39424 , RIbb2d888_64);
not \U$39082 ( \39425 , \39337 );
or \U$39083 ( \39426 , \39424 , \39425 );
and \U$39084 ( \39427 , RIbb2d900_63, \39168 );
not \U$39085 ( \39428 , RIbb2d900_63);
and \U$39086 ( \39429 , \39428 , \12349 );
or \U$39087 ( \39430 , \39427 , \39429 );
nand \U$39088 ( \39431 , \39430 , \17275 );
nand \U$39089 ( \39432 , \39426 , \39431 );
not \U$39090 ( \39433 , \39432 );
not \U$39091 ( \39434 , \39433 );
or \U$39092 ( \39435 , \39423 , \39434 );
not \U$39093 ( \39436 , \26834 );
not \U$39094 ( \39437 , \39310 );
or \U$39095 ( \39438 , \39436 , \39437 );
not \U$39096 ( \39439 , RIbb2d9f0_61);
not \U$39097 ( \39440 , \13546 );
or \U$39098 ( \39441 , \39439 , \39440 );
nand \U$39099 ( \39442 , \15055 , \21449 );
nand \U$39100 ( \39443 , \39441 , \39442 );
nand \U$39101 ( \39444 , \39443 , \16541 );
nand \U$39102 ( \39445 , \39438 , \39444 );
nand \U$39103 ( \39446 , \39435 , \39445 );
nand \U$39104 ( \39447 , \39432 , \39421 );
nand \U$39105 ( \39448 , \39446 , \39447 );
or \U$39106 ( \39449 , \39412 , \39448 );
not \U$39107 ( \39450 , \14613 );
and \U$39108 ( \39451 , RIbb2dcc0_55, \32984 );
not \U$39109 ( \39452 , RIbb2dcc0_55);
and \U$39110 ( \39453 , \39452 , \18093 );
or \U$39111 ( \39454 , \39451 , \39453 );
not \U$39112 ( \39455 , \39454 );
or \U$39113 ( \39456 , \39450 , \39455 );
nand \U$39114 ( \39457 , \39219 , \15181 );
nand \U$39115 ( \39458 , \39456 , \39457 );
not \U$39116 ( \39459 , \39458 );
not \U$39117 ( \39460 , \17397 );
not \U$39118 ( \39461 , \39324 );
or \U$39119 ( \39462 , \39460 , \39461 );
and \U$39120 ( \39463 , RIbb2dbd0_57, \15756 );
not \U$39121 ( \39464 , RIbb2dbd0_57);
and \U$39122 ( \39465 , \39464 , \15755 );
nor \U$39123 ( \39466 , \39463 , \39465 );
nand \U$39124 ( \39467 , \39466 , \19101 );
nand \U$39125 ( \39468 , \39462 , \39467 );
not \U$39126 ( \39469 , \39468 );
or \U$39127 ( \39470 , \39459 , \39469 );
or \U$39128 ( \39471 , \39468 , \39458 );
and \U$39129 ( \39472 , \17506 , \12168 );
not \U$39130 ( \39473 , \12690 );
and \U$39131 ( \39474 , RIbb2dea0_51, \17745 );
not \U$39132 ( \39475 , RIbb2dea0_51);
and \U$39133 ( \39476 , \39475 , \28621 );
or \U$39134 ( \39477 , \39474 , \39476 );
not \U$39135 ( \39478 , \39477 );
or \U$39136 ( \39479 , \39473 , \39478 );
nand \U$39137 ( \39480 , \39274 , \12692 );
nand \U$39138 ( \39481 , \39479 , \39480 );
xor \U$39139 ( \39482 , \39472 , \39481 );
not \U$39140 ( \39483 , \13459 );
not \U$39141 ( \39484 , \39285 );
or \U$39142 ( \39485 , \39483 , \39484 );
not \U$39143 ( \39486 , RIbb2ddb0_53);
not \U$39144 ( \39487 , \17750 );
or \U$39145 ( \39488 , \39486 , \39487 );
nand \U$39146 ( \39489 , \16704 , \16210 );
nand \U$39147 ( \39490 , \39488 , \39489 );
nand \U$39148 ( \39491 , \39490 , \17562 );
nand \U$39149 ( \39492 , \39485 , \39491 );
and \U$39150 ( \39493 , \39482 , \39492 );
and \U$39151 ( \39494 , \39472 , \39481 );
or \U$39152 ( \39495 , \39493 , \39494 );
nand \U$39153 ( \39496 , \39471 , \39495 );
nand \U$39154 ( \39497 , \39470 , \39496 );
nand \U$39155 ( \39498 , \39449 , \39497 );
nand \U$39156 ( \39499 , \39448 , \39412 );
nand \U$39157 ( \39500 , \39498 , \39499 );
and \U$39158 ( \39501 , \39410 , \39500 );
and \U$39159 ( \39502 , \39407 , \39409 );
or \U$39160 ( \39503 , \39501 , \39502 );
not \U$39161 ( \39504 , \39503 );
xor \U$39162 ( \39505 , \39402 , \39504 );
not \U$39163 ( \39506 , \39345 );
and \U$39164 ( \39507 , \39261 , \39347 );
not \U$39165 ( \39508 , \39261 );
and \U$39166 ( \39509 , \39508 , \39263 );
nor \U$39167 ( \39510 , \39507 , \39509 );
not \U$39168 ( \39511 , \39510 );
and \U$39169 ( \39512 , \39506 , \39511 );
and \U$39170 ( \39513 , \39345 , \39510 );
nor \U$39171 ( \39514 , \39512 , \39513 );
and \U$39172 ( \39515 , \39505 , \39514 );
and \U$39173 ( \39516 , \39402 , \39504 );
or \U$39174 ( \39517 , \39515 , \39516 );
nand \U$39175 ( \39518 , \39400 , \39517 );
not \U$39176 ( \39519 , \39518 );
xor \U$39177 ( \39520 , \39266 , \39315 );
xor \U$39178 ( \39521 , \39520 , \39342 );
not \U$39179 ( \39522 , \39521 );
xor \U$39180 ( \39523 , \39290 , \39301 );
xor \U$39181 ( \39524 , \39523 , \39312 );
not \U$39182 ( \39525 , \39524 );
xor \U$39183 ( \39526 , \39318 , \39328 );
xor \U$39184 ( \39527 , \39526 , \39339 );
not \U$39185 ( \39528 , \39527 );
or \U$39186 ( \39529 , \39525 , \39528 );
not \U$39187 ( \39530 , \39524 );
not \U$39188 ( \39531 , \39530 );
not \U$39189 ( \39532 , \39527 );
not \U$39190 ( \39533 , \39532 );
or \U$39191 ( \39534 , \39531 , \39533 );
or \U$39192 ( \39535 , RIbb2de28_52, RIbb2ddb0_53);
nand \U$39193 ( \39536 , \39535 , \17506 );
and \U$39194 ( \39537 , RIbb2de28_52, RIbb2ddb0_53);
nor \U$39195 ( \39538 , \39537 , \21882 );
and \U$39196 ( \39539 , \39536 , \39538 );
not \U$39197 ( \39540 , \12691 );
not \U$39198 ( \39541 , \39477 );
or \U$39199 ( \39542 , \39540 , \39541 );
and \U$39200 ( \39543 , RIbb2dea0_51, \19064 );
not \U$39201 ( \39544 , RIbb2dea0_51);
and \U$39202 ( \39545 , \39544 , \20747 );
nor \U$39203 ( \39546 , \39543 , \39545 );
nand \U$39204 ( \39547 , \39546 , \12690 );
nand \U$39205 ( \39548 , \39542 , \39547 );
and \U$39206 ( \39549 , \39539 , \39548 );
not \U$39207 ( \39550 , \15182 );
not \U$39208 ( \39551 , \39454 );
or \U$39209 ( \39552 , \39550 , \39551 );
and \U$39210 ( \39553 , RIbb2dcc0_55, \35763 );
not \U$39211 ( \39554 , RIbb2dcc0_55);
and \U$39212 ( \39555 , \39554 , \36811 );
or \U$39213 ( \39556 , \39553 , \39555 );
nand \U$39214 ( \39557 , \39556 , \14613 );
nand \U$39215 ( \39558 , \39552 , \39557 );
xor \U$39216 ( \39559 , \39549 , \39558 );
not \U$39217 ( \39560 , \15738 );
not \U$39218 ( \39561 , \39466 );
or \U$39219 ( \39562 , \39560 , \39561 );
not \U$39220 ( \39563 , RIbb2dbd0_57);
not \U$39221 ( \39564 , \16577 );
or \U$39222 ( \39565 , \39563 , \39564 );
nand \U$39223 ( \39566 , \16576 , \14602 );
nand \U$39224 ( \39567 , \39565 , \39566 );
nand \U$39225 ( \39568 , \39567 , \16674 );
nand \U$39226 ( \39569 , \39562 , \39568 );
and \U$39227 ( \39570 , \39559 , \39569 );
and \U$39228 ( \39571 , \39549 , \39558 );
or \U$39229 ( \39572 , \39570 , \39571 );
not \U$39230 ( \39573 , \39572 );
xor \U$39231 ( \39574 , \39267 , \39276 );
xor \U$39232 ( \39575 , \39574 , \39287 );
not \U$39233 ( \39576 , \39575 );
nand \U$39234 ( \39577 , \39573 , \39576 );
not \U$39235 ( \39578 , \39577 );
xor \U$39236 ( \39579 , \39472 , \39481 );
xor \U$39237 ( \39580 , \39579 , \39492 );
not \U$39238 ( \39581 , \18717 );
not \U$39239 ( \39582 , RIbb2d9f0_61);
not \U$39240 ( \39583 , \35682 );
or \U$39241 ( \39584 , \39582 , \39583 );
nand \U$39242 ( \39585 , \37489 , \16254 );
nand \U$39243 ( \39586 , \39584 , \39585 );
not \U$39244 ( \39587 , \39586 );
or \U$39245 ( \39588 , \39581 , \39587 );
nand \U$39246 ( \39589 , \39443 , \16533 );
nand \U$39247 ( \39590 , \39588 , \39589 );
xor \U$39248 ( \39591 , \39580 , \39590 );
not \U$39249 ( \39592 , \17470 );
not \U$39250 ( \39593 , \39417 );
or \U$39251 ( \39594 , \39592 , \39593 );
xnor \U$39252 ( \39595 , RIbb2dae0_59, \37560 );
nand \U$39253 ( \39596 , \39595 , \16271 );
nand \U$39254 ( \39597 , \39594 , \39596 );
and \U$39255 ( \39598 , \39591 , \39597 );
and \U$39256 ( \39599 , \39580 , \39590 );
or \U$39257 ( \39600 , \39598 , \39599 );
not \U$39258 ( \39601 , \39600 );
or \U$39259 ( \39602 , \39578 , \39601 );
nand \U$39260 ( \39603 , \39572 , \39575 );
nand \U$39261 ( \39604 , \39602 , \39603 );
nand \U$39262 ( \39605 , \39534 , \39604 );
nand \U$39263 ( \39606 , \39529 , \39605 );
not \U$39264 ( \39607 , \39606 );
nand \U$39265 ( \39608 , \39522 , \39607 );
not \U$39266 ( \39609 , \39608 );
xor \U$39267 ( \39610 , \39407 , \39409 );
xor \U$39268 ( \39611 , \39610 , \39500 );
not \U$39269 ( \39612 , \39611 );
or \U$39270 ( \39613 , \39609 , \39612 );
nand \U$39271 ( \39614 , \39521 , \39606 );
nand \U$39272 ( \39615 , \39613 , \39614 );
not \U$39273 ( \39616 , \39615 );
xor \U$39274 ( \39617 , \39402 , \39504 );
xor \U$39275 ( \39618 , \39617 , \39514 );
nand \U$39276 ( \39619 , \39616 , \39618 );
not \U$39277 ( \39620 , \39619 );
xor \U$39278 ( \39621 , \39521 , \39607 );
xor \U$39279 ( \39622 , \39621 , \39611 );
xor \U$39280 ( \39623 , \39412 , \39497 );
xnor \U$39281 ( \39624 , \39623 , \39448 );
xor \U$39282 ( \39625 , \39495 , \39458 );
xnor \U$39283 ( \39626 , \39625 , \39468 );
xor \U$39284 ( \39627 , \39539 , \39548 );
not \U$39285 ( \39628 , \13459 );
not \U$39286 ( \39629 , \39490 );
or \U$39287 ( \39630 , \39628 , \39629 );
and \U$39288 ( \39631 , \12681 , \16820 );
not \U$39289 ( \39632 , \12681 );
and \U$39290 ( \39633 , \39632 , \16821 );
nor \U$39291 ( \39634 , \39631 , \39633 );
nand \U$39292 ( \39635 , \39634 , \17562 );
nand \U$39293 ( \39636 , \39630 , \39635 );
xor \U$39294 ( \39637 , \39627 , \39636 );
not \U$39295 ( \39638 , \15181 );
not \U$39296 ( \39639 , \39556 );
or \U$39297 ( \39640 , \39638 , \39639 );
not \U$39298 ( \39641 , RIbb2dcc0_55);
not \U$39299 ( \39642 , \17768 );
or \U$39300 ( \39643 , \39641 , \39642 );
not \U$39301 ( \39644 , RIbb2dcc0_55);
nand \U$39302 ( \39645 , \39644 , \16706 );
nand \U$39303 ( \39646 , \39643 , \39645 );
nand \U$39304 ( \39647 , \39646 , \14613 );
nand \U$39305 ( \39648 , \39640 , \39647 );
and \U$39306 ( \39649 , \39637 , \39648 );
and \U$39307 ( \39650 , \39627 , \39636 );
or \U$39308 ( \39651 , \39649 , \39650 );
not \U$39309 ( \39652 , \17275 );
not \U$39310 ( \39653 , RIbb2d900_63);
not \U$39311 ( \39654 , \15761 );
or \U$39312 ( \39655 , \39653 , \39654 );
nand \U$39313 ( \39656 , \13474 , \17270 );
nand \U$39314 ( \39657 , \39655 , \39656 );
not \U$39315 ( \39658 , \39657 );
or \U$39316 ( \39659 , \39652 , \39658 );
nand \U$39317 ( \39660 , \39430 , RIbb2d888_64);
nand \U$39318 ( \39661 , \39659 , \39660 );
xor \U$39319 ( \39662 , \39651 , \39661 );
xor \U$39320 ( \39663 , \39549 , \39558 );
xor \U$39321 ( \39664 , \39663 , \39569 );
and \U$39322 ( \39665 , \39662 , \39664 );
and \U$39323 ( \39666 , \39651 , \39661 );
or \U$39324 ( \39667 , \39665 , \39666 );
not \U$39325 ( \39668 , \39667 );
xor \U$39326 ( \39669 , \39626 , \39668 );
not \U$39327 ( \39670 , \39445 );
not \U$39328 ( \39671 , \39433 );
or \U$39329 ( \39672 , \39670 , \39671 );
or \U$39330 ( \39673 , \39433 , \39445 );
nand \U$39331 ( \39674 , \39672 , \39673 );
and \U$39332 ( \39675 , \39674 , \39422 );
not \U$39333 ( \39676 , \39674 );
and \U$39334 ( \39677 , \39676 , \39421 );
nor \U$39335 ( \39678 , \39675 , \39677 );
and \U$39336 ( \39679 , \39669 , \39678 );
and \U$39337 ( \39680 , \39626 , \39668 );
or \U$39338 ( \39681 , \39679 , \39680 );
xor \U$39339 ( \39682 , \39624 , \39681 );
and \U$39340 ( \39683 , \39527 , \39524 );
not \U$39341 ( \39684 , \39527 );
and \U$39342 ( \39685 , \39684 , \39530 );
nor \U$39343 ( \39686 , \39683 , \39685 );
not \U$39344 ( \39687 , \39604 );
and \U$39345 ( \39688 , \39686 , \39687 );
not \U$39346 ( \39689 , \39686 );
and \U$39347 ( \39690 , \39689 , \39604 );
nor \U$39348 ( \39691 , \39688 , \39690 );
and \U$39349 ( \39692 , \39682 , \39691 );
and \U$39350 ( \39693 , \39624 , \39681 );
or \U$39351 ( \39694 , \39692 , \39693 );
nand \U$39352 ( \39695 , \39622 , \39694 );
not \U$39353 ( \39696 , \39695 );
xor \U$39354 ( \39697 , \39624 , \39681 );
xor \U$39355 ( \39698 , \39697 , \39691 );
xor \U$39356 ( \39699 , \39626 , \39668 );
xor \U$39357 ( \39700 , \39699 , \39678 );
and \U$39358 ( \39701 , \39572 , \39575 );
not \U$39359 ( \39702 , \39572 );
and \U$39360 ( \39703 , \39702 , \39576 );
or \U$39361 ( \39704 , \39701 , \39703 );
xor \U$39362 ( \39705 , \39704 , \39600 );
nand \U$39363 ( \39706 , \39700 , \39705 );
not \U$39364 ( \39707 , \17100 );
not \U$39365 ( \39708 , \39567 );
or \U$39366 ( \39709 , \39707 , \39708 );
not \U$39367 ( \39710 , RIbb2dbd0_57);
not \U$39368 ( \39711 , \16748 );
or \U$39369 ( \39712 , \39710 , \39711 );
nand \U$39370 ( \39713 , \16751 , \15741 );
nand \U$39371 ( \39714 , \39712 , \39713 );
nand \U$39372 ( \39715 , \39714 , \16674 );
nand \U$39373 ( \39716 , \39709 , \39715 );
and \U$39374 ( \39717 , \17506 , \12692 );
not \U$39375 ( \39718 , \13459 );
not \U$39376 ( \39719 , \39634 );
or \U$39377 ( \39720 , \39718 , \39719 );
not \U$39378 ( \39721 , RIbb2ddb0_53);
not \U$39379 ( \39722 , \17745 );
or \U$39380 ( \39723 , \39721 , \39722 );
nand \U$39381 ( \39724 , \38079 , \13463 );
nand \U$39382 ( \39725 , \39723 , \39724 );
not \U$39383 ( \39726 , \39725 );
or \U$39384 ( \39727 , \39726 , \13466 );
nand \U$39385 ( \39728 , \39720 , \39727 );
xor \U$39386 ( \39729 , \39717 , \39728 );
not \U$39387 ( \39730 , \15181 );
not \U$39388 ( \39731 , \39646 );
or \U$39389 ( \39732 , \39730 , \39731 );
not \U$39390 ( \39733 , RIbb2dcc0_55);
not \U$39391 ( \39734 , \17750 );
or \U$39392 ( \39735 , \39733 , \39734 );
not \U$39393 ( \39736 , RIbb2dcc0_55);
nand \U$39394 ( \39737 , \39736 , \18920 );
nand \U$39395 ( \39738 , \39735 , \39737 );
nand \U$39396 ( \39739 , \39738 , \14613 );
nand \U$39397 ( \39740 , \39732 , \39739 );
and \U$39398 ( \39741 , \39729 , \39740 );
and \U$39399 ( \39742 , \39717 , \39728 );
or \U$39400 ( \39743 , \39741 , \39742 );
xor \U$39401 ( \39744 , \39716 , \39743 );
not \U$39402 ( \39745 , \16533 );
not \U$39403 ( \39746 , \39586 );
or \U$39404 ( \39747 , \39745 , \39746 );
not \U$39405 ( \39748 , RIbb2d9f0_61);
not \U$39406 ( \39749 , \14528 );
or \U$39407 ( \39750 , \39748 , \39749 );
nand \U$39408 ( \39751 , \14527 , \16254 );
nand \U$39409 ( \39752 , \39750 , \39751 );
nand \U$39410 ( \39753 , \39752 , \18717 );
nand \U$39411 ( \39754 , \39747 , \39753 );
and \U$39412 ( \39755 , \39744 , \39754 );
and \U$39413 ( \39756 , \39716 , \39743 );
or \U$39414 ( \39757 , \39755 , \39756 );
xor \U$39415 ( \39758 , \39580 , \39590 );
xor \U$39416 ( \39759 , \39758 , \39597 );
xor \U$39417 ( \39760 , \39757 , \39759 );
xor \U$39418 ( \39761 , \39627 , \39636 );
xor \U$39419 ( \39762 , \39761 , \39648 );
not \U$39420 ( \39763 , RIbb2d888_64);
not \U$39421 ( \39764 , \39657 );
or \U$39422 ( \39765 , \39763 , \39764 );
not \U$39423 ( \39766 , RIbb2d900_63);
not \U$39424 ( \39767 , \13546 );
or \U$39425 ( \39768 , \39766 , \39767 );
nand \U$39426 ( \39769 , \15055 , \33296 );
nand \U$39427 ( \39770 , \39768 , \39769 );
nand \U$39428 ( \39771 , \39770 , \17275 );
nand \U$39429 ( \39772 , \39765 , \39771 );
xor \U$39430 ( \39773 , \39762 , \39772 );
not \U$39431 ( \39774 , \17470 );
not \U$39432 ( \39775 , \39595 );
or \U$39433 ( \39776 , \39774 , \39775 );
and \U$39434 ( \39777 , RIbb2dae0_59, \16568 );
not \U$39435 ( \39778 , RIbb2dae0_59);
and \U$39436 ( \39779 , \39778 , \15755 );
nor \U$39437 ( \39780 , \39777 , \39779 );
nand \U$39438 ( \39781 , \39780 , \16271 );
nand \U$39439 ( \39782 , \39776 , \39781 );
and \U$39440 ( \39783 , \39773 , \39782 );
and \U$39441 ( \39784 , \39762 , \39772 );
or \U$39442 ( \39785 , \39783 , \39784 );
and \U$39443 ( \39786 , \39760 , \39785 );
and \U$39444 ( \39787 , \39757 , \39759 );
or \U$39445 ( \39788 , \39786 , \39787 );
and \U$39446 ( \39789 , \39706 , \39788 );
nor \U$39447 ( \39790 , \39700 , \39705 );
nor \U$39448 ( \39791 , \39789 , \39790 );
nor \U$39449 ( \39792 , \39698 , \39791 );
not \U$39450 ( \39793 , \39792 );
or \U$39451 ( \39794 , \39696 , \39793 );
or \U$39452 ( \39795 , \39622 , \39694 );
nand \U$39453 ( \39796 , \39794 , \39795 );
not \U$39454 ( \39797 , \39796 );
or \U$39455 ( \39798 , \39620 , \39797 );
not \U$39456 ( \39799 , \39618 );
nand \U$39457 ( \39800 , \39799 , \39615 );
nand \U$39458 ( \39801 , \39798 , \39800 );
not \U$39459 ( \39802 , \39801 );
or \U$39460 ( \39803 , \39519 , \39802 );
or \U$39461 ( \39804 , \39400 , \39517 );
nand \U$39462 ( \39805 , \39803 , \39804 );
and \U$39463 ( \39806 , \39398 , \39805 );
not \U$39464 ( \39807 , \39396 );
nand \U$39465 ( \39808 , \39807 , \39393 );
not \U$39466 ( \39809 , \39808 );
not \U$39467 ( \39810 , \39252 );
nor \U$39468 ( \39811 , \39254 , \39356 );
not \U$39469 ( \39812 , \39811 );
or \U$39470 ( \39813 , \39810 , \39812 );
or \U$39471 ( \39814 , \39043 , \39251 );
nand \U$39472 ( \39815 , \39813 , \39814 );
nand \U$39473 ( \39816 , \39815 , \39397 );
not \U$39474 ( \39817 , \39816 );
or \U$39475 ( \39818 , \39809 , \39817 );
buf \U$39476 ( \39819 , \39384 );
nand \U$39477 ( \39820 , \39818 , \39819 );
not \U$39478 ( \39821 , \39383 );
nand \U$39479 ( \39822 , \39821 , \39373 );
nand \U$39480 ( \39823 , \39820 , \39822 );
nor \U$39481 ( \39824 , \39806 , \39823 );
xor \U$39482 ( \39825 , \39757 , \39759 );
xor \U$39483 ( \39826 , \39825 , \39785 );
not \U$39484 ( \39827 , \39826 );
xor \U$39485 ( \39828 , \39651 , \39661 );
xor \U$39486 ( \39829 , \39828 , \39664 );
not \U$39487 ( \39830 , \39829 );
not \U$39488 ( \39831 , \16257 );
not \U$39489 ( \39832 , \39780 );
or \U$39490 ( \39833 , \39831 , \39832 );
and \U$39491 ( \39834 , RIbb2dae0_59, \15824 );
not \U$39492 ( \39835 , RIbb2dae0_59);
and \U$39493 ( \39836 , \39835 , \15825 );
or \U$39494 ( \39837 , \39834 , \39836 );
nand \U$39495 ( \39838 , \39837 , \16271 );
nand \U$39496 ( \39839 , \39833 , \39838 );
not \U$39497 ( \39840 , \15738 );
not \U$39498 ( \39841 , \39714 );
or \U$39499 ( \39842 , \39840 , \39841 );
and \U$39500 ( \39843 , RIbb2dbd0_57, \32993 );
not \U$39501 ( \39844 , RIbb2dbd0_57);
and \U$39502 ( \39845 , \39844 , \19831 );
or \U$39503 ( \39846 , \39843 , \39845 );
nand \U$39504 ( \39847 , \39846 , \16674 );
nand \U$39505 ( \39848 , \39842 , \39847 );
or \U$39506 ( \39849 , \39839 , \39848 );
or \U$39507 ( \39850 , RIbb2dd38_54, RIbb2dcc0_55);
nand \U$39508 ( \39851 , \39850 , \17506 );
and \U$39509 ( \39852 , RIbb2dd38_54, RIbb2dcc0_55);
nor \U$39510 ( \39853 , \39852 , \13463 );
and \U$39511 ( \39854 , \39851 , \39853 );
not \U$39512 ( \39855 , \13459 );
not \U$39513 ( \39856 , \39725 );
or \U$39514 ( \39857 , \39855 , \39856 );
or \U$39515 ( \39858 , \17506 , \16210 );
or \U$39516 ( \39859 , \19063 , RIbb2ddb0_53);
nand \U$39517 ( \39860 , \39858 , \39859 );
nand \U$39518 ( \39861 , \39860 , \13467 );
nand \U$39519 ( \39862 , \39857 , \39861 );
and \U$39520 ( \39863 , \39854 , \39862 );
nand \U$39521 ( \39864 , \39849 , \39863 );
nand \U$39522 ( \39865 , \39839 , \39848 );
nand \U$39523 ( \39866 , \39864 , \39865 );
xor \U$39524 ( \39867 , \39716 , \39743 );
xor \U$39525 ( \39868 , \39867 , \39754 );
xor \U$39526 ( \39869 , \39866 , \39868 );
xor \U$39527 ( \39870 , \39717 , \39728 );
xor \U$39528 ( \39871 , \39870 , \39740 );
not \U$39529 ( \39872 , \17275 );
not \U$39530 ( \39873 , RIbb2d900_63);
not \U$39531 ( \39874 , \35682 );
or \U$39532 ( \39875 , \39873 , \39874 );
nand \U$39533 ( \39876 , \35685 , \17262 );
nand \U$39534 ( \39877 , \39875 , \39876 );
not \U$39535 ( \39878 , \39877 );
or \U$39536 ( \39879 , \39872 , \39878 );
nand \U$39537 ( \39880 , \39770 , RIbb2d888_64);
nand \U$39538 ( \39881 , \39879 , \39880 );
xor \U$39539 ( \39882 , \39871 , \39881 );
not \U$39540 ( \39883 , \26834 );
not \U$39541 ( \39884 , \39752 );
or \U$39542 ( \39885 , \39883 , \39884 );
not \U$39543 ( \39886 , RIbb2d9f0_61);
not \U$39544 ( \39887 , \37559 );
not \U$39545 ( \39888 , \39887 );
or \U$39546 ( \39889 , \39886 , \39888 );
nand \U$39547 ( \39890 , \37559 , \16254 );
nand \U$39548 ( \39891 , \39889 , \39890 );
nand \U$39549 ( \39892 , \39891 , \16541 );
nand \U$39550 ( \39893 , \39885 , \39892 );
and \U$39551 ( \39894 , \39882 , \39893 );
and \U$39552 ( \39895 , \39871 , \39881 );
or \U$39553 ( \39896 , \39894 , \39895 );
and \U$39554 ( \39897 , \39869 , \39896 );
and \U$39555 ( \39898 , \39866 , \39868 );
or \U$39556 ( \39899 , \39897 , \39898 );
not \U$39557 ( \39900 , \39899 );
and \U$39558 ( \39901 , \39830 , \39900 );
or \U$39559 ( \39902 , \39827 , \39901 );
nand \U$39560 ( \39903 , \39899 , \39829 );
nand \U$39561 ( \39904 , \39902 , \39903 );
not \U$39562 ( \39905 , \39788 );
not \U$39563 ( \39906 , \39705 );
and \U$39564 ( \39907 , \39905 , \39906 );
and \U$39565 ( \39908 , \39788 , \39705 );
nor \U$39566 ( \39909 , \39907 , \39908 );
xor \U$39567 ( \39910 , \39909 , \39700 );
or \U$39568 ( \39911 , \39904 , \39910 );
not \U$39569 ( \39912 , \39911 );
xor \U$39570 ( \39913 , \39762 , \39772 );
xor \U$39571 ( \39914 , \39913 , \39782 );
not \U$39572 ( \39915 , \39914 );
xor \U$39573 ( \39916 , \39854 , \39862 );
not \U$39574 ( \39917 , \15181 );
not \U$39575 ( \39918 , \39738 );
or \U$39576 ( \39919 , \39917 , \39918 );
and \U$39577 ( \39920 , RIbb2dcc0_55, \16818 );
not \U$39578 ( \39921 , RIbb2dcc0_55);
and \U$39579 ( \39922 , \39921 , \16820 );
nor \U$39580 ( \39923 , \39920 , \39922 );
nand \U$39581 ( \39924 , \39923 , \14613 );
nand \U$39582 ( \39925 , \39919 , \39924 );
xor \U$39583 ( \39926 , \39916 , \39925 );
not \U$39584 ( \39927 , \15738 );
not \U$39585 ( \39928 , \39846 );
or \U$39586 ( \39929 , \39927 , \39928 );
not \U$39587 ( \39930 , RIbb2dbd0_57);
not \U$39588 ( \39931 , \16555 );
or \U$39589 ( \39932 , \39930 , \39931 );
nand \U$39590 ( \39933 , \16706 , \15741 );
nand \U$39591 ( \39934 , \39932 , \39933 );
nand \U$39592 ( \39935 , \39934 , \19101 );
nand \U$39593 ( \39936 , \39929 , \39935 );
and \U$39594 ( \39937 , \39926 , \39936 );
and \U$39595 ( \39938 , \39916 , \39925 );
or \U$39596 ( \39939 , \39937 , \39938 );
not \U$39597 ( \39940 , \39939 );
xor \U$39598 ( \39941 , \39863 , \39848 );
xnor \U$39599 ( \39942 , \39941 , \39839 );
nand \U$39600 ( \39943 , \39940 , \39942 );
not \U$39601 ( \39944 , \39943 );
not \U$39602 ( \39945 , \16533 );
not \U$39603 ( \39946 , \39891 );
or \U$39604 ( \39947 , \39945 , \39946 );
not \U$39605 ( \39948 , RIbb2d9f0_61);
not \U$39606 ( \39949 , \21665 );
or \U$39607 ( \39950 , \39948 , \39949 );
nand \U$39608 ( \39951 , \15756 , \19746 );
nand \U$39609 ( \39952 , \39950 , \39951 );
nand \U$39610 ( \39953 , \39952 , \16541 );
nand \U$39611 ( \39954 , \39947 , \39953 );
not \U$39612 ( \39955 , \16257 );
not \U$39613 ( \39956 , \39837 );
or \U$39614 ( \39957 , \39955 , \39956 );
and \U$39615 ( \39958 , RIbb2dae0_59, \32984 );
not \U$39616 ( \39959 , RIbb2dae0_59);
and \U$39617 ( \39960 , \39959 , \16856 );
or \U$39618 ( \39961 , \39958 , \39960 );
nand \U$39619 ( \39962 , \39961 , \16271 );
nand \U$39620 ( \39963 , \39957 , \39962 );
or \U$39621 ( \39964 , \39954 , \39963 );
and \U$39622 ( \39965 , \17506 , \13459 );
not \U$39623 ( \39966 , \14613 );
and \U$39624 ( \39967 , RIbb2dcc0_55, \19841 );
not \U$39625 ( \39968 , RIbb2dcc0_55);
and \U$39626 ( \39969 , \39968 , \17745 );
nor \U$39627 ( \39970 , \39967 , \39969 );
not \U$39628 ( \39971 , \39970 );
or \U$39629 ( \39972 , \39966 , \39971 );
nand \U$39630 ( \39973 , \39923 , \15181 );
nand \U$39631 ( \39974 , \39972 , \39973 );
xor \U$39632 ( \39975 , \39965 , \39974 );
not \U$39633 ( \39976 , \15746 );
and \U$39634 ( \39977 , \17411 , \17750 );
not \U$39635 ( \39978 , \17411 );
and \U$39636 ( \39979 , \39978 , \16704 );
nor \U$39637 ( \39980 , \39977 , \39979 );
not \U$39638 ( \39981 , \39980 );
or \U$39639 ( \39982 , \39976 , \39981 );
nand \U$39640 ( \39983 , \39934 , \15738 );
nand \U$39641 ( \39984 , \39982 , \39983 );
and \U$39642 ( \39985 , \39975 , \39984 );
and \U$39643 ( \39986 , \39965 , \39974 );
or \U$39644 ( \39987 , \39985 , \39986 );
nand \U$39645 ( \39988 , \39964 , \39987 );
nand \U$39646 ( \39989 , \39954 , \39963 );
nand \U$39647 ( \39990 , \39988 , \39989 );
not \U$39648 ( \39991 , \39990 );
or \U$39649 ( \39992 , \39944 , \39991 );
not \U$39650 ( \39993 , \39942 );
nand \U$39651 ( \39994 , \39993 , \39939 );
nand \U$39652 ( \39995 , \39992 , \39994 );
not \U$39653 ( \39996 , \39995 );
nand \U$39654 ( \39997 , \39915 , \39996 );
not \U$39655 ( \39998 , \39997 );
xor \U$39656 ( \39999 , \39866 , \39868 );
xor \U$39657 ( \40000 , \39999 , \39896 );
not \U$39658 ( \40001 , \40000 );
or \U$39659 ( \40002 , \39998 , \40001 );
nand \U$39660 ( \40003 , \39914 , \39995 );
nand \U$39661 ( \40004 , \40002 , \40003 );
not \U$39662 ( \40005 , \40004 );
xor \U$39663 ( \40006 , \39830 , \39900 );
and \U$39664 ( \40007 , \40006 , \39827 );
not \U$39665 ( \40008 , \40006 );
and \U$39666 ( \40009 , \40008 , \39826 );
nor \U$39667 ( \40010 , \40007 , \40009 );
nand \U$39668 ( \40011 , \40005 , \40010 );
not \U$39669 ( \40012 , \40011 );
not \U$39670 ( \40013 , \15181 );
not \U$39671 ( \40014 , \39970 );
or \U$39672 ( \40015 , \40013 , \40014 );
and \U$39673 ( \40016 , RIbb2dcc0_55, \17506 );
not \U$39674 ( \40017 , RIbb2dcc0_55);
and \U$39675 ( \40018 , \40017 , \20747 );
nor \U$39676 ( \40019 , \40016 , \40018 );
nand \U$39677 ( \40020 , \40019 , \14612 );
nand \U$39678 ( \40021 , \40015 , \40020 );
or \U$39679 ( \40022 , RIbb2dc48_56, RIbb2dbd0_57);
nand \U$39680 ( \40023 , \40022 , \17506 );
and \U$39681 ( \40024 , RIbb2dc48_56, RIbb2dbd0_57);
nor \U$39682 ( \40025 , \40024 , \18174 );
and \U$39683 ( \40026 , \40023 , \40025 );
and \U$39684 ( \40027 , \40021 , \40026 );
not \U$39685 ( \40028 , \16257 );
not \U$39686 ( \40029 , \39961 );
or \U$39687 ( \40030 , \40028 , \40029 );
and \U$39688 ( \40031 , RIbb2dae0_59, \37964 );
not \U$39689 ( \40032 , RIbb2dae0_59);
and \U$39690 ( \40033 , \40032 , \36811 );
or \U$39691 ( \40034 , \40031 , \40033 );
nand \U$39692 ( \40035 , \40034 , \16271 );
nand \U$39693 ( \40036 , \40030 , \40035 );
xor \U$39694 ( \40037 , \40027 , \40036 );
not \U$39695 ( \40038 , \16533 );
not \U$39696 ( \40039 , \39952 );
or \U$39697 ( \40040 , \40038 , \40039 );
and \U$39698 ( \40041 , \16254 , \15824 );
not \U$39699 ( \40042 , \16254 );
and \U$39700 ( \40043 , \40042 , \16575 );
nor \U$39701 ( \40044 , \40041 , \40043 );
nand \U$39702 ( \40045 , \40044 , \16541 );
nand \U$39703 ( \40046 , \40040 , \40045 );
xnor \U$39704 ( \40047 , \40037 , \40046 );
not \U$39705 ( \40048 , \40047 );
not \U$39706 ( \40049 , \40048 );
not \U$39707 ( \40050 , RIbb2d888_64);
not \U$39708 ( \40051 , RIbb2d900_63);
not \U$39709 ( \40052 , \39887 );
or \U$39710 ( \40053 , \40051 , \40052 );
nand \U$39711 ( \40054 , \37559 , \17262 );
nand \U$39712 ( \40055 , \40053 , \40054 );
not \U$39713 ( \40056 , \40055 );
or \U$39714 ( \40057 , \40050 , \40056 );
xor \U$39715 ( \40058 , RIbb2d900_63, \23098 );
nand \U$39716 ( \40059 , \40058 , \17275 );
nand \U$39717 ( \40060 , \40057 , \40059 );
not \U$39718 ( \40061 , \16257 );
not \U$39719 ( \40062 , \40034 );
or \U$39720 ( \40063 , \40061 , \40062 );
not \U$39721 ( \40064 , \16555 );
not \U$39722 ( \40065 , RIbb2dae0_59);
or \U$39723 ( \40066 , \40064 , \40065 );
not \U$39724 ( \40067 , RIbb2dae0_59);
nand \U$39725 ( \40068 , \40067 , \16706 );
nand \U$39726 ( \40069 , \40066 , \40068 );
nand \U$39727 ( \40070 , \40069 , \16271 );
nand \U$39728 ( \40071 , \40063 , \40070 );
or \U$39729 ( \40072 , \40060 , \40071 );
not \U$39730 ( \40073 , \40072 );
and \U$39731 ( \40074 , \17506 , \15181 );
not \U$39732 ( \40075 , \15738 );
and \U$39733 ( \40076 , RIbb2dbd0_57, \17529 );
not \U$39734 ( \40077 , RIbb2dbd0_57);
and \U$39735 ( \40078 , \40077 , \35466 );
nor \U$39736 ( \40079 , \40076 , \40078 );
not \U$39737 ( \40080 , \40079 );
or \U$39738 ( \40081 , \40075 , \40080 );
not \U$39739 ( \40082 , RIbb2dbd0_57);
not \U$39740 ( \40083 , \17519 );
or \U$39741 ( \40084 , \40082 , \40083 );
nand \U$39742 ( \40085 , \17518 , \17411 );
nand \U$39743 ( \40086 , \40084 , \40085 );
nand \U$39744 ( \40087 , \40086 , \15746 );
nand \U$39745 ( \40088 , \40081 , \40087 );
xor \U$39746 ( \40089 , \40074 , \40088 );
not \U$39747 ( \40090 , \16256 );
not \U$39748 ( \40091 , \40069 );
or \U$39749 ( \40092 , \40090 , \40091 );
not \U$39750 ( \40093 , RIbb2dae0_59);
not \U$39751 ( \40094 , \17750 );
or \U$39752 ( \40095 , \40093 , \40094 );
not \U$39753 ( \40096 , RIbb2dae0_59);
nand \U$39754 ( \40097 , \40096 , \18920 );
nand \U$39755 ( \40098 , \40095 , \40097 );
nand \U$39756 ( \40099 , \16270 , \40098 );
nand \U$39757 ( \40100 , \40092 , \40099 );
and \U$39758 ( \40101 , \40089 , \40100 );
and \U$39759 ( \40102 , \40074 , \40088 );
or \U$39760 ( \40103 , \40101 , \40102 );
not \U$39761 ( \40104 , \40103 );
or \U$39762 ( \40105 , \40073 , \40104 );
nand \U$39763 ( \40106 , \40060 , \40071 );
nand \U$39764 ( \40107 , \40105 , \40106 );
not \U$39765 ( \40108 , \40107 );
nand \U$39766 ( \40109 , \40049 , \40108 );
not \U$39767 ( \40110 , \40109 );
xor \U$39768 ( \40111 , \39965 , \39974 );
xor \U$39769 ( \40112 , \40111 , \39984 );
not \U$39770 ( \40113 , RIbb2d888_64);
not \U$39771 ( \40114 , RIbb2d900_63);
not \U$39772 ( \40115 , \14528 );
or \U$39773 ( \40116 , \40114 , \40115 );
nand \U$39774 ( \40117 , \14527 , \17270 );
nand \U$39775 ( \40118 , \40116 , \40117 );
not \U$39776 ( \40119 , \40118 );
or \U$39777 ( \40120 , \40113 , \40119 );
nand \U$39778 ( \40121 , \40055 , \17275 );
nand \U$39779 ( \40122 , \40120 , \40121 );
xor \U$39780 ( \40123 , \40112 , \40122 );
not \U$39781 ( \40124 , \15738 );
not \U$39782 ( \40125 , \39980 );
or \U$39783 ( \40126 , \40124 , \40125 );
nand \U$39784 ( \40127 , \40079 , \16674 );
nand \U$39785 ( \40128 , \40126 , \40127 );
not \U$39786 ( \40129 , \40128 );
not \U$39787 ( \40130 , \16533 );
not \U$39788 ( \40131 , \40044 );
or \U$39789 ( \40132 , \40130 , \40131 );
not \U$39790 ( \40133 , RIbb2d9f0_61);
not \U$39791 ( \40134 , \16748 );
or \U$39792 ( \40135 , \40133 , \40134 );
not \U$39793 ( \40136 , \16747 );
nand \U$39794 ( \40137 , \40136 , \16254 );
nand \U$39795 ( \40138 , \40135 , \40137 );
nand \U$39796 ( \40139 , \40138 , \16541 );
nand \U$39797 ( \40140 , \40132 , \40139 );
not \U$39798 ( \40141 , \40140 );
or \U$39799 ( \40142 , \40129 , \40141 );
or \U$39800 ( \40143 , \40140 , \40128 );
xnor \U$39801 ( \40144 , \40021 , \40026 );
not \U$39802 ( \40145 , \40144 );
nand \U$39803 ( \40146 , \40143 , \40145 );
nand \U$39804 ( \40147 , \40142 , \40146 );
xor \U$39805 ( \40148 , \40123 , \40147 );
not \U$39806 ( \40149 , \40148 );
or \U$39807 ( \40150 , \40110 , \40149 );
nand \U$39808 ( \40151 , \40107 , \40048 );
nand \U$39809 ( \40152 , \40150 , \40151 );
not \U$39810 ( \40153 , \40152 );
xor \U$39811 ( \40154 , \39963 , \39987 );
xnor \U$39812 ( \40155 , \40154 , \39954 );
or \U$39813 ( \40156 , \40122 , \40112 );
nand \U$39814 ( \40157 , \40156 , \40147 );
nand \U$39815 ( \40158 , \40122 , \40112 );
and \U$39816 ( \40159 , \40157 , \40158 );
xor \U$39817 ( \40160 , \40155 , \40159 );
xor \U$39818 ( \40161 , \39916 , \39925 );
xor \U$39819 ( \40162 , \40161 , \39936 );
not \U$39820 ( \40163 , \17275 );
not \U$39821 ( \40164 , \40118 );
or \U$39822 ( \40165 , \40163 , \40164 );
nand \U$39823 ( \40166 , \39877 , RIbb2d888_64);
nand \U$39824 ( \40167 , \40165 , \40166 );
xor \U$39825 ( \40168 , \40162 , \40167 );
or \U$39826 ( \40169 , \40036 , \40046 );
nand \U$39827 ( \40170 , \40169 , \40027 );
nand \U$39828 ( \40171 , \40046 , \40036 );
nand \U$39829 ( \40172 , \40170 , \40171 );
xnor \U$39830 ( \40173 , \40168 , \40172 );
xor \U$39831 ( \40174 , \40160 , \40173 );
nand \U$39832 ( \40175 , \40153 , \40174 );
not \U$39833 ( \40176 , \40175 );
not \U$39834 ( \40177 , \15738 );
nor \U$39835 ( \40178 , \40177 , \20747 );
and \U$39836 ( \40179 , RIbb2dae0_59, \26050 );
not \U$39837 ( \40180 , RIbb2dae0_59);
and \U$39838 ( \40181 , \40180 , \17529 );
or \U$39839 ( \40182 , \40179 , \40181 );
not \U$39840 ( \40183 , \40182 );
not \U$39841 ( \40184 , \16256 );
or \U$39842 ( \40185 , \40183 , \40184 );
and \U$39843 ( \40186 , RIbb2dae0_59, \35598 );
not \U$39844 ( \40187 , RIbb2dae0_59);
and \U$39845 ( \40188 , \40187 , \17745 );
nor \U$39846 ( \40189 , \40186 , \40188 );
nand \U$39847 ( \40190 , \16270 , \40189 );
nand \U$39848 ( \40191 , \40185 , \40190 );
xor \U$39849 ( \40192 , \40178 , \40191 );
not \U$39850 ( \40193 , \16541 );
not \U$39851 ( \40194 , RIbb2d9f0_61);
not \U$39852 ( \40195 , \17750 );
or \U$39853 ( \40196 , \40194 , \40195 );
not \U$39854 ( \40197 , RIbb2d9f0_61);
nand \U$39855 ( \40198 , \40197 , \18923 );
nand \U$39856 ( \40199 , \40196 , \40198 );
not \U$39857 ( \40200 , \40199 );
or \U$39858 ( \40201 , \40193 , \40200 );
not \U$39859 ( \40202 , RIbb2d9f0_61);
not \U$39860 ( \40203 , \17768 );
or \U$39861 ( \40204 , \40202 , \40203 );
nand \U$39862 ( \40205 , \16706 , \16254 );
nand \U$39863 ( \40206 , \40204 , \40205 );
nand \U$39864 ( \40207 , \40206 , \16533 );
nand \U$39865 ( \40208 , \40201 , \40207 );
and \U$39866 ( \40209 , \40192 , \40208 );
and \U$39867 ( \40210 , \40178 , \40191 );
or \U$39868 ( \40211 , \40209 , \40210 );
not \U$39869 ( \40212 , \40211 );
not \U$39870 ( \40213 , \17274 );
and \U$39871 ( \40214 , RIbb2d900_63, \16751 );
not \U$39872 ( \40215 , RIbb2d900_63);
and \U$39873 ( \40216 , \40215 , \16748 );
nor \U$39874 ( \40217 , \40214 , \40216 );
not \U$39875 ( \40218 , \40217 );
or \U$39876 ( \40219 , \40213 , \40218 );
not \U$39877 ( \40220 , RIbb2d900_63);
not \U$39878 ( \40221 , \20716 );
or \U$39879 ( \40222 , \40220 , \40221 );
nand \U$39880 ( \40223 , \16575 , \17262 );
nand \U$39881 ( \40224 , \40222 , \40223 );
nand \U$39882 ( \40225 , \40224 , RIbb2d888_64);
nand \U$39883 ( \40226 , \40219 , \40225 );
not \U$39884 ( \40227 , \40226 );
nand \U$39885 ( \40228 , \40212 , \40227 );
not \U$39886 ( \40229 , \40228 );
not \U$39887 ( \40230 , \16256 );
not \U$39888 ( \40231 , \40098 );
or \U$39889 ( \40232 , \40230 , \40231 );
nand \U$39890 ( \40233 , \40182 , \16270 );
nand \U$39891 ( \40234 , \40232 , \40233 );
or \U$39892 ( \40235 , RIbb2db58_58, RIbb2dae0_59);
nand \U$39893 ( \40236 , \40235 , \17506 );
and \U$39894 ( \40237 , RIbb2db58_58, RIbb2dae0_59);
nor \U$39895 ( \40238 , \40237 , \17097 );
and \U$39896 ( \40239 , \40236 , \40238 );
not \U$39897 ( \40240 , \15738 );
not \U$39898 ( \40241 , \40086 );
or \U$39899 ( \40242 , \40240 , \40241 );
or \U$39900 ( \40243 , \17506 , \14602 );
or \U$39901 ( \40244 , \19063 , RIbb2dbd0_57);
nand \U$39902 ( \40245 , \40243 , \40244 );
nand \U$39903 ( \40246 , \40245 , \15746 );
nand \U$39904 ( \40247 , \40242 , \40246 );
xor \U$39905 ( \40248 , \40239 , \40247 );
xor \U$39906 ( \40249 , \40234 , \40248 );
not \U$39907 ( \40250 , \16533 );
and \U$39908 ( \40251 , RIbb2d9f0_61, \19831 );
not \U$39909 ( \40252 , RIbb2d9f0_61);
and \U$39910 ( \40253 , \40252 , \27577 );
nor \U$39911 ( \40254 , \40251 , \40253 );
not \U$39912 ( \40255 , \40254 );
or \U$39913 ( \40256 , \40250 , \40255 );
nand \U$39914 ( \40257 , \40206 , \16541 );
nand \U$39915 ( \40258 , \40256 , \40257 );
xor \U$39916 ( \40259 , \40249 , \40258 );
not \U$39917 ( \40260 , \40259 );
or \U$39918 ( \40261 , \40229 , \40260 );
nand \U$39919 ( \40262 , \40211 , \40226 );
nand \U$39920 ( \40263 , \40261 , \40262 );
xor \U$39921 ( \40264 , \40074 , \40088 );
xor \U$39922 ( \40265 , \40264 , \40100 );
xor \U$39923 ( \40266 , \40234 , \40248 );
and \U$39924 ( \40267 , \40266 , \40258 );
and \U$39925 ( \40268 , \40234 , \40248 );
or \U$39926 ( \40269 , \40267 , \40268 );
xor \U$39927 ( \40270 , \40265 , \40269 );
nand \U$39928 ( \40271 , \40247 , \40239 );
not \U$39929 ( \40272 , \16541 );
not \U$39930 ( \40273 , \40254 );
or \U$39931 ( \40274 , \40272 , \40273 );
nand \U$39932 ( \40275 , \40138 , \16533 );
nand \U$39933 ( \40276 , \40274 , \40275 );
xor \U$39934 ( \40277 , \40271 , \40276 );
not \U$39935 ( \40278 , RIbb2d888_64);
not \U$39936 ( \40279 , \40058 );
or \U$39937 ( \40280 , \40278 , \40279 );
nand \U$39938 ( \40281 , \40224 , \17274 );
nand \U$39939 ( \40282 , \40280 , \40281 );
xnor \U$39940 ( \40283 , \40277 , \40282 );
xor \U$39941 ( \40284 , \40270 , \40283 );
xor \U$39942 ( \40285 , \40263 , \40284 );
not \U$39943 ( \40286 , RIbb2d888_64);
not \U$39944 ( \40287 , \40217 );
or \U$39945 ( \40288 , \40286 , \40287 );
not \U$39946 ( \40289 , RIbb2d900_63);
not \U$39947 ( \40290 , \27577 );
or \U$39948 ( \40291 , \40289 , \40290 );
nand \U$39949 ( \40292 , \16829 , \19721 );
nand \U$39950 ( \40293 , \40291 , \40292 );
nand \U$39951 ( \40294 , \40293 , \17273 );
nand \U$39952 ( \40295 , \40288 , \40294 );
or \U$39953 ( \40296 , RIbb2da68_60, RIbb2d9f0_61);
nand \U$39954 ( \40297 , \40296 , \19064 );
and \U$39955 ( \40298 , RIbb2da68_60, RIbb2d9f0_61);
nor \U$39956 ( \40299 , \40298 , \17024 );
and \U$39957 ( \40300 , \40297 , \40299 );
not \U$39958 ( \40301 , \16256 );
not \U$39959 ( \40302 , \40189 );
or \U$39960 ( \40303 , \40301 , \40302 );
and \U$39961 ( \40304 , RIbb2dae0_59, \17506 );
not \U$39962 ( \40305 , RIbb2dae0_59);
and \U$39963 ( \40306 , \40305 , \20747 );
nor \U$39964 ( \40307 , \40304 , \40306 );
nand \U$39965 ( \40308 , \40307 , \16270 );
nand \U$39966 ( \40309 , \40303 , \40308 );
and \U$39967 ( \40310 , \40300 , \40309 );
nor \U$39968 ( \40311 , \40295 , \40310 );
xor \U$39969 ( \40312 , \40178 , \40191 );
xor \U$39970 ( \40313 , \40312 , \40208 );
not \U$39971 ( \40314 , \40313 );
or \U$39972 ( \40315 , \40311 , \40314 );
nand \U$39973 ( \40316 , \40295 , \40310 );
nand \U$39974 ( \40317 , \40315 , \40316 );
not \U$39975 ( \40318 , \40317 );
xor \U$39976 ( \40319 , \40227 , \40211 );
xor \U$39977 ( \40320 , \40259 , \40319 );
nand \U$39978 ( \40321 , \40318 , \40320 );
or \U$39979 ( \40322 , \18929 , \21654 );
not \U$39980 ( \40323 , \16532 );
not \U$39981 ( \40324 , RIbb2d9f0_61);
not \U$39982 ( \40325 , \16819 );
or \U$39983 ( \40326 , \40324 , \40325 );
nand \U$39984 ( \40327 , \17529 , \19746 );
nand \U$39985 ( \40328 , \40326 , \40327 );
not \U$39986 ( \40329 , \40328 );
or \U$39987 ( \40330 , \40323 , \40329 );
not \U$39988 ( \40331 , RIbb2d9f0_61);
not \U$39989 ( \40332 , \20552 );
or \U$39990 ( \40333 , \40331 , \40332 );
nand \U$39991 ( \40334 , \26129 , \19746 );
nand \U$39992 ( \40335 , \40333 , \40334 );
nand \U$39993 ( \40336 , \40335 , \16540 );
nand \U$39994 ( \40337 , \40330 , \40336 );
xor \U$39995 ( \40338 , \40322 , \40337 );
not \U$39996 ( \40339 , \17273 );
and \U$39997 ( \40340 , RIbb2d900_63, \17751 );
not \U$39998 ( \40341 , RIbb2d900_63);
and \U$39999 ( \40342 , \40341 , \18924 );
nor \U$40000 ( \40343 , \40340 , \40342 );
not \U$40001 ( \40344 , \40343 );
or \U$40002 ( \40345 , \40339 , \40344 );
xor \U$40003 ( \40346 , RIbb2d900_63, \16706 );
nand \U$40004 ( \40347 , \40346 , RIbb2d888_64);
nand \U$40005 ( \40348 , \40345 , \40347 );
xor \U$40006 ( \40349 , \40338 , \40348 );
or \U$40007 ( \40350 , RIbb2d978_62, RIbb2d900_63);
nand \U$40008 ( \40351 , \40350 , \17506 );
and \U$40009 ( \40352 , RIbb2d978_62, RIbb2d900_63);
nor \U$40010 ( \40353 , \40352 , \16537 );
nand \U$40011 ( \40354 , \40351 , \40353 );
not \U$40012 ( \40355 , \40354 );
not \U$40013 ( \40356 , \16532 );
not \U$40014 ( \40357 , \40335 );
or \U$40015 ( \40358 , \40356 , \40357 );
or \U$40016 ( \40359 , \19064 , \16254 );
or \U$40017 ( \40360 , \19063 , RIbb2d9f0_61);
nand \U$40018 ( \40361 , \40359 , \40360 );
nand \U$40019 ( \40362 , \40361 , \16540 );
nand \U$40020 ( \40363 , \40358 , \40362 );
nand \U$40021 ( \40364 , \40355 , \40363 );
nand \U$40022 ( \40365 , \40349 , \40364 );
not \U$40023 ( \40366 , RIbb2d888_64);
not \U$40024 ( \40367 , \40343 );
or \U$40025 ( \40368 , \40366 , \40367 );
and \U$40026 ( \40369 , RIbb2d900_63, \16818 );
not \U$40027 ( \40370 , RIbb2d900_63);
and \U$40028 ( \40371 , \40370 , \16819 );
nor \U$40029 ( \40372 , \40369 , \40371 );
nand \U$40030 ( \40373 , \40372 , \17273 );
nand \U$40031 ( \40374 , \40368 , \40373 );
not \U$40032 ( \40375 , \40354 );
not \U$40033 ( \40376 , \40363 );
or \U$40034 ( \40377 , \40375 , \40376 );
or \U$40035 ( \40378 , \40363 , \40354 );
nand \U$40036 ( \40379 , \40377 , \40378 );
nor \U$40037 ( \40380 , \40374 , \40379 );
and \U$40038 ( \40381 , \17506 , \16532 );
not \U$40039 ( \40382 , RIbb2d888_64);
not \U$40040 ( \40383 , \40372 );
or \U$40041 ( \40384 , \40382 , \40383 );
and \U$40042 ( \40385 , RIbb2d900_63, \17517 );
not \U$40043 ( \40386 , RIbb2d900_63);
and \U$40044 ( \40387 , \40386 , \17744 );
nor \U$40045 ( \40388 , \40385 , \40387 );
nand \U$40046 ( \40389 , \40388 , \17273 );
nand \U$40047 ( \40390 , \40384 , \40389 );
xor \U$40048 ( \40391 , \40381 , \40390 );
not \U$40049 ( \40392 , RIbb2d888_64);
not \U$40050 ( \40393 , \40388 );
or \U$40051 ( \40394 , \40392 , \40393 );
nand \U$40052 ( \40395 , \19063 , \17273 );
nand \U$40053 ( \40396 , \40394 , \40395 );
not \U$40054 ( \40397 , \40396 );
nand \U$40055 ( \40398 , \17506 , RIbb2d888_64);
nand \U$40056 ( \40399 , \40398 , RIbb2d900_63);
nor \U$40057 ( \40400 , \40397 , \40399 );
and \U$40058 ( \40401 , \40391 , \40400 );
and \U$40059 ( \40402 , \40381 , \40390 );
or \U$40060 ( \40403 , \40401 , \40402 );
not \U$40061 ( \40404 , \40403 );
or \U$40062 ( \40405 , \40380 , \40404 );
nand \U$40063 ( \40406 , \40374 , \40379 );
nand \U$40064 ( \40407 , \40405 , \40406 );
nand \U$40065 ( \40408 , \40365 , \40407 );
or \U$40066 ( \40409 , \40349 , \40364 );
nand \U$40067 ( \40410 , \40408 , \40409 );
not \U$40068 ( \40411 , \40410 );
not \U$40069 ( \40412 , \16533 );
not \U$40070 ( \40413 , \40199 );
or \U$40071 ( \40414 , \40412 , \40413 );
nand \U$40072 ( \40415 , \40328 , \16541 );
nand \U$40073 ( \40416 , \40414 , \40415 );
xor \U$40074 ( \40417 , \40300 , \40309 );
xor \U$40075 ( \40418 , \40416 , \40417 );
not \U$40076 ( \40419 , RIbb2d888_64);
not \U$40077 ( \40420 , \40293 );
or \U$40078 ( \40421 , \40419 , \40420 );
nand \U$40079 ( \40422 , \40346 , \17273 );
nand \U$40080 ( \40423 , \40421 , \40422 );
xor \U$40081 ( \40424 , \40418 , \40423 );
not \U$40082 ( \40425 , \40322 );
nand \U$40083 ( \40426 , \40425 , \40348 );
not \U$40084 ( \40427 , \40348 );
nand \U$40085 ( \40428 , \40427 , \40322 );
nand \U$40086 ( \40429 , \40428 , \40337 );
nand \U$40087 ( \40430 , \40426 , \40429 );
nor \U$40088 ( \40431 , \40424 , \40430 );
or \U$40089 ( \40432 , \40411 , \40431 );
nand \U$40090 ( \40433 , \40430 , \40424 );
nand \U$40091 ( \40434 , \40432 , \40433 );
xor \U$40092 ( \40435 , \40416 , \40417 );
and \U$40093 ( \40436 , \40435 , \40423 );
and \U$40094 ( \40437 , \40416 , \40417 );
or \U$40095 ( \40438 , \40436 , \40437 );
not \U$40096 ( \40439 , \40438 );
xor \U$40097 ( \40440 , \40310 , \40295 );
xnor \U$40098 ( \40441 , \40440 , \40313 );
nand \U$40099 ( \40442 , \40439 , \40441 );
nand \U$40100 ( \40443 , \40434 , \40442 );
not \U$40101 ( \40444 , \40441 );
nand \U$40102 ( \40445 , \40444 , \40438 );
nand \U$40103 ( \40446 , \40443 , \40445 );
nand \U$40104 ( \40447 , \40321 , \40446 );
not \U$40105 ( \40448 , \40320 );
nand \U$40106 ( \40449 , \40448 , \40317 );
nand \U$40107 ( \40450 , \40447 , \40449 );
and \U$40108 ( \40451 , \40285 , \40450 );
and \U$40109 ( \40452 , \40263 , \40284 );
or \U$40110 ( \40453 , \40451 , \40452 );
xor \U$40111 ( \40454 , \40265 , \40269 );
and \U$40112 ( \40455 , \40454 , \40283 );
and \U$40113 ( \40456 , \40265 , \40269 );
or \U$40114 ( \40457 , \40455 , \40456 );
not \U$40115 ( \40458 , \40457 );
xor \U$40116 ( \40459 , \40128 , \40144 );
xor \U$40117 ( \40460 , \40459 , \40140 );
or \U$40118 ( \40461 , \40282 , \40276 );
not \U$40119 ( \40462 , \40271 );
nand \U$40120 ( \40463 , \40461 , \40462 );
nand \U$40121 ( \40464 , \40282 , \40276 );
and \U$40122 ( \40465 , \40463 , \40464 );
xor \U$40123 ( \40466 , \40460 , \40465 );
xor \U$40124 ( \40467 , \40071 , \40103 );
xnor \U$40125 ( \40468 , \40467 , \40060 );
xor \U$40126 ( \40469 , \40466 , \40468 );
nand \U$40127 ( \40470 , \40458 , \40469 );
nand \U$40128 ( \40471 , \40453 , \40470 );
not \U$40129 ( \40472 , \40469 );
nand \U$40130 ( \40473 , \40472 , \40457 );
nand \U$40131 ( \40474 , \40471 , \40473 );
not \U$40132 ( \40475 , \40108 );
not \U$40133 ( \40476 , \40048 );
or \U$40134 ( \40477 , \40475 , \40476 );
nand \U$40135 ( \40478 , \40107 , \40047 );
nand \U$40136 ( \40479 , \40477 , \40478 );
xnor \U$40137 ( \40480 , \40479 , \40148 );
xor \U$40138 ( \40481 , \40460 , \40465 );
and \U$40139 ( \40482 , \40481 , \40468 );
and \U$40140 ( \40483 , \40460 , \40465 );
or \U$40141 ( \40484 , \40482 , \40483 );
nand \U$40142 ( \40485 , \40480 , \40484 );
nand \U$40143 ( \40486 , \40474 , \40485 );
or \U$40144 ( \40487 , \40480 , \40484 );
nand \U$40145 ( \40488 , \40486 , \40487 );
not \U$40146 ( \40489 , \40488 );
or \U$40147 ( \40490 , \40176 , \40489 );
not \U$40148 ( \40491 , \40174 );
nand \U$40149 ( \40492 , \40491 , \40152 );
nand \U$40150 ( \40493 , \40490 , \40492 );
not \U$40151 ( \40494 , \40493 );
xor \U$40152 ( \40495 , \39871 , \39881 );
xor \U$40153 ( \40496 , \40495 , \39893 );
not \U$40154 ( \40497 , \40496 );
not \U$40155 ( \40498 , \40497 );
xor \U$40156 ( \40499 , \39939 , \39993 );
xnor \U$40157 ( \40500 , \40499 , \39990 );
not \U$40158 ( \40501 , \40500 );
or \U$40159 ( \40502 , \40498 , \40501 );
not \U$40160 ( \40503 , \40162 );
not \U$40161 ( \40504 , \40167 );
or \U$40162 ( \40505 , \40503 , \40504 );
or \U$40163 ( \40506 , \40167 , \40162 );
nand \U$40164 ( \40507 , \40506 , \40172 );
nand \U$40165 ( \40508 , \40505 , \40507 );
nand \U$40166 ( \40509 , \40502 , \40508 );
not \U$40167 ( \40510 , \40500 );
nand \U$40168 ( \40511 , \40510 , \40496 );
nand \U$40169 ( \40512 , \40509 , \40511 );
not \U$40170 ( \40513 , \40512 );
not \U$40171 ( \40514 , \39914 );
not \U$40172 ( \40515 , \39996 );
or \U$40173 ( \40516 , \40514 , \40515 );
or \U$40174 ( \40517 , \39996 , \39914 );
nand \U$40175 ( \40518 , \40516 , \40517 );
xnor \U$40176 ( \40519 , \40000 , \40518 );
nand \U$40177 ( \40520 , \40513 , \40519 );
not \U$40178 ( \40521 , \40508 );
not \U$40179 ( \40522 , \40497 );
or \U$40180 ( \40523 , \40521 , \40522 );
not \U$40181 ( \40524 , \40508 );
nand \U$40182 ( \40525 , \40524 , \40496 );
nand \U$40183 ( \40526 , \40523 , \40525 );
and \U$40184 ( \40527 , \40526 , \40500 );
not \U$40185 ( \40528 , \40526 );
and \U$40186 ( \40529 , \40528 , \40510 );
nor \U$40187 ( \40530 , \40527 , \40529 );
xor \U$40188 ( \40531 , \40155 , \40159 );
and \U$40189 ( \40532 , \40531 , \40173 );
and \U$40190 ( \40533 , \40155 , \40159 );
or \U$40191 ( \40534 , \40532 , \40533 );
nand \U$40192 ( \40535 , \40530 , \40534 );
and \U$40193 ( \40536 , \40520 , \40535 );
not \U$40194 ( \40537 , \40536 );
or \U$40195 ( \40538 , \40494 , \40537 );
nor \U$40196 ( \40539 , \40530 , \40534 );
nand \U$40197 ( \40540 , \40520 , \40539 );
not \U$40198 ( \40541 , \40519 );
nand \U$40199 ( \40542 , \40541 , \40512 );
and \U$40200 ( \40543 , \40540 , \40542 );
nand \U$40201 ( \40544 , \40538 , \40543 );
not \U$40202 ( \40545 , \40544 );
or \U$40203 ( \40546 , \40012 , \40545 );
not \U$40204 ( \40547 , \40010 );
nand \U$40205 ( \40548 , \40547 , \40004 );
nand \U$40206 ( \40549 , \40546 , \40548 );
not \U$40207 ( \40550 , \40549 );
or \U$40208 ( \40551 , \39912 , \40550 );
nand \U$40209 ( \40552 , \39910 , \39904 );
nand \U$40210 ( \40553 , \40551 , \40552 );
nand \U$40211 ( \40554 , \39518 , \39619 );
buf \U$40212 ( \40555 , \39695 );
nand \U$40213 ( \40556 , \39791 , \39698 );
nand \U$40214 ( \40557 , \40555 , \40556 );
nor \U$40215 ( \40558 , \40554 , \40557 );
nand \U$40216 ( \40559 , \39398 , \40553 , \40558 );
nand \U$40217 ( \40560 , \39824 , \40559 );
nand \U$40218 ( \40561 , \38562 , \38632 );
and \U$40219 ( \40562 , \38652 , \40561 );
and \U$40220 ( \40563 , \40562 , \38753 , \38394 );
nand \U$40221 ( \40564 , \40560 , \40563 );
nand \U$40222 ( \40565 , \38756 , \40564 );
and \U$40223 ( \40566 , \36638 , \36845 );
not \U$40224 ( \40567 , \36638 );
and \U$40225 ( \40568 , \40567 , \36844 );
nor \U$40226 ( \40569 , \40566 , \40568 );
xnor \U$40227 ( \40570 , \36636 , \40569 );
buf \U$40228 ( \40571 , \40570 );
xor \U$40229 ( \40572 , \36458 , \36474 );
xor \U$40230 ( \40573 , \40572 , \36492 );
or \U$40231 ( \40574 , \40571 , \40573 );
xor \U$40232 ( \40575 , \36723 , \36725 );
xor \U$40233 ( \40576 , \40575 , \36841 );
not \U$40234 ( \40577 , \40576 );
not \U$40235 ( \40578 , \38673 );
nand \U$40236 ( \40579 , \40578 , \38678 );
not \U$40237 ( \40580 , \40579 );
not \U$40238 ( \40581 , \38671 );
or \U$40239 ( \40582 , \40580 , \40581 );
nand \U$40240 ( \40583 , \38673 , \38675 );
nand \U$40241 ( \40584 , \40582 , \40583 );
xor \U$40242 ( \40585 , \36641 , \36685 );
xor \U$40243 ( \40586 , \40585 , \36720 );
buf \U$40244 ( \40587 , \40586 );
or \U$40245 ( \40588 , \40584 , \40587 );
xor \U$40246 ( \40589 , \38723 , \38728 );
and \U$40247 ( \40590 , \40589 , \38733 );
and \U$40248 ( \40591 , \38723 , \38728 );
or \U$40249 ( \40592 , \40590 , \40591 );
nand \U$40250 ( \40593 , \40588 , \40592 );
nand \U$40251 ( \40594 , \40584 , \40587 );
nand \U$40252 ( \40595 , \40593 , \40594 );
not \U$40253 ( \40596 , \40595 );
nand \U$40254 ( \40597 , \40577 , \40596 );
not \U$40255 ( \40598 , \40597 );
xor \U$40256 ( \40599 , \36620 , \36630 );
xor \U$40257 ( \40600 , \40599 , \36633 );
not \U$40258 ( \40601 , \40600 );
or \U$40259 ( \40602 , \40598 , \40601 );
nand \U$40260 ( \40603 , \40576 , \40595 );
nand \U$40261 ( \40604 , \40602 , \40603 );
nand \U$40262 ( \40605 , \40574 , \40604 );
nand \U$40263 ( \40606 , \40571 , \40573 );
nand \U$40264 ( \40607 , \40605 , \40606 );
not \U$40265 ( \40608 , \40607 );
xor \U$40266 ( \40609 , \36856 , \36855 );
xnor \U$40267 ( \40610 , \40609 , \36617 );
nand \U$40268 ( \40611 , \40608 , \40610 );
xor \U$40269 ( \40612 , \40573 , \40570 );
xnor \U$40270 ( \40613 , \40612 , \40604 );
xor \U$40271 ( \40614 , \36728 , \36766 );
xnor \U$40272 ( \40615 , \40614 , \36839 );
not \U$40273 ( \40616 , \40615 );
xor \U$40274 ( \40617 , \36624 , \36627 );
xnor \U$40275 ( \40618 , \40617 , \36622 );
not \U$40276 ( \40619 , \40618 );
or \U$40277 ( \40620 , \40616 , \40619 );
not \U$40278 ( \40621 , \38708 );
not \U$40279 ( \40622 , \38714 );
or \U$40280 ( \40623 , \40621 , \40622 );
or \U$40281 ( \40624 , \38714 , \38708 );
nand \U$40282 ( \40625 , \40624 , \38717 );
nand \U$40283 ( \40626 , \40623 , \40625 );
nand \U$40284 ( \40627 , \40620 , \40626 );
not \U$40285 ( \40628 , \40618 );
not \U$40286 ( \40629 , \40615 );
nand \U$40287 ( \40630 , \40628 , \40629 );
and \U$40288 ( \40631 , \40627 , \40630 );
not \U$40289 ( \40632 , \40592 );
and \U$40290 ( \40633 , \40586 , \40632 );
not \U$40291 ( \40634 , \40586 );
and \U$40292 ( \40635 , \40634 , \40592 );
or \U$40293 ( \40636 , \40633 , \40635 );
not \U$40294 ( \40637 , \40584 );
and \U$40295 ( \40638 , \40636 , \40637 );
not \U$40296 ( \40639 , \40636 );
and \U$40297 ( \40640 , \40639 , \40584 );
nor \U$40298 ( \40641 , \40638 , \40640 );
not \U$40299 ( \40642 , \40641 );
not \U$40300 ( \40643 , \40642 );
not \U$40301 ( \40644 , \38721 );
not \U$40302 ( \40645 , \40644 );
not \U$40303 ( \40646 , \38739 );
or \U$40304 ( \40647 , \40645 , \40646 );
or \U$40305 ( \40648 , \38739 , \40644 );
nand \U$40306 ( \40649 , \40648 , \38734 );
nand \U$40307 ( \40650 , \40647 , \40649 );
not \U$40308 ( \40651 , \40650 );
or \U$40309 ( \40652 , \40643 , \40651 );
not \U$40310 ( \40653 , \40641 );
not \U$40311 ( \40654 , \40650 );
not \U$40312 ( \40655 , \40654 );
or \U$40313 ( \40656 , \40653 , \40655 );
nor \U$40314 ( \40657 , \38689 , \38681 );
or \U$40315 ( \40658 , \40657 , \38695 );
nand \U$40316 ( \40659 , \38689 , \38681 );
nand \U$40317 ( \40660 , \40658 , \40659 );
nand \U$40318 ( \40661 , \40656 , \40660 );
nand \U$40319 ( \40662 , \40652 , \40661 );
not \U$40320 ( \40663 , \40662 );
xor \U$40321 ( \40664 , \40631 , \40663 );
not \U$40322 ( \40665 , \40576 );
not \U$40323 ( \40666 , \40596 );
and \U$40324 ( \40667 , \40665 , \40666 );
and \U$40325 ( \40668 , \40576 , \40596 );
nor \U$40326 ( \40669 , \40667 , \40668 );
and \U$40327 ( \40670 , \40600 , \40669 );
not \U$40328 ( \40671 , \40600 );
not \U$40329 ( \40672 , \40669 );
and \U$40330 ( \40673 , \40671 , \40672 );
nor \U$40331 ( \40674 , \40670 , \40673 );
and \U$40332 ( \40675 , \40664 , \40674 );
and \U$40333 ( \40676 , \40631 , \40663 );
or \U$40334 ( \40677 , \40675 , \40676 );
nand \U$40335 ( \40678 , \40613 , \40677 );
nand \U$40336 ( \40679 , \40611 , \40678 );
xor \U$40337 ( \40680 , \40631 , \40663 );
xor \U$40338 ( \40681 , \40680 , \40674 );
not \U$40339 ( \40682 , \40681 );
not \U$40340 ( \40683 , \40615 );
not \U$40341 ( \40684 , \40626 );
or \U$40342 ( \40685 , \40683 , \40684 );
or \U$40343 ( \40686 , \40626 , \40615 );
nand \U$40344 ( \40687 , \40685 , \40686 );
and \U$40345 ( \40688 , \40687 , \40618 );
not \U$40346 ( \40689 , \40687 );
and \U$40347 ( \40690 , \40689 , \40628 );
nor \U$40348 ( \40691 , \40688 , \40690 );
not \U$40349 ( \40692 , \38718 );
not \U$40350 ( \40693 , \38740 );
or \U$40351 ( \40694 , \40692 , \40693 );
nand \U$40352 ( \40695 , \40694 , \38750 );
not \U$40353 ( \40696 , \38740 );
nand \U$40354 ( \40697 , \40696 , \38719 );
nand \U$40355 ( \40698 , \40695 , \40697 );
not \U$40356 ( \40699 , \40698 );
xor \U$40357 ( \40700 , \40691 , \40699 );
not \U$40358 ( \40701 , \40641 );
not \U$40359 ( \40702 , \40650 );
or \U$40360 ( \40703 , \40701 , \40702 );
or \U$40361 ( \40704 , \40650 , \40641 );
nand \U$40362 ( \40705 , \40703 , \40704 );
not \U$40363 ( \40706 , \40660 );
and \U$40364 ( \40707 , \40705 , \40706 );
not \U$40365 ( \40708 , \40705 );
and \U$40366 ( \40709 , \40708 , \40660 );
nor \U$40367 ( \40710 , \40707 , \40709 );
and \U$40368 ( \40711 , \40700 , \40710 );
and \U$40369 ( \40712 , \40691 , \40699 );
or \U$40370 ( \40713 , \40711 , \40712 );
not \U$40371 ( \40714 , \40713 );
or \U$40372 ( \40715 , \40682 , \40714 );
or \U$40373 ( \40716 , \38703 , \38696 );
nand \U$40374 ( \40717 , \40716 , \38751 );
nand \U$40375 ( \40718 , \38703 , \38696 );
nand \U$40376 ( \40719 , \40717 , \40718 );
not \U$40377 ( \40720 , \40719 );
xor \U$40378 ( \40721 , \40691 , \40699 );
xor \U$40379 ( \40722 , \40721 , \40710 );
nand \U$40380 ( \40723 , \40720 , \40722 );
nand \U$40381 ( \40724 , \40715 , \40723 );
nor \U$40382 ( \40725 , \40679 , \40724 );
nand \U$40383 ( \40726 , \40565 , \40725 );
not \U$40384 ( \40727 , \40726 );
and \U$40385 ( \40728 , \35286 , \35446 , \37385 , \40727 );
not \U$40386 ( \40729 , \37230 );
nand \U$40387 ( \40730 , \36614 , \36858 );
not \U$40388 ( \40731 , \40730 );
nand \U$40389 ( \40732 , \37031 , \36864 );
not \U$40390 ( \40733 , \40732 );
or \U$40391 ( \40734 , \40731 , \40733 );
nand \U$40392 ( \40735 , \40734 , \37033 );
and \U$40393 ( \40736 , \37241 , \37242 );
not \U$40394 ( \40737 , \37241 );
and \U$40395 ( \40738 , \40737 , \37212 );
nor \U$40396 ( \40739 , \40736 , \40738 );
nor \U$40397 ( \40740 , \40739 , \37234 );
or \U$40398 ( \40741 , \40735 , \40740 );
nand \U$40399 ( \40742 , \40739 , \37234 );
nand \U$40400 ( \40743 , \40741 , \40742 );
not \U$40401 ( \40744 , \40743 );
or \U$40402 ( \40745 , \40729 , \40744 );
or \U$40403 ( \40746 , \37201 , \37229 );
nand \U$40404 ( \40747 , \40745 , \40746 );
and \U$40405 ( \40748 , \37374 , \37382 , \37331 , \37344 );
nand \U$40406 ( \40749 , \40747 , \40748 );
not \U$40407 ( \40750 , \40749 );
not \U$40408 ( \40751 , \37382 );
not \U$40409 ( \40752 , \37374 );
not \U$40410 ( \40753 , \37330 );
nor \U$40411 ( \40754 , \37333 , \37343 );
not \U$40412 ( \40755 , \40754 );
or \U$40413 ( \40756 , \40753 , \40755 );
not \U$40414 ( \40757 , \37316 );
not \U$40415 ( \40758 , \37329 );
nand \U$40416 ( \40759 , \40757 , \40758 );
nand \U$40417 ( \40760 , \40756 , \40759 );
not \U$40418 ( \40761 , \40760 );
or \U$40419 ( \40762 , \40752 , \40761 );
not \U$40420 ( \40763 , \37369 );
not \U$40421 ( \40764 , \37373 );
nand \U$40422 ( \40765 , \40763 , \40764 );
nand \U$40423 ( \40766 , \40762 , \40765 );
not \U$40424 ( \40767 , \40766 );
or \U$40425 ( \40768 , \40751 , \40767 );
not \U$40426 ( \40769 , \37377 );
not \U$40427 ( \40770 , \37381 );
nand \U$40428 ( \40771 , \40769 , \40770 );
nand \U$40429 ( \40772 , \40768 , \40771 );
not \U$40430 ( \40773 , \40772 );
not \U$40431 ( \40774 , \40773 );
or \U$40432 ( \40775 , \40750 , \40774 );
nand \U$40433 ( \40776 , \35284 , \35445 );
not \U$40434 ( \40777 , \40776 );
nand \U$40435 ( \40778 , \40775 , \40777 );
buf \U$40436 ( \40779 , \35414 );
not \U$40437 ( \40780 , \40779 );
and \U$40438 ( \40781 , \35431 , \35434 );
not \U$40439 ( \40782 , \35438 );
not \U$40440 ( \40783 , \35442 );
nand \U$40441 ( \40784 , \40782 , \40783 );
or \U$40442 ( \40785 , \40781 , \40784 );
or \U$40443 ( \40786 , \35434 , \35431 );
nand \U$40444 ( \40787 , \40785 , \40786 );
not \U$40445 ( \40788 , \40787 );
or \U$40446 ( \40789 , \40780 , \40788 );
or \U$40447 ( \40790 , \35380 , \35413 );
nand \U$40448 ( \40791 , \40789 , \40790 );
buf \U$40449 ( \40792 , \35370 );
and \U$40450 ( \40793 , \40791 , \40792 );
not \U$40451 ( \40794 , \35157 );
nor \U$40452 ( \40795 , \40794 , \35282 );
not \U$40453 ( \40796 , \40795 );
not \U$40454 ( \40797 , \35445 );
or \U$40455 ( \40798 , \40796 , \40797 );
or \U$40456 ( \40799 , \35295 , \35369 );
nand \U$40457 ( \40800 , \40798 , \40799 );
nor \U$40458 ( \40801 , \40793 , \40800 );
nand \U$40459 ( \40802 , \40778 , \40801 );
nor \U$40460 ( \40803 , \40728 , \40802 );
nor \U$40461 ( \40804 , \35285 , \37384 );
not \U$40462 ( \40805 , \40611 );
not \U$40463 ( \40806 , \40678 );
nand \U$40464 ( \40807 , \40681 , \40713 );
not \U$40465 ( \40808 , \40719 );
nor \U$40466 ( \40809 , \40808 , \40722 );
nand \U$40467 ( \40810 , \40807 , \40809 );
not \U$40468 ( \40811 , \40681 );
not \U$40469 ( \40812 , \40713 );
nand \U$40470 ( \40813 , \40811 , \40812 );
nand \U$40471 ( \40814 , \40810 , \40813 );
not \U$40472 ( \40815 , \40814 );
or \U$40473 ( \40816 , \40806 , \40815 );
not \U$40474 ( \40817 , \40613 );
not \U$40475 ( \40818 , \40677 );
nand \U$40476 ( \40819 , \40817 , \40818 );
nand \U$40477 ( \40820 , \40816 , \40819 );
not \U$40478 ( \40821 , \40820 );
or \U$40479 ( \40822 , \40805 , \40821 );
not \U$40480 ( \40823 , \40610 );
nand \U$40481 ( \40824 , \40823 , \40607 );
nand \U$40482 ( \40825 , \40822 , \40824 );
not \U$40483 ( \40826 , \40825 );
not \U$40484 ( \40827 , \40826 );
and \U$40485 ( \40828 , \40804 , \35446 , \40827 );
nand \U$40486 ( \40829 , \34755 , \34759 );
not \U$40487 ( \40830 , \40829 );
not \U$40488 ( \40831 , \34622 );
nor \U$40489 ( \40832 , \34762 , \35151 );
not \U$40490 ( \40833 , \40832 );
or \U$40491 ( \40834 , \40831 , \40833 );
not \U$40492 ( \40835 , \34253 );
not \U$40493 ( \40836 , \34621 );
nand \U$40494 ( \40837 , \40835 , \40836 );
nand \U$40495 ( \40838 , \40834 , \40837 );
not \U$40496 ( \40839 , \40838 );
or \U$40497 ( \40840 , \40830 , \40839 );
or \U$40498 ( \40841 , \34755 , \34759 );
nand \U$40499 ( \40842 , \40840 , \40841 );
buf \U$40500 ( \40843 , \35283 );
and \U$40501 ( \40844 , \35446 , \40842 , \40843 );
nor \U$40502 ( \40845 , \40828 , \40844 );
nand \U$40503 ( \40846 , \40803 , \40845 );
and \U$40504 ( \40847 , \32721 , \32550 );
not \U$40505 ( \40848 , \31723 );
not \U$40506 ( \40849 , \29851 );
not \U$40507 ( \40850 , \28361 );
not \U$40508 ( \40851 , \28922 );
nand \U$40509 ( \40852 , \40850 , \40851 );
and \U$40510 ( \40853 , \29364 , \40852 );
buf \U$40511 ( \40854 , \29361 );
nand \U$40512 ( \40855 , \40849 , \40853 , \40854 );
nor \U$40513 ( \40856 , \40848 , \40855 );
nand \U$40514 ( \40857 , \40846 , \40847 , \40856 );
nand \U$40515 ( \40858 , \32723 , \32744 , \40857 );
buf \U$40516 ( \40859 , \24550 );
not \U$40517 ( \40860 , \24558 );
or \U$40518 ( \40861 , \23833 , \24545 );
and \U$40519 ( \40862 , \22870 , \40859 , \40860 , \40861 );
and \U$40520 ( \40863 , \20630 , \21548 );
nand \U$40521 ( \40864 , \40862 , \40863 , \24580 , \24585 );
not \U$40522 ( \40865 , \40864 );
and \U$40523 ( \40866 , \25578 , \40858 , \40865 );
nor \U$40524 ( \40867 , \25615 , \40866 );
not \U$40525 ( \40868 , \40867 );
not \U$40526 ( \40869 , \40868 );
or \U$40527 ( \40870 , \16141 , \40869 );
not \U$40528 ( \40871 , \16127 );
not \U$40529 ( \40872 , \16139 );
and \U$40530 ( \40873 , \14463 , \15229 );
and \U$40531 ( \40874 , \15359 , \15886 );
or \U$40532 ( \40875 , \40873 , \40874 );
nand \U$40533 ( \40876 , \40875 , \15230 );
or \U$40534 ( \40877 , \40876 , \15356 );
nand \U$40535 ( \40878 , \15351 , \15355 );
nand \U$40536 ( \40879 , \40877 , \40878 );
not \U$40537 ( \40880 , \40879 );
or \U$40538 ( \40881 , \40872 , \40880 );
not \U$40539 ( \40882 , \16138 );
nand \U$40540 ( \40883 , \40882 , \16131 );
nand \U$40541 ( \40884 , \40881 , \40883 );
not \U$40542 ( \40885 , \40884 );
or \U$40543 ( \40886 , \40871 , \40885 );
not \U$40544 ( \40887 , \16126 );
not \U$40545 ( \40888 , \16114 );
not \U$40546 ( \40889 , \16096 );
and \U$40547 ( \40890 , \16060 , \15997 );
not \U$40548 ( \40891 , \40890 );
or \U$40549 ( \40892 , \40889 , \40891 );
not \U$40550 ( \40893 , \16090 );
not \U$40551 ( \40894 , \16095 );
nand \U$40552 ( \40895 , \40893 , \40894 );
nand \U$40553 ( \40896 , \40892 , \40895 );
not \U$40554 ( \40897 , \40896 );
or \U$40555 ( \40898 , \40888 , \40897 );
not \U$40556 ( \40899 , \16109 );
not \U$40557 ( \40900 , \16113 );
nand \U$40558 ( \40901 , \40899 , \40900 );
nand \U$40559 ( \40902 , \40898 , \40901 );
not \U$40560 ( \40903 , \40902 );
or \U$40561 ( \40904 , \40887 , \40903 );
not \U$40562 ( \40905 , \16125 );
nand \U$40563 ( \40906 , \40905 , \16122 );
nand \U$40564 ( \40907 , \40904 , \40906 );
not \U$40565 ( \40908 , \40907 );
nand \U$40566 ( \40909 , \40886 , \40908 );
buf \U$40567 ( \40910 , \11947 );
and \U$40568 ( \40911 , \40909 , \40910 );
not \U$40569 ( \40912 , \9637 );
not \U$40570 ( \40913 , \9582 );
nand \U$40571 ( \40914 , \40913 , \9528 );
or \U$40572 ( \40915 , \40912 , \40914 );
not \U$40573 ( \40916 , \9636 );
nand \U$40574 ( \40917 , \40916 , \9591 );
nand \U$40575 ( \40918 , \40915 , \40917 );
not \U$40576 ( \40919 , \9643 );
nand \U$40577 ( \40920 , \40919 , \9673 );
and \U$40578 ( \40921 , \40918 , \40920 );
not \U$40579 ( \40922 , \9643 );
nor \U$40580 ( \40923 , \40922 , \9673 );
nor \U$40581 ( \40924 , \40921 , \40923 );
not \U$40582 ( \40925 , \40924 );
not \U$40583 ( \40926 , \11924 );
not \U$40584 ( \40927 , \11896 );
nand \U$40585 ( \40928 , \40926 , \40927 );
not \U$40586 ( \40929 , \40928 );
nor \U$40587 ( \40930 , \11430 , \11890 );
not \U$40588 ( \40931 , \40930 );
not \U$40589 ( \40932 , \11427 );
or \U$40590 ( \40933 , \40931 , \40932 );
not \U$40591 ( \40934 , \10809 );
not \U$40592 ( \40935 , \11426 );
nand \U$40593 ( \40936 , \40934 , \40935 );
nand \U$40594 ( \40937 , \40933 , \40936 );
nand \U$40595 ( \40938 , \40937 , \11925 );
not \U$40596 ( \40939 , \40938 );
or \U$40597 ( \40940 , \40929 , \40939 );
not \U$40598 ( \40941 , \11935 );
nand \U$40599 ( \40942 , \40940 , \40941 );
nand \U$40600 ( \40943 , \11928 , \11934 );
nand \U$40601 ( \40944 , \40942 , \40943 );
nand \U$40602 ( \40945 , \40944 , \9675 );
not \U$40603 ( \40946 , \40945 );
or \U$40604 ( \40947 , \40925 , \40946 );
nand \U$40605 ( \40948 , \40947 , \11946 );
not \U$40606 ( \40949 , \11945 );
nand \U$40607 ( \40950 , \40949 , \11942 );
nand \U$40608 ( \40951 , \40948 , \40950 );
nor \U$40609 ( \40952 , \40911 , \40951 );
nand \U$40610 ( \40953 , \40870 , \40952 );
not \U$40611 ( \40954 , \40953 );
or \U$40612 ( \40955 , \8301 , \40954 );
not \U$40613 ( \40956 , \8298 );
not \U$40614 ( \40957 , \40956 );
not \U$40615 ( \40958 , \8290 );
not \U$40616 ( \40959 , \8178 );
not \U$40617 ( \40960 , \5823 );
not \U$40618 ( \40961 , \7545 );
not \U$40619 ( \40962 , \6572 );
and \U$40620 ( \40963 , \6903 , \7532 );
nand \U$40621 ( \40964 , \40963 , \6900 );
buf \U$40622 ( \40965 , \6575 );
nand \U$40623 ( \40966 , \40965 , \6898 );
nand \U$40624 ( \40967 , \40964 , \40966 );
not \U$40625 ( \40968 , \40967 );
or \U$40626 ( \40969 , \40962 , \40968 );
not \U$40627 ( \40970 , \6571 );
nand \U$40628 ( \40971 , \40970 , \6550 );
nand \U$40629 ( \40972 , \40969 , \40971 );
not \U$40630 ( \40973 , \40972 );
or \U$40631 ( \40974 , \40961 , \40973 );
nand \U$40632 ( \40975 , \7544 , \7542 );
nand \U$40633 ( \40976 , \40974 , \40975 );
not \U$40634 ( \40977 , \40976 );
or \U$40635 ( \40978 , \40960 , \40977 );
not \U$40636 ( \40979 , \5821 );
nand \U$40637 ( \40980 , \5109 , \4865 );
not \U$40638 ( \40981 , \40980 );
nand \U$40639 ( \40982 , \40981 , \5370 );
not \U$40640 ( \40983 , \5369 );
nand \U$40641 ( \40984 , \40983 , \5114 );
nand \U$40642 ( \40985 , \40982 , \40984 );
not \U$40643 ( \40986 , \40985 );
or \U$40644 ( \40987 , \40979 , \40986 );
or \U$40645 ( \40988 , \5816 , \5820 );
nand \U$40646 ( \40989 , \40987 , \40988 );
buf \U$40647 ( \40990 , \5814 );
and \U$40648 ( \40991 , \40989 , \40990 );
and \U$40649 ( \40992 , \5788 , \5813 );
nor \U$40650 ( \40993 , \40991 , \40992 );
nand \U$40651 ( \40994 , \40978 , \40993 );
not \U$40652 ( \40995 , \40994 );
or \U$40653 ( \40996 , \40959 , \40995 );
not \U$40654 ( \40997 , \8126 );
not \U$40655 ( \40998 , \8150 );
nand \U$40656 ( \40999 , \8171 , \8175 );
or \U$40657 ( \41000 , \8168 , \40999 );
nand \U$40658 ( \41001 , \8165 , \8167 );
nand \U$40659 ( \41002 , \41000 , \41001 );
not \U$40660 ( \41003 , \41002 );
or \U$40661 ( \41004 , \40998 , \41003 );
not \U$40662 ( \41005 , \8149 );
nand \U$40663 ( \41006 , \41005 , \8146 );
nand \U$40664 ( \41007 , \41004 , \41006 );
not \U$40665 ( \41008 , \41007 );
or \U$40666 ( \41009 , \40997 , \41008 );
nand \U$40667 ( \41010 , \8085 , \8125 );
nand \U$40668 ( \41011 , \41009 , \41010 );
not \U$40669 ( \41012 , \41011 );
nand \U$40670 ( \41013 , \40996 , \41012 );
not \U$40671 ( \41014 , \41013 );
or \U$40672 ( \41015 , \40958 , \41014 );
nand \U$40673 ( \41016 , \8266 , \8269 );
buf \U$40674 ( \41017 , \8261 );
or \U$40675 ( \41018 , \41016 , \41017 );
nand \U$40676 ( \41019 , \8246 , \8260 );
nand \U$40677 ( \41020 , \41018 , \41019 );
not \U$40678 ( \41021 , \8289 );
and \U$40679 ( \41022 , \41020 , \41021 );
and \U$40680 ( \41023 , \8284 , \8288 );
nor \U$40681 ( \41024 , \41022 , \41023 );
nand \U$40682 ( \41025 , \41015 , \41024 );
not \U$40683 ( \41026 , \41025 );
or \U$40684 ( \41027 , \40957 , \41026 );
nand \U$40685 ( \41028 , \8295 , \8297 );
nand \U$40686 ( \41029 , \41027 , \41028 );
not \U$40687 ( \41030 , \41029 );
nand \U$40688 ( \41031 , \40955 , \41030 );
not \U$40689 ( \41032 , \41031 );
or \U$40690 ( \41033 , \2907 , \41032 );
not \U$40691 ( \41034 , \2905 );
not \U$40692 ( \41035 , \2634 );
not \U$40693 ( \41036 , \2641 );
nand \U$40694 ( \41037 , \2192 , \2316 );
or \U$40695 ( \41038 , \41037 , \2431 );
nand \U$40696 ( \41039 , \2426 , \2430 );
nand \U$40697 ( \41040 , \41038 , \41039 );
not \U$40698 ( \41041 , \41040 );
or \U$40699 ( \41042 , \41036 , \41041 );
nand \U$40700 ( \41043 , \2640 , \2636 );
nand \U$40701 ( \41044 , \41042 , \41043 );
not \U$40702 ( \41045 , \41044 );
or \U$40703 ( \41046 , \41035 , \41045 );
nand \U$40704 ( \41047 , \2615 , \2633 );
nand \U$40705 ( \41048 , \41046 , \41047 );
not \U$40706 ( \41049 , \41048 );
or \U$40707 ( \41050 , \41034 , \41049 );
nand \U$40708 ( \41051 , \2729 , \2733 );
or \U$40709 ( \41052 , \41051 , \2824 );
nand \U$40710 ( \41053 , \2823 , \2738 );
nand \U$40711 ( \41054 , \41052 , \41053 );
and \U$40712 ( \41055 , \41054 , \2904 );
and \U$40713 ( \41056 , \2829 , \2903 );
nor \U$40714 ( \41057 , \41055 , \41056 );
nand \U$40715 ( \41058 , \41050 , \41057 );
not \U$40716 ( \41059 , \41058 );
nand \U$40717 ( \41060 , \41033 , \41059 );
xor \U$40718 ( \41061 , \2833 , \2883 );
and \U$40719 ( \41062 , \41061 , \2902 );
and \U$40720 ( \41063 , \2833 , \2883 );
or \U$40721 ( \41064 , \41062 , \41063 );
or \U$40722 ( \41065 , \2843 , \1771 );
or \U$40723 ( \41066 , \2133 , \1524 );
nand \U$40724 ( \41067 , \41065 , \41066 );
not \U$40725 ( \41068 , \41067 );
and \U$40726 ( \41069 , \1733 , \1394 );
xor \U$40727 ( \41070 , \41068 , \41069 );
not \U$40728 ( \41071 , \1147 );
and \U$40729 ( \41072 , \1477 , RIbb2f430_5);
not \U$40730 ( \41073 , \1477 );
and \U$40731 ( \41074 , \41073 , \1898 );
nor \U$40732 ( \41075 , \41072 , \41074 );
not \U$40733 ( \41076 , \41075 );
or \U$40734 ( \41077 , \41071 , \41076 );
not \U$40735 ( \41078 , \2851 );
or \U$40736 ( \41079 , \41078 , \1621 );
nand \U$40737 ( \41080 , \41077 , \41079 );
xor \U$40738 ( \41081 , \41070 , \41080 );
xor \U$40739 ( \41082 , \2839 , \2845 );
and \U$40740 ( \41083 , \41082 , \2855 );
and \U$40741 ( \41084 , \2839 , \2845 );
or \U$40742 ( \41085 , \41083 , \41084 );
xor \U$40743 ( \41086 , \2863 , \2871 );
and \U$40744 ( \41087 , \41086 , \2881 );
and \U$40745 ( \41088 , \2863 , \2871 );
or \U$40746 ( \41089 , \41087 , \41088 );
xor \U$40747 ( \41090 , \41085 , \41089 );
xor \U$40748 ( \41091 , \41081 , \41090 );
not \U$40749 ( \41092 , \1430 );
not \U$40750 ( \41093 , \2859 );
or \U$40751 ( \41094 , \41092 , \41093 );
xor \U$40752 ( \41095 , \1394 , \1042 );
nand \U$40753 ( \41096 , \41095 , \1376 );
nand \U$40754 ( \41097 , \41094 , \41096 );
not \U$40755 ( \41098 , \1294 );
and \U$40756 ( \41099 , \1291 , \953 );
not \U$40757 ( \41100 , \1291 );
and \U$40758 ( \41101 , \41100 , \957 );
nor \U$40759 ( \41102 , \41099 , \41101 );
not \U$40760 ( \41103 , \41102 );
or \U$40761 ( \41104 , \41098 , \41103 );
nand \U$40762 ( \41105 , \2878 , \1265 );
nand \U$40763 ( \41106 , \41104 , \41105 );
xor \U$40764 ( \41107 , \41097 , \41106 );
not \U$40765 ( \41108 , \1737 );
and \U$40766 ( \41109 , \1581 , RIbb2f340_7);
not \U$40767 ( \41110 , \1581 );
and \U$40768 ( \41111 , \41110 , \1734 );
nor \U$40769 ( \41112 , \41109 , \41111 );
not \U$40770 ( \41113 , \41112 );
or \U$40771 ( \41114 , \41108 , \41113 );
or \U$40772 ( \41115 , \2869 , \1703 );
nand \U$40773 ( \41116 , \41114 , \41115 );
xor \U$40774 ( \41117 , \41107 , \41116 );
xor \U$40775 ( \41118 , \2753 , \2886 );
and \U$40776 ( \41119 , \41118 , \2891 );
and \U$40777 ( \41120 , \2753 , \2886 );
or \U$40778 ( \41121 , \41119 , \41120 );
xor \U$40779 ( \41122 , \41117 , \41121 );
xor \U$40780 ( \41123 , \2837 , \2856 );
and \U$40781 ( \41124 , \41123 , \2882 );
and \U$40782 ( \41125 , \2837 , \2856 );
or \U$40783 ( \41126 , \41124 , \41125 );
xor \U$40784 ( \41127 , \41122 , \41126 );
xor \U$40785 ( \41128 , \41091 , \41127 );
xor \U$40786 ( \41129 , \2753 , \2886 );
xor \U$40787 ( \41130 , \41129 , \2891 );
and \U$40788 ( \41131 , \2896 , \41130 );
xor \U$40789 ( \41132 , \2753 , \2886 );
xor \U$40790 ( \41133 , \41132 , \2891 );
and \U$40791 ( \41134 , \2900 , \41133 );
and \U$40792 ( \41135 , \2896 , \2900 );
or \U$40793 ( \41136 , \41131 , \41134 , \41135 );
xor \U$40794 ( \41137 , \41128 , \41136 );
or \U$40795 ( \41138 , \41064 , \41137 );
nand \U$40796 ( \41139 , \41064 , \41137 );
nand \U$40797 ( \41140 , \41138 , \41139 );
xor \U$40798 ( \41141 , \41060 , \41140 );
xor \U$40799 ( \41142 , RIbb345c0_231, RIbb34bd8_244);
and \U$40800 ( \41143 , RIbb336c0_199, RIbb34278_224);
not \U$40801 ( \41144 , RIbb336c0_199);
not \U$40802 ( \41145 , RIbb34278_224);
and \U$40803 ( \41146 , \41144 , \41145 );
nor \U$40804 ( \41147 , \41143 , \41146 );
xor \U$40805 ( \41148 , \41142 , \41147 );
not \U$40806 ( \41149 , RIbb338a0_203);
nand \U$40807 ( \41150 , \41149 , RIbb34db8_248);
not \U$40808 ( \41151 , RIbb34db8_248);
nand \U$40809 ( \41152 , \41151 , RIbb338a0_203);
nand \U$40810 ( \41153 , \41150 , \41152 );
not \U$40811 ( \41154 , \41153 );
not \U$40812 ( \41155 , RIbb33a08_206);
and \U$40813 ( \41156 , RIbb34098_220, \41155 );
not \U$40814 ( \41157 , RIbb34098_220);
and \U$40815 ( \41158 , \41157 , RIbb33a08_206);
nor \U$40816 ( \41159 , \41156 , \41158 );
not \U$40817 ( \41160 , \41159 );
or \U$40818 ( \41161 , \41154 , \41160 );
or \U$40819 ( \41162 , \41159 , \41153 );
nand \U$40820 ( \41163 , \41161 , \41162 );
xor \U$40821 ( \41164 , \41148 , \41163 );
xnor \U$40822 ( \41165 , RIbb34110_221, RIbb33990_205);
not \U$40823 ( \41166 , \41165 );
and \U$40824 ( \41167 , RIbb347a0_235, RIbb34cc8_246);
not \U$40825 ( \41168 , RIbb347a0_235);
not \U$40826 ( \41169 , RIbb34cc8_246);
and \U$40827 ( \41170 , \41168 , \41169 );
nor \U$40828 ( \41171 , \41167 , \41170 );
not \U$40829 ( \41172 , \41171 );
and \U$40830 ( \41173 , \41166 , \41172 );
and \U$40831 ( \41174 , \41165 , \41171 );
nor \U$40832 ( \41175 , \41173 , \41174 );
not \U$40833 ( \41176 , RIbb33c60_211);
not \U$40834 ( \41177 , RIbb34d40_247);
not \U$40835 ( \41178 , \41177 );
or \U$40836 ( \41179 , \41176 , \41178 );
not \U$40837 ( \41180 , RIbb33c60_211);
nand \U$40838 ( \41181 , \41180 , RIbb34d40_247);
nand \U$40839 ( \41182 , \41179 , \41181 );
not \U$40840 ( \41183 , \41182 );
not \U$40841 ( \41184 , RIbb33d50_213);
and \U$40842 ( \41185 , RIbb33f30_217, \41184 );
not \U$40843 ( \41186 , RIbb33f30_217);
and \U$40844 ( \41187 , \41186 , RIbb33d50_213);
nor \U$40845 ( \41188 , \41185 , \41187 );
not \U$40846 ( \41189 , \41188 );
or \U$40847 ( \41190 , \41183 , \41189 );
or \U$40848 ( \41191 , \41188 , \41182 );
nand \U$40849 ( \41192 , \41190 , \41191 );
xor \U$40850 ( \41193 , \41175 , \41192 );
xor \U$40851 ( \41194 , \41164 , \41193 );
not \U$40852 ( \41195 , \41194 );
not \U$40853 ( \41196 , RIbb34548_230);
nand \U$40854 ( \41197 , \41196 , RIbb34ea8_250);
not \U$40855 ( \41198 , RIbb34ea8_250);
nand \U$40856 ( \41199 , \41198 , RIbb34548_230);
nand \U$40857 ( \41200 , \41197 , \41199 );
not \U$40858 ( \41201 , \41200 );
xnor \U$40859 ( \41202 , RIbb34908_238, RIbb33a80_207);
not \U$40860 ( \41203 , \41202 );
or \U$40861 ( \41204 , \41201 , \41203 );
or \U$40862 ( \41205 , \41202 , \41200 );
nand \U$40863 ( \41206 , \41204 , \41205 );
not \U$40864 ( \41207 , \41206 );
xor \U$40865 ( \41208 , RIbb334e0_195, RIbb35010_253);
xor \U$40866 ( \41209 , RIbb33738_200, RIbb349f8_240);
xor \U$40867 ( \41210 , \41208 , \41209 );
nand \U$40868 ( \41211 , \41207 , \41210 );
not \U$40869 ( \41212 , \41210 );
nand \U$40870 ( \41213 , \41212 , \41206 );
nand \U$40871 ( \41214 , \41211 , \41213 );
xor \U$40872 ( \41215 , RIbb33918_204, RIbb34980_239);
and \U$40873 ( \41216 , RIbb33828_202, RIbb34188_222);
not \U$40874 ( \41217 , RIbb33828_202);
not \U$40875 ( \41218 , RIbb34188_222);
and \U$40876 ( \41219 , \41217 , \41218 );
nor \U$40877 ( \41220 , \41216 , \41219 );
xor \U$40878 ( \41221 , \41215 , \41220 );
not \U$40879 ( \41222 , RIbb34728_234);
nand \U$40880 ( \41223 , \41222 , RIbb35088_254);
not \U$40881 ( \41224 , RIbb35088_254);
nand \U$40882 ( \41225 , \41224 , RIbb34728_234);
nand \U$40883 ( \41226 , \41223 , \41225 );
not \U$40884 ( \41227 , \41226 );
not \U$40885 ( \41228 , RIbb34638_232);
and \U$40886 ( \41229 , RIbb346b0_233, \41228 );
not \U$40887 ( \41230 , RIbb346b0_233);
and \U$40888 ( \41231 , \41230 , RIbb34638_232);
nor \U$40889 ( \41232 , \41229 , \41231 );
not \U$40890 ( \41233 , \41232 );
or \U$40891 ( \41234 , \41227 , \41233 );
or \U$40892 ( \41235 , \41232 , \41226 );
nand \U$40893 ( \41236 , \41234 , \41235 );
xor \U$40894 ( \41237 , \41221 , \41236 );
xor \U$40895 ( \41238 , \41214 , \41237 );
not \U$40896 ( \41239 , \41238 );
or \U$40897 ( \41240 , \41195 , \41239 );
or \U$40898 ( \41241 , \41194 , \41238 );
nand \U$40899 ( \41242 , \41240 , \41241 );
not \U$40900 ( \41243 , \41242 );
xor \U$40901 ( \41244 , RIbb34458_228, RIbb34ae8_242);
xor \U$40902 ( \41245 , RIbb33b70_209, RIbb33fa8_218);
xnor \U$40903 ( \41246 , \41244 , \41245 );
xor \U$40904 ( \41247 , RIbb33558_196, RIbb34e30_249);
xor \U$40905 ( \41248 , RIbb33af8_208, RIbb34020_219);
xor \U$40906 ( \41249 , \41247 , \41248 );
xor \U$40907 ( \41250 , \41246 , \41249 );
not \U$40908 ( \41251 , RIbb333f0_193);
not \U$40909 ( \41252 , RIbb35178_256);
not \U$40910 ( \41253 , \41252 );
or \U$40911 ( \41254 , \41251 , \41253 );
not \U$40912 ( \41255 , RIbb333f0_193);
nand \U$40913 ( \41256 , \41255 , RIbb35178_256);
nand \U$40914 ( \41257 , \41254 , \41256 );
not \U$40915 ( \41258 , \41257 );
xnor \U$40916 ( \41259 , RIbb343e0_227, RIbb34368_226);
not \U$40917 ( \41260 , \41259 );
or \U$40918 ( \41261 , \41258 , \41260 );
or \U$40919 ( \41262 , \41259 , \41257 );
nand \U$40920 ( \41263 , \41261 , \41262 );
not \U$40921 ( \41264 , \41263 );
xnor \U$40922 ( \41265 , RIbb34a70_241, RIbb335d0_197);
not \U$40923 ( \41266 , \41265 );
xor \U$40924 ( \41267 , RIbb344d0_229, RIbb34b60_243);
not \U$40925 ( \41268 , \41267 );
and \U$40926 ( \41269 , \41266 , \41268 );
and \U$40927 ( \41270 , \41265 , \41267 );
nor \U$40928 ( \41271 , \41269 , \41270 );
not \U$40929 ( \41272 , \41271 );
or \U$40930 ( \41273 , \41264 , \41272 );
or \U$40931 ( \41274 , \41271 , \41263 );
nand \U$40932 ( \41275 , \41273 , \41274 );
xor \U$40933 ( \41276 , \41250 , \41275 );
xor \U$40934 ( \41277 , RIbb33be8_210, RIbb34f98_252);
xor \U$40935 ( \41278 , RIbb33cd8_212, RIbb34890_237);
xor \U$40936 ( \41279 , \41277 , \41278 );
not \U$40937 ( \41280 , \41279 );
not \U$40938 ( \41281 , \41280 );
not \U$40939 ( \41282 , RIbb33648_198);
and \U$40940 ( \41283 , RIbb342f0_225, \41282 );
not \U$40941 ( \41284 , RIbb342f0_225);
and \U$40942 ( \41285 , \41284 , RIbb33648_198);
nor \U$40943 ( \41286 , \41283 , \41285 );
xor \U$40944 ( \41287 , RIbb34c50_245, RIbb34f20_251);
xor \U$40945 ( \41288 , \41286 , \41287 );
not \U$40946 ( \41289 , \41288 );
not \U$40947 ( \41290 , \41289 );
or \U$40948 ( \41291 , \41281 , \41290 );
nand \U$40949 ( \41292 , \41288 , \41279 );
nand \U$40950 ( \41293 , \41291 , \41292 );
xnor \U$40951 ( \41294 , RIbb33468_194, RIbb35100_255);
and \U$40952 ( \41295 , RIbb337b0_201, RIbb34200_223);
not \U$40953 ( \41296 , RIbb337b0_201);
not \U$40954 ( \41297 , RIbb34200_223);
and \U$40955 ( \41298 , \41296 , \41297 );
nor \U$40956 ( \41299 , \41295 , \41298 );
xor \U$40957 ( \41300 , \41294 , \41299 );
and \U$40958 ( \41301 , RIbb33eb8_216, RIbb34818_236);
not \U$40959 ( \41302 , RIbb33eb8_216);
not \U$40960 ( \41303 , RIbb34818_236);
and \U$40961 ( \41304 , \41302 , \41303 );
nor \U$40962 ( \41305 , \41301 , \41304 );
and \U$40963 ( \41306 , RIbb33dc8_214, RIbb33e40_215);
not \U$40964 ( \41307 , RIbb33dc8_214);
not \U$40965 ( \41308 , RIbb33e40_215);
and \U$40966 ( \41309 , \41307 , \41308 );
nor \U$40967 ( \41310 , \41306 , \41309 );
xor \U$40968 ( \41311 , \41305 , \41310 );
xor \U$40969 ( \41312 , \41300 , \41311 );
xnor \U$40970 ( \41313 , \41293 , \41312 );
and \U$40971 ( \41314 , \41276 , \41313 );
nor \U$40972 ( \41315 , \41276 , \41313 );
nor \U$40973 ( \41316 , \41314 , \41315 );
not \U$40974 ( \41317 , \41316 );
or \U$40975 ( \41318 , \41243 , \41317 );
or \U$40976 ( \41319 , \41316 , \41242 );
nand \U$40977 ( \41320 , \41318 , \41319 );
not \U$40978 ( \41321 , \41320 );
buf \U$40979 ( \41322 , \41321 );
buf \U$40980 ( \41323 , \41322 );
nor \U$40981 ( \41324 , \41141 , \41323 );
buf \U$40982 ( \41325 , \41324 );
not \U$40983 ( \41326 , \2825 );
not \U$40984 ( \41327 , \2642 );
not \U$40985 ( \41328 , \8300 );
nor \U$40986 ( \41329 , \41327 , \41328 );
not \U$40987 ( \41330 , \41329 );
buf \U$40988 ( \41331 , \40953 );
not \U$40989 ( \41332 , \41331 );
or \U$40990 ( \41333 , \41330 , \41332 );
and \U$40991 ( \41334 , \2642 , \41029 );
nor \U$40992 ( \41335 , \41334 , \41048 );
nand \U$40993 ( \41336 , \41333 , \41335 );
not \U$40994 ( \41337 , \41336 );
or \U$40995 ( \41338 , \41326 , \41337 );
not \U$40996 ( \41339 , \41054 );
nand \U$40997 ( \41340 , \41338 , \41339 );
not \U$40998 ( \41341 , \2904 );
nor \U$40999 ( \41342 , \41341 , \41056 );
xnor \U$41000 ( \41343 , \41340 , \41342 );
buf \U$41001 ( \41344 , \41320 );
not \U$41002 ( \41345 , \41344 );
nor \U$41003 ( \41346 , \41343 , \41345 );
buf \U$41004 ( \41347 , \41346 );
or \U$41005 ( \41348 , \2729 , \2733 );
nand \U$41006 ( \41349 , \41348 , \41051 );
xor \U$41007 ( \41350 , \41336 , \41349 );
nor \U$41008 ( \41351 , \41350 , \41323 );
buf \U$41009 ( \41352 , \41351 );
not \U$41010 ( \41353 , \2317 );
not \U$41011 ( \41354 , \41353 );
not \U$41012 ( \41355 , \41031 );
or \U$41013 ( \41356 , \41354 , \41355 );
nand \U$41014 ( \41357 , \41356 , \41037 );
not \U$41015 ( \41358 , \2431 );
nand \U$41016 ( \41359 , \41358 , \41039 );
xor \U$41017 ( \41360 , \41357 , \41359 );
nor \U$41018 ( \41361 , \41360 , \41323 );
buf \U$41019 ( \41362 , \41361 );
not \U$41020 ( \41363 , \8291 );
not \U$41021 ( \41364 , \41363 );
not \U$41022 ( \41365 , \7547 );
not \U$41023 ( \41366 , \40953 );
or \U$41024 ( \41367 , \41365 , \41366 );
buf \U$41025 ( \41368 , \40994 );
not \U$41026 ( \41369 , \41368 );
nand \U$41027 ( \41370 , \41367 , \41369 );
not \U$41028 ( \41371 , \41370 );
or \U$41029 ( \41372 , \41364 , \41371 );
and \U$41030 ( \41373 , \41011 , \8290 );
not \U$41031 ( \41374 , \41024 );
nor \U$41032 ( \41375 , \41373 , \41374 );
nand \U$41033 ( \41376 , \41372 , \41375 );
nand \U$41034 ( \41377 , \40956 , \41028 );
xor \U$41035 ( \41378 , \41376 , \41377 );
nor \U$41036 ( \41379 , \41378 , \41323 );
buf \U$41037 ( \41380 , \41379 );
not \U$41038 ( \41381 , \5821 );
nor \U$41039 ( \41382 , \7546 , \5371 );
not \U$41040 ( \41383 , \41382 );
not \U$41041 ( \41384 , \41331 );
or \U$41042 ( \41385 , \41383 , \41384 );
buf \U$41043 ( \41386 , \40976 );
not \U$41044 ( \41387 , \5371 );
and \U$41045 ( \41388 , \41386 , \41387 );
buf \U$41046 ( \41389 , \40985 );
nor \U$41047 ( \41390 , \41388 , \41389 );
nand \U$41048 ( \41391 , \41385 , \41390 );
not \U$41049 ( \41392 , \41391 );
or \U$41050 ( \41393 , \41381 , \41392 );
nand \U$41051 ( \41394 , \41393 , \40988 );
not \U$41052 ( \41395 , \40992 );
nand \U$41053 ( \41396 , \41395 , \40990 );
xor \U$41054 ( \41397 , \41394 , \41396 );
nor \U$41055 ( \41398 , \41397 , \41323 );
buf \U$41056 ( \41399 , \41398 );
not \U$41057 ( \41400 , \7546 );
not \U$41058 ( \41401 , \41400 );
not \U$41059 ( \41402 , \41331 );
or \U$41060 ( \41403 , \41401 , \41402 );
not \U$41061 ( \41404 , \41386 );
nand \U$41062 ( \41405 , \41403 , \41404 );
nand \U$41063 ( \41406 , \5110 , \40980 );
xor \U$41064 ( \41407 , \41405 , \41406 );
nor \U$41065 ( \41408 , \41407 , \41345 );
buf \U$41066 ( \41409 , \41408 );
not \U$41067 ( \41410 , \7535 );
buf \U$41068 ( \41411 , \41331 );
not \U$41069 ( \41412 , \41411 );
or \U$41070 ( \41413 , \41410 , \41412 );
not \U$41071 ( \41414 , \40972 );
nand \U$41072 ( \41415 , \41413 , \41414 );
nand \U$41073 ( \41416 , \7545 , \40975 );
xor \U$41074 ( \41417 , \41415 , \41416 );
nor \U$41075 ( \41418 , \41417 , \41345 );
buf \U$41076 ( \41419 , \41418 );
not \U$41077 ( \41420 , \7533 );
not \U$41078 ( \41421 , \41411 );
or \U$41079 ( \41422 , \41420 , \41421 );
not \U$41080 ( \41423 , \40963 );
nand \U$41081 ( \41424 , \41422 , \41423 );
nand \U$41082 ( \41425 , \6901 , \40966 );
xor \U$41083 ( \41426 , \41424 , \41425 );
buf \U$41084 ( \41427 , \41344 );
not \U$41085 ( \41428 , \41427 );
nor \U$41086 ( \41429 , \41426 , \41428 );
buf \U$41087 ( \41430 , \41429 );
not \U$41088 ( \41431 , \9583 );
nor \U$41089 ( \41432 , \41431 , \40912 );
not \U$41090 ( \41433 , \41432 );
and \U$41091 ( \41434 , \11936 , \11892 );
not \U$41092 ( \41435 , \41434 );
and \U$41093 ( \41436 , \15888 , \16127 , \16139 );
not \U$41094 ( \41437 , \41436 );
not \U$41095 ( \41438 , \40867 );
not \U$41096 ( \41439 , \41438 );
or \U$41097 ( \41440 , \41437 , \41439 );
not \U$41098 ( \41441 , \40909 );
nand \U$41099 ( \41442 , \41440 , \41441 );
not \U$41100 ( \41443 , \41442 );
or \U$41101 ( \41444 , \41435 , \41443 );
not \U$41102 ( \41445 , \40944 );
nand \U$41103 ( \41446 , \41444 , \41445 );
not \U$41104 ( \41447 , \41446 );
or \U$41105 ( \41448 , \41433 , \41447 );
not \U$41106 ( \41449 , \40918 );
nand \U$41107 ( \41450 , \41448 , \41449 );
not \U$41108 ( \41451 , \40923 );
nand \U$41109 ( \41452 , \41451 , \40920 );
xor \U$41110 ( \41453 , \41450 , \41452 );
nor \U$41111 ( \41454 , \41453 , \41428 );
buf \U$41112 ( \41455 , \41454 );
not \U$41113 ( \41456 , \9583 );
not \U$41114 ( \41457 , \41446 );
or \U$41115 ( \41458 , \41456 , \41457 );
nand \U$41116 ( \41459 , \41458 , \40914 );
nand \U$41117 ( \41460 , \40917 , \9637 );
xor \U$41118 ( \41461 , \41459 , \41460 );
nor \U$41119 ( \41462 , \41461 , \41428 );
buf \U$41120 ( \41463 , \41462 );
nand \U$41121 ( \41464 , \9583 , \40914 );
xor \U$41122 ( \41465 , \41446 , \41464 );
nor \U$41123 ( \41466 , \41465 , \41428 );
buf \U$41124 ( \41467 , \41466 );
not \U$41125 ( \41468 , \11925 );
not \U$41126 ( \41469 , \11892 );
not \U$41127 ( \41470 , \41442 );
or \U$41128 ( \41471 , \41469 , \41470 );
not \U$41129 ( \41472 , \40937 );
nand \U$41130 ( \41473 , \41471 , \41472 );
not \U$41131 ( \41474 , \41473 );
or \U$41132 ( \41475 , \41468 , \41474 );
nand \U$41133 ( \41476 , \41475 , \40928 );
nand \U$41134 ( \41477 , \40941 , \40943 );
xor \U$41135 ( \41478 , \41476 , \41477 );
nor \U$41136 ( \41479 , \41478 , \41428 );
buf \U$41137 ( \41480 , \41479 );
not \U$41138 ( \41481 , \11891 );
not \U$41139 ( \41482 , \41442 );
or \U$41140 ( \41483 , \41481 , \41482 );
not \U$41141 ( \41484 , \40930 );
nand \U$41142 ( \41485 , \41483 , \41484 );
nand \U$41143 ( \41486 , \40936 , \11428 );
xor \U$41144 ( \41487 , \41485 , \41486 );
nor \U$41145 ( \41488 , \41487 , \41428 );
buf \U$41146 ( \41489 , \41488 );
nand \U$41147 ( \41490 , \41484 , \11891 );
not \U$41148 ( \41491 , \41490 );
not \U$41149 ( \41492 , \41442 );
or \U$41150 ( \41493 , \41491 , \41492 );
or \U$41151 ( \41494 , \41442 , \41490 );
nand \U$41152 ( \41495 , \41493 , \41494 );
and \U$41153 ( \41496 , \41495 , \41427 );
buf \U$41154 ( \41497 , \41496 );
not \U$41155 ( \41498 , \16114 );
and \U$41156 ( \41499 , \16061 , \16096 );
not \U$41157 ( \41500 , \41499 );
and \U$41158 ( \41501 , \15888 , \16139 );
not \U$41159 ( \41502 , \41501 );
not \U$41160 ( \41503 , \41438 );
or \U$41161 ( \41504 , \41502 , \41503 );
not \U$41162 ( \41505 , \40884 );
nand \U$41163 ( \41506 , \41504 , \41505 );
not \U$41164 ( \41507 , \41506 );
or \U$41165 ( \41508 , \41500 , \41507 );
not \U$41166 ( \41509 , \40896 );
nand \U$41167 ( \41510 , \41508 , \41509 );
not \U$41168 ( \41511 , \41510 );
or \U$41169 ( \41512 , \41498 , \41511 );
nand \U$41170 ( \41513 , \41512 , \40901 );
nand \U$41171 ( \41514 , \16126 , \40906 );
xor \U$41172 ( \41515 , \41513 , \41514 );
nor \U$41173 ( \41516 , \41515 , \41428 );
buf \U$41174 ( \41517 , \41516 );
not \U$41175 ( \41518 , \16061 );
not \U$41176 ( \41519 , \41506 );
or \U$41177 ( \41520 , \41518 , \41519 );
not \U$41178 ( \41521 , \40890 );
nand \U$41179 ( \41522 , \41520 , \41521 );
nand \U$41180 ( \41523 , \40895 , \16096 );
xor \U$41181 ( \41524 , \41522 , \41523 );
nor \U$41182 ( \41525 , \41524 , \41428 );
buf \U$41183 ( \41526 , \41525 );
nand \U$41184 ( \41527 , \16061 , \41521 );
not \U$41185 ( \41528 , \41527 );
not \U$41186 ( \41529 , \41506 );
or \U$41187 ( \41530 , \41528 , \41529 );
or \U$41188 ( \41531 , \41506 , \41527 );
nand \U$41189 ( \41532 , \41530 , \41531 );
and \U$41190 ( \41533 , \41532 , \41427 );
buf \U$41191 ( \41534 , \41533 );
and \U$41192 ( \41535 , \15230 , \15887 );
not \U$41193 ( \41536 , \41535 );
buf \U$41194 ( \41537 , \41438 );
not \U$41195 ( \41538 , \41537 );
or \U$41196 ( \41539 , \41536 , \41538 );
nand \U$41197 ( \41540 , \41539 , \40876 );
nand \U$41198 ( \41541 , \40878 , \15357 );
xor \U$41199 ( \41542 , \41540 , \41541 );
nor \U$41200 ( \41543 , \41542 , \41345 );
buf \U$41201 ( \41544 , \41543 );
not \U$41202 ( \41545 , \15887 );
not \U$41203 ( \41546 , \41537 );
or \U$41204 ( \41547 , \41545 , \41546 );
not \U$41205 ( \41548 , \40874 );
nand \U$41206 ( \41549 , \41547 , \41548 );
not \U$41207 ( \41550 , \40873 );
nand \U$41208 ( \41551 , \41550 , \15230 );
xor \U$41209 ( \41552 , \41549 , \41551 );
nor \U$41210 ( \41553 , \41552 , \41345 );
buf \U$41211 ( \41554 , \41553 );
and \U$41212 ( \41555 , \41548 , \15887 );
xor \U$41213 ( \41556 , \41537 , \41555 );
and \U$41214 ( \41557 , \41556 , \41427 );
buf \U$41215 ( \41558 , \41557 );
buf \U$41216 ( \41559 , \25536 );
not \U$41217 ( \41560 , \41559 );
not \U$41218 ( \41561 , \25510 );
not \U$41219 ( \41562 , \41561 );
not \U$41220 ( \41563 , \25584 );
buf \U$41221 ( \41564 , \25154 );
buf \U$41222 ( \41565 , \25565 );
and \U$41223 ( \41566 , \41563 , \41564 , \41565 , \25577 );
not \U$41224 ( \41567 , \41566 );
not \U$41225 ( \41568 , \40865 );
buf \U$41226 ( \41569 , \40858 );
not \U$41227 ( \41570 , \41569 );
or \U$41228 ( \41571 , \41568 , \41570 );
buf \U$41229 ( \41572 , \24588 );
nand \U$41230 ( \41573 , \41571 , \41572 );
not \U$41231 ( \41574 , \41573 );
or \U$41232 ( \41575 , \41567 , \41574 );
not \U$41233 ( \41576 , \25577 );
buf \U$41234 ( \41577 , \25587 );
not \U$41235 ( \41578 , \41577 );
not \U$41236 ( \41579 , \41565 );
or \U$41237 ( \41580 , \41578 , \41579 );
buf \U$41238 ( \41581 , \25590 );
nand \U$41239 ( \41582 , \41580 , \41581 );
not \U$41240 ( \41583 , \41582 );
or \U$41241 ( \41584 , \41576 , \41583 );
nand \U$41242 ( \41585 , \41584 , \25591 );
not \U$41243 ( \41586 , \41585 );
nand \U$41244 ( \41587 , \41575 , \41586 );
not \U$41245 ( \41588 , \41587 );
or \U$41246 ( \41589 , \41562 , \41588 );
not \U$41247 ( \41590 , \25601 );
nand \U$41248 ( \41591 , \41589 , \41590 );
not \U$41249 ( \41592 , \41591 );
or \U$41250 ( \41593 , \41560 , \41592 );
buf \U$41251 ( \41594 , \25604 );
nand \U$41252 ( \41595 , \41593 , \41594 );
nand \U$41253 ( \41596 , \25612 , \25607 );
xor \U$41254 ( \41597 , \41595 , \41596 );
nor \U$41255 ( \41598 , \41597 , \41345 );
buf \U$41256 ( \41599 , \41598 );
and \U$41257 ( \41600 , \41563 , \41564 , \41565 );
not \U$41258 ( \41601 , \41600 );
not \U$41259 ( \41602 , \41573 );
or \U$41260 ( \41603 , \41601 , \41602 );
not \U$41261 ( \41604 , \41582 );
nand \U$41262 ( \41605 , \41603 , \41604 );
nand \U$41263 ( \41606 , \25577 , \25591 );
xor \U$41264 ( \41607 , \41605 , \41606 );
not \U$41265 ( \41608 , \41322 );
not \U$41266 ( \41609 , \41608 );
nor \U$41267 ( \41610 , \41607 , \41609 );
buf \U$41268 ( \41611 , \41610 );
not \U$41269 ( \41612 , \25155 );
not \U$41270 ( \41613 , \41573 );
or \U$41271 ( \41614 , \41612 , \41613 );
not \U$41272 ( \41615 , \41577 );
nand \U$41273 ( \41616 , \41614 , \41615 );
nand \U$41274 ( \41617 , \41565 , \41581 );
xor \U$41275 ( \41618 , \41616 , \41617 );
nor \U$41276 ( \41619 , \41618 , \41609 );
buf \U$41277 ( \41620 , \41619 );
not \U$41278 ( \41621 , \41564 );
not \U$41279 ( \41622 , \41573 );
or \U$41280 ( \41623 , \41621 , \41622 );
buf \U$41281 ( \41624 , \25583 );
nand \U$41282 ( \41625 , \41623 , \41624 );
nand \U$41283 ( \41626 , \41563 , \25586 );
xor \U$41284 ( \41627 , \41625 , \41626 );
nor \U$41285 ( \41628 , \41627 , \41323 );
buf \U$41286 ( \41629 , \41628 );
nand \U$41287 ( \41630 , \41624 , \41564 );
xnor \U$41288 ( \41631 , \41630 , \41573 );
not \U$41289 ( \41632 , \41322 );
not \U$41290 ( \41633 , \41632 );
not \U$41291 ( \41634 , \41633 );
and \U$41292 ( \41635 , \41631 , \41634 );
buf \U$41293 ( \41636 , \41635 );
buf \U$41294 ( \41637 , \24580 );
and \U$41295 ( \41638 , \40863 , \41637 );
not \U$41296 ( \41639 , \41638 );
not \U$41297 ( \41640 , \40862 );
buf \U$41298 ( \41641 , \41569 );
not \U$41299 ( \41642 , \41641 );
or \U$41300 ( \41643 , \41640 , \41642 );
not \U$41301 ( \41644 , \24567 );
nand \U$41302 ( \41645 , \41643 , \41644 );
not \U$41303 ( \41646 , \41645 );
or \U$41304 ( \41647 , \41639 , \41646 );
buf \U$41305 ( \41648 , \24579 );
and \U$41306 ( \41649 , \41648 , \41637 );
not \U$41307 ( \41650 , \24583 );
nor \U$41308 ( \41651 , \41649 , \41650 );
nand \U$41309 ( \41652 , \41647 , \41651 );
not \U$41310 ( \41653 , \24586 );
nand \U$41311 ( \41654 , \41653 , \24571 );
xor \U$41312 ( \41655 , \41652 , \41654 );
nor \U$41313 ( \41656 , \41655 , \41428 );
buf \U$41314 ( \41657 , \41656 );
not \U$41315 ( \41658 , \21549 );
not \U$41316 ( \41659 , \41658 );
not \U$41317 ( \41660 , \41645 );
or \U$41318 ( \41661 , \41659 , \41660 );
not \U$41319 ( \41662 , \24573 );
nand \U$41320 ( \41663 , \41661 , \41662 );
not \U$41321 ( \41664 , \20631 );
nand \U$41322 ( \41665 , \41664 , \24578 );
xor \U$41323 ( \41666 , \41663 , \41665 );
nor \U$41324 ( \41667 , \41666 , \41323 );
buf \U$41325 ( \41668 , \41667 );
buf \U$41326 ( \41669 , \40860 );
not \U$41327 ( \41670 , \41669 );
buf \U$41328 ( \41671 , \40861 );
and \U$41329 ( \41672 , \40859 , \41671 );
not \U$41330 ( \41673 , \41672 );
not \U$41331 ( \41674 , \41641 );
or \U$41332 ( \41675 , \41673 , \41674 );
buf \U$41333 ( \41676 , \24551 );
nand \U$41334 ( \41677 , \41675 , \41676 );
not \U$41335 ( \41678 , \41677 );
or \U$41336 ( \41679 , \41670 , \41678 );
nand \U$41337 ( \41680 , \41679 , \24560 );
nand \U$41338 ( \41681 , \24566 , \22870 );
xor \U$41339 ( \41682 , \41680 , \41681 );
nor \U$41340 ( \41683 , \41682 , \41609 );
buf \U$41341 ( \41684 , \41683 );
nand \U$41342 ( \41685 , \41669 , \24560 );
xor \U$41343 ( \41686 , \41677 , \41685 );
nor \U$41344 ( \41687 , \41686 , \41345 );
buf \U$41345 ( \41688 , \41687 );
not \U$41346 ( \41689 , \41671 );
not \U$41347 ( \41690 , \41641 );
or \U$41348 ( \41691 , \41689 , \41690 );
buf \U$41349 ( \41692 , \24546 );
nand \U$41350 ( \41693 , \41691 , \41692 );
not \U$41351 ( \41694 , \23818 );
not \U$41352 ( \41695 , \24548 );
not \U$41353 ( \41696 , \41695 );
or \U$41354 ( \41697 , \41694 , \41696 );
nand \U$41355 ( \41698 , \41697 , \40859 );
xor \U$41356 ( \41699 , \41693 , \41698 );
nor \U$41357 ( \41700 , \41699 , \41323 );
buf \U$41358 ( \41701 , \41700 );
nand \U$41359 ( \41702 , \41692 , \41671 );
not \U$41360 ( \41703 , \41702 );
and \U$41361 ( \41704 , \41641 , \41703 );
not \U$41362 ( \41705 , \41641 );
and \U$41363 ( \41706 , \41705 , \41702 );
nor \U$41364 ( \41707 , \41704 , \41706 );
not \U$41365 ( \41708 , \41707 );
nor \U$41366 ( \41709 , \41708 , \41609 );
buf \U$41367 ( \41710 , \41709 );
not \U$41368 ( \41711 , RIbb2f610_1);
nor \U$41369 ( \41712 , \41711 , \41608 );
not \U$41370 ( \41713 , \41712 );
not \U$41371 ( \41714 , \32726 );
buf \U$41372 ( \41715 , \32687 );
and \U$41373 ( \41716 , \32643 , \41715 );
not \U$41374 ( \41717 , \41716 );
not \U$41375 ( \41718 , \32550 );
not \U$41376 ( \41719 , \40856 );
buf \U$41377 ( \41720 , \40846 );
not \U$41378 ( \41721 , \41720 );
or \U$41379 ( \41722 , \41719 , \41721 );
not \U$41380 ( \41723 , \31737 );
nand \U$41381 ( \41724 , \41722 , \41723 );
not \U$41382 ( \41725 , \41724 );
or \U$41383 ( \41726 , \41718 , \41725 );
not \U$41384 ( \41727 , \32571 );
nand \U$41385 ( \41728 , \41726 , \41727 );
not \U$41386 ( \41729 , \41728 );
or \U$41387 ( \41730 , \41717 , \41729 );
not \U$41388 ( \41731 , \32735 );
nand \U$41389 ( \41732 , \41730 , \41731 );
not \U$41390 ( \41733 , \41732 );
or \U$41391 ( \41734 , \41714 , \41733 );
nand \U$41392 ( \41735 , \41734 , \32738 );
nand \U$41393 ( \41736 , \32742 , \32724 );
not \U$41394 ( \41737 , \41736 );
and \U$41395 ( \41738 , \41735 , \41737 );
not \U$41396 ( \41739 , \41735 );
and \U$41397 ( \41740 , \41739 , \41736 );
nor \U$41398 ( \41741 , \41738 , \41740 );
not \U$41399 ( \41742 , \41345 );
nand \U$41400 ( \41743 , \41741 , \41742 );
nand \U$41401 ( \41744 , \41713 , \41743 );
buf \U$41402 ( \41745 , \41744 );
not \U$41403 ( \41746 , RIbb2f520_3);
nor \U$41404 ( \41747 , \41746 , \41608 );
not \U$41405 ( \41748 , \41747 );
not \U$41406 ( \41749 , \32643 );
not \U$41407 ( \41750 , \41728 );
or \U$41408 ( \41751 , \41749 , \41750 );
not \U$41409 ( \41752 , \32729 );
nand \U$41410 ( \41753 , \41751 , \41752 );
nand \U$41411 ( \41754 , \32734 , \41715 );
not \U$41412 ( \41755 , \41754 );
and \U$41413 ( \41756 , \41753 , \41755 );
not \U$41414 ( \41757 , \41753 );
and \U$41415 ( \41758 , \41757 , \41754 );
nor \U$41416 ( \41759 , \41756 , \41758 );
nand \U$41417 ( \41760 , \41759 , \41427 );
nand \U$41418 ( \41761 , \41748 , \41760 );
buf \U$41419 ( \41762 , \41761 );
nand \U$41420 ( \41763 , \41752 , \32643 );
xnor \U$41421 ( \41764 , \41763 , \41728 );
and \U$41422 ( \41765 , \41608 , \41764 );
not \U$41423 ( \41766 , \41608 );
and \U$41424 ( \41767 , \41766 , RIbb2f4a8_4);
or \U$41425 ( \41768 , \41765 , \41767 );
buf \U$41426 ( \41769 , \41768 );
not \U$41427 ( \41770 , RIbb2f430_5);
nor \U$41428 ( \41771 , \41770 , \41608 );
not \U$41429 ( \41772 , \41771 );
not \U$41430 ( \41773 , \32401 );
buf \U$41431 ( \41774 , \32539 );
buf \U$41432 ( \41775 , \32549 );
and \U$41433 ( \41776 , \41774 , \41775 );
not \U$41434 ( \41777 , \41776 );
not \U$41435 ( \41778 , \41724 );
or \U$41436 ( \41779 , \41777 , \41778 );
not \U$41437 ( \41780 , \32559 );
nand \U$41438 ( \41781 , \41779 , \41780 );
not \U$41439 ( \41782 , \41781 );
or \U$41440 ( \41783 , \41773 , \41782 );
buf \U$41441 ( \41784 , \32564 );
nand \U$41442 ( \41785 , \41783 , \41784 );
nand \U$41443 ( \41786 , \32570 , \32566 );
not \U$41444 ( \41787 , \41786 );
and \U$41445 ( \41788 , \41785 , \41787 );
not \U$41446 ( \41789 , \41785 );
and \U$41447 ( \41790 , \41789 , \41786 );
nor \U$41448 ( \41791 , \41788 , \41790 );
nand \U$41449 ( \41792 , \41791 , \41427 );
nand \U$41450 ( \41793 , \41772 , \41792 );
buf \U$41451 ( \41794 , \41793 );
not \U$41452 ( \41795 , RIbb2f3b8_6);
nor \U$41453 ( \41796 , \41795 , \41344 );
not \U$41454 ( \41797 , \41796 );
nand \U$41455 ( \41798 , \41784 , \32401 );
not \U$41456 ( \41799 , \41798 );
not \U$41457 ( \41800 , \41781 );
or \U$41458 ( \41801 , \41799 , \41800 );
or \U$41459 ( \41802 , \41781 , \41798 );
nand \U$41460 ( \41803 , \41801 , \41802 );
nand \U$41461 ( \41804 , \41803 , \41742 );
nand \U$41462 ( \41805 , \41797 , \41804 );
buf \U$41463 ( \41806 , \41805 );
not \U$41464 ( \41807 , RIbb2f340_7);
nor \U$41465 ( \41808 , \41807 , \41608 );
not \U$41466 ( \41809 , \41808 );
not \U$41467 ( \41810 , \41775 );
not \U$41468 ( \41811 , \41724 );
or \U$41469 ( \41812 , \41810 , \41811 );
not \U$41470 ( \41813 , \32554 );
nand \U$41471 ( \41814 , \41812 , \41813 );
nand \U$41472 ( \41815 , \32558 , \41774 );
not \U$41473 ( \41816 , \41815 );
and \U$41474 ( \41817 , \41814 , \41816 );
not \U$41475 ( \41818 , \41814 );
and \U$41476 ( \41819 , \41818 , \41815 );
nor \U$41477 ( \41820 , \41817 , \41819 );
nand \U$41478 ( \41821 , \41820 , \41427 );
nand \U$41479 ( \41822 , \41809 , \41821 );
buf \U$41480 ( \41823 , \41822 );
and \U$41481 ( \41824 , \41322 , RIbb2f2c8_8);
not \U$41482 ( \41825 , \41322 );
nand \U$41483 ( \41826 , \41813 , \41775 );
not \U$41484 ( \41827 , \41826 );
buf \U$41485 ( \41828 , \41724 );
not \U$41486 ( \41829 , \41828 );
or \U$41487 ( \41830 , \41827 , \41829 );
or \U$41488 ( \41831 , \41828 , \41826 );
nand \U$41489 ( \41832 , \41830 , \41831 );
and \U$41490 ( \41833 , \41825 , \41832 );
or \U$41491 ( \41834 , \41824 , \41833 );
buf \U$41492 ( \41835 , \41834 );
not \U$41493 ( \41836 , RIbb2f250_9);
nor \U$41494 ( \41837 , \41836 , \41608 );
not \U$41495 ( \41838 , \41837 );
buf \U$41496 ( \41839 , \31303 );
not \U$41497 ( \41840 , \41839 );
not \U$41498 ( \41841 , \30838 );
not \U$41499 ( \41842 , \41841 );
not \U$41500 ( \41843 , \40855 );
not \U$41501 ( \41844 , \41843 );
not \U$41502 ( \41845 , \41720 );
or \U$41503 ( \41846 , \41844 , \41845 );
not \U$41504 ( \41847 , \29852 );
nand \U$41505 ( \41848 , \41846 , \41847 );
not \U$41506 ( \41849 , \41848 );
or \U$41507 ( \41850 , \41842 , \41849 );
buf \U$41508 ( \41851 , \31729 );
not \U$41509 ( \41852 , \41851 );
nor \U$41510 ( \41853 , \41852 , \31727 );
nand \U$41511 ( \41854 , \41850 , \41853 );
not \U$41512 ( \41855 , \41854 );
or \U$41513 ( \41856 , \41840 , \41855 );
buf \U$41514 ( \41857 , \31728 );
nand \U$41515 ( \41858 , \41856 , \41857 );
nand \U$41516 ( \41859 , \31721 , \31734 );
not \U$41517 ( \41860 , \41859 );
and \U$41518 ( \41861 , \41858 , \41860 );
not \U$41519 ( \41862 , \41858 );
and \U$41520 ( \41863 , \41862 , \41859 );
nor \U$41521 ( \41864 , \41861 , \41863 );
nand \U$41522 ( \41865 , \41864 , \41427 );
nand \U$41523 ( \41866 , \41838 , \41865 );
buf \U$41524 ( \41867 , \41866 );
not \U$41525 ( \41868 , RIbb2f1d8_10);
nor \U$41526 ( \41869 , \41868 , \41344 );
not \U$41527 ( \41870 , \41869 );
nand \U$41528 ( \41871 , \41857 , \41839 );
not \U$41529 ( \41872 , \41871 );
and \U$41530 ( \41873 , \41854 , \41872 );
not \U$41531 ( \41874 , \41854 );
and \U$41532 ( \41875 , \41874 , \41871 );
nor \U$41533 ( \41876 , \41873 , \41875 );
not \U$41534 ( \41877 , \41345 );
nand \U$41535 ( \41878 , \41876 , \41877 );
nand \U$41536 ( \41879 , \41870 , \41878 );
buf \U$41537 ( \41880 , \41879 );
not \U$41538 ( \41881 , RIbb2f160_11);
nor \U$41539 ( \41882 , \41881 , \41608 );
not \U$41540 ( \41883 , \41882 );
not \U$41541 ( \41884 , \30837 );
not \U$41542 ( \41885 , \41848 );
or \U$41543 ( \41886 , \41884 , \41885 );
buf \U$41544 ( \41887 , \31726 );
nand \U$41545 ( \41888 , \41886 , \41887 );
and \U$41546 ( \41889 , \41851 , \30828 );
and \U$41547 ( \41890 , \41888 , \41889 );
not \U$41548 ( \41891 , \41888 );
not \U$41549 ( \41892 , \41889 );
and \U$41550 ( \41893 , \41891 , \41892 );
nor \U$41551 ( \41894 , \41890 , \41893 );
nand \U$41552 ( \41895 , \41894 , \41427 );
nand \U$41553 ( \41896 , \41883 , \41895 );
buf \U$41554 ( \41897 , \41896 );
and \U$41555 ( \41898 , \41322 , RIbb2f0e8_12);
not \U$41556 ( \41899 , \41322 );
nand \U$41557 ( \41900 , \41887 , \30837 );
not \U$41558 ( \41901 , \41900 );
not \U$41559 ( \41902 , \41848 );
or \U$41560 ( \41903 , \41901 , \41902 );
or \U$41561 ( \41904 , \41900 , \41848 );
nand \U$41562 ( \41905 , \41903 , \41904 );
and \U$41563 ( \41906 , \41899 , \41905 );
or \U$41564 ( \41907 , \41898 , \41906 );
buf \U$41565 ( \41908 , \41907 );
not \U$41566 ( \41909 , RIbb2f070_13);
nor \U$41567 ( \41910 , \41909 , \41608 );
not \U$41568 ( \41911 , \41910 );
not \U$41569 ( \41912 , \40854 );
not \U$41570 ( \41913 , \40853 );
buf \U$41571 ( \41914 , \41720 );
not \U$41572 ( \41915 , \41914 );
or \U$41573 ( \41916 , \41913 , \41915 );
buf \U$41574 ( \41917 , \29364 );
nand \U$41575 ( \41918 , \28924 , \41917 );
nand \U$41576 ( \41919 , \41916 , \41918 );
not \U$41577 ( \41920 , \41919 );
or \U$41578 ( \41921 , \41912 , \41920 );
buf \U$41579 ( \41922 , \29847 );
nand \U$41580 ( \41923 , \41921 , \41922 );
nand \U$41581 ( \41924 , \40849 , \29846 );
not \U$41582 ( \41925 , \41924 );
and \U$41583 ( \41926 , \41923 , \41925 );
not \U$41584 ( \41927 , \41923 );
and \U$41585 ( \41928 , \41927 , \41924 );
nor \U$41586 ( \41929 , \41926 , \41928 );
nand \U$41587 ( \41930 , \41929 , \41608 );
nand \U$41588 ( \41931 , \41911 , \41930 );
buf \U$41589 ( \41932 , \41931 );
not \U$41590 ( \41933 , \41608 );
nand \U$41591 ( \41934 , \40854 , \41922 );
not \U$41592 ( \41935 , \41934 );
not \U$41593 ( \41936 , \41919 );
or \U$41594 ( \41937 , \41935 , \41936 );
or \U$41595 ( \41938 , \41934 , \41919 );
nand \U$41596 ( \41939 , \41937 , \41938 );
not \U$41597 ( \41940 , \41939 );
or \U$41598 ( \41941 , \41933 , \41940 );
nand \U$41599 ( \41942 , \41322 , RIbb2eff8_14);
nand \U$41600 ( \41943 , \41941 , \41942 );
buf \U$41601 ( \41944 , \41943 );
and \U$41602 ( \41945 , \41609 , \2356 );
not \U$41603 ( \41946 , \41609 );
not \U$41604 ( \41947 , \40852 );
not \U$41605 ( \41948 , \41720 );
or \U$41606 ( \41949 , \41947 , \41948 );
buf \U$41607 ( \41950 , \28923 );
nand \U$41608 ( \41951 , \41949 , \41950 );
nand \U$41609 ( \41952 , \28357 , \27928 );
nand \U$41610 ( \41953 , \41952 , \41917 );
xor \U$41611 ( \41954 , \41951 , \41953 );
and \U$41612 ( \41955 , \41946 , \41954 );
nor \U$41613 ( \41956 , \41945 , \41955 );
buf \U$41614 ( \41957 , \41956 );
not \U$41615 ( \41958 , \41608 );
not \U$41616 ( \41959 , \41720 );
nand \U$41617 ( \41960 , \41950 , \40852 );
not \U$41618 ( \41961 , \41960 );
or \U$41619 ( \41962 , \41959 , \41961 );
or \U$41620 ( \41963 , \41914 , \41960 );
nand \U$41621 ( \41964 , \41962 , \41963 );
not \U$41622 ( \41965 , \41964 );
or \U$41623 ( \41966 , \41958 , \41965 );
nand \U$41624 ( \41967 , \41322 , RIbb2ef08_16);
nand \U$41625 ( \41968 , \41966 , \41967 );
buf \U$41626 ( \41969 , \41968 );
not \U$41627 ( \41970 , RIbb2ee90_17);
nor \U$41628 ( \41971 , \41970 , \41608 );
not \U$41629 ( \41972 , \41971 );
nand \U$41630 ( \41973 , \40799 , \40792 );
not \U$41631 ( \41974 , \41973 );
not \U$41632 ( \41975 , \40779 );
not \U$41633 ( \41976 , \35444 );
not \U$41634 ( \41977 , \41976 );
not \U$41635 ( \41978 , \35286 );
not \U$41636 ( \41979 , \37385 );
nand \U$41637 ( \41980 , \40826 , \40726 );
not \U$41638 ( \41981 , \41980 );
or \U$41639 ( \41982 , \41979 , \41981 );
and \U$41640 ( \41983 , \40773 , \40749 );
nand \U$41641 ( \41984 , \41982 , \41983 );
not \U$41642 ( \41985 , \41984 );
or \U$41643 ( \41986 , \41978 , \41985 );
not \U$41644 ( \41987 , \40843 );
not \U$41645 ( \41988 , \40842 );
or \U$41646 ( \41989 , \41987 , \41988 );
not \U$41647 ( \41990 , \40795 );
nand \U$41648 ( \41991 , \41989 , \41990 );
not \U$41649 ( \41992 , \41991 );
nand \U$41650 ( \41993 , \41986 , \41992 );
not \U$41651 ( \41994 , \41993 );
or \U$41652 ( \41995 , \41977 , \41994 );
not \U$41653 ( \41996 , \40787 );
nand \U$41654 ( \41997 , \41995 , \41996 );
not \U$41655 ( \41998 , \41997 );
or \U$41656 ( \41999 , \41975 , \41998 );
nand \U$41657 ( \42000 , \41999 , \40790 );
not \U$41658 ( \42001 , \42000 );
or \U$41659 ( \42002 , \41974 , \42001 );
or \U$41660 ( \42003 , \42000 , \41973 );
nand \U$41661 ( \42004 , \42002 , \42003 );
nand \U$41662 ( \42005 , \42004 , \41427 );
nand \U$41663 ( \42006 , \41972 , \42005 );
buf \U$41664 ( \42007 , \42006 );
not \U$41665 ( \42008 , RIbb2ee18_18);
nor \U$41666 ( \42009 , \42008 , \41344 );
not \U$41667 ( \42010 , \42009 );
nand \U$41668 ( \42011 , \40790 , \40779 );
not \U$41669 ( \42012 , \42011 );
not \U$41670 ( \42013 , \41997 );
or \U$41671 ( \42014 , \42012 , \42013 );
or \U$41672 ( \42015 , \41997 , \42011 );
nand \U$41673 ( \42016 , \42014 , \42015 );
nand \U$41674 ( \42017 , \42016 , \41608 );
nand \U$41675 ( \42018 , \42010 , \42017 );
buf \U$41676 ( \42019 , \42018 );
not \U$41677 ( \42020 , RIbb2eda0_19);
nor \U$41678 ( \42021 , \42020 , \41608 );
not \U$41679 ( \42022 , \42021 );
buf \U$41680 ( \42023 , \35443 );
not \U$41681 ( \42024 , \42023 );
not \U$41682 ( \42025 , \41993 );
or \U$41683 ( \42026 , \42024 , \42025 );
buf \U$41684 ( \42027 , \40784 );
nand \U$41685 ( \42028 , \42026 , \42027 );
not \U$41686 ( \42029 , \40781 );
nand \U$41687 ( \42030 , \42029 , \40786 );
not \U$41688 ( \42031 , \42030 );
and \U$41689 ( \42032 , \42028 , \42031 );
not \U$41690 ( \42033 , \42028 );
and \U$41691 ( \42034 , \42033 , \42030 );
nor \U$41692 ( \42035 , \42032 , \42034 );
nand \U$41693 ( \42036 , \42035 , \41742 );
nand \U$41694 ( \42037 , \42022 , \42036 );
buf \U$41695 ( \42038 , \42037 );
not \U$41696 ( \42039 , RIbb2ed28_20);
nor \U$41697 ( \42040 , \42039 , \41608 );
not \U$41698 ( \42041 , \42040 );
nand \U$41699 ( \42042 , \42027 , \42023 );
not \U$41700 ( \42043 , \42042 );
not \U$41701 ( \42044 , \41993 );
or \U$41702 ( \42045 , \42043 , \42044 );
or \U$41703 ( \42046 , \42042 , \41993 );
nand \U$41704 ( \42047 , \42045 , \42046 );
nand \U$41705 ( \42048 , \41742 , \42047 );
nand \U$41706 ( \42049 , \42041 , \42048 );
buf \U$41707 ( \42050 , \42049 );
not \U$41708 ( \42051 , RIbb2ecb0_21);
nor \U$41709 ( \42052 , \42051 , \41608 );
not \U$41710 ( \42053 , \42052 );
not \U$41711 ( \42054 , \40829 );
buf \U$41712 ( \42055 , \34622 );
and \U$41713 ( \42056 , \42055 , \35152 );
not \U$41714 ( \42057 , \42056 );
not \U$41715 ( \42058 , \41984 );
or \U$41716 ( \42059 , \42057 , \42058 );
not \U$41717 ( \42060 , \40838 );
nand \U$41718 ( \42061 , \42059 , \42060 );
not \U$41719 ( \42062 , \42061 );
or \U$41720 ( \42063 , \42054 , \42062 );
buf \U$41721 ( \42064 , \40841 );
nand \U$41722 ( \42065 , \42063 , \42064 );
nand \U$41723 ( \42066 , \40843 , \41990 );
not \U$41724 ( \42067 , \42066 );
and \U$41725 ( \42068 , \42065 , \42067 );
not \U$41726 ( \42069 , \42065 );
and \U$41727 ( \42070 , \42069 , \42066 );
nor \U$41728 ( \42071 , \42068 , \42070 );
nand \U$41729 ( \42072 , \42071 , \41742 );
nand \U$41730 ( \42073 , \42053 , \42072 );
buf \U$41731 ( \42074 , \42073 );
not \U$41732 ( \42075 , RIbb2ec38_22);
nor \U$41733 ( \42076 , \42075 , \41427 );
not \U$41734 ( \42077 , \42076 );
nand \U$41735 ( \42078 , \42064 , \40829 );
not \U$41736 ( \42079 , \42078 );
and \U$41737 ( \42080 , \42061 , \42079 );
not \U$41738 ( \42081 , \42061 );
and \U$41739 ( \42082 , \42081 , \42078 );
nor \U$41740 ( \42083 , \42080 , \42082 );
nand \U$41741 ( \42084 , \42083 , \41427 );
nand \U$41742 ( \42085 , \42077 , \42084 );
buf \U$41743 ( \42086 , \42085 );
not \U$41744 ( \42087 , RIbb2ebc0_23);
nor \U$41745 ( \42088 , \42087 , \41608 );
not \U$41746 ( \42089 , \42088 );
not \U$41747 ( \42090 , \35152 );
not \U$41748 ( \42091 , \41984 );
or \U$41749 ( \42092 , \42090 , \42091 );
not \U$41750 ( \42093 , \40832 );
nand \U$41751 ( \42094 , \42092 , \42093 );
nand \U$41752 ( \42095 , \42055 , \40837 );
not \U$41753 ( \42096 , \42095 );
and \U$41754 ( \42097 , \42094 , \42096 );
not \U$41755 ( \42098 , \42094 );
and \U$41756 ( \42099 , \42098 , \42095 );
nor \U$41757 ( \42100 , \42097 , \42099 );
nand \U$41758 ( \42101 , \42100 , \41427 );
nand \U$41759 ( \42102 , \42089 , \42101 );
buf \U$41760 ( \42103 , \42102 );
not \U$41761 ( \42104 , RIbb2eb48_24);
nor \U$41762 ( \42105 , \42104 , \41427 );
not \U$41763 ( \42106 , \42105 );
nand \U$41764 ( \42107 , \42093 , \35152 );
not \U$41765 ( \42108 , \42107 );
and \U$41766 ( \42109 , \41984 , \42108 );
not \U$41767 ( \42110 , \41984 );
and \U$41768 ( \42111 , \42110 , \42107 );
nor \U$41769 ( \42112 , \42109 , \42111 );
not \U$41770 ( \42113 , \41345 );
nand \U$41771 ( \42114 , \42112 , \42113 );
nand \U$41772 ( \42115 , \42106 , \42114 );
buf \U$41773 ( \42116 , \42115 );
not \U$41774 ( \42117 , RIbb2ead0_25);
nor \U$41775 ( \42118 , \42117 , \41344 );
not \U$41776 ( \42119 , \42118 );
nand \U$41777 ( \42120 , \40771 , \37383 );
not \U$41778 ( \42121 , \42120 );
not \U$41779 ( \42122 , \37375 );
not \U$41780 ( \42123 , \37345 );
not \U$41781 ( \42124 , \37248 );
not \U$41782 ( \42125 , \41980 );
or \U$41783 ( \42126 , \42124 , \42125 );
not \U$41784 ( \42127 , \40747 );
nand \U$41785 ( \42128 , \42126 , \42127 );
not \U$41786 ( \42129 , \42128 );
or \U$41787 ( \42130 , \42123 , \42129 );
not \U$41788 ( \42131 , \40760 );
nand \U$41789 ( \42132 , \42130 , \42131 );
not \U$41790 ( \42133 , \42132 );
or \U$41791 ( \42134 , \42122 , \42133 );
nand \U$41792 ( \42135 , \42134 , \40765 );
not \U$41793 ( \42136 , \42135 );
or \U$41794 ( \42137 , \42121 , \42136 );
or \U$41795 ( \42138 , \42135 , \42120 );
nand \U$41796 ( \42139 , \42137 , \42138 );
nand \U$41797 ( \42140 , \42139 , \41427 );
nand \U$41798 ( \42141 , \42119 , \42140 );
buf \U$41799 ( \42142 , \42141 );
not \U$41800 ( \42143 , RIbb2ea58_26);
nor \U$41801 ( \42144 , \42143 , \41608 );
not \U$41802 ( \42145 , \42144 );
and \U$41803 ( \42146 , \40765 , \37375 );
xor \U$41804 ( \42147 , \42146 , \42132 );
nand \U$41805 ( \42148 , \42147 , \42113 );
nand \U$41806 ( \42149 , \42145 , \42148 );
buf \U$41807 ( \42150 , \42149 );
not \U$41808 ( \42151 , RIbb2e9e0_27);
nor \U$41809 ( \42152 , \42151 , \41427 );
not \U$41810 ( \42153 , \42152 );
nand \U$41811 ( \42154 , \40759 , \37331 );
not \U$41812 ( \42155 , \42154 );
not \U$41813 ( \42156 , \37344 );
not \U$41814 ( \42157 , \42128 );
or \U$41815 ( \42158 , \42156 , \42157 );
not \U$41816 ( \42159 , \40754 );
nand \U$41817 ( \42160 , \42158 , \42159 );
not \U$41818 ( \42161 , \42160 );
or \U$41819 ( \42162 , \42155 , \42161 );
or \U$41820 ( \42163 , \42160 , \42154 );
nand \U$41821 ( \42164 , \42162 , \42163 );
nand \U$41822 ( \42165 , \42164 , \41877 );
nand \U$41823 ( \42166 , \42153 , \42165 );
buf \U$41824 ( \42167 , \42166 );
not \U$41825 ( \42168 , RIbb2e968_28);
nor \U$41826 ( \42169 , \42168 , \41427 );
not \U$41827 ( \42170 , \42169 );
nand \U$41828 ( \42171 , \37344 , \42159 );
xnor \U$41829 ( \42172 , \42171 , \42128 );
nand \U$41830 ( \42173 , \42113 , \42172 );
nand \U$41831 ( \42174 , \42170 , \42173 );
buf \U$41832 ( \42175 , \42174 );
not \U$41833 ( \42176 , RIbb2e8f0_29);
nor \U$41834 ( \42177 , \42176 , \41344 );
not \U$41835 ( \42178 , \42177 );
nand \U$41836 ( \42179 , \40746 , \37230 );
not \U$41837 ( \42180 , \42179 );
not \U$41838 ( \42181 , \37247 );
not \U$41839 ( \42182 , \37034 );
not \U$41840 ( \42183 , \41980 );
or \U$41841 ( \42184 , \42182 , \42183 );
nand \U$41842 ( \42185 , \42184 , \40735 );
not \U$41843 ( \42186 , \42185 );
or \U$41844 ( \42187 , \42181 , \42186 );
nand \U$41845 ( \42188 , \42187 , \40742 );
not \U$41846 ( \42189 , \42188 );
or \U$41847 ( \42190 , \42180 , \42189 );
or \U$41848 ( \42191 , \42188 , \42179 );
nand \U$41849 ( \42192 , \42190 , \42191 );
nand \U$41850 ( \42193 , \42192 , \41427 );
nand \U$41851 ( \42194 , \42178 , \42193 );
buf \U$41852 ( \42195 , \42194 );
not \U$41853 ( \42196 , RIbb2e878_30);
nor \U$41854 ( \42197 , \42196 , \41427 );
not \U$41855 ( \42198 , \42197 );
nand \U$41856 ( \42199 , \37247 , \40742 );
not \U$41857 ( \42200 , \42199 );
not \U$41858 ( \42201 , \42185 );
or \U$41859 ( \42202 , \42200 , \42201 );
or \U$41860 ( \42203 , \42185 , \42199 );
nand \U$41861 ( \42204 , \42202 , \42203 );
nand \U$41862 ( \42205 , \42204 , \42113 );
nand \U$41863 ( \42206 , \42198 , \42205 );
buf \U$41864 ( \42207 , \42206 );
not \U$41865 ( \42208 , RIbb2e800_31);
nor \U$41866 ( \42209 , \42208 , \41427 );
not \U$41867 ( \42210 , \42209 );
nand \U$41868 ( \42211 , \37033 , \40732 );
not \U$41869 ( \42212 , \42211 );
not \U$41870 ( \42213 , \36860 );
not \U$41871 ( \42214 , \41980 );
or \U$41872 ( \42215 , \42213 , \42214 );
buf \U$41873 ( \42216 , \40730 );
nand \U$41874 ( \42217 , \42215 , \42216 );
not \U$41875 ( \42218 , \42217 );
or \U$41876 ( \42219 , \42212 , \42218 );
or \U$41877 ( \42220 , \42217 , \42211 );
nand \U$41878 ( \42221 , \42219 , \42220 );
nand \U$41879 ( \42222 , \42221 , \41742 );
nand \U$41880 ( \42223 , \42210 , \42222 );
buf \U$41881 ( \42224 , \42223 );
not \U$41882 ( \42225 , RIbb2e788_32);
nor \U$41883 ( \42226 , \42225 , \41608 );
not \U$41884 ( \42227 , \42226 );
nand \U$41885 ( \42228 , \42216 , \36860 );
not \U$41886 ( \42229 , \42228 );
not \U$41887 ( \42230 , \41980 );
or \U$41888 ( \42231 , \42229 , \42230 );
or \U$41889 ( \42232 , \42228 , \41980 );
nand \U$41890 ( \42233 , \42231 , \42232 );
nand \U$41891 ( \42234 , \42233 , \41877 );
nand \U$41892 ( \42235 , \42227 , \42234 );
buf \U$41893 ( \42236 , \42235 );
not \U$41894 ( \42237 , RIbb2e710_33);
nor \U$41895 ( \42238 , \42237 , \41427 );
not \U$41896 ( \42239 , \42238 );
not \U$41897 ( \42240 , \40678 );
not \U$41898 ( \42241 , \40724 );
not \U$41899 ( \42242 , \42241 );
buf \U$41900 ( \42243 , \40565 );
not \U$41901 ( \42244 , \42243 );
or \U$41902 ( \42245 , \42242 , \42244 );
not \U$41903 ( \42246 , \40814 );
nand \U$41904 ( \42247 , \42245 , \42246 );
not \U$41905 ( \42248 , \42247 );
or \U$41906 ( \42249 , \42240 , \42248 );
nand \U$41907 ( \42250 , \42249 , \40819 );
nand \U$41908 ( \42251 , \40824 , \40611 );
not \U$41909 ( \42252 , \42251 );
and \U$41910 ( \42253 , \42250 , \42252 );
not \U$41911 ( \42254 , \42250 );
and \U$41912 ( \42255 , \42254 , \42251 );
nor \U$41913 ( \42256 , \42253 , \42255 );
nand \U$41914 ( \42257 , \42256 , \42113 );
nand \U$41915 ( \42258 , \42239 , \42257 );
buf \U$41916 ( \42259 , \42258 );
not \U$41917 ( \42260 , RIbb2e698_34);
nor \U$41918 ( \42261 , \42260 , \41427 );
not \U$41919 ( \42262 , \42261 );
nand \U$41920 ( \42263 , \40819 , \40678 );
not \U$41921 ( \42264 , \42263 );
and \U$41922 ( \42265 , \42247 , \42264 );
not \U$41923 ( \42266 , \42247 );
and \U$41924 ( \42267 , \42266 , \42263 );
nor \U$41925 ( \42268 , \42265 , \42267 );
nand \U$41926 ( \42269 , \42268 , \41877 );
nand \U$41927 ( \42270 , \42262 , \42269 );
buf \U$41928 ( \42271 , \42270 );
not \U$41929 ( \42272 , RIbb2e620_35);
nor \U$41930 ( \42273 , \42272 , \41427 );
not \U$41931 ( \42274 , \42273 );
not \U$41932 ( \42275 , \40723 );
not \U$41933 ( \42276 , \42243 );
or \U$41934 ( \42277 , \42275 , \42276 );
not \U$41935 ( \42278 , \40809 );
nand \U$41936 ( \42279 , \42277 , \42278 );
nand \U$41937 ( \42280 , \40813 , \40807 );
not \U$41938 ( \42281 , \42280 );
and \U$41939 ( \42282 , \42279 , \42281 );
not \U$41940 ( \42283 , \42279 );
and \U$41941 ( \42284 , \42283 , \42280 );
nor \U$41942 ( \42285 , \42282 , \42284 );
nand \U$41943 ( \42286 , \42285 , \41877 );
nand \U$41944 ( \42287 , \42274 , \42286 );
buf \U$41945 ( \42288 , \42287 );
not \U$41946 ( \42289 , RIbb2e5a8_36);
nor \U$41947 ( \42290 , \42289 , \41427 );
not \U$41948 ( \42291 , \42290 );
nand \U$41949 ( \42292 , \42278 , \40723 );
not \U$41950 ( \42293 , \42292 );
and \U$41951 ( \42294 , \42243 , \42293 );
not \U$41952 ( \42295 , \42243 );
and \U$41953 ( \42296 , \42295 , \42292 );
nor \U$41954 ( \42297 , \42294 , \42296 );
nand \U$41955 ( \42298 , \42297 , \42113 );
nand \U$41956 ( \42299 , \42291 , \42298 );
buf \U$41957 ( \42300 , \42299 );
not \U$41958 ( \42301 , RIbb2e530_37);
nor \U$41959 ( \42302 , \42301 , \41608 );
not \U$41960 ( \42303 , \42302 );
not \U$41961 ( \42304 , \38394 );
not \U$41962 ( \42305 , \40562 );
buf \U$41963 ( \42306 , \40560 );
not \U$41964 ( \42307 , \42306 );
or \U$41965 ( \42308 , \42305 , \42307 );
not \U$41966 ( \42309 , \38657 );
nand \U$41967 ( \42310 , \42308 , \42309 );
not \U$41968 ( \42311 , \42310 );
or \U$41969 ( \42312 , \42304 , \42311 );
nand \U$41970 ( \42313 , \42312 , \38662 );
not \U$41971 ( \42314 , \38755 );
nand \U$41972 ( \42315 , \42314 , \38753 );
not \U$41973 ( \42316 , \42315 );
and \U$41974 ( \42317 , \42313 , \42316 );
not \U$41975 ( \42318 , \42313 );
and \U$41976 ( \42319 , \42318 , \42315 );
nor \U$41977 ( \42320 , \42317 , \42319 );
nand \U$41978 ( \42321 , \42320 , \41877 );
nand \U$41979 ( \42322 , \42303 , \42321 );
buf \U$41980 ( \42323 , \42322 );
not \U$41981 ( \42324 , RIbb2e4b8_38);
nor \U$41982 ( \42325 , \42324 , \41427 );
not \U$41983 ( \42326 , \42325 );
nand \U$41984 ( \42327 , \38662 , \38394 );
not \U$41985 ( \42328 , \42327 );
not \U$41986 ( \42329 , \42310 );
or \U$41987 ( \42330 , \42328 , \42329 );
or \U$41988 ( \42331 , \42310 , \42327 );
nand \U$41989 ( \42332 , \42330 , \42331 );
nand \U$41990 ( \42333 , \41742 , \42332 );
nand \U$41991 ( \42334 , \42326 , \42333 );
buf \U$41992 ( \42335 , \42334 );
not \U$41993 ( \42336 , RIbb2e440_39);
nor \U$41994 ( \42337 , \42336 , \41608 );
not \U$41995 ( \42338 , \42337 );
not \U$41996 ( \42339 , \40561 );
not \U$41997 ( \42340 , \42306 );
or \U$41998 ( \42341 , \42339 , \42340 );
buf \U$41999 ( \42342 , \38633 );
not \U$42000 ( \42343 , \42342 );
nand \U$42001 ( \42344 , \42341 , \42343 );
nand \U$42002 ( \42345 , \38656 , \38652 );
not \U$42003 ( \42346 , \42345 );
and \U$42004 ( \42347 , \42344 , \42346 );
not \U$42005 ( \42348 , \42344 );
and \U$42006 ( \42349 , \42348 , \42345 );
nor \U$42007 ( \42350 , \42347 , \42349 );
nand \U$42008 ( \42351 , \42350 , \42113 );
nand \U$42009 ( \42352 , \42338 , \42351 );
buf \U$42010 ( \42353 , \42352 );
not \U$42011 ( \42354 , RIbb2e3c8_40);
nor \U$42012 ( \42355 , \42354 , \41427 );
not \U$42013 ( \42356 , \42355 );
nand \U$42014 ( \42357 , \42343 , \40561 );
not \U$42015 ( \42358 , \42357 );
and \U$42016 ( \42359 , \42306 , \42358 );
not \U$42017 ( \42360 , \42306 );
and \U$42018 ( \42361 , \42360 , \42357 );
nor \U$42019 ( \42362 , \42359 , \42361 );
nand \U$42020 ( \42363 , \42362 , \42113 );
nand \U$42021 ( \42364 , \42356 , \42363 );
buf \U$42022 ( \42365 , \42364 );
not \U$42023 ( \42366 , RIbb2e350_41);
nor \U$42024 ( \42367 , \42366 , \41427 );
not \U$42025 ( \42368 , \42367 );
buf \U$42026 ( \42369 , \39397 );
not \U$42027 ( \42370 , \42369 );
not \U$42028 ( \42371 , \39359 );
and \U$42029 ( \42372 , \40553 , \40558 );
or \U$42030 ( \42373 , \42372 , \39805 );
not \U$42031 ( \42374 , \42373 );
or \U$42032 ( \42375 , \42371 , \42374 );
not \U$42033 ( \42376 , \39815 );
nand \U$42034 ( \42377 , \42375 , \42376 );
not \U$42035 ( \42378 , \42377 );
or \U$42036 ( \42379 , \42370 , \42378 );
nand \U$42037 ( \42380 , \42379 , \39808 );
nand \U$42038 ( \42381 , \39819 , \39822 );
not \U$42039 ( \42382 , \42381 );
and \U$42040 ( \42383 , \42380 , \42382 );
not \U$42041 ( \42384 , \42380 );
and \U$42042 ( \42385 , \42384 , \42381 );
nor \U$42043 ( \42386 , \42383 , \42385 );
nand \U$42044 ( \42387 , \42386 , \41427 );
nand \U$42045 ( \42388 , \42368 , \42387 );
buf \U$42046 ( \42389 , \42388 );
and \U$42047 ( \42390 , \41322 , RIbb2e2d8_42);
not \U$42048 ( \42391 , \41322 );
nand \U$42049 ( \42392 , \39808 , \42369 );
not \U$42050 ( \42393 , \42392 );
and \U$42051 ( \42394 , \42377 , \42393 );
not \U$42052 ( \42395 , \42377 );
and \U$42053 ( \42396 , \42395 , \42392 );
nor \U$42054 ( \42397 , \42394 , \42396 );
and \U$42055 ( \42398 , \42391 , \42397 );
or \U$42056 ( \42399 , \42390 , \42398 );
buf \U$42057 ( \42400 , \42399 );
and \U$42058 ( \42401 , \41322 , RIbb2e260_43);
not \U$42059 ( \42402 , \41322 );
not \U$42060 ( \42403 , \39357 );
not \U$42061 ( \42404 , \42373 );
or \U$42062 ( \42405 , \42403 , \42404 );
not \U$42063 ( \42406 , \39811 );
nand \U$42064 ( \42407 , \42405 , \42406 );
nand \U$42065 ( \42408 , \39814 , \39252 );
not \U$42066 ( \42409 , \42408 );
and \U$42067 ( \42410 , \42407 , \42409 );
not \U$42068 ( \42411 , \42407 );
and \U$42069 ( \42412 , \42411 , \42408 );
nor \U$42070 ( \42413 , \42410 , \42412 );
and \U$42071 ( \42414 , \42402 , \42413 );
or \U$42072 ( \42415 , \42401 , \42414 );
buf \U$42073 ( \42416 , \42415 );
not \U$42074 ( \42417 , \41608 );
and \U$42075 ( \42418 , \42406 , \39357 );
xor \U$42076 ( \42419 , \42373 , \42418 );
not \U$42077 ( \42420 , \42419 );
or \U$42078 ( \42421 , \42417 , \42420 );
nand \U$42079 ( \42422 , \41609 , RIbb2e1e8_44);
nand \U$42080 ( \42423 , \42421 , \42422 );
buf \U$42081 ( \42424 , \42423 );
and \U$42082 ( \42425 , \41322 , RIbb2e170_45);
not \U$42083 ( \42426 , \41322 );
not \U$42084 ( \42427 , \39619 );
not \U$42085 ( \42428 , \40557 );
not \U$42086 ( \42429 , \42428 );
not \U$42087 ( \42430 , \40553 );
or \U$42088 ( \42431 , \42429 , \42430 );
not \U$42089 ( \42432 , \39796 );
nand \U$42090 ( \42433 , \42431 , \42432 );
not \U$42091 ( \42434 , \42433 );
or \U$42092 ( \42435 , \42427 , \42434 );
nand \U$42093 ( \42436 , \42435 , \39800 );
nand \U$42094 ( \42437 , \39518 , \39804 );
not \U$42095 ( \42438 , \42437 );
and \U$42096 ( \42439 , \42436 , \42438 );
not \U$42097 ( \42440 , \42436 );
and \U$42098 ( \42441 , \42440 , \42437 );
nor \U$42099 ( \42442 , \42439 , \42441 );
and \U$42100 ( \42443 , \42426 , \42442 );
or \U$42101 ( \42444 , \42425 , \42443 );
buf \U$42102 ( \42445 , \42444 );
not \U$42103 ( \42446 , \41608 );
nand \U$42104 ( \42447 , \39619 , \39800 );
not \U$42105 ( \42448 , \42447 );
not \U$42106 ( \42449 , \42433 );
or \U$42107 ( \42450 , \42448 , \42449 );
or \U$42108 ( \42451 , \42447 , \42433 );
nand \U$42109 ( \42452 , \42450 , \42451 );
not \U$42110 ( \42453 , \42452 );
or \U$42111 ( \42454 , \42446 , \42453 );
nand \U$42112 ( \42455 , \41609 , RIbb2e0f8_46);
nand \U$42113 ( \42456 , \42454 , \42455 );
buf \U$42114 ( \42457 , \42456 );
not \U$42115 ( \42458 , \41608 );
nand \U$42116 ( \42459 , \39795 , \40555 );
not \U$42117 ( \42460 , \42459 );
not \U$42118 ( \42461 , \40556 );
not \U$42119 ( \42462 , \40553 );
or \U$42120 ( \42463 , \42461 , \42462 );
not \U$42121 ( \42464 , \39792 );
nand \U$42122 ( \42465 , \42463 , \42464 );
not \U$42123 ( \42466 , \42465 );
or \U$42124 ( \42467 , \42460 , \42466 );
or \U$42125 ( \42468 , \42459 , \42465 );
nand \U$42126 ( \42469 , \42467 , \42468 );
not \U$42127 ( \42470 , \42469 );
or \U$42128 ( \42471 , \42458 , \42470 );
nand \U$42129 ( \42472 , RIbb2e080_47, \41345 );
nand \U$42130 ( \42473 , \42471 , \42472 );
buf \U$42131 ( \42474 , \42473 );
and \U$42132 ( \42475 , \41322 , RIbb2e008_48);
not \U$42133 ( \42476 , \41322 );
nand \U$42134 ( \42477 , \42464 , \40556 );
not \U$42135 ( \42478 , \42477 );
and \U$42136 ( \42479 , \40553 , \42478 );
not \U$42137 ( \42480 , \40553 );
and \U$42138 ( \42481 , \42480 , \42477 );
nor \U$42139 ( \42482 , \42479 , \42481 );
and \U$42140 ( \42483 , \42476 , \42482 );
or \U$42141 ( \42484 , \42475 , \42483 );
buf \U$42142 ( \42485 , \42484 );
and \U$42143 ( \42486 , \41345 , RIbb2df90_49);
not \U$42144 ( \42487 , \41345 );
nand \U$42145 ( \42488 , \39911 , \40552 );
xnor \U$42146 ( \42489 , \40549 , \42488 );
and \U$42147 ( \42490 , \42487 , \42489 );
or \U$42148 ( \42491 , \42486 , \42490 );
buf \U$42149 ( \42492 , \42491 );
nand \U$42150 ( \42493 , \40548 , \40011 );
xnor \U$42151 ( \42494 , \40544 , \42493 );
and \U$42152 ( \42495 , \41344 , \42494 );
not \U$42153 ( \42496 , \41344 );
and \U$42154 ( \42497 , \42496 , RIbb2df18_50);
or \U$42155 ( \42498 , \42495 , \42497 );
buf \U$42156 ( \42499 , \42498 );
not \U$42157 ( \42500 , \40535 );
not \U$42158 ( \42501 , \40493 );
or \U$42159 ( \42502 , \42500 , \42501 );
not \U$42160 ( \42503 , \40539 );
nand \U$42161 ( \42504 , \42502 , \42503 );
nand \U$42162 ( \42505 , \40542 , \40520 );
xnor \U$42163 ( \42506 , \42504 , \42505 );
and \U$42164 ( \42507 , \41344 , \42506 );
not \U$42165 ( \42508 , \41344 );
and \U$42166 ( \42509 , \42508 , RIbb2dea0_51);
or \U$42167 ( \42510 , \42507 , \42509 );
buf \U$42168 ( \42511 , \42510 );
not \U$42169 ( \42512 , \41608 );
nand \U$42170 ( \42513 , \42503 , \40535 );
xnor \U$42171 ( \42514 , \40493 , \42513 );
not \U$42172 ( \42515 , \42514 );
or \U$42173 ( \42516 , \42512 , \42515 );
nand \U$42174 ( \42517 , \41322 , RIbb2de28_52);
nand \U$42175 ( \42518 , \42516 , \42517 );
buf \U$42176 ( \42519 , \42518 );
not \U$42177 ( \42520 , \41608 );
not \U$42178 ( \42521 , \40488 );
nand \U$42179 ( \42522 , \40492 , \40175 );
not \U$42180 ( \42523 , \42522 );
or \U$42181 ( \42524 , \42521 , \42523 );
or \U$42182 ( \42525 , \40488 , \42522 );
nand \U$42183 ( \42526 , \42524 , \42525 );
not \U$42184 ( \42527 , \42526 );
or \U$42185 ( \42528 , \42520 , \42527 );
not \U$42186 ( \42529 , \41322 );
not \U$42187 ( \42530 , \42529 );
nand \U$42188 ( \42531 , RIbb2ddb0_53, \42530 );
nand \U$42189 ( \42532 , \42528 , \42531 );
buf \U$42190 ( \42533 , \42532 );
nand \U$42191 ( \42534 , \40487 , \40485 );
xnor \U$42192 ( \42535 , \42534 , \40474 );
and \U$42193 ( \42536 , \41344 , \42535 );
not \U$42194 ( \42537 , \41344 );
and \U$42195 ( \42538 , \42537 , RIbb2dd38_54);
or \U$42196 ( \42539 , \42536 , \42538 );
buf \U$42197 ( \42540 , \42539 );
endmodule

