//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RIb559478_125,RIb55f760_53,RIb55f6e8_54,RIb55f670_55,RIb5594f0_124,RIb559388_127,RIb55f850_51,RIb55f7d8_52,RIb559400_126,
        RIb559310_128,RIb55f8c8_50,RIb55f940_49,RIb55da50_115,RIb55f2b0_63,RIb55f238_64,RIb55dac8_114,RIb55d960_117,RIb55f3a0_61,RIb55f328_62,
        RIb55d9d8_116,RIb55d870_119,RIb55f490_59,RIb55f418_60,RIb55d8e8_118,RIb55d780_121,RIb55f580_57,RIb55f508_58,RIb55d7f8_120,RIb55d690_123,
        RIb55f5f8_56,RIb55d708_122,RIb55db40_113,RIb55dbb8_112,RIb55fa30_47,RIb55f9b8_48,RIb55dc30_111,RIb55dca8_110,RIb55fb20_45,RIb55faa8_46,
        RIb55dd20_109,RIb55dd98_108,RIb55fc10_43,RIb55fb98_44,RIb55de10_107,RIb55fc88_42,RIb55fd00_41,RIb55de88_106,RIb55df00_105,RIb55df78_104,
        RIb55fdf0_39,RIb55fd78_40,RIb55dff0_103,RIb55e068_102,RIb55fee0_37,RIb55fe68_38,RIb55e0e0_101,RIb55e158_100,RIb55ffd0_35,RIb55ff58_36,
        RIb55e1d0_99,RIb55e248_98,RIb5600c0_33,RIb560048_34,RIb55e2c0_97,RIb55e338_96,RIb5601b0_31,RIb560138_32,RIb55e3b0_95,RIb55e428_94,
        RIb5602a0_29,RIb560228_30,RIb55e4a0_93,RIb560318_28,RIb560390_27,RIb55e518_92,RIb55e590_91,RIb55e608_90,RIb560480_25,RIb560408_26,
        RIb55e680_89,RIb55e6f8_88,RIb560570_23,RIb5604f8_24,RIb55e770_87,RIb55e7e8_86,RIb560660_21,RIb5605e8_22,RIb55e860_85,RIb55e8d8_84,
        RIb560750_19,RIb5606d8_20,RIb55e950_83,RIb55e9c8_82,RIb560840_17,RIb5607c8_18,RIb55ea40_81,RIb5608b8_16,RIb560930_15,RIb55eab8_80,
        RIb55eb30_79,RIb5609a8_14,RIb560a20_13,RIb55eba8_78,RIb55ec20_77,RIb560a98_12,RIb560b10_11,RIb55ec98_76,RIb55ed10_75,RIb55ed88_74,
        RIb560c00_9,RIb560b88_10,RIb55ee00_73,RIb560c78_8,RIb560cf0_7,RIb55ee78_72,RIb55eef0_71,RIb55ef68_70,RIb560de0_5,RIb560d68_6,
        RIb55efe0_69,RIb55f058_68,RIb560ed0_3,RIb560e58_4,RIb55f0d0_67,RIb560f48_2,RIb560fc0_1,RIb55f148_66,RIb55f1c0_65,R_81_7e072f0);
input RIb559478_125,RIb55f760_53,RIb55f6e8_54,RIb55f670_55,RIb5594f0_124,RIb559388_127,RIb55f850_51,RIb55f7d8_52,RIb559400_126,
        RIb559310_128,RIb55f8c8_50,RIb55f940_49,RIb55da50_115,RIb55f2b0_63,RIb55f238_64,RIb55dac8_114,RIb55d960_117,RIb55f3a0_61,RIb55f328_62,
        RIb55d9d8_116,RIb55d870_119,RIb55f490_59,RIb55f418_60,RIb55d8e8_118,RIb55d780_121,RIb55f580_57,RIb55f508_58,RIb55d7f8_120,RIb55d690_123,
        RIb55f5f8_56,RIb55d708_122,RIb55db40_113,RIb55dbb8_112,RIb55fa30_47,RIb55f9b8_48,RIb55dc30_111,RIb55dca8_110,RIb55fb20_45,RIb55faa8_46,
        RIb55dd20_109,RIb55dd98_108,RIb55fc10_43,RIb55fb98_44,RIb55de10_107,RIb55fc88_42,RIb55fd00_41,RIb55de88_106,RIb55df00_105,RIb55df78_104,
        RIb55fdf0_39,RIb55fd78_40,RIb55dff0_103,RIb55e068_102,RIb55fee0_37,RIb55fe68_38,RIb55e0e0_101,RIb55e158_100,RIb55ffd0_35,RIb55ff58_36,
        RIb55e1d0_99,RIb55e248_98,RIb5600c0_33,RIb560048_34,RIb55e2c0_97,RIb55e338_96,RIb5601b0_31,RIb560138_32,RIb55e3b0_95,RIb55e428_94,
        RIb5602a0_29,RIb560228_30,RIb55e4a0_93,RIb560318_28,RIb560390_27,RIb55e518_92,RIb55e590_91,RIb55e608_90,RIb560480_25,RIb560408_26,
        RIb55e680_89,RIb55e6f8_88,RIb560570_23,RIb5604f8_24,RIb55e770_87,RIb55e7e8_86,RIb560660_21,RIb5605e8_22,RIb55e860_85,RIb55e8d8_84,
        RIb560750_19,RIb5606d8_20,RIb55e950_83,RIb55e9c8_82,RIb560840_17,RIb5607c8_18,RIb55ea40_81,RIb5608b8_16,RIb560930_15,RIb55eab8_80,
        RIb55eb30_79,RIb5609a8_14,RIb560a20_13,RIb55eba8_78,RIb55ec20_77,RIb560a98_12,RIb560b10_11,RIb55ec98_76,RIb55ed10_75,RIb55ed88_74,
        RIb560c00_9,RIb560b88_10,RIb55ee00_73,RIb560c78_8,RIb560cf0_7,RIb55ee78_72,RIb55eef0_71,RIb55ef68_70,RIb560de0_5,RIb560d68_6,
        RIb55efe0_69,RIb55f058_68,RIb560ed0_3,RIb560e58_4,RIb55f0d0_67,RIb560f48_2,RIb560fc0_1,RIb55f148_66,RIb55f1c0_65;
output R_81_7e072f0;

wire \130 , \131_N$1 , \132_ZERO , \133_ONE , \134 , \135 , \136 , \137 , \138 ,
         \139 , \140 , \141 , \142 , \143 , \144 , \145 , \146 , \147 , \148 ,
         \149 , \150 , \151 , \152 , \153 , \154 , \155 , \156 , \157 , \158 ,
         \159 , \160 , \161 , \162 , \163 , \164 , \165 , \166 , \167 , \168 ,
         \169 , \170 , \171 , \172 , \173 , \174 , \175 , \176 , \177 , \178 ,
         \179 , \180 , \181 , \182 , \183 , \184 , \185 , \186 , \187 , \188 ,
         \189 , \190 , \191 , \192 , \193 , \194 , \195 , \196 , \197 , \198 ,
         \199 , \200 , \201 , \202 , \203 , \204 , \205 , \206 , \207 , \208 ,
         \209 , \210 , \211 , \212 , \213 , \214 , \215 , \216 , \217 , \218 ,
         \219 , \220 , \221 , \222 , \223 , \224 , \225 , \226 , \227 , \228 ,
         \229 , \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 , \238 ,
         \239 , \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 , \248 ,
         \249 , \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 , \258 ,
         \259 , \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 , \268 ,
         \269 , \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 , \278 ,
         \279 , \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 , \288 ,
         \289 , \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 , \298 ,
         \299 , \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 , \308 ,
         \309 , \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 , \318 ,
         \319 , \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 , \328 ,
         \329 , \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 , \338 ,
         \339 , \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 , \348 ,
         \349 , \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 ,
         \359 , \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 ,
         \369 , \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 ,
         \379 , \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 ,
         \389 , \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 ,
         \399 , \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 ,
         \409 , \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 ,
         \419 , \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 ,
         \429 , \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 ,
         \439 , \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 ,
         \449 , \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 ,
         \459 , \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 ,
         \469 , \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 ,
         \479 , \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 ,
         \489 , \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 ,
         \499 , \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 ,
         \509 , \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 ,
         \519 , \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 ,
         \529 , \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 ,
         \539 , \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 ,
         \549 , \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 ,
         \559 , \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 ,
         \569 , \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 ,
         \579 , \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 ,
         \589 , \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 ,
         \599 , \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 ,
         \609 , \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 ,
         \619 , \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 ,
         \629 , \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 ,
         \639 , \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 ,
         \649 , \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 ,
         \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 ,
         \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 ,
         \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 ,
         \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 ,
         \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 ,
         \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 ,
         \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 ,
         \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 ,
         \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 ,
         \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 ,
         \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 ,
         \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 ,
         \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 ,
         \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 ,
         \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 ,
         \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 ,
         \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 ,
         \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 ,
         \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 ,
         \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 ,
         \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 ,
         \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 ,
         \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 ,
         \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 ,
         \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 ,
         \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 ,
         \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 ,
         \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 ,
         \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 ,
         \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 ,
         \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 ,
         \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 ,
         \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 ,
         \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 , \998 ,
         \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 ,
         \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 ,
         \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 ,
         \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 ,
         \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 ,
         \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 ,
         \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 ,
         \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 ,
         \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 ,
         \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 ,
         \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 ,
         \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 ,
         \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 ,
         \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 ,
         \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 ,
         \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 ,
         \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 ,
         \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 ,
         \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 ,
         \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 ,
         \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 ,
         \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 ,
         \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 ,
         \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 ,
         \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 ,
         \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 ,
         \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 ,
         \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 ,
         \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 ,
         \1289 , \1290 , \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 ,
         \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 ,
         \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 ,
         \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 ,
         \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 ,
         \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 ,
         \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 ,
         \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 ,
         \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 ,
         \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 ,
         \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 ,
         \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 ,
         \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 ,
         \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 ,
         \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 ,
         \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 ,
         \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 ,
         \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 ,
         \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 ,
         \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 ,
         \1489 , \1490 , \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 ,
         \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 ,
         \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 ,
         \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 ,
         \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 ,
         \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 ,
         \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 ,
         \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 ,
         \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 ,
         \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 ,
         \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 ,
         \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 ,
         \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 ,
         \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 ,
         \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 ,
         \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 ,
         \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 ,
         \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 ,
         \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 ,
         \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 ,
         \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 ,
         \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 ,
         \1709 , \1710 , \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 ,
         \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 ,
         \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 ,
         \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 ,
         \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 ,
         \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 ,
         \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 ,
         \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 ,
         \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 ,
         \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 ,
         \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 ,
         \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 ,
         \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 ,
         \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 ,
         \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 ,
         \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 ,
         \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 ,
         \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 ,
         \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 ,
         \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 ,
         \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 ,
         \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 ,
         \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 ,
         \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 ,
         \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 ,
         \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 ,
         \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 ,
         \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 ,
         \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 ,
         \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 ,
         \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 ,
         \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 ,
         \2029 , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 ,
         \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 ,
         \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 ,
         \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 ,
         \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 ,
         \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 ,
         \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 ,
         \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 ,
         \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 ,
         \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 ,
         \2129 , \2130 , \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 ,
         \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 ,
         \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 ,
         \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 ,
         \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 ,
         \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 ,
         \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 ,
         \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 ,
         \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 ,
         \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 ,
         \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 ,
         \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 ,
         \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 ,
         \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 ,
         \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 ,
         \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 ,
         \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 ,
         \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 ,
         \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 ,
         \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 ,
         \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 ,
         \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 ,
         \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 ,
         \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 ,
         \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 ,
         \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 ,
         \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 ,
         \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 ,
         \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 ,
         \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 ,
         \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 ,
         \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 ,
         \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 ,
         \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 ,
         \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 ,
         \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 ,
         \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 ,
         \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 ,
         \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 ,
         \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 ,
         \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 ,
         \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 ,
         \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 ,
         \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 ,
         \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 ,
         \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 ,
         \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 ,
         \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 ,
         \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 ,
         \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 ,
         \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 ,
         \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 ,
         \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 ,
         \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 ,
         \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 ,
         \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 ,
         \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 ,
         \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 ,
         \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 ,
         \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 ,
         \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 ,
         \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 ,
         \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 ,
         \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 ,
         \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 ,
         \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 ,
         \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 ,
         \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 ,
         \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 ,
         \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 ,
         \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 ,
         \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 ,
         \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 ,
         \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 ,
         \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 ,
         \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 ,
         \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 ,
         \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 ,
         \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 ,
         \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 ,
         \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 ,
         \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 ,
         \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 ,
         \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 ,
         \2969 , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 ,
         \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 ,
         \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 ,
         \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 ,
         \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 ,
         \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 ,
         \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 ,
         \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 ,
         \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 ,
         \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 ,
         \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 ,
         \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 ,
         \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 ,
         \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 ,
         \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 ,
         \3119 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 ,
         \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 ,
         \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 ,
         \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 ,
         \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 ,
         \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 ,
         \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 ,
         \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 ,
         \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 ,
         \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 ,
         \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 ,
         \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 ,
         \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 ,
         \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 ,
         \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 ,
         \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 ,
         \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 ,
         \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 ,
         \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 ,
         \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 ,
         \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 ,
         \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 ,
         \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 ,
         \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 ,
         \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 ,
         \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 ,
         \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 ,
         \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 ,
         \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 ,
         \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 ,
         \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 ,
         \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 ,
         \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 ,
         \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 ,
         \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 ,
         \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 ,
         \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 ,
         \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 ,
         \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 ,
         \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 ,
         \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 ,
         \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 ,
         \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 ,
         \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 ,
         \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 ,
         \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 ,
         \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 ,
         \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 ,
         \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 ,
         \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 ,
         \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 ,
         \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 ,
         \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 ,
         \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 ,
         \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 ,
         \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 ,
         \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 ,
         \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 ,
         \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 ,
         \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 ,
         \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 ,
         \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 ,
         \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 ,
         \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 ,
         \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 ,
         \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 ,
         \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 ,
         \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 ,
         \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 ,
         \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 ,
         \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 ,
         \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 ,
         \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 ,
         \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 ,
         \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 ,
         \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 ,
         \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 ,
         \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 ,
         \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 ,
         \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 ,
         \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 ,
         \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 ,
         \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 ,
         \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 ,
         \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 ,
         \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 ,
         \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 ,
         \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 ,
         \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 ,
         \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 ,
         \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 ,
         \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 ,
         \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 ,
         \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 ,
         \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 ,
         \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 ,
         \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 ,
         \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 ,
         \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 ,
         \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 ,
         \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 ,
         \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 ,
         \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 ,
         \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 ,
         \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 ,
         \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 ,
         \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 ,
         \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 ,
         \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 ,
         \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 ,
         \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 ,
         \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 ,
         \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 ,
         \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 ,
         \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 ,
         \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 ,
         \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 ,
         \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 ,
         \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 ,
         \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 ,
         \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 ,
         \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 ,
         \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 ,
         \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 ,
         \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 ,
         \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 ,
         \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 ,
         \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 ,
         \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 ,
         \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 ,
         \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 ,
         \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 ,
         \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 ,
         \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 ,
         \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 ,
         \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 ,
         \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 ,
         \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 ,
         \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 ,
         \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 ,
         \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 ,
         \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 ,
         \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 ,
         \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 ,
         \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 ,
         \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 ,
         \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 ,
         \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 ,
         \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 ,
         \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 ,
         \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 ,
         \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 ,
         \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 ,
         \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 ,
         \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 ,
         \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 ,
         \4679 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 ,
         \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 ,
         \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 ,
         \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 ,
         \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 ,
         \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 ,
         \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 ,
         \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 ,
         \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 ,
         \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 ,
         \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 ,
         \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 ,
         \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 ,
         \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 ,
         \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 ,
         \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 ,
         \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 ,
         \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 ,
         \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 ,
         \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 ,
         \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 ,
         \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 ,
         \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 ,
         \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 ,
         \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 ,
         \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 ,
         \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 ,
         \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 ,
         \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 ,
         \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 ,
         \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 ,
         \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 ,
         \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 ,
         \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 ,
         \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 ,
         \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 ,
         \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 ,
         \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 ,
         \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 ,
         \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 ,
         \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 ,
         \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 ,
         \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 ,
         \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 ,
         \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 ,
         \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 ,
         \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 ,
         \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 ,
         \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 ,
         \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 ,
         \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 ,
         \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 ,
         \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 ,
         \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 ,
         \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 ,
         \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 ,
         \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 ,
         \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 ,
         \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 ,
         \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 ,
         \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 ,
         \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 ,
         \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 ,
         \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 ,
         \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 ,
         \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 ,
         \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 ,
         \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 ,
         \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 ,
         \5369 , \5370 , \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 ,
         \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 ,
         \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 ,
         \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 ,
         \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 ,
         \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 ,
         \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 ,
         \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 ,
         \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 ,
         \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 ,
         \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 ,
         \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 ,
         \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 ,
         \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 ,
         \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 ,
         \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 ,
         \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 ,
         \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 ,
         \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 ,
         \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 ,
         \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 ,
         \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 ,
         \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 ,
         \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 ,
         \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 ,
         \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 ,
         \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 ,
         \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 ,
         \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 ,
         \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 ,
         \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 ,
         \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 ,
         \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 ,
         \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 ,
         \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 ,
         \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 ,
         \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 ,
         \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 ,
         \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 ,
         \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 ,
         \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 ,
         \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 ,
         \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 ,
         \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 ,
         \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818 ,
         \5819 , \5820 , \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 ,
         \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 ,
         \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 ,
         \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 ,
         \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 ,
         \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 ,
         \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 ,
         \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 ,
         \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 ,
         \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 ,
         \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 ,
         \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 ,
         \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 ,
         \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 ,
         \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 ,
         \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 ,
         \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 ,
         \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 ,
         \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 ,
         \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 ,
         \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 ,
         \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 ,
         \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 ,
         \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 ,
         \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 ,
         \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 ,
         \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 ,
         \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 ,
         \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 ,
         \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 ,
         \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 ,
         \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 ,
         \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 ,
         \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 ,
         \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 ,
         \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 ,
         \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 ,
         \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 ,
         \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 ,
         \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 ,
         \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 ,
         \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 ,
         \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 ,
         \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 ,
         \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 ,
         \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 ,
         \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 ,
         \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 ,
         \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 ,
         \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 ,
         \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 ,
         \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 ,
         \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 ,
         \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 ,
         \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 ,
         \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 ,
         \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 ,
         \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 ,
         \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 ,
         \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 ,
         \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 ,
         \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 ,
         \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 ,
         \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 ,
         \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 ,
         \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 ,
         \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 ,
         \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 ,
         \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 ,
         \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 ,
         \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 ,
         \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 ,
         \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 ,
         \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 ,
         \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 ,
         \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 ,
         \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 ,
         \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 ,
         \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 ,
         \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 ,
         \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 ,
         \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 ,
         \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 ,
         \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 ,
         \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 ,
         \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 ,
         \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 ,
         \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 ,
         \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 ,
         \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 ,
         \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 ,
         \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 ,
         \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 ,
         \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 ,
         \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 ,
         \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 ,
         \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 ,
         \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 ,
         \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 ,
         \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 ,
         \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 ,
         \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 ,
         \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 ,
         \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 ,
         \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 ,
         \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 ,
         \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 ,
         \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 ,
         \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 ,
         \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 ,
         \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 ,
         \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 ,
         \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 ,
         \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 ,
         \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 ,
         \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 ,
         \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 ,
         \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 ,
         \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 ,
         \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 ,
         \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 ,
         \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 ,
         \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 ,
         \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 ,
         \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 ,
         \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 ,
         \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 ,
         \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 ,
         \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 ,
         \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 ,
         \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 ,
         \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 ,
         \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 ,
         \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 ,
         \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 ,
         \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 ,
         \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 ,
         \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 ,
         \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 ,
         \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 ,
         \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 ,
         \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 ,
         \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 ,
         \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 ,
         \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 ,
         \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 ,
         \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 ,
         \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 ,
         \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 ,
         \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 ,
         \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 ,
         \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 ,
         \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 ,
         \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 ,
         \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 ,
         \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 ,
         \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 ,
         \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 ,
         \7399 , \7400 , \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 ,
         \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 ,
         \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 ,
         \7429 , \7430 , \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 ,
         \7439 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 ,
         \7449 , \7450 , \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 ,
         \7459 , \7460 , \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 ,
         \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 ,
         \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 ,
         \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 ,
         \7499 , \7500 , \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 ,
         \7509 , \7510 , \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 ,
         \7519 , \7520 , \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 ,
         \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 ,
         \7539 , \7540 , \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 ,
         \7549 , \7550 , \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 ,
         \7559 , \7560 , \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 ,
         \7569 , \7570 , \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 ,
         \7579 , \7580 , \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 ,
         \7589 , \7590 , \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 ,
         \7599 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 ,
         \7609 , \7610 , \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 ,
         \7619 , \7620 , \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 ,
         \7629 , \7630 , \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 ,
         \7639 , \7640 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 ,
         \7649 , \7650 , \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 ,
         \7659 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 ,
         \7669 , \7670 , \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 ,
         \7679 , \7680 , \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 ,
         \7689 , \7690 , \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 ,
         \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 ,
         \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 ,
         \7719 , \7720 , \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 ,
         \7729 , \7730 , \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 ,
         \7739 , \7740 , \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 ,
         \7749 , \7750 , \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 ,
         \7759 , \7760 , \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 , \7768 ,
         \7769 , \7770 , \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 ,
         \7779 , \7780 , \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 ,
         \7789 , \7790 , \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 ,
         \7799 , \7800 , \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 ,
         \7809 , \7810 , \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 ,
         \7819 , \7820 , \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 ,
         \7829 , \7830 , \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 ,
         \7839 , \7840 , \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 ,
         \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 ,
         \7859 , \7860 , \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 , \7868 ,
         \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 ,
         \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 ,
         \7889 , \7890 , \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 ,
         \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 ,
         \7909 , \7910 , \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 , \7918 ,
         \7919 , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 ,
         \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 ,
         \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 ,
         \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 ,
         \7959 , \7960 , \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 ,
         \7969 , \7970 , \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 ,
         \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 ,
         \7989 , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 ,
         \7999 , \8000 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 ,
         \8009 , \8010 , \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 ,
         \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 ,
         \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 ,
         \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 ,
         \8049 , \8050 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 , \8058 ,
         \8059 , \8060 , \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 ,
         \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 ,
         \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 ,
         \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 ,
         \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 ,
         \8109 , \8110 , \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 ,
         \8119 , \8120 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 ,
         \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 ,
         \8139 , \8140 , \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 ,
         \8149 , \8150 , \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 , \8158 ,
         \8159 , \8160 , \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 ,
         \8169 , \8170 , \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 , \8178 ,
         \8179 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 ,
         \8189 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 ,
         \8199 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208 ,
         \8209 , \8210 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 ,
         \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 , \8228 ,
         \8229 , \8230 , \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 ,
         \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 ,
         \8249 , \8250 , \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 ,
         \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 ,
         \8269 , \8270 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 ,
         \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 ,
         \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 , \8298 ,
         \8299 , \8300 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 ,
         \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318 ,
         \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 ,
         \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 , \8338 ,
         \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 ,
         \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 ,
         \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 ,
         \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 ,
         \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 ,
         \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 ,
         \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 ,
         \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 ,
         \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 ,
         \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 ,
         \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 ,
         \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 ,
         \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 ,
         \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 ,
         \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 , \8488 ,
         \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 ,
         \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 , \8508 ,
         \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 ,
         \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 , \8528 ,
         \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 ,
         \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 , \8548 ,
         \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 ,
         \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 ,
         \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 ,
         \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 ,
         \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 ,
         \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 ,
         \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 ,
         \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 ,
         \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 ,
         \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 ,
         \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 ,
         \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 ,
         \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 ,
         \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 ,
         \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 ,
         \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 ,
         \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 ,
         \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 ,
         \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 ,
         \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 ,
         \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 , \8758 ,
         \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 ,
         \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 ,
         \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 ,
         \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 ,
         \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 ,
         \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 ,
         \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 ,
         \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 ,
         \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 ,
         \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 ,
         \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 , \8868 ,
         \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 ,
         \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 ,
         \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 , \8898 ,
         \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 ,
         \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918 ,
         \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 , \8928 ,
         \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 ,
         \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 ,
         \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 , \8958 ,
         \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 ,
         \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 ,
         \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 ,
         \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 ,
         \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 , \9008 ,
         \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 ,
         \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 ,
         \9029 , \9030 , \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 , \9038 ,
         \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048 ,
         \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 ,
         \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 ,
         \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 , \9078 ,
         \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 ,
         \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 , \9098 ,
         \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 , \9108 ,
         \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 , \9118 ,
         \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 , \9128 ,
         \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 , \9138 ,
         \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 , \9148 ,
         \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 , \9158 ,
         \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 , \9168 ,
         \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 , \9178 ,
         \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 , \9188 ,
         \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 , \9198 ,
         \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 , \9208 ,
         \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 , \9218 ,
         \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 , \9228 ,
         \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 , \9238 ,
         \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 , \9248 ,
         \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 , \9258 ,
         \9259 , \9260 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 , \9268 ,
         \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 , \9278 ,
         \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 , \9288 ,
         \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 , \9298 ,
         \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 , \9308 ,
         \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 , \9318 ,
         \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 , \9328 ,
         \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 , \9338 ,
         \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 , \9348 ,
         \9349 , \9350 , \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 , \9358 ,
         \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 , \9368 ,
         \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 , \9378 ,
         \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 , \9388 ,
         \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 , \9398 ,
         \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 , \9408 ,
         \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 , \9418 ,
         \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 , \9428 ,
         \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 , \9438 ,
         \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 , \9448 ,
         \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 , \9458 ,
         \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 , \9468 ,
         \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 , \9478 ,
         \9479 , \9480 , \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 , \9488 ,
         \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 , \9498 ,
         \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 , \9508 ,
         \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 , \9518 ,
         \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 , \9528 ,
         \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 , \9538 ,
         \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 , \9548 ,
         \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 , \9558 ,
         \9559 , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 , \9568 ,
         \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 , \9578 ,
         \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 , \9588 ,
         \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 , \9598 ,
         \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 , \9608 ,
         \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 , \9618 ,
         \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 , \9628 ,
         \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 , \9638 ,
         \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 , \9648 ,
         \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 ,
         \9659 , \9660 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 , \9668 ,
         \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 ,
         \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 ,
         \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 , \9698 ,
         \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 ,
         \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 , \9718 ,
         \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 ,
         \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 , \9738 ,
         \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 ,
         \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 ,
         \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 , \9768 ,
         \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 ,
         \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 ,
         \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 ,
         \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 ,
         \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 ,
         \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 ,
         \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 ,
         \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 ,
         \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 ,
         \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 ,
         \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 ,
         \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 ,
         \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 ,
         \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 ,
         \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 ,
         \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 ,
         \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 ,
         \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 ,
         \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 ,
         \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 ,
         \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 ,
         \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 ,
         \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 ,
         \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 ,
         \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 ,
         \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 ,
         \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 ,
         \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 ,
         \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 , \10058 ,
         \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 ,
         \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 ,
         \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 ,
         \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 ,
         \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 ,
         \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 ,
         \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 ,
         \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 ,
         \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 ,
         \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 ,
         \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 ,
         \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 ,
         \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 ,
         \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 ,
         \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 ,
         \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 ,
         \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 ,
         \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 ,
         \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 ,
         \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 ,
         \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 , \10268 ,
         \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 ,
         \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 ,
         \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 ,
         \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 ,
         \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 ,
         \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 ,
         \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 ,
         \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 , \10348 ,
         \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 ,
         \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 , \10368 ,
         \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 ,
         \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 ,
         \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 , \10398 ,
         \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 ,
         \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 ,
         \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 ,
         \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 ,
         \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 ,
         \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 ,
         \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 ,
         \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 ,
         \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 ,
         \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 ,
         \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 ,
         \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 ,
         \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 ,
         \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 ,
         \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 ,
         \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 ,
         \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 ,
         \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 ,
         \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 ,
         \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 ,
         \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 ,
         \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 , \10618 ,
         \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 ,
         \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 ,
         \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 ,
         \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 , \10658 ,
         \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 ,
         \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 ,
         \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 ,
         \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 ,
         \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 ,
         \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 ,
         \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 ,
         \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 ,
         \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 ,
         \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 ,
         \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 ,
         \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 ,
         \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 ,
         \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 ,
         \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 ,
         \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 ,
         \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 ,
         \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 ,
         \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 ,
         \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 ,
         \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 ,
         \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 ,
         \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 ,
         \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 ,
         \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 ,
         \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 ,
         \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 ,
         \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 ,
         \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 ,
         \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 , \10958 ,
         \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 ,
         \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 ,
         \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 , \10988 ,
         \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 ,
         \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 ,
         \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 ,
         \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 ,
         \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 ,
         \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 ,
         \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 ,
         \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 ,
         \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 ,
         \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 ,
         \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 ,
         \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 ,
         \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 ,
         \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 ,
         \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 ,
         \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 ,
         \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 ,
         \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 ,
         \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 ,
         \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 ,
         \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 ,
         \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 ,
         \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 ,
         \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 ,
         \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 ,
         \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 ,
         \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 ,
         \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11268 ,
         \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 , \11278 ,
         \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 ,
         \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 ,
         \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 , \11308 ,
         \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 ,
         \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 ,
         \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 ,
         \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 ,
         \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 ,
         \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 ,
         \11369 , \11370 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 ,
         \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 ,
         \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 ,
         \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 ,
         \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 ,
         \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 ,
         \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 , \11438 ,
         \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 ,
         \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 ,
         \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 ,
         \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 ,
         \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 ,
         \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 ,
         \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 ,
         \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 ,
         \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 ,
         \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 ,
         \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 ,
         \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 ,
         \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 , \11568 ,
         \11569 , \11570 , \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 , \11578 ,
         \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 , \11588 ,
         \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 , \11598 ,
         \11599 , \11600 , \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 , \11608 ,
         \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 ,
         \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 ,
         \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 ,
         \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 ,
         \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 ,
         \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 ,
         \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 ,
         \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 ,
         \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 ,
         \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 ,
         \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 ,
         \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 ,
         \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 , \11738 ,
         \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 ,
         \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 ,
         \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 ,
         \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 ,
         \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 ,
         \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 ,
         \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 ,
         \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 ,
         \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 ,
         \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 ,
         \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 ,
         \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 ,
         \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 , \11868 ,
         \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 ,
         \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 ,
         \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 ,
         \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 ,
         \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 ,
         \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 ,
         \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 ,
         \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 ,
         \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 ,
         \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 ,
         \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 ,
         \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 ,
         \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 ,
         \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 , \12008 ,
         \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 ,
         \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 ,
         \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 ,
         \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 ,
         \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 ,
         \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 ,
         \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 ,
         \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 ,
         \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 ,
         \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 ,
         \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 ,
         \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 ,
         \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 ,
         \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 , \12148 ,
         \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 ,
         \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 ,
         \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 , \12178 ,
         \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 ,
         \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 ,
         \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 ,
         \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 ,
         \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 ,
         \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 ,
         \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 , \12248 ,
         \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 ,
         \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 ,
         \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 ,
         \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 ,
         \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 ,
         \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 ,
         \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 ,
         \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 ,
         \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 ,
         \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 ,
         \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 ,
         \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 ,
         \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 ,
         \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 ,
         \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 ,
         \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 ,
         \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 ,
         \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 ,
         \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 ,
         \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 ,
         \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 ,
         \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 ,
         \12469 , \12470 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 , \12478 ,
         \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 ,
         \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 ,
         \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 ,
         \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 ,
         \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 ,
         \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 ,
         \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 ,
         \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 ,
         \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 ,
         \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 ,
         \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 ,
         \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 ,
         \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 ,
         \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 ,
         \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 , \12628 ,
         \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 ,
         \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 ,
         \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 ,
         \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 ,
         \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 ,
         \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 ,
         \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 ,
         \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 ,
         \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 ,
         \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 , \12728 ,
         \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 ,
         \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 ,
         \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 ,
         \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 ,
         \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 , \12778 ,
         \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 ,
         \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 ,
         \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 ,
         \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 ,
         \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 ,
         \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 ,
         \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 ,
         \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 ,
         \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 ,
         \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 ,
         \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 ,
         \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 ,
         \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 ,
         \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 ,
         \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 ,
         \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 ,
         \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 ,
         \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 ,
         \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 ,
         \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978 ,
         \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 ,
         \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 ,
         \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 ,
         \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 , \13018 ,
         \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 ,
         \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 ,
         \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 ,
         \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 ,
         \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 ,
         \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 ,
         \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 ,
         \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 ,
         \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 ,
         \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 ,
         \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 ,
         \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 ,
         \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 ,
         \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 ,
         \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 ,
         \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 ,
         \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 , \13188 ,
         \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 ,
         \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 ,
         \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 , \13218 ,
         \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 ,
         \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 ,
         \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 ,
         \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 ,
         \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 ,
         \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 ,
         \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 ,
         \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 ,
         \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 ,
         \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 , \13318 ,
         \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 ,
         \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 ,
         \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 ,
         \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 , \13358 ,
         \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 ,
         \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 , \13378 ,
         \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 ,
         \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 ,
         \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 , \13408 ,
         \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 ,
         \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 ,
         \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 ,
         \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 ,
         \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 ,
         \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 ,
         \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 , \13478 ,
         \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 ,
         \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 , \13498 ,
         \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 ,
         \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 ,
         \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 , \13528 ,
         \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 ,
         \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 , \13548 ,
         \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 ,
         \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 ,
         \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 ,
         \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 ,
         \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 ,
         \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 ,
         \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 ,
         \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 ,
         \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 ,
         \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 ,
         \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 ,
         \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 ,
         \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 ,
         \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 ,
         \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 ,
         \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 ,
         \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 ,
         \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 ,
         \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 , \13738 ,
         \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 ,
         \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 , \13758 ,
         \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 ,
         \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 ,
         \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 ,
         \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 ,
         \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 ,
         \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 ,
         \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 ,
         \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 ,
         \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 ,
         \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 ,
         \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 ,
         \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 ,
         \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 ,
         \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 ,
         \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 ,
         \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 ,
         \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 ,
         \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 ,
         \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 ,
         \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 , \13958 ,
         \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 ,
         \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 ,
         \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 ,
         \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 ,
         \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 ,
         \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 ,
         \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 , \14028 ,
         \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 ,
         \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 ,
         \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 ,
         \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 ,
         \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 , \14078 ,
         \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 ,
         \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 ,
         \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 ,
         \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 ,
         \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 ,
         \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 ,
         \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 ,
         \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 ,
         \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 ,
         \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 ,
         \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 ,
         \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 ,
         \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 ,
         \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 ,
         \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 ,
         \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 ,
         \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 ,
         \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 ,
         \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 ,
         \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 ,
         \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 ,
         \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 ,
         \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 ,
         \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 ,
         \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 ,
         \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 ,
         \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 , \14348 ,
         \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 ,
         \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 ,
         \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 ,
         \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 ,
         \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 ,
         \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 ,
         \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 ,
         \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 ,
         \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 ,
         \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 ,
         \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 ,
         \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 ,
         \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 ,
         \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 ,
         \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 ,
         \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 ,
         \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 ,
         \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 ,
         \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 ,
         \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 ,
         \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 ,
         \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 ,
         \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 ,
         \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 ,
         \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 ,
         \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 ,
         \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 , \14618 ,
         \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 ,
         \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 ,
         \14639 , \14640 , \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 , \14648 ,
         \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 ,
         \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 ,
         \14669 , \14670 , \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 ,
         \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 ,
         \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 ,
         \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 ,
         \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 ,
         \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 ,
         \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 ,
         \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 ,
         \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 ,
         \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 ,
         \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 ,
         \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 ,
         \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 ,
         \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 ,
         \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 ,
         \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 ,
         \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 ,
         \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 ,
         \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 ,
         \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 ,
         \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 ,
         \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 ,
         \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 ,
         \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 ,
         \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 ,
         \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 ,
         \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 ,
         \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 ,
         \14949 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 , \14958 ,
         \14959 , \14960 , \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 ,
         \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 ,
         \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 , \14988 ,
         \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 ,
         \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 ,
         \15009 , \15010 , \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 , \15018 ,
         \15019 , \15020 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 ,
         \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 ,
         \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 , \15048 ,
         \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 ,
         \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 ,
         \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 ,
         \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 ,
         \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 ,
         \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 ,
         \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 ,
         \15119 , \15120 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 ,
         \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 ,
         \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 ,
         \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 ,
         \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 ,
         \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 ,
         \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 ,
         \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 ,
         \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 ,
         \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 ,
         \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 ,
         \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 ,
         \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 ,
         \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 ,
         \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 ,
         \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 ,
         \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 , \15288 ,
         \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 ,
         \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 ,
         \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 , \15318 ,
         \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 ,
         \15329 , \15330 , \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 , \15338 ,
         \15339 , \15340 , \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 ,
         \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 ,
         \15359 , \15360 , \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 , \15368 ,
         \15369 , \15370 , \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 ,
         \15379 , \15380 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 ,
         \15389 , \15390 , \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 ,
         \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 ,
         \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 ,
         \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 ,
         \15429 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 ,
         \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 ,
         \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 ,
         \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 ,
         \15469 , \15470 , \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 ,
         \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 ,
         \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 ,
         \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 ,
         \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 ,
         \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 ,
         \15529 , \15530 , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 ,
         \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 ,
         \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 , \15558 ,
         \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 ,
         \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 ,
         \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 ,
         \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 ,
         \15599 , \15600 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 , \15608 ,
         \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 ,
         \15619 , \15620 , \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 ,
         \15629 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 ,
         \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 ,
         \15649 , \15650 , \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 , \15658 ,
         \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 ,
         \15669 , \15670 , \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 ,
         \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 ,
         \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 ,
         \15699 , \15700 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 , \15708 ,
         \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 ,
         \15719 , \15720 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 ,
         \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 ,
         \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 ,
         \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 ,
         \15759 , \15760 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 ,
         \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 ,
         \15779 , \15780 , \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 , \15788 ,
         \15789 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 ,
         \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 ,
         \15809 , \15810 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 ,
         \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 ,
         \15829 , \15830 , \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 ,
         \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 ,
         \15849 , \15850 , \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 ,
         \15859 , \15860 , \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 ,
         \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 ,
         \15879 , \15880 , \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 ,
         \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 ,
         \15899 , \15900 , \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 ,
         \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 ,
         \15919 , \15920 , \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 ,
         \15929 , \15930 , \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 , \15938 ,
         \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 ,
         \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 ,
         \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 ,
         \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 ,
         \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 , \15988 ,
         \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 ,
         \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 ,
         \16009 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 ,
         \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 ,
         \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 ,
         \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 ,
         \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 ,
         \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 ,
         \16069 , \16070 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 ,
         \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 ,
         \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 ,
         \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 ,
         \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 ,
         \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 ,
         \16129 , \16130 , \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 ,
         \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 ,
         \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 ,
         \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 ,
         \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 ,
         \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 ,
         \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 , \16198 ,
         \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 ,
         \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 ,
         \16219 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 ,
         \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 ,
         \16239 , \16240 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 ,
         \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 ,
         \16259 , \16260 , \16261 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 ,
         \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 ,
         \16279 , \16280 , \16281 , \16282 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 ,
         \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 ,
         \16299 , \16300 , \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 ,
         \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 ,
         \16319 , \16320 , \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 ,
         \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 ,
         \16339 , \16340 , \16341 , \16342 , \16343 , \16344 , \16345 , \16346 , \16347 , \16348 ,
         \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 ,
         \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 ,
         \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 ,
         \16379 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 ,
         \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 ,
         \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 , \16408 ,
         \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 ,
         \16419 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 ,
         \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 ,
         \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448 ,
         \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 ,
         \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 ,
         \16469 , \16470 , \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 ,
         \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 ,
         \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 ,
         \16499 , \16500 , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 ,
         \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 ,
         \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 ,
         \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 ,
         \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 ,
         \16549 , \16550 , \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 , \16558 ,
         \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 ,
         \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 ,
         \16579 , \16580 , \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 ,
         \16589 , \16590 , \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 ,
         \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 ,
         \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 ,
         \16619 , \16620 , \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 ,
         \16629 , \16630 , \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 , \16638 ,
         \16639 , \16640 , \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 ,
         \16649 , \16650 , \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 ,
         \16659 , \16660 , \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 ,
         \16669 , \16670 , \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 , \16678 ,
         \16679 , \16680 , \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 , \16688 ,
         \16689 , \16690 , \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 ,
         \16699 , \16700 , \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 ,
         \16709 , \16710 , \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 , \16718 ,
         \16719 , \16720 , \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 , \16728 ,
         \16729 , \16730 , \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 ,
         \16739 , \16740 , \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 , \16748 ,
         \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 ,
         \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 ,
         \16769 , \16770 , \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 ,
         \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 ,
         \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 ,
         \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 ,
         \16809 , \16810 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 ,
         \16819 , \16820 , \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 , \16828 ,
         \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 ,
         \16839 , \16840 , \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 ,
         \16849 , \16850 , \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 , \16858 ,
         \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 ,
         \16869 , \16870 , \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 ,
         \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 ,
         \16889 , \16890 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 ,
         \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 ,
         \16909 , \16910 , \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 , \16918 ,
         \16919 , \16920 , \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 , \16928 ,
         \16929 , \16930 , \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 ,
         \16939 , \16940 , \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 , \16948 ,
         \16949 , \16950 , \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 ,
         \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 ,
         \16969 , \16970 , \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 ,
         \16979 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 ,
         \16989 , \16990 , \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 , \16998 ,
         \16999 , \17000 , \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 ,
         \17009 , \17010 , \17011 , \17012 , \17013 , \17014 , \17015 , \17016 , \17017 , \17018 ,
         \17019 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 ,
         \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 , \17038 ,
         \17039 , \17040 , \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 ,
         \17049 , \17050 , \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 ,
         \17059 , \17060 , \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 ,
         \17069 , \17070 , \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 , \17078 ,
         \17079 , \17080 , \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 , \17088 ,
         \17089 , \17090 , \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 ,
         \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 ,
         \17109 , \17110 , \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 ,
         \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 ,
         \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 , \17138 ,
         \17139 , \17140 , \17141 , \17142 , \17143 , \17144 , \17145 , \17146 , \17147 , \17148 ,
         \17149 , \17150 , \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 , \17158 ,
         \17159 , \17160 , \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 , \17168 ,
         \17169 , \17170 , \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 , \17178 ,
         \17179 , \17180 , \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188 ,
         \17189 , \17190 , \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 , \17198 ,
         \17199 , \17200 , \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 ,
         \17209 , \17210 , \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 ,
         \17219 , \17220 , \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 , \17228 ,
         \17229 , \17230 , \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 , \17238 ,
         \17239 , \17240 , \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 , \17248 ,
         \17249 , \17250 , \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 , \17258 ,
         \17259 , \17260 , \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 , \17268 ,
         \17269 , \17270 , \17271 , \17272 , \17273 , \17274 , \17275 , \17276 , \17277 , \17278 ,
         \17279 , \17280 , \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 , \17288 ,
         \17289 , \17290 , \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 , \17298 ,
         \17299 , \17300 , \17301 , \17302 , \17303 , \17304 , \17305 , \17306 , \17307 , \17308 ,
         \17309 , \17310 , \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 , \17318 ,
         \17319 , \17320 , \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 , \17328 ,
         \17329 , \17330 , \17331 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 , \17338 ,
         \17339 , \17340 , \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 , \17348 ,
         \17349 , \17350 , \17351 , \17352 , \17353 , \17354 , \17355 , \17356 , \17357 , \17358 ,
         \17359 , \17360 , \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 , \17368 ,
         \17369 , \17370 , \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 , \17378 ,
         \17379 , \17380 , \17381 , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 , \17388 ,
         \17389 , \17390 , \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 , \17398 ,
         \17399 , \17400 , \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 , \17408 ,
         \17409 , \17410 , \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 , \17418 ,
         \17419 , \17420 , \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 , \17428 ,
         \17429 , \17430 , \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 , \17438 ,
         \17439 , \17440 , \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 , \17448 ,
         \17449 , \17450 , \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 , \17458 ,
         \17459 , \17460 , \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 , \17468 ,
         \17469 , \17470 , \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 , \17478 ,
         \17479 , \17480 , \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 , \17488 ,
         \17489 , \17490 , \17491 , \17492 , \17493 , \17494 , \17495 , \17496 , \17497 , \17498 ,
         \17499 , \17500 , \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 , \17508 ,
         \17509 , \17510 , \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 , \17518 ,
         \17519 , \17520 , \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 , \17528 ,
         \17529 , \17530 , \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 , \17538 ,
         \17539 , \17540 , \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 , \17548 ,
         \17549 , \17550 , \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 , \17558 ,
         \17559 , \17560 , \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 , \17568 ,
         \17569 , \17570 , \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 , \17578 ,
         \17579 , \17580 , \17581 , \17582 , \17583 , \17584 , \17585 , \17586 , \17587 , \17588 ,
         \17589 , \17590 , \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 , \17598 ,
         \17599 , \17600 , \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 , \17608 ,
         \17609 , \17610 , \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 , \17618 ,
         \17619 , \17620 , \17621 , \17622 , \17623 , \17624 , \17625 , \17626 , \17627 , \17628 ,
         \17629 , \17630 , \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 , \17638 ,
         \17639 , \17640 , \17641 , \17642 , \17643 , \17644 , \17645 , \17646 , \17647 , \17648 ,
         \17649 , \17650 , \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 , \17658 ,
         \17659 , \17660 , \17661 , \17662 , \17663 , \17664 , \17665 , \17666 , \17667 , \17668 ,
         \17669 , \17670 , \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 , \17678 ,
         \17679 , \17680 , \17681 , \17682 , \17683 , \17684 , \17685 , \17686 , \17687 , \17688 ,
         \17689 , \17690 , \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 , \17698 ,
         \17699 , \17700 , \17701 , \17702 , \17703 , \17704 , \17705 , \17706 , \17707 , \17708 ,
         \17709 , \17710 , \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 , \17718 ,
         \17719 , \17720 , \17721 , \17722 , \17723 , \17724 , \17725 , \17726 , \17727 , \17728 ,
         \17729 , \17730 , \17731 , \17732 , \17733 , \17734 , \17735 , \17736 , \17737 , \17738 ,
         \17739 , \17740 , \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 , \17748 ,
         \17749 , \17750 , \17751 , \17752 , \17753 , \17754 , \17755 , \17756 , \17757 , \17758 ,
         \17759 , \17760 , \17761 , \17762 , \17763 , \17764 , \17765 , \17766 , \17767 , \17768 ,
         \17769 , \17770 , \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 , \17778 ,
         \17779 , \17780 , \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 , \17788 ,
         \17789 , \17790 , \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 , \17798 ,
         \17799 , \17800 , \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 , \17808 ,
         \17809 , \17810 , \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 , \17818 ,
         \17819 , \17820 , \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 , \17828 ,
         \17829 , \17830 , \17831 , \17832 , \17833 , \17834 , \17835 , \17836 , \17837 , \17838 ,
         \17839 , \17840 , \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 , \17848 ,
         \17849 , \17850 , \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 , \17858 ,
         \17859 , \17860 , \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 , \17868 ,
         \17869 , \17870 , \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 , \17878 ,
         \17879 , \17880 , \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 , \17888 ,
         \17889 , \17890 , \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 , \17898 ,
         \17899 , \17900 , \17901 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 , \17908 ,
         \17909 , \17910 , \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 , \17918 ,
         \17919 , \17920 , \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 , \17928 ,
         \17929 , \17930 , \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 , \17938 ,
         \17939 , \17940 , \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 , \17948 ,
         \17949 , \17950 , \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 , \17958 ,
         \17959 , \17960 , \17961 , \17962 , \17963 , \17964 , \17965 , \17966 , \17967 , \17968 ,
         \17969 , \17970 , \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 , \17978 ,
         \17979 , \17980 , \17981 , \17982 , \17983 , \17984 , \17985 , \17986 , \17987 , \17988 ,
         \17989 , \17990 , \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 , \17998 ,
         \17999 , \18000 , \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 , \18008 ,
         \18009 , \18010 , \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 , \18018 ,
         \18019 , \18020 , \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 , \18028 ,
         \18029 , \18030 , \18031 , \18032 , \18033 , \18034 , \18035 , \18036 , \18037 , \18038 ,
         \18039 , \18040 , \18041 , \18042 , \18043 , \18044 , \18045 , \18046 , \18047 , \18048 ,
         \18049 , \18050 , \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 , \18058 ,
         \18059 , \18060 , \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 , \18068 ,
         \18069 , \18070 , \18071 , \18072 , \18073 , \18074 , \18075 , \18076 , \18077 , \18078 ,
         \18079 , \18080 , \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 , \18088 ,
         \18089 , \18090 , \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 , \18098 ,
         \18099 , \18100 , \18101 , \18102 , \18103 , \18104 , \18105 , \18106 , \18107 , \18108 ,
         \18109 , \18110 , \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 , \18118 ,
         \18119 , \18120 , \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 , \18128 ,
         \18129 , \18130 , \18131 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 , \18138 ,
         \18139 , \18140 , \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 , \18148 ,
         \18149 , \18150 , \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 , \18158 ,
         \18159 , \18160 , \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 , \18168 ,
         \18169 , \18170 , \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 , \18178 ,
         \18179 , \18180 , \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 , \18188 ,
         \18189 , \18190 , \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 , \18198 ,
         \18199 , \18200 , \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 , \18208 ,
         \18209 , \18210 , \18211 , \18212 , \18213 , \18214 , \18215 , \18216 , \18217 , \18218 ,
         \18219 , \18220 , \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 , \18228 ,
         \18229 , \18230 , \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 , \18238 ,
         \18239 , \18240 , \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 , \18248 ,
         \18249 , \18250 , \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 , \18258 ,
         \18259 , \18260 , \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 , \18268 ,
         \18269 , \18270 , \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 , \18278 ,
         \18279 , \18280 , \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 , \18288 ,
         \18289 , \18290 , \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 , \18298 ,
         \18299 , \18300 , \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 , \18308 ,
         \18309 , \18310 , \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 , \18318 ,
         \18319 , \18320 , \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 , \18328 ,
         \18329 , \18330 , \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 , \18338 ,
         \18339 , \18340 , \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 , \18348 ,
         \18349 , \18350 , \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 , \18358 ,
         \18359 , \18360 , \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 , \18368 ,
         \18369 , \18370 , \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 , \18378 ,
         \18379 , \18380 , \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 , \18388 ,
         \18389 , \18390 , \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 , \18398 ,
         \18399 , \18400 , \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 , \18408 ,
         \18409 , \18410 , \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 , \18418 ,
         \18419 , \18420 , \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 , \18428 ,
         \18429 , \18430 , \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 , \18438 ,
         \18439 , \18440 , \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 , \18448 ,
         \18449 , \18450 , \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 , \18458 ,
         \18459 , \18460 , \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 , \18468 ,
         \18469 , \18470 , \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 , \18478 ,
         \18479 , \18480 , \18481 , \18482 , \18483 , \18484 , \18485 , \18486 , \18487 , \18488 ,
         \18489 , \18490 , \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 , \18498 ,
         \18499 , \18500 , \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 , \18508 ,
         \18509 , \18510 , \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 , \18518 ,
         \18519 , \18520 , \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 , \18528 ,
         \18529 , \18530 , \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 , \18538 ,
         \18539 , \18540 , \18541 , \18542 , \18543 , \18544 , \18545 , \18546 , \18547 , \18548 ,
         \18549 , \18550 , \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 , \18558 ,
         \18559 , \18560 , \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 , \18568 ,
         \18569 , \18570 , \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 , \18578 ,
         \18579 , \18580 , \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 , \18588 ,
         \18589 , \18590 , \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 , \18598 ,
         \18599 , \18600 , \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 , \18608 ,
         \18609 , \18610 , \18611 , \18612 , \18613 , \18614 , \18615 , \18616 , \18617 , \18618 ,
         \18619 , \18620 , \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 , \18628 ,
         \18629 , \18630 , \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 , \18638 ,
         \18639 , \18640 , \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 , \18648 ,
         \18649 , \18650 , \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 , \18658 ,
         \18659 , \18660 , \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 , \18668 ,
         \18669 , \18670 , \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 , \18678 ,
         \18679 , \18680 , \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 , \18688 ,
         \18689 , \18690 , \18691 , \18692 , \18693 , \18694 , \18695 , \18696 , \18697 , \18698 ,
         \18699 , \18700 , \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 , \18708 ,
         \18709 , \18710 , \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717 , \18718 ,
         \18719 , \18720 , \18721 , \18722 , \18723 , \18724 , \18725 , \18726 , \18727 , \18728 ,
         \18729 , \18730 , \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 , \18738 ,
         \18739 , \18740 , \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 , \18748 ,
         \18749 , \18750 , \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 , \18758 ,
         \18759 , \18760 , \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 , \18768 ,
         \18769 , \18770 , \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 , \18778 ,
         \18779 , \18780 , \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 , \18788 ,
         \18789 , \18790 , \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 , \18798 ,
         \18799 , \18800 , \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 , \18808 ,
         \18809 , \18810 , \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 , \18818 ,
         \18819 , \18820 , \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 , \18828 ,
         \18829 , \18830 , \18831 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 , \18838 ,
         \18839 , \18840 , \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 , \18848 ,
         \18849 , \18850 , \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 , \18858 ,
         \18859 , \18860 , \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 , \18868 ,
         \18869 , \18870 , \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 , \18878 ,
         \18879 , \18880 , \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887 , \18888 ,
         \18889 , \18890 , \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 , \18898 ,
         \18899 , \18900 , \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 , \18908 ,
         \18909 , \18910 , \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 , \18918 ,
         \18919 , \18920 , \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 , \18928 ,
         \18929 , \18930 , \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 , \18938 ,
         \18939 , \18940 , \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 , \18948 ,
         \18949 , \18950 , \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 , \18958 ,
         \18959 , \18960 , \18961 , \18962 , \18963 , \18964 , \18965 , \18966 , \18967 , \18968 ,
         \18969 , \18970 , \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 , \18978 ,
         \18979 , \18980 , \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 , \18988 ,
         \18989 , \18990 , \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 , \18998 ,
         \18999 , \19000 , \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 , \19008 ,
         \19009 , \19010 , \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 , \19018 ,
         \19019 , \19020 , \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 , \19028 ,
         \19029 , \19030 , \19031 , \19032 , \19033 , \19034 , \19035 , \19036 , \19037 , \19038 ,
         \19039 , \19040 , \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 , \19048 ,
         \19049 , \19050 , \19051 , \19052 , \19053 , \19054 , \19055 , \19056 , \19057 , \19058 ,
         \19059 , \19060 , \19061 , \19062 , \19063 , \19064 , \19065 , \19066 , \19067 , \19068 ,
         \19069 , \19070 , \19071 , \19072 , \19073 , \19074 , \19075 , \19076 , \19077 , \19078 ,
         \19079 , \19080 , \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 , \19088 ,
         \19089 , \19090 , \19091 , \19092 , \19093 , \19094 , \19095 , \19096 , \19097 , \19098 ,
         \19099 , \19100 , \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 , \19108 ,
         \19109 , \19110 , \19111 , \19112 , \19113 , \19114 , \19115 , \19116 , \19117 , \19118 ,
         \19119 , \19120 , \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 , \19128 ,
         \19129 , \19130 , \19131 , \19132 , \19133 , \19134 , \19135 , \19136 , \19137 , \19138 ,
         \19139 , \19140 , \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 , \19148 ,
         \19149 , \19150 , \19151 , \19152 , \19153 , \19154 , \19155 , \19156 , \19157 , \19158 ,
         \19159 , \19160 , \19161 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 , \19168 ,
         \19169 , \19170 , \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 , \19178 ,
         \19179 , \19180 , \19181 , \19182 , \19183 , \19184 , \19185 , \19186 , \19187 , \19188 ,
         \19189 , \19190 , \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 , \19198 ,
         \19199 , \19200 , \19201 , \19202 , \19203 , \19204 , \19205 , \19206 , \19207 , \19208 ,
         \19209 , \19210 , \19211 , \19212 , \19213 , \19214 , \19215 , \19216 , \19217 , \19218 ,
         \19219 , \19220 , \19221 , \19222 , \19223 , \19224 , \19225 , \19226 , \19227 , \19228 ,
         \19229 , \19230 , \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 , \19238 ,
         \19239 , \19240 , \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 , \19248 ,
         \19249 , \19250 , \19251 , \19252 , \19253 , \19254 , \19255 , \19256 , \19257 , \19258 ,
         \19259 , \19260 , \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 , \19268 ,
         \19269 , \19270 , \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 , \19278 ,
         \19279 , \19280 , \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 , \19288 ,
         \19289 , \19290 , \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 , \19298 ,
         \19299 , \19300 , \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 , \19308 ,
         \19309 , \19310 , \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 , \19318 ,
         \19319 , \19320 , \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 , \19328 ,
         \19329 , \19330 , \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 , \19338 ,
         \19339 , \19340 , \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 , \19348 ,
         \19349 , \19350 , \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 , \19358 ,
         \19359 , \19360 , \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 , \19368 ,
         \19369 , \19370 , \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 , \19378 ,
         \19379 , \19380 , \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 , \19388 ,
         \19389 , \19390 , \19391 , \19392 , \19393 , \19394 , \19395 , \19396 , \19397 , \19398 ,
         \19399 , \19400 , \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 , \19408 ,
         \19409 , \19410 , \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 , \19418 ,
         \19419 , \19420 , \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 , \19428 ,
         \19429 , \19430 , \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 , \19438 ,
         \19439 , \19440 , \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 , \19448 ,
         \19449 , \19450 , \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 , \19458 ,
         \19459 , \19460 , \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 , \19468 ,
         \19469 , \19470 , \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 , \19478 ,
         \19479 , \19480 , \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 , \19488 ,
         \19489 , \19490 , \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 , \19498 ,
         \19499 , \19500 , \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 , \19508 ,
         \19509 , \19510 , \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 , \19518 ,
         \19519 , \19520 , \19521 , \19522 , \19523 , \19524 , \19525 , \19526 , \19527 , \19528 ,
         \19529 , \19530 , \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 , \19538 ,
         \19539 , \19540 , \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 , \19548 ,
         \19549 , \19550 , \19551 , \19552 , \19553 , \19554 , \19555 , \19556 , \19557 , \19558 ,
         \19559 , \19560 , \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 , \19568 ,
         \19569 , \19570 , \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 , \19578 ,
         \19579 , \19580 , \19581 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 , \19588 ,
         \19589 , \19590 , \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 , \19598 ,
         \19599 , \19600 , \19601 , \19602 , \19603 , \19604 , \19605 , \19606 , \19607 , \19608 ,
         \19609 , \19610 , \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 , \19618 ,
         \19619 , \19620 , \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 , \19628 ,
         \19629 , \19630 , \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 , \19638 ,
         \19639 , \19640 , \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 , \19648 ,
         \19649 , \19650 , \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 , \19658 ,
         \19659 , \19660 , \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 , \19668 ,
         \19669 , \19670 , \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 , \19678 ,
         \19679 , \19680 , \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 , \19688 ,
         \19689 , \19690 , \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 , \19698 ,
         \19699 , \19700 , \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 , \19708 ,
         \19709 , \19710 , \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 , \19718 ,
         \19719 , \19720 , \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 , \19728 ,
         \19729 , \19730 , \19731 , \19732 , \19733 , \19734 , \19735 , \19736 , \19737 , \19738 ,
         \19739 , \19740 , \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 , \19748 ,
         \19749 , \19750 , \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 , \19758 ,
         \19759 , \19760 , \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 , \19768 ,
         \19769 , \19770 , \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 , \19778 ,
         \19779 , \19780 , \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 , \19788 ,
         \19789 , \19790 , \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 , \19798 ,
         \19799 , \19800 , \19801 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 , \19808 ,
         \19809 , \19810 , \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 , \19818 ,
         \19819 , \19820 , \19821 , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 , \19828 ,
         \19829 , \19830 , \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 , \19838 ,
         \19839 , \19840 , \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 , \19848 ,
         \19849 , \19850 , \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 , \19858 ,
         \19859 , \19860 , \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 , \19868 ,
         \19869 , \19870 , \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 , \19878 ,
         \19879 , \19880 , \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 , \19888 ,
         \19889 , \19890 , \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 , \19898 ,
         \19899 , \19900 , \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 , \19908 ,
         \19909 , \19910 , \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 , \19918 ,
         \19919 , \19920 , \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 , \19928 ,
         \19929 , \19930 , \19931 , \19932 , \19933 , \19934 , \19935 , \19936 , \19937 , \19938 ,
         \19939 , \19940 , \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 , \19948 ,
         \19949 , \19950 , \19951 , \19952 , \19953 , \19954 , \19955 , \19956 , \19957 , \19958 ,
         \19959 , \19960 , \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 , \19968 ,
         \19969 , \19970 , \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 , \19978 ,
         \19979 , \19980 , \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 , \19988 ,
         \19989 , \19990 , \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 , \19998 ,
         \19999 , \20000 , \20001 , \20002 , \20003 , \20004 , \20005 , \20006 , \20007 , \20008 ,
         \20009 , \20010 , \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 , \20018 ,
         \20019 , \20020 , \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 , \20028 ,
         \20029 , \20030 , \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 , \20038 ,
         \20039 , \20040 , \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 , \20048 ,
         \20049 , \20050 , \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 , \20058 ,
         \20059 , \20060 , \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 , \20068 ,
         \20069 , \20070 , \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 , \20078 ,
         \20079 , \20080 , \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 , \20088 ,
         \20089 , \20090 , \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 , \20098 ,
         \20099 , \20100 , \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 , \20108 ,
         \20109 , \20110 , \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 , \20118 ,
         \20119 , \20120 , \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 , \20128 ,
         \20129 , \20130 , \20131 , \20132 , \20133 , \20134 , \20135 , \20136 , \20137 , \20138 ,
         \20139 , \20140 , \20141 , \20142 , \20143 , \20144 , \20145 , \20146 , \20147 , \20148 ,
         \20149 , \20150 , \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , \20157 , \20158 ,
         \20159 , \20160 , \20161 , \20162 , \20163 , \20164 , \20165 , \20166 , \20167 , \20168 ,
         \20169 , \20170 , \20171 , \20172 , \20173 , \20174 , \20175 , \20176 , \20177 , \20178 ,
         \20179 , \20180 , \20181 , \20182 , \20183 , \20184 , \20185 , \20186 , \20187 , \20188 ,
         \20189 , \20190 , \20191 , \20192 , \20193 , \20194 , \20195 , \20196 , \20197 , \20198 ,
         \20199 , \20200 , \20201 , \20202 , \20203 , \20204 , \20205 , \20206 , \20207 , \20208 ,
         \20209 , \20210 , \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 , \20218 ,
         \20219 , \20220 , \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 , \20228 ,
         \20229 , \20230 , \20231 , \20232 , \20233 , \20234 , \20235 , \20236 , \20237 , \20238 ,
         \20239 , \20240 , \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 , \20248 ,
         \20249 , \20250 , \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 , \20258 ,
         \20259 , \20260 , \20261 , \20262 , \20263 , \20264 , \20265 , \20266 , \20267 , \20268 ,
         \20269 , \20270 , \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 , \20278 ,
         \20279 , \20280 , \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 , \20288 ,
         \20289 , \20290 , \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 , \20298 ,
         \20299 , \20300 , \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 , \20308 ,
         \20309 , \20310 , \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 , \20318 ,
         \20319 , \20320 , \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 , \20328 ,
         \20329 , \20330 , \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 , \20338 ,
         \20339 , \20340 , \20341 , \20342 , \20343 , \20344 , \20345 , \20346 , \20347 , \20348 ,
         \20349 , \20350 , \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 , \20358 ,
         \20359 , \20360 , \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 , \20368 ,
         \20369 , \20370 , \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 , \20378 ,
         \20379 , \20380 , \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 , \20388 ,
         \20389 , \20390 , \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 , \20398 ,
         \20399 , \20400 , \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 , \20408 ,
         \20409 , \20410 , \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 , \20418 ,
         \20419 , \20420 , \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 , \20428 ,
         \20429 , \20430 , \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 , \20438 ,
         \20439 , \20440 , \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 , \20448 ,
         \20449 , \20450 , \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457 , \20458 ,
         \20459 , \20460 , \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 , \20468 ,
         \20469 , \20470 , \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 , \20478 ,
         \20479 , \20480 , \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 , \20488 ,
         \20489 , \20490 , \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 , \20498 ,
         \20499 , \20500 , \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 , \20508 ,
         \20509 , \20510 , \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 , \20518 ,
         \20519 , \20520 , \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 , \20528 ,
         \20529 , \20530 , \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 , \20538 ,
         \20539 , \20540 , \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 , \20548 ,
         \20549 , \20550 , \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 , \20558 ,
         \20559 , \20560 , \20561 , \20562 , \20563 , \20564 , \20565 , \20566 , \20567 , \20568 ,
         \20569 , \20570 , \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 , \20578 ,
         \20579 , \20580 , \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 , \20588 ,
         \20589 , \20590 , \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 , \20598 ,
         \20599 , \20600 , \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 , \20608 ,
         \20609 , \20610 , \20611 , \20612 , \20613 , \20614 , \20615 , \20616 , \20617 , \20618 ,
         \20619 , \20620 , \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 , \20628 ,
         \20629 , \20630 , \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 , \20638 ,
         \20639 , \20640 , \20641 , \20642 , \20643 , \20644 , \20645 , \20646 , \20647 , \20648 ,
         \20649 , \20650 , \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 , \20658 ,
         \20659 , \20660 , \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 , \20668 ,
         \20669 , \20670 , \20671 , \20672 , \20673 , \20674 , \20675 , \20676 , \20677 , \20678 ,
         \20679 , \20680 , \20681 , \20682 , \20683 , \20684 , \20685 , \20686 , \20687 , \20688 ,
         \20689 , \20690 , \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 , \20698 ,
         \20699 , \20700 , \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 , \20708 ,
         \20709 , \20710 , \20711 , \20712 , \20713 , \20714 , \20715 , \20716 , \20717 , \20718 ,
         \20719 , \20720 , \20721 , \20722 , \20723 , \20724 , \20725 , \20726 , \20727 , \20728 ,
         \20729 , \20730 , \20731 , \20732 , \20733 , \20734 , \20735 , \20736 , \20737 , \20738 ,
         \20739 , \20740 , \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 , \20748 ,
         \20749 , \20750 , \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 , \20758 ,
         \20759 , \20760 , \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 , \20768 ,
         \20769 , \20770 , \20771 , \20772 , \20773 , \20774 , \20775 , \20776 , \20777 , \20778 ,
         \20779 , \20780 , \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 , \20788 ,
         \20789 , \20790 , \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 , \20798 ,
         \20799 , \20800 , \20801 , \20802 , \20803 , \20804 , \20805 , \20806 , \20807 , \20808 ,
         \20809 , \20810 , \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 , \20818 ,
         \20819 , \20820 , \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 , \20828 ,
         \20829 , \20830 , \20831 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 , \20838 ,
         \20839 , \20840 , \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 , \20848 ,
         \20849 , \20850 , \20851 , \20852 , \20853 , \20854 , \20855 , \20856 , \20857 , \20858 ,
         \20859 , \20860 , \20861 , \20862 , \20863 , \20864 , \20865 , \20866 , \20867 , \20868 ,
         \20869 , \20870 , \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 , \20878 ,
         \20879 , \20880 , \20881 , \20882 , \20883 , \20884 , \20885 , \20886 , \20887 , \20888 ,
         \20889 , \20890 , \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 , \20898 ,
         \20899 , \20900 , \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 , \20908 ,
         \20909 , \20910 , \20911 , \20912 , \20913 , \20914 , \20915 , \20916 , \20917 , \20918 ,
         \20919 , \20920 , \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 , \20928 ,
         \20929 , \20930 , \20931 , \20932 , \20933 , \20934 , \20935 , \20936 , \20937 , \20938 ,
         \20939 , \20940 , \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 , \20948 ,
         \20949 , \20950 , \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 , \20958 ,
         \20959 , \20960 , \20961 , \20962 , \20963 , \20964 , \20965 , \20966 , \20967 , \20968 ,
         \20969 , \20970 , \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 , \20978 ,
         \20979 , \20980 , \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 , \20988 ,
         \20989 , \20990 , \20991 , \20992 , \20993 , \20994 , \20995 , \20996 , \20997 , \20998 ,
         \20999 , \21000 , \21001 , \21002 , \21003 , \21004 , \21005 , \21006 , \21007 , \21008 ,
         \21009 , \21010 , \21011 , \21012 , \21013 , \21014 , \21015 , \21016 , \21017 , \21018 ,
         \21019 , \21020 , \21021 , \21022 , \21023 , \21024 , \21025 , \21026 , \21027 , \21028 ,
         \21029 , \21030 , \21031 , \21032 , \21033 , \21034 , \21035 , \21036 , \21037 , \21038 ,
         \21039 , \21040 , \21041 , \21042 , \21043 , \21044 , \21045 , \21046 , \21047 , \21048 ,
         \21049 , \21050 , \21051 , \21052 , \21053 , \21054 , \21055 , \21056 , \21057 , \21058 ,
         \21059 , \21060 , \21061 , \21062 , \21063 , \21064 , \21065 , \21066 , \21067 , \21068 ,
         \21069 , \21070 , \21071 , \21072 , \21073 , \21074 , \21075 , \21076 , \21077 , \21078 ,
         \21079 , \21080 , \21081 , \21082 , \21083 , \21084 , \21085 , \21086 , \21087 , \21088 ,
         \21089 , \21090 , \21091 , \21092 , \21093 , \21094 , \21095 , \21096 , \21097 , \21098 ,
         \21099 , \21100 , \21101 , \21102 , \21103 , \21104 , \21105 , \21106 , \21107 , \21108 ,
         \21109 , \21110 , \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 , \21118 ,
         \21119 , \21120 , \21121 , \21122 , \21123 , \21124 , \21125 , \21126 , \21127 , \21128 ,
         \21129 , \21130 , \21131 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 , \21138 ,
         \21139 , \21140 , \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 , \21148 ,
         \21149 , \21150 , \21151 , \21152 , \21153 , \21154 , \21155 , \21156 , \21157 , \21158 ,
         \21159 , \21160 , \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 , \21168 ,
         \21169 , \21170 , \21171 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 , \21178 ,
         \21179 , \21180 , \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 , \21188 ,
         \21189 , \21190 , \21191 , \21192 , \21193 , \21194 , \21195 , \21196 , \21197 , \21198 ,
         \21199 , \21200 , \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207 , \21208 ,
         \21209 , \21210 , \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 , \21218 ,
         \21219 , \21220 , \21221 , \21222 , \21223 , \21224 , \21225 , \21226 , \21227 , \21228 ,
         \21229 , \21230 , \21231 , \21232 , \21233 , \21234 , \21235 , \21236 , \21237 , \21238 ,
         \21239 , \21240 , \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 , \21248 ,
         \21249 , \21250 , \21251 , \21252 , \21253 , \21254 , \21255 , \21256 , \21257 , \21258 ,
         \21259 , \21260 , \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 , \21268 ,
         \21269 , \21270 , \21271 , \21272 , \21273 , \21274 , \21275 , \21276 , \21277 , \21278 ,
         \21279 , \21280 , \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 , \21288 ,
         \21289 , \21290 , \21291 , \21292 , \21293 , \21294 , \21295 , \21296 , \21297 , \21298 ,
         \21299 , \21300 , \21301 , \21302 , \21303 , \21304 , \21305 , \21306 , \21307 , \21308 ,
         \21309 , \21310 , \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 , \21318 ,
         \21319 , \21320 , \21321 , \21322 , \21323 , \21324 , \21325 , \21326 , \21327 , \21328 ,
         \21329 , \21330 , \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 , \21338 ,
         \21339 , \21340 , \21341 , \21342 , \21343 , \21344 , \21345 , \21346 , \21347 , \21348 ,
         \21349 , \21350 , \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 , \21358 ,
         \21359 , \21360 , \21361 , \21362 , \21363 , \21364 , \21365 , \21366 , \21367 , \21368 ,
         \21369 , \21370 , \21371 , \21372 , \21373 , \21374 , \21375 , \21376 , \21377 , \21378 ,
         \21379 , \21380 , \21381 , \21382 , \21383 , \21384 , \21385 , \21386 , \21387 , \21388 ,
         \21389 , \21390 , \21391 , \21392 , \21393 , \21394 , \21395 , \21396 , \21397 , \21398 ,
         \21399 , \21400 , \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 , \21408 ,
         \21409 , \21410 , \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 , \21418 ,
         \21419 , \21420 , \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 , \21428 ,
         \21429 , \21430 , \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 , \21438 ,
         \21439 , \21440 , \21441 , \21442 , \21443 , \21444 , \21445 , \21446 , \21447 , \21448 ,
         \21449 , \21450 , \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 , \21458 ,
         \21459 , \21460 , \21461 , \21462 , \21463 , \21464 , \21465 , \21466 , \21467 , \21468 ,
         \21469 , \21470 , \21471 , \21472 , \21473 , \21474 , \21475 , \21476 , \21477 , \21478 ,
         \21479 , \21480 , \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 , \21488 ,
         \21489 , \21490 , \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 , \21498 ,
         \21499 , \21500 , \21501 , \21502 , \21503 , \21504 , \21505 , \21506 , \21507 , \21508 ,
         \21509 , \21510 , \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517 , \21518 ,
         \21519 , \21520 , \21521 , \21522 , \21523 , \21524 , \21525 , \21526 , \21527 , \21528 ,
         \21529 , \21530 , \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 , \21538 ,
         \21539 , \21540 , \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 , \21548 ,
         \21549 , \21550 , \21551 , \21552 , \21553 , \21554 , \21555 , \21556 , \21557 , \21558 ,
         \21559 , \21560 , \21561 , \21562 , \21563 , \21564 , \21565 , \21566 , \21567 , \21568 ,
         \21569 , \21570 , \21571 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 , \21578 ,
         \21579 , \21580 , \21581 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 , \21588 ,
         \21589 , \21590 , \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 , \21598 ,
         \21599 , \21600 , \21601 , \21602 , \21603 , \21604 , \21605 , \21606 , \21607 , \21608 ,
         \21609 , \21610 , \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 , \21618 ,
         \21619 , \21620 , \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 , \21628 ,
         \21629 , \21630 , \21631 , \21632 , \21633 , \21634 , \21635 , \21636 , \21637 , \21638 ,
         \21639 , \21640 , \21641 , \21642 , \21643 , \21644 , \21645 , \21646 , \21647 , \21648 ,
         \21649 , \21650 , \21651 , \21652 , \21653 , \21654 , \21655 , \21656 , \21657 , \21658 ,
         \21659 , \21660 , \21661 , \21662 , \21663 , \21664 , \21665 , \21666 , \21667 , \21668 ,
         \21669 , \21670 , \21671 , \21672 , \21673 , \21674 , \21675 , \21676 , \21677 , \21678 ,
         \21679 , \21680 , \21681 , \21682 , \21683 , \21684 , \21685 , \21686 , \21687 , \21688 ,
         \21689 , \21690 , \21691 , \21692 , \21693 , \21694 , \21695 , \21696 , \21697 , \21698 ,
         \21699 , \21700 , \21701 , \21702 , \21703 , \21704 , \21705 , \21706 , \21707 , \21708 ,
         \21709 , \21710 , \21711 , \21712 , \21713 , \21714 , \21715 , \21716 , \21717 , \21718 ,
         \21719 , \21720 , \21721 , \21722 , \21723 , \21724 , \21725 , \21726 , \21727 , \21728 ,
         \21729 , \21730 , \21731 , \21732 , \21733 , \21734 , \21735 , \21736 , \21737 , \21738 ,
         \21739 , \21740 , \21741 , \21742 , \21743 , \21744 , \21745 , \21746 , \21747 , \21748 ,
         \21749 , \21750 , \21751 , \21752 , \21753 , \21754 , \21755 , \21756 , \21757 , \21758 ,
         \21759 , \21760 , \21761 , \21762 , \21763 , \21764 , \21765 , \21766 , \21767 , \21768 ,
         \21769 , \21770 , \21771 , \21772 , \21773 , \21774 , \21775 , \21776 , \21777 , \21778 ,
         \21779 , \21780 , \21781 , \21782 , \21783 , \21784 , \21785 , \21786 , \21787 , \21788 ,
         \21789 , \21790 , \21791 , \21792 , \21793 , \21794 , \21795 , \21796 , \21797 , \21798 ,
         \21799 , \21800 , \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 ,
         \21809 , \21810 , \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 ,
         \21819 , \21820 , \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 , \21828 ,
         \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 ,
         \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 ,
         \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 ,
         \21859 , \21860 , \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 , \21868 ,
         \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 ,
         \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 ,
         \21889 , \21890 , \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 , \21898 ,
         \21899 , \21900 , \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 , \21908 ,
         \21909 , \21910 , \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 , \21918 ,
         \21919 , \21920 , \21921 , \21922 , \21923 , \21924 , \21925 , \21926 , \21927 , \21928 ,
         \21929 , \21930 , \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937_nR56af , \21938 ;
buf \U$labaj2213 ( R_81_7e072f0, \21938 );
buf \U$2 ( \134 , RIb559478_125);
buf \U$3 ( \135 , RIb55f760_53);
buf \U$4 ( \136 , RIb55f6e8_54);
xor \U$5 ( \137 , \135 , \136 );
buf \U$6 ( \138 , RIb55f670_55);
xor \U$7 ( \139 , \136 , \138 );
not \U$8 ( \140 , \139 );
and \U$9 ( \141 , \137 , \140 );
and \U$10 ( \142 , \134 , \141 );
buf \U$11 ( \143 , RIb5594f0_124);
and \U$12 ( \144 , \143 , \139 );
nor \U$13 ( \145 , \142 , \144 );
and \U$14 ( \146 , \136 , \138 );
not \U$15 ( \147 , \146 );
and \U$16 ( \148 , \135 , \147 );
xnor \U$17 ( \149 , \145 , \148 );
buf \U$18 ( \150 , RIb559388_127);
buf \U$19 ( \151 , RIb55f850_51);
buf \U$20 ( \152 , RIb55f7d8_52);
xor \U$21 ( \153 , \151 , \152 );
xor \U$22 ( \154 , \152 , \135 );
not \U$23 ( \155 , \154 );
and \U$24 ( \156 , \153 , \155 );
and \U$25 ( \157 , \150 , \156 );
buf \U$26 ( \158 , RIb559400_126);
and \U$27 ( \159 , \158 , \154 );
nor \U$28 ( \160 , \157 , \159 );
and \U$29 ( \161 , \152 , \135 );
not \U$30 ( \162 , \161 );
and \U$31 ( \163 , \151 , \162 );
xnor \U$32 ( \164 , \160 , \163 );
and \U$33 ( \165 , \149 , \164 );
buf \U$34 ( \166 , RIb559310_128);
buf \U$35 ( \167 , RIb55f8c8_50);
xor \U$36 ( \168 , \167 , \151 );
nand \U$37 ( \169 , \166 , \168 );
buf \U$38 ( \170 , RIb55f940_49);
and \U$39 ( \171 , \167 , \151 );
not \U$40 ( \172 , \171 );
and \U$41 ( \173 , \170 , \172 );
xnor \U$42 ( \174 , \169 , \173 );
and \U$43 ( \175 , \164 , \174 );
and \U$44 ( \176 , \149 , \174 );
or \U$45 ( \177 , \165 , \175 , \176 );
buf \U$46 ( \178 , RIb55da50_115);
buf \U$47 ( \179 , RIb55f2b0_63);
buf \U$48 ( \180 , RIb55f238_64);
xor \U$49 ( \181 , \179 , \180 );
not \U$50 ( \182 , \180 );
and \U$51 ( \183 , \181 , \182 );
and \U$52 ( \184 , \178 , \183 );
buf \U$53 ( \185 , RIb55dac8_114);
and \U$54 ( \186 , \185 , \180 );
nor \U$55 ( \187 , \184 , \186 );
xnor \U$56 ( \188 , \187 , \179 );
buf \U$57 ( \189 , RIb55d960_117);
buf \U$58 ( \190 , RIb55f3a0_61);
buf \U$59 ( \191 , RIb55f328_62);
xor \U$60 ( \192 , \190 , \191 );
xor \U$61 ( \193 , \191 , \179 );
not \U$62 ( \194 , \193 );
and \U$63 ( \195 , \192 , \194 );
and \U$64 ( \196 , \189 , \195 );
buf \U$65 ( \197 , RIb55d9d8_116);
and \U$66 ( \198 , \197 , \193 );
nor \U$67 ( \199 , \196 , \198 );
and \U$68 ( \200 , \191 , \179 );
not \U$69 ( \201 , \200 );
and \U$70 ( \202 , \190 , \201 );
xnor \U$71 ( \203 , \199 , \202 );
and \U$72 ( \204 , \188 , \203 );
and \U$73 ( \205 , \203 , \173 );
and \U$74 ( \206 , \188 , \173 );
or \U$75 ( \207 , \204 , \205 , \206 );
and \U$76 ( \208 , \177 , \207 );
buf \U$77 ( \209 , RIb55d870_119);
buf \U$78 ( \210 , RIb55f490_59);
buf \U$79 ( \211 , RIb55f418_60);
xor \U$80 ( \212 , \210 , \211 );
xor \U$81 ( \213 , \211 , \190 );
not \U$82 ( \214 , \213 );
and \U$83 ( \215 , \212 , \214 );
and \U$84 ( \216 , \209 , \215 );
buf \U$85 ( \217 , RIb55d8e8_118);
and \U$86 ( \218 , \217 , \213 );
nor \U$87 ( \219 , \216 , \218 );
and \U$88 ( \220 , \211 , \190 );
not \U$89 ( \221 , \220 );
and \U$90 ( \222 , \210 , \221 );
xnor \U$91 ( \223 , \219 , \222 );
buf \U$92 ( \224 , RIb55d780_121);
buf \U$93 ( \225 , RIb55f580_57);
buf \U$94 ( \226 , RIb55f508_58);
xor \U$95 ( \227 , \225 , \226 );
xor \U$96 ( \228 , \226 , \210 );
not \U$97 ( \229 , \228 );
and \U$98 ( \230 , \227 , \229 );
and \U$99 ( \231 , \224 , \230 );
buf \U$100 ( \232 , RIb55d7f8_120);
and \U$101 ( \233 , \232 , \228 );
nor \U$102 ( \234 , \231 , \233 );
and \U$103 ( \235 , \226 , \210 );
not \U$104 ( \236 , \235 );
and \U$105 ( \237 , \225 , \236 );
xnor \U$106 ( \238 , \234 , \237 );
and \U$107 ( \239 , \223 , \238 );
buf \U$108 ( \240 , RIb55d690_123);
buf \U$109 ( \241 , RIb55f5f8_56);
xor \U$110 ( \242 , \138 , \241 );
xor \U$111 ( \243 , \241 , \225 );
not \U$112 ( \244 , \243 );
and \U$113 ( \245 , \242 , \244 );
and \U$114 ( \246 , \240 , \245 );
buf \U$115 ( \247 , RIb55d708_122);
and \U$116 ( \248 , \247 , \243 );
nor \U$117 ( \249 , \246 , \248 );
and \U$118 ( \250 , \241 , \225 );
not \U$119 ( \251 , \250 );
and \U$120 ( \252 , \138 , \251 );
xnor \U$121 ( \253 , \249 , \252 );
and \U$122 ( \254 , \238 , \253 );
and \U$123 ( \255 , \223 , \253 );
or \U$124 ( \256 , \239 , \254 , \255 );
and \U$125 ( \257 , \207 , \256 );
and \U$126 ( \258 , \177 , \256 );
or \U$127 ( \259 , \208 , \257 , \258 );
and \U$128 ( \260 , \185 , \183 );
buf \U$129 ( \261 , RIb55db40_113);
and \U$130 ( \262 , \261 , \180 );
nor \U$131 ( \263 , \260 , \262 );
xnor \U$132 ( \264 , \263 , \179 );
and \U$133 ( \265 , \197 , \195 );
and \U$134 ( \266 , \178 , \193 );
nor \U$135 ( \267 , \265 , \266 );
xnor \U$136 ( \268 , \267 , \202 );
xor \U$137 ( \269 , \264 , \268 );
and \U$138 ( \270 , \217 , \215 );
and \U$139 ( \271 , \189 , \213 );
nor \U$140 ( \272 , \270 , \271 );
xnor \U$141 ( \273 , \272 , \222 );
xor \U$142 ( \274 , \269 , \273 );
and \U$143 ( \275 , \232 , \230 );
and \U$144 ( \276 , \209 , \228 );
nor \U$145 ( \277 , \275 , \276 );
xnor \U$146 ( \278 , \277 , \237 );
and \U$147 ( \279 , \247 , \245 );
and \U$148 ( \280 , \224 , \243 );
nor \U$149 ( \281 , \279 , \280 );
xnor \U$150 ( \282 , \281 , \252 );
xor \U$151 ( \283 , \278 , \282 );
and \U$152 ( \284 , \143 , \141 );
and \U$153 ( \285 , \240 , \139 );
nor \U$154 ( \286 , \284 , \285 );
xnor \U$155 ( \287 , \286 , \148 );
xor \U$156 ( \288 , \283 , \287 );
and \U$157 ( \289 , \274 , \288 );
and \U$158 ( \290 , \158 , \156 );
and \U$159 ( \291 , \134 , \154 );
nor \U$160 ( \292 , \290 , \291 );
xnor \U$161 ( \293 , \292 , \163 );
xor \U$162 ( \294 , \170 , \167 );
not \U$163 ( \295 , \168 );
and \U$164 ( \296 , \294 , \295 );
and \U$165 ( \297 , \166 , \296 );
and \U$166 ( \298 , \150 , \168 );
nor \U$167 ( \299 , \297 , \298 );
xnor \U$168 ( \300 , \299 , \173 );
xor \U$169 ( \301 , \293 , \300 );
and \U$170 ( \302 , \288 , \301 );
and \U$171 ( \303 , \274 , \301 );
or \U$172 ( \304 , \289 , \302 , \303 );
and \U$173 ( \305 , \259 , \304 );
and \U$174 ( \306 , \261 , \183 );
buf \U$175 ( \307 , RIb55dbb8_112);
and \U$176 ( \308 , \307 , \180 );
nor \U$177 ( \309 , \306 , \308 );
xnor \U$178 ( \310 , \309 , \179 );
and \U$179 ( \311 , \178 , \195 );
and \U$180 ( \312 , \185 , \193 );
nor \U$181 ( \313 , \311 , \312 );
xnor \U$182 ( \314 , \313 , \202 );
xor \U$183 ( \315 , \310 , \314 );
buf \U$184 ( \316 , RIb55fa30_47);
buf \U$185 ( \317 , RIb55f9b8_48);
and \U$186 ( \318 , \317 , \170 );
not \U$187 ( \319 , \318 );
and \U$188 ( \320 , \316 , \319 );
xor \U$189 ( \321 , \315 , \320 );
and \U$190 ( \322 , \304 , \321 );
and \U$191 ( \323 , \259 , \321 );
or \U$192 ( \324 , \305 , \322 , \323 );
and \U$193 ( \325 , \264 , \268 );
and \U$194 ( \326 , \268 , \273 );
and \U$195 ( \327 , \264 , \273 );
or \U$196 ( \328 , \325 , \326 , \327 );
and \U$197 ( \329 , \278 , \282 );
and \U$198 ( \330 , \282 , \287 );
and \U$199 ( \331 , \278 , \287 );
or \U$200 ( \332 , \329 , \330 , \331 );
xor \U$201 ( \333 , \328 , \332 );
and \U$202 ( \334 , \293 , \300 );
xor \U$203 ( \335 , \333 , \334 );
xor \U$204 ( \336 , \317 , \170 );
nand \U$205 ( \337 , \166 , \336 );
xnor \U$206 ( \338 , \337 , \320 );
and \U$207 ( \339 , \189 , \215 );
and \U$208 ( \340 , \197 , \213 );
nor \U$209 ( \341 , \339 , \340 );
xnor \U$210 ( \342 , \341 , \222 );
and \U$211 ( \343 , \209 , \230 );
and \U$212 ( \344 , \217 , \228 );
nor \U$213 ( \345 , \343 , \344 );
xnor \U$214 ( \346 , \345 , \237 );
xor \U$215 ( \347 , \342 , \346 );
and \U$216 ( \348 , \224 , \245 );
and \U$217 ( \349 , \232 , \243 );
nor \U$218 ( \350 , \348 , \349 );
xnor \U$219 ( \351 , \350 , \252 );
xor \U$220 ( \352 , \347 , \351 );
xor \U$221 ( \353 , \338 , \352 );
and \U$222 ( \354 , \240 , \141 );
and \U$223 ( \355 , \247 , \139 );
nor \U$224 ( \356 , \354 , \355 );
xnor \U$225 ( \357 , \356 , \148 );
and \U$226 ( \358 , \134 , \156 );
and \U$227 ( \359 , \143 , \154 );
nor \U$228 ( \360 , \358 , \359 );
xnor \U$229 ( \361 , \360 , \163 );
xor \U$230 ( \362 , \357 , \361 );
and \U$231 ( \363 , \150 , \296 );
and \U$232 ( \364 , \158 , \168 );
nor \U$233 ( \365 , \363 , \364 );
xnor \U$234 ( \366 , \365 , \173 );
xor \U$235 ( \367 , \362 , \366 );
xor \U$236 ( \368 , \353 , \367 );
and \U$237 ( \369 , \335 , \368 );
and \U$238 ( \370 , \324 , \369 );
and \U$239 ( \371 , \342 , \346 );
and \U$240 ( \372 , \346 , \351 );
and \U$241 ( \373 , \342 , \351 );
or \U$242 ( \374 , \371 , \372 , \373 );
and \U$243 ( \375 , \310 , \314 );
and \U$244 ( \376 , \314 , \320 );
and \U$245 ( \377 , \310 , \320 );
or \U$246 ( \378 , \375 , \376 , \377 );
xor \U$247 ( \379 , \374 , \378 );
and \U$248 ( \380 , \357 , \361 );
and \U$249 ( \381 , \361 , \366 );
and \U$250 ( \382 , \357 , \366 );
or \U$251 ( \383 , \380 , \381 , \382 );
xor \U$252 ( \384 , \379 , \383 );
and \U$253 ( \385 , \369 , \384 );
and \U$254 ( \386 , \324 , \384 );
or \U$255 ( \387 , \370 , \385 , \386 );
and \U$256 ( \388 , \328 , \332 );
and \U$257 ( \389 , \332 , \334 );
and \U$258 ( \390 , \328 , \334 );
or \U$259 ( \391 , \388 , \389 , \390 );
and \U$260 ( \392 , \338 , \352 );
and \U$261 ( \393 , \352 , \367 );
and \U$262 ( \394 , \338 , \367 );
or \U$263 ( \395 , \392 , \393 , \394 );
and \U$264 ( \396 , \391 , \395 );
and \U$265 ( \397 , \217 , \230 );
and \U$266 ( \398 , \189 , \228 );
nor \U$267 ( \399 , \397 , \398 );
xnor \U$268 ( \400 , \399 , \237 );
and \U$269 ( \401 , \232 , \245 );
and \U$270 ( \402 , \209 , \243 );
nor \U$271 ( \403 , \401 , \402 );
xnor \U$272 ( \404 , \403 , \252 );
xor \U$273 ( \405 , \400 , \404 );
and \U$274 ( \406 , \247 , \141 );
and \U$275 ( \407 , \224 , \139 );
nor \U$276 ( \408 , \406 , \407 );
xnor \U$277 ( \409 , \408 , \148 );
xor \U$278 ( \410 , \405 , \409 );
and \U$279 ( \411 , \307 , \183 );
buf \U$280 ( \412 , RIb55dc30_111);
and \U$281 ( \413 , \412 , \180 );
nor \U$282 ( \414 , \411 , \413 );
xnor \U$283 ( \415 , \414 , \179 );
and \U$284 ( \416 , \185 , \195 );
and \U$285 ( \417 , \261 , \193 );
nor \U$286 ( \418 , \416 , \417 );
xnor \U$287 ( \419 , \418 , \202 );
xor \U$288 ( \420 , \415 , \419 );
and \U$289 ( \421 , \197 , \215 );
and \U$290 ( \422 , \178 , \213 );
nor \U$291 ( \423 , \421 , \422 );
xnor \U$292 ( \424 , \423 , \222 );
xor \U$293 ( \425 , \420 , \424 );
xor \U$294 ( \426 , \410 , \425 );
and \U$295 ( \427 , \143 , \156 );
and \U$296 ( \428 , \240 , \154 );
nor \U$297 ( \429 , \427 , \428 );
xnor \U$298 ( \430 , \429 , \163 );
and \U$299 ( \431 , \158 , \296 );
and \U$300 ( \432 , \134 , \168 );
nor \U$301 ( \433 , \431 , \432 );
xnor \U$302 ( \434 , \433 , \173 );
xor \U$303 ( \435 , \430 , \434 );
xor \U$304 ( \436 , \316 , \317 );
not \U$305 ( \437 , \336 );
and \U$306 ( \438 , \436 , \437 );
and \U$307 ( \439 , \166 , \438 );
and \U$308 ( \440 , \150 , \336 );
nor \U$309 ( \441 , \439 , \440 );
xnor \U$310 ( \442 , \441 , \320 );
xor \U$311 ( \443 , \435 , \442 );
xor \U$312 ( \444 , \426 , \443 );
and \U$313 ( \445 , \395 , \444 );
and \U$314 ( \446 , \391 , \444 );
or \U$315 ( \447 , \396 , \445 , \446 );
and \U$316 ( \448 , \374 , \378 );
and \U$317 ( \449 , \378 , \383 );
and \U$318 ( \450 , \374 , \383 );
or \U$319 ( \451 , \448 , \449 , \450 );
and \U$320 ( \452 , \410 , \425 );
and \U$321 ( \453 , \425 , \443 );
and \U$322 ( \454 , \410 , \443 );
or \U$323 ( \455 , \452 , \453 , \454 );
xor \U$324 ( \456 , \451 , \455 );
and \U$325 ( \457 , \178 , \215 );
and \U$326 ( \458 , \185 , \213 );
nor \U$327 ( \459 , \457 , \458 );
xnor \U$328 ( \460 , \459 , \222 );
and \U$329 ( \461 , \189 , \230 );
and \U$330 ( \462 , \197 , \228 );
nor \U$331 ( \463 , \461 , \462 );
xnor \U$332 ( \464 , \463 , \237 );
xor \U$333 ( \465 , \460 , \464 );
and \U$334 ( \466 , \209 , \245 );
and \U$335 ( \467 , \217 , \243 );
nor \U$336 ( \468 , \466 , \467 );
xnor \U$337 ( \469 , \468 , \252 );
xor \U$338 ( \470 , \465 , \469 );
xor \U$339 ( \471 , \456 , \470 );
xor \U$340 ( \472 , \447 , \471 );
and \U$341 ( \473 , \412 , \183 );
buf \U$342 ( \474 , RIb55dca8_110);
and \U$343 ( \475 , \474 , \180 );
nor \U$344 ( \476 , \473 , \475 );
xnor \U$345 ( \477 , \476 , \179 );
and \U$346 ( \478 , \261 , \195 );
and \U$347 ( \479 , \307 , \193 );
nor \U$348 ( \480 , \478 , \479 );
xnor \U$349 ( \481 , \480 , \202 );
xor \U$350 ( \482 , \477 , \481 );
buf \U$351 ( \483 , RIb55fb20_45);
buf \U$352 ( \484 , RIb55faa8_46);
and \U$353 ( \485 , \484 , \316 );
not \U$354 ( \486 , \485 );
and \U$355 ( \487 , \483 , \486 );
xor \U$356 ( \488 , \482 , \487 );
and \U$357 ( \489 , \400 , \404 );
and \U$358 ( \490 , \404 , \409 );
and \U$359 ( \491 , \400 , \409 );
or \U$360 ( \492 , \489 , \490 , \491 );
and \U$361 ( \493 , \415 , \419 );
and \U$362 ( \494 , \419 , \424 );
and \U$363 ( \495 , \415 , \424 );
or \U$364 ( \496 , \493 , \494 , \495 );
xor \U$365 ( \497 , \492 , \496 );
and \U$366 ( \498 , \430 , \434 );
and \U$367 ( \499 , \434 , \442 );
and \U$368 ( \500 , \430 , \442 );
or \U$369 ( \501 , \498 , \499 , \500 );
xor \U$370 ( \502 , \497 , \501 );
xor \U$371 ( \503 , \488 , \502 );
and \U$372 ( \504 , \150 , \438 );
and \U$373 ( \505 , \158 , \336 );
nor \U$374 ( \506 , \504 , \505 );
xnor \U$375 ( \507 , \506 , \320 );
xor \U$376 ( \508 , \484 , \316 );
nand \U$377 ( \509 , \166 , \508 );
xnor \U$378 ( \510 , \509 , \487 );
xor \U$379 ( \511 , \507 , \510 );
and \U$380 ( \512 , \224 , \141 );
and \U$381 ( \513 , \232 , \139 );
nor \U$382 ( \514 , \512 , \513 );
xnor \U$383 ( \515 , \514 , \148 );
and \U$384 ( \516 , \240 , \156 );
and \U$385 ( \517 , \247 , \154 );
nor \U$386 ( \518 , \516 , \517 );
xnor \U$387 ( \519 , \518 , \163 );
xor \U$388 ( \520 , \515 , \519 );
and \U$389 ( \521 , \134 , \296 );
and \U$390 ( \522 , \143 , \168 );
nor \U$391 ( \523 , \521 , \522 );
xnor \U$392 ( \524 , \523 , \173 );
xor \U$393 ( \525 , \520 , \524 );
xor \U$394 ( \526 , \511 , \525 );
xor \U$395 ( \527 , \503 , \526 );
xor \U$396 ( \528 , \472 , \527 );
xor \U$397 ( \529 , \387 , \528 );
xor \U$398 ( \530 , \324 , \369 );
xor \U$399 ( \531 , \530 , \384 );
xor \U$400 ( \532 , \391 , \395 );
xor \U$401 ( \533 , \532 , \444 );
and \U$402 ( \534 , \531 , \533 );
xor \U$403 ( \535 , \529 , \534 );
xor \U$404 ( \536 , \531 , \533 );
and \U$405 ( \537 , \197 , \183 );
and \U$406 ( \538 , \178 , \180 );
nor \U$407 ( \539 , \537 , \538 );
xnor \U$408 ( \540 , \539 , \179 );
and \U$409 ( \541 , \217 , \195 );
and \U$410 ( \542 , \189 , \193 );
nor \U$411 ( \543 , \541 , \542 );
xnor \U$412 ( \544 , \543 , \202 );
and \U$413 ( \545 , \540 , \544 );
and \U$414 ( \546 , \232 , \215 );
and \U$415 ( \547 , \209 , \213 );
nor \U$416 ( \548 , \546 , \547 );
xnor \U$417 ( \549 , \548 , \222 );
and \U$418 ( \550 , \544 , \549 );
and \U$419 ( \551 , \540 , \549 );
or \U$420 ( \552 , \545 , \550 , \551 );
and \U$421 ( \553 , \247 , \230 );
and \U$422 ( \554 , \224 , \228 );
nor \U$423 ( \555 , \553 , \554 );
xnor \U$424 ( \556 , \555 , \237 );
and \U$425 ( \557 , \143 , \245 );
and \U$426 ( \558 , \240 , \243 );
nor \U$427 ( \559 , \557 , \558 );
xnor \U$428 ( \560 , \559 , \252 );
and \U$429 ( \561 , \556 , \560 );
and \U$430 ( \562 , \158 , \141 );
and \U$431 ( \563 , \134 , \139 );
nor \U$432 ( \564 , \562 , \563 );
xnor \U$433 ( \565 , \564 , \148 );
and \U$434 ( \566 , \560 , \565 );
and \U$435 ( \567 , \556 , \565 );
or \U$436 ( \568 , \561 , \566 , \567 );
and \U$437 ( \569 , \552 , \568 );
xor \U$438 ( \570 , \149 , \164 );
xor \U$439 ( \571 , \570 , \174 );
and \U$440 ( \572 , \568 , \571 );
and \U$441 ( \573 , \552 , \571 );
or \U$442 ( \574 , \569 , \572 , \573 );
xor \U$443 ( \575 , \188 , \203 );
xor \U$444 ( \576 , \575 , \173 );
xor \U$445 ( \577 , \223 , \238 );
xor \U$446 ( \578 , \577 , \253 );
and \U$447 ( \579 , \576 , \578 );
and \U$448 ( \580 , \574 , \579 );
xor \U$449 ( \581 , \274 , \288 );
xor \U$450 ( \582 , \581 , \301 );
and \U$451 ( \583 , \579 , \582 );
and \U$452 ( \584 , \574 , \582 );
or \U$453 ( \585 , \580 , \583 , \584 );
xor \U$454 ( \586 , \259 , \304 );
xor \U$455 ( \587 , \586 , \321 );
and \U$456 ( \588 , \585 , \587 );
xor \U$457 ( \589 , \335 , \368 );
and \U$458 ( \590 , \587 , \589 );
and \U$459 ( \591 , \585 , \589 );
or \U$460 ( \592 , \588 , \590 , \591 );
and \U$461 ( \593 , \536 , \592 );
xor \U$462 ( \594 , \536 , \592 );
xor \U$463 ( \595 , \585 , \587 );
xor \U$464 ( \596 , \595 , \589 );
and \U$465 ( \597 , \189 , \183 );
and \U$466 ( \598 , \197 , \180 );
nor \U$467 ( \599 , \597 , \598 );
xnor \U$468 ( \600 , \599 , \179 );
and \U$469 ( \601 , \209 , \195 );
and \U$470 ( \602 , \217 , \193 );
nor \U$471 ( \603 , \601 , \602 );
xnor \U$472 ( \604 , \603 , \202 );
and \U$473 ( \605 , \600 , \604 );
and \U$474 ( \606 , \604 , \163 );
and \U$475 ( \607 , \600 , \163 );
or \U$476 ( \608 , \605 , \606 , \607 );
and \U$477 ( \609 , \224 , \215 );
and \U$478 ( \610 , \232 , \213 );
nor \U$479 ( \611 , \609 , \610 );
xnor \U$480 ( \612 , \611 , \222 );
and \U$481 ( \613 , \240 , \230 );
and \U$482 ( \614 , \247 , \228 );
nor \U$483 ( \615 , \613 , \614 );
xnor \U$484 ( \616 , \615 , \237 );
and \U$485 ( \617 , \612 , \616 );
and \U$486 ( \618 , \134 , \245 );
and \U$487 ( \619 , \143 , \243 );
nor \U$488 ( \620 , \618 , \619 );
xnor \U$489 ( \621 , \620 , \252 );
and \U$490 ( \622 , \616 , \621 );
and \U$491 ( \623 , \612 , \621 );
or \U$492 ( \624 , \617 , \622 , \623 );
and \U$493 ( \625 , \608 , \624 );
and \U$494 ( \626 , \166 , \156 );
and \U$495 ( \627 , \150 , \154 );
nor \U$496 ( \628 , \626 , \627 );
xnor \U$497 ( \629 , \628 , \163 );
and \U$498 ( \630 , \624 , \629 );
and \U$499 ( \631 , \608 , \629 );
or \U$500 ( \632 , \625 , \630 , \631 );
xor \U$501 ( \633 , \552 , \568 );
xor \U$502 ( \634 , \633 , \571 );
and \U$503 ( \635 , \632 , \634 );
xor \U$504 ( \636 , \576 , \578 );
and \U$505 ( \637 , \634 , \636 );
and \U$506 ( \638 , \632 , \636 );
or \U$507 ( \639 , \635 , \637 , \638 );
xor \U$508 ( \640 , \177 , \207 );
xor \U$509 ( \641 , \640 , \256 );
and \U$510 ( \642 , \639 , \641 );
xor \U$511 ( \643 , \574 , \579 );
xor \U$512 ( \644 , \643 , \582 );
and \U$513 ( \645 , \641 , \644 );
and \U$514 ( \646 , \639 , \644 );
or \U$515 ( \647 , \642 , \645 , \646 );
and \U$516 ( \648 , \596 , \647 );
xor \U$517 ( \649 , \596 , \647 );
xor \U$518 ( \650 , \639 , \641 );
xor \U$519 ( \651 , \650 , \644 );
and \U$520 ( \652 , \143 , \230 );
and \U$521 ( \653 , \240 , \228 );
nor \U$522 ( \654 , \652 , \653 );
xnor \U$523 ( \655 , \654 , \237 );
and \U$524 ( \656 , \158 , \245 );
and \U$525 ( \657 , \134 , \243 );
nor \U$526 ( \658 , \656 , \657 );
xnor \U$527 ( \659 , \658 , \252 );
and \U$528 ( \660 , \655 , \659 );
and \U$529 ( \661 , \166 , \141 );
and \U$530 ( \662 , \150 , \139 );
nor \U$531 ( \663 , \661 , \662 );
xnor \U$532 ( \664 , \663 , \148 );
and \U$533 ( \665 , \659 , \664 );
and \U$534 ( \666 , \655 , \664 );
or \U$535 ( \667 , \660 , \665 , \666 );
and \U$536 ( \668 , \217 , \183 );
and \U$537 ( \669 , \189 , \180 );
nor \U$538 ( \670 , \668 , \669 );
xnor \U$539 ( \671 , \670 , \179 );
and \U$540 ( \672 , \232 , \195 );
and \U$541 ( \673 , \209 , \193 );
nor \U$542 ( \674 , \672 , \673 );
xnor \U$543 ( \675 , \674 , \202 );
and \U$544 ( \676 , \671 , \675 );
and \U$545 ( \677 , \247 , \215 );
and \U$546 ( \678 , \224 , \213 );
nor \U$547 ( \679 , \677 , \678 );
xnor \U$548 ( \680 , \679 , \222 );
and \U$549 ( \681 , \675 , \680 );
and \U$550 ( \682 , \671 , \680 );
or \U$551 ( \683 , \676 , \681 , \682 );
and \U$552 ( \684 , \667 , \683 );
and \U$553 ( \685 , \150 , \141 );
and \U$554 ( \686 , \158 , \139 );
nor \U$555 ( \687 , \685 , \686 );
xnor \U$556 ( \688 , \687 , \148 );
and \U$557 ( \689 , \683 , \688 );
and \U$558 ( \690 , \667 , \688 );
or \U$559 ( \691 , \684 , \689 , \690 );
nand \U$560 ( \692 , \166 , \154 );
xnor \U$561 ( \693 , \692 , \163 );
xor \U$562 ( \694 , \600 , \604 );
xor \U$563 ( \695 , \694 , \163 );
and \U$564 ( \696 , \693 , \695 );
xor \U$565 ( \697 , \612 , \616 );
xor \U$566 ( \698 , \697 , \621 );
and \U$567 ( \699 , \695 , \698 );
and \U$568 ( \700 , \693 , \698 );
or \U$569 ( \701 , \696 , \699 , \700 );
and \U$570 ( \702 , \691 , \701 );
xor \U$571 ( \703 , \556 , \560 );
xor \U$572 ( \704 , \703 , \565 );
and \U$573 ( \705 , \701 , \704 );
and \U$574 ( \706 , \691 , \704 );
or \U$575 ( \707 , \702 , \705 , \706 );
xor \U$576 ( \708 , \540 , \544 );
xor \U$577 ( \709 , \708 , \549 );
xor \U$578 ( \710 , \608 , \624 );
xor \U$579 ( \711 , \710 , \629 );
and \U$580 ( \712 , \709 , \711 );
and \U$581 ( \713 , \707 , \712 );
xor \U$582 ( \714 , \632 , \634 );
xor \U$583 ( \715 , \714 , \636 );
and \U$584 ( \716 , \712 , \715 );
and \U$585 ( \717 , \707 , \715 );
or \U$586 ( \718 , \713 , \716 , \717 );
and \U$587 ( \719 , \651 , \718 );
xor \U$588 ( \720 , \651 , \718 );
xor \U$589 ( \721 , \707 , \712 );
xor \U$590 ( \722 , \721 , \715 );
and \U$591 ( \723 , \240 , \215 );
and \U$592 ( \724 , \247 , \213 );
nor \U$593 ( \725 , \723 , \724 );
xnor \U$594 ( \726 , \725 , \222 );
and \U$595 ( \727 , \134 , \230 );
and \U$596 ( \728 , \143 , \228 );
nor \U$597 ( \729 , \727 , \728 );
xnor \U$598 ( \730 , \729 , \237 );
and \U$599 ( \731 , \726 , \730 );
and \U$600 ( \732 , \150 , \245 );
and \U$601 ( \733 , \158 , \243 );
nor \U$602 ( \734 , \732 , \733 );
xnor \U$603 ( \735 , \734 , \252 );
and \U$604 ( \736 , \730 , \735 );
and \U$605 ( \737 , \726 , \735 );
or \U$606 ( \738 , \731 , \736 , \737 );
and \U$607 ( \739 , \209 , \183 );
and \U$608 ( \740 , \217 , \180 );
nor \U$609 ( \741 , \739 , \740 );
xnor \U$610 ( \742 , \741 , \179 );
and \U$611 ( \743 , \224 , \195 );
and \U$612 ( \744 , \232 , \193 );
nor \U$613 ( \745 , \743 , \744 );
xnor \U$614 ( \746 , \745 , \202 );
and \U$615 ( \747 , \742 , \746 );
and \U$616 ( \748 , \746 , \148 );
and \U$617 ( \749 , \742 , \148 );
or \U$618 ( \750 , \747 , \748 , \749 );
and \U$619 ( \751 , \738 , \750 );
xor \U$620 ( \752 , \655 , \659 );
xor \U$621 ( \753 , \752 , \664 );
and \U$622 ( \754 , \750 , \753 );
and \U$623 ( \755 , \738 , \753 );
or \U$624 ( \756 , \751 , \754 , \755 );
xor \U$625 ( \757 , \667 , \683 );
xor \U$626 ( \758 , \757 , \688 );
and \U$627 ( \759 , \756 , \758 );
xor \U$628 ( \760 , \693 , \695 );
xor \U$629 ( \761 , \760 , \698 );
and \U$630 ( \762 , \758 , \761 );
and \U$631 ( \763 , \756 , \761 );
or \U$632 ( \764 , \759 , \762 , \763 );
xor \U$633 ( \765 , \691 , \701 );
xor \U$634 ( \766 , \765 , \704 );
and \U$635 ( \767 , \764 , \766 );
xor \U$636 ( \768 , \709 , \711 );
and \U$637 ( \769 , \766 , \768 );
and \U$638 ( \770 , \764 , \768 );
or \U$639 ( \771 , \767 , \769 , \770 );
and \U$640 ( \772 , \722 , \771 );
xor \U$641 ( \773 , \722 , \771 );
xor \U$642 ( \774 , \764 , \766 );
xor \U$643 ( \775 , \774 , \768 );
and \U$644 ( \776 , \232 , \183 );
and \U$645 ( \777 , \209 , \180 );
nor \U$646 ( \778 , \776 , \777 );
xnor \U$647 ( \779 , \778 , \179 );
and \U$648 ( \780 , \247 , \195 );
and \U$649 ( \781 , \224 , \193 );
nor \U$650 ( \782 , \780 , \781 );
xnor \U$651 ( \783 , \782 , \202 );
and \U$652 ( \784 , \779 , \783 );
and \U$653 ( \785 , \143 , \215 );
and \U$654 ( \786 , \240 , \213 );
nor \U$655 ( \787 , \785 , \786 );
xnor \U$656 ( \788 , \787 , \222 );
and \U$657 ( \789 , \783 , \788 );
and \U$658 ( \790 , \779 , \788 );
or \U$659 ( \791 , \784 , \789 , \790 );
nand \U$660 ( \792 , \166 , \139 );
xnor \U$661 ( \793 , \792 , \148 );
and \U$662 ( \794 , \791 , \793 );
xor \U$663 ( \795 , \726 , \730 );
xor \U$664 ( \796 , \795 , \735 );
and \U$665 ( \797 , \793 , \796 );
and \U$666 ( \798 , \791 , \796 );
or \U$667 ( \799 , \794 , \797 , \798 );
xor \U$668 ( \800 , \671 , \675 );
xor \U$669 ( \801 , \800 , \680 );
and \U$670 ( \802 , \799 , \801 );
xor \U$671 ( \803 , \738 , \750 );
xor \U$672 ( \804 , \803 , \753 );
and \U$673 ( \805 , \801 , \804 );
and \U$674 ( \806 , \799 , \804 );
or \U$675 ( \807 , \802 , \805 , \806 );
xor \U$676 ( \808 , \756 , \758 );
xor \U$677 ( \809 , \808 , \761 );
and \U$678 ( \810 , \807 , \809 );
and \U$679 ( \811 , \775 , \810 );
xor \U$680 ( \812 , \775 , \810 );
xor \U$681 ( \813 , \807 , \809 );
and \U$682 ( \814 , \134 , \215 );
and \U$683 ( \815 , \143 , \213 );
nor \U$684 ( \816 , \814 , \815 );
xnor \U$685 ( \817 , \816 , \222 );
and \U$686 ( \818 , \150 , \230 );
and \U$687 ( \819 , \158 , \228 );
nor \U$688 ( \820 , \818 , \819 );
xnor \U$689 ( \821 , \820 , \237 );
and \U$690 ( \822 , \817 , \821 );
nand \U$691 ( \823 , \166 , \243 );
xnor \U$692 ( \824 , \823 , \252 );
and \U$693 ( \825 , \821 , \824 );
and \U$694 ( \826 , \817 , \824 );
or \U$695 ( \827 , \822 , \825 , \826 );
and \U$696 ( \828 , \224 , \183 );
and \U$697 ( \829 , \232 , \180 );
nor \U$698 ( \830 , \828 , \829 );
xnor \U$699 ( \831 , \830 , \179 );
and \U$700 ( \832 , \240 , \195 );
and \U$701 ( \833 , \247 , \193 );
nor \U$702 ( \834 , \832 , \833 );
xnor \U$703 ( \835 , \834 , \202 );
and \U$704 ( \836 , \831 , \835 );
and \U$705 ( \837 , \835 , \252 );
and \U$706 ( \838 , \831 , \252 );
or \U$707 ( \839 , \836 , \837 , \838 );
and \U$708 ( \840 , \827 , \839 );
and \U$709 ( \841 , \158 , \230 );
and \U$710 ( \842 , \134 , \228 );
nor \U$711 ( \843 , \841 , \842 );
xnor \U$712 ( \844 , \843 , \237 );
and \U$713 ( \845 , \839 , \844 );
and \U$714 ( \846 , \827 , \844 );
or \U$715 ( \847 , \840 , \845 , \846 );
and \U$716 ( \848 , \166 , \245 );
and \U$717 ( \849 , \150 , \243 );
nor \U$718 ( \850 , \848 , \849 );
xnor \U$719 ( \851 , \850 , \252 );
xor \U$720 ( \852 , \779 , \783 );
xor \U$721 ( \853 , \852 , \788 );
and \U$722 ( \854 , \851 , \853 );
and \U$723 ( \855 , \847 , \854 );
xor \U$724 ( \856 , \742 , \746 );
xor \U$725 ( \857 , \856 , \148 );
and \U$726 ( \858 , \854 , \857 );
and \U$727 ( \859 , \847 , \857 );
or \U$728 ( \860 , \855 , \858 , \859 );
xor \U$729 ( \861 , \799 , \801 );
xor \U$730 ( \862 , \861 , \804 );
and \U$731 ( \863 , \860 , \862 );
and \U$732 ( \864 , \813 , \863 );
xor \U$733 ( \865 , \813 , \863 );
xor \U$734 ( \866 , \860 , \862 );
xor \U$735 ( \867 , \791 , \793 );
xor \U$736 ( \868 , \867 , \796 );
xor \U$737 ( \869 , \847 , \854 );
xor \U$738 ( \870 , \869 , \857 );
and \U$739 ( \871 , \868 , \870 );
and \U$740 ( \872 , \866 , \871 );
xor \U$741 ( \873 , \866 , \871 );
xor \U$742 ( \874 , \868 , \870 );
and \U$743 ( \875 , \247 , \183 );
and \U$744 ( \876 , \224 , \180 );
nor \U$745 ( \877 , \875 , \876 );
xnor \U$746 ( \878 , \877 , \179 );
and \U$747 ( \879 , \143 , \195 );
and \U$748 ( \880 , \240 , \193 );
nor \U$749 ( \881 , \879 , \880 );
xnor \U$750 ( \882 , \881 , \202 );
and \U$751 ( \883 , \878 , \882 );
and \U$752 ( \884 , \158 , \215 );
and \U$753 ( \885 , \134 , \213 );
nor \U$754 ( \886 , \884 , \885 );
xnor \U$755 ( \887 , \886 , \222 );
and \U$756 ( \888 , \882 , \887 );
and \U$757 ( \889 , \878 , \887 );
or \U$758 ( \890 , \883 , \888 , \889 );
xor \U$759 ( \891 , \817 , \821 );
xor \U$760 ( \892 , \891 , \824 );
and \U$761 ( \893 , \890 , \892 );
xor \U$762 ( \894 , \831 , \835 );
xor \U$763 ( \895 , \894 , \252 );
and \U$764 ( \896 , \892 , \895 );
and \U$765 ( \897 , \890 , \895 );
or \U$766 ( \898 , \893 , \896 , \897 );
xor \U$767 ( \899 , \827 , \839 );
xor \U$768 ( \900 , \899 , \844 );
and \U$769 ( \901 , \898 , \900 );
xor \U$770 ( \902 , \851 , \853 );
and \U$771 ( \903 , \900 , \902 );
and \U$772 ( \904 , \898 , \902 );
or \U$773 ( \905 , \901 , \903 , \904 );
and \U$774 ( \906 , \874 , \905 );
xor \U$775 ( \907 , \874 , \905 );
xor \U$776 ( \908 , \898 , \900 );
xor \U$777 ( \909 , \908 , \902 );
and \U$778 ( \910 , \240 , \183 );
and \U$779 ( \911 , \247 , \180 );
nor \U$780 ( \912 , \910 , \911 );
xnor \U$781 ( \913 , \912 , \179 );
and \U$782 ( \914 , \134 , \195 );
and \U$783 ( \915 , \143 , \193 );
nor \U$784 ( \916 , \914 , \915 );
xnor \U$785 ( \917 , \916 , \202 );
and \U$786 ( \918 , \913 , \917 );
and \U$787 ( \919 , \917 , \237 );
and \U$788 ( \920 , \913 , \237 );
or \U$789 ( \921 , \918 , \919 , \920 );
and \U$790 ( \922 , \150 , \215 );
and \U$791 ( \923 , \158 , \213 );
nor \U$792 ( \924 , \922 , \923 );
xnor \U$793 ( \925 , \924 , \222 );
nand \U$794 ( \926 , \166 , \228 );
xnor \U$795 ( \927 , \926 , \237 );
and \U$796 ( \928 , \925 , \927 );
and \U$797 ( \929 , \921 , \928 );
and \U$798 ( \930 , \166 , \230 );
and \U$799 ( \931 , \150 , \228 );
nor \U$800 ( \932 , \930 , \931 );
xnor \U$801 ( \933 , \932 , \237 );
and \U$802 ( \934 , \928 , \933 );
and \U$803 ( \935 , \921 , \933 );
or \U$804 ( \936 , \929 , \934 , \935 );
xor \U$805 ( \937 , \890 , \892 );
xor \U$806 ( \938 , \937 , \895 );
and \U$807 ( \939 , \936 , \938 );
and \U$808 ( \940 , \909 , \939 );
xor \U$809 ( \941 , \909 , \939 );
xor \U$810 ( \942 , \936 , \938 );
xor \U$811 ( \943 , \878 , \882 );
xor \U$812 ( \944 , \943 , \887 );
xor \U$813 ( \945 , \921 , \928 );
xor \U$814 ( \946 , \945 , \933 );
and \U$815 ( \947 , \944 , \946 );
and \U$816 ( \948 , \942 , \947 );
xor \U$817 ( \949 , \942 , \947 );
xor \U$818 ( \950 , \944 , \946 );
and \U$819 ( \951 , \143 , \183 );
and \U$820 ( \952 , \240 , \180 );
nor \U$821 ( \953 , \951 , \952 );
xnor \U$822 ( \954 , \953 , \179 );
and \U$823 ( \955 , \158 , \195 );
and \U$824 ( \956 , \134 , \193 );
nor \U$825 ( \957 , \955 , \956 );
xnor \U$826 ( \958 , \957 , \202 );
and \U$827 ( \959 , \954 , \958 );
and \U$828 ( \960 , \166 , \215 );
and \U$829 ( \961 , \150 , \213 );
nor \U$830 ( \962 , \960 , \961 );
xnor \U$831 ( \963 , \962 , \222 );
and \U$832 ( \964 , \958 , \963 );
and \U$833 ( \965 , \954 , \963 );
or \U$834 ( \966 , \959 , \964 , \965 );
xor \U$835 ( \967 , \913 , \917 );
xor \U$836 ( \968 , \967 , \237 );
and \U$837 ( \969 , \966 , \968 );
xor \U$838 ( \970 , \925 , \927 );
and \U$839 ( \971 , \968 , \970 );
and \U$840 ( \972 , \966 , \970 );
or \U$841 ( \973 , \969 , \971 , \972 );
and \U$842 ( \974 , \950 , \973 );
xor \U$843 ( \975 , \950 , \973 );
xor \U$844 ( \976 , \966 , \968 );
xor \U$845 ( \977 , \976 , \970 );
and \U$846 ( \978 , \134 , \183 );
and \U$847 ( \979 , \143 , \180 );
nor \U$848 ( \980 , \978 , \979 );
xnor \U$849 ( \981 , \980 , \179 );
and \U$850 ( \982 , \150 , \195 );
and \U$851 ( \983 , \158 , \193 );
nor \U$852 ( \984 , \982 , \983 );
xnor \U$853 ( \985 , \984 , \202 );
and \U$854 ( \986 , \981 , \985 );
and \U$855 ( \987 , \985 , \222 );
and \U$856 ( \988 , \981 , \222 );
or \U$857 ( \989 , \986 , \987 , \988 );
xor \U$858 ( \990 , \954 , \958 );
xor \U$859 ( \991 , \990 , \963 );
and \U$860 ( \992 , \989 , \991 );
and \U$861 ( \993 , \977 , \992 );
xor \U$862 ( \994 , \977 , \992 );
xor \U$863 ( \995 , \989 , \991 );
nand \U$864 ( \996 , \166 , \213 );
xnor \U$865 ( \997 , \996 , \222 );
xor \U$866 ( \998 , \981 , \985 );
xor \U$867 ( \999 , \998 , \222 );
and \U$868 ( \1000 , \997 , \999 );
and \U$869 ( \1001 , \995 , \1000 );
xor \U$870 ( \1002 , \995 , \1000 );
xor \U$871 ( \1003 , \997 , \999 );
and \U$872 ( \1004 , \158 , \183 );
and \U$873 ( \1005 , \134 , \180 );
nor \U$874 ( \1006 , \1004 , \1005 );
xnor \U$875 ( \1007 , \1006 , \179 );
and \U$876 ( \1008 , \166 , \195 );
and \U$877 ( \1009 , \150 , \193 );
nor \U$878 ( \1010 , \1008 , \1009 );
xnor \U$879 ( \1011 , \1010 , \202 );
and \U$880 ( \1012 , \1007 , \1011 );
and \U$881 ( \1013 , \1003 , \1012 );
xor \U$882 ( \1014 , \1003 , \1012 );
xor \U$883 ( \1015 , \1007 , \1011 );
and \U$884 ( \1016 , \150 , \183 );
and \U$885 ( \1017 , \158 , \180 );
nor \U$886 ( \1018 , \1016 , \1017 );
xnor \U$887 ( \1019 , \1018 , \179 );
and \U$888 ( \1020 , \1019 , \202 );
and \U$889 ( \1021 , \1015 , \1020 );
xor \U$890 ( \1022 , \1015 , \1020 );
nand \U$891 ( \1023 , \166 , \193 );
xnor \U$892 ( \1024 , \1023 , \202 );
xor \U$893 ( \1025 , \1019 , \202 );
and \U$894 ( \1026 , \1024 , \1025 );
xor \U$895 ( \1027 , \1024 , \1025 );
and \U$896 ( \1028 , \166 , \183 );
and \U$897 ( \1029 , \150 , \180 );
nor \U$898 ( \1030 , \1028 , \1029 );
xnor \U$899 ( \1031 , \1030 , \179 );
nand \U$900 ( \1032 , \166 , \180 );
xnor \U$901 ( \1033 , \1032 , \179 );
and \U$902 ( \1034 , \1033 , \179 );
and \U$903 ( \1035 , \1031 , \1034 );
and \U$904 ( \1036 , \1027 , \1035 );
or \U$905 ( \1037 , \1026 , \1036 );
and \U$906 ( \1038 , \1022 , \1037 );
or \U$907 ( \1039 , \1021 , \1038 );
and \U$908 ( \1040 , \1014 , \1039 );
or \U$909 ( \1041 , \1013 , \1040 );
and \U$910 ( \1042 , \1002 , \1041 );
or \U$911 ( \1043 , \1001 , \1042 );
and \U$912 ( \1044 , \994 , \1043 );
or \U$913 ( \1045 , \993 , \1044 );
and \U$914 ( \1046 , \975 , \1045 );
or \U$915 ( \1047 , \974 , \1046 );
and \U$916 ( \1048 , \949 , \1047 );
or \U$917 ( \1049 , \948 , \1048 );
and \U$918 ( \1050 , \941 , \1049 );
or \U$919 ( \1051 , \940 , \1050 );
and \U$920 ( \1052 , \907 , \1051 );
or \U$921 ( \1053 , \906 , \1052 );
and \U$922 ( \1054 , \873 , \1053 );
or \U$923 ( \1055 , \872 , \1054 );
and \U$924 ( \1056 , \865 , \1055 );
or \U$925 ( \1057 , \864 , \1056 );
and \U$926 ( \1058 , \812 , \1057 );
or \U$927 ( \1059 , \811 , \1058 );
and \U$928 ( \1060 , \773 , \1059 );
or \U$929 ( \1061 , \772 , \1060 );
and \U$930 ( \1062 , \720 , \1061 );
or \U$931 ( \1063 , \719 , \1062 );
and \U$932 ( \1064 , \649 , \1063 );
or \U$933 ( \1065 , \648 , \1064 );
and \U$934 ( \1066 , \594 , \1065 );
or \U$935 ( \1067 , \593 , \1066 );
xor \U$936 ( \1068 , \535 , \1067 );
buf \U$937 ( \1069 , \1068 );
buf \U$938 ( \1070 , \1069 );
and \U$939 ( \1071 , \447 , \471 );
and \U$940 ( \1072 , \471 , \527 );
and \U$941 ( \1073 , \447 , \527 );
or \U$942 ( \1074 , \1071 , \1072 , \1073 );
and \U$943 ( \1075 , \451 , \455 );
and \U$944 ( \1076 , \455 , \470 );
and \U$945 ( \1077 , \451 , \470 );
or \U$946 ( \1078 , \1075 , \1076 , \1077 );
and \U$947 ( \1079 , \488 , \502 );
and \U$948 ( \1080 , \502 , \526 );
and \U$949 ( \1081 , \488 , \526 );
or \U$950 ( \1082 , \1079 , \1080 , \1081 );
xor \U$951 ( \1083 , \1078 , \1082 );
xor \U$952 ( \1084 , \483 , \484 );
not \U$953 ( \1085 , \508 );
and \U$954 ( \1086 , \1084 , \1085 );
and \U$955 ( \1087 , \166 , \1086 );
and \U$956 ( \1088 , \150 , \508 );
nor \U$957 ( \1089 , \1087 , \1088 );
xnor \U$958 ( \1090 , \1089 , \487 );
and \U$959 ( \1091 , \247 , \156 );
and \U$960 ( \1092 , \224 , \154 );
nor \U$961 ( \1093 , \1091 , \1092 );
xnor \U$962 ( \1094 , \1093 , \163 );
and \U$963 ( \1095 , \143 , \296 );
and \U$964 ( \1096 , \240 , \168 );
nor \U$965 ( \1097 , \1095 , \1096 );
xnor \U$966 ( \1098 , \1097 , \173 );
xor \U$967 ( \1099 , \1094 , \1098 );
and \U$968 ( \1100 , \158 , \438 );
and \U$969 ( \1101 , \134 , \336 );
nor \U$970 ( \1102 , \1100 , \1101 );
xnor \U$971 ( \1103 , \1102 , \320 );
xor \U$972 ( \1104 , \1099 , \1103 );
xor \U$973 ( \1105 , \1090 , \1104 );
and \U$974 ( \1106 , \197 , \230 );
and \U$975 ( \1107 , \178 , \228 );
nor \U$976 ( \1108 , \1106 , \1107 );
xnor \U$977 ( \1109 , \1108 , \237 );
and \U$978 ( \1110 , \217 , \245 );
and \U$979 ( \1111 , \189 , \243 );
nor \U$980 ( \1112 , \1110 , \1111 );
xnor \U$981 ( \1113 , \1112 , \252 );
xor \U$982 ( \1114 , \1109 , \1113 );
and \U$983 ( \1115 , \232 , \141 );
and \U$984 ( \1116 , \209 , \139 );
nor \U$985 ( \1117 , \1115 , \1116 );
xnor \U$986 ( \1118 , \1117 , \148 );
xor \U$987 ( \1119 , \1114 , \1118 );
xor \U$988 ( \1120 , \1105 , \1119 );
xor \U$989 ( \1121 , \1083 , \1120 );
xor \U$990 ( \1122 , \1074 , \1121 );
and \U$991 ( \1123 , \477 , \481 );
and \U$992 ( \1124 , \481 , \487 );
and \U$993 ( \1125 , \477 , \487 );
or \U$994 ( \1126 , \1123 , \1124 , \1125 );
and \U$995 ( \1127 , \515 , \519 );
and \U$996 ( \1128 , \519 , \524 );
and \U$997 ( \1129 , \515 , \524 );
or \U$998 ( \1130 , \1127 , \1128 , \1129 );
xor \U$999 ( \1131 , \1126 , \1130 );
and \U$1000 ( \1132 , \460 , \464 );
and \U$1001 ( \1133 , \464 , \469 );
and \U$1002 ( \1134 , \460 , \469 );
or \U$1003 ( \1135 , \1132 , \1133 , \1134 );
xor \U$1004 ( \1136 , \1131 , \1135 );
and \U$1005 ( \1137 , \492 , \496 );
and \U$1006 ( \1138 , \496 , \501 );
and \U$1007 ( \1139 , \492 , \501 );
or \U$1008 ( \1140 , \1137 , \1138 , \1139 );
and \U$1009 ( \1141 , \507 , \510 );
and \U$1010 ( \1142 , \510 , \525 );
and \U$1011 ( \1143 , \507 , \525 );
or \U$1012 ( \1144 , \1141 , \1142 , \1143 );
xor \U$1013 ( \1145 , \1140 , \1144 );
and \U$1014 ( \1146 , \474 , \183 );
buf \U$1015 ( \1147 , RIb55dd20_109);
and \U$1016 ( \1148 , \1147 , \180 );
nor \U$1017 ( \1149 , \1146 , \1148 );
xnor \U$1018 ( \1150 , \1149 , \179 );
and \U$1019 ( \1151 , \307 , \195 );
and \U$1020 ( \1152 , \412 , \193 );
nor \U$1021 ( \1153 , \1151 , \1152 );
xnor \U$1022 ( \1154 , \1153 , \202 );
xor \U$1023 ( \1155 , \1150 , \1154 );
and \U$1024 ( \1156 , \185 , \215 );
and \U$1025 ( \1157 , \261 , \213 );
nor \U$1026 ( \1158 , \1156 , \1157 );
xnor \U$1027 ( \1159 , \1158 , \222 );
xor \U$1028 ( \1160 , \1155 , \1159 );
xor \U$1029 ( \1161 , \1145 , \1160 );
xor \U$1030 ( \1162 , \1136 , \1161 );
xor \U$1031 ( \1163 , \1122 , \1162 );
and \U$1032 ( \1164 , \387 , \528 );
xor \U$1033 ( \1165 , \1163 , \1164 );
and \U$1034 ( \1166 , \529 , \534 );
and \U$1035 ( \1167 , \535 , \1067 );
or \U$1036 ( \1168 , \1166 , \1167 );
xor \U$1037 ( \1169 , \1165 , \1168 );
buf \U$1038 ( \1170 , \1169 );
buf \U$1039 ( \1171 , \1170 );
and \U$1040 ( \1172 , \1078 , \1082 );
and \U$1041 ( \1173 , \1082 , \1120 );
and \U$1042 ( \1174 , \1078 , \1120 );
or \U$1043 ( \1175 , \1172 , \1173 , \1174 );
and \U$1044 ( \1176 , \1136 , \1161 );
xor \U$1045 ( \1177 , \1175 , \1176 );
and \U$1046 ( \1178 , \1140 , \1144 );
and \U$1047 ( \1179 , \1144 , \1160 );
and \U$1048 ( \1180 , \1140 , \1160 );
or \U$1049 ( \1181 , \1178 , \1179 , \1180 );
and \U$1050 ( \1182 , \1126 , \1130 );
and \U$1051 ( \1183 , \1130 , \1135 );
and \U$1052 ( \1184 , \1126 , \1135 );
or \U$1053 ( \1185 , \1182 , \1183 , \1184 );
and \U$1054 ( \1186 , \1090 , \1104 );
and \U$1055 ( \1187 , \1104 , \1119 );
and \U$1056 ( \1188 , \1090 , \1119 );
or \U$1057 ( \1189 , \1186 , \1187 , \1188 );
xor \U$1058 ( \1190 , \1185 , \1189 );
and \U$1059 ( \1191 , \1147 , \183 );
buf \U$1060 ( \1192 , RIb55dd98_108);
and \U$1061 ( \1193 , \1192 , \180 );
nor \U$1062 ( \1194 , \1191 , \1193 );
xnor \U$1063 ( \1195 , \1194 , \179 );
and \U$1064 ( \1196 , \412 , \195 );
and \U$1065 ( \1197 , \474 , \193 );
nor \U$1066 ( \1198 , \1196 , \1197 );
xnor \U$1067 ( \1199 , \1198 , \202 );
xor \U$1068 ( \1200 , \1195 , \1199 );
buf \U$1069 ( \1201 , RIb55fc10_43);
buf \U$1070 ( \1202 , RIb55fb98_44);
and \U$1071 ( \1203 , \1202 , \483 );
not \U$1072 ( \1204 , \1203 );
and \U$1073 ( \1205 , \1201 , \1204 );
xor \U$1074 ( \1206 , \1200 , \1205 );
xor \U$1075 ( \1207 , \1190 , \1206 );
xor \U$1076 ( \1208 , \1181 , \1207 );
and \U$1077 ( \1209 , \1094 , \1098 );
and \U$1078 ( \1210 , \1098 , \1103 );
and \U$1079 ( \1211 , \1094 , \1103 );
or \U$1080 ( \1212 , \1209 , \1210 , \1211 );
and \U$1081 ( \1213 , \1150 , \1154 );
and \U$1082 ( \1214 , \1154 , \1159 );
and \U$1083 ( \1215 , \1150 , \1159 );
or \U$1084 ( \1216 , \1213 , \1214 , \1215 );
xor \U$1085 ( \1217 , \1212 , \1216 );
and \U$1086 ( \1218 , \1109 , \1113 );
and \U$1087 ( \1219 , \1113 , \1118 );
and \U$1088 ( \1220 , \1109 , \1118 );
or \U$1089 ( \1221 , \1218 , \1219 , \1220 );
xor \U$1090 ( \1222 , \1217 , \1221 );
and \U$1091 ( \1223 , \261 , \215 );
and \U$1092 ( \1224 , \307 , \213 );
nor \U$1093 ( \1225 , \1223 , \1224 );
xnor \U$1094 ( \1226 , \1225 , \222 );
and \U$1095 ( \1227 , \178 , \230 );
and \U$1096 ( \1228 , \185 , \228 );
nor \U$1097 ( \1229 , \1227 , \1228 );
xnor \U$1098 ( \1230 , \1229 , \237 );
xor \U$1099 ( \1231 , \1226 , \1230 );
and \U$1100 ( \1232 , \189 , \245 );
and \U$1101 ( \1233 , \197 , \243 );
nor \U$1102 ( \1234 , \1232 , \1233 );
xnor \U$1103 ( \1235 , \1234 , \252 );
xor \U$1104 ( \1236 , \1231 , \1235 );
and \U$1105 ( \1237 , \134 , \438 );
and \U$1106 ( \1238 , \143 , \336 );
nor \U$1107 ( \1239 , \1237 , \1238 );
xnor \U$1108 ( \1240 , \1239 , \320 );
and \U$1109 ( \1241 , \150 , \1086 );
and \U$1110 ( \1242 , \158 , \508 );
nor \U$1111 ( \1243 , \1241 , \1242 );
xnor \U$1112 ( \1244 , \1243 , \487 );
xor \U$1113 ( \1245 , \1240 , \1244 );
xor \U$1114 ( \1246 , \1202 , \483 );
nand \U$1115 ( \1247 , \166 , \1246 );
xnor \U$1116 ( \1248 , \1247 , \1205 );
xor \U$1117 ( \1249 , \1245 , \1248 );
xor \U$1118 ( \1250 , \1236 , \1249 );
and \U$1119 ( \1251 , \209 , \141 );
and \U$1120 ( \1252 , \217 , \139 );
nor \U$1121 ( \1253 , \1251 , \1252 );
xnor \U$1122 ( \1254 , \1253 , \148 );
and \U$1123 ( \1255 , \224 , \156 );
and \U$1124 ( \1256 , \232 , \154 );
nor \U$1125 ( \1257 , \1255 , \1256 );
xnor \U$1126 ( \1258 , \1257 , \163 );
xor \U$1127 ( \1259 , \1254 , \1258 );
and \U$1128 ( \1260 , \240 , \296 );
and \U$1129 ( \1261 , \247 , \168 );
nor \U$1130 ( \1262 , \1260 , \1261 );
xnor \U$1131 ( \1263 , \1262 , \173 );
xor \U$1132 ( \1264 , \1259 , \1263 );
xor \U$1133 ( \1265 , \1250 , \1264 );
xor \U$1134 ( \1266 , \1222 , \1265 );
xor \U$1135 ( \1267 , \1208 , \1266 );
xor \U$1136 ( \1268 , \1177 , \1267 );
and \U$1137 ( \1269 , \1074 , \1121 );
and \U$1138 ( \1270 , \1121 , \1162 );
and \U$1139 ( \1271 , \1074 , \1162 );
or \U$1140 ( \1272 , \1269 , \1270 , \1271 );
xor \U$1141 ( \1273 , \1268 , \1272 );
and \U$1142 ( \1274 , \1163 , \1164 );
and \U$1143 ( \1275 , \1165 , \1168 );
or \U$1144 ( \1276 , \1274 , \1275 );
xor \U$1145 ( \1277 , \1273 , \1276 );
buf \U$1146 ( \1278 , \1277 );
buf \U$1147 ( \1279 , \1278 );
and \U$1148 ( \1280 , \1181 , \1207 );
and \U$1149 ( \1281 , \1207 , \1266 );
and \U$1150 ( \1282 , \1181 , \1266 );
or \U$1151 ( \1283 , \1280 , \1281 , \1282 );
and \U$1152 ( \1284 , \1185 , \1189 );
and \U$1153 ( \1285 , \1189 , \1206 );
and \U$1154 ( \1286 , \1185 , \1206 );
or \U$1155 ( \1287 , \1284 , \1285 , \1286 );
and \U$1156 ( \1288 , \1222 , \1265 );
xor \U$1157 ( \1289 , \1287 , \1288 );
and \U$1158 ( \1290 , \1240 , \1244 );
and \U$1159 ( \1291 , \1244 , \1248 );
and \U$1160 ( \1292 , \1240 , \1248 );
or \U$1161 ( \1293 , \1290 , \1291 , \1292 );
and \U$1162 ( \1294 , \158 , \1086 );
and \U$1163 ( \1295 , \134 , \508 );
nor \U$1164 ( \1296 , \1294 , \1295 );
xnor \U$1165 ( \1297 , \1296 , \487 );
xor \U$1166 ( \1298 , \1293 , \1297 );
xor \U$1167 ( \1299 , \1201 , \1202 );
not \U$1168 ( \1300 , \1246 );
and \U$1169 ( \1301 , \1299 , \1300 );
and \U$1170 ( \1302 , \166 , \1301 );
and \U$1171 ( \1303 , \150 , \1246 );
nor \U$1172 ( \1304 , \1302 , \1303 );
xnor \U$1173 ( \1305 , \1304 , \1205 );
xor \U$1174 ( \1306 , \1298 , \1305 );
xor \U$1175 ( \1307 , \1289 , \1306 );
xor \U$1176 ( \1308 , \1283 , \1307 );
and \U$1177 ( \1309 , \1195 , \1199 );
and \U$1178 ( \1310 , \1199 , \1205 );
and \U$1179 ( \1311 , \1195 , \1205 );
or \U$1180 ( \1312 , \1309 , \1310 , \1311 );
and \U$1181 ( \1313 , \1226 , \1230 );
and \U$1182 ( \1314 , \1230 , \1235 );
and \U$1183 ( \1315 , \1226 , \1235 );
or \U$1184 ( \1316 , \1313 , \1314 , \1315 );
xor \U$1185 ( \1317 , \1312 , \1316 );
and \U$1186 ( \1318 , \1254 , \1258 );
and \U$1187 ( \1319 , \1258 , \1263 );
and \U$1188 ( \1320 , \1254 , \1263 );
or \U$1189 ( \1321 , \1318 , \1319 , \1320 );
xor \U$1190 ( \1322 , \1317 , \1321 );
and \U$1191 ( \1323 , \1212 , \1216 );
and \U$1192 ( \1324 , \1216 , \1221 );
and \U$1193 ( \1325 , \1212 , \1221 );
or \U$1194 ( \1326 , \1323 , \1324 , \1325 );
and \U$1195 ( \1327 , \1236 , \1249 );
and \U$1196 ( \1328 , \1249 , \1264 );
and \U$1197 ( \1329 , \1236 , \1264 );
or \U$1198 ( \1330 , \1327 , \1328 , \1329 );
xor \U$1199 ( \1331 , \1326 , \1330 );
and \U$1200 ( \1332 , \1192 , \183 );
buf \U$1201 ( \1333 , RIb55de10_107);
and \U$1202 ( \1334 , \1333 , \180 );
nor \U$1203 ( \1335 , \1332 , \1334 );
xnor \U$1204 ( \1336 , \1335 , \179 );
and \U$1205 ( \1337 , \474 , \195 );
and \U$1206 ( \1338 , \1147 , \193 );
nor \U$1207 ( \1339 , \1337 , \1338 );
xnor \U$1208 ( \1340 , \1339 , \202 );
xor \U$1209 ( \1341 , \1336 , \1340 );
and \U$1210 ( \1342 , \307 , \215 );
and \U$1211 ( \1343 , \412 , \213 );
nor \U$1212 ( \1344 , \1342 , \1343 );
xnor \U$1213 ( \1345 , \1344 , \222 );
xor \U$1214 ( \1346 , \1341 , \1345 );
and \U$1215 ( \1347 , \232 , \156 );
and \U$1216 ( \1348 , \209 , \154 );
nor \U$1217 ( \1349 , \1347 , \1348 );
xnor \U$1218 ( \1350 , \1349 , \163 );
and \U$1219 ( \1351 , \247 , \296 );
and \U$1220 ( \1352 , \224 , \168 );
nor \U$1221 ( \1353 , \1351 , \1352 );
xnor \U$1222 ( \1354 , \1353 , \173 );
xor \U$1223 ( \1355 , \1350 , \1354 );
and \U$1224 ( \1356 , \143 , \438 );
and \U$1225 ( \1357 , \240 , \336 );
nor \U$1226 ( \1358 , \1356 , \1357 );
xnor \U$1227 ( \1359 , \1358 , \320 );
xor \U$1228 ( \1360 , \1355 , \1359 );
xor \U$1229 ( \1361 , \1346 , \1360 );
and \U$1230 ( \1362 , \185 , \230 );
and \U$1231 ( \1363 , \261 , \228 );
nor \U$1232 ( \1364 , \1362 , \1363 );
xnor \U$1233 ( \1365 , \1364 , \237 );
and \U$1234 ( \1366 , \197 , \245 );
and \U$1235 ( \1367 , \178 , \243 );
nor \U$1236 ( \1368 , \1366 , \1367 );
xnor \U$1237 ( \1369 , \1368 , \252 );
xor \U$1238 ( \1370 , \1365 , \1369 );
and \U$1239 ( \1371 , \217 , \141 );
and \U$1240 ( \1372 , \189 , \139 );
nor \U$1241 ( \1373 , \1371 , \1372 );
xnor \U$1242 ( \1374 , \1373 , \148 );
xor \U$1243 ( \1375 , \1370 , \1374 );
xor \U$1244 ( \1376 , \1361 , \1375 );
xor \U$1245 ( \1377 , \1331 , \1376 );
xor \U$1246 ( \1378 , \1322 , \1377 );
xor \U$1247 ( \1379 , \1308 , \1378 );
and \U$1248 ( \1380 , \1175 , \1176 );
and \U$1249 ( \1381 , \1176 , \1267 );
and \U$1250 ( \1382 , \1175 , \1267 );
or \U$1251 ( \1383 , \1380 , \1381 , \1382 );
xor \U$1252 ( \1384 , \1379 , \1383 );
and \U$1253 ( \1385 , \1268 , \1272 );
and \U$1254 ( \1386 , \1273 , \1276 );
or \U$1255 ( \1387 , \1385 , \1386 );
xor \U$1256 ( \1388 , \1384 , \1387 );
buf \U$1257 ( \1389 , \1388 );
buf \U$1258 ( \1390 , \1389 );
and \U$1259 ( \1391 , \1287 , \1288 );
and \U$1260 ( \1392 , \1288 , \1306 );
and \U$1261 ( \1393 , \1287 , \1306 );
or \U$1262 ( \1394 , \1391 , \1392 , \1393 );
and \U$1263 ( \1395 , \1322 , \1377 );
xor \U$1264 ( \1396 , \1394 , \1395 );
and \U$1265 ( \1397 , \1326 , \1330 );
and \U$1266 ( \1398 , \1330 , \1376 );
and \U$1267 ( \1399 , \1326 , \1376 );
or \U$1268 ( \1400 , \1397 , \1398 , \1399 );
and \U$1269 ( \1401 , \1293 , \1297 );
and \U$1270 ( \1402 , \1297 , \1305 );
and \U$1271 ( \1403 , \1293 , \1305 );
or \U$1272 ( \1404 , \1401 , \1402 , \1403 );
and \U$1273 ( \1405 , \1312 , \1316 );
and \U$1274 ( \1406 , \1316 , \1321 );
and \U$1275 ( \1407 , \1312 , \1321 );
or \U$1276 ( \1408 , \1405 , \1406 , \1407 );
xor \U$1277 ( \1409 , \1404 , \1408 );
and \U$1278 ( \1410 , \1346 , \1360 );
and \U$1279 ( \1411 , \1360 , \1375 );
and \U$1280 ( \1412 , \1346 , \1375 );
or \U$1281 ( \1413 , \1410 , \1411 , \1412 );
xor \U$1282 ( \1414 , \1409 , \1413 );
xor \U$1283 ( \1415 , \1400 , \1414 );
and \U$1284 ( \1416 , \1336 , \1340 );
and \U$1285 ( \1417 , \1340 , \1345 );
and \U$1286 ( \1418 , \1336 , \1345 );
or \U$1287 ( \1419 , \1416 , \1417 , \1418 );
and \U$1288 ( \1420 , \1350 , \1354 );
and \U$1289 ( \1421 , \1354 , \1359 );
and \U$1290 ( \1422 , \1350 , \1359 );
or \U$1291 ( \1423 , \1420 , \1421 , \1422 );
xor \U$1292 ( \1424 , \1419 , \1423 );
and \U$1293 ( \1425 , \1365 , \1369 );
and \U$1294 ( \1426 , \1369 , \1374 );
and \U$1295 ( \1427 , \1365 , \1374 );
or \U$1296 ( \1428 , \1425 , \1426 , \1427 );
xor \U$1297 ( \1429 , \1424 , \1428 );
buf \U$1298 ( \1430 , RIb55fc88_42);
xor \U$1299 ( \1431 , \1430 , \1201 );
nand \U$1300 ( \1432 , \166 , \1431 );
buf \U$1301 ( \1433 , RIb55fd00_41);
and \U$1302 ( \1434 , \1430 , \1201 );
not \U$1303 ( \1435 , \1434 );
and \U$1304 ( \1436 , \1433 , \1435 );
xnor \U$1305 ( \1437 , \1432 , \1436 );
and \U$1306 ( \1438 , \189 , \141 );
and \U$1307 ( \1439 , \197 , \139 );
nor \U$1308 ( \1440 , \1438 , \1439 );
xnor \U$1309 ( \1441 , \1440 , \148 );
and \U$1310 ( \1442 , \209 , \156 );
and \U$1311 ( \1443 , \217 , \154 );
nor \U$1312 ( \1444 , \1442 , \1443 );
xnor \U$1313 ( \1445 , \1444 , \163 );
xor \U$1314 ( \1446 , \1441 , \1445 );
and \U$1315 ( \1447 , \224 , \296 );
and \U$1316 ( \1448 , \232 , \168 );
nor \U$1317 ( \1449 , \1447 , \1448 );
xnor \U$1318 ( \1450 , \1449 , \173 );
xor \U$1319 ( \1451 , \1446 , \1450 );
xor \U$1320 ( \1452 , \1437 , \1451 );
and \U$1321 ( \1453 , \240 , \438 );
and \U$1322 ( \1454 , \247 , \336 );
nor \U$1323 ( \1455 , \1453 , \1454 );
xnor \U$1324 ( \1456 , \1455 , \320 );
and \U$1325 ( \1457 , \134 , \1086 );
and \U$1326 ( \1458 , \143 , \508 );
nor \U$1327 ( \1459 , \1457 , \1458 );
xnor \U$1328 ( \1460 , \1459 , \487 );
xor \U$1329 ( \1461 , \1456 , \1460 );
and \U$1330 ( \1462 , \150 , \1301 );
and \U$1331 ( \1463 , \158 , \1246 );
nor \U$1332 ( \1464 , \1462 , \1463 );
xnor \U$1333 ( \1465 , \1464 , \1205 );
xor \U$1334 ( \1466 , \1461 , \1465 );
xor \U$1335 ( \1467 , \1452 , \1466 );
xor \U$1336 ( \1468 , \1429 , \1467 );
and \U$1337 ( \1469 , \412 , \215 );
and \U$1338 ( \1470 , \474 , \213 );
nor \U$1339 ( \1471 , \1469 , \1470 );
xnor \U$1340 ( \1472 , \1471 , \222 );
and \U$1341 ( \1473 , \261 , \230 );
and \U$1342 ( \1474 , \307 , \228 );
nor \U$1343 ( \1475 , \1473 , \1474 );
xnor \U$1344 ( \1476 , \1475 , \237 );
xor \U$1345 ( \1477 , \1472 , \1476 );
and \U$1346 ( \1478 , \178 , \245 );
and \U$1347 ( \1479 , \185 , \243 );
nor \U$1348 ( \1480 , \1478 , \1479 );
xnor \U$1349 ( \1481 , \1480 , \252 );
xor \U$1350 ( \1482 , \1477 , \1481 );
and \U$1351 ( \1483 , \1333 , \183 );
buf \U$1352 ( \1484 , RIb55de88_106);
and \U$1353 ( \1485 , \1484 , \180 );
nor \U$1354 ( \1486 , \1483 , \1485 );
xnor \U$1355 ( \1487 , \1486 , \179 );
and \U$1356 ( \1488 , \1147 , \195 );
and \U$1357 ( \1489 , \1192 , \193 );
nor \U$1358 ( \1490 , \1488 , \1489 );
xnor \U$1359 ( \1491 , \1490 , \202 );
xor \U$1360 ( \1492 , \1487 , \1491 );
xor \U$1361 ( \1493 , \1492 , \1436 );
xor \U$1362 ( \1494 , \1482 , \1493 );
xor \U$1363 ( \1495 , \1468 , \1494 );
xor \U$1364 ( \1496 , \1415 , \1495 );
xor \U$1365 ( \1497 , \1396 , \1496 );
and \U$1366 ( \1498 , \1283 , \1307 );
and \U$1367 ( \1499 , \1307 , \1378 );
and \U$1368 ( \1500 , \1283 , \1378 );
or \U$1369 ( \1501 , \1498 , \1499 , \1500 );
xor \U$1370 ( \1502 , \1497 , \1501 );
and \U$1371 ( \1503 , \1379 , \1383 );
and \U$1372 ( \1504 , \1384 , \1387 );
or \U$1373 ( \1505 , \1503 , \1504 );
xor \U$1374 ( \1506 , \1502 , \1505 );
buf \U$1375 ( \1507 , \1506 );
buf \U$1376 ( \1508 , \1507 );
and \U$1377 ( \1509 , \1400 , \1414 );
and \U$1378 ( \1510 , \1414 , \1495 );
and \U$1379 ( \1511 , \1400 , \1495 );
or \U$1380 ( \1512 , \1509 , \1510 , \1511 );
and \U$1381 ( \1513 , \1419 , \1423 );
and \U$1382 ( \1514 , \1423 , \1428 );
and \U$1383 ( \1515 , \1419 , \1428 );
or \U$1384 ( \1516 , \1513 , \1514 , \1515 );
and \U$1385 ( \1517 , \1437 , \1451 );
and \U$1386 ( \1518 , \1451 , \1466 );
and \U$1387 ( \1519 , \1437 , \1466 );
or \U$1388 ( \1520 , \1517 , \1518 , \1519 );
xor \U$1389 ( \1521 , \1516 , \1520 );
and \U$1390 ( \1522 , \1482 , \1493 );
xor \U$1391 ( \1523 , \1521 , \1522 );
xor \U$1392 ( \1524 , \1512 , \1523 );
and \U$1393 ( \1525 , \1404 , \1408 );
and \U$1394 ( \1526 , \1408 , \1413 );
and \U$1395 ( \1527 , \1404 , \1413 );
or \U$1396 ( \1528 , \1525 , \1526 , \1527 );
and \U$1397 ( \1529 , \1429 , \1467 );
and \U$1398 ( \1530 , \1467 , \1494 );
and \U$1399 ( \1531 , \1429 , \1494 );
or \U$1400 ( \1532 , \1529 , \1530 , \1531 );
xor \U$1401 ( \1533 , \1528 , \1532 );
and \U$1402 ( \1534 , \1472 , \1476 );
and \U$1403 ( \1535 , \1476 , \1481 );
and \U$1404 ( \1536 , \1472 , \1481 );
or \U$1405 ( \1537 , \1534 , \1535 , \1536 );
and \U$1406 ( \1538 , \1441 , \1445 );
and \U$1407 ( \1539 , \1445 , \1450 );
and \U$1408 ( \1540 , \1441 , \1450 );
or \U$1409 ( \1541 , \1538 , \1539 , \1540 );
xor \U$1410 ( \1542 , \1537 , \1541 );
and \U$1411 ( \1543 , \1487 , \1491 );
and \U$1412 ( \1544 , \1491 , \1436 );
and \U$1413 ( \1545 , \1487 , \1436 );
or \U$1414 ( \1546 , \1543 , \1544 , \1545 );
xor \U$1415 ( \1547 , \1542 , \1546 );
and \U$1416 ( \1548 , \1456 , \1460 );
and \U$1417 ( \1549 , \1460 , \1465 );
and \U$1418 ( \1550 , \1456 , \1465 );
or \U$1419 ( \1551 , \1548 , \1549 , \1550 );
and \U$1420 ( \1552 , \217 , \156 );
and \U$1421 ( \1553 , \189 , \154 );
nor \U$1422 ( \1554 , \1552 , \1553 );
xnor \U$1423 ( \1555 , \1554 , \163 );
and \U$1424 ( \1556 , \232 , \296 );
and \U$1425 ( \1557 , \209 , \168 );
nor \U$1426 ( \1558 , \1556 , \1557 );
xnor \U$1427 ( \1559 , \1558 , \173 );
xor \U$1428 ( \1560 , \1555 , \1559 );
and \U$1429 ( \1561 , \247 , \438 );
and \U$1430 ( \1562 , \224 , \336 );
nor \U$1431 ( \1563 , \1561 , \1562 );
xnor \U$1432 ( \1564 , \1563 , \320 );
xor \U$1433 ( \1565 , \1560 , \1564 );
xor \U$1434 ( \1566 , \1551 , \1565 );
and \U$1435 ( \1567 , \143 , \1086 );
and \U$1436 ( \1568 , \240 , \508 );
nor \U$1437 ( \1569 , \1567 , \1568 );
xnor \U$1438 ( \1570 , \1569 , \487 );
and \U$1439 ( \1571 , \158 , \1301 );
and \U$1440 ( \1572 , \134 , \1246 );
nor \U$1441 ( \1573 , \1571 , \1572 );
xnor \U$1442 ( \1574 , \1573 , \1205 );
xor \U$1443 ( \1575 , \1570 , \1574 );
xor \U$1444 ( \1576 , \1433 , \1430 );
not \U$1445 ( \1577 , \1431 );
and \U$1446 ( \1578 , \1576 , \1577 );
and \U$1447 ( \1579 , \166 , \1578 );
and \U$1448 ( \1580 , \150 , \1431 );
nor \U$1449 ( \1581 , \1579 , \1580 );
xnor \U$1450 ( \1582 , \1581 , \1436 );
xor \U$1451 ( \1583 , \1575 , \1582 );
xor \U$1452 ( \1584 , \1566 , \1583 );
xor \U$1453 ( \1585 , \1547 , \1584 );
and \U$1454 ( \1586 , \307 , \230 );
and \U$1455 ( \1587 , \412 , \228 );
nor \U$1456 ( \1588 , \1586 , \1587 );
xnor \U$1457 ( \1589 , \1588 , \237 );
and \U$1458 ( \1590 , \185 , \245 );
and \U$1459 ( \1591 , \261 , \243 );
nor \U$1460 ( \1592 , \1590 , \1591 );
xnor \U$1461 ( \1593 , \1592 , \252 );
xor \U$1462 ( \1594 , \1589 , \1593 );
and \U$1463 ( \1595 , \197 , \141 );
and \U$1464 ( \1596 , \178 , \139 );
nor \U$1465 ( \1597 , \1595 , \1596 );
xnor \U$1466 ( \1598 , \1597 , \148 );
xor \U$1467 ( \1599 , \1594 , \1598 );
and \U$1468 ( \1600 , \1484 , \183 );
buf \U$1469 ( \1601 , RIb55df00_105);
and \U$1470 ( \1602 , \1601 , \180 );
nor \U$1471 ( \1603 , \1600 , \1602 );
xnor \U$1472 ( \1604 , \1603 , \179 );
and \U$1473 ( \1605 , \1192 , \195 );
and \U$1474 ( \1606 , \1333 , \193 );
nor \U$1475 ( \1607 , \1605 , \1606 );
xnor \U$1476 ( \1608 , \1607 , \202 );
xor \U$1477 ( \1609 , \1604 , \1608 );
and \U$1478 ( \1610 , \474 , \215 );
and \U$1479 ( \1611 , \1147 , \213 );
nor \U$1480 ( \1612 , \1610 , \1611 );
xnor \U$1481 ( \1613 , \1612 , \222 );
xor \U$1482 ( \1614 , \1609 , \1613 );
xor \U$1483 ( \1615 , \1599 , \1614 );
xor \U$1484 ( \1616 , \1585 , \1615 );
xor \U$1485 ( \1617 , \1533 , \1616 );
xor \U$1486 ( \1618 , \1524 , \1617 );
and \U$1487 ( \1619 , \1394 , \1395 );
and \U$1488 ( \1620 , \1395 , \1496 );
and \U$1489 ( \1621 , \1394 , \1496 );
or \U$1490 ( \1622 , \1619 , \1620 , \1621 );
xor \U$1491 ( \1623 , \1618 , \1622 );
and \U$1492 ( \1624 , \1497 , \1501 );
and \U$1493 ( \1625 , \1502 , \1505 );
or \U$1494 ( \1626 , \1624 , \1625 );
xor \U$1495 ( \1627 , \1623 , \1626 );
buf \U$1496 ( \1628 , \1627 );
buf \U$1497 ( \1629 , \1628 );
and \U$1498 ( \1630 , \1528 , \1532 );
and \U$1499 ( \1631 , \1532 , \1616 );
and \U$1500 ( \1632 , \1528 , \1616 );
or \U$1501 ( \1633 , \1630 , \1631 , \1632 );
and \U$1502 ( \1634 , \1537 , \1541 );
and \U$1503 ( \1635 , \1541 , \1546 );
and \U$1504 ( \1636 , \1537 , \1546 );
or \U$1505 ( \1637 , \1634 , \1635 , \1636 );
and \U$1506 ( \1638 , \1551 , \1565 );
and \U$1507 ( \1639 , \1565 , \1583 );
and \U$1508 ( \1640 , \1551 , \1583 );
or \U$1509 ( \1641 , \1638 , \1639 , \1640 );
xor \U$1510 ( \1642 , \1637 , \1641 );
and \U$1511 ( \1643 , \1599 , \1614 );
xor \U$1512 ( \1644 , \1642 , \1643 );
xor \U$1513 ( \1645 , \1633 , \1644 );
and \U$1514 ( \1646 , \1516 , \1520 );
and \U$1515 ( \1647 , \1520 , \1522 );
and \U$1516 ( \1648 , \1516 , \1522 );
or \U$1517 ( \1649 , \1646 , \1647 , \1648 );
and \U$1518 ( \1650 , \1547 , \1584 );
and \U$1519 ( \1651 , \1584 , \1615 );
and \U$1520 ( \1652 , \1547 , \1615 );
or \U$1521 ( \1653 , \1650 , \1651 , \1652 );
xor \U$1522 ( \1654 , \1649 , \1653 );
and \U$1523 ( \1655 , \1589 , \1593 );
and \U$1524 ( \1656 , \1593 , \1598 );
and \U$1525 ( \1657 , \1589 , \1598 );
or \U$1526 ( \1658 , \1655 , \1656 , \1657 );
and \U$1527 ( \1659 , \1555 , \1559 );
and \U$1528 ( \1660 , \1559 , \1564 );
and \U$1529 ( \1661 , \1555 , \1564 );
or \U$1530 ( \1662 , \1659 , \1660 , \1661 );
xor \U$1531 ( \1663 , \1658 , \1662 );
and \U$1532 ( \1664 , \1604 , \1608 );
and \U$1533 ( \1665 , \1608 , \1613 );
and \U$1534 ( \1666 , \1604 , \1613 );
or \U$1535 ( \1667 , \1664 , \1665 , \1666 );
xor \U$1536 ( \1668 , \1663 , \1667 );
and \U$1537 ( \1669 , \1147 , \215 );
and \U$1538 ( \1670 , \1192 , \213 );
nor \U$1539 ( \1671 , \1669 , \1670 );
xnor \U$1540 ( \1672 , \1671 , \222 );
and \U$1541 ( \1673 , \412 , \230 );
and \U$1542 ( \1674 , \474 , \228 );
nor \U$1543 ( \1675 , \1673 , \1674 );
xnor \U$1544 ( \1676 , \1675 , \237 );
xor \U$1545 ( \1677 , \1672 , \1676 );
and \U$1546 ( \1678 , \261 , \245 );
and \U$1547 ( \1679 , \307 , \243 );
nor \U$1548 ( \1680 , \1678 , \1679 );
xnor \U$1549 ( \1681 , \1680 , \252 );
xor \U$1550 ( \1682 , \1677 , \1681 );
and \U$1551 ( \1683 , \1601 , \183 );
buf \U$1552 ( \1684 , RIb55df78_104);
and \U$1553 ( \1685 , \1684 , \180 );
nor \U$1554 ( \1686 , \1683 , \1685 );
xnor \U$1555 ( \1687 , \1686 , \179 );
and \U$1556 ( \1688 , \1333 , \195 );
and \U$1557 ( \1689 , \1484 , \193 );
nor \U$1558 ( \1690 , \1688 , \1689 );
xnor \U$1559 ( \1691 , \1690 , \202 );
xor \U$1560 ( \1692 , \1687 , \1691 );
buf \U$1561 ( \1693 , RIb55fdf0_39);
buf \U$1562 ( \1694 , RIb55fd78_40);
and \U$1563 ( \1695 , \1694 , \1433 );
not \U$1564 ( \1696 , \1695 );
and \U$1565 ( \1697 , \1693 , \1696 );
xor \U$1566 ( \1698 , \1692 , \1697 );
xor \U$1567 ( \1699 , \1682 , \1698 );
and \U$1568 ( \1700 , \178 , \141 );
and \U$1569 ( \1701 , \185 , \139 );
nor \U$1570 ( \1702 , \1700 , \1701 );
xnor \U$1571 ( \1703 , \1702 , \148 );
and \U$1572 ( \1704 , \189 , \156 );
and \U$1573 ( \1705 , \197 , \154 );
nor \U$1574 ( \1706 , \1704 , \1705 );
xnor \U$1575 ( \1707 , \1706 , \163 );
xor \U$1576 ( \1708 , \1703 , \1707 );
and \U$1577 ( \1709 , \209 , \296 );
and \U$1578 ( \1710 , \217 , \168 );
nor \U$1579 ( \1711 , \1709 , \1710 );
xnor \U$1580 ( \1712 , \1711 , \173 );
xor \U$1581 ( \1713 , \1708 , \1712 );
xor \U$1582 ( \1714 , \1699 , \1713 );
xor \U$1583 ( \1715 , \1668 , \1714 );
and \U$1584 ( \1716 , \1570 , \1574 );
and \U$1585 ( \1717 , \1574 , \1582 );
and \U$1586 ( \1718 , \1570 , \1582 );
or \U$1587 ( \1719 , \1716 , \1717 , \1718 );
and \U$1588 ( \1720 , \224 , \438 );
and \U$1589 ( \1721 , \232 , \336 );
nor \U$1590 ( \1722 , \1720 , \1721 );
xnor \U$1591 ( \1723 , \1722 , \320 );
and \U$1592 ( \1724 , \240 , \1086 );
and \U$1593 ( \1725 , \247 , \508 );
nor \U$1594 ( \1726 , \1724 , \1725 );
xnor \U$1595 ( \1727 , \1726 , \487 );
xor \U$1596 ( \1728 , \1723 , \1727 );
and \U$1597 ( \1729 , \134 , \1301 );
and \U$1598 ( \1730 , \143 , \1246 );
nor \U$1599 ( \1731 , \1729 , \1730 );
xnor \U$1600 ( \1732 , \1731 , \1205 );
xor \U$1601 ( \1733 , \1728 , \1732 );
xor \U$1602 ( \1734 , \1719 , \1733 );
and \U$1603 ( \1735 , \150 , \1578 );
and \U$1604 ( \1736 , \158 , \1431 );
nor \U$1605 ( \1737 , \1735 , \1736 );
xnor \U$1606 ( \1738 , \1737 , \1436 );
xor \U$1607 ( \1739 , \1694 , \1433 );
nand \U$1608 ( \1740 , \166 , \1739 );
xnor \U$1609 ( \1741 , \1740 , \1697 );
xor \U$1610 ( \1742 , \1738 , \1741 );
xor \U$1611 ( \1743 , \1734 , \1742 );
xor \U$1612 ( \1744 , \1715 , \1743 );
xor \U$1613 ( \1745 , \1654 , \1744 );
xor \U$1614 ( \1746 , \1645 , \1745 );
and \U$1615 ( \1747 , \1512 , \1523 );
and \U$1616 ( \1748 , \1523 , \1617 );
and \U$1617 ( \1749 , \1512 , \1617 );
or \U$1618 ( \1750 , \1747 , \1748 , \1749 );
xor \U$1619 ( \1751 , \1746 , \1750 );
and \U$1620 ( \1752 , \1618 , \1622 );
and \U$1621 ( \1753 , \1623 , \1626 );
or \U$1622 ( \1754 , \1752 , \1753 );
xor \U$1623 ( \1755 , \1751 , \1754 );
buf \U$1624 ( \1756 , \1755 );
buf \U$1625 ( \1757 , \1756 );
and \U$1626 ( \1758 , \1649 , \1653 );
and \U$1627 ( \1759 , \1653 , \1744 );
and \U$1628 ( \1760 , \1649 , \1744 );
or \U$1629 ( \1761 , \1758 , \1759 , \1760 );
and \U$1630 ( \1762 , \1637 , \1641 );
and \U$1631 ( \1763 , \1641 , \1643 );
and \U$1632 ( \1764 , \1637 , \1643 );
or \U$1633 ( \1765 , \1762 , \1763 , \1764 );
and \U$1634 ( \1766 , \1668 , \1714 );
and \U$1635 ( \1767 , \1714 , \1743 );
and \U$1636 ( \1768 , \1668 , \1743 );
or \U$1637 ( \1769 , \1766 , \1767 , \1768 );
xor \U$1638 ( \1770 , \1765 , \1769 );
and \U$1639 ( \1771 , \1672 , \1676 );
and \U$1640 ( \1772 , \1676 , \1681 );
and \U$1641 ( \1773 , \1672 , \1681 );
or \U$1642 ( \1774 , \1771 , \1772 , \1773 );
and \U$1643 ( \1775 , \1687 , \1691 );
and \U$1644 ( \1776 , \1691 , \1697 );
and \U$1645 ( \1777 , \1687 , \1697 );
or \U$1646 ( \1778 , \1775 , \1776 , \1777 );
xor \U$1647 ( \1779 , \1774 , \1778 );
and \U$1648 ( \1780 , \1703 , \1707 );
and \U$1649 ( \1781 , \1707 , \1712 );
and \U$1650 ( \1782 , \1703 , \1712 );
or \U$1651 ( \1783 , \1780 , \1781 , \1782 );
xor \U$1652 ( \1784 , \1779 , \1783 );
xor \U$1653 ( \1785 , \1770 , \1784 );
xor \U$1654 ( \1786 , \1761 , \1785 );
and \U$1655 ( \1787 , \1658 , \1662 );
and \U$1656 ( \1788 , \1662 , \1667 );
and \U$1657 ( \1789 , \1658 , \1667 );
or \U$1658 ( \1790 , \1787 , \1788 , \1789 );
and \U$1659 ( \1791 , \1682 , \1698 );
and \U$1660 ( \1792 , \1698 , \1713 );
and \U$1661 ( \1793 , \1682 , \1713 );
or \U$1662 ( \1794 , \1791 , \1792 , \1793 );
xor \U$1663 ( \1795 , \1790 , \1794 );
and \U$1664 ( \1796 , \1719 , \1733 );
and \U$1665 ( \1797 , \1733 , \1742 );
and \U$1666 ( \1798 , \1719 , \1742 );
or \U$1667 ( \1799 , \1796 , \1797 , \1798 );
xor \U$1668 ( \1800 , \1795 , \1799 );
and \U$1669 ( \1801 , \1684 , \183 );
buf \U$1670 ( \1802 , RIb55dff0_103);
and \U$1671 ( \1803 , \1802 , \180 );
nor \U$1672 ( \1804 , \1801 , \1803 );
xnor \U$1673 ( \1805 , \1804 , \179 );
and \U$1674 ( \1806 , \1484 , \195 );
and \U$1675 ( \1807 , \1601 , \193 );
nor \U$1676 ( \1808 , \1806 , \1807 );
xnor \U$1677 ( \1809 , \1808 , \202 );
xor \U$1678 ( \1810 , \1805 , \1809 );
and \U$1679 ( \1811 , \1192 , \215 );
and \U$1680 ( \1812 , \1333 , \213 );
nor \U$1681 ( \1813 , \1811 , \1812 );
xnor \U$1682 ( \1814 , \1813 , \222 );
xor \U$1683 ( \1815 , \1810 , \1814 );
and \U$1684 ( \1816 , \1723 , \1727 );
and \U$1685 ( \1817 , \1727 , \1732 );
and \U$1686 ( \1818 , \1723 , \1732 );
or \U$1687 ( \1819 , \1816 , \1817 , \1818 );
and \U$1688 ( \1820 , \1738 , \1741 );
xor \U$1689 ( \1821 , \1819 , \1820 );
xor \U$1690 ( \1822 , \1693 , \1694 );
not \U$1691 ( \1823 , \1739 );
and \U$1692 ( \1824 , \1822 , \1823 );
and \U$1693 ( \1825 , \166 , \1824 );
and \U$1694 ( \1826 , \150 , \1739 );
nor \U$1695 ( \1827 , \1825 , \1826 );
xnor \U$1696 ( \1828 , \1827 , \1697 );
xor \U$1697 ( \1829 , \1821 , \1828 );
xor \U$1698 ( \1830 , \1815 , \1829 );
and \U$1699 ( \1831 , \474 , \230 );
and \U$1700 ( \1832 , \1147 , \228 );
nor \U$1701 ( \1833 , \1831 , \1832 );
xnor \U$1702 ( \1834 , \1833 , \237 );
and \U$1703 ( \1835 , \307 , \245 );
and \U$1704 ( \1836 , \412 , \243 );
nor \U$1705 ( \1837 , \1835 , \1836 );
xnor \U$1706 ( \1838 , \1837 , \252 );
xor \U$1707 ( \1839 , \1834 , \1838 );
and \U$1708 ( \1840 , \185 , \141 );
and \U$1709 ( \1841 , \261 , \139 );
nor \U$1710 ( \1842 , \1840 , \1841 );
xnor \U$1711 ( \1843 , \1842 , \148 );
xor \U$1712 ( \1844 , \1839 , \1843 );
and \U$1713 ( \1845 , \247 , \1086 );
and \U$1714 ( \1846 , \224 , \508 );
nor \U$1715 ( \1847 , \1845 , \1846 );
xnor \U$1716 ( \1848 , \1847 , \487 );
and \U$1717 ( \1849 , \143 , \1301 );
and \U$1718 ( \1850 , \240 , \1246 );
nor \U$1719 ( \1851 , \1849 , \1850 );
xnor \U$1720 ( \1852 , \1851 , \1205 );
xor \U$1721 ( \1853 , \1848 , \1852 );
and \U$1722 ( \1854 , \158 , \1578 );
and \U$1723 ( \1855 , \134 , \1431 );
nor \U$1724 ( \1856 , \1854 , \1855 );
xnor \U$1725 ( \1857 , \1856 , \1436 );
xor \U$1726 ( \1858 , \1853 , \1857 );
xor \U$1727 ( \1859 , \1844 , \1858 );
and \U$1728 ( \1860 , \197 , \156 );
and \U$1729 ( \1861 , \178 , \154 );
nor \U$1730 ( \1862 , \1860 , \1861 );
xnor \U$1731 ( \1863 , \1862 , \163 );
and \U$1732 ( \1864 , \217 , \296 );
and \U$1733 ( \1865 , \189 , \168 );
nor \U$1734 ( \1866 , \1864 , \1865 );
xnor \U$1735 ( \1867 , \1866 , \173 );
xor \U$1736 ( \1868 , \1863 , \1867 );
and \U$1737 ( \1869 , \232 , \438 );
and \U$1738 ( \1870 , \209 , \336 );
nor \U$1739 ( \1871 , \1869 , \1870 );
xnor \U$1740 ( \1872 , \1871 , \320 );
xor \U$1741 ( \1873 , \1868 , \1872 );
xor \U$1742 ( \1874 , \1859 , \1873 );
xor \U$1743 ( \1875 , \1830 , \1874 );
xor \U$1744 ( \1876 , \1800 , \1875 );
xor \U$1745 ( \1877 , \1786 , \1876 );
and \U$1746 ( \1878 , \1633 , \1644 );
and \U$1747 ( \1879 , \1644 , \1745 );
and \U$1748 ( \1880 , \1633 , \1745 );
or \U$1749 ( \1881 , \1878 , \1879 , \1880 );
xor \U$1750 ( \1882 , \1877 , \1881 );
and \U$1751 ( \1883 , \1746 , \1750 );
and \U$1752 ( \1884 , \1751 , \1754 );
or \U$1753 ( \1885 , \1883 , \1884 );
xor \U$1754 ( \1886 , \1882 , \1885 );
buf \U$1755 ( \1887 , \1886 );
buf \U$1756 ( \1888 , \1887 );
and \U$1757 ( \1889 , \1765 , \1769 );
and \U$1758 ( \1890 , \1769 , \1784 );
and \U$1759 ( \1891 , \1765 , \1784 );
or \U$1760 ( \1892 , \1889 , \1890 , \1891 );
and \U$1761 ( \1893 , \1800 , \1875 );
xor \U$1762 ( \1894 , \1892 , \1893 );
and \U$1763 ( \1895 , \1774 , \1778 );
and \U$1764 ( \1896 , \1778 , \1783 );
and \U$1765 ( \1897 , \1774 , \1783 );
or \U$1766 ( \1898 , \1895 , \1896 , \1897 );
and \U$1767 ( \1899 , \1819 , \1820 );
and \U$1768 ( \1900 , \1820 , \1828 );
and \U$1769 ( \1901 , \1819 , \1828 );
or \U$1770 ( \1902 , \1899 , \1900 , \1901 );
xor \U$1771 ( \1903 , \1898 , \1902 );
and \U$1772 ( \1904 , \1844 , \1858 );
and \U$1773 ( \1905 , \1858 , \1873 );
and \U$1774 ( \1906 , \1844 , \1873 );
or \U$1775 ( \1907 , \1904 , \1905 , \1906 );
xor \U$1776 ( \1908 , \1903 , \1907 );
xor \U$1777 ( \1909 , \1894 , \1908 );
and \U$1778 ( \1910 , \1790 , \1794 );
and \U$1779 ( \1911 , \1794 , \1799 );
and \U$1780 ( \1912 , \1790 , \1799 );
or \U$1781 ( \1913 , \1910 , \1911 , \1912 );
and \U$1782 ( \1914 , \1815 , \1829 );
and \U$1783 ( \1915 , \1829 , \1874 );
and \U$1784 ( \1916 , \1815 , \1874 );
or \U$1785 ( \1917 , \1914 , \1915 , \1916 );
xor \U$1786 ( \1918 , \1913 , \1917 );
and \U$1787 ( \1919 , \1834 , \1838 );
and \U$1788 ( \1920 , \1838 , \1843 );
and \U$1789 ( \1921 , \1834 , \1843 );
or \U$1790 ( \1922 , \1919 , \1920 , \1921 );
and \U$1791 ( \1923 , \1805 , \1809 );
and \U$1792 ( \1924 , \1809 , \1814 );
and \U$1793 ( \1925 , \1805 , \1814 );
or \U$1794 ( \1926 , \1923 , \1924 , \1925 );
xor \U$1795 ( \1927 , \1922 , \1926 );
and \U$1796 ( \1928 , \1863 , \1867 );
and \U$1797 ( \1929 , \1867 , \1872 );
and \U$1798 ( \1930 , \1863 , \1872 );
or \U$1799 ( \1931 , \1928 , \1929 , \1930 );
xor \U$1800 ( \1932 , \1927 , \1931 );
and \U$1801 ( \1933 , \261 , \141 );
and \U$1802 ( \1934 , \307 , \139 );
nor \U$1803 ( \1935 , \1933 , \1934 );
xnor \U$1804 ( \1936 , \1935 , \148 );
and \U$1805 ( \1937 , \178 , \156 );
and \U$1806 ( \1938 , \185 , \154 );
nor \U$1807 ( \1939 , \1937 , \1938 );
xnor \U$1808 ( \1940 , \1939 , \163 );
xor \U$1809 ( \1941 , \1936 , \1940 );
and \U$1810 ( \1942 , \189 , \296 );
and \U$1811 ( \1943 , \197 , \168 );
nor \U$1812 ( \1944 , \1942 , \1943 );
xnor \U$1813 ( \1945 , \1944 , \173 );
xor \U$1814 ( \1946 , \1941 , \1945 );
and \U$1815 ( \1947 , \1802 , \183 );
buf \U$1816 ( \1948 , RIb55e068_102);
and \U$1817 ( \1949 , \1948 , \180 );
nor \U$1818 ( \1950 , \1947 , \1949 );
xnor \U$1819 ( \1951 , \1950 , \179 );
and \U$1820 ( \1952 , \1601 , \195 );
and \U$1821 ( \1953 , \1684 , \193 );
nor \U$1822 ( \1954 , \1952 , \1953 );
xnor \U$1823 ( \1955 , \1954 , \202 );
xor \U$1824 ( \1956 , \1951 , \1955 );
buf \U$1825 ( \1957 , RIb55fee0_37);
buf \U$1826 ( \1958 , RIb55fe68_38);
and \U$1827 ( \1959 , \1958 , \1693 );
not \U$1828 ( \1960 , \1959 );
and \U$1829 ( \1961 , \1957 , \1960 );
xor \U$1830 ( \1962 , \1956 , \1961 );
xor \U$1831 ( \1963 , \1946 , \1962 );
and \U$1832 ( \1964 , \1333 , \215 );
and \U$1833 ( \1965 , \1484 , \213 );
nor \U$1834 ( \1966 , \1964 , \1965 );
xnor \U$1835 ( \1967 , \1966 , \222 );
and \U$1836 ( \1968 , \1147 , \230 );
and \U$1837 ( \1969 , \1192 , \228 );
nor \U$1838 ( \1970 , \1968 , \1969 );
xnor \U$1839 ( \1971 , \1970 , \237 );
xor \U$1840 ( \1972 , \1967 , \1971 );
and \U$1841 ( \1973 , \412 , \245 );
and \U$1842 ( \1974 , \474 , \243 );
nor \U$1843 ( \1975 , \1973 , \1974 );
xnor \U$1844 ( \1976 , \1975 , \252 );
xor \U$1845 ( \1977 , \1972 , \1976 );
xor \U$1846 ( \1978 , \1963 , \1977 );
xor \U$1847 ( \1979 , \1932 , \1978 );
and \U$1848 ( \1980 , \1848 , \1852 );
and \U$1849 ( \1981 , \1852 , \1857 );
and \U$1850 ( \1982 , \1848 , \1857 );
or \U$1851 ( \1983 , \1980 , \1981 , \1982 );
and \U$1852 ( \1984 , \209 , \438 );
and \U$1853 ( \1985 , \217 , \336 );
nor \U$1854 ( \1986 , \1984 , \1985 );
xnor \U$1855 ( \1987 , \1986 , \320 );
and \U$1856 ( \1988 , \224 , \1086 );
and \U$1857 ( \1989 , \232 , \508 );
nor \U$1858 ( \1990 , \1988 , \1989 );
xnor \U$1859 ( \1991 , \1990 , \487 );
xor \U$1860 ( \1992 , \1987 , \1991 );
and \U$1861 ( \1993 , \240 , \1301 );
and \U$1862 ( \1994 , \247 , \1246 );
nor \U$1863 ( \1995 , \1993 , \1994 );
xnor \U$1864 ( \1996 , \1995 , \1205 );
xor \U$1865 ( \1997 , \1992 , \1996 );
xor \U$1866 ( \1998 , \1983 , \1997 );
and \U$1867 ( \1999 , \134 , \1578 );
and \U$1868 ( \2000 , \143 , \1431 );
nor \U$1869 ( \2001 , \1999 , \2000 );
xnor \U$1870 ( \2002 , \2001 , \1436 );
and \U$1871 ( \2003 , \150 , \1824 );
and \U$1872 ( \2004 , \158 , \1739 );
nor \U$1873 ( \2005 , \2003 , \2004 );
xnor \U$1874 ( \2006 , \2005 , \1697 );
xor \U$1875 ( \2007 , \2002 , \2006 );
xor \U$1876 ( \2008 , \1958 , \1693 );
nand \U$1877 ( \2009 , \166 , \2008 );
xnor \U$1878 ( \2010 , \2009 , \1961 );
xor \U$1879 ( \2011 , \2007 , \2010 );
xor \U$1880 ( \2012 , \1998 , \2011 );
xor \U$1881 ( \2013 , \1979 , \2012 );
xor \U$1882 ( \2014 , \1918 , \2013 );
xor \U$1883 ( \2015 , \1909 , \2014 );
and \U$1884 ( \2016 , \1761 , \1785 );
and \U$1885 ( \2017 , \1785 , \1876 );
and \U$1886 ( \2018 , \1761 , \1876 );
or \U$1887 ( \2019 , \2016 , \2017 , \2018 );
xor \U$1888 ( \2020 , \2015 , \2019 );
and \U$1889 ( \2021 , \1877 , \1881 );
and \U$1890 ( \2022 , \1882 , \1885 );
or \U$1891 ( \2023 , \2021 , \2022 );
xor \U$1892 ( \2024 , \2020 , \2023 );
buf \U$1893 ( \2025 , \2024 );
buf \U$1894 ( \2026 , \2025 );
and \U$1895 ( \2027 , \1892 , \1893 );
and \U$1896 ( \2028 , \1893 , \1908 );
and \U$1897 ( \2029 , \1892 , \1908 );
or \U$1898 ( \2030 , \2027 , \2028 , \2029 );
and \U$1899 ( \2031 , \1913 , \1917 );
and \U$1900 ( \2032 , \1917 , \2013 );
and \U$1901 ( \2033 , \1913 , \2013 );
or \U$1902 ( \2034 , \2031 , \2032 , \2033 );
and \U$1903 ( \2035 , \1898 , \1902 );
and \U$1904 ( \2036 , \1902 , \1907 );
and \U$1905 ( \2037 , \1898 , \1907 );
or \U$1906 ( \2038 , \2035 , \2036 , \2037 );
and \U$1907 ( \2039 , \1932 , \1978 );
and \U$1908 ( \2040 , \1978 , \2012 );
and \U$1909 ( \2041 , \1932 , \2012 );
or \U$1910 ( \2042 , \2039 , \2040 , \2041 );
xor \U$1911 ( \2043 , \2038 , \2042 );
and \U$1912 ( \2044 , \1987 , \1991 );
and \U$1913 ( \2045 , \1991 , \1996 );
and \U$1914 ( \2046 , \1987 , \1996 );
or \U$1915 ( \2047 , \2044 , \2045 , \2046 );
and \U$1916 ( \2048 , \2002 , \2006 );
and \U$1917 ( \2049 , \2006 , \2010 );
and \U$1918 ( \2050 , \2002 , \2010 );
or \U$1919 ( \2051 , \2048 , \2049 , \2050 );
xor \U$1920 ( \2052 , \2047 , \2051 );
and \U$1921 ( \2053 , \158 , \1824 );
and \U$1922 ( \2054 , \134 , \1739 );
nor \U$1923 ( \2055 , \2053 , \2054 );
xnor \U$1924 ( \2056 , \2055 , \1697 );
xor \U$1925 ( \2057 , \2052 , \2056 );
xor \U$1926 ( \2058 , \2043 , \2057 );
xor \U$1927 ( \2059 , \2034 , \2058 );
and \U$1928 ( \2060 , \1936 , \1940 );
and \U$1929 ( \2061 , \1940 , \1945 );
and \U$1930 ( \2062 , \1936 , \1945 );
or \U$1931 ( \2063 , \2060 , \2061 , \2062 );
and \U$1932 ( \2064 , \1951 , \1955 );
and \U$1933 ( \2065 , \1955 , \1961 );
and \U$1934 ( \2066 , \1951 , \1961 );
or \U$1935 ( \2067 , \2064 , \2065 , \2066 );
xor \U$1936 ( \2068 , \2063 , \2067 );
and \U$1937 ( \2069 , \1967 , \1971 );
and \U$1938 ( \2070 , \1971 , \1976 );
and \U$1939 ( \2071 , \1967 , \1976 );
or \U$1940 ( \2072 , \2069 , \2070 , \2071 );
xor \U$1941 ( \2073 , \2068 , \2072 );
and \U$1942 ( \2074 , \1922 , \1926 );
and \U$1943 ( \2075 , \1926 , \1931 );
and \U$1944 ( \2076 , \1922 , \1931 );
or \U$1945 ( \2077 , \2074 , \2075 , \2076 );
and \U$1946 ( \2078 , \1946 , \1962 );
and \U$1947 ( \2079 , \1962 , \1977 );
and \U$1948 ( \2080 , \1946 , \1977 );
or \U$1949 ( \2081 , \2078 , \2079 , \2080 );
xor \U$1950 ( \2082 , \2077 , \2081 );
and \U$1951 ( \2083 , \1983 , \1997 );
and \U$1952 ( \2084 , \1997 , \2011 );
and \U$1953 ( \2085 , \1983 , \2011 );
or \U$1954 ( \2086 , \2083 , \2084 , \2085 );
xor \U$1955 ( \2087 , \2082 , \2086 );
xor \U$1956 ( \2088 , \2073 , \2087 );
and \U$1957 ( \2089 , \1948 , \183 );
buf \U$1958 ( \2090 , RIb55e0e0_101);
and \U$1959 ( \2091 , \2090 , \180 );
nor \U$1960 ( \2092 , \2089 , \2091 );
xnor \U$1961 ( \2093 , \2092 , \179 );
and \U$1962 ( \2094 , \1684 , \195 );
and \U$1963 ( \2095 , \1802 , \193 );
nor \U$1964 ( \2096 , \2094 , \2095 );
xnor \U$1965 ( \2097 , \2096 , \202 );
xor \U$1966 ( \2098 , \2093 , \2097 );
and \U$1967 ( \2099 , \1484 , \215 );
and \U$1968 ( \2100 , \1601 , \213 );
nor \U$1969 ( \2101 , \2099 , \2100 );
xnor \U$1970 ( \2102 , \2101 , \222 );
xor \U$1971 ( \2103 , \2098 , \2102 );
and \U$1972 ( \2104 , \1192 , \230 );
and \U$1973 ( \2105 , \1333 , \228 );
nor \U$1974 ( \2106 , \2104 , \2105 );
xnor \U$1975 ( \2107 , \2106 , \237 );
and \U$1976 ( \2108 , \474 , \245 );
and \U$1977 ( \2109 , \1147 , \243 );
nor \U$1978 ( \2110 , \2108 , \2109 );
xnor \U$1979 ( \2111 , \2110 , \252 );
xor \U$1980 ( \2112 , \2107 , \2111 );
and \U$1981 ( \2113 , \307 , \141 );
and \U$1982 ( \2114 , \412 , \139 );
nor \U$1983 ( \2115 , \2113 , \2114 );
xnor \U$1984 ( \2116 , \2115 , \148 );
xor \U$1985 ( \2117 , \2112 , \2116 );
xor \U$1986 ( \2118 , \2103 , \2117 );
xor \U$1987 ( \2119 , \1957 , \1958 );
not \U$1988 ( \2120 , \2008 );
and \U$1989 ( \2121 , \2119 , \2120 );
and \U$1990 ( \2122 , \166 , \2121 );
and \U$1991 ( \2123 , \150 , \2008 );
nor \U$1992 ( \2124 , \2122 , \2123 );
xnor \U$1993 ( \2125 , \2124 , \1961 );
and \U$1994 ( \2126 , \232 , \1086 );
and \U$1995 ( \2127 , \209 , \508 );
nor \U$1996 ( \2128 , \2126 , \2127 );
xnor \U$1997 ( \2129 , \2128 , \487 );
and \U$1998 ( \2130 , \247 , \1301 );
and \U$1999 ( \2131 , \224 , \1246 );
nor \U$2000 ( \2132 , \2130 , \2131 );
xnor \U$2001 ( \2133 , \2132 , \1205 );
xor \U$2002 ( \2134 , \2129 , \2133 );
and \U$2003 ( \2135 , \143 , \1578 );
and \U$2004 ( \2136 , \240 , \1431 );
nor \U$2005 ( \2137 , \2135 , \2136 );
xnor \U$2006 ( \2138 , \2137 , \1436 );
xor \U$2007 ( \2139 , \2134 , \2138 );
xor \U$2008 ( \2140 , \2125 , \2139 );
and \U$2009 ( \2141 , \185 , \156 );
and \U$2010 ( \2142 , \261 , \154 );
nor \U$2011 ( \2143 , \2141 , \2142 );
xnor \U$2012 ( \2144 , \2143 , \163 );
and \U$2013 ( \2145 , \197 , \296 );
and \U$2014 ( \2146 , \178 , \168 );
nor \U$2015 ( \2147 , \2145 , \2146 );
xnor \U$2016 ( \2148 , \2147 , \173 );
xor \U$2017 ( \2149 , \2144 , \2148 );
and \U$2018 ( \2150 , \217 , \438 );
and \U$2019 ( \2151 , \189 , \336 );
nor \U$2020 ( \2152 , \2150 , \2151 );
xnor \U$2021 ( \2153 , \2152 , \320 );
xor \U$2022 ( \2154 , \2149 , \2153 );
xor \U$2023 ( \2155 , \2140 , \2154 );
xor \U$2024 ( \2156 , \2118 , \2155 );
xor \U$2025 ( \2157 , \2088 , \2156 );
xor \U$2026 ( \2158 , \2059 , \2157 );
xor \U$2027 ( \2159 , \2030 , \2158 );
and \U$2028 ( \2160 , \1909 , \2014 );
xor \U$2029 ( \2161 , \2159 , \2160 );
and \U$2030 ( \2162 , \2015 , \2019 );
and \U$2031 ( \2163 , \2020 , \2023 );
or \U$2032 ( \2164 , \2162 , \2163 );
xor \U$2033 ( \2165 , \2161 , \2164 );
buf \U$2034 ( \2166 , \2165 );
buf \U$2035 ( \2167 , \2166 );
and \U$2036 ( \2168 , \2034 , \2058 );
and \U$2037 ( \2169 , \2058 , \2157 );
and \U$2038 ( \2170 , \2034 , \2157 );
or \U$2039 ( \2171 , \2168 , \2169 , \2170 );
and \U$2040 ( \2172 , \2038 , \2042 );
and \U$2041 ( \2173 , \2042 , \2057 );
and \U$2042 ( \2174 , \2038 , \2057 );
or \U$2043 ( \2175 , \2172 , \2173 , \2174 );
and \U$2044 ( \2176 , \2073 , \2087 );
and \U$2045 ( \2177 , \2087 , \2156 );
and \U$2046 ( \2178 , \2073 , \2156 );
or \U$2047 ( \2179 , \2176 , \2177 , \2178 );
xor \U$2048 ( \2180 , \2175 , \2179 );
and \U$2049 ( \2181 , \2090 , \183 );
buf \U$2050 ( \2182 , RIb55e158_100);
and \U$2051 ( \2183 , \2182 , \180 );
nor \U$2052 ( \2184 , \2181 , \2183 );
xnor \U$2053 ( \2185 , \2184 , \179 );
and \U$2054 ( \2186 , \1802 , \195 );
and \U$2055 ( \2187 , \1948 , \193 );
nor \U$2056 ( \2188 , \2186 , \2187 );
xnor \U$2057 ( \2189 , \2188 , \202 );
xor \U$2058 ( \2190 , \2185 , \2189 );
buf \U$2059 ( \2191 , RIb55ffd0_35);
buf \U$2060 ( \2192 , RIb55ff58_36);
and \U$2061 ( \2193 , \2192 , \1957 );
not \U$2062 ( \2194 , \2193 );
and \U$2063 ( \2195 , \2191 , \2194 );
xor \U$2064 ( \2196 , \2190 , \2195 );
and \U$2065 ( \2197 , \412 , \141 );
and \U$2066 ( \2198 , \474 , \139 );
nor \U$2067 ( \2199 , \2197 , \2198 );
xnor \U$2068 ( \2200 , \2199 , \148 );
and \U$2069 ( \2201 , \261 , \156 );
and \U$2070 ( \2202 , \307 , \154 );
nor \U$2071 ( \2203 , \2201 , \2202 );
xnor \U$2072 ( \2204 , \2203 , \163 );
xor \U$2073 ( \2205 , \2200 , \2204 );
and \U$2074 ( \2206 , \178 , \296 );
and \U$2075 ( \2207 , \185 , \168 );
nor \U$2076 ( \2208 , \2206 , \2207 );
xnor \U$2077 ( \2209 , \2208 , \173 );
xor \U$2078 ( \2210 , \2205 , \2209 );
and \U$2079 ( \2211 , \1601 , \215 );
and \U$2080 ( \2212 , \1684 , \213 );
nor \U$2081 ( \2213 , \2211 , \2212 );
xnor \U$2082 ( \2214 , \2213 , \222 );
and \U$2083 ( \2215 , \1333 , \230 );
and \U$2084 ( \2216 , \1484 , \228 );
nor \U$2085 ( \2217 , \2215 , \2216 );
xnor \U$2086 ( \2218 , \2217 , \237 );
xor \U$2087 ( \2219 , \2214 , \2218 );
and \U$2088 ( \2220 , \1147 , \245 );
and \U$2089 ( \2221 , \1192 , \243 );
nor \U$2090 ( \2222 , \2220 , \2221 );
xnor \U$2091 ( \2223 , \2222 , \252 );
xor \U$2092 ( \2224 , \2219 , \2223 );
xor \U$2093 ( \2225 , \2210 , \2224 );
and \U$2094 ( \2226 , \189 , \438 );
and \U$2095 ( \2227 , \197 , \336 );
nor \U$2096 ( \2228 , \2226 , \2227 );
xnor \U$2097 ( \2229 , \2228 , \320 );
and \U$2098 ( \2230 , \209 , \1086 );
and \U$2099 ( \2231 , \217 , \508 );
nor \U$2100 ( \2232 , \2230 , \2231 );
xnor \U$2101 ( \2233 , \2232 , \487 );
xor \U$2102 ( \2234 , \2229 , \2233 );
and \U$2103 ( \2235 , \224 , \1301 );
and \U$2104 ( \2236 , \232 , \1246 );
nor \U$2105 ( \2237 , \2235 , \2236 );
xnor \U$2106 ( \2238 , \2237 , \1205 );
xor \U$2107 ( \2239 , \2234 , \2238 );
xor \U$2108 ( \2240 , \2225 , \2239 );
xor \U$2109 ( \2241 , \2196 , \2240 );
and \U$2110 ( \2242 , \2129 , \2133 );
and \U$2111 ( \2243 , \2133 , \2138 );
and \U$2112 ( \2244 , \2129 , \2138 );
or \U$2113 ( \2245 , \2242 , \2243 , \2244 );
xor \U$2114 ( \2246 , \2192 , \1957 );
nand \U$2115 ( \2247 , \166 , \2246 );
xnor \U$2116 ( \2248 , \2247 , \2195 );
xor \U$2117 ( \2249 , \2245 , \2248 );
and \U$2118 ( \2250 , \240 , \1578 );
and \U$2119 ( \2251 , \247 , \1431 );
nor \U$2120 ( \2252 , \2250 , \2251 );
xnor \U$2121 ( \2253 , \2252 , \1436 );
and \U$2122 ( \2254 , \134 , \1824 );
and \U$2123 ( \2255 , \143 , \1739 );
nor \U$2124 ( \2256 , \2254 , \2255 );
xnor \U$2125 ( \2257 , \2256 , \1697 );
xor \U$2126 ( \2258 , \2253 , \2257 );
and \U$2127 ( \2259 , \150 , \2121 );
and \U$2128 ( \2260 , \158 , \2008 );
nor \U$2129 ( \2261 , \2259 , \2260 );
xnor \U$2130 ( \2262 , \2261 , \1961 );
xor \U$2131 ( \2263 , \2258 , \2262 );
xor \U$2132 ( \2264 , \2249 , \2263 );
xor \U$2133 ( \2265 , \2241 , \2264 );
xor \U$2134 ( \2266 , \2180 , \2265 );
xor \U$2135 ( \2267 , \2171 , \2266 );
and \U$2136 ( \2268 , \2047 , \2051 );
and \U$2137 ( \2269 , \2051 , \2056 );
and \U$2138 ( \2270 , \2047 , \2056 );
or \U$2139 ( \2271 , \2268 , \2269 , \2270 );
and \U$2140 ( \2272 , \2063 , \2067 );
and \U$2141 ( \2273 , \2067 , \2072 );
and \U$2142 ( \2274 , \2063 , \2072 );
or \U$2143 ( \2275 , \2272 , \2273 , \2274 );
xor \U$2144 ( \2276 , \2271 , \2275 );
and \U$2145 ( \2277 , \2125 , \2139 );
and \U$2146 ( \2278 , \2139 , \2154 );
and \U$2147 ( \2279 , \2125 , \2154 );
or \U$2148 ( \2280 , \2277 , \2278 , \2279 );
xor \U$2149 ( \2281 , \2276 , \2280 );
and \U$2150 ( \2282 , \2077 , \2081 );
and \U$2151 ( \2283 , \2081 , \2086 );
and \U$2152 ( \2284 , \2077 , \2086 );
or \U$2153 ( \2285 , \2282 , \2283 , \2284 );
and \U$2154 ( \2286 , \2103 , \2117 );
and \U$2155 ( \2287 , \2117 , \2155 );
and \U$2156 ( \2288 , \2103 , \2155 );
or \U$2157 ( \2289 , \2286 , \2287 , \2288 );
xor \U$2158 ( \2290 , \2285 , \2289 );
and \U$2159 ( \2291 , \2093 , \2097 );
and \U$2160 ( \2292 , \2097 , \2102 );
and \U$2161 ( \2293 , \2093 , \2102 );
or \U$2162 ( \2294 , \2291 , \2292 , \2293 );
and \U$2163 ( \2295 , \2144 , \2148 );
and \U$2164 ( \2296 , \2148 , \2153 );
and \U$2165 ( \2297 , \2144 , \2153 );
or \U$2166 ( \2298 , \2295 , \2296 , \2297 );
xor \U$2167 ( \2299 , \2294 , \2298 );
and \U$2168 ( \2300 , \2107 , \2111 );
and \U$2169 ( \2301 , \2111 , \2116 );
and \U$2170 ( \2302 , \2107 , \2116 );
or \U$2171 ( \2303 , \2300 , \2301 , \2302 );
xor \U$2172 ( \2304 , \2299 , \2303 );
xor \U$2173 ( \2305 , \2290 , \2304 );
xor \U$2174 ( \2306 , \2281 , \2305 );
xor \U$2175 ( \2307 , \2267 , \2306 );
and \U$2176 ( \2308 , \2030 , \2158 );
xor \U$2177 ( \2309 , \2307 , \2308 );
and \U$2178 ( \2310 , \2159 , \2160 );
and \U$2179 ( \2311 , \2161 , \2164 );
or \U$2180 ( \2312 , \2310 , \2311 );
xor \U$2181 ( \2313 , \2309 , \2312 );
buf \U$2182 ( \2314 , \2313 );
buf \U$2183 ( \2315 , \2314 );
and \U$2184 ( \2316 , \2175 , \2179 );
and \U$2185 ( \2317 , \2179 , \2265 );
and \U$2186 ( \2318 , \2175 , \2265 );
or \U$2187 ( \2319 , \2316 , \2317 , \2318 );
and \U$2188 ( \2320 , \2281 , \2305 );
xor \U$2189 ( \2321 , \2319 , \2320 );
and \U$2190 ( \2322 , \2285 , \2289 );
and \U$2191 ( \2323 , \2289 , \2304 );
and \U$2192 ( \2324 , \2285 , \2304 );
or \U$2193 ( \2325 , \2322 , \2323 , \2324 );
and \U$2194 ( \2326 , \2271 , \2275 );
and \U$2195 ( \2327 , \2275 , \2280 );
and \U$2196 ( \2328 , \2271 , \2280 );
or \U$2197 ( \2329 , \2326 , \2327 , \2328 );
and \U$2198 ( \2330 , \2196 , \2240 );
and \U$2199 ( \2331 , \2240 , \2264 );
and \U$2200 ( \2332 , \2196 , \2264 );
or \U$2201 ( \2333 , \2330 , \2331 , \2332 );
xor \U$2202 ( \2334 , \2329 , \2333 );
and \U$2203 ( \2335 , \2200 , \2204 );
and \U$2204 ( \2336 , \2204 , \2209 );
and \U$2205 ( \2337 , \2200 , \2209 );
or \U$2206 ( \2338 , \2335 , \2336 , \2337 );
and \U$2207 ( \2339 , \2214 , \2218 );
and \U$2208 ( \2340 , \2218 , \2223 );
and \U$2209 ( \2341 , \2214 , \2223 );
or \U$2210 ( \2342 , \2339 , \2340 , \2341 );
xor \U$2211 ( \2343 , \2338 , \2342 );
and \U$2212 ( \2344 , \2185 , \2189 );
and \U$2213 ( \2345 , \2189 , \2195 );
and \U$2214 ( \2346 , \2185 , \2195 );
or \U$2215 ( \2347 , \2344 , \2345 , \2346 );
xor \U$2216 ( \2348 , \2343 , \2347 );
xor \U$2217 ( \2349 , \2334 , \2348 );
xor \U$2218 ( \2350 , \2325 , \2349 );
and \U$2219 ( \2351 , \2294 , \2298 );
and \U$2220 ( \2352 , \2298 , \2303 );
and \U$2221 ( \2353 , \2294 , \2303 );
or \U$2222 ( \2354 , \2351 , \2352 , \2353 );
and \U$2223 ( \2355 , \2210 , \2224 );
and \U$2224 ( \2356 , \2224 , \2239 );
and \U$2225 ( \2357 , \2210 , \2239 );
or \U$2226 ( \2358 , \2355 , \2356 , \2357 );
xor \U$2227 ( \2359 , \2354 , \2358 );
and \U$2228 ( \2360 , \2245 , \2248 );
and \U$2229 ( \2361 , \2248 , \2263 );
and \U$2230 ( \2362 , \2245 , \2263 );
or \U$2231 ( \2363 , \2360 , \2361 , \2362 );
xor \U$2232 ( \2364 , \2359 , \2363 );
and \U$2233 ( \2365 , \2182 , \183 );
buf \U$2234 ( \2366 , RIb55e1d0_99);
and \U$2235 ( \2367 , \2366 , \180 );
nor \U$2236 ( \2368 , \2365 , \2367 );
xnor \U$2237 ( \2369 , \2368 , \179 );
and \U$2238 ( \2370 , \1948 , \195 );
and \U$2239 ( \2371 , \2090 , \193 );
nor \U$2240 ( \2372 , \2370 , \2371 );
xnor \U$2241 ( \2373 , \2372 , \202 );
xor \U$2242 ( \2374 , \2369 , \2373 );
and \U$2243 ( \2375 , \1684 , \215 );
and \U$2244 ( \2376 , \1802 , \213 );
nor \U$2245 ( \2377 , \2375 , \2376 );
xnor \U$2246 ( \2378 , \2377 , \222 );
xor \U$2247 ( \2379 , \2374 , \2378 );
and \U$2248 ( \2380 , \2229 , \2233 );
and \U$2249 ( \2381 , \2233 , \2238 );
and \U$2250 ( \2382 , \2229 , \2238 );
or \U$2251 ( \2383 , \2380 , \2381 , \2382 );
and \U$2252 ( \2384 , \2253 , \2257 );
and \U$2253 ( \2385 , \2257 , \2262 );
and \U$2254 ( \2386 , \2253 , \2262 );
or \U$2255 ( \2387 , \2384 , \2385 , \2386 );
xor \U$2256 ( \2388 , \2383 , \2387 );
and \U$2257 ( \2389 , \143 , \1824 );
and \U$2258 ( \2390 , \240 , \1739 );
nor \U$2259 ( \2391 , \2389 , \2390 );
xnor \U$2260 ( \2392 , \2391 , \1697 );
and \U$2261 ( \2393 , \158 , \2121 );
and \U$2262 ( \2394 , \134 , \2008 );
nor \U$2263 ( \2395 , \2393 , \2394 );
xnor \U$2264 ( \2396 , \2395 , \1961 );
xor \U$2265 ( \2397 , \2392 , \2396 );
xor \U$2266 ( \2398 , \2191 , \2192 );
not \U$2267 ( \2399 , \2246 );
and \U$2268 ( \2400 , \2398 , \2399 );
and \U$2269 ( \2401 , \166 , \2400 );
and \U$2270 ( \2402 , \150 , \2246 );
nor \U$2271 ( \2403 , \2401 , \2402 );
xnor \U$2272 ( \2404 , \2403 , \2195 );
xor \U$2273 ( \2405 , \2397 , \2404 );
xor \U$2274 ( \2406 , \2388 , \2405 );
xor \U$2275 ( \2407 , \2379 , \2406 );
and \U$2276 ( \2408 , \307 , \156 );
and \U$2277 ( \2409 , \412 , \154 );
nor \U$2278 ( \2410 , \2408 , \2409 );
xnor \U$2279 ( \2411 , \2410 , \163 );
and \U$2280 ( \2412 , \185 , \296 );
and \U$2281 ( \2413 , \261 , \168 );
nor \U$2282 ( \2414 , \2412 , \2413 );
xnor \U$2283 ( \2415 , \2414 , \173 );
xor \U$2284 ( \2416 , \2411 , \2415 );
and \U$2285 ( \2417 , \197 , \438 );
and \U$2286 ( \2418 , \178 , \336 );
nor \U$2287 ( \2419 , \2417 , \2418 );
xnor \U$2288 ( \2420 , \2419 , \320 );
xor \U$2289 ( \2421 , \2416 , \2420 );
and \U$2290 ( \2422 , \1484 , \230 );
and \U$2291 ( \2423 , \1601 , \228 );
nor \U$2292 ( \2424 , \2422 , \2423 );
xnor \U$2293 ( \2425 , \2424 , \237 );
and \U$2294 ( \2426 , \1192 , \245 );
and \U$2295 ( \2427 , \1333 , \243 );
nor \U$2296 ( \2428 , \2426 , \2427 );
xnor \U$2297 ( \2429 , \2428 , \252 );
xor \U$2298 ( \2430 , \2425 , \2429 );
and \U$2299 ( \2431 , \474 , \141 );
and \U$2300 ( \2432 , \1147 , \139 );
nor \U$2301 ( \2433 , \2431 , \2432 );
xnor \U$2302 ( \2434 , \2433 , \148 );
xor \U$2303 ( \2435 , \2430 , \2434 );
xor \U$2304 ( \2436 , \2421 , \2435 );
and \U$2305 ( \2437 , \217 , \1086 );
and \U$2306 ( \2438 , \189 , \508 );
nor \U$2307 ( \2439 , \2437 , \2438 );
xnor \U$2308 ( \2440 , \2439 , \487 );
and \U$2309 ( \2441 , \232 , \1301 );
and \U$2310 ( \2442 , \209 , \1246 );
nor \U$2311 ( \2443 , \2441 , \2442 );
xnor \U$2312 ( \2444 , \2443 , \1205 );
xor \U$2313 ( \2445 , \2440 , \2444 );
and \U$2314 ( \2446 , \247 , \1578 );
and \U$2315 ( \2447 , \224 , \1431 );
nor \U$2316 ( \2448 , \2446 , \2447 );
xnor \U$2317 ( \2449 , \2448 , \1436 );
xor \U$2318 ( \2450 , \2445 , \2449 );
xor \U$2319 ( \2451 , \2436 , \2450 );
xor \U$2320 ( \2452 , \2407 , \2451 );
xor \U$2321 ( \2453 , \2364 , \2452 );
xor \U$2322 ( \2454 , \2350 , \2453 );
xor \U$2323 ( \2455 , \2321 , \2454 );
and \U$2324 ( \2456 , \2171 , \2266 );
and \U$2325 ( \2457 , \2266 , \2306 );
and \U$2326 ( \2458 , \2171 , \2306 );
or \U$2327 ( \2459 , \2456 , \2457 , \2458 );
xor \U$2328 ( \2460 , \2455 , \2459 );
and \U$2329 ( \2461 , \2307 , \2308 );
and \U$2330 ( \2462 , \2309 , \2312 );
or \U$2331 ( \2463 , \2461 , \2462 );
xor \U$2332 ( \2464 , \2460 , \2463 );
buf \U$2333 ( \2465 , \2464 );
buf \U$2334 ( \2466 , \2465 );
and \U$2335 ( \2467 , \2325 , \2349 );
and \U$2336 ( \2468 , \2349 , \2453 );
and \U$2337 ( \2469 , \2325 , \2453 );
or \U$2338 ( \2470 , \2467 , \2468 , \2469 );
and \U$2339 ( \2471 , \2329 , \2333 );
and \U$2340 ( \2472 , \2333 , \2348 );
and \U$2341 ( \2473 , \2329 , \2348 );
or \U$2342 ( \2474 , \2471 , \2472 , \2473 );
and \U$2343 ( \2475 , \2364 , \2452 );
xor \U$2344 ( \2476 , \2474 , \2475 );
and \U$2345 ( \2477 , \2392 , \2396 );
and \U$2346 ( \2478 , \2396 , \2404 );
and \U$2347 ( \2479 , \2392 , \2404 );
or \U$2348 ( \2480 , \2477 , \2478 , \2479 );
and \U$2349 ( \2481 , \2440 , \2444 );
and \U$2350 ( \2482 , \2444 , \2449 );
and \U$2351 ( \2483 , \2440 , \2449 );
or \U$2352 ( \2484 , \2481 , \2482 , \2483 );
xor \U$2353 ( \2485 , \2480 , \2484 );
and \U$2354 ( \2486 , \150 , \2400 );
and \U$2355 ( \2487 , \158 , \2246 );
nor \U$2356 ( \2488 , \2486 , \2487 );
xnor \U$2357 ( \2489 , \2488 , \2195 );
xor \U$2358 ( \2490 , \2485 , \2489 );
and \U$2359 ( \2491 , \1802 , \215 );
and \U$2360 ( \2492 , \1948 , \213 );
nor \U$2361 ( \2493 , \2491 , \2492 );
xnor \U$2362 ( \2494 , \2493 , \222 );
and \U$2363 ( \2495 , \1601 , \230 );
and \U$2364 ( \2496 , \1684 , \228 );
nor \U$2365 ( \2497 , \2495 , \2496 );
xnor \U$2366 ( \2498 , \2497 , \237 );
xor \U$2367 ( \2499 , \2494 , \2498 );
and \U$2368 ( \2500 , \1333 , \245 );
and \U$2369 ( \2501 , \1484 , \243 );
nor \U$2370 ( \2502 , \2500 , \2501 );
xnor \U$2371 ( \2503 , \2502 , \252 );
xor \U$2372 ( \2504 , \2499 , \2503 );
and \U$2373 ( \2505 , \1147 , \141 );
and \U$2374 ( \2506 , \1192 , \139 );
nor \U$2375 ( \2507 , \2505 , \2506 );
xnor \U$2376 ( \2508 , \2507 , \148 );
and \U$2377 ( \2509 , \412 , \156 );
and \U$2378 ( \2510 , \474 , \154 );
nor \U$2379 ( \2511 , \2509 , \2510 );
xnor \U$2380 ( \2512 , \2511 , \163 );
xor \U$2381 ( \2513 , \2508 , \2512 );
and \U$2382 ( \2514 , \261 , \296 );
and \U$2383 ( \2515 , \307 , \168 );
nor \U$2384 ( \2516 , \2514 , \2515 );
xnor \U$2385 ( \2517 , \2516 , \173 );
xor \U$2386 ( \2518 , \2513 , \2517 );
xor \U$2387 ( \2519 , \2504 , \2518 );
and \U$2388 ( \2520 , \2366 , \183 );
buf \U$2389 ( \2521 , RIb55e248_98);
and \U$2390 ( \2522 , \2521 , \180 );
nor \U$2391 ( \2523 , \2520 , \2522 );
xnor \U$2392 ( \2524 , \2523 , \179 );
and \U$2393 ( \2525 , \2090 , \195 );
and \U$2394 ( \2526 , \2182 , \193 );
nor \U$2395 ( \2527 , \2525 , \2526 );
xnor \U$2396 ( \2528 , \2527 , \202 );
xor \U$2397 ( \2529 , \2524 , \2528 );
buf \U$2398 ( \2530 , RIb5600c0_33);
buf \U$2399 ( \2531 , RIb560048_34);
and \U$2400 ( \2532 , \2531 , \2191 );
not \U$2401 ( \2533 , \2532 );
and \U$2402 ( \2534 , \2530 , \2533 );
xor \U$2403 ( \2535 , \2529 , \2534 );
xor \U$2404 ( \2536 , \2519 , \2535 );
xor \U$2405 ( \2537 , \2490 , \2536 );
xor \U$2406 ( \2538 , \2531 , \2191 );
nand \U$2407 ( \2539 , \166 , \2538 );
xnor \U$2408 ( \2540 , \2539 , \2534 );
and \U$2409 ( \2541 , \224 , \1578 );
and \U$2410 ( \2542 , \232 , \1431 );
nor \U$2411 ( \2543 , \2541 , \2542 );
xnor \U$2412 ( \2544 , \2543 , \1436 );
and \U$2413 ( \2545 , \240 , \1824 );
and \U$2414 ( \2546 , \247 , \1739 );
nor \U$2415 ( \2547 , \2545 , \2546 );
xnor \U$2416 ( \2548 , \2547 , \1697 );
xor \U$2417 ( \2549 , \2544 , \2548 );
and \U$2418 ( \2550 , \134 , \2121 );
and \U$2419 ( \2551 , \143 , \2008 );
nor \U$2420 ( \2552 , \2550 , \2551 );
xnor \U$2421 ( \2553 , \2552 , \1961 );
xor \U$2422 ( \2554 , \2549 , \2553 );
xor \U$2423 ( \2555 , \2540 , \2554 );
and \U$2424 ( \2556 , \178 , \438 );
and \U$2425 ( \2557 , \185 , \336 );
nor \U$2426 ( \2558 , \2556 , \2557 );
xnor \U$2427 ( \2559 , \2558 , \320 );
and \U$2428 ( \2560 , \189 , \1086 );
and \U$2429 ( \2561 , \197 , \508 );
nor \U$2430 ( \2562 , \2560 , \2561 );
xnor \U$2431 ( \2563 , \2562 , \487 );
xor \U$2432 ( \2564 , \2559 , \2563 );
and \U$2433 ( \2565 , \209 , \1301 );
and \U$2434 ( \2566 , \217 , \1246 );
nor \U$2435 ( \2567 , \2565 , \2566 );
xnor \U$2436 ( \2568 , \2567 , \1205 );
xor \U$2437 ( \2569 , \2564 , \2568 );
xor \U$2438 ( \2570 , \2555 , \2569 );
xor \U$2439 ( \2571 , \2537 , \2570 );
xor \U$2440 ( \2572 , \2476 , \2571 );
xor \U$2441 ( \2573 , \2470 , \2572 );
and \U$2442 ( \2574 , \2338 , \2342 );
and \U$2443 ( \2575 , \2342 , \2347 );
and \U$2444 ( \2576 , \2338 , \2347 );
or \U$2445 ( \2577 , \2574 , \2575 , \2576 );
and \U$2446 ( \2578 , \2383 , \2387 );
and \U$2447 ( \2579 , \2387 , \2405 );
and \U$2448 ( \2580 , \2383 , \2405 );
or \U$2449 ( \2581 , \2578 , \2579 , \2580 );
xor \U$2450 ( \2582 , \2577 , \2581 );
and \U$2451 ( \2583 , \2421 , \2435 );
and \U$2452 ( \2584 , \2435 , \2450 );
and \U$2453 ( \2585 , \2421 , \2450 );
or \U$2454 ( \2586 , \2583 , \2584 , \2585 );
xor \U$2455 ( \2587 , \2582 , \2586 );
and \U$2456 ( \2588 , \2354 , \2358 );
and \U$2457 ( \2589 , \2358 , \2363 );
and \U$2458 ( \2590 , \2354 , \2363 );
or \U$2459 ( \2591 , \2588 , \2589 , \2590 );
and \U$2460 ( \2592 , \2379 , \2406 );
and \U$2461 ( \2593 , \2406 , \2451 );
and \U$2462 ( \2594 , \2379 , \2451 );
or \U$2463 ( \2595 , \2592 , \2593 , \2594 );
xor \U$2464 ( \2596 , \2591 , \2595 );
and \U$2465 ( \2597 , \2411 , \2415 );
and \U$2466 ( \2598 , \2415 , \2420 );
and \U$2467 ( \2599 , \2411 , \2420 );
or \U$2468 ( \2600 , \2597 , \2598 , \2599 );
and \U$2469 ( \2601 , \2425 , \2429 );
and \U$2470 ( \2602 , \2429 , \2434 );
and \U$2471 ( \2603 , \2425 , \2434 );
or \U$2472 ( \2604 , \2601 , \2602 , \2603 );
xor \U$2473 ( \2605 , \2600 , \2604 );
and \U$2474 ( \2606 , \2369 , \2373 );
and \U$2475 ( \2607 , \2373 , \2378 );
and \U$2476 ( \2608 , \2369 , \2378 );
or \U$2477 ( \2609 , \2606 , \2607 , \2608 );
xor \U$2478 ( \2610 , \2605 , \2609 );
xor \U$2479 ( \2611 , \2596 , \2610 );
xor \U$2480 ( \2612 , \2587 , \2611 );
xor \U$2481 ( \2613 , \2573 , \2612 );
and \U$2482 ( \2614 , \2319 , \2320 );
and \U$2483 ( \2615 , \2320 , \2454 );
and \U$2484 ( \2616 , \2319 , \2454 );
or \U$2485 ( \2617 , \2614 , \2615 , \2616 );
xor \U$2486 ( \2618 , \2613 , \2617 );
and \U$2487 ( \2619 , \2455 , \2459 );
and \U$2488 ( \2620 , \2460 , \2463 );
or \U$2489 ( \2621 , \2619 , \2620 );
xor \U$2490 ( \2622 , \2618 , \2621 );
buf \U$2491 ( \2623 , \2622 );
buf \U$2492 ( \2624 , \2623 );
and \U$2493 ( \2625 , \2474 , \2475 );
and \U$2494 ( \2626 , \2475 , \2571 );
and \U$2495 ( \2627 , \2474 , \2571 );
or \U$2496 ( \2628 , \2625 , \2626 , \2627 );
and \U$2497 ( \2629 , \2587 , \2611 );
xor \U$2498 ( \2630 , \2628 , \2629 );
and \U$2499 ( \2631 , \2591 , \2595 );
and \U$2500 ( \2632 , \2595 , \2610 );
and \U$2501 ( \2633 , \2591 , \2610 );
or \U$2502 ( \2634 , \2631 , \2632 , \2633 );
and \U$2503 ( \2635 , \2577 , \2581 );
and \U$2504 ( \2636 , \2581 , \2586 );
and \U$2505 ( \2637 , \2577 , \2586 );
or \U$2506 ( \2638 , \2635 , \2636 , \2637 );
and \U$2507 ( \2639 , \2490 , \2536 );
and \U$2508 ( \2640 , \2536 , \2570 );
and \U$2509 ( \2641 , \2490 , \2570 );
or \U$2510 ( \2642 , \2639 , \2640 , \2641 );
xor \U$2511 ( \2643 , \2638 , \2642 );
and \U$2512 ( \2644 , \2494 , \2498 );
and \U$2513 ( \2645 , \2498 , \2503 );
and \U$2514 ( \2646 , \2494 , \2503 );
or \U$2515 ( \2647 , \2644 , \2645 , \2646 );
and \U$2516 ( \2648 , \2508 , \2512 );
and \U$2517 ( \2649 , \2512 , \2517 );
and \U$2518 ( \2650 , \2508 , \2517 );
or \U$2519 ( \2651 , \2648 , \2649 , \2650 );
xor \U$2520 ( \2652 , \2647 , \2651 );
and \U$2521 ( \2653 , \2524 , \2528 );
and \U$2522 ( \2654 , \2528 , \2534 );
and \U$2523 ( \2655 , \2524 , \2534 );
or \U$2524 ( \2656 , \2653 , \2654 , \2655 );
xor \U$2525 ( \2657 , \2652 , \2656 );
and \U$2526 ( \2658 , \2544 , \2548 );
and \U$2527 ( \2659 , \2548 , \2553 );
and \U$2528 ( \2660 , \2544 , \2553 );
or \U$2529 ( \2661 , \2658 , \2659 , \2660 );
and \U$2530 ( \2662 , \2559 , \2563 );
and \U$2531 ( \2663 , \2563 , \2568 );
and \U$2532 ( \2664 , \2559 , \2568 );
or \U$2533 ( \2665 , \2662 , \2663 , \2664 );
xor \U$2534 ( \2666 , \2661 , \2665 );
xor \U$2535 ( \2667 , \2530 , \2531 );
not \U$2536 ( \2668 , \2538 );
and \U$2537 ( \2669 , \2667 , \2668 );
and \U$2538 ( \2670 , \166 , \2669 );
and \U$2539 ( \2671 , \150 , \2538 );
nor \U$2540 ( \2672 , \2670 , \2671 );
xnor \U$2541 ( \2673 , \2672 , \2534 );
xor \U$2542 ( \2674 , \2666 , \2673 );
xor \U$2543 ( \2675 , \2657 , \2674 );
and \U$2544 ( \2676 , \197 , \1086 );
and \U$2545 ( \2677 , \178 , \508 );
nor \U$2546 ( \2678 , \2676 , \2677 );
xnor \U$2547 ( \2679 , \2678 , \487 );
and \U$2548 ( \2680 , \217 , \1301 );
and \U$2549 ( \2681 , \189 , \1246 );
nor \U$2550 ( \2682 , \2680 , \2681 );
xnor \U$2551 ( \2683 , \2682 , \1205 );
xor \U$2552 ( \2684 , \2679 , \2683 );
and \U$2553 ( \2685 , \232 , \1578 );
and \U$2554 ( \2686 , \209 , \1431 );
nor \U$2555 ( \2687 , \2685 , \2686 );
xnor \U$2556 ( \2688 , \2687 , \1436 );
xor \U$2557 ( \2689 , \2684 , \2688 );
and \U$2558 ( \2690 , \247 , \1824 );
and \U$2559 ( \2691 , \224 , \1739 );
nor \U$2560 ( \2692 , \2690 , \2691 );
xnor \U$2561 ( \2693 , \2692 , \1697 );
and \U$2562 ( \2694 , \143 , \2121 );
and \U$2563 ( \2695 , \240 , \2008 );
nor \U$2564 ( \2696 , \2694 , \2695 );
xnor \U$2565 ( \2697 , \2696 , \1961 );
xor \U$2566 ( \2698 , \2693 , \2697 );
and \U$2567 ( \2699 , \158 , \2400 );
and \U$2568 ( \2700 , \134 , \2246 );
nor \U$2569 ( \2701 , \2699 , \2700 );
xnor \U$2570 ( \2702 , \2701 , \2195 );
xor \U$2571 ( \2703 , \2698 , \2702 );
xor \U$2572 ( \2704 , \2689 , \2703 );
and \U$2573 ( \2705 , \474 , \156 );
and \U$2574 ( \2706 , \1147 , \154 );
nor \U$2575 ( \2707 , \2705 , \2706 );
xnor \U$2576 ( \2708 , \2707 , \163 );
and \U$2577 ( \2709 , \307 , \296 );
and \U$2578 ( \2710 , \412 , \168 );
nor \U$2579 ( \2711 , \2709 , \2710 );
xnor \U$2580 ( \2712 , \2711 , \173 );
xor \U$2581 ( \2713 , \2708 , \2712 );
and \U$2582 ( \2714 , \185 , \438 );
and \U$2583 ( \2715 , \261 , \336 );
nor \U$2584 ( \2716 , \2714 , \2715 );
xnor \U$2585 ( \2717 , \2716 , \320 );
xor \U$2586 ( \2718 , \2713 , \2717 );
xor \U$2587 ( \2719 , \2704 , \2718 );
xor \U$2588 ( \2720 , \2675 , \2719 );
xor \U$2589 ( \2721 , \2643 , \2720 );
xor \U$2590 ( \2722 , \2634 , \2721 );
and \U$2591 ( \2723 , \2600 , \2604 );
and \U$2592 ( \2724 , \2604 , \2609 );
and \U$2593 ( \2725 , \2600 , \2609 );
or \U$2594 ( \2726 , \2723 , \2724 , \2725 );
and \U$2595 ( \2727 , \2480 , \2484 );
and \U$2596 ( \2728 , \2484 , \2489 );
and \U$2597 ( \2729 , \2480 , \2489 );
or \U$2598 ( \2730 , \2727 , \2728 , \2729 );
xor \U$2599 ( \2731 , \2726 , \2730 );
and \U$2600 ( \2732 , \2540 , \2554 );
and \U$2601 ( \2733 , \2554 , \2569 );
and \U$2602 ( \2734 , \2540 , \2569 );
or \U$2603 ( \2735 , \2732 , \2733 , \2734 );
xor \U$2604 ( \2736 , \2731 , \2735 );
and \U$2605 ( \2737 , \2504 , \2518 );
and \U$2606 ( \2738 , \2518 , \2535 );
and \U$2607 ( \2739 , \2504 , \2535 );
or \U$2608 ( \2740 , \2737 , \2738 , \2739 );
and \U$2609 ( \2741 , \1684 , \230 );
and \U$2610 ( \2742 , \1802 , \228 );
nor \U$2611 ( \2743 , \2741 , \2742 );
xnor \U$2612 ( \2744 , \2743 , \237 );
and \U$2613 ( \2745 , \1484 , \245 );
and \U$2614 ( \2746 , \1601 , \243 );
nor \U$2615 ( \2747 , \2745 , \2746 );
xnor \U$2616 ( \2748 , \2747 , \252 );
xor \U$2617 ( \2749 , \2744 , \2748 );
and \U$2618 ( \2750 , \1192 , \141 );
and \U$2619 ( \2751 , \1333 , \139 );
nor \U$2620 ( \2752 , \2750 , \2751 );
xnor \U$2621 ( \2753 , \2752 , \148 );
xor \U$2622 ( \2754 , \2749 , \2753 );
xor \U$2623 ( \2755 , \2740 , \2754 );
and \U$2624 ( \2756 , \2521 , \183 );
buf \U$2625 ( \2757 , RIb55e2c0_97);
and \U$2626 ( \2758 , \2757 , \180 );
nor \U$2627 ( \2759 , \2756 , \2758 );
xnor \U$2628 ( \2760 , \2759 , \179 );
and \U$2629 ( \2761 , \2182 , \195 );
and \U$2630 ( \2762 , \2366 , \193 );
nor \U$2631 ( \2763 , \2761 , \2762 );
xnor \U$2632 ( \2764 , \2763 , \202 );
xor \U$2633 ( \2765 , \2760 , \2764 );
and \U$2634 ( \2766 , \1948 , \215 );
and \U$2635 ( \2767 , \2090 , \213 );
nor \U$2636 ( \2768 , \2766 , \2767 );
xnor \U$2637 ( \2769 , \2768 , \222 );
xor \U$2638 ( \2770 , \2765 , \2769 );
xor \U$2639 ( \2771 , \2755 , \2770 );
xor \U$2640 ( \2772 , \2736 , \2771 );
xor \U$2641 ( \2773 , \2722 , \2772 );
xor \U$2642 ( \2774 , \2630 , \2773 );
and \U$2643 ( \2775 , \2470 , \2572 );
and \U$2644 ( \2776 , \2572 , \2612 );
and \U$2645 ( \2777 , \2470 , \2612 );
or \U$2646 ( \2778 , \2775 , \2776 , \2777 );
xor \U$2647 ( \2779 , \2774 , \2778 );
and \U$2648 ( \2780 , \2613 , \2617 );
and \U$2649 ( \2781 , \2618 , \2621 );
or \U$2650 ( \2782 , \2780 , \2781 );
xor \U$2651 ( \2783 , \2779 , \2782 );
buf \U$2652 ( \2784 , \2783 );
buf \U$2653 ( \2785 , \2784 );
and \U$2654 ( \2786 , \2634 , \2721 );
and \U$2655 ( \2787 , \2721 , \2772 );
and \U$2656 ( \2788 , \2634 , \2772 );
or \U$2657 ( \2789 , \2786 , \2787 , \2788 );
and \U$2658 ( \2790 , \2726 , \2730 );
and \U$2659 ( \2791 , \2730 , \2735 );
and \U$2660 ( \2792 , \2726 , \2735 );
or \U$2661 ( \2793 , \2790 , \2791 , \2792 );
and \U$2662 ( \2794 , \2740 , \2754 );
and \U$2663 ( \2795 , \2754 , \2770 );
and \U$2664 ( \2796 , \2740 , \2770 );
or \U$2665 ( \2797 , \2794 , \2795 , \2796 );
xor \U$2666 ( \2798 , \2793 , \2797 );
and \U$2667 ( \2799 , \2657 , \2674 );
and \U$2668 ( \2800 , \2674 , \2719 );
and \U$2669 ( \2801 , \2657 , \2719 );
or \U$2670 ( \2802 , \2799 , \2800 , \2801 );
xor \U$2671 ( \2803 , \2798 , \2802 );
xor \U$2672 ( \2804 , \2789 , \2803 );
and \U$2673 ( \2805 , \2638 , \2642 );
and \U$2674 ( \2806 , \2642 , \2720 );
and \U$2675 ( \2807 , \2638 , \2720 );
or \U$2676 ( \2808 , \2805 , \2806 , \2807 );
and \U$2677 ( \2809 , \2736 , \2771 );
xor \U$2678 ( \2810 , \2808 , \2809 );
and \U$2679 ( \2811 , \2647 , \2651 );
and \U$2680 ( \2812 , \2651 , \2656 );
and \U$2681 ( \2813 , \2647 , \2656 );
or \U$2682 ( \2814 , \2811 , \2812 , \2813 );
and \U$2683 ( \2815 , \2661 , \2665 );
and \U$2684 ( \2816 , \2665 , \2673 );
and \U$2685 ( \2817 , \2661 , \2673 );
or \U$2686 ( \2818 , \2815 , \2816 , \2817 );
xor \U$2687 ( \2819 , \2814 , \2818 );
and \U$2688 ( \2820 , \2689 , \2703 );
and \U$2689 ( \2821 , \2703 , \2718 );
and \U$2690 ( \2822 , \2689 , \2718 );
or \U$2691 ( \2823 , \2820 , \2821 , \2822 );
xor \U$2692 ( \2824 , \2819 , \2823 );
and \U$2693 ( \2825 , \2757 , \183 );
buf \U$2694 ( \2826 , RIb55e338_96);
and \U$2695 ( \2827 , \2826 , \180 );
nor \U$2696 ( \2828 , \2825 , \2827 );
xnor \U$2697 ( \2829 , \2828 , \179 );
and \U$2698 ( \2830 , \2366 , \195 );
and \U$2699 ( \2831 , \2521 , \193 );
nor \U$2700 ( \2832 , \2830 , \2831 );
xnor \U$2701 ( \2833 , \2832 , \202 );
xor \U$2702 ( \2834 , \2829 , \2833 );
buf \U$2703 ( \2835 , RIb5601b0_31);
buf \U$2704 ( \2836 , RIb560138_32);
and \U$2705 ( \2837 , \2836 , \2530 );
not \U$2706 ( \2838 , \2837 );
and \U$2707 ( \2839 , \2835 , \2838 );
xor \U$2708 ( \2840 , \2834 , \2839 );
and \U$2709 ( \2841 , \2090 , \215 );
and \U$2710 ( \2842 , \2182 , \213 );
nor \U$2711 ( \2843 , \2841 , \2842 );
xnor \U$2712 ( \2844 , \2843 , \222 );
and \U$2713 ( \2845 , \1802 , \230 );
and \U$2714 ( \2846 , \1948 , \228 );
nor \U$2715 ( \2847 , \2845 , \2846 );
xnor \U$2716 ( \2848 , \2847 , \237 );
xor \U$2717 ( \2849 , \2844 , \2848 );
and \U$2718 ( \2850 , \1601 , \245 );
and \U$2719 ( \2851 , \1684 , \243 );
nor \U$2720 ( \2852 , \2850 , \2851 );
xnor \U$2721 ( \2853 , \2852 , \252 );
xor \U$2722 ( \2854 , \2849 , \2853 );
xor \U$2723 ( \2855 , \2840 , \2854 );
and \U$2724 ( \2856 , \209 , \1578 );
and \U$2725 ( \2857 , \217 , \1431 );
nor \U$2726 ( \2858 , \2856 , \2857 );
xnor \U$2727 ( \2859 , \2858 , \1436 );
and \U$2728 ( \2860 , \224 , \1824 );
and \U$2729 ( \2861 , \232 , \1739 );
nor \U$2730 ( \2862 , \2860 , \2861 );
xnor \U$2731 ( \2863 , \2862 , \1697 );
xor \U$2732 ( \2864 , \2859 , \2863 );
and \U$2733 ( \2865 , \240 , \2121 );
and \U$2734 ( \2866 , \247 , \2008 );
nor \U$2735 ( \2867 , \2865 , \2866 );
xnor \U$2736 ( \2868 , \2867 , \1961 );
xor \U$2737 ( \2869 , \2864 , \2868 );
and \U$2738 ( \2870 , \1333 , \141 );
and \U$2739 ( \2871 , \1484 , \139 );
nor \U$2740 ( \2872 , \2870 , \2871 );
xnor \U$2741 ( \2873 , \2872 , \148 );
and \U$2742 ( \2874 , \1147 , \156 );
and \U$2743 ( \2875 , \1192 , \154 );
nor \U$2744 ( \2876 , \2874 , \2875 );
xnor \U$2745 ( \2877 , \2876 , \163 );
xor \U$2746 ( \2878 , \2873 , \2877 );
and \U$2747 ( \2879 , \412 , \296 );
and \U$2748 ( \2880 , \474 , \168 );
nor \U$2749 ( \2881 , \2879 , \2880 );
xnor \U$2750 ( \2882 , \2881 , \173 );
xor \U$2751 ( \2883 , \2878 , \2882 );
xor \U$2752 ( \2884 , \2869 , \2883 );
and \U$2753 ( \2885 , \261 , \438 );
and \U$2754 ( \2886 , \307 , \336 );
nor \U$2755 ( \2887 , \2885 , \2886 );
xnor \U$2756 ( \2888 , \2887 , \320 );
and \U$2757 ( \2889 , \178 , \1086 );
and \U$2758 ( \2890 , \185 , \508 );
nor \U$2759 ( \2891 , \2889 , \2890 );
xnor \U$2760 ( \2892 , \2891 , \487 );
xor \U$2761 ( \2893 , \2888 , \2892 );
and \U$2762 ( \2894 , \189 , \1301 );
and \U$2763 ( \2895 , \197 , \1246 );
nor \U$2764 ( \2896 , \2894 , \2895 );
xnor \U$2765 ( \2897 , \2896 , \1205 );
xor \U$2766 ( \2898 , \2893 , \2897 );
xor \U$2767 ( \2899 , \2884 , \2898 );
xor \U$2768 ( \2900 , \2855 , \2899 );
xor \U$2769 ( \2901 , \2824 , \2900 );
and \U$2770 ( \2902 , \2744 , \2748 );
and \U$2771 ( \2903 , \2748 , \2753 );
and \U$2772 ( \2904 , \2744 , \2753 );
or \U$2773 ( \2905 , \2902 , \2903 , \2904 );
and \U$2774 ( \2906 , \2760 , \2764 );
and \U$2775 ( \2907 , \2764 , \2769 );
and \U$2776 ( \2908 , \2760 , \2769 );
or \U$2777 ( \2909 , \2906 , \2907 , \2908 );
xor \U$2778 ( \2910 , \2905 , \2909 );
and \U$2779 ( \2911 , \2708 , \2712 );
and \U$2780 ( \2912 , \2712 , \2717 );
and \U$2781 ( \2913 , \2708 , \2717 );
or \U$2782 ( \2914 , \2911 , \2912 , \2913 );
xor \U$2783 ( \2915 , \2910 , \2914 );
and \U$2784 ( \2916 , \2679 , \2683 );
and \U$2785 ( \2917 , \2683 , \2688 );
and \U$2786 ( \2918 , \2679 , \2688 );
or \U$2787 ( \2919 , \2916 , \2917 , \2918 );
and \U$2788 ( \2920 , \2693 , \2697 );
and \U$2789 ( \2921 , \2697 , \2702 );
and \U$2790 ( \2922 , \2693 , \2702 );
or \U$2791 ( \2923 , \2920 , \2921 , \2922 );
xor \U$2792 ( \2924 , \2919 , \2923 );
and \U$2793 ( \2925 , \134 , \2400 );
and \U$2794 ( \2926 , \143 , \2246 );
nor \U$2795 ( \2927 , \2925 , \2926 );
xnor \U$2796 ( \2928 , \2927 , \2195 );
and \U$2797 ( \2929 , \150 , \2669 );
and \U$2798 ( \2930 , \158 , \2538 );
nor \U$2799 ( \2931 , \2929 , \2930 );
xnor \U$2800 ( \2932 , \2931 , \2534 );
xor \U$2801 ( \2933 , \2928 , \2932 );
xor \U$2802 ( \2934 , \2836 , \2530 );
nand \U$2803 ( \2935 , \166 , \2934 );
xnor \U$2804 ( \2936 , \2935 , \2839 );
xor \U$2805 ( \2937 , \2933 , \2936 );
xor \U$2806 ( \2938 , \2924 , \2937 );
xor \U$2807 ( \2939 , \2915 , \2938 );
xor \U$2808 ( \2940 , \2901 , \2939 );
xor \U$2809 ( \2941 , \2810 , \2940 );
xor \U$2810 ( \2942 , \2804 , \2941 );
and \U$2811 ( \2943 , \2628 , \2629 );
and \U$2812 ( \2944 , \2629 , \2773 );
and \U$2813 ( \2945 , \2628 , \2773 );
or \U$2814 ( \2946 , \2943 , \2944 , \2945 );
xor \U$2815 ( \2947 , \2942 , \2946 );
and \U$2816 ( \2948 , \2774 , \2778 );
and \U$2817 ( \2949 , \2779 , \2782 );
or \U$2818 ( \2950 , \2948 , \2949 );
xor \U$2819 ( \2951 , \2947 , \2950 );
buf \U$2820 ( \2952 , \2951 );
buf \U$2821 ( \2953 , \2952 );
and \U$2822 ( \2954 , \2808 , \2809 );
and \U$2823 ( \2955 , \2809 , \2940 );
and \U$2824 ( \2956 , \2808 , \2940 );
or \U$2825 ( \2957 , \2954 , \2955 , \2956 );
and \U$2826 ( \2958 , \2814 , \2818 );
and \U$2827 ( \2959 , \2818 , \2823 );
and \U$2828 ( \2960 , \2814 , \2823 );
or \U$2829 ( \2961 , \2958 , \2959 , \2960 );
and \U$2830 ( \2962 , \2840 , \2854 );
and \U$2831 ( \2963 , \2854 , \2899 );
and \U$2832 ( \2964 , \2840 , \2899 );
or \U$2833 ( \2965 , \2962 , \2963 , \2964 );
xor \U$2834 ( \2966 , \2961 , \2965 );
and \U$2835 ( \2967 , \2915 , \2938 );
xor \U$2836 ( \2968 , \2966 , \2967 );
xor \U$2837 ( \2969 , \2957 , \2968 );
and \U$2838 ( \2970 , \2793 , \2797 );
and \U$2839 ( \2971 , \2797 , \2802 );
and \U$2840 ( \2972 , \2793 , \2802 );
or \U$2841 ( \2973 , \2970 , \2971 , \2972 );
and \U$2842 ( \2974 , \2824 , \2900 );
and \U$2843 ( \2975 , \2900 , \2939 );
and \U$2844 ( \2976 , \2824 , \2939 );
or \U$2845 ( \2977 , \2974 , \2975 , \2976 );
xor \U$2846 ( \2978 , \2973 , \2977 );
and \U$2847 ( \2979 , \2873 , \2877 );
and \U$2848 ( \2980 , \2877 , \2882 );
and \U$2849 ( \2981 , \2873 , \2882 );
or \U$2850 ( \2982 , \2979 , \2980 , \2981 );
and \U$2851 ( \2983 , \2829 , \2833 );
and \U$2852 ( \2984 , \2833 , \2839 );
and \U$2853 ( \2985 , \2829 , \2839 );
or \U$2854 ( \2986 , \2983 , \2984 , \2985 );
xor \U$2855 ( \2987 , \2982 , \2986 );
and \U$2856 ( \2988 , \2844 , \2848 );
and \U$2857 ( \2989 , \2848 , \2853 );
and \U$2858 ( \2990 , \2844 , \2853 );
or \U$2859 ( \2991 , \2988 , \2989 , \2990 );
xor \U$2860 ( \2992 , \2987 , \2991 );
and \U$2861 ( \2993 , \2905 , \2909 );
and \U$2862 ( \2994 , \2909 , \2914 );
and \U$2863 ( \2995 , \2905 , \2914 );
or \U$2864 ( \2996 , \2993 , \2994 , \2995 );
and \U$2865 ( \2997 , \2869 , \2883 );
and \U$2866 ( \2998 , \2883 , \2898 );
and \U$2867 ( \2999 , \2869 , \2898 );
or \U$2868 ( \3000 , \2997 , \2998 , \2999 );
xor \U$2869 ( \3001 , \2996 , \3000 );
and \U$2870 ( \3002 , \2919 , \2923 );
and \U$2871 ( \3003 , \2923 , \2937 );
and \U$2872 ( \3004 , \2919 , \2937 );
or \U$2873 ( \3005 , \3002 , \3003 , \3004 );
xor \U$2874 ( \3006 , \3001 , \3005 );
xor \U$2875 ( \3007 , \2992 , \3006 );
and \U$2876 ( \3008 , \2859 , \2863 );
and \U$2877 ( \3009 , \2863 , \2868 );
and \U$2878 ( \3010 , \2859 , \2868 );
or \U$2879 ( \3011 , \3008 , \3009 , \3010 );
and \U$2880 ( \3012 , \2928 , \2932 );
and \U$2881 ( \3013 , \2932 , \2936 );
and \U$2882 ( \3014 , \2928 , \2936 );
or \U$2883 ( \3015 , \3012 , \3013 , \3014 );
xor \U$2884 ( \3016 , \3011 , \3015 );
and \U$2885 ( \3017 , \2888 , \2892 );
and \U$2886 ( \3018 , \2892 , \2897 );
and \U$2887 ( \3019 , \2888 , \2897 );
or \U$2888 ( \3020 , \3017 , \3018 , \3019 );
xor \U$2889 ( \3021 , \3016 , \3020 );
and \U$2890 ( \3022 , \1192 , \156 );
and \U$2891 ( \3023 , \1333 , \154 );
nor \U$2892 ( \3024 , \3022 , \3023 );
xnor \U$2893 ( \3025 , \3024 , \163 );
and \U$2894 ( \3026 , \474 , \296 );
and \U$2895 ( \3027 , \1147 , \168 );
nor \U$2896 ( \3028 , \3026 , \3027 );
xnor \U$2897 ( \3029 , \3028 , \173 );
xor \U$2898 ( \3030 , \3025 , \3029 );
and \U$2899 ( \3031 , \307 , \438 );
and \U$2900 ( \3032 , \412 , \336 );
nor \U$2901 ( \3033 , \3031 , \3032 );
xnor \U$2902 ( \3034 , \3033 , \320 );
xor \U$2903 ( \3035 , \3030 , \3034 );
and \U$2904 ( \3036 , \2826 , \183 );
buf \U$2905 ( \3037 , RIb55e3b0_95);
and \U$2906 ( \3038 , \3037 , \180 );
nor \U$2907 ( \3039 , \3036 , \3038 );
xnor \U$2908 ( \3040 , \3039 , \179 );
and \U$2909 ( \3041 , \2521 , \195 );
and \U$2910 ( \3042 , \2757 , \193 );
nor \U$2911 ( \3043 , \3041 , \3042 );
xnor \U$2912 ( \3044 , \3043 , \202 );
xor \U$2913 ( \3045 , \3040 , \3044 );
and \U$2914 ( \3046 , \2182 , \215 );
and \U$2915 ( \3047 , \2366 , \213 );
nor \U$2916 ( \3048 , \3046 , \3047 );
xnor \U$2917 ( \3049 , \3048 , \222 );
xor \U$2918 ( \3050 , \3045 , \3049 );
xor \U$2919 ( \3051 , \3035 , \3050 );
and \U$2920 ( \3052 , \1948 , \230 );
and \U$2921 ( \3053 , \2090 , \228 );
nor \U$2922 ( \3054 , \3052 , \3053 );
xnor \U$2923 ( \3055 , \3054 , \237 );
and \U$2924 ( \3056 , \1684 , \245 );
and \U$2925 ( \3057 , \1802 , \243 );
nor \U$2926 ( \3058 , \3056 , \3057 );
xnor \U$2927 ( \3059 , \3058 , \252 );
xor \U$2928 ( \3060 , \3055 , \3059 );
and \U$2929 ( \3061 , \1484 , \141 );
and \U$2930 ( \3062 , \1601 , \139 );
nor \U$2931 ( \3063 , \3061 , \3062 );
xnor \U$2932 ( \3064 , \3063 , \148 );
xor \U$2933 ( \3065 , \3060 , \3064 );
xor \U$2934 ( \3066 , \3051 , \3065 );
xor \U$2935 ( \3067 , \3021 , \3066 );
and \U$2936 ( \3068 , \232 , \1824 );
and \U$2937 ( \3069 , \209 , \1739 );
nor \U$2938 ( \3070 , \3068 , \3069 );
xnor \U$2939 ( \3071 , \3070 , \1697 );
and \U$2940 ( \3072 , \247 , \2121 );
and \U$2941 ( \3073 , \224 , \2008 );
nor \U$2942 ( \3074 , \3072 , \3073 );
xnor \U$2943 ( \3075 , \3074 , \1961 );
xor \U$2944 ( \3076 , \3071 , \3075 );
and \U$2945 ( \3077 , \143 , \2400 );
and \U$2946 ( \3078 , \240 , \2246 );
nor \U$2947 ( \3079 , \3077 , \3078 );
xnor \U$2948 ( \3080 , \3079 , \2195 );
xor \U$2949 ( \3081 , \3076 , \3080 );
and \U$2950 ( \3082 , \185 , \1086 );
and \U$2951 ( \3083 , \261 , \508 );
nor \U$2952 ( \3084 , \3082 , \3083 );
xnor \U$2953 ( \3085 , \3084 , \487 );
and \U$2954 ( \3086 , \197 , \1301 );
and \U$2955 ( \3087 , \178 , \1246 );
nor \U$2956 ( \3088 , \3086 , \3087 );
xnor \U$2957 ( \3089 , \3088 , \1205 );
xor \U$2958 ( \3090 , \3085 , \3089 );
and \U$2959 ( \3091 , \217 , \1578 );
and \U$2960 ( \3092 , \189 , \1431 );
nor \U$2961 ( \3093 , \3091 , \3092 );
xnor \U$2962 ( \3094 , \3093 , \1436 );
xor \U$2963 ( \3095 , \3090 , \3094 );
xor \U$2964 ( \3096 , \3081 , \3095 );
and \U$2965 ( \3097 , \158 , \2669 );
and \U$2966 ( \3098 , \134 , \2538 );
nor \U$2967 ( \3099 , \3097 , \3098 );
xnor \U$2968 ( \3100 , \3099 , \2534 );
xor \U$2969 ( \3101 , \2835 , \2836 );
not \U$2970 ( \3102 , \2934 );
and \U$2971 ( \3103 , \3101 , \3102 );
and \U$2972 ( \3104 , \166 , \3103 );
and \U$2973 ( \3105 , \150 , \2934 );
nor \U$2974 ( \3106 , \3104 , \3105 );
xnor \U$2975 ( \3107 , \3106 , \2839 );
xor \U$2976 ( \3108 , \3100 , \3107 );
xor \U$2977 ( \3109 , \3096 , \3108 );
xor \U$2978 ( \3110 , \3067 , \3109 );
xor \U$2979 ( \3111 , \3007 , \3110 );
xor \U$2980 ( \3112 , \2978 , \3111 );
xor \U$2981 ( \3113 , \2969 , \3112 );
and \U$2982 ( \3114 , \2789 , \2803 );
and \U$2983 ( \3115 , \2803 , \2941 );
and \U$2984 ( \3116 , \2789 , \2941 );
or \U$2985 ( \3117 , \3114 , \3115 , \3116 );
xor \U$2986 ( \3118 , \3113 , \3117 );
and \U$2987 ( \3119 , \2942 , \2946 );
and \U$2988 ( \3120 , \2947 , \2950 );
or \U$2989 ( \3121 , \3119 , \3120 );
xor \U$2990 ( \3122 , \3118 , \3121 );
buf \U$2991 ( \3123 , \3122 );
buf \U$2992 ( \3124 , \3123 );
and \U$2993 ( \3125 , \2973 , \2977 );
and \U$2994 ( \3126 , \2977 , \3111 );
and \U$2995 ( \3127 , \2973 , \3111 );
or \U$2996 ( \3128 , \3125 , \3126 , \3127 );
and \U$2997 ( \3129 , \2961 , \2965 );
and \U$2998 ( \3130 , \2965 , \2967 );
and \U$2999 ( \3131 , \2961 , \2967 );
or \U$3000 ( \3132 , \3129 , \3130 , \3131 );
and \U$3001 ( \3133 , \2992 , \3006 );
and \U$3002 ( \3134 , \3006 , \3110 );
and \U$3003 ( \3135 , \2992 , \3110 );
or \U$3004 ( \3136 , \3133 , \3134 , \3135 );
xor \U$3005 ( \3137 , \3132 , \3136 );
and \U$3006 ( \3138 , \3035 , \3050 );
and \U$3007 ( \3139 , \3050 , \3065 );
and \U$3008 ( \3140 , \3035 , \3065 );
or \U$3009 ( \3141 , \3138 , \3139 , \3140 );
and \U$3010 ( \3142 , \3037 , \183 );
buf \U$3011 ( \3143 , RIb55e428_94);
and \U$3012 ( \3144 , \3143 , \180 );
nor \U$3013 ( \3145 , \3142 , \3144 );
xnor \U$3014 ( \3146 , \3145 , \179 );
and \U$3015 ( \3147 , \2757 , \195 );
and \U$3016 ( \3148 , \2826 , \193 );
nor \U$3017 ( \3149 , \3147 , \3148 );
xnor \U$3018 ( \3150 , \3149 , \202 );
xor \U$3019 ( \3151 , \3146 , \3150 );
buf \U$3020 ( \3152 , RIb5602a0_29);
buf \U$3021 ( \3153 , RIb560228_30);
and \U$3022 ( \3154 , \3153 , \2835 );
not \U$3023 ( \3155 , \3154 );
and \U$3024 ( \3156 , \3152 , \3155 );
xor \U$3025 ( \3157 , \3151 , \3156 );
xor \U$3026 ( \3158 , \3141 , \3157 );
and \U$3027 ( \3159 , \2366 , \215 );
and \U$3028 ( \3160 , \2521 , \213 );
nor \U$3029 ( \3161 , \3159 , \3160 );
xnor \U$3030 ( \3162 , \3161 , \222 );
and \U$3031 ( \3163 , \2090 , \230 );
and \U$3032 ( \3164 , \2182 , \228 );
nor \U$3033 ( \3165 , \3163 , \3164 );
xnor \U$3034 ( \3166 , \3165 , \237 );
xor \U$3035 ( \3167 , \3162 , \3166 );
and \U$3036 ( \3168 , \1802 , \245 );
and \U$3037 ( \3169 , \1948 , \243 );
nor \U$3038 ( \3170 , \3168 , \3169 );
xnor \U$3039 ( \3171 , \3170 , \252 );
xor \U$3040 ( \3172 , \3167 , \3171 );
and \U$3041 ( \3173 , \412 , \438 );
and \U$3042 ( \3174 , \474 , \336 );
nor \U$3043 ( \3175 , \3173 , \3174 );
xnor \U$3044 ( \3176 , \3175 , \320 );
and \U$3045 ( \3177 , \261 , \1086 );
and \U$3046 ( \3178 , \307 , \508 );
nor \U$3047 ( \3179 , \3177 , \3178 );
xnor \U$3048 ( \3180 , \3179 , \487 );
xor \U$3049 ( \3181 , \3176 , \3180 );
and \U$3050 ( \3182 , \178 , \1301 );
and \U$3051 ( \3183 , \185 , \1246 );
nor \U$3052 ( \3184 , \3182 , \3183 );
xnor \U$3053 ( \3185 , \3184 , \1205 );
xor \U$3054 ( \3186 , \3181 , \3185 );
xor \U$3055 ( \3187 , \3172 , \3186 );
and \U$3056 ( \3188 , \1601 , \141 );
and \U$3057 ( \3189 , \1684 , \139 );
nor \U$3058 ( \3190 , \3188 , \3189 );
xnor \U$3059 ( \3191 , \3190 , \148 );
and \U$3060 ( \3192 , \1333 , \156 );
and \U$3061 ( \3193 , \1484 , \154 );
nor \U$3062 ( \3194 , \3192 , \3193 );
xnor \U$3063 ( \3195 , \3194 , \163 );
xor \U$3064 ( \3196 , \3191 , \3195 );
and \U$3065 ( \3197 , \1147 , \296 );
and \U$3066 ( \3198 , \1192 , \168 );
nor \U$3067 ( \3199 , \3197 , \3198 );
xnor \U$3068 ( \3200 , \3199 , \173 );
xor \U$3069 ( \3201 , \3196 , \3200 );
xor \U$3070 ( \3202 , \3187 , \3201 );
xor \U$3071 ( \3203 , \3158 , \3202 );
xor \U$3072 ( \3204 , \3137 , \3203 );
xor \U$3073 ( \3205 , \3128 , \3204 );
and \U$3074 ( \3206 , \3011 , \3015 );
and \U$3075 ( \3207 , \3015 , \3020 );
and \U$3076 ( \3208 , \3011 , \3020 );
or \U$3077 ( \3209 , \3206 , \3207 , \3208 );
and \U$3078 ( \3210 , \2982 , \2986 );
and \U$3079 ( \3211 , \2986 , \2991 );
and \U$3080 ( \3212 , \2982 , \2991 );
or \U$3081 ( \3213 , \3210 , \3211 , \3212 );
xor \U$3082 ( \3214 , \3209 , \3213 );
and \U$3083 ( \3215 , \3081 , \3095 );
and \U$3084 ( \3216 , \3095 , \3108 );
and \U$3085 ( \3217 , \3081 , \3108 );
or \U$3086 ( \3218 , \3215 , \3216 , \3217 );
xor \U$3087 ( \3219 , \3214 , \3218 );
and \U$3088 ( \3220 , \2996 , \3000 );
and \U$3089 ( \3221 , \3000 , \3005 );
and \U$3090 ( \3222 , \2996 , \3005 );
or \U$3091 ( \3223 , \3220 , \3221 , \3222 );
and \U$3092 ( \3224 , \3021 , \3066 );
and \U$3093 ( \3225 , \3066 , \3109 );
and \U$3094 ( \3226 , \3021 , \3109 );
or \U$3095 ( \3227 , \3224 , \3225 , \3226 );
xor \U$3096 ( \3228 , \3223 , \3227 );
and \U$3097 ( \3229 , \3025 , \3029 );
and \U$3098 ( \3230 , \3029 , \3034 );
and \U$3099 ( \3231 , \3025 , \3034 );
or \U$3100 ( \3232 , \3229 , \3230 , \3231 );
and \U$3101 ( \3233 , \3040 , \3044 );
and \U$3102 ( \3234 , \3044 , \3049 );
and \U$3103 ( \3235 , \3040 , \3049 );
or \U$3104 ( \3236 , \3233 , \3234 , \3235 );
xor \U$3105 ( \3237 , \3232 , \3236 );
and \U$3106 ( \3238 , \3055 , \3059 );
and \U$3107 ( \3239 , \3059 , \3064 );
and \U$3108 ( \3240 , \3055 , \3064 );
or \U$3109 ( \3241 , \3238 , \3239 , \3240 );
xor \U$3110 ( \3242 , \3237 , \3241 );
and \U$3111 ( \3243 , \3071 , \3075 );
and \U$3112 ( \3244 , \3075 , \3080 );
and \U$3113 ( \3245 , \3071 , \3080 );
or \U$3114 ( \3246 , \3243 , \3244 , \3245 );
and \U$3115 ( \3247 , \3085 , \3089 );
and \U$3116 ( \3248 , \3089 , \3094 );
and \U$3117 ( \3249 , \3085 , \3094 );
or \U$3118 ( \3250 , \3247 , \3248 , \3249 );
xor \U$3119 ( \3251 , \3246 , \3250 );
and \U$3120 ( \3252 , \3100 , \3107 );
xor \U$3121 ( \3253 , \3251 , \3252 );
xor \U$3122 ( \3254 , \3242 , \3253 );
xor \U$3123 ( \3255 , \3153 , \2835 );
nand \U$3124 ( \3256 , \166 , \3255 );
xnor \U$3125 ( \3257 , \3256 , \3156 );
and \U$3126 ( \3258 , \189 , \1578 );
and \U$3127 ( \3259 , \197 , \1431 );
nor \U$3128 ( \3260 , \3258 , \3259 );
xnor \U$3129 ( \3261 , \3260 , \1436 );
and \U$3130 ( \3262 , \209 , \1824 );
and \U$3131 ( \3263 , \217 , \1739 );
nor \U$3132 ( \3264 , \3262 , \3263 );
xnor \U$3133 ( \3265 , \3264 , \1697 );
xor \U$3134 ( \3266 , \3261 , \3265 );
and \U$3135 ( \3267 , \224 , \2121 );
and \U$3136 ( \3268 , \232 , \2008 );
nor \U$3137 ( \3269 , \3267 , \3268 );
xnor \U$3138 ( \3270 , \3269 , \1961 );
xor \U$3139 ( \3271 , \3266 , \3270 );
xor \U$3140 ( \3272 , \3257 , \3271 );
and \U$3141 ( \3273 , \240 , \2400 );
and \U$3142 ( \3274 , \247 , \2246 );
nor \U$3143 ( \3275 , \3273 , \3274 );
xnor \U$3144 ( \3276 , \3275 , \2195 );
and \U$3145 ( \3277 , \134 , \2669 );
and \U$3146 ( \3278 , \143 , \2538 );
nor \U$3147 ( \3279 , \3277 , \3278 );
xnor \U$3148 ( \3280 , \3279 , \2534 );
xor \U$3149 ( \3281 , \3276 , \3280 );
and \U$3150 ( \3282 , \150 , \3103 );
and \U$3151 ( \3283 , \158 , \2934 );
nor \U$3152 ( \3284 , \3282 , \3283 );
xnor \U$3153 ( \3285 , \3284 , \2839 );
xor \U$3154 ( \3286 , \3281 , \3285 );
xor \U$3155 ( \3287 , \3272 , \3286 );
xor \U$3156 ( \3288 , \3254 , \3287 );
xor \U$3157 ( \3289 , \3228 , \3288 );
xor \U$3158 ( \3290 , \3219 , \3289 );
xor \U$3159 ( \3291 , \3205 , \3290 );
and \U$3160 ( \3292 , \2957 , \2968 );
and \U$3161 ( \3293 , \2968 , \3112 );
and \U$3162 ( \3294 , \2957 , \3112 );
or \U$3163 ( \3295 , \3292 , \3293 , \3294 );
xor \U$3164 ( \3296 , \3291 , \3295 );
and \U$3165 ( \3297 , \3113 , \3117 );
and \U$3166 ( \3298 , \3118 , \3121 );
or \U$3167 ( \3299 , \3297 , \3298 );
xor \U$3168 ( \3300 , \3296 , \3299 );
buf \U$3169 ( \3301 , \3300 );
buf \U$3170 ( \3302 , \3301 );
and \U$3171 ( \3303 , \3132 , \3136 );
and \U$3172 ( \3304 , \3136 , \3203 );
and \U$3173 ( \3305 , \3132 , \3203 );
or \U$3174 ( \3306 , \3303 , \3304 , \3305 );
and \U$3175 ( \3307 , \3219 , \3289 );
xor \U$3176 ( \3308 , \3306 , \3307 );
and \U$3177 ( \3309 , \3223 , \3227 );
and \U$3178 ( \3310 , \3227 , \3288 );
and \U$3179 ( \3311 , \3223 , \3288 );
or \U$3180 ( \3312 , \3309 , \3310 , \3311 );
and \U$3181 ( \3313 , \3209 , \3213 );
and \U$3182 ( \3314 , \3213 , \3218 );
and \U$3183 ( \3315 , \3209 , \3218 );
or \U$3184 ( \3316 , \3313 , \3314 , \3315 );
and \U$3185 ( \3317 , \3141 , \3157 );
and \U$3186 ( \3318 , \3157 , \3202 );
and \U$3187 ( \3319 , \3141 , \3202 );
or \U$3188 ( \3320 , \3317 , \3318 , \3319 );
xor \U$3189 ( \3321 , \3316 , \3320 );
and \U$3190 ( \3322 , \3242 , \3253 );
and \U$3191 ( \3323 , \3253 , \3287 );
and \U$3192 ( \3324 , \3242 , \3287 );
or \U$3193 ( \3325 , \3322 , \3323 , \3324 );
xor \U$3194 ( \3326 , \3321 , \3325 );
xor \U$3195 ( \3327 , \3312 , \3326 );
and \U$3196 ( \3328 , \3232 , \3236 );
and \U$3197 ( \3329 , \3236 , \3241 );
and \U$3198 ( \3330 , \3232 , \3241 );
or \U$3199 ( \3331 , \3328 , \3329 , \3330 );
and \U$3200 ( \3332 , \3246 , \3250 );
and \U$3201 ( \3333 , \3250 , \3252 );
and \U$3202 ( \3334 , \3246 , \3252 );
or \U$3203 ( \3335 , \3332 , \3333 , \3334 );
xor \U$3204 ( \3336 , \3331 , \3335 );
and \U$3205 ( \3337 , \3257 , \3271 );
and \U$3206 ( \3338 , \3271 , \3286 );
and \U$3207 ( \3339 , \3257 , \3286 );
or \U$3208 ( \3340 , \3337 , \3338 , \3339 );
xor \U$3209 ( \3341 , \3336 , \3340 );
and \U$3210 ( \3342 , \3172 , \3186 );
and \U$3211 ( \3343 , \3186 , \3201 );
and \U$3212 ( \3344 , \3172 , \3201 );
or \U$3213 ( \3345 , \3342 , \3343 , \3344 );
and \U$3214 ( \3346 , \143 , \2669 );
and \U$3215 ( \3347 , \240 , \2538 );
nor \U$3216 ( \3348 , \3346 , \3347 );
xnor \U$3217 ( \3349 , \3348 , \2534 );
and \U$3218 ( \3350 , \158 , \3103 );
and \U$3219 ( \3351 , \134 , \2934 );
nor \U$3220 ( \3352 , \3350 , \3351 );
xnor \U$3221 ( \3353 , \3352 , \2839 );
xor \U$3222 ( \3354 , \3349 , \3353 );
xor \U$3223 ( \3355 , \3152 , \3153 );
not \U$3224 ( \3356 , \3255 );
and \U$3225 ( \3357 , \3355 , \3356 );
and \U$3226 ( \3358 , \166 , \3357 );
and \U$3227 ( \3359 , \150 , \3255 );
nor \U$3228 ( \3360 , \3358 , \3359 );
xnor \U$3229 ( \3361 , \3360 , \3156 );
xor \U$3230 ( \3362 , \3354 , \3361 );
and \U$3231 ( \3363 , \217 , \1824 );
and \U$3232 ( \3364 , \189 , \1739 );
nor \U$3233 ( \3365 , \3363 , \3364 );
xnor \U$3234 ( \3366 , \3365 , \1697 );
and \U$3235 ( \3367 , \232 , \2121 );
and \U$3236 ( \3368 , \209 , \2008 );
nor \U$3237 ( \3369 , \3367 , \3368 );
xnor \U$3238 ( \3370 , \3369 , \1961 );
xor \U$3239 ( \3371 , \3366 , \3370 );
and \U$3240 ( \3372 , \247 , \2400 );
and \U$3241 ( \3373 , \224 , \2246 );
nor \U$3242 ( \3374 , \3372 , \3373 );
xnor \U$3243 ( \3375 , \3374 , \2195 );
xor \U$3244 ( \3376 , \3371 , \3375 );
xor \U$3245 ( \3377 , \3362 , \3376 );
and \U$3246 ( \3378 , \307 , \1086 );
and \U$3247 ( \3379 , \412 , \508 );
nor \U$3248 ( \3380 , \3378 , \3379 );
xnor \U$3249 ( \3381 , \3380 , \487 );
and \U$3250 ( \3382 , \185 , \1301 );
and \U$3251 ( \3383 , \261 , \1246 );
nor \U$3252 ( \3384 , \3382 , \3383 );
xnor \U$3253 ( \3385 , \3384 , \1205 );
xor \U$3254 ( \3386 , \3381 , \3385 );
and \U$3255 ( \3387 , \197 , \1578 );
and \U$3256 ( \3388 , \178 , \1431 );
nor \U$3257 ( \3389 , \3387 , \3388 );
xnor \U$3258 ( \3390 , \3389 , \1436 );
xor \U$3259 ( \3391 , \3386 , \3390 );
xor \U$3260 ( \3392 , \3377 , \3391 );
xor \U$3261 ( \3393 , \3345 , \3392 );
and \U$3262 ( \3394 , \3143 , \183 );
buf \U$3263 ( \3395 , RIb55e4a0_93);
and \U$3264 ( \3396 , \3395 , \180 );
nor \U$3265 ( \3397 , \3394 , \3396 );
xnor \U$3266 ( \3398 , \3397 , \179 );
and \U$3267 ( \3399 , \2826 , \195 );
and \U$3268 ( \3400 , \3037 , \193 );
nor \U$3269 ( \3401 , \3399 , \3400 );
xnor \U$3270 ( \3402 , \3401 , \202 );
xor \U$3271 ( \3403 , \3398 , \3402 );
and \U$3272 ( \3404 , \2521 , \215 );
and \U$3273 ( \3405 , \2757 , \213 );
nor \U$3274 ( \3406 , \3404 , \3405 );
xnor \U$3275 ( \3407 , \3406 , \222 );
xor \U$3276 ( \3408 , \3403 , \3407 );
and \U$3277 ( \3409 , \2182 , \230 );
and \U$3278 ( \3410 , \2366 , \228 );
nor \U$3279 ( \3411 , \3409 , \3410 );
xnor \U$3280 ( \3412 , \3411 , \237 );
and \U$3281 ( \3413 , \1948 , \245 );
and \U$3282 ( \3414 , \2090 , \243 );
nor \U$3283 ( \3415 , \3413 , \3414 );
xnor \U$3284 ( \3416 , \3415 , \252 );
xor \U$3285 ( \3417 , \3412 , \3416 );
and \U$3286 ( \3418 , \1684 , \141 );
and \U$3287 ( \3419 , \1802 , \139 );
nor \U$3288 ( \3420 , \3418 , \3419 );
xnor \U$3289 ( \3421 , \3420 , \148 );
xor \U$3290 ( \3422 , \3417 , \3421 );
xor \U$3291 ( \3423 , \3408 , \3422 );
and \U$3292 ( \3424 , \1484 , \156 );
and \U$3293 ( \3425 , \1601 , \154 );
nor \U$3294 ( \3426 , \3424 , \3425 );
xnor \U$3295 ( \3427 , \3426 , \163 );
and \U$3296 ( \3428 , \1192 , \296 );
and \U$3297 ( \3429 , \1333 , \168 );
nor \U$3298 ( \3430 , \3428 , \3429 );
xnor \U$3299 ( \3431 , \3430 , \173 );
xor \U$3300 ( \3432 , \3427 , \3431 );
and \U$3301 ( \3433 , \474 , \438 );
and \U$3302 ( \3434 , \1147 , \336 );
nor \U$3303 ( \3435 , \3433 , \3434 );
xnor \U$3304 ( \3436 , \3435 , \320 );
xor \U$3305 ( \3437 , \3432 , \3436 );
xor \U$3306 ( \3438 , \3423 , \3437 );
xor \U$3307 ( \3439 , \3393 , \3438 );
xor \U$3308 ( \3440 , \3341 , \3439 );
and \U$3309 ( \3441 , \3146 , \3150 );
and \U$3310 ( \3442 , \3150 , \3156 );
and \U$3311 ( \3443 , \3146 , \3156 );
or \U$3312 ( \3444 , \3441 , \3442 , \3443 );
and \U$3313 ( \3445 , \3162 , \3166 );
and \U$3314 ( \3446 , \3166 , \3171 );
and \U$3315 ( \3447 , \3162 , \3171 );
or \U$3316 ( \3448 , \3445 , \3446 , \3447 );
xor \U$3317 ( \3449 , \3444 , \3448 );
and \U$3318 ( \3450 , \3191 , \3195 );
and \U$3319 ( \3451 , \3195 , \3200 );
and \U$3320 ( \3452 , \3191 , \3200 );
or \U$3321 ( \3453 , \3450 , \3451 , \3452 );
xor \U$3322 ( \3454 , \3449 , \3453 );
and \U$3323 ( \3455 , \3176 , \3180 );
and \U$3324 ( \3456 , \3180 , \3185 );
and \U$3325 ( \3457 , \3176 , \3185 );
or \U$3326 ( \3458 , \3455 , \3456 , \3457 );
and \U$3327 ( \3459 , \3261 , \3265 );
and \U$3328 ( \3460 , \3265 , \3270 );
and \U$3329 ( \3461 , \3261 , \3270 );
or \U$3330 ( \3462 , \3459 , \3460 , \3461 );
xor \U$3331 ( \3463 , \3458 , \3462 );
and \U$3332 ( \3464 , \3276 , \3280 );
and \U$3333 ( \3465 , \3280 , \3285 );
and \U$3334 ( \3466 , \3276 , \3285 );
or \U$3335 ( \3467 , \3464 , \3465 , \3466 );
xor \U$3336 ( \3468 , \3463 , \3467 );
xor \U$3337 ( \3469 , \3454 , \3468 );
xor \U$3338 ( \3470 , \3440 , \3469 );
xor \U$3339 ( \3471 , \3327 , \3470 );
xor \U$3340 ( \3472 , \3308 , \3471 );
and \U$3341 ( \3473 , \3128 , \3204 );
and \U$3342 ( \3474 , \3204 , \3290 );
and \U$3343 ( \3475 , \3128 , \3290 );
or \U$3344 ( \3476 , \3473 , \3474 , \3475 );
xor \U$3345 ( \3477 , \3472 , \3476 );
and \U$3346 ( \3478 , \3291 , \3295 );
and \U$3347 ( \3479 , \3296 , \3299 );
or \U$3348 ( \3480 , \3478 , \3479 );
xor \U$3349 ( \3481 , \3477 , \3480 );
buf \U$3350 ( \3482 , \3481 );
buf \U$3351 ( \3483 , \3482 );
and \U$3352 ( \3484 , \3312 , \3326 );
and \U$3353 ( \3485 , \3326 , \3470 );
and \U$3354 ( \3486 , \3312 , \3470 );
or \U$3355 ( \3487 , \3484 , \3485 , \3486 );
and \U$3356 ( \3488 , \3331 , \3335 );
and \U$3357 ( \3489 , \3335 , \3340 );
and \U$3358 ( \3490 , \3331 , \3340 );
or \U$3359 ( \3491 , \3488 , \3489 , \3490 );
and \U$3360 ( \3492 , \3345 , \3392 );
and \U$3361 ( \3493 , \3392 , \3438 );
and \U$3362 ( \3494 , \3345 , \3438 );
or \U$3363 ( \3495 , \3492 , \3493 , \3494 );
xor \U$3364 ( \3496 , \3491 , \3495 );
and \U$3365 ( \3497 , \3454 , \3468 );
xor \U$3366 ( \3498 , \3496 , \3497 );
xor \U$3367 ( \3499 , \3487 , \3498 );
and \U$3368 ( \3500 , \3316 , \3320 );
and \U$3369 ( \3501 , \3320 , \3325 );
and \U$3370 ( \3502 , \3316 , \3325 );
or \U$3371 ( \3503 , \3500 , \3501 , \3502 );
and \U$3372 ( \3504 , \3341 , \3439 );
and \U$3373 ( \3505 , \3439 , \3469 );
and \U$3374 ( \3506 , \3341 , \3469 );
or \U$3375 ( \3507 , \3504 , \3505 , \3506 );
xor \U$3376 ( \3508 , \3503 , \3507 );
and \U$3377 ( \3509 , \3444 , \3448 );
and \U$3378 ( \3510 , \3448 , \3453 );
and \U$3379 ( \3511 , \3444 , \3453 );
or \U$3380 ( \3512 , \3509 , \3510 , \3511 );
and \U$3381 ( \3513 , \3458 , \3462 );
and \U$3382 ( \3514 , \3462 , \3467 );
and \U$3383 ( \3515 , \3458 , \3467 );
or \U$3384 ( \3516 , \3513 , \3514 , \3515 );
xor \U$3385 ( \3517 , \3512 , \3516 );
and \U$3386 ( \3518 , \3362 , \3376 );
and \U$3387 ( \3519 , \3376 , \3391 );
and \U$3388 ( \3520 , \3362 , \3391 );
or \U$3389 ( \3521 , \3518 , \3519 , \3520 );
xor \U$3390 ( \3522 , \3517 , \3521 );
and \U$3391 ( \3523 , \3398 , \3402 );
and \U$3392 ( \3524 , \3402 , \3407 );
and \U$3393 ( \3525 , \3398 , \3407 );
or \U$3394 ( \3526 , \3523 , \3524 , \3525 );
and \U$3395 ( \3527 , \3412 , \3416 );
and \U$3396 ( \3528 , \3416 , \3421 );
and \U$3397 ( \3529 , \3412 , \3421 );
or \U$3398 ( \3530 , \3527 , \3528 , \3529 );
xor \U$3399 ( \3531 , \3526 , \3530 );
and \U$3400 ( \3532 , \3427 , \3431 );
and \U$3401 ( \3533 , \3431 , \3436 );
and \U$3402 ( \3534 , \3427 , \3436 );
or \U$3403 ( \3535 , \3532 , \3533 , \3534 );
xor \U$3404 ( \3536 , \3531 , \3535 );
and \U$3405 ( \3537 , \3349 , \3353 );
and \U$3406 ( \3538 , \3353 , \3361 );
and \U$3407 ( \3539 , \3349 , \3361 );
or \U$3408 ( \3540 , \3537 , \3538 , \3539 );
and \U$3409 ( \3541 , \3366 , \3370 );
and \U$3410 ( \3542 , \3370 , \3375 );
and \U$3411 ( \3543 , \3366 , \3375 );
or \U$3412 ( \3544 , \3541 , \3542 , \3543 );
xor \U$3413 ( \3545 , \3540 , \3544 );
and \U$3414 ( \3546 , \3381 , \3385 );
and \U$3415 ( \3547 , \3385 , \3390 );
and \U$3416 ( \3548 , \3381 , \3390 );
or \U$3417 ( \3549 , \3546 , \3547 , \3548 );
xor \U$3418 ( \3550 , \3545 , \3549 );
xor \U$3419 ( \3551 , \3536 , \3550 );
and \U$3420 ( \3552 , \150 , \3357 );
and \U$3421 ( \3553 , \158 , \3255 );
nor \U$3422 ( \3554 , \3552 , \3553 );
xnor \U$3423 ( \3555 , \3554 , \3156 );
buf \U$3424 ( \3556 , RIb560318_28);
xor \U$3425 ( \3557 , \3556 , \3152 );
nand \U$3426 ( \3558 , \166 , \3557 );
buf \U$3427 ( \3559 , RIb560390_27);
and \U$3428 ( \3560 , \3556 , \3152 );
not \U$3429 ( \3561 , \3560 );
and \U$3430 ( \3562 , \3559 , \3561 );
xnor \U$3431 ( \3563 , \3558 , \3562 );
xor \U$3432 ( \3564 , \3555 , \3563 );
and \U$3433 ( \3565 , \224 , \2400 );
and \U$3434 ( \3566 , \232 , \2246 );
nor \U$3435 ( \3567 , \3565 , \3566 );
xnor \U$3436 ( \3568 , \3567 , \2195 );
and \U$3437 ( \3569 , \240 , \2669 );
and \U$3438 ( \3570 , \247 , \2538 );
nor \U$3439 ( \3571 , \3569 , \3570 );
xnor \U$3440 ( \3572 , \3571 , \2534 );
xor \U$3441 ( \3573 , \3568 , \3572 );
and \U$3442 ( \3574 , \134 , \3103 );
and \U$3443 ( \3575 , \143 , \2934 );
nor \U$3444 ( \3576 , \3574 , \3575 );
xnor \U$3445 ( \3577 , \3576 , \2839 );
xor \U$3446 ( \3578 , \3573 , \3577 );
xor \U$3447 ( \3579 , \3564 , \3578 );
xor \U$3448 ( \3580 , \3551 , \3579 );
xor \U$3449 ( \3581 , \3522 , \3580 );
and \U$3450 ( \3582 , \3408 , \3422 );
and \U$3451 ( \3583 , \3422 , \3437 );
and \U$3452 ( \3584 , \3408 , \3437 );
or \U$3453 ( \3585 , \3582 , \3583 , \3584 );
and \U$3454 ( \3586 , \1802 , \141 );
and \U$3455 ( \3587 , \1948 , \139 );
nor \U$3456 ( \3588 , \3586 , \3587 );
xnor \U$3457 ( \3589 , \3588 , \148 );
and \U$3458 ( \3590 , \1601 , \156 );
and \U$3459 ( \3591 , \1684 , \154 );
nor \U$3460 ( \3592 , \3590 , \3591 );
xnor \U$3461 ( \3593 , \3592 , \163 );
xor \U$3462 ( \3594 , \3589 , \3593 );
and \U$3463 ( \3595 , \1333 , \296 );
and \U$3464 ( \3596 , \1484 , \168 );
nor \U$3465 ( \3597 , \3595 , \3596 );
xnor \U$3466 ( \3598 , \3597 , \173 );
xor \U$3467 ( \3599 , \3594 , \3598 );
and \U$3468 ( \3600 , \1147 , \438 );
and \U$3469 ( \3601 , \1192 , \336 );
nor \U$3470 ( \3602 , \3600 , \3601 );
xnor \U$3471 ( \3603 , \3602 , \320 );
and \U$3472 ( \3604 , \412 , \1086 );
and \U$3473 ( \3605 , \474 , \508 );
nor \U$3474 ( \3606 , \3604 , \3605 );
xnor \U$3475 ( \3607 , \3606 , \487 );
xor \U$3476 ( \3608 , \3603 , \3607 );
and \U$3477 ( \3609 , \261 , \1301 );
and \U$3478 ( \3610 , \307 , \1246 );
nor \U$3479 ( \3611 , \3609 , \3610 );
xnor \U$3480 ( \3612 , \3611 , \1205 );
xor \U$3481 ( \3613 , \3608 , \3612 );
xor \U$3482 ( \3614 , \3599 , \3613 );
and \U$3483 ( \3615 , \178 , \1578 );
and \U$3484 ( \3616 , \185 , \1431 );
nor \U$3485 ( \3617 , \3615 , \3616 );
xnor \U$3486 ( \3618 , \3617 , \1436 );
and \U$3487 ( \3619 , \189 , \1824 );
and \U$3488 ( \3620 , \197 , \1739 );
nor \U$3489 ( \3621 , \3619 , \3620 );
xnor \U$3490 ( \3622 , \3621 , \1697 );
xor \U$3491 ( \3623 , \3618 , \3622 );
and \U$3492 ( \3624 , \209 , \2121 );
and \U$3493 ( \3625 , \217 , \2008 );
nor \U$3494 ( \3626 , \3624 , \3625 );
xnor \U$3495 ( \3627 , \3626 , \1961 );
xor \U$3496 ( \3628 , \3623 , \3627 );
xor \U$3497 ( \3629 , \3614 , \3628 );
xor \U$3498 ( \3630 , \3585 , \3629 );
and \U$3499 ( \3631 , \2757 , \215 );
and \U$3500 ( \3632 , \2826 , \213 );
nor \U$3501 ( \3633 , \3631 , \3632 );
xnor \U$3502 ( \3634 , \3633 , \222 );
and \U$3503 ( \3635 , \2366 , \230 );
and \U$3504 ( \3636 , \2521 , \228 );
nor \U$3505 ( \3637 , \3635 , \3636 );
xnor \U$3506 ( \3638 , \3637 , \237 );
xor \U$3507 ( \3639 , \3634 , \3638 );
and \U$3508 ( \3640 , \2090 , \245 );
and \U$3509 ( \3641 , \2182 , \243 );
nor \U$3510 ( \3642 , \3640 , \3641 );
xnor \U$3511 ( \3643 , \3642 , \252 );
xor \U$3512 ( \3644 , \3639 , \3643 );
and \U$3513 ( \3645 , \3395 , \183 );
buf \U$3514 ( \3646 , RIb55e518_92);
and \U$3515 ( \3647 , \3646 , \180 );
nor \U$3516 ( \3648 , \3645 , \3647 );
xnor \U$3517 ( \3649 , \3648 , \179 );
and \U$3518 ( \3650 , \3037 , \195 );
and \U$3519 ( \3651 , \3143 , \193 );
nor \U$3520 ( \3652 , \3650 , \3651 );
xnor \U$3521 ( \3653 , \3652 , \202 );
xor \U$3522 ( \3654 , \3649 , \3653 );
xor \U$3523 ( \3655 , \3654 , \3562 );
xor \U$3524 ( \3656 , \3644 , \3655 );
xor \U$3525 ( \3657 , \3630 , \3656 );
xor \U$3526 ( \3658 , \3581 , \3657 );
xor \U$3527 ( \3659 , \3508 , \3658 );
xor \U$3528 ( \3660 , \3499 , \3659 );
and \U$3529 ( \3661 , \3306 , \3307 );
and \U$3530 ( \3662 , \3307 , \3471 );
and \U$3531 ( \3663 , \3306 , \3471 );
or \U$3532 ( \3664 , \3661 , \3662 , \3663 );
xor \U$3533 ( \3665 , \3660 , \3664 );
and \U$3534 ( \3666 , \3472 , \3476 );
and \U$3535 ( \3667 , \3477 , \3480 );
or \U$3536 ( \3668 , \3666 , \3667 );
xor \U$3537 ( \3669 , \3665 , \3668 );
buf \U$3538 ( \3670 , \3669 );
buf \U$3539 ( \3671 , \3670 );
and \U$3540 ( \3672 , \3503 , \3507 );
and \U$3541 ( \3673 , \3507 , \3658 );
and \U$3542 ( \3674 , \3503 , \3658 );
or \U$3543 ( \3675 , \3672 , \3673 , \3674 );
and \U$3544 ( \3676 , \3491 , \3495 );
and \U$3545 ( \3677 , \3495 , \3497 );
and \U$3546 ( \3678 , \3491 , \3497 );
or \U$3547 ( \3679 , \3676 , \3677 , \3678 );
and \U$3548 ( \3680 , \3522 , \3580 );
and \U$3549 ( \3681 , \3580 , \3657 );
and \U$3550 ( \3682 , \3522 , \3657 );
or \U$3551 ( \3683 , \3680 , \3681 , \3682 );
xor \U$3552 ( \3684 , \3679 , \3683 );
and \U$3553 ( \3685 , \3526 , \3530 );
and \U$3554 ( \3686 , \3530 , \3535 );
and \U$3555 ( \3687 , \3526 , \3535 );
or \U$3556 ( \3688 , \3685 , \3686 , \3687 );
and \U$3557 ( \3689 , \3540 , \3544 );
and \U$3558 ( \3690 , \3544 , \3549 );
and \U$3559 ( \3691 , \3540 , \3549 );
or \U$3560 ( \3692 , \3689 , \3690 , \3691 );
xor \U$3561 ( \3693 , \3688 , \3692 );
and \U$3562 ( \3694 , \3555 , \3563 );
and \U$3563 ( \3695 , \3563 , \3578 );
and \U$3564 ( \3696 , \3555 , \3578 );
or \U$3565 ( \3697 , \3694 , \3695 , \3696 );
xor \U$3566 ( \3698 , \3693 , \3697 );
xor \U$3567 ( \3699 , \3684 , \3698 );
xor \U$3568 ( \3700 , \3675 , \3699 );
and \U$3569 ( \3701 , \3512 , \3516 );
and \U$3570 ( \3702 , \3516 , \3521 );
and \U$3571 ( \3703 , \3512 , \3521 );
or \U$3572 ( \3704 , \3701 , \3702 , \3703 );
and \U$3573 ( \3705 , \3536 , \3550 );
and \U$3574 ( \3706 , \3550 , \3579 );
and \U$3575 ( \3707 , \3536 , \3579 );
or \U$3576 ( \3708 , \3705 , \3706 , \3707 );
xor \U$3577 ( \3709 , \3704 , \3708 );
and \U$3578 ( \3710 , \3585 , \3629 );
and \U$3579 ( \3711 , \3629 , \3656 );
and \U$3580 ( \3712 , \3585 , \3656 );
or \U$3581 ( \3713 , \3710 , \3711 , \3712 );
xor \U$3582 ( \3714 , \3709 , \3713 );
and \U$3583 ( \3715 , \3589 , \3593 );
and \U$3584 ( \3716 , \3593 , \3598 );
and \U$3585 ( \3717 , \3589 , \3598 );
or \U$3586 ( \3718 , \3715 , \3716 , \3717 );
and \U$3587 ( \3719 , \3634 , \3638 );
and \U$3588 ( \3720 , \3638 , \3643 );
and \U$3589 ( \3721 , \3634 , \3643 );
or \U$3590 ( \3722 , \3719 , \3720 , \3721 );
xor \U$3591 ( \3723 , \3718 , \3722 );
and \U$3592 ( \3724 , \3649 , \3653 );
and \U$3593 ( \3725 , \3653 , \3562 );
and \U$3594 ( \3726 , \3649 , \3562 );
or \U$3595 ( \3727 , \3724 , \3725 , \3726 );
xor \U$3596 ( \3728 , \3723 , \3727 );
and \U$3597 ( \3729 , \3599 , \3613 );
and \U$3598 ( \3730 , \3613 , \3628 );
and \U$3599 ( \3731 , \3599 , \3628 );
or \U$3600 ( \3732 , \3729 , \3730 , \3731 );
and \U$3601 ( \3733 , \3644 , \3655 );
xor \U$3602 ( \3734 , \3732 , \3733 );
and \U$3603 ( \3735 , \3646 , \183 );
buf \U$3604 ( \3736 , RIb55e590_91);
and \U$3605 ( \3737 , \3736 , \180 );
nor \U$3606 ( \3738 , \3735 , \3737 );
xnor \U$3607 ( \3739 , \3738 , \179 );
and \U$3608 ( \3740 , \3143 , \195 );
and \U$3609 ( \3741 , \3395 , \193 );
nor \U$3610 ( \3742 , \3740 , \3741 );
xnor \U$3611 ( \3743 , \3742 , \202 );
xor \U$3612 ( \3744 , \3739 , \3743 );
and \U$3613 ( \3745 , \2826 , \215 );
and \U$3614 ( \3746 , \3037 , \213 );
nor \U$3615 ( \3747 , \3745 , \3746 );
xnor \U$3616 ( \3748 , \3747 , \222 );
xor \U$3617 ( \3749 , \3744 , \3748 );
xor \U$3618 ( \3750 , \3734 , \3749 );
xor \U$3619 ( \3751 , \3728 , \3750 );
and \U$3620 ( \3752 , \3568 , \3572 );
and \U$3621 ( \3753 , \3572 , \3577 );
and \U$3622 ( \3754 , \3568 , \3577 );
or \U$3623 ( \3755 , \3752 , \3753 , \3754 );
and \U$3624 ( \3756 , \3603 , \3607 );
and \U$3625 ( \3757 , \3607 , \3612 );
and \U$3626 ( \3758 , \3603 , \3612 );
or \U$3627 ( \3759 , \3756 , \3757 , \3758 );
xor \U$3628 ( \3760 , \3755 , \3759 );
and \U$3629 ( \3761 , \3618 , \3622 );
and \U$3630 ( \3762 , \3622 , \3627 );
and \U$3631 ( \3763 , \3618 , \3627 );
or \U$3632 ( \3764 , \3761 , \3762 , \3763 );
xor \U$3633 ( \3765 , \3760 , \3764 );
and \U$3634 ( \3766 , \1684 , \156 );
and \U$3635 ( \3767 , \1802 , \154 );
nor \U$3636 ( \3768 , \3766 , \3767 );
xnor \U$3637 ( \3769 , \3768 , \163 );
and \U$3638 ( \3770 , \1484 , \296 );
and \U$3639 ( \3771 , \1601 , \168 );
nor \U$3640 ( \3772 , \3770 , \3771 );
xnor \U$3641 ( \3773 , \3772 , \173 );
xor \U$3642 ( \3774 , \3769 , \3773 );
and \U$3643 ( \3775 , \1192 , \438 );
and \U$3644 ( \3776 , \1333 , \336 );
nor \U$3645 ( \3777 , \3775 , \3776 );
xnor \U$3646 ( \3778 , \3777 , \320 );
xor \U$3647 ( \3779 , \3774 , \3778 );
and \U$3648 ( \3780 , \474 , \1086 );
and \U$3649 ( \3781 , \1147 , \508 );
nor \U$3650 ( \3782 , \3780 , \3781 );
xnor \U$3651 ( \3783 , \3782 , \487 );
and \U$3652 ( \3784 , \307 , \1301 );
and \U$3653 ( \3785 , \412 , \1246 );
nor \U$3654 ( \3786 , \3784 , \3785 );
xnor \U$3655 ( \3787 , \3786 , \1205 );
xor \U$3656 ( \3788 , \3783 , \3787 );
and \U$3657 ( \3789 , \185 , \1578 );
and \U$3658 ( \3790 , \261 , \1431 );
nor \U$3659 ( \3791 , \3789 , \3790 );
xnor \U$3660 ( \3792 , \3791 , \1436 );
xor \U$3661 ( \3793 , \3788 , \3792 );
xor \U$3662 ( \3794 , \3779 , \3793 );
and \U$3663 ( \3795 , \2521 , \230 );
and \U$3664 ( \3796 , \2757 , \228 );
nor \U$3665 ( \3797 , \3795 , \3796 );
xnor \U$3666 ( \3798 , \3797 , \237 );
and \U$3667 ( \3799 , \2182 , \245 );
and \U$3668 ( \3800 , \2366 , \243 );
nor \U$3669 ( \3801 , \3799 , \3800 );
xnor \U$3670 ( \3802 , \3801 , \252 );
xor \U$3671 ( \3803 , \3798 , \3802 );
and \U$3672 ( \3804 , \1948 , \141 );
and \U$3673 ( \3805 , \2090 , \139 );
nor \U$3674 ( \3806 , \3804 , \3805 );
xnor \U$3675 ( \3807 , \3806 , \148 );
xor \U$3676 ( \3808 , \3803 , \3807 );
xor \U$3677 ( \3809 , \3794 , \3808 );
xor \U$3678 ( \3810 , \3765 , \3809 );
xor \U$3679 ( \3811 , \3559 , \3556 );
not \U$3680 ( \3812 , \3557 );
and \U$3681 ( \3813 , \3811 , \3812 );
and \U$3682 ( \3814 , \166 , \3813 );
and \U$3683 ( \3815 , \150 , \3557 );
nor \U$3684 ( \3816 , \3814 , \3815 );
xnor \U$3685 ( \3817 , \3816 , \3562 );
and \U$3686 ( \3818 , \247 , \2669 );
and \U$3687 ( \3819 , \224 , \2538 );
nor \U$3688 ( \3820 , \3818 , \3819 );
xnor \U$3689 ( \3821 , \3820 , \2534 );
and \U$3690 ( \3822 , \143 , \3103 );
and \U$3691 ( \3823 , \240 , \2934 );
nor \U$3692 ( \3824 , \3822 , \3823 );
xnor \U$3693 ( \3825 , \3824 , \2839 );
xor \U$3694 ( \3826 , \3821 , \3825 );
and \U$3695 ( \3827 , \158 , \3357 );
and \U$3696 ( \3828 , \134 , \3255 );
nor \U$3697 ( \3829 , \3827 , \3828 );
xnor \U$3698 ( \3830 , \3829 , \3156 );
xor \U$3699 ( \3831 , \3826 , \3830 );
xor \U$3700 ( \3832 , \3817 , \3831 );
and \U$3701 ( \3833 , \197 , \1824 );
and \U$3702 ( \3834 , \178 , \1739 );
nor \U$3703 ( \3835 , \3833 , \3834 );
xnor \U$3704 ( \3836 , \3835 , \1697 );
and \U$3705 ( \3837 , \217 , \2121 );
and \U$3706 ( \3838 , \189 , \2008 );
nor \U$3707 ( \3839 , \3837 , \3838 );
xnor \U$3708 ( \3840 , \3839 , \1961 );
xor \U$3709 ( \3841 , \3836 , \3840 );
and \U$3710 ( \3842 , \232 , \2400 );
and \U$3711 ( \3843 , \209 , \2246 );
nor \U$3712 ( \3844 , \3842 , \3843 );
xnor \U$3713 ( \3845 , \3844 , \2195 );
xor \U$3714 ( \3846 , \3841 , \3845 );
xor \U$3715 ( \3847 , \3832 , \3846 );
xor \U$3716 ( \3848 , \3810 , \3847 );
xor \U$3717 ( \3849 , \3751 , \3848 );
xor \U$3718 ( \3850 , \3714 , \3849 );
xor \U$3719 ( \3851 , \3700 , \3850 );
and \U$3720 ( \3852 , \3487 , \3498 );
and \U$3721 ( \3853 , \3498 , \3659 );
and \U$3722 ( \3854 , \3487 , \3659 );
or \U$3723 ( \3855 , \3852 , \3853 , \3854 );
xor \U$3724 ( \3856 , \3851 , \3855 );
and \U$3725 ( \3857 , \3660 , \3664 );
and \U$3726 ( \3858 , \3665 , \3668 );
or \U$3727 ( \3859 , \3857 , \3858 );
xor \U$3728 ( \3860 , \3856 , \3859 );
buf \U$3729 ( \3861 , \3860 );
buf \U$3730 ( \3862 , \3861 );
and \U$3731 ( \3863 , \3679 , \3683 );
and \U$3732 ( \3864 , \3683 , \3698 );
and \U$3733 ( \3865 , \3679 , \3698 );
or \U$3734 ( \3866 , \3863 , \3864 , \3865 );
and \U$3735 ( \3867 , \3714 , \3849 );
xor \U$3736 ( \3868 , \3866 , \3867 );
and \U$3737 ( \3869 , \3688 , \3692 );
and \U$3738 ( \3870 , \3692 , \3697 );
and \U$3739 ( \3871 , \3688 , \3697 );
or \U$3740 ( \3872 , \3869 , \3870 , \3871 );
and \U$3741 ( \3873 , \3732 , \3733 );
and \U$3742 ( \3874 , \3733 , \3749 );
and \U$3743 ( \3875 , \3732 , \3749 );
or \U$3744 ( \3876 , \3873 , \3874 , \3875 );
xor \U$3745 ( \3877 , \3872 , \3876 );
and \U$3746 ( \3878 , \3765 , \3809 );
and \U$3747 ( \3879 , \3809 , \3847 );
and \U$3748 ( \3880 , \3765 , \3847 );
or \U$3749 ( \3881 , \3878 , \3879 , \3880 );
xor \U$3750 ( \3882 , \3877 , \3881 );
xor \U$3751 ( \3883 , \3868 , \3882 );
and \U$3752 ( \3884 , \3704 , \3708 );
and \U$3753 ( \3885 , \3708 , \3713 );
and \U$3754 ( \3886 , \3704 , \3713 );
or \U$3755 ( \3887 , \3884 , \3885 , \3886 );
and \U$3756 ( \3888 , \3728 , \3750 );
and \U$3757 ( \3889 , \3750 , \3848 );
and \U$3758 ( \3890 , \3728 , \3848 );
or \U$3759 ( \3891 , \3888 , \3889 , \3890 );
xor \U$3760 ( \3892 , \3887 , \3891 );
and \U$3761 ( \3893 , \3718 , \3722 );
and \U$3762 ( \3894 , \3722 , \3727 );
and \U$3763 ( \3895 , \3718 , \3727 );
or \U$3764 ( \3896 , \3893 , \3894 , \3895 );
and \U$3765 ( \3897 , \3755 , \3759 );
and \U$3766 ( \3898 , \3759 , \3764 );
and \U$3767 ( \3899 , \3755 , \3764 );
or \U$3768 ( \3900 , \3897 , \3898 , \3899 );
xor \U$3769 ( \3901 , \3896 , \3900 );
and \U$3770 ( \3902 , \3817 , \3831 );
and \U$3771 ( \3903 , \3831 , \3846 );
and \U$3772 ( \3904 , \3817 , \3846 );
or \U$3773 ( \3905 , \3902 , \3903 , \3904 );
xor \U$3774 ( \3906 , \3901 , \3905 );
and \U$3775 ( \3907 , \3779 , \3793 );
and \U$3776 ( \3908 , \3793 , \3808 );
and \U$3777 ( \3909 , \3779 , \3808 );
or \U$3778 ( \3910 , \3907 , \3908 , \3909 );
and \U$3779 ( \3911 , \3736 , \183 );
buf \U$3780 ( \3912 , RIb55e608_90);
and \U$3781 ( \3913 , \3912 , \180 );
nor \U$3782 ( \3914 , \3911 , \3913 );
xnor \U$3783 ( \3915 , \3914 , \179 );
and \U$3784 ( \3916 , \3395 , \195 );
and \U$3785 ( \3917 , \3646 , \193 );
nor \U$3786 ( \3918 , \3916 , \3917 );
xnor \U$3787 ( \3919 , \3918 , \202 );
xor \U$3788 ( \3920 , \3915 , \3919 );
buf \U$3789 ( \3921 , RIb560480_25);
buf \U$3790 ( \3922 , RIb560408_26);
and \U$3791 ( \3923 , \3922 , \3559 );
not \U$3792 ( \3924 , \3923 );
and \U$3793 ( \3925 , \3921 , \3924 );
xor \U$3794 ( \3926 , \3920 , \3925 );
xor \U$3795 ( \3927 , \3910 , \3926 );
and \U$3796 ( \3928 , \1333 , \438 );
and \U$3797 ( \3929 , \1484 , \336 );
nor \U$3798 ( \3930 , \3928 , \3929 );
xnor \U$3799 ( \3931 , \3930 , \320 );
and \U$3800 ( \3932 , \1147 , \1086 );
and \U$3801 ( \3933 , \1192 , \508 );
nor \U$3802 ( \3934 , \3932 , \3933 );
xnor \U$3803 ( \3935 , \3934 , \487 );
xor \U$3804 ( \3936 , \3931 , \3935 );
and \U$3805 ( \3937 , \412 , \1301 );
and \U$3806 ( \3938 , \474 , \1246 );
nor \U$3807 ( \3939 , \3937 , \3938 );
xnor \U$3808 ( \3940 , \3939 , \1205 );
xor \U$3809 ( \3941 , \3936 , \3940 );
and \U$3810 ( \3942 , \2090 , \141 );
and \U$3811 ( \3943 , \2182 , \139 );
nor \U$3812 ( \3944 , \3942 , \3943 );
xnor \U$3813 ( \3945 , \3944 , \148 );
and \U$3814 ( \3946 , \1802 , \156 );
and \U$3815 ( \3947 , \1948 , \154 );
nor \U$3816 ( \3948 , \3946 , \3947 );
xnor \U$3817 ( \3949 , \3948 , \163 );
xor \U$3818 ( \3950 , \3945 , \3949 );
and \U$3819 ( \3951 , \1601 , \296 );
and \U$3820 ( \3952 , \1684 , \168 );
nor \U$3821 ( \3953 , \3951 , \3952 );
xnor \U$3822 ( \3954 , \3953 , \173 );
xor \U$3823 ( \3955 , \3950 , \3954 );
xor \U$3824 ( \3956 , \3941 , \3955 );
and \U$3825 ( \3957 , \3037 , \215 );
and \U$3826 ( \3958 , \3143 , \213 );
nor \U$3827 ( \3959 , \3957 , \3958 );
xnor \U$3828 ( \3960 , \3959 , \222 );
and \U$3829 ( \3961 , \2757 , \230 );
and \U$3830 ( \3962 , \2826 , \228 );
nor \U$3831 ( \3963 , \3961 , \3962 );
xnor \U$3832 ( \3964 , \3963 , \237 );
xor \U$3833 ( \3965 , \3960 , \3964 );
and \U$3834 ( \3966 , \2366 , \245 );
and \U$3835 ( \3967 , \2521 , \243 );
nor \U$3836 ( \3968 , \3966 , \3967 );
xnor \U$3837 ( \3969 , \3968 , \252 );
xor \U$3838 ( \3970 , \3965 , \3969 );
xor \U$3839 ( \3971 , \3956 , \3970 );
xor \U$3840 ( \3972 , \3927 , \3971 );
xor \U$3841 ( \3973 , \3906 , \3972 );
and \U$3842 ( \3974 , \3821 , \3825 );
and \U$3843 ( \3975 , \3825 , \3830 );
and \U$3844 ( \3976 , \3821 , \3830 );
or \U$3845 ( \3977 , \3974 , \3975 , \3976 );
and \U$3846 ( \3978 , \3783 , \3787 );
and \U$3847 ( \3979 , \3787 , \3792 );
and \U$3848 ( \3980 , \3783 , \3792 );
or \U$3849 ( \3981 , \3978 , \3979 , \3980 );
xor \U$3850 ( \3982 , \3977 , \3981 );
and \U$3851 ( \3983 , \3836 , \3840 );
and \U$3852 ( \3984 , \3840 , \3845 );
and \U$3853 ( \3985 , \3836 , \3845 );
or \U$3854 ( \3986 , \3983 , \3984 , \3985 );
xor \U$3855 ( \3987 , \3982 , \3986 );
and \U$3856 ( \3988 , \3769 , \3773 );
and \U$3857 ( \3989 , \3773 , \3778 );
and \U$3858 ( \3990 , \3769 , \3778 );
or \U$3859 ( \3991 , \3988 , \3989 , \3990 );
and \U$3860 ( \3992 , \3798 , \3802 );
and \U$3861 ( \3993 , \3802 , \3807 );
and \U$3862 ( \3994 , \3798 , \3807 );
or \U$3863 ( \3995 , \3992 , \3993 , \3994 );
xor \U$3864 ( \3996 , \3991 , \3995 );
and \U$3865 ( \3997 , \3739 , \3743 );
and \U$3866 ( \3998 , \3743 , \3748 );
and \U$3867 ( \3999 , \3739 , \3748 );
or \U$3868 ( \4000 , \3997 , \3998 , \3999 );
xor \U$3869 ( \4001 , \3996 , \4000 );
xor \U$3870 ( \4002 , \3987 , \4001 );
and \U$3871 ( \4003 , \134 , \3357 );
and \U$3872 ( \4004 , \143 , \3255 );
nor \U$3873 ( \4005 , \4003 , \4004 );
xnor \U$3874 ( \4006 , \4005 , \3156 );
and \U$3875 ( \4007 , \150 , \3813 );
and \U$3876 ( \4008 , \158 , \3557 );
nor \U$3877 ( \4009 , \4007 , \4008 );
xnor \U$3878 ( \4010 , \4009 , \3562 );
xor \U$3879 ( \4011 , \4006 , \4010 );
xor \U$3880 ( \4012 , \3922 , \3559 );
nand \U$3881 ( \4013 , \166 , \4012 );
xnor \U$3882 ( \4014 , \4013 , \3925 );
xor \U$3883 ( \4015 , \4011 , \4014 );
and \U$3884 ( \4016 , \209 , \2400 );
and \U$3885 ( \4017 , \217 , \2246 );
nor \U$3886 ( \4018 , \4016 , \4017 );
xnor \U$3887 ( \4019 , \4018 , \2195 );
and \U$3888 ( \4020 , \224 , \2669 );
and \U$3889 ( \4021 , \232 , \2538 );
nor \U$3890 ( \4022 , \4020 , \4021 );
xnor \U$3891 ( \4023 , \4022 , \2534 );
xor \U$3892 ( \4024 , \4019 , \4023 );
and \U$3893 ( \4025 , \240 , \3103 );
and \U$3894 ( \4026 , \247 , \2934 );
nor \U$3895 ( \4027 , \4025 , \4026 );
xnor \U$3896 ( \4028 , \4027 , \2839 );
xor \U$3897 ( \4029 , \4024 , \4028 );
xor \U$3898 ( \4030 , \4015 , \4029 );
and \U$3899 ( \4031 , \261 , \1578 );
and \U$3900 ( \4032 , \307 , \1431 );
nor \U$3901 ( \4033 , \4031 , \4032 );
xnor \U$3902 ( \4034 , \4033 , \1436 );
and \U$3903 ( \4035 , \178 , \1824 );
and \U$3904 ( \4036 , \185 , \1739 );
nor \U$3905 ( \4037 , \4035 , \4036 );
xnor \U$3906 ( \4038 , \4037 , \1697 );
xor \U$3907 ( \4039 , \4034 , \4038 );
and \U$3908 ( \4040 , \189 , \2121 );
and \U$3909 ( \4041 , \197 , \2008 );
nor \U$3910 ( \4042 , \4040 , \4041 );
xnor \U$3911 ( \4043 , \4042 , \1961 );
xor \U$3912 ( \4044 , \4039 , \4043 );
xor \U$3913 ( \4045 , \4030 , \4044 );
xor \U$3914 ( \4046 , \4002 , \4045 );
xor \U$3915 ( \4047 , \3973 , \4046 );
xor \U$3916 ( \4048 , \3892 , \4047 );
xor \U$3917 ( \4049 , \3883 , \4048 );
and \U$3918 ( \4050 , \3675 , \3699 );
and \U$3919 ( \4051 , \3699 , \3850 );
and \U$3920 ( \4052 , \3675 , \3850 );
or \U$3921 ( \4053 , \4050 , \4051 , \4052 );
xor \U$3922 ( \4054 , \4049 , \4053 );
and \U$3923 ( \4055 , \3851 , \3855 );
and \U$3924 ( \4056 , \3856 , \3859 );
or \U$3925 ( \4057 , \4055 , \4056 );
xor \U$3926 ( \4058 , \4054 , \4057 );
buf \U$3927 ( \4059 , \4058 );
buf \U$3928 ( \4060 , \4059 );
and \U$3929 ( \4061 , \3866 , \3867 );
and \U$3930 ( \4062 , \3867 , \3882 );
and \U$3931 ( \4063 , \3866 , \3882 );
or \U$3932 ( \4064 , \4061 , \4062 , \4063 );
and \U$3933 ( \4065 , \3887 , \3891 );
and \U$3934 ( \4066 , \3891 , \4047 );
and \U$3935 ( \4067 , \3887 , \4047 );
or \U$3936 ( \4068 , \4065 , \4066 , \4067 );
and \U$3937 ( \4069 , \3896 , \3900 );
and \U$3938 ( \4070 , \3900 , \3905 );
and \U$3939 ( \4071 , \3896 , \3905 );
or \U$3940 ( \4072 , \4069 , \4070 , \4071 );
and \U$3941 ( \4073 , \3910 , \3926 );
and \U$3942 ( \4074 , \3926 , \3971 );
and \U$3943 ( \4075 , \3910 , \3971 );
or \U$3944 ( \4076 , \4073 , \4074 , \4075 );
xor \U$3945 ( \4077 , \4072 , \4076 );
and \U$3946 ( \4078 , \3987 , \4001 );
and \U$3947 ( \4079 , \4001 , \4045 );
and \U$3948 ( \4080 , \3987 , \4045 );
or \U$3949 ( \4081 , \4078 , \4079 , \4080 );
xor \U$3950 ( \4082 , \4077 , \4081 );
xor \U$3951 ( \4083 , \4068 , \4082 );
and \U$3952 ( \4084 , \3872 , \3876 );
and \U$3953 ( \4085 , \3876 , \3881 );
and \U$3954 ( \4086 , \3872 , \3881 );
or \U$3955 ( \4087 , \4084 , \4085 , \4086 );
and \U$3956 ( \4088 , \3906 , \3972 );
and \U$3957 ( \4089 , \3972 , \4046 );
and \U$3958 ( \4090 , \3906 , \4046 );
or \U$3959 ( \4091 , \4088 , \4089 , \4090 );
xor \U$3960 ( \4092 , \4087 , \4091 );
and \U$3961 ( \4093 , \3977 , \3981 );
and \U$3962 ( \4094 , \3981 , \3986 );
and \U$3963 ( \4095 , \3977 , \3986 );
or \U$3964 ( \4096 , \4093 , \4094 , \4095 );
and \U$3965 ( \4097 , \3991 , \3995 );
and \U$3966 ( \4098 , \3995 , \4000 );
and \U$3967 ( \4099 , \3991 , \4000 );
or \U$3968 ( \4100 , \4097 , \4098 , \4099 );
xor \U$3969 ( \4101 , \4096 , \4100 );
and \U$3970 ( \4102 , \4015 , \4029 );
and \U$3971 ( \4103 , \4029 , \4044 );
and \U$3972 ( \4104 , \4015 , \4044 );
or \U$3973 ( \4105 , \4102 , \4103 , \4104 );
xor \U$3974 ( \4106 , \4101 , \4105 );
and \U$3975 ( \4107 , \3915 , \3919 );
and \U$3976 ( \4108 , \3919 , \3925 );
and \U$3977 ( \4109 , \3915 , \3925 );
or \U$3978 ( \4110 , \4107 , \4108 , \4109 );
and \U$3979 ( \4111 , \3945 , \3949 );
and \U$3980 ( \4112 , \3949 , \3954 );
and \U$3981 ( \4113 , \3945 , \3954 );
or \U$3982 ( \4114 , \4111 , \4112 , \4113 );
xor \U$3983 ( \4115 , \4110 , \4114 );
and \U$3984 ( \4116 , \3960 , \3964 );
and \U$3985 ( \4117 , \3964 , \3969 );
and \U$3986 ( \4118 , \3960 , \3969 );
or \U$3987 ( \4119 , \4116 , \4117 , \4118 );
xor \U$3988 ( \4120 , \4115 , \4119 );
and \U$3989 ( \4121 , \4006 , \4010 );
and \U$3990 ( \4122 , \4010 , \4014 );
and \U$3991 ( \4123 , \4006 , \4014 );
or \U$3992 ( \4124 , \4121 , \4122 , \4123 );
and \U$3993 ( \4125 , \158 , \3813 );
and \U$3994 ( \4126 , \134 , \3557 );
nor \U$3995 ( \4127 , \4125 , \4126 );
xnor \U$3996 ( \4128 , \4127 , \3562 );
xor \U$3997 ( \4129 , \4124 , \4128 );
xor \U$3998 ( \4130 , \3921 , \3922 );
not \U$3999 ( \4131 , \4012 );
and \U$4000 ( \4132 , \4130 , \4131 );
and \U$4001 ( \4133 , \166 , \4132 );
and \U$4002 ( \4134 , \150 , \4012 );
nor \U$4003 ( \4135 , \4133 , \4134 );
xnor \U$4004 ( \4136 , \4135 , \3925 );
xor \U$4005 ( \4137 , \4129 , \4136 );
xor \U$4006 ( \4138 , \4120 , \4137 );
and \U$4007 ( \4139 , \3931 , \3935 );
and \U$4008 ( \4140 , \3935 , \3940 );
and \U$4009 ( \4141 , \3931 , \3940 );
or \U$4010 ( \4142 , \4139 , \4140 , \4141 );
and \U$4011 ( \4143 , \4019 , \4023 );
and \U$4012 ( \4144 , \4023 , \4028 );
and \U$4013 ( \4145 , \4019 , \4028 );
or \U$4014 ( \4146 , \4143 , \4144 , \4145 );
xor \U$4015 ( \4147 , \4142 , \4146 );
and \U$4016 ( \4148 , \4034 , \4038 );
and \U$4017 ( \4149 , \4038 , \4043 );
and \U$4018 ( \4150 , \4034 , \4043 );
or \U$4019 ( \4151 , \4148 , \4149 , \4150 );
xor \U$4020 ( \4152 , \4147 , \4151 );
xor \U$4021 ( \4153 , \4138 , \4152 );
xor \U$4022 ( \4154 , \4106 , \4153 );
and \U$4023 ( \4155 , \3941 , \3955 );
and \U$4024 ( \4156 , \3955 , \3970 );
and \U$4025 ( \4157 , \3941 , \3970 );
or \U$4026 ( \4158 , \4155 , \4156 , \4157 );
and \U$4027 ( \4159 , \3912 , \183 );
buf \U$4028 ( \4160 , RIb55e680_89);
and \U$4029 ( \4161 , \4160 , \180 );
nor \U$4030 ( \4162 , \4159 , \4161 );
xnor \U$4031 ( \4163 , \4162 , \179 );
and \U$4032 ( \4164 , \3646 , \195 );
and \U$4033 ( \4165 , \3736 , \193 );
nor \U$4034 ( \4166 , \4164 , \4165 );
xnor \U$4035 ( \4167 , \4166 , \202 );
xor \U$4036 ( \4168 , \4163 , \4167 );
and \U$4037 ( \4169 , \3143 , \215 );
and \U$4038 ( \4170 , \3395 , \213 );
nor \U$4039 ( \4171 , \4169 , \4170 );
xnor \U$4040 ( \4172 , \4171 , \222 );
xor \U$4041 ( \4173 , \4168 , \4172 );
and \U$4042 ( \4174 , \2826 , \230 );
and \U$4043 ( \4175 , \3037 , \228 );
nor \U$4044 ( \4176 , \4174 , \4175 );
xnor \U$4045 ( \4177 , \4176 , \237 );
and \U$4046 ( \4178 , \2521 , \245 );
and \U$4047 ( \4179 , \2757 , \243 );
nor \U$4048 ( \4180 , \4178 , \4179 );
xnor \U$4049 ( \4181 , \4180 , \252 );
xor \U$4050 ( \4182 , \4177 , \4181 );
and \U$4051 ( \4183 , \2182 , \141 );
and \U$4052 ( \4184 , \2366 , \139 );
nor \U$4053 ( \4185 , \4183 , \4184 );
xnor \U$4054 ( \4186 , \4185 , \148 );
xor \U$4055 ( \4187 , \4182 , \4186 );
xor \U$4056 ( \4188 , \4173 , \4187 );
and \U$4057 ( \4189 , \1948 , \156 );
and \U$4058 ( \4190 , \2090 , \154 );
nor \U$4059 ( \4191 , \4189 , \4190 );
xnor \U$4060 ( \4192 , \4191 , \163 );
and \U$4061 ( \4193 , \1684 , \296 );
and \U$4062 ( \4194 , \1802 , \168 );
nor \U$4063 ( \4195 , \4193 , \4194 );
xnor \U$4064 ( \4196 , \4195 , \173 );
xor \U$4065 ( \4197 , \4192 , \4196 );
and \U$4066 ( \4198 , \1484 , \438 );
and \U$4067 ( \4199 , \1601 , \336 );
nor \U$4068 ( \4200 , \4198 , \4199 );
xnor \U$4069 ( \4201 , \4200 , \320 );
xor \U$4070 ( \4202 , \4197 , \4201 );
xor \U$4071 ( \4203 , \4188 , \4202 );
xor \U$4072 ( \4204 , \4158 , \4203 );
and \U$4073 ( \4205 , \185 , \1824 );
and \U$4074 ( \4206 , \261 , \1739 );
nor \U$4075 ( \4207 , \4205 , \4206 );
xnor \U$4076 ( \4208 , \4207 , \1697 );
and \U$4077 ( \4209 , \197 , \2121 );
and \U$4078 ( \4210 , \178 , \2008 );
nor \U$4079 ( \4211 , \4209 , \4210 );
xnor \U$4080 ( \4212 , \4211 , \1961 );
xor \U$4081 ( \4213 , \4208 , \4212 );
and \U$4082 ( \4214 , \217 , \2400 );
and \U$4083 ( \4215 , \189 , \2246 );
nor \U$4084 ( \4216 , \4214 , \4215 );
xnor \U$4085 ( \4217 , \4216 , \2195 );
xor \U$4086 ( \4218 , \4213 , \4217 );
and \U$4087 ( \4219 , \1192 , \1086 );
and \U$4088 ( \4220 , \1333 , \508 );
nor \U$4089 ( \4221 , \4219 , \4220 );
xnor \U$4090 ( \4222 , \4221 , \487 );
and \U$4091 ( \4223 , \474 , \1301 );
and \U$4092 ( \4224 , \1147 , \1246 );
nor \U$4093 ( \4225 , \4223 , \4224 );
xnor \U$4094 ( \4226 , \4225 , \1205 );
xor \U$4095 ( \4227 , \4222 , \4226 );
and \U$4096 ( \4228 , \307 , \1578 );
and \U$4097 ( \4229 , \412 , \1431 );
nor \U$4098 ( \4230 , \4228 , \4229 );
xnor \U$4099 ( \4231 , \4230 , \1436 );
xor \U$4100 ( \4232 , \4227 , \4231 );
xor \U$4101 ( \4233 , \4218 , \4232 );
and \U$4102 ( \4234 , \232 , \2669 );
and \U$4103 ( \4235 , \209 , \2538 );
nor \U$4104 ( \4236 , \4234 , \4235 );
xnor \U$4105 ( \4237 , \4236 , \2534 );
and \U$4106 ( \4238 , \247 , \3103 );
and \U$4107 ( \4239 , \224 , \2934 );
nor \U$4108 ( \4240 , \4238 , \4239 );
xnor \U$4109 ( \4241 , \4240 , \2839 );
xor \U$4110 ( \4242 , \4237 , \4241 );
and \U$4111 ( \4243 , \143 , \3357 );
and \U$4112 ( \4244 , \240 , \3255 );
nor \U$4113 ( \4245 , \4243 , \4244 );
xnor \U$4114 ( \4246 , \4245 , \3156 );
xor \U$4115 ( \4247 , \4242 , \4246 );
xor \U$4116 ( \4248 , \4233 , \4247 );
xor \U$4117 ( \4249 , \4204 , \4248 );
xor \U$4118 ( \4250 , \4154 , \4249 );
xor \U$4119 ( \4251 , \4092 , \4250 );
xor \U$4120 ( \4252 , \4083 , \4251 );
xor \U$4121 ( \4253 , \4064 , \4252 );
and \U$4122 ( \4254 , \3883 , \4048 );
xor \U$4123 ( \4255 , \4253 , \4254 );
and \U$4124 ( \4256 , \4049 , \4053 );
and \U$4125 ( \4257 , \4054 , \4057 );
or \U$4126 ( \4258 , \4256 , \4257 );
xor \U$4127 ( \4259 , \4255 , \4258 );
buf \U$4128 ( \4260 , \4259 );
buf \U$4129 ( \4261 , \4260 );
and \U$4130 ( \4262 , \4068 , \4082 );
and \U$4131 ( \4263 , \4082 , \4251 );
and \U$4132 ( \4264 , \4068 , \4251 );
or \U$4133 ( \4265 , \4262 , \4263 , \4264 );
and \U$4134 ( \4266 , \4087 , \4091 );
and \U$4135 ( \4267 , \4091 , \4250 );
and \U$4136 ( \4268 , \4087 , \4250 );
or \U$4137 ( \4269 , \4266 , \4267 , \4268 );
and \U$4138 ( \4270 , \4072 , \4076 );
and \U$4139 ( \4271 , \4076 , \4081 );
and \U$4140 ( \4272 , \4072 , \4081 );
or \U$4141 ( \4273 , \4270 , \4271 , \4272 );
and \U$4142 ( \4274 , \4106 , \4153 );
and \U$4143 ( \4275 , \4153 , \4249 );
and \U$4144 ( \4276 , \4106 , \4249 );
or \U$4145 ( \4277 , \4274 , \4275 , \4276 );
xor \U$4146 ( \4278 , \4273 , \4277 );
and \U$4147 ( \4279 , \4173 , \4187 );
and \U$4148 ( \4280 , \4187 , \4202 );
and \U$4149 ( \4281 , \4173 , \4202 );
or \U$4150 ( \4282 , \4279 , \4280 , \4281 );
and \U$4151 ( \4283 , \4218 , \4232 );
and \U$4152 ( \4284 , \4232 , \4247 );
and \U$4153 ( \4285 , \4218 , \4247 );
or \U$4154 ( \4286 , \4283 , \4284 , \4285 );
xor \U$4155 ( \4287 , \4282 , \4286 );
and \U$4156 ( \4288 , \3395 , \215 );
and \U$4157 ( \4289 , \3646 , \213 );
nor \U$4158 ( \4290 , \4288 , \4289 );
xnor \U$4159 ( \4291 , \4290 , \222 );
and \U$4160 ( \4292 , \3037 , \230 );
and \U$4161 ( \4293 , \3143 , \228 );
nor \U$4162 ( \4294 , \4292 , \4293 );
xnor \U$4163 ( \4295 , \4294 , \237 );
xor \U$4164 ( \4296 , \4291 , \4295 );
and \U$4165 ( \4297 , \2757 , \245 );
and \U$4166 ( \4298 , \2826 , \243 );
nor \U$4167 ( \4299 , \4297 , \4298 );
xnor \U$4168 ( \4300 , \4299 , \252 );
xor \U$4169 ( \4301 , \4296 , \4300 );
xor \U$4170 ( \4302 , \4287 , \4301 );
xor \U$4171 ( \4303 , \4278 , \4302 );
xor \U$4172 ( \4304 , \4269 , \4303 );
and \U$4173 ( \4305 , \4110 , \4114 );
and \U$4174 ( \4306 , \4114 , \4119 );
and \U$4175 ( \4307 , \4110 , \4119 );
or \U$4176 ( \4308 , \4305 , \4306 , \4307 );
and \U$4177 ( \4309 , \4124 , \4128 );
and \U$4178 ( \4310 , \4128 , \4136 );
and \U$4179 ( \4311 , \4124 , \4136 );
or \U$4180 ( \4312 , \4309 , \4310 , \4311 );
xor \U$4181 ( \4313 , \4308 , \4312 );
and \U$4182 ( \4314 , \4142 , \4146 );
and \U$4183 ( \4315 , \4146 , \4151 );
and \U$4184 ( \4316 , \4142 , \4151 );
or \U$4185 ( \4317 , \4314 , \4315 , \4316 );
xor \U$4186 ( \4318 , \4313 , \4317 );
and \U$4187 ( \4319 , \4096 , \4100 );
and \U$4188 ( \4320 , \4100 , \4105 );
and \U$4189 ( \4321 , \4096 , \4105 );
or \U$4190 ( \4322 , \4319 , \4320 , \4321 );
and \U$4191 ( \4323 , \4120 , \4137 );
and \U$4192 ( \4324 , \4137 , \4152 );
and \U$4193 ( \4325 , \4120 , \4152 );
or \U$4194 ( \4326 , \4323 , \4324 , \4325 );
xor \U$4195 ( \4327 , \4322 , \4326 );
and \U$4196 ( \4328 , \4158 , \4203 );
and \U$4197 ( \4329 , \4203 , \4248 );
and \U$4198 ( \4330 , \4158 , \4248 );
or \U$4199 ( \4331 , \4328 , \4329 , \4330 );
xor \U$4200 ( \4332 , \4327 , \4331 );
xor \U$4201 ( \4333 , \4318 , \4332 );
and \U$4202 ( \4334 , \4163 , \4167 );
and \U$4203 ( \4335 , \4167 , \4172 );
and \U$4204 ( \4336 , \4163 , \4172 );
or \U$4205 ( \4337 , \4334 , \4335 , \4336 );
and \U$4206 ( \4338 , \4177 , \4181 );
and \U$4207 ( \4339 , \4181 , \4186 );
and \U$4208 ( \4340 , \4177 , \4186 );
or \U$4209 ( \4341 , \4338 , \4339 , \4340 );
xor \U$4210 ( \4342 , \4337 , \4341 );
and \U$4211 ( \4343 , \4192 , \4196 );
and \U$4212 ( \4344 , \4196 , \4201 );
and \U$4213 ( \4345 , \4192 , \4201 );
or \U$4214 ( \4346 , \4343 , \4344 , \4345 );
xor \U$4215 ( \4347 , \4342 , \4346 );
and \U$4216 ( \4348 , \4208 , \4212 );
and \U$4217 ( \4349 , \4212 , \4217 );
and \U$4218 ( \4350 , \4208 , \4217 );
or \U$4219 ( \4351 , \4348 , \4349 , \4350 );
and \U$4220 ( \4352 , \4222 , \4226 );
and \U$4221 ( \4353 , \4226 , \4231 );
and \U$4222 ( \4354 , \4222 , \4231 );
or \U$4223 ( \4355 , \4352 , \4353 , \4354 );
xor \U$4224 ( \4356 , \4351 , \4355 );
and \U$4225 ( \4357 , \4237 , \4241 );
and \U$4226 ( \4358 , \4241 , \4246 );
and \U$4227 ( \4359 , \4237 , \4246 );
or \U$4228 ( \4360 , \4357 , \4358 , \4359 );
xor \U$4229 ( \4361 , \4356 , \4360 );
xor \U$4230 ( \4362 , \4347 , \4361 );
and \U$4231 ( \4363 , \4160 , \183 );
buf \U$4232 ( \4364 , RIb55e6f8_88);
and \U$4233 ( \4365 , \4364 , \180 );
nor \U$4234 ( \4366 , \4363 , \4365 );
xnor \U$4235 ( \4367 , \4366 , \179 );
and \U$4236 ( \4368 , \3736 , \195 );
and \U$4237 ( \4369 , \3912 , \193 );
nor \U$4238 ( \4370 , \4368 , \4369 );
xnor \U$4239 ( \4371 , \4370 , \202 );
xor \U$4240 ( \4372 , \4367 , \4371 );
buf \U$4241 ( \4373 , RIb560570_23);
buf \U$4242 ( \4374 , RIb5604f8_24);
and \U$4243 ( \4375 , \4374 , \3921 );
not \U$4244 ( \4376 , \4375 );
and \U$4245 ( \4377 , \4373 , \4376 );
xor \U$4246 ( \4378 , \4372 , \4377 );
and \U$4247 ( \4379 , \2366 , \141 );
and \U$4248 ( \4380 , \2521 , \139 );
nor \U$4249 ( \4381 , \4379 , \4380 );
xnor \U$4250 ( \4382 , \4381 , \148 );
and \U$4251 ( \4383 , \2090 , \156 );
and \U$4252 ( \4384 , \2182 , \154 );
nor \U$4253 ( \4385 , \4383 , \4384 );
xnor \U$4254 ( \4386 , \4385 , \163 );
xor \U$4255 ( \4387 , \4382 , \4386 );
and \U$4256 ( \4388 , \1802 , \296 );
and \U$4257 ( \4389 , \1948 , \168 );
nor \U$4258 ( \4390 , \4388 , \4389 );
xnor \U$4259 ( \4391 , \4390 , \173 );
xor \U$4260 ( \4392 , \4387 , \4391 );
and \U$4261 ( \4393 , \1601 , \438 );
and \U$4262 ( \4394 , \1684 , \336 );
nor \U$4263 ( \4395 , \4393 , \4394 );
xnor \U$4264 ( \4396 , \4395 , \320 );
and \U$4265 ( \4397 , \1333 , \1086 );
and \U$4266 ( \4398 , \1484 , \508 );
nor \U$4267 ( \4399 , \4397 , \4398 );
xnor \U$4268 ( \4400 , \4399 , \487 );
xor \U$4269 ( \4401 , \4396 , \4400 );
and \U$4270 ( \4402 , \1147 , \1301 );
and \U$4271 ( \4403 , \1192 , \1246 );
nor \U$4272 ( \4404 , \4402 , \4403 );
xnor \U$4273 ( \4405 , \4404 , \1205 );
xor \U$4274 ( \4406 , \4401 , \4405 );
xor \U$4275 ( \4407 , \4392 , \4406 );
and \U$4276 ( \4408 , \412 , \1578 );
and \U$4277 ( \4409 , \474 , \1431 );
nor \U$4278 ( \4410 , \4408 , \4409 );
xnor \U$4279 ( \4411 , \4410 , \1436 );
and \U$4280 ( \4412 , \261 , \1824 );
and \U$4281 ( \4413 , \307 , \1739 );
nor \U$4282 ( \4414 , \4412 , \4413 );
xnor \U$4283 ( \4415 , \4414 , \1697 );
xor \U$4284 ( \4416 , \4411 , \4415 );
and \U$4285 ( \4417 , \178 , \2121 );
and \U$4286 ( \4418 , \185 , \2008 );
nor \U$4287 ( \4419 , \4417 , \4418 );
xnor \U$4288 ( \4420 , \4419 , \1961 );
xor \U$4289 ( \4421 , \4416 , \4420 );
xor \U$4290 ( \4422 , \4407 , \4421 );
xor \U$4291 ( \4423 , \4378 , \4422 );
xor \U$4292 ( \4424 , \4374 , \3921 );
nand \U$4293 ( \4425 , \166 , \4424 );
xnor \U$4294 ( \4426 , \4425 , \4377 );
and \U$4295 ( \4427 , \189 , \2400 );
and \U$4296 ( \4428 , \197 , \2246 );
nor \U$4297 ( \4429 , \4427 , \4428 );
xnor \U$4298 ( \4430 , \4429 , \2195 );
and \U$4299 ( \4431 , \209 , \2669 );
and \U$4300 ( \4432 , \217 , \2538 );
nor \U$4301 ( \4433 , \4431 , \4432 );
xnor \U$4302 ( \4434 , \4433 , \2534 );
xor \U$4303 ( \4435 , \4430 , \4434 );
and \U$4304 ( \4436 , \224 , \3103 );
and \U$4305 ( \4437 , \232 , \2934 );
nor \U$4306 ( \4438 , \4436 , \4437 );
xnor \U$4307 ( \4439 , \4438 , \2839 );
xor \U$4308 ( \4440 , \4435 , \4439 );
xor \U$4309 ( \4441 , \4426 , \4440 );
and \U$4310 ( \4442 , \240 , \3357 );
and \U$4311 ( \4443 , \247 , \3255 );
nor \U$4312 ( \4444 , \4442 , \4443 );
xnor \U$4313 ( \4445 , \4444 , \3156 );
and \U$4314 ( \4446 , \134 , \3813 );
and \U$4315 ( \4447 , \143 , \3557 );
nor \U$4316 ( \4448 , \4446 , \4447 );
xnor \U$4317 ( \4449 , \4448 , \3562 );
xor \U$4318 ( \4450 , \4445 , \4449 );
and \U$4319 ( \4451 , \150 , \4132 );
and \U$4320 ( \4452 , \158 , \4012 );
nor \U$4321 ( \4453 , \4451 , \4452 );
xnor \U$4322 ( \4454 , \4453 , \3925 );
xor \U$4323 ( \4455 , \4450 , \4454 );
xor \U$4324 ( \4456 , \4441 , \4455 );
xor \U$4325 ( \4457 , \4423 , \4456 );
xor \U$4326 ( \4458 , \4362 , \4457 );
xor \U$4327 ( \4459 , \4333 , \4458 );
xor \U$4328 ( \4460 , \4304 , \4459 );
xor \U$4329 ( \4461 , \4265 , \4460 );
and \U$4330 ( \4462 , \4064 , \4252 );
xor \U$4331 ( \4463 , \4461 , \4462 );
and \U$4332 ( \4464 , \4253 , \4254 );
and \U$4333 ( \4465 , \4255 , \4258 );
or \U$4334 ( \4466 , \4464 , \4465 );
xor \U$4335 ( \4467 , \4463 , \4466 );
buf \U$4336 ( \4468 , \4467 );
buf \U$4337 ( \4469 , \4468 );
and \U$4338 ( \4470 , \4269 , \4303 );
and \U$4339 ( \4471 , \4303 , \4459 );
and \U$4340 ( \4472 , \4269 , \4459 );
or \U$4341 ( \4473 , \4470 , \4471 , \4472 );
and \U$4342 ( \4474 , \4273 , \4277 );
and \U$4343 ( \4475 , \4277 , \4302 );
and \U$4344 ( \4476 , \4273 , \4302 );
or \U$4345 ( \4477 , \4474 , \4475 , \4476 );
and \U$4346 ( \4478 , \4318 , \4332 );
and \U$4347 ( \4479 , \4332 , \4458 );
and \U$4348 ( \4480 , \4318 , \4458 );
or \U$4349 ( \4481 , \4478 , \4479 , \4480 );
xor \U$4350 ( \4482 , \4477 , \4481 );
and \U$4351 ( \4483 , \4308 , \4312 );
and \U$4352 ( \4484 , \4312 , \4317 );
and \U$4353 ( \4485 , \4308 , \4317 );
or \U$4354 ( \4486 , \4483 , \4484 , \4485 );
and \U$4355 ( \4487 , \4282 , \4286 );
and \U$4356 ( \4488 , \4286 , \4301 );
and \U$4357 ( \4489 , \4282 , \4301 );
or \U$4358 ( \4490 , \4487 , \4488 , \4489 );
xor \U$4359 ( \4491 , \4486 , \4490 );
and \U$4360 ( \4492 , \4378 , \4422 );
and \U$4361 ( \4493 , \4422 , \4456 );
and \U$4362 ( \4494 , \4378 , \4456 );
or \U$4363 ( \4495 , \4492 , \4493 , \4494 );
xor \U$4364 ( \4496 , \4491 , \4495 );
xor \U$4365 ( \4497 , \4482 , \4496 );
xor \U$4366 ( \4498 , \4473 , \4497 );
and \U$4367 ( \4499 , \4322 , \4326 );
and \U$4368 ( \4500 , \4326 , \4331 );
and \U$4369 ( \4501 , \4322 , \4331 );
or \U$4370 ( \4502 , \4499 , \4500 , \4501 );
and \U$4371 ( \4503 , \4347 , \4361 );
and \U$4372 ( \4504 , \4361 , \4457 );
and \U$4373 ( \4505 , \4347 , \4457 );
or \U$4374 ( \4506 , \4503 , \4504 , \4505 );
xor \U$4375 ( \4507 , \4502 , \4506 );
and \U$4376 ( \4508 , \4337 , \4341 );
and \U$4377 ( \4509 , \4341 , \4346 );
and \U$4378 ( \4510 , \4337 , \4346 );
or \U$4379 ( \4511 , \4508 , \4509 , \4510 );
and \U$4380 ( \4512 , \4351 , \4355 );
and \U$4381 ( \4513 , \4355 , \4360 );
and \U$4382 ( \4514 , \4351 , \4360 );
or \U$4383 ( \4515 , \4512 , \4513 , \4514 );
xor \U$4384 ( \4516 , \4511 , \4515 );
and \U$4385 ( \4517 , \4426 , \4440 );
and \U$4386 ( \4518 , \4440 , \4455 );
and \U$4387 ( \4519 , \4426 , \4455 );
or \U$4388 ( \4520 , \4517 , \4518 , \4519 );
xor \U$4389 ( \4521 , \4516 , \4520 );
and \U$4390 ( \4522 , \4382 , \4386 );
and \U$4391 ( \4523 , \4386 , \4391 );
and \U$4392 ( \4524 , \4382 , \4391 );
or \U$4393 ( \4525 , \4522 , \4523 , \4524 );
and \U$4394 ( \4526 , \4291 , \4295 );
and \U$4395 ( \4527 , \4295 , \4300 );
and \U$4396 ( \4528 , \4291 , \4300 );
or \U$4397 ( \4529 , \4526 , \4527 , \4528 );
xor \U$4398 ( \4530 , \4525 , \4529 );
and \U$4399 ( \4531 , \4367 , \4371 );
and \U$4400 ( \4532 , \4371 , \4377 );
and \U$4401 ( \4533 , \4367 , \4377 );
or \U$4402 ( \4534 , \4531 , \4532 , \4533 );
xor \U$4403 ( \4535 , \4530 , \4534 );
and \U$4404 ( \4536 , \4430 , \4434 );
and \U$4405 ( \4537 , \4434 , \4439 );
and \U$4406 ( \4538 , \4430 , \4439 );
or \U$4407 ( \4539 , \4536 , \4537 , \4538 );
and \U$4408 ( \4540 , \4396 , \4400 );
and \U$4409 ( \4541 , \4400 , \4405 );
and \U$4410 ( \4542 , \4396 , \4405 );
or \U$4411 ( \4543 , \4540 , \4541 , \4542 );
xor \U$4412 ( \4544 , \4539 , \4543 );
and \U$4413 ( \4545 , \4411 , \4415 );
and \U$4414 ( \4546 , \4415 , \4420 );
and \U$4415 ( \4547 , \4411 , \4420 );
or \U$4416 ( \4548 , \4545 , \4546 , \4547 );
xor \U$4417 ( \4549 , \4544 , \4548 );
xor \U$4418 ( \4550 , \4535 , \4549 );
and \U$4419 ( \4551 , \4445 , \4449 );
and \U$4420 ( \4552 , \4449 , \4454 );
and \U$4421 ( \4553 , \4445 , \4454 );
or \U$4422 ( \4554 , \4551 , \4552 , \4553 );
and \U$4423 ( \4555 , \217 , \2669 );
and \U$4424 ( \4556 , \189 , \2538 );
nor \U$4425 ( \4557 , \4555 , \4556 );
xnor \U$4426 ( \4558 , \4557 , \2534 );
and \U$4427 ( \4559 , \232 , \3103 );
and \U$4428 ( \4560 , \209 , \2934 );
nor \U$4429 ( \4561 , \4559 , \4560 );
xnor \U$4430 ( \4562 , \4561 , \2839 );
xor \U$4431 ( \4563 , \4558 , \4562 );
and \U$4432 ( \4564 , \247 , \3357 );
and \U$4433 ( \4565 , \224 , \3255 );
nor \U$4434 ( \4566 , \4564 , \4565 );
xnor \U$4435 ( \4567 , \4566 , \3156 );
xor \U$4436 ( \4568 , \4563 , \4567 );
xor \U$4437 ( \4569 , \4554 , \4568 );
and \U$4438 ( \4570 , \143 , \3813 );
and \U$4439 ( \4571 , \240 , \3557 );
nor \U$4440 ( \4572 , \4570 , \4571 );
xnor \U$4441 ( \4573 , \4572 , \3562 );
and \U$4442 ( \4574 , \158 , \4132 );
and \U$4443 ( \4575 , \134 , \4012 );
nor \U$4444 ( \4576 , \4574 , \4575 );
xnor \U$4445 ( \4577 , \4576 , \3925 );
xor \U$4446 ( \4578 , \4573 , \4577 );
xor \U$4447 ( \4579 , \4373 , \4374 );
not \U$4448 ( \4580 , \4424 );
and \U$4449 ( \4581 , \4579 , \4580 );
and \U$4450 ( \4582 , \166 , \4581 );
and \U$4451 ( \4583 , \150 , \4424 );
nor \U$4452 ( \4584 , \4582 , \4583 );
xnor \U$4453 ( \4585 , \4584 , \4377 );
xor \U$4454 ( \4586 , \4578 , \4585 );
xor \U$4455 ( \4587 , \4569 , \4586 );
xor \U$4456 ( \4588 , \4550 , \4587 );
xor \U$4457 ( \4589 , \4521 , \4588 );
and \U$4458 ( \4590 , \4392 , \4406 );
and \U$4459 ( \4591 , \4406 , \4421 );
and \U$4460 ( \4592 , \4392 , \4421 );
or \U$4461 ( \4593 , \4590 , \4591 , \4592 );
and \U$4462 ( \4594 , \307 , \1824 );
and \U$4463 ( \4595 , \412 , \1739 );
nor \U$4464 ( \4596 , \4594 , \4595 );
xnor \U$4465 ( \4597 , \4596 , \1697 );
and \U$4466 ( \4598 , \185 , \2121 );
and \U$4467 ( \4599 , \261 , \2008 );
nor \U$4468 ( \4600 , \4598 , \4599 );
xnor \U$4469 ( \4601 , \4600 , \1961 );
xor \U$4470 ( \4602 , \4597 , \4601 );
and \U$4471 ( \4603 , \197 , \2400 );
and \U$4472 ( \4604 , \178 , \2246 );
nor \U$4473 ( \4605 , \4603 , \4604 );
xnor \U$4474 ( \4606 , \4605 , \2195 );
xor \U$4475 ( \4607 , \4602 , \4606 );
and \U$4476 ( \4608 , \2182 , \156 );
and \U$4477 ( \4609 , \2366 , \154 );
nor \U$4478 ( \4610 , \4608 , \4609 );
xnor \U$4479 ( \4611 , \4610 , \163 );
and \U$4480 ( \4612 , \1948 , \296 );
and \U$4481 ( \4613 , \2090 , \168 );
nor \U$4482 ( \4614 , \4612 , \4613 );
xnor \U$4483 ( \4615 , \4614 , \173 );
xor \U$4484 ( \4616 , \4611 , \4615 );
and \U$4485 ( \4617 , \1684 , \438 );
and \U$4486 ( \4618 , \1802 , \336 );
nor \U$4487 ( \4619 , \4617 , \4618 );
xnor \U$4488 ( \4620 , \4619 , \320 );
xor \U$4489 ( \4621 , \4616 , \4620 );
xor \U$4490 ( \4622 , \4607 , \4621 );
and \U$4491 ( \4623 , \1484 , \1086 );
and \U$4492 ( \4624 , \1601 , \508 );
nor \U$4493 ( \4625 , \4623 , \4624 );
xnor \U$4494 ( \4626 , \4625 , \487 );
and \U$4495 ( \4627 , \1192 , \1301 );
and \U$4496 ( \4628 , \1333 , \1246 );
nor \U$4497 ( \4629 , \4627 , \4628 );
xnor \U$4498 ( \4630 , \4629 , \1205 );
xor \U$4499 ( \4631 , \4626 , \4630 );
and \U$4500 ( \4632 , \474 , \1578 );
and \U$4501 ( \4633 , \1147 , \1431 );
nor \U$4502 ( \4634 , \4632 , \4633 );
xnor \U$4503 ( \4635 , \4634 , \1436 );
xor \U$4504 ( \4636 , \4631 , \4635 );
xor \U$4505 ( \4637 , \4622 , \4636 );
xor \U$4506 ( \4638 , \4593 , \4637 );
and \U$4507 ( \4639 , \3143 , \230 );
and \U$4508 ( \4640 , \3395 , \228 );
nor \U$4509 ( \4641 , \4639 , \4640 );
xnor \U$4510 ( \4642 , \4641 , \237 );
and \U$4511 ( \4643 , \2826 , \245 );
and \U$4512 ( \4644 , \3037 , \243 );
nor \U$4513 ( \4645 , \4643 , \4644 );
xnor \U$4514 ( \4646 , \4645 , \252 );
xor \U$4515 ( \4647 , \4642 , \4646 );
and \U$4516 ( \4648 , \2521 , \141 );
and \U$4517 ( \4649 , \2757 , \139 );
nor \U$4518 ( \4650 , \4648 , \4649 );
xnor \U$4519 ( \4651 , \4650 , \148 );
xor \U$4520 ( \4652 , \4647 , \4651 );
and \U$4521 ( \4653 , \4364 , \183 );
buf \U$4522 ( \4654 , RIb55e770_87);
and \U$4523 ( \4655 , \4654 , \180 );
nor \U$4524 ( \4656 , \4653 , \4655 );
xnor \U$4525 ( \4657 , \4656 , \179 );
and \U$4526 ( \4658 , \3912 , \195 );
and \U$4527 ( \4659 , \4160 , \193 );
nor \U$4528 ( \4660 , \4658 , \4659 );
xnor \U$4529 ( \4661 , \4660 , \202 );
xor \U$4530 ( \4662 , \4657 , \4661 );
and \U$4531 ( \4663 , \3646 , \215 );
and \U$4532 ( \4664 , \3736 , \213 );
nor \U$4533 ( \4665 , \4663 , \4664 );
xnor \U$4534 ( \4666 , \4665 , \222 );
xor \U$4535 ( \4667 , \4662 , \4666 );
xor \U$4536 ( \4668 , \4652 , \4667 );
xor \U$4537 ( \4669 , \4638 , \4668 );
xor \U$4538 ( \4670 , \4589 , \4669 );
xor \U$4539 ( \4671 , \4507 , \4670 );
xor \U$4540 ( \4672 , \4498 , \4671 );
and \U$4541 ( \4673 , \4265 , \4460 );
xor \U$4542 ( \4674 , \4672 , \4673 );
and \U$4543 ( \4675 , \4461 , \4462 );
and \U$4544 ( \4676 , \4463 , \4466 );
or \U$4545 ( \4677 , \4675 , \4676 );
xor \U$4546 ( \4678 , \4674 , \4677 );
buf \U$4547 ( \4679 , \4678 );
buf \U$4548 ( \4680 , \4679 );
and \U$4549 ( \4681 , \4477 , \4481 );
and \U$4550 ( \4682 , \4481 , \4496 );
and \U$4551 ( \4683 , \4477 , \4496 );
or \U$4552 ( \4684 , \4681 , \4682 , \4683 );
and \U$4553 ( \4685 , \4502 , \4506 );
and \U$4554 ( \4686 , \4506 , \4670 );
and \U$4555 ( \4687 , \4502 , \4670 );
or \U$4556 ( \4688 , \4685 , \4686 , \4687 );
and \U$4557 ( \4689 , \4486 , \4490 );
and \U$4558 ( \4690 , \4490 , \4495 );
and \U$4559 ( \4691 , \4486 , \4495 );
or \U$4560 ( \4692 , \4689 , \4690 , \4691 );
and \U$4561 ( \4693 , \4521 , \4588 );
and \U$4562 ( \4694 , \4588 , \4669 );
and \U$4563 ( \4695 , \4521 , \4669 );
or \U$4564 ( \4696 , \4693 , \4694 , \4695 );
xor \U$4565 ( \4697 , \4692 , \4696 );
and \U$4566 ( \4698 , \4525 , \4529 );
and \U$4567 ( \4699 , \4529 , \4534 );
and \U$4568 ( \4700 , \4525 , \4534 );
or \U$4569 ( \4701 , \4698 , \4699 , \4700 );
and \U$4570 ( \4702 , \4539 , \4543 );
and \U$4571 ( \4703 , \4543 , \4548 );
and \U$4572 ( \4704 , \4539 , \4548 );
or \U$4573 ( \4705 , \4702 , \4703 , \4704 );
xor \U$4574 ( \4706 , \4701 , \4705 );
and \U$4575 ( \4707 , \4554 , \4568 );
and \U$4576 ( \4708 , \4568 , \4586 );
and \U$4577 ( \4709 , \4554 , \4586 );
or \U$4578 ( \4710 , \4707 , \4708 , \4709 );
xor \U$4579 ( \4711 , \4706 , \4710 );
xor \U$4580 ( \4712 , \4697 , \4711 );
xor \U$4581 ( \4713 , \4688 , \4712 );
and \U$4582 ( \4714 , \4511 , \4515 );
and \U$4583 ( \4715 , \4515 , \4520 );
and \U$4584 ( \4716 , \4511 , \4520 );
or \U$4585 ( \4717 , \4714 , \4715 , \4716 );
and \U$4586 ( \4718 , \4535 , \4549 );
and \U$4587 ( \4719 , \4549 , \4587 );
and \U$4588 ( \4720 , \4535 , \4587 );
or \U$4589 ( \4721 , \4718 , \4719 , \4720 );
xor \U$4590 ( \4722 , \4717 , \4721 );
and \U$4591 ( \4723 , \4593 , \4637 );
and \U$4592 ( \4724 , \4637 , \4668 );
and \U$4593 ( \4725 , \4593 , \4668 );
or \U$4594 ( \4726 , \4723 , \4724 , \4725 );
xor \U$4595 ( \4727 , \4722 , \4726 );
and \U$4596 ( \4728 , \4611 , \4615 );
and \U$4597 ( \4729 , \4615 , \4620 );
and \U$4598 ( \4730 , \4611 , \4620 );
or \U$4599 ( \4731 , \4728 , \4729 , \4730 );
and \U$4600 ( \4732 , \4642 , \4646 );
and \U$4601 ( \4733 , \4646 , \4651 );
and \U$4602 ( \4734 , \4642 , \4651 );
or \U$4603 ( \4735 , \4732 , \4733 , \4734 );
xor \U$4604 ( \4736 , \4731 , \4735 );
and \U$4605 ( \4737 , \4657 , \4661 );
and \U$4606 ( \4738 , \4661 , \4666 );
and \U$4607 ( \4739 , \4657 , \4666 );
or \U$4608 ( \4740 , \4737 , \4738 , \4739 );
xor \U$4609 ( \4741 , \4736 , \4740 );
and \U$4610 ( \4742 , \4607 , \4621 );
and \U$4611 ( \4743 , \4621 , \4636 );
and \U$4612 ( \4744 , \4607 , \4636 );
or \U$4613 ( \4745 , \4742 , \4743 , \4744 );
and \U$4614 ( \4746 , \4652 , \4667 );
xor \U$4615 ( \4747 , \4745 , \4746 );
and \U$4616 ( \4748 , \4654 , \183 );
buf \U$4617 ( \4749 , RIb55e7e8_86);
and \U$4618 ( \4750 , \4749 , \180 );
nor \U$4619 ( \4751 , \4748 , \4750 );
xnor \U$4620 ( \4752 , \4751 , \179 );
and \U$4621 ( \4753 , \4160 , \195 );
and \U$4622 ( \4754 , \4364 , \193 );
nor \U$4623 ( \4755 , \4753 , \4754 );
xnor \U$4624 ( \4756 , \4755 , \202 );
xor \U$4625 ( \4757 , \4752 , \4756 );
buf \U$4626 ( \4758 , RIb560660_21);
buf \U$4627 ( \4759 , RIb5605e8_22);
and \U$4628 ( \4760 , \4759 , \4373 );
not \U$4629 ( \4761 , \4760 );
and \U$4630 ( \4762 , \4758 , \4761 );
xor \U$4631 ( \4763 , \4757 , \4762 );
and \U$4632 ( \4764 , \2757 , \141 );
and \U$4633 ( \4765 , \2826 , \139 );
nor \U$4634 ( \4766 , \4764 , \4765 );
xnor \U$4635 ( \4767 , \4766 , \148 );
and \U$4636 ( \4768 , \2366 , \156 );
and \U$4637 ( \4769 , \2521 , \154 );
nor \U$4638 ( \4770 , \4768 , \4769 );
xnor \U$4639 ( \4771 , \4770 , \163 );
xor \U$4640 ( \4772 , \4767 , \4771 );
and \U$4641 ( \4773 , \2090 , \296 );
and \U$4642 ( \4774 , \2182 , \168 );
nor \U$4643 ( \4775 , \4773 , \4774 );
xnor \U$4644 ( \4776 , \4775 , \173 );
xor \U$4645 ( \4777 , \4772 , \4776 );
xor \U$4646 ( \4778 , \4763 , \4777 );
and \U$4647 ( \4779 , \3736 , \215 );
and \U$4648 ( \4780 , \3912 , \213 );
nor \U$4649 ( \4781 , \4779 , \4780 );
xnor \U$4650 ( \4782 , \4781 , \222 );
and \U$4651 ( \4783 , \3395 , \230 );
and \U$4652 ( \4784 , \3646 , \228 );
nor \U$4653 ( \4785 , \4783 , \4784 );
xnor \U$4654 ( \4786 , \4785 , \237 );
xor \U$4655 ( \4787 , \4782 , \4786 );
and \U$4656 ( \4788 , \3037 , \245 );
and \U$4657 ( \4789 , \3143 , \243 );
nor \U$4658 ( \4790 , \4788 , \4789 );
xnor \U$4659 ( \4791 , \4790 , \252 );
xor \U$4660 ( \4792 , \4787 , \4791 );
xor \U$4661 ( \4793 , \4778 , \4792 );
xor \U$4662 ( \4794 , \4747 , \4793 );
xor \U$4663 ( \4795 , \4741 , \4794 );
and \U$4664 ( \4796 , \4597 , \4601 );
and \U$4665 ( \4797 , \4601 , \4606 );
and \U$4666 ( \4798 , \4597 , \4606 );
or \U$4667 ( \4799 , \4796 , \4797 , \4798 );
and \U$4668 ( \4800 , \4558 , \4562 );
and \U$4669 ( \4801 , \4562 , \4567 );
and \U$4670 ( \4802 , \4558 , \4567 );
or \U$4671 ( \4803 , \4800 , \4801 , \4802 );
xor \U$4672 ( \4804 , \4799 , \4803 );
and \U$4673 ( \4805 , \4626 , \4630 );
and \U$4674 ( \4806 , \4630 , \4635 );
and \U$4675 ( \4807 , \4626 , \4635 );
or \U$4676 ( \4808 , \4805 , \4806 , \4807 );
xor \U$4677 ( \4809 , \4804 , \4808 );
and \U$4678 ( \4810 , \178 , \2400 );
and \U$4679 ( \4811 , \185 , \2246 );
nor \U$4680 ( \4812 , \4810 , \4811 );
xnor \U$4681 ( \4813 , \4812 , \2195 );
and \U$4682 ( \4814 , \189 , \2669 );
and \U$4683 ( \4815 , \197 , \2538 );
nor \U$4684 ( \4816 , \4814 , \4815 );
xnor \U$4685 ( \4817 , \4816 , \2534 );
xor \U$4686 ( \4818 , \4813 , \4817 );
and \U$4687 ( \4819 , \209 , \3103 );
and \U$4688 ( \4820 , \217 , \2934 );
nor \U$4689 ( \4821 , \4819 , \4820 );
xnor \U$4690 ( \4822 , \4821 , \2839 );
xor \U$4691 ( \4823 , \4818 , \4822 );
and \U$4692 ( \4824 , \1802 , \438 );
and \U$4693 ( \4825 , \1948 , \336 );
nor \U$4694 ( \4826 , \4824 , \4825 );
xnor \U$4695 ( \4827 , \4826 , \320 );
and \U$4696 ( \4828 , \1601 , \1086 );
and \U$4697 ( \4829 , \1684 , \508 );
nor \U$4698 ( \4830 , \4828 , \4829 );
xnor \U$4699 ( \4831 , \4830 , \487 );
xor \U$4700 ( \4832 , \4827 , \4831 );
and \U$4701 ( \4833 , \1333 , \1301 );
and \U$4702 ( \4834 , \1484 , \1246 );
nor \U$4703 ( \4835 , \4833 , \4834 );
xnor \U$4704 ( \4836 , \4835 , \1205 );
xor \U$4705 ( \4837 , \4832 , \4836 );
xor \U$4706 ( \4838 , \4823 , \4837 );
and \U$4707 ( \4839 , \1147 , \1578 );
and \U$4708 ( \4840 , \1192 , \1431 );
nor \U$4709 ( \4841 , \4839 , \4840 );
xnor \U$4710 ( \4842 , \4841 , \1436 );
and \U$4711 ( \4843 , \412 , \1824 );
and \U$4712 ( \4844 , \474 , \1739 );
nor \U$4713 ( \4845 , \4843 , \4844 );
xnor \U$4714 ( \4846 , \4845 , \1697 );
xor \U$4715 ( \4847 , \4842 , \4846 );
and \U$4716 ( \4848 , \261 , \2121 );
and \U$4717 ( \4849 , \307 , \2008 );
nor \U$4718 ( \4850 , \4848 , \4849 );
xnor \U$4719 ( \4851 , \4850 , \1961 );
xor \U$4720 ( \4852 , \4847 , \4851 );
xor \U$4721 ( \4853 , \4838 , \4852 );
xor \U$4722 ( \4854 , \4809 , \4853 );
and \U$4723 ( \4855 , \4573 , \4577 );
and \U$4724 ( \4856 , \4577 , \4585 );
and \U$4725 ( \4857 , \4573 , \4585 );
or \U$4726 ( \4858 , \4855 , \4856 , \4857 );
and \U$4727 ( \4859 , \224 , \3357 );
and \U$4728 ( \4860 , \232 , \3255 );
nor \U$4729 ( \4861 , \4859 , \4860 );
xnor \U$4730 ( \4862 , \4861 , \3156 );
and \U$4731 ( \4863 , \240 , \3813 );
and \U$4732 ( \4864 , \247 , \3557 );
nor \U$4733 ( \4865 , \4863 , \4864 );
xnor \U$4734 ( \4866 , \4865 , \3562 );
xor \U$4735 ( \4867 , \4862 , \4866 );
and \U$4736 ( \4868 , \134 , \4132 );
and \U$4737 ( \4869 , \143 , \4012 );
nor \U$4738 ( \4870 , \4868 , \4869 );
xnor \U$4739 ( \4871 , \4870 , \3925 );
xor \U$4740 ( \4872 , \4867 , \4871 );
xor \U$4741 ( \4873 , \4858 , \4872 );
and \U$4742 ( \4874 , \150 , \4581 );
and \U$4743 ( \4875 , \158 , \4424 );
nor \U$4744 ( \4876 , \4874 , \4875 );
xnor \U$4745 ( \4877 , \4876 , \4377 );
xor \U$4746 ( \4878 , \4759 , \4373 );
nand \U$4747 ( \4879 , \166 , \4878 );
xnor \U$4748 ( \4880 , \4879 , \4762 );
xor \U$4749 ( \4881 , \4877 , \4880 );
xor \U$4750 ( \4882 , \4873 , \4881 );
xor \U$4751 ( \4883 , \4854 , \4882 );
xor \U$4752 ( \4884 , \4795 , \4883 );
xor \U$4753 ( \4885 , \4727 , \4884 );
xor \U$4754 ( \4886 , \4713 , \4885 );
xor \U$4755 ( \4887 , \4684 , \4886 );
and \U$4756 ( \4888 , \4473 , \4497 );
and \U$4757 ( \4889 , \4497 , \4671 );
and \U$4758 ( \4890 , \4473 , \4671 );
or \U$4759 ( \4891 , \4888 , \4889 , \4890 );
xor \U$4760 ( \4892 , \4887 , \4891 );
and \U$4761 ( \4893 , \4672 , \4673 );
and \U$4762 ( \4894 , \4674 , \4677 );
or \U$4763 ( \4895 , \4893 , \4894 );
xor \U$4764 ( \4896 , \4892 , \4895 );
buf \U$4765 ( \4897 , \4896 );
buf \U$4766 ( \4898 , \4897 );
and \U$4767 ( \4899 , \4688 , \4712 );
and \U$4768 ( \4900 , \4712 , \4885 );
and \U$4769 ( \4901 , \4688 , \4885 );
or \U$4770 ( \4902 , \4899 , \4900 , \4901 );
and \U$4771 ( \4903 , \4717 , \4721 );
and \U$4772 ( \4904 , \4721 , \4726 );
and \U$4773 ( \4905 , \4717 , \4726 );
or \U$4774 ( \4906 , \4903 , \4904 , \4905 );
and \U$4775 ( \4907 , \4741 , \4794 );
and \U$4776 ( \4908 , \4794 , \4883 );
and \U$4777 ( \4909 , \4741 , \4883 );
or \U$4778 ( \4910 , \4907 , \4908 , \4909 );
xor \U$4779 ( \4911 , \4906 , \4910 );
and \U$4780 ( \4912 , \4763 , \4777 );
and \U$4781 ( \4913 , \4777 , \4792 );
and \U$4782 ( \4914 , \4763 , \4792 );
or \U$4783 ( \4915 , \4912 , \4913 , \4914 );
and \U$4784 ( \4916 , \4823 , \4837 );
and \U$4785 ( \4917 , \4837 , \4852 );
and \U$4786 ( \4918 , \4823 , \4852 );
or \U$4787 ( \4919 , \4916 , \4917 , \4918 );
xor \U$4788 ( \4920 , \4915 , \4919 );
and \U$4789 ( \4921 , \4749 , \183 );
buf \U$4790 ( \4922 , RIb55e860_85);
and \U$4791 ( \4923 , \4922 , \180 );
nor \U$4792 ( \4924 , \4921 , \4923 );
xnor \U$4793 ( \4925 , \4924 , \179 );
and \U$4794 ( \4926 , \4364 , \195 );
and \U$4795 ( \4927 , \4654 , \193 );
nor \U$4796 ( \4928 , \4926 , \4927 );
xnor \U$4797 ( \4929 , \4928 , \202 );
xor \U$4798 ( \4930 , \4925 , \4929 );
and \U$4799 ( \4931 , \3912 , \215 );
and \U$4800 ( \4932 , \4160 , \213 );
nor \U$4801 ( \4933 , \4931 , \4932 );
xnor \U$4802 ( \4934 , \4933 , \222 );
xor \U$4803 ( \4935 , \4930 , \4934 );
xor \U$4804 ( \4936 , \4920 , \4935 );
xor \U$4805 ( \4937 , \4911 , \4936 );
xor \U$4806 ( \4938 , \4902 , \4937 );
and \U$4807 ( \4939 , \4692 , \4696 );
and \U$4808 ( \4940 , \4696 , \4711 );
and \U$4809 ( \4941 , \4692 , \4711 );
or \U$4810 ( \4942 , \4939 , \4940 , \4941 );
and \U$4811 ( \4943 , \4727 , \4884 );
xor \U$4812 ( \4944 , \4942 , \4943 );
and \U$4813 ( \4945 , \4799 , \4803 );
and \U$4814 ( \4946 , \4803 , \4808 );
and \U$4815 ( \4947 , \4799 , \4808 );
or \U$4816 ( \4948 , \4945 , \4946 , \4947 );
and \U$4817 ( \4949 , \4731 , \4735 );
and \U$4818 ( \4950 , \4735 , \4740 );
and \U$4819 ( \4951 , \4731 , \4740 );
or \U$4820 ( \4952 , \4949 , \4950 , \4951 );
xor \U$4821 ( \4953 , \4948 , \4952 );
and \U$4822 ( \4954 , \4858 , \4872 );
and \U$4823 ( \4955 , \4872 , \4881 );
and \U$4824 ( \4956 , \4858 , \4881 );
or \U$4825 ( \4957 , \4954 , \4955 , \4956 );
xor \U$4826 ( \4958 , \4953 , \4957 );
and \U$4827 ( \4959 , \4701 , \4705 );
and \U$4828 ( \4960 , \4705 , \4710 );
and \U$4829 ( \4961 , \4701 , \4710 );
or \U$4830 ( \4962 , \4959 , \4960 , \4961 );
and \U$4831 ( \4963 , \4745 , \4746 );
and \U$4832 ( \4964 , \4746 , \4793 );
and \U$4833 ( \4965 , \4745 , \4793 );
or \U$4834 ( \4966 , \4963 , \4964 , \4965 );
xor \U$4835 ( \4967 , \4962 , \4966 );
and \U$4836 ( \4968 , \4809 , \4853 );
and \U$4837 ( \4969 , \4853 , \4882 );
and \U$4838 ( \4970 , \4809 , \4882 );
or \U$4839 ( \4971 , \4968 , \4969 , \4970 );
xor \U$4840 ( \4972 , \4967 , \4971 );
xor \U$4841 ( \4973 , \4958 , \4972 );
and \U$4842 ( \4974 , \4813 , \4817 );
and \U$4843 ( \4975 , \4817 , \4822 );
and \U$4844 ( \4976 , \4813 , \4822 );
or \U$4845 ( \4977 , \4974 , \4975 , \4976 );
and \U$4846 ( \4978 , \4827 , \4831 );
and \U$4847 ( \4979 , \4831 , \4836 );
and \U$4848 ( \4980 , \4827 , \4836 );
or \U$4849 ( \4981 , \4978 , \4979 , \4980 );
xor \U$4850 ( \4982 , \4977 , \4981 );
and \U$4851 ( \4983 , \4842 , \4846 );
and \U$4852 ( \4984 , \4846 , \4851 );
and \U$4853 ( \4985 , \4842 , \4851 );
or \U$4854 ( \4986 , \4983 , \4984 , \4985 );
xor \U$4855 ( \4987 , \4982 , \4986 );
and \U$4856 ( \4988 , \4752 , \4756 );
and \U$4857 ( \4989 , \4756 , \4762 );
and \U$4858 ( \4990 , \4752 , \4762 );
or \U$4859 ( \4991 , \4988 , \4989 , \4990 );
and \U$4860 ( \4992 , \4767 , \4771 );
and \U$4861 ( \4993 , \4771 , \4776 );
and \U$4862 ( \4994 , \4767 , \4776 );
or \U$4863 ( \4995 , \4992 , \4993 , \4994 );
xor \U$4864 ( \4996 , \4991 , \4995 );
and \U$4865 ( \4997 , \4782 , \4786 );
and \U$4866 ( \4998 , \4786 , \4791 );
and \U$4867 ( \4999 , \4782 , \4791 );
or \U$4868 ( \5000 , \4997 , \4998 , \4999 );
xor \U$4869 ( \5001 , \4996 , \5000 );
xor \U$4870 ( \5002 , \4987 , \5001 );
and \U$4871 ( \5003 , \4862 , \4866 );
and \U$4872 ( \5004 , \4866 , \4871 );
and \U$4873 ( \5005 , \4862 , \4871 );
or \U$4874 ( \5006 , \5003 , \5004 , \5005 );
and \U$4875 ( \5007 , \4877 , \4880 );
xor \U$4876 ( \5008 , \5006 , \5007 );
xor \U$4877 ( \5009 , \4758 , \4759 );
not \U$4878 ( \5010 , \4878 );
and \U$4879 ( \5011 , \5009 , \5010 );
and \U$4880 ( \5012 , \166 , \5011 );
and \U$4881 ( \5013 , \150 , \4878 );
nor \U$4882 ( \5014 , \5012 , \5013 );
xnor \U$4883 ( \5015 , \5014 , \4762 );
xor \U$4884 ( \5016 , \5008 , \5015 );
and \U$4885 ( \5017 , \3646 , \230 );
and \U$4886 ( \5018 , \3736 , \228 );
nor \U$4887 ( \5019 , \5017 , \5018 );
xnor \U$4888 ( \5020 , \5019 , \237 );
and \U$4889 ( \5021 , \3143 , \245 );
and \U$4890 ( \5022 , \3395 , \243 );
nor \U$4891 ( \5023 , \5021 , \5022 );
xnor \U$4892 ( \5024 , \5023 , \252 );
xor \U$4893 ( \5025 , \5020 , \5024 );
and \U$4894 ( \5026 , \2826 , \141 );
and \U$4895 ( \5027 , \3037 , \139 );
nor \U$4896 ( \5028 , \5026 , \5027 );
xnor \U$4897 ( \5029 , \5028 , \148 );
xor \U$4898 ( \5030 , \5025 , \5029 );
and \U$4899 ( \5031 , \1684 , \1086 );
and \U$4900 ( \5032 , \1802 , \508 );
nor \U$4901 ( \5033 , \5031 , \5032 );
xnor \U$4902 ( \5034 , \5033 , \487 );
and \U$4903 ( \5035 , \1484 , \1301 );
and \U$4904 ( \5036 , \1601 , \1246 );
nor \U$4905 ( \5037 , \5035 , \5036 );
xnor \U$4906 ( \5038 , \5037 , \1205 );
xor \U$4907 ( \5039 , \5034 , \5038 );
and \U$4908 ( \5040 , \1192 , \1578 );
and \U$4909 ( \5041 , \1333 , \1431 );
nor \U$4910 ( \5042 , \5040 , \5041 );
xnor \U$4911 ( \5043 , \5042 , \1436 );
xor \U$4912 ( \5044 , \5039 , \5043 );
xor \U$4913 ( \5045 , \5030 , \5044 );
and \U$4914 ( \5046 , \2521 , \156 );
and \U$4915 ( \5047 , \2757 , \154 );
nor \U$4916 ( \5048 , \5046 , \5047 );
xnor \U$4917 ( \5049 , \5048 , \163 );
and \U$4918 ( \5050 , \2182 , \296 );
and \U$4919 ( \5051 , \2366 , \168 );
nor \U$4920 ( \5052 , \5050 , \5051 );
xnor \U$4921 ( \5053 , \5052 , \173 );
xor \U$4922 ( \5054 , \5049 , \5053 );
and \U$4923 ( \5055 , \1948 , \438 );
and \U$4924 ( \5056 , \2090 , \336 );
nor \U$4925 ( \5057 , \5055 , \5056 );
xnor \U$4926 ( \5058 , \5057 , \320 );
xor \U$4927 ( \5059 , \5054 , \5058 );
xor \U$4928 ( \5060 , \5045 , \5059 );
xor \U$4929 ( \5061 , \5016 , \5060 );
and \U$4930 ( \5062 , \474 , \1824 );
and \U$4931 ( \5063 , \1147 , \1739 );
nor \U$4932 ( \5064 , \5062 , \5063 );
xnor \U$4933 ( \5065 , \5064 , \1697 );
and \U$4934 ( \5066 , \307 , \2121 );
and \U$4935 ( \5067 , \412 , \2008 );
nor \U$4936 ( \5068 , \5066 , \5067 );
xnor \U$4937 ( \5069 , \5068 , \1961 );
xor \U$4938 ( \5070 , \5065 , \5069 );
and \U$4939 ( \5071 , \185 , \2400 );
and \U$4940 ( \5072 , \261 , \2246 );
nor \U$4941 ( \5073 , \5071 , \5072 );
xnor \U$4942 ( \5074 , \5073 , \2195 );
xor \U$4943 ( \5075 , \5070 , \5074 );
and \U$4944 ( \5076 , \247 , \3813 );
and \U$4945 ( \5077 , \224 , \3557 );
nor \U$4946 ( \5078 , \5076 , \5077 );
xnor \U$4947 ( \5079 , \5078 , \3562 );
and \U$4948 ( \5080 , \143 , \4132 );
and \U$4949 ( \5081 , \240 , \4012 );
nor \U$4950 ( \5082 , \5080 , \5081 );
xnor \U$4951 ( \5083 , \5082 , \3925 );
xor \U$4952 ( \5084 , \5079 , \5083 );
and \U$4953 ( \5085 , \158 , \4581 );
and \U$4954 ( \5086 , \134 , \4424 );
nor \U$4955 ( \5087 , \5085 , \5086 );
xnor \U$4956 ( \5088 , \5087 , \4377 );
xor \U$4957 ( \5089 , \5084 , \5088 );
xor \U$4958 ( \5090 , \5075 , \5089 );
and \U$4959 ( \5091 , \197 , \2669 );
and \U$4960 ( \5092 , \178 , \2538 );
nor \U$4961 ( \5093 , \5091 , \5092 );
xnor \U$4962 ( \5094 , \5093 , \2534 );
and \U$4963 ( \5095 , \217 , \3103 );
and \U$4964 ( \5096 , \189 , \2934 );
nor \U$4965 ( \5097 , \5095 , \5096 );
xnor \U$4966 ( \5098 , \5097 , \2839 );
xor \U$4967 ( \5099 , \5094 , \5098 );
and \U$4968 ( \5100 , \232 , \3357 );
and \U$4969 ( \5101 , \209 , \3255 );
nor \U$4970 ( \5102 , \5100 , \5101 );
xnor \U$4971 ( \5103 , \5102 , \3156 );
xor \U$4972 ( \5104 , \5099 , \5103 );
xor \U$4973 ( \5105 , \5090 , \5104 );
xor \U$4974 ( \5106 , \5061 , \5105 );
xor \U$4975 ( \5107 , \5002 , \5106 );
xor \U$4976 ( \5108 , \4973 , \5107 );
xor \U$4977 ( \5109 , \4944 , \5108 );
xor \U$4978 ( \5110 , \4938 , \5109 );
and \U$4979 ( \5111 , \4684 , \4886 );
xor \U$4980 ( \5112 , \5110 , \5111 );
and \U$4981 ( \5113 , \4887 , \4891 );
and \U$4982 ( \5114 , \4892 , \4895 );
or \U$4983 ( \5115 , \5113 , \5114 );
xor \U$4984 ( \5116 , \5112 , \5115 );
buf \U$4985 ( \5117 , \5116 );
buf \U$4986 ( \5118 , \5117 );
and \U$4987 ( \5119 , \4942 , \4943 );
and \U$4988 ( \5120 , \4943 , \5108 );
and \U$4989 ( \5121 , \4942 , \5108 );
or \U$4990 ( \5122 , \5119 , \5120 , \5121 );
and \U$4991 ( \5123 , \4906 , \4910 );
and \U$4992 ( \5124 , \4910 , \4936 );
and \U$4993 ( \5125 , \4906 , \4936 );
or \U$4994 ( \5126 , \5123 , \5124 , \5125 );
and \U$4995 ( \5127 , \4958 , \4972 );
and \U$4996 ( \5128 , \4972 , \5107 );
and \U$4997 ( \5129 , \4958 , \5107 );
or \U$4998 ( \5130 , \5127 , \5128 , \5129 );
xor \U$4999 ( \5131 , \5126 , \5130 );
and \U$5000 ( \5132 , \4925 , \4929 );
and \U$5001 ( \5133 , \4929 , \4934 );
and \U$5002 ( \5134 , \4925 , \4934 );
or \U$5003 ( \5135 , \5132 , \5133 , \5134 );
and \U$5004 ( \5136 , \5020 , \5024 );
and \U$5005 ( \5137 , \5024 , \5029 );
and \U$5006 ( \5138 , \5020 , \5029 );
or \U$5007 ( \5139 , \5136 , \5137 , \5138 );
xor \U$5008 ( \5140 , \5135 , \5139 );
and \U$5009 ( \5141 , \5049 , \5053 );
and \U$5010 ( \5142 , \5053 , \5058 );
and \U$5011 ( \5143 , \5049 , \5058 );
or \U$5012 ( \5144 , \5141 , \5142 , \5143 );
xor \U$5013 ( \5145 , \5140 , \5144 );
and \U$5014 ( \5146 , \5030 , \5044 );
and \U$5015 ( \5147 , \5044 , \5059 );
and \U$5016 ( \5148 , \5030 , \5059 );
or \U$5017 ( \5149 , \5146 , \5147 , \5148 );
and \U$5018 ( \5150 , \5075 , \5089 );
and \U$5019 ( \5151 , \5089 , \5104 );
and \U$5020 ( \5152 , \5075 , \5104 );
or \U$5021 ( \5153 , \5150 , \5151 , \5152 );
xor \U$5022 ( \5154 , \5149 , \5153 );
and \U$5023 ( \5155 , \4922 , \183 );
buf \U$5024 ( \5156 , RIb55e8d8_84);
and \U$5025 ( \5157 , \5156 , \180 );
nor \U$5026 ( \5158 , \5155 , \5157 );
xnor \U$5027 ( \5159 , \5158 , \179 );
and \U$5028 ( \5160 , \4654 , \195 );
and \U$5029 ( \5161 , \4749 , \193 );
nor \U$5030 ( \5162 , \5160 , \5161 );
xnor \U$5031 ( \5163 , \5162 , \202 );
xor \U$5032 ( \5164 , \5159 , \5163 );
buf \U$5033 ( \5165 , RIb560750_19);
buf \U$5034 ( \5166 , RIb5606d8_20);
and \U$5035 ( \5167 , \5166 , \4758 );
not \U$5036 ( \5168 , \5167 );
and \U$5037 ( \5169 , \5165 , \5168 );
xor \U$5038 ( \5170 , \5164 , \5169 );
and \U$5039 ( \5171 , \3037 , \141 );
and \U$5040 ( \5172 , \3143 , \139 );
nor \U$5041 ( \5173 , \5171 , \5172 );
xnor \U$5042 ( \5174 , \5173 , \148 );
and \U$5043 ( \5175 , \2757 , \156 );
and \U$5044 ( \5176 , \2826 , \154 );
nor \U$5045 ( \5177 , \5175 , \5176 );
xnor \U$5046 ( \5178 , \5177 , \163 );
xor \U$5047 ( \5179 , \5174 , \5178 );
and \U$5048 ( \5180 , \2366 , \296 );
and \U$5049 ( \5181 , \2521 , \168 );
nor \U$5050 ( \5182 , \5180 , \5181 );
xnor \U$5051 ( \5183 , \5182 , \173 );
xor \U$5052 ( \5184 , \5179 , \5183 );
xor \U$5053 ( \5185 , \5170 , \5184 );
and \U$5054 ( \5186 , \4160 , \215 );
and \U$5055 ( \5187 , \4364 , \213 );
nor \U$5056 ( \5188 , \5186 , \5187 );
xnor \U$5057 ( \5189 , \5188 , \222 );
and \U$5058 ( \5190 , \3736 , \230 );
and \U$5059 ( \5191 , \3912 , \228 );
nor \U$5060 ( \5192 , \5190 , \5191 );
xnor \U$5061 ( \5193 , \5192 , \237 );
xor \U$5062 ( \5194 , \5189 , \5193 );
and \U$5063 ( \5195 , \3395 , \245 );
and \U$5064 ( \5196 , \3646 , \243 );
nor \U$5065 ( \5197 , \5195 , \5196 );
xnor \U$5066 ( \5198 , \5197 , \252 );
xor \U$5067 ( \5199 , \5194 , \5198 );
xor \U$5068 ( \5200 , \5185 , \5199 );
xor \U$5069 ( \5201 , \5154 , \5200 );
xor \U$5070 ( \5202 , \5145 , \5201 );
and \U$5071 ( \5203 , \5065 , \5069 );
and \U$5072 ( \5204 , \5069 , \5074 );
and \U$5073 ( \5205 , \5065 , \5074 );
or \U$5074 ( \5206 , \5203 , \5204 , \5205 );
and \U$5075 ( \5207 , \5094 , \5098 );
and \U$5076 ( \5208 , \5098 , \5103 );
and \U$5077 ( \5209 , \5094 , \5103 );
or \U$5078 ( \5210 , \5207 , \5208 , \5209 );
xor \U$5079 ( \5211 , \5206 , \5210 );
and \U$5080 ( \5212 , \5034 , \5038 );
and \U$5081 ( \5213 , \5038 , \5043 );
and \U$5082 ( \5214 , \5034 , \5043 );
or \U$5083 ( \5215 , \5212 , \5213 , \5214 );
xor \U$5084 ( \5216 , \5211 , \5215 );
and \U$5085 ( \5217 , \2090 , \438 );
and \U$5086 ( \5218 , \2182 , \336 );
nor \U$5087 ( \5219 , \5217 , \5218 );
xnor \U$5088 ( \5220 , \5219 , \320 );
and \U$5089 ( \5221 , \1802 , \1086 );
and \U$5090 ( \5222 , \1948 , \508 );
nor \U$5091 ( \5223 , \5221 , \5222 );
xnor \U$5092 ( \5224 , \5223 , \487 );
xor \U$5093 ( \5225 , \5220 , \5224 );
and \U$5094 ( \5226 , \1601 , \1301 );
and \U$5095 ( \5227 , \1684 , \1246 );
nor \U$5096 ( \5228 , \5226 , \5227 );
xnor \U$5097 ( \5229 , \5228 , \1205 );
xor \U$5098 ( \5230 , \5225 , \5229 );
and \U$5099 ( \5231 , \1333 , \1578 );
and \U$5100 ( \5232 , \1484 , \1431 );
nor \U$5101 ( \5233 , \5231 , \5232 );
xnor \U$5102 ( \5234 , \5233 , \1436 );
and \U$5103 ( \5235 , \1147 , \1824 );
and \U$5104 ( \5236 , \1192 , \1739 );
nor \U$5105 ( \5237 , \5235 , \5236 );
xnor \U$5106 ( \5238 , \5237 , \1697 );
xor \U$5107 ( \5239 , \5234 , \5238 );
and \U$5108 ( \5240 , \412 , \2121 );
and \U$5109 ( \5241 , \474 , \2008 );
nor \U$5110 ( \5242 , \5240 , \5241 );
xnor \U$5111 ( \5243 , \5242 , \1961 );
xor \U$5112 ( \5244 , \5239 , \5243 );
xor \U$5113 ( \5245 , \5230 , \5244 );
and \U$5114 ( \5246 , \261 , \2400 );
and \U$5115 ( \5247 , \307 , \2246 );
nor \U$5116 ( \5248 , \5246 , \5247 );
xnor \U$5117 ( \5249 , \5248 , \2195 );
and \U$5118 ( \5250 , \178 , \2669 );
and \U$5119 ( \5251 , \185 , \2538 );
nor \U$5120 ( \5252 , \5250 , \5251 );
xnor \U$5121 ( \5253 , \5252 , \2534 );
xor \U$5122 ( \5254 , \5249 , \5253 );
and \U$5123 ( \5255 , \189 , \3103 );
and \U$5124 ( \5256 , \197 , \2934 );
nor \U$5125 ( \5257 , \5255 , \5256 );
xnor \U$5126 ( \5258 , \5257 , \2839 );
xor \U$5127 ( \5259 , \5254 , \5258 );
xor \U$5128 ( \5260 , \5245 , \5259 );
xor \U$5129 ( \5261 , \5216 , \5260 );
and \U$5130 ( \5262 , \5079 , \5083 );
and \U$5131 ( \5263 , \5083 , \5088 );
and \U$5132 ( \5264 , \5079 , \5088 );
or \U$5133 ( \5265 , \5262 , \5263 , \5264 );
and \U$5134 ( \5266 , \134 , \4581 );
and \U$5135 ( \5267 , \143 , \4424 );
nor \U$5136 ( \5268 , \5266 , \5267 );
xnor \U$5137 ( \5269 , \5268 , \4377 );
and \U$5138 ( \5270 , \150 , \5011 );
and \U$5139 ( \5271 , \158 , \4878 );
nor \U$5140 ( \5272 , \5270 , \5271 );
xnor \U$5141 ( \5273 , \5272 , \4762 );
xor \U$5142 ( \5274 , \5269 , \5273 );
xor \U$5143 ( \5275 , \5166 , \4758 );
nand \U$5144 ( \5276 , \166 , \5275 );
xnor \U$5145 ( \5277 , \5276 , \5169 );
xor \U$5146 ( \5278 , \5274 , \5277 );
xor \U$5147 ( \5279 , \5265 , \5278 );
and \U$5148 ( \5280 , \209 , \3357 );
and \U$5149 ( \5281 , \217 , \3255 );
nor \U$5150 ( \5282 , \5280 , \5281 );
xnor \U$5151 ( \5283 , \5282 , \3156 );
and \U$5152 ( \5284 , \224 , \3813 );
and \U$5153 ( \5285 , \232 , \3557 );
nor \U$5154 ( \5286 , \5284 , \5285 );
xnor \U$5155 ( \5287 , \5286 , \3562 );
xor \U$5156 ( \5288 , \5283 , \5287 );
and \U$5157 ( \5289 , \240 , \4132 );
and \U$5158 ( \5290 , \247 , \4012 );
nor \U$5159 ( \5291 , \5289 , \5290 );
xnor \U$5160 ( \5292 , \5291 , \3925 );
xor \U$5161 ( \5293 , \5288 , \5292 );
xor \U$5162 ( \5294 , \5279 , \5293 );
xor \U$5163 ( \5295 , \5261 , \5294 );
xor \U$5164 ( \5296 , \5202 , \5295 );
xor \U$5165 ( \5297 , \5131 , \5296 );
xor \U$5166 ( \5298 , \5122 , \5297 );
and \U$5167 ( \5299 , \4948 , \4952 );
and \U$5168 ( \5300 , \4952 , \4957 );
and \U$5169 ( \5301 , \4948 , \4957 );
or \U$5170 ( \5302 , \5299 , \5300 , \5301 );
and \U$5171 ( \5303 , \4915 , \4919 );
and \U$5172 ( \5304 , \4919 , \4935 );
and \U$5173 ( \5305 , \4915 , \4935 );
or \U$5174 ( \5306 , \5303 , \5304 , \5305 );
xor \U$5175 ( \5307 , \5302 , \5306 );
and \U$5176 ( \5308 , \5016 , \5060 );
and \U$5177 ( \5309 , \5060 , \5105 );
and \U$5178 ( \5310 , \5016 , \5105 );
or \U$5179 ( \5311 , \5308 , \5309 , \5310 );
xor \U$5180 ( \5312 , \5307 , \5311 );
and \U$5181 ( \5313 , \4962 , \4966 );
and \U$5182 ( \5314 , \4966 , \4971 );
and \U$5183 ( \5315 , \4962 , \4971 );
or \U$5184 ( \5316 , \5313 , \5314 , \5315 );
and \U$5185 ( \5317 , \4987 , \5001 );
and \U$5186 ( \5318 , \5001 , \5106 );
and \U$5187 ( \5319 , \4987 , \5106 );
or \U$5188 ( \5320 , \5317 , \5318 , \5319 );
xor \U$5189 ( \5321 , \5316 , \5320 );
and \U$5190 ( \5322 , \4977 , \4981 );
and \U$5191 ( \5323 , \4981 , \4986 );
and \U$5192 ( \5324 , \4977 , \4986 );
or \U$5193 ( \5325 , \5322 , \5323 , \5324 );
and \U$5194 ( \5326 , \4991 , \4995 );
and \U$5195 ( \5327 , \4995 , \5000 );
and \U$5196 ( \5328 , \4991 , \5000 );
or \U$5197 ( \5329 , \5326 , \5327 , \5328 );
xor \U$5198 ( \5330 , \5325 , \5329 );
and \U$5199 ( \5331 , \5006 , \5007 );
and \U$5200 ( \5332 , \5007 , \5015 );
and \U$5201 ( \5333 , \5006 , \5015 );
or \U$5202 ( \5334 , \5331 , \5332 , \5333 );
xor \U$5203 ( \5335 , \5330 , \5334 );
xor \U$5204 ( \5336 , \5321 , \5335 );
xor \U$5205 ( \5337 , \5312 , \5336 );
xor \U$5206 ( \5338 , \5298 , \5337 );
and \U$5207 ( \5339 , \4902 , \4937 );
and \U$5208 ( \5340 , \4937 , \5109 );
and \U$5209 ( \5341 , \4902 , \5109 );
or \U$5210 ( \5342 , \5339 , \5340 , \5341 );
xor \U$5211 ( \5343 , \5338 , \5342 );
and \U$5212 ( \5344 , \5110 , \5111 );
and \U$5213 ( \5345 , \5112 , \5115 );
or \U$5214 ( \5346 , \5344 , \5345 );
xor \U$5215 ( \5347 , \5343 , \5346 );
buf \U$5216 ( \5348 , \5347 );
buf \U$5217 ( \5349 , \5348 );
and \U$5218 ( \5350 , \5126 , \5130 );
and \U$5219 ( \5351 , \5130 , \5296 );
and \U$5220 ( \5352 , \5126 , \5296 );
or \U$5221 ( \5353 , \5350 , \5351 , \5352 );
and \U$5222 ( \5354 , \5312 , \5336 );
xor \U$5223 ( \5355 , \5353 , \5354 );
and \U$5224 ( \5356 , \5316 , \5320 );
and \U$5225 ( \5357 , \5320 , \5335 );
and \U$5226 ( \5358 , \5316 , \5335 );
or \U$5227 ( \5359 , \5356 , \5357 , \5358 );
and \U$5228 ( \5360 , \5302 , \5306 );
and \U$5229 ( \5361 , \5306 , \5311 );
and \U$5230 ( \5362 , \5302 , \5311 );
or \U$5231 ( \5363 , \5360 , \5361 , \5362 );
and \U$5232 ( \5364 , \5145 , \5201 );
and \U$5233 ( \5365 , \5201 , \5295 );
and \U$5234 ( \5366 , \5145 , \5295 );
or \U$5235 ( \5367 , \5364 , \5365 , \5366 );
xor \U$5236 ( \5368 , \5363 , \5367 );
and \U$5237 ( \5369 , \5135 , \5139 );
and \U$5238 ( \5370 , \5139 , \5144 );
and \U$5239 ( \5371 , \5135 , \5144 );
or \U$5240 ( \5372 , \5369 , \5370 , \5371 );
and \U$5241 ( \5373 , \5206 , \5210 );
and \U$5242 ( \5374 , \5210 , \5215 );
and \U$5243 ( \5375 , \5206 , \5215 );
or \U$5244 ( \5376 , \5373 , \5374 , \5375 );
xor \U$5245 ( \5377 , \5372 , \5376 );
and \U$5246 ( \5378 , \5265 , \5278 );
and \U$5247 ( \5379 , \5278 , \5293 );
and \U$5248 ( \5380 , \5265 , \5293 );
or \U$5249 ( \5381 , \5378 , \5379 , \5380 );
xor \U$5250 ( \5382 , \5377 , \5381 );
xor \U$5251 ( \5383 , \5368 , \5382 );
xor \U$5252 ( \5384 , \5359 , \5383 );
and \U$5253 ( \5385 , \5325 , \5329 );
and \U$5254 ( \5386 , \5329 , \5334 );
and \U$5255 ( \5387 , \5325 , \5334 );
or \U$5256 ( \5388 , \5385 , \5386 , \5387 );
and \U$5257 ( \5389 , \5149 , \5153 );
and \U$5258 ( \5390 , \5153 , \5200 );
and \U$5259 ( \5391 , \5149 , \5200 );
or \U$5260 ( \5392 , \5389 , \5390 , \5391 );
xor \U$5261 ( \5393 , \5388 , \5392 );
and \U$5262 ( \5394 , \5216 , \5260 );
and \U$5263 ( \5395 , \5260 , \5294 );
and \U$5264 ( \5396 , \5216 , \5294 );
or \U$5265 ( \5397 , \5394 , \5395 , \5396 );
xor \U$5266 ( \5398 , \5393 , \5397 );
and \U$5267 ( \5399 , \5159 , \5163 );
and \U$5268 ( \5400 , \5163 , \5169 );
and \U$5269 ( \5401 , \5159 , \5169 );
or \U$5270 ( \5402 , \5399 , \5400 , \5401 );
and \U$5271 ( \5403 , \5174 , \5178 );
and \U$5272 ( \5404 , \5178 , \5183 );
and \U$5273 ( \5405 , \5174 , \5183 );
or \U$5274 ( \5406 , \5403 , \5404 , \5405 );
xor \U$5275 ( \5407 , \5402 , \5406 );
and \U$5276 ( \5408 , \5189 , \5193 );
and \U$5277 ( \5409 , \5193 , \5198 );
and \U$5278 ( \5410 , \5189 , \5198 );
or \U$5279 ( \5411 , \5408 , \5409 , \5410 );
xor \U$5280 ( \5412 , \5407 , \5411 );
and \U$5281 ( \5413 , \5220 , \5224 );
and \U$5282 ( \5414 , \5224 , \5229 );
and \U$5283 ( \5415 , \5220 , \5229 );
or \U$5284 ( \5416 , \5413 , \5414 , \5415 );
and \U$5285 ( \5417 , \5234 , \5238 );
and \U$5286 ( \5418 , \5238 , \5243 );
and \U$5287 ( \5419 , \5234 , \5243 );
or \U$5288 ( \5420 , \5417 , \5418 , \5419 );
xor \U$5289 ( \5421 , \5416 , \5420 );
and \U$5290 ( \5422 , \5249 , \5253 );
and \U$5291 ( \5423 , \5253 , \5258 );
and \U$5292 ( \5424 , \5249 , \5258 );
or \U$5293 ( \5425 , \5422 , \5423 , \5424 );
xor \U$5294 ( \5426 , \5421 , \5425 );
xor \U$5295 ( \5427 , \5412 , \5426 );
and \U$5296 ( \5428 , \5269 , \5273 );
and \U$5297 ( \5429 , \5273 , \5277 );
and \U$5298 ( \5430 , \5269 , \5277 );
or \U$5299 ( \5431 , \5428 , \5429 , \5430 );
and \U$5300 ( \5432 , \5283 , \5287 );
and \U$5301 ( \5433 , \5287 , \5292 );
and \U$5302 ( \5434 , \5283 , \5292 );
or \U$5303 ( \5435 , \5432 , \5433 , \5434 );
xor \U$5304 ( \5436 , \5431 , \5435 );
and \U$5305 ( \5437 , \158 , \5011 );
and \U$5306 ( \5438 , \134 , \4878 );
nor \U$5307 ( \5439 , \5437 , \5438 );
xnor \U$5308 ( \5440 , \5439 , \4762 );
xor \U$5309 ( \5441 , \5436 , \5440 );
xor \U$5310 ( \5442 , \5427 , \5441 );
and \U$5311 ( \5443 , \5230 , \5244 );
and \U$5312 ( \5444 , \5244 , \5259 );
and \U$5313 ( \5445 , \5230 , \5259 );
or \U$5314 ( \5446 , \5443 , \5444 , \5445 );
and \U$5315 ( \5447 , \5170 , \5184 );
and \U$5316 ( \5448 , \5184 , \5199 );
and \U$5317 ( \5449 , \5170 , \5199 );
or \U$5318 ( \5450 , \5447 , \5448 , \5449 );
xor \U$5319 ( \5451 , \5446 , \5450 );
and \U$5320 ( \5452 , \3912 , \230 );
and \U$5321 ( \5453 , \4160 , \228 );
nor \U$5322 ( \5454 , \5452 , \5453 );
xnor \U$5323 ( \5455 , \5454 , \237 );
and \U$5324 ( \5456 , \3646 , \245 );
and \U$5325 ( \5457 , \3736 , \243 );
nor \U$5326 ( \5458 , \5456 , \5457 );
xnor \U$5327 ( \5459 , \5458 , \252 );
xor \U$5328 ( \5460 , \5455 , \5459 );
and \U$5329 ( \5461 , \3143 , \141 );
and \U$5330 ( \5462 , \3395 , \139 );
nor \U$5331 ( \5463 , \5461 , \5462 );
xnor \U$5332 ( \5464 , \5463 , \148 );
xor \U$5333 ( \5465 , \5460 , \5464 );
xor \U$5334 ( \5466 , \5451 , \5465 );
xor \U$5335 ( \5467 , \5442 , \5466 );
and \U$5336 ( \5468 , \5156 , \183 );
buf \U$5337 ( \5469 , RIb55e950_83);
and \U$5338 ( \5470 , \5469 , \180 );
nor \U$5339 ( \5471 , \5468 , \5470 );
xnor \U$5340 ( \5472 , \5471 , \179 );
and \U$5341 ( \5473 , \4749 , \195 );
and \U$5342 ( \5474 , \4922 , \193 );
nor \U$5343 ( \5475 , \5473 , \5474 );
xnor \U$5344 ( \5476 , \5475 , \202 );
xor \U$5345 ( \5477 , \5472 , \5476 );
and \U$5346 ( \5478 , \4364 , \215 );
and \U$5347 ( \5479 , \4654 , \213 );
nor \U$5348 ( \5480 , \5478 , \5479 );
xnor \U$5349 ( \5481 , \5480 , \222 );
xor \U$5350 ( \5482 , \5477 , \5481 );
xor \U$5351 ( \5483 , \5165 , \5166 );
not \U$5352 ( \5484 , \5275 );
and \U$5353 ( \5485 , \5483 , \5484 );
and \U$5354 ( \5486 , \166 , \5485 );
and \U$5355 ( \5487 , \150 , \5275 );
nor \U$5356 ( \5488 , \5486 , \5487 );
xnor \U$5357 ( \5489 , \5488 , \5169 );
and \U$5358 ( \5490 , \185 , \2669 );
and \U$5359 ( \5491 , \261 , \2538 );
nor \U$5360 ( \5492 , \5490 , \5491 );
xnor \U$5361 ( \5493 , \5492 , \2534 );
and \U$5362 ( \5494 , \197 , \3103 );
and \U$5363 ( \5495 , \178 , \2934 );
nor \U$5364 ( \5496 , \5494 , \5495 );
xnor \U$5365 ( \5497 , \5496 , \2839 );
xor \U$5366 ( \5498 , \5493 , \5497 );
and \U$5367 ( \5499 , \217 , \3357 );
and \U$5368 ( \5500 , \189 , \3255 );
nor \U$5369 ( \5501 , \5499 , \5500 );
xnor \U$5370 ( \5502 , \5501 , \3156 );
xor \U$5371 ( \5503 , \5498 , \5502 );
xor \U$5372 ( \5504 , \5489 , \5503 );
and \U$5373 ( \5505 , \232 , \3813 );
and \U$5374 ( \5506 , \209 , \3557 );
nor \U$5375 ( \5507 , \5505 , \5506 );
xnor \U$5376 ( \5508 , \5507 , \3562 );
and \U$5377 ( \5509 , \247 , \4132 );
and \U$5378 ( \5510 , \224 , \4012 );
nor \U$5379 ( \5511 , \5509 , \5510 );
xnor \U$5380 ( \5512 , \5511 , \3925 );
xor \U$5381 ( \5513 , \5508 , \5512 );
and \U$5382 ( \5514 , \143 , \4581 );
and \U$5383 ( \5515 , \240 , \4424 );
nor \U$5384 ( \5516 , \5514 , \5515 );
xnor \U$5385 ( \5517 , \5516 , \4377 );
xor \U$5386 ( \5518 , \5513 , \5517 );
xor \U$5387 ( \5519 , \5504 , \5518 );
xor \U$5388 ( \5520 , \5482 , \5519 );
and \U$5389 ( \5521 , \1948 , \1086 );
and \U$5390 ( \5522 , \2090 , \508 );
nor \U$5391 ( \5523 , \5521 , \5522 );
xnor \U$5392 ( \5524 , \5523 , \487 );
and \U$5393 ( \5525 , \1684 , \1301 );
and \U$5394 ( \5526 , \1802 , \1246 );
nor \U$5395 ( \5527 , \5525 , \5526 );
xnor \U$5396 ( \5528 , \5527 , \1205 );
xor \U$5397 ( \5529 , \5524 , \5528 );
and \U$5398 ( \5530 , \1484 , \1578 );
and \U$5399 ( \5531 , \1601 , \1431 );
nor \U$5400 ( \5532 , \5530 , \5531 );
xnor \U$5401 ( \5533 , \5532 , \1436 );
xor \U$5402 ( \5534 , \5529 , \5533 );
and \U$5403 ( \5535 , \1192 , \1824 );
and \U$5404 ( \5536 , \1333 , \1739 );
nor \U$5405 ( \5537 , \5535 , \5536 );
xnor \U$5406 ( \5538 , \5537 , \1697 );
and \U$5407 ( \5539 , \474 , \2121 );
and \U$5408 ( \5540 , \1147 , \2008 );
nor \U$5409 ( \5541 , \5539 , \5540 );
xnor \U$5410 ( \5542 , \5541 , \1961 );
xor \U$5411 ( \5543 , \5538 , \5542 );
and \U$5412 ( \5544 , \307 , \2400 );
and \U$5413 ( \5545 , \412 , \2246 );
nor \U$5414 ( \5546 , \5544 , \5545 );
xnor \U$5415 ( \5547 , \5546 , \2195 );
xor \U$5416 ( \5548 , \5543 , \5547 );
xor \U$5417 ( \5549 , \5534 , \5548 );
and \U$5418 ( \5550 , \2826 , \156 );
and \U$5419 ( \5551 , \3037 , \154 );
nor \U$5420 ( \5552 , \5550 , \5551 );
xnor \U$5421 ( \5553 , \5552 , \163 );
and \U$5422 ( \5554 , \2521 , \296 );
and \U$5423 ( \5555 , \2757 , \168 );
nor \U$5424 ( \5556 , \5554 , \5555 );
xnor \U$5425 ( \5557 , \5556 , \173 );
xor \U$5426 ( \5558 , \5553 , \5557 );
and \U$5427 ( \5559 , \2182 , \438 );
and \U$5428 ( \5560 , \2366 , \336 );
nor \U$5429 ( \5561 , \5559 , \5560 );
xnor \U$5430 ( \5562 , \5561 , \320 );
xor \U$5431 ( \5563 , \5558 , \5562 );
xor \U$5432 ( \5564 , \5549 , \5563 );
xor \U$5433 ( \5565 , \5520 , \5564 );
xor \U$5434 ( \5566 , \5467 , \5565 );
xor \U$5435 ( \5567 , \5398 , \5566 );
xor \U$5436 ( \5568 , \5384 , \5567 );
xor \U$5437 ( \5569 , \5355 , \5568 );
and \U$5438 ( \5570 , \5122 , \5297 );
and \U$5439 ( \5571 , \5297 , \5337 );
and \U$5440 ( \5572 , \5122 , \5337 );
or \U$5441 ( \5573 , \5570 , \5571 , \5572 );
xor \U$5442 ( \5574 , \5569 , \5573 );
and \U$5443 ( \5575 , \5338 , \5342 );
and \U$5444 ( \5576 , \5343 , \5346 );
or \U$5445 ( \5577 , \5575 , \5576 );
xor \U$5446 ( \5578 , \5574 , \5577 );
buf \U$5447 ( \5579 , \5578 );
buf \U$5448 ( \5580 , \5579 );
and \U$5449 ( \5581 , \5359 , \5383 );
and \U$5450 ( \5582 , \5383 , \5567 );
and \U$5451 ( \5583 , \5359 , \5567 );
or \U$5452 ( \5584 , \5581 , \5582 , \5583 );
and \U$5453 ( \5585 , \5363 , \5367 );
and \U$5454 ( \5586 , \5367 , \5382 );
and \U$5455 ( \5587 , \5363 , \5382 );
or \U$5456 ( \5588 , \5585 , \5586 , \5587 );
and \U$5457 ( \5589 , \5398 , \5566 );
xor \U$5458 ( \5590 , \5588 , \5589 );
and \U$5459 ( \5591 , \5412 , \5426 );
and \U$5460 ( \5592 , \5426 , \5441 );
and \U$5461 ( \5593 , \5412 , \5441 );
or \U$5462 ( \5594 , \5591 , \5592 , \5593 );
and \U$5463 ( \5595 , \5524 , \5528 );
and \U$5464 ( \5596 , \5528 , \5533 );
and \U$5465 ( \5597 , \5524 , \5533 );
or \U$5466 ( \5598 , \5595 , \5596 , \5597 );
and \U$5467 ( \5599 , \5538 , \5542 );
and \U$5468 ( \5600 , \5542 , \5547 );
and \U$5469 ( \5601 , \5538 , \5547 );
or \U$5470 ( \5602 , \5599 , \5600 , \5601 );
xor \U$5471 ( \5603 , \5598 , \5602 );
and \U$5472 ( \5604 , \5493 , \5497 );
and \U$5473 ( \5605 , \5497 , \5502 );
and \U$5474 ( \5606 , \5493 , \5502 );
or \U$5475 ( \5607 , \5604 , \5605 , \5606 );
xor \U$5476 ( \5608 , \5603 , \5607 );
xor \U$5477 ( \5609 , \5594 , \5608 );
and \U$5478 ( \5610 , \5455 , \5459 );
and \U$5479 ( \5611 , \5459 , \5464 );
and \U$5480 ( \5612 , \5455 , \5464 );
or \U$5481 ( \5613 , \5610 , \5611 , \5612 );
and \U$5482 ( \5614 , \5553 , \5557 );
and \U$5483 ( \5615 , \5557 , \5562 );
and \U$5484 ( \5616 , \5553 , \5562 );
or \U$5485 ( \5617 , \5614 , \5615 , \5616 );
xor \U$5486 ( \5618 , \5613 , \5617 );
and \U$5487 ( \5619 , \5472 , \5476 );
and \U$5488 ( \5620 , \5476 , \5481 );
and \U$5489 ( \5621 , \5472 , \5481 );
or \U$5490 ( \5622 , \5619 , \5620 , \5621 );
xor \U$5491 ( \5623 , \5618 , \5622 );
xor \U$5492 ( \5624 , \5609 , \5623 );
xor \U$5493 ( \5625 , \5590 , \5624 );
xor \U$5494 ( \5626 , \5584 , \5625 );
and \U$5495 ( \5627 , \5372 , \5376 );
and \U$5496 ( \5628 , \5376 , \5381 );
and \U$5497 ( \5629 , \5372 , \5381 );
or \U$5498 ( \5630 , \5627 , \5628 , \5629 );
and \U$5499 ( \5631 , \5446 , \5450 );
and \U$5500 ( \5632 , \5450 , \5465 );
and \U$5501 ( \5633 , \5446 , \5465 );
or \U$5502 ( \5634 , \5631 , \5632 , \5633 );
xor \U$5503 ( \5635 , \5630 , \5634 );
and \U$5504 ( \5636 , \5482 , \5519 );
and \U$5505 ( \5637 , \5519 , \5564 );
and \U$5506 ( \5638 , \5482 , \5564 );
or \U$5507 ( \5639 , \5636 , \5637 , \5638 );
xor \U$5508 ( \5640 , \5635 , \5639 );
and \U$5509 ( \5641 , \5388 , \5392 );
and \U$5510 ( \5642 , \5392 , \5397 );
and \U$5511 ( \5643 , \5388 , \5397 );
or \U$5512 ( \5644 , \5641 , \5642 , \5643 );
and \U$5513 ( \5645 , \5442 , \5466 );
and \U$5514 ( \5646 , \5466 , \5565 );
and \U$5515 ( \5647 , \5442 , \5565 );
or \U$5516 ( \5648 , \5645 , \5646 , \5647 );
xor \U$5517 ( \5649 , \5644 , \5648 );
and \U$5518 ( \5650 , \5402 , \5406 );
and \U$5519 ( \5651 , \5406 , \5411 );
and \U$5520 ( \5652 , \5402 , \5411 );
or \U$5521 ( \5653 , \5650 , \5651 , \5652 );
and \U$5522 ( \5654 , \5416 , \5420 );
and \U$5523 ( \5655 , \5420 , \5425 );
and \U$5524 ( \5656 , \5416 , \5425 );
or \U$5525 ( \5657 , \5654 , \5655 , \5656 );
xor \U$5526 ( \5658 , \5653 , \5657 );
and \U$5527 ( \5659 , \5431 , \5435 );
and \U$5528 ( \5660 , \5435 , \5440 );
and \U$5529 ( \5661 , \5431 , \5440 );
or \U$5530 ( \5662 , \5659 , \5660 , \5661 );
xor \U$5531 ( \5663 , \5658 , \5662 );
and \U$5532 ( \5664 , \5489 , \5503 );
and \U$5533 ( \5665 , \5503 , \5518 );
and \U$5534 ( \5666 , \5489 , \5518 );
or \U$5535 ( \5667 , \5664 , \5665 , \5666 );
and \U$5536 ( \5668 , \5534 , \5548 );
and \U$5537 ( \5669 , \5548 , \5563 );
and \U$5538 ( \5670 , \5534 , \5563 );
or \U$5539 ( \5671 , \5668 , \5669 , \5670 );
xor \U$5540 ( \5672 , \5667 , \5671 );
and \U$5541 ( \5673 , \5469 , \183 );
buf \U$5542 ( \5674 , RIb55e9c8_82);
and \U$5543 ( \5675 , \5674 , \180 );
nor \U$5544 ( \5676 , \5673 , \5675 );
xnor \U$5545 ( \5677 , \5676 , \179 );
and \U$5546 ( \5678 , \4922 , \195 );
and \U$5547 ( \5679 , \5156 , \193 );
nor \U$5548 ( \5680 , \5678 , \5679 );
xnor \U$5549 ( \5681 , \5680 , \202 );
xor \U$5550 ( \5682 , \5677 , \5681 );
buf \U$5551 ( \5683 , RIb560840_17);
buf \U$5552 ( \5684 , RIb5607c8_18);
and \U$5553 ( \5685 , \5684 , \5165 );
not \U$5554 ( \5686 , \5685 );
and \U$5555 ( \5687 , \5683 , \5686 );
xor \U$5556 ( \5688 , \5682 , \5687 );
xor \U$5557 ( \5689 , \5672 , \5688 );
xor \U$5558 ( \5690 , \5663 , \5689 );
and \U$5559 ( \5691 , \5508 , \5512 );
and \U$5560 ( \5692 , \5512 , \5517 );
and \U$5561 ( \5693 , \5508 , \5517 );
or \U$5562 ( \5694 , \5691 , \5692 , \5693 );
xor \U$5563 ( \5695 , \5684 , \5165 );
nand \U$5564 ( \5696 , \166 , \5695 );
xnor \U$5565 ( \5697 , \5696 , \5687 );
xor \U$5566 ( \5698 , \5694 , \5697 );
and \U$5567 ( \5699 , \240 , \4581 );
and \U$5568 ( \5700 , \247 , \4424 );
nor \U$5569 ( \5701 , \5699 , \5700 );
xnor \U$5570 ( \5702 , \5701 , \4377 );
and \U$5571 ( \5703 , \134 , \5011 );
and \U$5572 ( \5704 , \143 , \4878 );
nor \U$5573 ( \5705 , \5703 , \5704 );
xnor \U$5574 ( \5706 , \5705 , \4762 );
xor \U$5575 ( \5707 , \5702 , \5706 );
and \U$5576 ( \5708 , \150 , \5485 );
and \U$5577 ( \5709 , \158 , \5275 );
nor \U$5578 ( \5710 , \5708 , \5709 );
xnor \U$5579 ( \5711 , \5710 , \5169 );
xor \U$5580 ( \5712 , \5707 , \5711 );
xor \U$5581 ( \5713 , \5698 , \5712 );
and \U$5582 ( \5714 , \412 , \2400 );
and \U$5583 ( \5715 , \474 , \2246 );
nor \U$5584 ( \5716 , \5714 , \5715 );
xnor \U$5585 ( \5717 , \5716 , \2195 );
and \U$5586 ( \5718 , \261 , \2669 );
and \U$5587 ( \5719 , \307 , \2538 );
nor \U$5588 ( \5720 , \5718 , \5719 );
xnor \U$5589 ( \5721 , \5720 , \2534 );
xor \U$5590 ( \5722 , \5717 , \5721 );
and \U$5591 ( \5723 , \178 , \3103 );
and \U$5592 ( \5724 , \185 , \2934 );
nor \U$5593 ( \5725 , \5723 , \5724 );
xnor \U$5594 ( \5726 , \5725 , \2839 );
xor \U$5595 ( \5727 , \5722 , \5726 );
and \U$5596 ( \5728 , \189 , \3357 );
and \U$5597 ( \5729 , \197 , \3255 );
nor \U$5598 ( \5730 , \5728 , \5729 );
xnor \U$5599 ( \5731 , \5730 , \3156 );
and \U$5600 ( \5732 , \209 , \3813 );
and \U$5601 ( \5733 , \217 , \3557 );
nor \U$5602 ( \5734 , \5732 , \5733 );
xnor \U$5603 ( \5735 , \5734 , \3562 );
xor \U$5604 ( \5736 , \5731 , \5735 );
and \U$5605 ( \5737 , \224 , \4132 );
and \U$5606 ( \5738 , \232 , \4012 );
nor \U$5607 ( \5739 , \5737 , \5738 );
xnor \U$5608 ( \5740 , \5739 , \3925 );
xor \U$5609 ( \5741 , \5736 , \5740 );
xor \U$5610 ( \5742 , \5727 , \5741 );
and \U$5611 ( \5743 , \1601 , \1578 );
and \U$5612 ( \5744 , \1684 , \1431 );
nor \U$5613 ( \5745 , \5743 , \5744 );
xnor \U$5614 ( \5746 , \5745 , \1436 );
and \U$5615 ( \5747 , \1333 , \1824 );
and \U$5616 ( \5748 , \1484 , \1739 );
nor \U$5617 ( \5749 , \5747 , \5748 );
xnor \U$5618 ( \5750 , \5749 , \1697 );
xor \U$5619 ( \5751 , \5746 , \5750 );
and \U$5620 ( \5752 , \1147 , \2121 );
and \U$5621 ( \5753 , \1192 , \2008 );
nor \U$5622 ( \5754 , \5752 , \5753 );
xnor \U$5623 ( \5755 , \5754 , \1961 );
xor \U$5624 ( \5756 , \5751 , \5755 );
xor \U$5625 ( \5757 , \5742 , \5756 );
xor \U$5626 ( \5758 , \5713 , \5757 );
and \U$5627 ( \5759 , \4654 , \215 );
and \U$5628 ( \5760 , \4749 , \213 );
nor \U$5629 ( \5761 , \5759 , \5760 );
xnor \U$5630 ( \5762 , \5761 , \222 );
and \U$5631 ( \5763 , \4160 , \230 );
and \U$5632 ( \5764 , \4364 , \228 );
nor \U$5633 ( \5765 , \5763 , \5764 );
xnor \U$5634 ( \5766 , \5765 , \237 );
xor \U$5635 ( \5767 , \5762 , \5766 );
and \U$5636 ( \5768 , \3736 , \245 );
and \U$5637 ( \5769 , \3912 , \243 );
nor \U$5638 ( \5770 , \5768 , \5769 );
xnor \U$5639 ( \5771 , \5770 , \252 );
xor \U$5640 ( \5772 , \5767 , \5771 );
and \U$5641 ( \5773 , \2366 , \438 );
and \U$5642 ( \5774 , \2521 , \336 );
nor \U$5643 ( \5775 , \5773 , \5774 );
xnor \U$5644 ( \5776 , \5775 , \320 );
and \U$5645 ( \5777 , \2090 , \1086 );
and \U$5646 ( \5778 , \2182 , \508 );
nor \U$5647 ( \5779 , \5777 , \5778 );
xnor \U$5648 ( \5780 , \5779 , \487 );
xor \U$5649 ( \5781 , \5776 , \5780 );
and \U$5650 ( \5782 , \1802 , \1301 );
and \U$5651 ( \5783 , \1948 , \1246 );
nor \U$5652 ( \5784 , \5782 , \5783 );
xnor \U$5653 ( \5785 , \5784 , \1205 );
xor \U$5654 ( \5786 , \5781 , \5785 );
xor \U$5655 ( \5787 , \5772 , \5786 );
and \U$5656 ( \5788 , \3395 , \141 );
and \U$5657 ( \5789 , \3646 , \139 );
nor \U$5658 ( \5790 , \5788 , \5789 );
xnor \U$5659 ( \5791 , \5790 , \148 );
and \U$5660 ( \5792 , \3037 , \156 );
and \U$5661 ( \5793 , \3143 , \154 );
nor \U$5662 ( \5794 , \5792 , \5793 );
xnor \U$5663 ( \5795 , \5794 , \163 );
xor \U$5664 ( \5796 , \5791 , \5795 );
and \U$5665 ( \5797 , \2757 , \296 );
and \U$5666 ( \5798 , \2826 , \168 );
nor \U$5667 ( \5799 , \5797 , \5798 );
xnor \U$5668 ( \5800 , \5799 , \173 );
xor \U$5669 ( \5801 , \5796 , \5800 );
xor \U$5670 ( \5802 , \5787 , \5801 );
xor \U$5671 ( \5803 , \5758 , \5802 );
xor \U$5672 ( \5804 , \5690 , \5803 );
xor \U$5673 ( \5805 , \5649 , \5804 );
xor \U$5674 ( \5806 , \5640 , \5805 );
xor \U$5675 ( \5807 , \5626 , \5806 );
and \U$5676 ( \5808 , \5353 , \5354 );
and \U$5677 ( \5809 , \5354 , \5568 );
and \U$5678 ( \5810 , \5353 , \5568 );
or \U$5679 ( \5811 , \5808 , \5809 , \5810 );
xor \U$5680 ( \5812 , \5807 , \5811 );
and \U$5681 ( \5813 , \5569 , \5573 );
and \U$5682 ( \5814 , \5574 , \5577 );
or \U$5683 ( \5815 , \5813 , \5814 );
xor \U$5684 ( \5816 , \5812 , \5815 );
buf \U$5685 ( \5817 , \5816 );
buf \U$5686 ( \5818 , \5817 );
and \U$5687 ( \5819 , \5588 , \5589 );
and \U$5688 ( \5820 , \5589 , \5624 );
and \U$5689 ( \5821 , \5588 , \5624 );
or \U$5690 ( \5822 , \5819 , \5820 , \5821 );
and \U$5691 ( \5823 , \5640 , \5805 );
xor \U$5692 ( \5824 , \5822 , \5823 );
and \U$5693 ( \5825 , \5644 , \5648 );
and \U$5694 ( \5826 , \5648 , \5804 );
and \U$5695 ( \5827 , \5644 , \5804 );
or \U$5696 ( \5828 , \5825 , \5826 , \5827 );
and \U$5697 ( \5829 , \5630 , \5634 );
and \U$5698 ( \5830 , \5634 , \5639 );
and \U$5699 ( \5831 , \5630 , \5639 );
or \U$5700 ( \5832 , \5829 , \5830 , \5831 );
and \U$5701 ( \5833 , \5594 , \5608 );
and \U$5702 ( \5834 , \5608 , \5623 );
and \U$5703 ( \5835 , \5594 , \5623 );
or \U$5704 ( \5836 , \5833 , \5834 , \5835 );
xor \U$5705 ( \5837 , \5832 , \5836 );
and \U$5706 ( \5838 , \5663 , \5689 );
and \U$5707 ( \5839 , \5689 , \5803 );
and \U$5708 ( \5840 , \5663 , \5803 );
or \U$5709 ( \5841 , \5838 , \5839 , \5840 );
xor \U$5710 ( \5842 , \5837 , \5841 );
xor \U$5711 ( \5843 , \5828 , \5842 );
and \U$5712 ( \5844 , \5653 , \5657 );
and \U$5713 ( \5845 , \5657 , \5662 );
and \U$5714 ( \5846 , \5653 , \5662 );
or \U$5715 ( \5847 , \5844 , \5845 , \5846 );
and \U$5716 ( \5848 , \5667 , \5671 );
and \U$5717 ( \5849 , \5671 , \5688 );
and \U$5718 ( \5850 , \5667 , \5688 );
or \U$5719 ( \5851 , \5848 , \5849 , \5850 );
xor \U$5720 ( \5852 , \5847 , \5851 );
and \U$5721 ( \5853 , \5713 , \5757 );
and \U$5722 ( \5854 , \5757 , \5802 );
and \U$5723 ( \5855 , \5713 , \5802 );
or \U$5724 ( \5856 , \5853 , \5854 , \5855 );
xor \U$5725 ( \5857 , \5852 , \5856 );
and \U$5726 ( \5858 , \5717 , \5721 );
and \U$5727 ( \5859 , \5721 , \5726 );
and \U$5728 ( \5860 , \5717 , \5726 );
or \U$5729 ( \5861 , \5858 , \5859 , \5860 );
and \U$5730 ( \5862 , \5746 , \5750 );
and \U$5731 ( \5863 , \5750 , \5755 );
and \U$5732 ( \5864 , \5746 , \5755 );
or \U$5733 ( \5865 , \5862 , \5863 , \5864 );
xor \U$5734 ( \5866 , \5861 , \5865 );
and \U$5735 ( \5867 , \5776 , \5780 );
and \U$5736 ( \5868 , \5780 , \5785 );
and \U$5737 ( \5869 , \5776 , \5785 );
or \U$5738 ( \5870 , \5867 , \5868 , \5869 );
xor \U$5739 ( \5871 , \5866 , \5870 );
and \U$5740 ( \5872 , \5762 , \5766 );
and \U$5741 ( \5873 , \5766 , \5771 );
and \U$5742 ( \5874 , \5762 , \5771 );
or \U$5743 ( \5875 , \5872 , \5873 , \5874 );
and \U$5744 ( \5876 , \5677 , \5681 );
and \U$5745 ( \5877 , \5681 , \5687 );
and \U$5746 ( \5878 , \5677 , \5687 );
or \U$5747 ( \5879 , \5876 , \5877 , \5878 );
xor \U$5748 ( \5880 , \5875 , \5879 );
and \U$5749 ( \5881 , \5791 , \5795 );
and \U$5750 ( \5882 , \5795 , \5800 );
and \U$5751 ( \5883 , \5791 , \5800 );
or \U$5752 ( \5884 , \5881 , \5882 , \5883 );
xor \U$5753 ( \5885 , \5880 , \5884 );
xor \U$5754 ( \5886 , \5871 , \5885 );
and \U$5755 ( \5887 , \217 , \3813 );
and \U$5756 ( \5888 , \189 , \3557 );
nor \U$5757 ( \5889 , \5887 , \5888 );
xnor \U$5758 ( \5890 , \5889 , \3562 );
and \U$5759 ( \5891 , \232 , \4132 );
and \U$5760 ( \5892 , \209 , \4012 );
nor \U$5761 ( \5893 , \5891 , \5892 );
xnor \U$5762 ( \5894 , \5893 , \3925 );
xor \U$5763 ( \5895 , \5890 , \5894 );
and \U$5764 ( \5896 , \247 , \4581 );
and \U$5765 ( \5897 , \224 , \4424 );
nor \U$5766 ( \5898 , \5896 , \5897 );
xnor \U$5767 ( \5899 , \5898 , \4377 );
xor \U$5768 ( \5900 , \5895 , \5899 );
and \U$5769 ( \5901 , \1484 , \1824 );
and \U$5770 ( \5902 , \1601 , \1739 );
nor \U$5771 ( \5903 , \5901 , \5902 );
xnor \U$5772 ( \5904 , \5903 , \1697 );
and \U$5773 ( \5905 , \1192 , \2121 );
and \U$5774 ( \5906 , \1333 , \2008 );
nor \U$5775 ( \5907 , \5905 , \5906 );
xnor \U$5776 ( \5908 , \5907 , \1961 );
xor \U$5777 ( \5909 , \5904 , \5908 );
and \U$5778 ( \5910 , \474 , \2400 );
and \U$5779 ( \5911 , \1147 , \2246 );
nor \U$5780 ( \5912 , \5910 , \5911 );
xnor \U$5781 ( \5913 , \5912 , \2195 );
xor \U$5782 ( \5914 , \5909 , \5913 );
xor \U$5783 ( \5915 , \5900 , \5914 );
and \U$5784 ( \5916 , \307 , \2669 );
and \U$5785 ( \5917 , \412 , \2538 );
nor \U$5786 ( \5918 , \5916 , \5917 );
xnor \U$5787 ( \5919 , \5918 , \2534 );
and \U$5788 ( \5920 , \185 , \3103 );
and \U$5789 ( \5921 , \261 , \2934 );
nor \U$5790 ( \5922 , \5920 , \5921 );
xnor \U$5791 ( \5923 , \5922 , \2839 );
xor \U$5792 ( \5924 , \5919 , \5923 );
and \U$5793 ( \5925 , \197 , \3357 );
and \U$5794 ( \5926 , \178 , \3255 );
nor \U$5795 ( \5927 , \5925 , \5926 );
xnor \U$5796 ( \5928 , \5927 , \3156 );
xor \U$5797 ( \5929 , \5924 , \5928 );
xor \U$5798 ( \5930 , \5915 , \5929 );
and \U$5799 ( \5931 , \4364 , \230 );
and \U$5800 ( \5932 , \4654 , \228 );
nor \U$5801 ( \5933 , \5931 , \5932 );
xnor \U$5802 ( \5934 , \5933 , \237 );
and \U$5803 ( \5935 , \3912 , \245 );
and \U$5804 ( \5936 , \4160 , \243 );
nor \U$5805 ( \5937 , \5935 , \5936 );
xnor \U$5806 ( \5938 , \5937 , \252 );
xor \U$5807 ( \5939 , \5934 , \5938 );
and \U$5808 ( \5940 , \3646 , \141 );
and \U$5809 ( \5941 , \3736 , \139 );
nor \U$5810 ( \5942 , \5940 , \5941 );
xnor \U$5811 ( \5943 , \5942 , \148 );
xor \U$5812 ( \5944 , \5939 , \5943 );
and \U$5813 ( \5945 , \2182 , \1086 );
and \U$5814 ( \5946 , \2366 , \508 );
nor \U$5815 ( \5947 , \5945 , \5946 );
xnor \U$5816 ( \5948 , \5947 , \487 );
and \U$5817 ( \5949 , \1948 , \1301 );
and \U$5818 ( \5950 , \2090 , \1246 );
nor \U$5819 ( \5951 , \5949 , \5950 );
xnor \U$5820 ( \5952 , \5951 , \1205 );
xor \U$5821 ( \5953 , \5948 , \5952 );
and \U$5822 ( \5954 , \1684 , \1578 );
and \U$5823 ( \5955 , \1802 , \1431 );
nor \U$5824 ( \5956 , \5954 , \5955 );
xnor \U$5825 ( \5957 , \5956 , \1436 );
xor \U$5826 ( \5958 , \5953 , \5957 );
xor \U$5827 ( \5959 , \5944 , \5958 );
and \U$5828 ( \5960 , \3143 , \156 );
and \U$5829 ( \5961 , \3395 , \154 );
nor \U$5830 ( \5962 , \5960 , \5961 );
xnor \U$5831 ( \5963 , \5962 , \163 );
and \U$5832 ( \5964 , \2826 , \296 );
and \U$5833 ( \5965 , \3037 , \168 );
nor \U$5834 ( \5966 , \5964 , \5965 );
xnor \U$5835 ( \5967 , \5966 , \173 );
xor \U$5836 ( \5968 , \5963 , \5967 );
and \U$5837 ( \5969 , \2521 , \438 );
and \U$5838 ( \5970 , \2757 , \336 );
nor \U$5839 ( \5971 , \5969 , \5970 );
xnor \U$5840 ( \5972 , \5971 , \320 );
xor \U$5841 ( \5973 , \5968 , \5972 );
xor \U$5842 ( \5974 , \5959 , \5973 );
xor \U$5843 ( \5975 , \5930 , \5974 );
and \U$5844 ( \5976 , \5731 , \5735 );
and \U$5845 ( \5977 , \5735 , \5740 );
and \U$5846 ( \5978 , \5731 , \5740 );
or \U$5847 ( \5979 , \5976 , \5977 , \5978 );
and \U$5848 ( \5980 , \5702 , \5706 );
and \U$5849 ( \5981 , \5706 , \5711 );
and \U$5850 ( \5982 , \5702 , \5711 );
or \U$5851 ( \5983 , \5980 , \5981 , \5982 );
xor \U$5852 ( \5984 , \5979 , \5983 );
and \U$5853 ( \5985 , \143 , \5011 );
and \U$5854 ( \5986 , \240 , \4878 );
nor \U$5855 ( \5987 , \5985 , \5986 );
xnor \U$5856 ( \5988 , \5987 , \4762 );
and \U$5857 ( \5989 , \158 , \5485 );
and \U$5858 ( \5990 , \134 , \5275 );
nor \U$5859 ( \5991 , \5989 , \5990 );
xnor \U$5860 ( \5992 , \5991 , \5169 );
xor \U$5861 ( \5993 , \5988 , \5992 );
xor \U$5862 ( \5994 , \5683 , \5684 );
not \U$5863 ( \5995 , \5695 );
and \U$5864 ( \5996 , \5994 , \5995 );
and \U$5865 ( \5997 , \166 , \5996 );
and \U$5866 ( \5998 , \150 , \5695 );
nor \U$5867 ( \5999 , \5997 , \5998 );
xnor \U$5868 ( \6000 , \5999 , \5687 );
xor \U$5869 ( \6001 , \5993 , \6000 );
xor \U$5870 ( \6002 , \5984 , \6001 );
xor \U$5871 ( \6003 , \5975 , \6002 );
xor \U$5872 ( \6004 , \5886 , \6003 );
xor \U$5873 ( \6005 , \5857 , \6004 );
and \U$5874 ( \6006 , \5598 , \5602 );
and \U$5875 ( \6007 , \5602 , \5607 );
and \U$5876 ( \6008 , \5598 , \5607 );
or \U$5877 ( \6009 , \6006 , \6007 , \6008 );
and \U$5878 ( \6010 , \5613 , \5617 );
and \U$5879 ( \6011 , \5617 , \5622 );
and \U$5880 ( \6012 , \5613 , \5622 );
or \U$5881 ( \6013 , \6010 , \6011 , \6012 );
xor \U$5882 ( \6014 , \6009 , \6013 );
and \U$5883 ( \6015 , \5694 , \5697 );
and \U$5884 ( \6016 , \5697 , \5712 );
and \U$5885 ( \6017 , \5694 , \5712 );
or \U$5886 ( \6018 , \6015 , \6016 , \6017 );
xor \U$5887 ( \6019 , \6014 , \6018 );
and \U$5888 ( \6020 , \5727 , \5741 );
and \U$5889 ( \6021 , \5741 , \5756 );
and \U$5890 ( \6022 , \5727 , \5756 );
or \U$5891 ( \6023 , \6020 , \6021 , \6022 );
and \U$5892 ( \6024 , \5772 , \5786 );
and \U$5893 ( \6025 , \5786 , \5801 );
and \U$5894 ( \6026 , \5772 , \5801 );
or \U$5895 ( \6027 , \6024 , \6025 , \6026 );
xor \U$5896 ( \6028 , \6023 , \6027 );
and \U$5897 ( \6029 , \5674 , \183 );
buf \U$5898 ( \6030 , RIb55ea40_81);
and \U$5899 ( \6031 , \6030 , \180 );
nor \U$5900 ( \6032 , \6029 , \6031 );
xnor \U$5901 ( \6033 , \6032 , \179 );
and \U$5902 ( \6034 , \5156 , \195 );
and \U$5903 ( \6035 , \5469 , \193 );
nor \U$5904 ( \6036 , \6034 , \6035 );
xnor \U$5905 ( \6037 , \6036 , \202 );
xor \U$5906 ( \6038 , \6033 , \6037 );
and \U$5907 ( \6039 , \4749 , \215 );
and \U$5908 ( \6040 , \4922 , \213 );
nor \U$5909 ( \6041 , \6039 , \6040 );
xnor \U$5910 ( \6042 , \6041 , \222 );
xor \U$5911 ( \6043 , \6038 , \6042 );
xor \U$5912 ( \6044 , \6028 , \6043 );
xor \U$5913 ( \6045 , \6019 , \6044 );
xor \U$5914 ( \6046 , \6005 , \6045 );
xor \U$5915 ( \6047 , \5843 , \6046 );
xor \U$5916 ( \6048 , \5824 , \6047 );
and \U$5917 ( \6049 , \5584 , \5625 );
and \U$5918 ( \6050 , \5625 , \5806 );
and \U$5919 ( \6051 , \5584 , \5806 );
or \U$5920 ( \6052 , \6049 , \6050 , \6051 );
xor \U$5921 ( \6053 , \6048 , \6052 );
and \U$5922 ( \6054 , \5807 , \5811 );
and \U$5923 ( \6055 , \5812 , \5815 );
or \U$5924 ( \6056 , \6054 , \6055 );
xor \U$5925 ( \6057 , \6053 , \6056 );
buf \U$5926 ( \6058 , \6057 );
buf \U$5927 ( \6059 , \6058 );
and \U$5928 ( \6060 , \5828 , \5842 );
and \U$5929 ( \6061 , \5842 , \6046 );
and \U$5930 ( \6062 , \5828 , \6046 );
or \U$5931 ( \6063 , \6060 , \6061 , \6062 );
and \U$5932 ( \6064 , \5847 , \5851 );
and \U$5933 ( \6065 , \5851 , \5856 );
and \U$5934 ( \6066 , \5847 , \5856 );
or \U$5935 ( \6067 , \6064 , \6065 , \6066 );
and \U$5936 ( \6068 , \5871 , \5885 );
and \U$5937 ( \6069 , \5885 , \6003 );
and \U$5938 ( \6070 , \5871 , \6003 );
or \U$5939 ( \6071 , \6068 , \6069 , \6070 );
xor \U$5940 ( \6072 , \6067 , \6071 );
and \U$5941 ( \6073 , \6019 , \6044 );
xor \U$5942 ( \6074 , \6072 , \6073 );
xor \U$5943 ( \6075 , \6063 , \6074 );
and \U$5944 ( \6076 , \5832 , \5836 );
and \U$5945 ( \6077 , \5836 , \5841 );
and \U$5946 ( \6078 , \5832 , \5841 );
or \U$5947 ( \6079 , \6076 , \6077 , \6078 );
and \U$5948 ( \6080 , \5857 , \6004 );
and \U$5949 ( \6081 , \6004 , \6045 );
and \U$5950 ( \6082 , \5857 , \6045 );
or \U$5951 ( \6083 , \6080 , \6081 , \6082 );
xor \U$5952 ( \6084 , \6079 , \6083 );
and \U$5953 ( \6085 , \6009 , \6013 );
and \U$5954 ( \6086 , \6013 , \6018 );
and \U$5955 ( \6087 , \6009 , \6018 );
or \U$5956 ( \6088 , \6085 , \6086 , \6087 );
and \U$5957 ( \6089 , \6023 , \6027 );
and \U$5958 ( \6090 , \6027 , \6043 );
and \U$5959 ( \6091 , \6023 , \6043 );
or \U$5960 ( \6092 , \6089 , \6090 , \6091 );
xor \U$5961 ( \6093 , \6088 , \6092 );
and \U$5962 ( \6094 , \5930 , \5974 );
and \U$5963 ( \6095 , \5974 , \6002 );
and \U$5964 ( \6096 , \5930 , \6002 );
or \U$5965 ( \6097 , \6094 , \6095 , \6096 );
xor \U$5966 ( \6098 , \6093 , \6097 );
and \U$5967 ( \6099 , \6033 , \6037 );
and \U$5968 ( \6100 , \6037 , \6042 );
and \U$5969 ( \6101 , \6033 , \6042 );
or \U$5970 ( \6102 , \6099 , \6100 , \6101 );
and \U$5971 ( \6103 , \5934 , \5938 );
and \U$5972 ( \6104 , \5938 , \5943 );
and \U$5973 ( \6105 , \5934 , \5943 );
or \U$5974 ( \6106 , \6103 , \6104 , \6105 );
xor \U$5975 ( \6107 , \6102 , \6106 );
and \U$5976 ( \6108 , \5963 , \5967 );
and \U$5977 ( \6109 , \5967 , \5972 );
and \U$5978 ( \6110 , \5963 , \5972 );
or \U$5979 ( \6111 , \6108 , \6109 , \6110 );
xor \U$5980 ( \6112 , \6107 , \6111 );
and \U$5981 ( \6113 , \5904 , \5908 );
and \U$5982 ( \6114 , \5908 , \5913 );
and \U$5983 ( \6115 , \5904 , \5913 );
or \U$5984 ( \6116 , \6113 , \6114 , \6115 );
and \U$5985 ( \6117 , \5919 , \5923 );
and \U$5986 ( \6118 , \5923 , \5928 );
and \U$5987 ( \6119 , \5919 , \5928 );
or \U$5988 ( \6120 , \6117 , \6118 , \6119 );
xor \U$5989 ( \6121 , \6116 , \6120 );
and \U$5990 ( \6122 , \5948 , \5952 );
and \U$5991 ( \6123 , \5952 , \5957 );
and \U$5992 ( \6124 , \5948 , \5957 );
or \U$5993 ( \6125 , \6122 , \6123 , \6124 );
xor \U$5994 ( \6126 , \6121 , \6125 );
xor \U$5995 ( \6127 , \6112 , \6126 );
and \U$5996 ( \6128 , \5890 , \5894 );
and \U$5997 ( \6129 , \5894 , \5899 );
and \U$5998 ( \6130 , \5890 , \5899 );
or \U$5999 ( \6131 , \6128 , \6129 , \6130 );
and \U$6000 ( \6132 , \5988 , \5992 );
and \U$6001 ( \6133 , \5992 , \6000 );
and \U$6002 ( \6134 , \5988 , \6000 );
or \U$6003 ( \6135 , \6132 , \6133 , \6134 );
xor \U$6004 ( \6136 , \6131 , \6135 );
and \U$6005 ( \6137 , \150 , \5996 );
and \U$6006 ( \6138 , \158 , \5695 );
nor \U$6007 ( \6139 , \6137 , \6138 );
xnor \U$6008 ( \6140 , \6139 , \5687 );
xor \U$6009 ( \6141 , \6136 , \6140 );
buf \U$6010 ( \6142 , RIb5608b8_16);
xor \U$6011 ( \6143 , \6142 , \5683 );
nand \U$6012 ( \6144 , \166 , \6143 );
buf \U$6013 ( \6145 , RIb560930_15);
and \U$6014 ( \6146 , \6142 , \5683 );
not \U$6015 ( \6147 , \6146 );
and \U$6016 ( \6148 , \6145 , \6147 );
xnor \U$6017 ( \6149 , \6144 , \6148 );
and \U$6018 ( \6150 , \178 , \3357 );
and \U$6019 ( \6151 , \185 , \3255 );
nor \U$6020 ( \6152 , \6150 , \6151 );
xnor \U$6021 ( \6153 , \6152 , \3156 );
and \U$6022 ( \6154 , \189 , \3813 );
and \U$6023 ( \6155 , \197 , \3557 );
nor \U$6024 ( \6156 , \6154 , \6155 );
xnor \U$6025 ( \6157 , \6156 , \3562 );
xor \U$6026 ( \6158 , \6153 , \6157 );
and \U$6027 ( \6159 , \209 , \4132 );
and \U$6028 ( \6160 , \217 , \4012 );
nor \U$6029 ( \6161 , \6159 , \6160 );
xnor \U$6030 ( \6162 , \6161 , \3925 );
xor \U$6031 ( \6163 , \6158 , \6162 );
xor \U$6032 ( \6164 , \6149 , \6163 );
and \U$6033 ( \6165 , \224 , \4581 );
and \U$6034 ( \6166 , \232 , \4424 );
nor \U$6035 ( \6167 , \6165 , \6166 );
xnor \U$6036 ( \6168 , \6167 , \4377 );
and \U$6037 ( \6169 , \240 , \5011 );
and \U$6038 ( \6170 , \247 , \4878 );
nor \U$6039 ( \6171 , \6169 , \6170 );
xnor \U$6040 ( \6172 , \6171 , \4762 );
xor \U$6041 ( \6173 , \6168 , \6172 );
and \U$6042 ( \6174 , \134 , \5485 );
and \U$6043 ( \6175 , \143 , \5275 );
nor \U$6044 ( \6176 , \6174 , \6175 );
xnor \U$6045 ( \6177 , \6176 , \5169 );
xor \U$6046 ( \6178 , \6173 , \6177 );
xor \U$6047 ( \6179 , \6164 , \6178 );
xor \U$6048 ( \6180 , \6141 , \6179 );
and \U$6049 ( \6181 , \1802 , \1578 );
and \U$6050 ( \6182 , \1948 , \1431 );
nor \U$6051 ( \6183 , \6181 , \6182 );
xnor \U$6052 ( \6184 , \6183 , \1436 );
and \U$6053 ( \6185 , \1601 , \1824 );
and \U$6054 ( \6186 , \1684 , \1739 );
nor \U$6055 ( \6187 , \6185 , \6186 );
xnor \U$6056 ( \6188 , \6187 , \1697 );
xor \U$6057 ( \6189 , \6184 , \6188 );
and \U$6058 ( \6190 , \1333 , \2121 );
and \U$6059 ( \6191 , \1484 , \2008 );
nor \U$6060 ( \6192 , \6190 , \6191 );
xnor \U$6061 ( \6193 , \6192 , \1961 );
xor \U$6062 ( \6194 , \6189 , \6193 );
and \U$6063 ( \6195 , \2757 , \438 );
and \U$6064 ( \6196 , \2826 , \336 );
nor \U$6065 ( \6197 , \6195 , \6196 );
xnor \U$6066 ( \6198 , \6197 , \320 );
and \U$6067 ( \6199 , \2366 , \1086 );
and \U$6068 ( \6200 , \2521 , \508 );
nor \U$6069 ( \6201 , \6199 , \6200 );
xnor \U$6070 ( \6202 , \6201 , \487 );
xor \U$6071 ( \6203 , \6198 , \6202 );
and \U$6072 ( \6204 , \2090 , \1301 );
and \U$6073 ( \6205 , \2182 , \1246 );
nor \U$6074 ( \6206 , \6204 , \6205 );
xnor \U$6075 ( \6207 , \6206 , \1205 );
xor \U$6076 ( \6208 , \6203 , \6207 );
xor \U$6077 ( \6209 , \6194 , \6208 );
and \U$6078 ( \6210 , \1147 , \2400 );
and \U$6079 ( \6211 , \1192 , \2246 );
nor \U$6080 ( \6212 , \6210 , \6211 );
xnor \U$6081 ( \6213 , \6212 , \2195 );
and \U$6082 ( \6214 , \412 , \2669 );
and \U$6083 ( \6215 , \474 , \2538 );
nor \U$6084 ( \6216 , \6214 , \6215 );
xnor \U$6085 ( \6217 , \6216 , \2534 );
xor \U$6086 ( \6218 , \6213 , \6217 );
and \U$6087 ( \6219 , \261 , \3103 );
and \U$6088 ( \6220 , \307 , \2934 );
nor \U$6089 ( \6221 , \6219 , \6220 );
xnor \U$6090 ( \6222 , \6221 , \2839 );
xor \U$6091 ( \6223 , \6218 , \6222 );
xor \U$6092 ( \6224 , \6209 , \6223 );
xor \U$6093 ( \6225 , \6180 , \6224 );
xor \U$6094 ( \6226 , \6127 , \6225 );
xor \U$6095 ( \6227 , \6098 , \6226 );
and \U$6096 ( \6228 , \5861 , \5865 );
and \U$6097 ( \6229 , \5865 , \5870 );
and \U$6098 ( \6230 , \5861 , \5870 );
or \U$6099 ( \6231 , \6228 , \6229 , \6230 );
and \U$6100 ( \6232 , \5875 , \5879 );
and \U$6101 ( \6233 , \5879 , \5884 );
and \U$6102 ( \6234 , \5875 , \5884 );
or \U$6103 ( \6235 , \6232 , \6233 , \6234 );
xor \U$6104 ( \6236 , \6231 , \6235 );
and \U$6105 ( \6237 , \5979 , \5983 );
and \U$6106 ( \6238 , \5983 , \6001 );
and \U$6107 ( \6239 , \5979 , \6001 );
or \U$6108 ( \6240 , \6237 , \6238 , \6239 );
xor \U$6109 ( \6241 , \6236 , \6240 );
and \U$6110 ( \6242 , \5900 , \5914 );
and \U$6111 ( \6243 , \5914 , \5929 );
and \U$6112 ( \6244 , \5900 , \5929 );
or \U$6113 ( \6245 , \6242 , \6243 , \6244 );
and \U$6114 ( \6246 , \5944 , \5958 );
and \U$6115 ( \6247 , \5958 , \5973 );
and \U$6116 ( \6248 , \5944 , \5973 );
or \U$6117 ( \6249 , \6246 , \6247 , \6248 );
xor \U$6118 ( \6250 , \6245 , \6249 );
and \U$6119 ( \6251 , \3736 , \141 );
and \U$6120 ( \6252 , \3912 , \139 );
nor \U$6121 ( \6253 , \6251 , \6252 );
xnor \U$6122 ( \6254 , \6253 , \148 );
and \U$6123 ( \6255 , \3395 , \156 );
and \U$6124 ( \6256 , \3646 , \154 );
nor \U$6125 ( \6257 , \6255 , \6256 );
xnor \U$6126 ( \6258 , \6257 , \163 );
xor \U$6127 ( \6259 , \6254 , \6258 );
and \U$6128 ( \6260 , \3037 , \296 );
and \U$6129 ( \6261 , \3143 , \168 );
nor \U$6130 ( \6262 , \6260 , \6261 );
xnor \U$6131 ( \6263 , \6262 , \173 );
xor \U$6132 ( \6264 , \6259 , \6263 );
and \U$6133 ( \6265 , \4922 , \215 );
and \U$6134 ( \6266 , \5156 , \213 );
nor \U$6135 ( \6267 , \6265 , \6266 );
xnor \U$6136 ( \6268 , \6267 , \222 );
and \U$6137 ( \6269 , \4654 , \230 );
and \U$6138 ( \6270 , \4749 , \228 );
nor \U$6139 ( \6271 , \6269 , \6270 );
xnor \U$6140 ( \6272 , \6271 , \237 );
xor \U$6141 ( \6273 , \6268 , \6272 );
and \U$6142 ( \6274 , \4160 , \245 );
and \U$6143 ( \6275 , \4364 , \243 );
nor \U$6144 ( \6276 , \6274 , \6275 );
xnor \U$6145 ( \6277 , \6276 , \252 );
xor \U$6146 ( \6278 , \6273 , \6277 );
xor \U$6147 ( \6279 , \6264 , \6278 );
and \U$6148 ( \6280 , \6030 , \183 );
buf \U$6149 ( \6281 , RIb55eab8_80);
and \U$6150 ( \6282 , \6281 , \180 );
nor \U$6151 ( \6283 , \6280 , \6282 );
xnor \U$6152 ( \6284 , \6283 , \179 );
and \U$6153 ( \6285 , \5469 , \195 );
and \U$6154 ( \6286 , \5674 , \193 );
nor \U$6155 ( \6287 , \6285 , \6286 );
xnor \U$6156 ( \6288 , \6287 , \202 );
xor \U$6157 ( \6289 , \6284 , \6288 );
xor \U$6158 ( \6290 , \6289 , \6148 );
xor \U$6159 ( \6291 , \6279 , \6290 );
xor \U$6160 ( \6292 , \6250 , \6291 );
xor \U$6161 ( \6293 , \6241 , \6292 );
xor \U$6162 ( \6294 , \6227 , \6293 );
xor \U$6163 ( \6295 , \6084 , \6294 );
xor \U$6164 ( \6296 , \6075 , \6295 );
and \U$6165 ( \6297 , \5822 , \5823 );
and \U$6166 ( \6298 , \5823 , \6047 );
and \U$6167 ( \6299 , \5822 , \6047 );
or \U$6168 ( \6300 , \6297 , \6298 , \6299 );
xor \U$6169 ( \6301 , \6296 , \6300 );
and \U$6170 ( \6302 , \6048 , \6052 );
and \U$6171 ( \6303 , \6053 , \6056 );
or \U$6172 ( \6304 , \6302 , \6303 );
xor \U$6173 ( \6305 , \6301 , \6304 );
buf \U$6174 ( \6306 , \6305 );
buf \U$6175 ( \6307 , \6306 );
and \U$6176 ( \6308 , \6079 , \6083 );
and \U$6177 ( \6309 , \6083 , \6294 );
and \U$6178 ( \6310 , \6079 , \6294 );
or \U$6179 ( \6311 , \6308 , \6309 , \6310 );
and \U$6180 ( \6312 , \6088 , \6092 );
and \U$6181 ( \6313 , \6092 , \6097 );
and \U$6182 ( \6314 , \6088 , \6097 );
or \U$6183 ( \6315 , \6312 , \6313 , \6314 );
and \U$6184 ( \6316 , \6112 , \6126 );
and \U$6185 ( \6317 , \6126 , \6225 );
and \U$6186 ( \6318 , \6112 , \6225 );
or \U$6187 ( \6319 , \6316 , \6317 , \6318 );
xor \U$6188 ( \6320 , \6315 , \6319 );
and \U$6189 ( \6321 , \6241 , \6292 );
xor \U$6190 ( \6322 , \6320 , \6321 );
xor \U$6191 ( \6323 , \6311 , \6322 );
and \U$6192 ( \6324 , \6067 , \6071 );
and \U$6193 ( \6325 , \6071 , \6073 );
and \U$6194 ( \6326 , \6067 , \6073 );
or \U$6195 ( \6327 , \6324 , \6325 , \6326 );
and \U$6196 ( \6328 , \6098 , \6226 );
and \U$6197 ( \6329 , \6226 , \6293 );
and \U$6198 ( \6330 , \6098 , \6293 );
or \U$6199 ( \6331 , \6328 , \6329 , \6330 );
xor \U$6200 ( \6332 , \6327 , \6331 );
and \U$6201 ( \6333 , \6131 , \6135 );
and \U$6202 ( \6334 , \6135 , \6140 );
and \U$6203 ( \6335 , \6131 , \6140 );
or \U$6204 ( \6336 , \6333 , \6334 , \6335 );
and \U$6205 ( \6337 , \6102 , \6106 );
and \U$6206 ( \6338 , \6106 , \6111 );
and \U$6207 ( \6339 , \6102 , \6111 );
or \U$6208 ( \6340 , \6337 , \6338 , \6339 );
xor \U$6209 ( \6341 , \6336 , \6340 );
and \U$6210 ( \6342 , \6116 , \6120 );
and \U$6211 ( \6343 , \6120 , \6125 );
and \U$6212 ( \6344 , \6116 , \6125 );
or \U$6213 ( \6345 , \6342 , \6343 , \6344 );
xor \U$6214 ( \6346 , \6341 , \6345 );
and \U$6215 ( \6347 , \6231 , \6235 );
and \U$6216 ( \6348 , \6235 , \6240 );
and \U$6217 ( \6349 , \6231 , \6240 );
or \U$6218 ( \6350 , \6347 , \6348 , \6349 );
and \U$6219 ( \6351 , \6245 , \6249 );
and \U$6220 ( \6352 , \6249 , \6291 );
and \U$6221 ( \6353 , \6245 , \6291 );
or \U$6222 ( \6354 , \6351 , \6352 , \6353 );
xor \U$6223 ( \6355 , \6350 , \6354 );
and \U$6224 ( \6356 , \6141 , \6179 );
and \U$6225 ( \6357 , \6179 , \6224 );
and \U$6226 ( \6358 , \6141 , \6224 );
or \U$6227 ( \6359 , \6356 , \6357 , \6358 );
xor \U$6228 ( \6360 , \6355 , \6359 );
xor \U$6229 ( \6361 , \6346 , \6360 );
and \U$6230 ( \6362 , \6264 , \6278 );
and \U$6231 ( \6363 , \6278 , \6290 );
and \U$6232 ( \6364 , \6264 , \6290 );
or \U$6233 ( \6365 , \6362 , \6363 , \6364 );
and \U$6234 ( \6366 , \6149 , \6163 );
and \U$6235 ( \6367 , \6163 , \6178 );
and \U$6236 ( \6368 , \6149 , \6178 );
or \U$6237 ( \6369 , \6366 , \6367 , \6368 );
xor \U$6238 ( \6370 , \6365 , \6369 );
and \U$6239 ( \6371 , \6194 , \6208 );
and \U$6240 ( \6372 , \6208 , \6223 );
and \U$6241 ( \6373 , \6194 , \6223 );
or \U$6242 ( \6374 , \6371 , \6372 , \6373 );
xor \U$6243 ( \6375 , \6370 , \6374 );
and \U$6244 ( \6376 , \6254 , \6258 );
and \U$6245 ( \6377 , \6258 , \6263 );
and \U$6246 ( \6378 , \6254 , \6263 );
or \U$6247 ( \6379 , \6376 , \6377 , \6378 );
and \U$6248 ( \6380 , \6268 , \6272 );
and \U$6249 ( \6381 , \6272 , \6277 );
and \U$6250 ( \6382 , \6268 , \6277 );
or \U$6251 ( \6383 , \6380 , \6381 , \6382 );
xor \U$6252 ( \6384 , \6379 , \6383 );
and \U$6253 ( \6385 , \6284 , \6288 );
and \U$6254 ( \6386 , \6288 , \6148 );
and \U$6255 ( \6387 , \6284 , \6148 );
or \U$6256 ( \6388 , \6385 , \6386 , \6387 );
xor \U$6257 ( \6389 , \6384 , \6388 );
and \U$6258 ( \6390 , \6153 , \6157 );
and \U$6259 ( \6391 , \6157 , \6162 );
and \U$6260 ( \6392 , \6153 , \6162 );
or \U$6261 ( \6393 , \6390 , \6391 , \6392 );
and \U$6262 ( \6394 , \6168 , \6172 );
and \U$6263 ( \6395 , \6172 , \6177 );
and \U$6264 ( \6396 , \6168 , \6177 );
or \U$6265 ( \6397 , \6394 , \6395 , \6396 );
xor \U$6266 ( \6398 , \6393 , \6397 );
xor \U$6267 ( \6399 , \6145 , \6142 );
not \U$6268 ( \6400 , \6143 );
and \U$6269 ( \6401 , \6399 , \6400 );
and \U$6270 ( \6402 , \166 , \6401 );
and \U$6271 ( \6403 , \150 , \6143 );
nor \U$6272 ( \6404 , \6402 , \6403 );
xnor \U$6273 ( \6405 , \6404 , \6148 );
xor \U$6274 ( \6406 , \6398 , \6405 );
xor \U$6275 ( \6407 , \6389 , \6406 );
and \U$6276 ( \6408 , \6184 , \6188 );
and \U$6277 ( \6409 , \6188 , \6193 );
and \U$6278 ( \6410 , \6184 , \6193 );
or \U$6279 ( \6411 , \6408 , \6409 , \6410 );
and \U$6280 ( \6412 , \6198 , \6202 );
and \U$6281 ( \6413 , \6202 , \6207 );
and \U$6282 ( \6414 , \6198 , \6207 );
or \U$6283 ( \6415 , \6412 , \6413 , \6414 );
xor \U$6284 ( \6416 , \6411 , \6415 );
and \U$6285 ( \6417 , \6213 , \6217 );
and \U$6286 ( \6418 , \6217 , \6222 );
and \U$6287 ( \6419 , \6213 , \6222 );
or \U$6288 ( \6420 , \6417 , \6418 , \6419 );
xor \U$6289 ( \6421 , \6416 , \6420 );
xor \U$6290 ( \6422 , \6407 , \6421 );
xor \U$6291 ( \6423 , \6375 , \6422 );
and \U$6292 ( \6424 , \247 , \5011 );
and \U$6293 ( \6425 , \224 , \4878 );
nor \U$6294 ( \6426 , \6424 , \6425 );
xnor \U$6295 ( \6427 , \6426 , \4762 );
and \U$6296 ( \6428 , \143 , \5485 );
and \U$6297 ( \6429 , \240 , \5275 );
nor \U$6298 ( \6430 , \6428 , \6429 );
xnor \U$6299 ( \6431 , \6430 , \5169 );
xor \U$6300 ( \6432 , \6427 , \6431 );
and \U$6301 ( \6433 , \158 , \5996 );
and \U$6302 ( \6434 , \134 , \5695 );
nor \U$6303 ( \6435 , \6433 , \6434 );
xnor \U$6304 ( \6436 , \6435 , \5687 );
xor \U$6305 ( \6437 , \6432 , \6436 );
and \U$6306 ( \6438 , \474 , \2669 );
and \U$6307 ( \6439 , \1147 , \2538 );
nor \U$6308 ( \6440 , \6438 , \6439 );
xnor \U$6309 ( \6441 , \6440 , \2534 );
and \U$6310 ( \6442 , \307 , \3103 );
and \U$6311 ( \6443 , \412 , \2934 );
nor \U$6312 ( \6444 , \6442 , \6443 );
xnor \U$6313 ( \6445 , \6444 , \2839 );
xor \U$6314 ( \6446 , \6441 , \6445 );
and \U$6315 ( \6447 , \185 , \3357 );
and \U$6316 ( \6448 , \261 , \3255 );
nor \U$6317 ( \6449 , \6447 , \6448 );
xnor \U$6318 ( \6450 , \6449 , \3156 );
xor \U$6319 ( \6451 , \6446 , \6450 );
xor \U$6320 ( \6452 , \6437 , \6451 );
and \U$6321 ( \6453 , \197 , \3813 );
and \U$6322 ( \6454 , \178 , \3557 );
nor \U$6323 ( \6455 , \6453 , \6454 );
xnor \U$6324 ( \6456 , \6455 , \3562 );
and \U$6325 ( \6457 , \217 , \4132 );
and \U$6326 ( \6458 , \189 , \4012 );
nor \U$6327 ( \6459 , \6457 , \6458 );
xnor \U$6328 ( \6460 , \6459 , \3925 );
xor \U$6329 ( \6461 , \6456 , \6460 );
and \U$6330 ( \6462 , \232 , \4581 );
and \U$6331 ( \6463 , \209 , \4424 );
nor \U$6332 ( \6464 , \6462 , \6463 );
xnor \U$6333 ( \6465 , \6464 , \4377 );
xor \U$6334 ( \6466 , \6461 , \6465 );
xor \U$6335 ( \6467 , \6452 , \6466 );
and \U$6336 ( \6468 , \1684 , \1824 );
and \U$6337 ( \6469 , \1802 , \1739 );
nor \U$6338 ( \6470 , \6468 , \6469 );
xnor \U$6339 ( \6471 , \6470 , \1697 );
and \U$6340 ( \6472 , \1484 , \2121 );
and \U$6341 ( \6473 , \1601 , \2008 );
nor \U$6342 ( \6474 , \6472 , \6473 );
xnor \U$6343 ( \6475 , \6474 , \1961 );
xor \U$6344 ( \6476 , \6471 , \6475 );
and \U$6345 ( \6477 , \1192 , \2400 );
and \U$6346 ( \6478 , \1333 , \2246 );
nor \U$6347 ( \6479 , \6477 , \6478 );
xnor \U$6348 ( \6480 , \6479 , \2195 );
xor \U$6349 ( \6481 , \6476 , \6480 );
and \U$6350 ( \6482 , \2521 , \1086 );
and \U$6351 ( \6483 , \2757 , \508 );
nor \U$6352 ( \6484 , \6482 , \6483 );
xnor \U$6353 ( \6485 , \6484 , \487 );
and \U$6354 ( \6486 , \2182 , \1301 );
and \U$6355 ( \6487 , \2366 , \1246 );
nor \U$6356 ( \6488 , \6486 , \6487 );
xnor \U$6357 ( \6489 , \6488 , \1205 );
xor \U$6358 ( \6490 , \6485 , \6489 );
and \U$6359 ( \6491 , \1948 , \1578 );
and \U$6360 ( \6492 , \2090 , \1431 );
nor \U$6361 ( \6493 , \6491 , \6492 );
xnor \U$6362 ( \6494 , \6493 , \1436 );
xor \U$6363 ( \6495 , \6490 , \6494 );
xor \U$6364 ( \6496 , \6481 , \6495 );
and \U$6365 ( \6497 , \3646 , \156 );
and \U$6366 ( \6498 , \3736 , \154 );
nor \U$6367 ( \6499 , \6497 , \6498 );
xnor \U$6368 ( \6500 , \6499 , \163 );
and \U$6369 ( \6501 , \3143 , \296 );
and \U$6370 ( \6502 , \3395 , \168 );
nor \U$6371 ( \6503 , \6501 , \6502 );
xnor \U$6372 ( \6504 , \6503 , \173 );
xor \U$6373 ( \6505 , \6500 , \6504 );
and \U$6374 ( \6506 , \2826 , \438 );
and \U$6375 ( \6507 , \3037 , \336 );
nor \U$6376 ( \6508 , \6506 , \6507 );
xnor \U$6377 ( \6509 , \6508 , \320 );
xor \U$6378 ( \6510 , \6505 , \6509 );
xor \U$6379 ( \6511 , \6496 , \6510 );
xor \U$6380 ( \6512 , \6467 , \6511 );
and \U$6381 ( \6513 , \6281 , \183 );
buf \U$6382 ( \6514 , RIb55eb30_79);
and \U$6383 ( \6515 , \6514 , \180 );
nor \U$6384 ( \6516 , \6513 , \6515 );
xnor \U$6385 ( \6517 , \6516 , \179 );
and \U$6386 ( \6518 , \5674 , \195 );
and \U$6387 ( \6519 , \6030 , \193 );
nor \U$6388 ( \6520 , \6518 , \6519 );
xnor \U$6389 ( \6521 , \6520 , \202 );
xor \U$6390 ( \6522 , \6517 , \6521 );
and \U$6391 ( \6523 , \5156 , \215 );
and \U$6392 ( \6524 , \5469 , \213 );
nor \U$6393 ( \6525 , \6523 , \6524 );
xnor \U$6394 ( \6526 , \6525 , \222 );
xor \U$6395 ( \6527 , \6522 , \6526 );
and \U$6396 ( \6528 , \4749 , \230 );
and \U$6397 ( \6529 , \4922 , \228 );
nor \U$6398 ( \6530 , \6528 , \6529 );
xnor \U$6399 ( \6531 , \6530 , \237 );
and \U$6400 ( \6532 , \4364 , \245 );
and \U$6401 ( \6533 , \4654 , \243 );
nor \U$6402 ( \6534 , \6532 , \6533 );
xnor \U$6403 ( \6535 , \6534 , \252 );
xor \U$6404 ( \6536 , \6531 , \6535 );
and \U$6405 ( \6537 , \3912 , \141 );
and \U$6406 ( \6538 , \4160 , \139 );
nor \U$6407 ( \6539 , \6537 , \6538 );
xnor \U$6408 ( \6540 , \6539 , \148 );
xor \U$6409 ( \6541 , \6536 , \6540 );
xor \U$6410 ( \6542 , \6527 , \6541 );
xor \U$6411 ( \6543 , \6512 , \6542 );
xor \U$6412 ( \6544 , \6423 , \6543 );
xor \U$6413 ( \6545 , \6361 , \6544 );
xor \U$6414 ( \6546 , \6332 , \6545 );
xor \U$6415 ( \6547 , \6323 , \6546 );
and \U$6416 ( \6548 , \6063 , \6074 );
and \U$6417 ( \6549 , \6074 , \6295 );
and \U$6418 ( \6550 , \6063 , \6295 );
or \U$6419 ( \6551 , \6548 , \6549 , \6550 );
xor \U$6420 ( \6552 , \6547 , \6551 );
and \U$6421 ( \6553 , \6296 , \6300 );
and \U$6422 ( \6554 , \6301 , \6304 );
or \U$6423 ( \6555 , \6553 , \6554 );
xor \U$6424 ( \6556 , \6552 , \6555 );
buf \U$6425 ( \6557 , \6556 );
buf \U$6426 ( \6558 , \6557 );
and \U$6427 ( \6559 , \6327 , \6331 );
and \U$6428 ( \6560 , \6331 , \6545 );
and \U$6429 ( \6561 , \6327 , \6545 );
or \U$6430 ( \6562 , \6559 , \6560 , \6561 );
and \U$6431 ( \6563 , \6350 , \6354 );
and \U$6432 ( \6564 , \6354 , \6359 );
and \U$6433 ( \6565 , \6350 , \6359 );
or \U$6434 ( \6566 , \6563 , \6564 , \6565 );
and \U$6435 ( \6567 , \6375 , \6422 );
and \U$6436 ( \6568 , \6422 , \6543 );
and \U$6437 ( \6569 , \6375 , \6543 );
or \U$6438 ( \6570 , \6567 , \6568 , \6569 );
xor \U$6439 ( \6571 , \6566 , \6570 );
and \U$6440 ( \6572 , \6437 , \6451 );
and \U$6441 ( \6573 , \6451 , \6466 );
and \U$6442 ( \6574 , \6437 , \6466 );
or \U$6443 ( \6575 , \6572 , \6573 , \6574 );
and \U$6444 ( \6576 , \6481 , \6495 );
and \U$6445 ( \6577 , \6495 , \6510 );
and \U$6446 ( \6578 , \6481 , \6510 );
or \U$6447 ( \6579 , \6576 , \6577 , \6578 );
xor \U$6448 ( \6580 , \6575 , \6579 );
and \U$6449 ( \6581 , \6527 , \6541 );
xor \U$6450 ( \6582 , \6580 , \6581 );
xor \U$6451 ( \6583 , \6571 , \6582 );
xor \U$6452 ( \6584 , \6562 , \6583 );
and \U$6453 ( \6585 , \6315 , \6319 );
and \U$6454 ( \6586 , \6319 , \6321 );
and \U$6455 ( \6587 , \6315 , \6321 );
or \U$6456 ( \6588 , \6585 , \6586 , \6587 );
and \U$6457 ( \6589 , \6346 , \6360 );
and \U$6458 ( \6590 , \6360 , \6544 );
and \U$6459 ( \6591 , \6346 , \6544 );
or \U$6460 ( \6592 , \6589 , \6590 , \6591 );
xor \U$6461 ( \6593 , \6588 , \6592 );
and \U$6462 ( \6594 , \6379 , \6383 );
and \U$6463 ( \6595 , \6383 , \6388 );
and \U$6464 ( \6596 , \6379 , \6388 );
or \U$6465 ( \6597 , \6594 , \6595 , \6596 );
and \U$6466 ( \6598 , \6393 , \6397 );
and \U$6467 ( \6599 , \6397 , \6405 );
and \U$6468 ( \6600 , \6393 , \6405 );
or \U$6469 ( \6601 , \6598 , \6599 , \6600 );
xor \U$6470 ( \6602 , \6597 , \6601 );
and \U$6471 ( \6603 , \6411 , \6415 );
and \U$6472 ( \6604 , \6415 , \6420 );
and \U$6473 ( \6605 , \6411 , \6420 );
or \U$6474 ( \6606 , \6603 , \6604 , \6605 );
xor \U$6475 ( \6607 , \6602 , \6606 );
and \U$6476 ( \6608 , \6365 , \6369 );
and \U$6477 ( \6609 , \6369 , \6374 );
and \U$6478 ( \6610 , \6365 , \6374 );
or \U$6479 ( \6611 , \6608 , \6609 , \6610 );
and \U$6480 ( \6612 , \6336 , \6340 );
and \U$6481 ( \6613 , \6340 , \6345 );
and \U$6482 ( \6614 , \6336 , \6345 );
or \U$6483 ( \6615 , \6612 , \6613 , \6614 );
xor \U$6484 ( \6616 , \6611 , \6615 );
and \U$6485 ( \6617 , \6467 , \6511 );
and \U$6486 ( \6618 , \6511 , \6542 );
and \U$6487 ( \6619 , \6467 , \6542 );
or \U$6488 ( \6620 , \6617 , \6618 , \6619 );
xor \U$6489 ( \6621 , \6616 , \6620 );
xor \U$6490 ( \6622 , \6607 , \6621 );
and \U$6491 ( \6623 , \6389 , \6406 );
and \U$6492 ( \6624 , \6406 , \6421 );
and \U$6493 ( \6625 , \6389 , \6421 );
or \U$6494 ( \6626 , \6623 , \6624 , \6625 );
and \U$6495 ( \6627 , \6500 , \6504 );
and \U$6496 ( \6628 , \6504 , \6509 );
and \U$6497 ( \6629 , \6500 , \6509 );
or \U$6498 ( \6630 , \6627 , \6628 , \6629 );
and \U$6499 ( \6631 , \6517 , \6521 );
and \U$6500 ( \6632 , \6521 , \6526 );
and \U$6501 ( \6633 , \6517 , \6526 );
or \U$6502 ( \6634 , \6631 , \6632 , \6633 );
xor \U$6503 ( \6635 , \6630 , \6634 );
and \U$6504 ( \6636 , \6531 , \6535 );
and \U$6505 ( \6637 , \6535 , \6540 );
and \U$6506 ( \6638 , \6531 , \6540 );
or \U$6507 ( \6639 , \6636 , \6637 , \6638 );
xor \U$6508 ( \6640 , \6635 , \6639 );
and \U$6509 ( \6641 , \6471 , \6475 );
and \U$6510 ( \6642 , \6475 , \6480 );
and \U$6511 ( \6643 , \6471 , \6480 );
or \U$6512 ( \6644 , \6641 , \6642 , \6643 );
and \U$6513 ( \6645 , \6485 , \6489 );
and \U$6514 ( \6646 , \6489 , \6494 );
and \U$6515 ( \6647 , \6485 , \6494 );
or \U$6516 ( \6648 , \6645 , \6646 , \6647 );
xor \U$6517 ( \6649 , \6644 , \6648 );
and \U$6518 ( \6650 , \6441 , \6445 );
and \U$6519 ( \6651 , \6445 , \6450 );
and \U$6520 ( \6652 , \6441 , \6450 );
or \U$6521 ( \6653 , \6650 , \6651 , \6652 );
xor \U$6522 ( \6654 , \6649 , \6653 );
xor \U$6523 ( \6655 , \6640 , \6654 );
and \U$6524 ( \6656 , \6427 , \6431 );
and \U$6525 ( \6657 , \6431 , \6436 );
and \U$6526 ( \6658 , \6427 , \6436 );
or \U$6527 ( \6659 , \6656 , \6657 , \6658 );
and \U$6528 ( \6660 , \6456 , \6460 );
and \U$6529 ( \6661 , \6460 , \6465 );
and \U$6530 ( \6662 , \6456 , \6465 );
or \U$6531 ( \6663 , \6660 , \6661 , \6662 );
xor \U$6532 ( \6664 , \6659 , \6663 );
and \U$6533 ( \6665 , \134 , \5996 );
and \U$6534 ( \6666 , \143 , \5695 );
nor \U$6535 ( \6667 , \6665 , \6666 );
xnor \U$6536 ( \6668 , \6667 , \5687 );
and \U$6537 ( \6669 , \150 , \6401 );
and \U$6538 ( \6670 , \158 , \6143 );
nor \U$6539 ( \6671 , \6669 , \6670 );
xnor \U$6540 ( \6672 , \6671 , \6148 );
xor \U$6541 ( \6673 , \6668 , \6672 );
buf \U$6542 ( \6674 , RIb5609a8_14);
xor \U$6543 ( \6675 , \6674 , \6145 );
nand \U$6544 ( \6676 , \166 , \6675 );
buf \U$6545 ( \6677 , RIb560a20_13);
and \U$6546 ( \6678 , \6674 , \6145 );
not \U$6547 ( \6679 , \6678 );
and \U$6548 ( \6680 , \6677 , \6679 );
xnor \U$6549 ( \6681 , \6676 , \6680 );
xor \U$6550 ( \6682 , \6673 , \6681 );
xor \U$6551 ( \6683 , \6664 , \6682 );
xor \U$6552 ( \6684 , \6655 , \6683 );
xor \U$6553 ( \6685 , \6626 , \6684 );
and \U$6554 ( \6686 , \261 , \3357 );
and \U$6555 ( \6687 , \307 , \3255 );
nor \U$6556 ( \6688 , \6686 , \6687 );
xnor \U$6557 ( \6689 , \6688 , \3156 );
and \U$6558 ( \6690 , \178 , \3813 );
and \U$6559 ( \6691 , \185 , \3557 );
nor \U$6560 ( \6692 , \6690 , \6691 );
xnor \U$6561 ( \6693 , \6692 , \3562 );
xor \U$6562 ( \6694 , \6689 , \6693 );
and \U$6563 ( \6695 , \189 , \4132 );
and \U$6564 ( \6696 , \197 , \4012 );
nor \U$6565 ( \6697 , \6695 , \6696 );
xnor \U$6566 ( \6698 , \6697 , \3925 );
xor \U$6567 ( \6699 , \6694 , \6698 );
and \U$6568 ( \6700 , \1333 , \2400 );
and \U$6569 ( \6701 , \1484 , \2246 );
nor \U$6570 ( \6702 , \6700 , \6701 );
xnor \U$6571 ( \6703 , \6702 , \2195 );
and \U$6572 ( \6704 , \1147 , \2669 );
and \U$6573 ( \6705 , \1192 , \2538 );
nor \U$6574 ( \6706 , \6704 , \6705 );
xnor \U$6575 ( \6707 , \6706 , \2534 );
xor \U$6576 ( \6708 , \6703 , \6707 );
and \U$6577 ( \6709 , \412 , \3103 );
and \U$6578 ( \6710 , \474 , \2934 );
nor \U$6579 ( \6711 , \6709 , \6710 );
xnor \U$6580 ( \6712 , \6711 , \2839 );
xor \U$6581 ( \6713 , \6708 , \6712 );
xor \U$6582 ( \6714 , \6699 , \6713 );
and \U$6583 ( \6715 , \209 , \4581 );
and \U$6584 ( \6716 , \217 , \4424 );
nor \U$6585 ( \6717 , \6715 , \6716 );
xnor \U$6586 ( \6718 , \6717 , \4377 );
and \U$6587 ( \6719 , \224 , \5011 );
and \U$6588 ( \6720 , \232 , \4878 );
nor \U$6589 ( \6721 , \6719 , \6720 );
xnor \U$6590 ( \6722 , \6721 , \4762 );
xor \U$6591 ( \6723 , \6718 , \6722 );
and \U$6592 ( \6724 , \240 , \5485 );
and \U$6593 ( \6725 , \247 , \5275 );
nor \U$6594 ( \6726 , \6724 , \6725 );
xnor \U$6595 ( \6727 , \6726 , \5169 );
xor \U$6596 ( \6728 , \6723 , \6727 );
xor \U$6597 ( \6729 , \6714 , \6728 );
and \U$6598 ( \6730 , \2090 , \1578 );
and \U$6599 ( \6731 , \2182 , \1431 );
nor \U$6600 ( \6732 , \6730 , \6731 );
xnor \U$6601 ( \6733 , \6732 , \1436 );
and \U$6602 ( \6734 , \1802 , \1824 );
and \U$6603 ( \6735 , \1948 , \1739 );
nor \U$6604 ( \6736 , \6734 , \6735 );
xnor \U$6605 ( \6737 , \6736 , \1697 );
xor \U$6606 ( \6738 , \6733 , \6737 );
and \U$6607 ( \6739 , \1601 , \2121 );
and \U$6608 ( \6740 , \1684 , \2008 );
nor \U$6609 ( \6741 , \6739 , \6740 );
xnor \U$6610 ( \6742 , \6741 , \1961 );
xor \U$6611 ( \6743 , \6738 , \6742 );
and \U$6612 ( \6744 , \3037 , \438 );
and \U$6613 ( \6745 , \3143 , \336 );
nor \U$6614 ( \6746 , \6744 , \6745 );
xnor \U$6615 ( \6747 , \6746 , \320 );
and \U$6616 ( \6748 , \2757 , \1086 );
and \U$6617 ( \6749 , \2826 , \508 );
nor \U$6618 ( \6750 , \6748 , \6749 );
xnor \U$6619 ( \6751 , \6750 , \487 );
xor \U$6620 ( \6752 , \6747 , \6751 );
and \U$6621 ( \6753 , \2366 , \1301 );
and \U$6622 ( \6754 , \2521 , \1246 );
nor \U$6623 ( \6755 , \6753 , \6754 );
xnor \U$6624 ( \6756 , \6755 , \1205 );
xor \U$6625 ( \6757 , \6752 , \6756 );
xor \U$6626 ( \6758 , \6743 , \6757 );
and \U$6627 ( \6759 , \4160 , \141 );
and \U$6628 ( \6760 , \4364 , \139 );
nor \U$6629 ( \6761 , \6759 , \6760 );
xnor \U$6630 ( \6762 , \6761 , \148 );
and \U$6631 ( \6763 , \3736 , \156 );
and \U$6632 ( \6764 , \3912 , \154 );
nor \U$6633 ( \6765 , \6763 , \6764 );
xnor \U$6634 ( \6766 , \6765 , \163 );
xor \U$6635 ( \6767 , \6762 , \6766 );
and \U$6636 ( \6768 , \3395 , \296 );
and \U$6637 ( \6769 , \3646 , \168 );
nor \U$6638 ( \6770 , \6768 , \6769 );
xnor \U$6639 ( \6771 , \6770 , \173 );
xor \U$6640 ( \6772 , \6767 , \6771 );
xor \U$6641 ( \6773 , \6758 , \6772 );
xor \U$6642 ( \6774 , \6729 , \6773 );
and \U$6643 ( \6775 , \5469 , \215 );
and \U$6644 ( \6776 , \5674 , \213 );
nor \U$6645 ( \6777 , \6775 , \6776 );
xnor \U$6646 ( \6778 , \6777 , \222 );
and \U$6647 ( \6779 , \4922 , \230 );
and \U$6648 ( \6780 , \5156 , \228 );
nor \U$6649 ( \6781 , \6779 , \6780 );
xnor \U$6650 ( \6782 , \6781 , \237 );
xor \U$6651 ( \6783 , \6778 , \6782 );
and \U$6652 ( \6784 , \4654 , \245 );
and \U$6653 ( \6785 , \4749 , \243 );
nor \U$6654 ( \6786 , \6784 , \6785 );
xnor \U$6655 ( \6787 , \6786 , \252 );
xor \U$6656 ( \6788 , \6783 , \6787 );
and \U$6657 ( \6789 , \6514 , \183 );
buf \U$6658 ( \6790 , RIb55eba8_78);
and \U$6659 ( \6791 , \6790 , \180 );
nor \U$6660 ( \6792 , \6789 , \6791 );
xnor \U$6661 ( \6793 , \6792 , \179 );
and \U$6662 ( \6794 , \6030 , \195 );
and \U$6663 ( \6795 , \6281 , \193 );
nor \U$6664 ( \6796 , \6794 , \6795 );
xnor \U$6665 ( \6797 , \6796 , \202 );
xor \U$6666 ( \6798 , \6793 , \6797 );
xor \U$6667 ( \6799 , \6798 , \6680 );
xor \U$6668 ( \6800 , \6788 , \6799 );
xor \U$6669 ( \6801 , \6774 , \6800 );
xor \U$6670 ( \6802 , \6685 , \6801 );
xor \U$6671 ( \6803 , \6622 , \6802 );
xor \U$6672 ( \6804 , \6593 , \6803 );
xor \U$6673 ( \6805 , \6584 , \6804 );
and \U$6674 ( \6806 , \6311 , \6322 );
and \U$6675 ( \6807 , \6322 , \6546 );
and \U$6676 ( \6808 , \6311 , \6546 );
or \U$6677 ( \6809 , \6806 , \6807 , \6808 );
xor \U$6678 ( \6810 , \6805 , \6809 );
and \U$6679 ( \6811 , \6547 , \6551 );
and \U$6680 ( \6812 , \6552 , \6555 );
or \U$6681 ( \6813 , \6811 , \6812 );
xor \U$6682 ( \6814 , \6810 , \6813 );
buf \U$6683 ( \6815 , \6814 );
buf \U$6684 ( \6816 , \6815 );
and \U$6685 ( \6817 , \6588 , \6592 );
and \U$6686 ( \6818 , \6592 , \6803 );
and \U$6687 ( \6819 , \6588 , \6803 );
or \U$6688 ( \6820 , \6817 , \6818 , \6819 );
and \U$6689 ( \6821 , \6611 , \6615 );
and \U$6690 ( \6822 , \6615 , \6620 );
and \U$6691 ( \6823 , \6611 , \6620 );
or \U$6692 ( \6824 , \6821 , \6822 , \6823 );
and \U$6693 ( \6825 , \6626 , \6684 );
and \U$6694 ( \6826 , \6684 , \6801 );
and \U$6695 ( \6827 , \6626 , \6801 );
or \U$6696 ( \6828 , \6825 , \6826 , \6827 );
xor \U$6697 ( \6829 , \6824 , \6828 );
and \U$6698 ( \6830 , \6699 , \6713 );
and \U$6699 ( \6831 , \6713 , \6728 );
and \U$6700 ( \6832 , \6699 , \6728 );
or \U$6701 ( \6833 , \6830 , \6831 , \6832 );
and \U$6702 ( \6834 , \6743 , \6757 );
and \U$6703 ( \6835 , \6757 , \6772 );
and \U$6704 ( \6836 , \6743 , \6772 );
or \U$6705 ( \6837 , \6834 , \6835 , \6836 );
xor \U$6706 ( \6838 , \6833 , \6837 );
and \U$6707 ( \6839 , \6788 , \6799 );
xor \U$6708 ( \6840 , \6838 , \6839 );
xor \U$6709 ( \6841 , \6829 , \6840 );
xor \U$6710 ( \6842 , \6820 , \6841 );
and \U$6711 ( \6843 , \6566 , \6570 );
and \U$6712 ( \6844 , \6570 , \6582 );
and \U$6713 ( \6845 , \6566 , \6582 );
or \U$6714 ( \6846 , \6843 , \6844 , \6845 );
and \U$6715 ( \6847 , \6607 , \6621 );
and \U$6716 ( \6848 , \6621 , \6802 );
and \U$6717 ( \6849 , \6607 , \6802 );
or \U$6718 ( \6850 , \6847 , \6848 , \6849 );
xor \U$6719 ( \6851 , \6846 , \6850 );
and \U$6720 ( \6852 , \6630 , \6634 );
and \U$6721 ( \6853 , \6634 , \6639 );
and \U$6722 ( \6854 , \6630 , \6639 );
or \U$6723 ( \6855 , \6852 , \6853 , \6854 );
and \U$6724 ( \6856 , \6644 , \6648 );
and \U$6725 ( \6857 , \6648 , \6653 );
and \U$6726 ( \6858 , \6644 , \6653 );
or \U$6727 ( \6859 , \6856 , \6857 , \6858 );
xor \U$6728 ( \6860 , \6855 , \6859 );
and \U$6729 ( \6861 , \6659 , \6663 );
and \U$6730 ( \6862 , \6663 , \6682 );
and \U$6731 ( \6863 , \6659 , \6682 );
or \U$6732 ( \6864 , \6861 , \6862 , \6863 );
xor \U$6733 ( \6865 , \6860 , \6864 );
and \U$6734 ( \6866 , \6597 , \6601 );
and \U$6735 ( \6867 , \6601 , \6606 );
and \U$6736 ( \6868 , \6597 , \6606 );
or \U$6737 ( \6869 , \6866 , \6867 , \6868 );
and \U$6738 ( \6870 , \6575 , \6579 );
and \U$6739 ( \6871 , \6579 , \6581 );
and \U$6740 ( \6872 , \6575 , \6581 );
or \U$6741 ( \6873 , \6870 , \6871 , \6872 );
xor \U$6742 ( \6874 , \6869 , \6873 );
and \U$6743 ( \6875 , \6729 , \6773 );
and \U$6744 ( \6876 , \6773 , \6800 );
and \U$6745 ( \6877 , \6729 , \6800 );
or \U$6746 ( \6878 , \6875 , \6876 , \6877 );
xor \U$6747 ( \6879 , \6874 , \6878 );
xor \U$6748 ( \6880 , \6865 , \6879 );
and \U$6749 ( \6881 , \6640 , \6654 );
and \U$6750 ( \6882 , \6654 , \6683 );
and \U$6751 ( \6883 , \6640 , \6683 );
or \U$6752 ( \6884 , \6881 , \6882 , \6883 );
and \U$6753 ( \6885 , \6733 , \6737 );
and \U$6754 ( \6886 , \6737 , \6742 );
and \U$6755 ( \6887 , \6733 , \6742 );
or \U$6756 ( \6888 , \6885 , \6886 , \6887 );
and \U$6757 ( \6889 , \6747 , \6751 );
and \U$6758 ( \6890 , \6751 , \6756 );
and \U$6759 ( \6891 , \6747 , \6756 );
or \U$6760 ( \6892 , \6889 , \6890 , \6891 );
xor \U$6761 ( \6893 , \6888 , \6892 );
and \U$6762 ( \6894 , \6703 , \6707 );
and \U$6763 ( \6895 , \6707 , \6712 );
and \U$6764 ( \6896 , \6703 , \6712 );
or \U$6765 ( \6897 , \6894 , \6895 , \6896 );
xor \U$6766 ( \6898 , \6893 , \6897 );
and \U$6767 ( \6899 , \6762 , \6766 );
and \U$6768 ( \6900 , \6766 , \6771 );
and \U$6769 ( \6901 , \6762 , \6771 );
or \U$6770 ( \6902 , \6899 , \6900 , \6901 );
and \U$6771 ( \6903 , \6778 , \6782 );
and \U$6772 ( \6904 , \6782 , \6787 );
and \U$6773 ( \6905 , \6778 , \6787 );
or \U$6774 ( \6906 , \6903 , \6904 , \6905 );
xor \U$6775 ( \6907 , \6902 , \6906 );
and \U$6776 ( \6908 , \6793 , \6797 );
and \U$6777 ( \6909 , \6797 , \6680 );
and \U$6778 ( \6910 , \6793 , \6680 );
or \U$6779 ( \6911 , \6908 , \6909 , \6910 );
xor \U$6780 ( \6912 , \6907 , \6911 );
xor \U$6781 ( \6913 , \6898 , \6912 );
and \U$6782 ( \6914 , \6689 , \6693 );
and \U$6783 ( \6915 , \6693 , \6698 );
and \U$6784 ( \6916 , \6689 , \6698 );
or \U$6785 ( \6917 , \6914 , \6915 , \6916 );
and \U$6786 ( \6918 , \6668 , \6672 );
and \U$6787 ( \6919 , \6672 , \6681 );
and \U$6788 ( \6920 , \6668 , \6681 );
or \U$6789 ( \6921 , \6918 , \6919 , \6920 );
xor \U$6790 ( \6922 , \6917 , \6921 );
and \U$6791 ( \6923 , \6718 , \6722 );
and \U$6792 ( \6924 , \6722 , \6727 );
and \U$6793 ( \6925 , \6718 , \6727 );
or \U$6794 ( \6926 , \6923 , \6924 , \6925 );
xor \U$6795 ( \6927 , \6922 , \6926 );
xor \U$6796 ( \6928 , \6913 , \6927 );
xor \U$6797 ( \6929 , \6884 , \6928 );
and \U$6798 ( \6930 , \3912 , \156 );
and \U$6799 ( \6931 , \4160 , \154 );
nor \U$6800 ( \6932 , \6930 , \6931 );
xnor \U$6801 ( \6933 , \6932 , \163 );
and \U$6802 ( \6934 , \3646 , \296 );
and \U$6803 ( \6935 , \3736 , \168 );
nor \U$6804 ( \6936 , \6934 , \6935 );
xnor \U$6805 ( \6937 , \6936 , \173 );
xor \U$6806 ( \6938 , \6933 , \6937 );
and \U$6807 ( \6939 , \3143 , \438 );
and \U$6808 ( \6940 , \3395 , \336 );
nor \U$6809 ( \6941 , \6939 , \6940 );
xnor \U$6810 ( \6942 , \6941 , \320 );
xor \U$6811 ( \6943 , \6938 , \6942 );
and \U$6812 ( \6944 , \6790 , \183 );
buf \U$6813 ( \6945 , RIb55ec20_77);
and \U$6814 ( \6946 , \6945 , \180 );
nor \U$6815 ( \6947 , \6944 , \6946 );
xnor \U$6816 ( \6948 , \6947 , \179 );
and \U$6817 ( \6949 , \6281 , \195 );
and \U$6818 ( \6950 , \6514 , \193 );
nor \U$6819 ( \6951 , \6949 , \6950 );
xnor \U$6820 ( \6952 , \6951 , \202 );
xor \U$6821 ( \6953 , \6948 , \6952 );
and \U$6822 ( \6954 , \5674 , \215 );
and \U$6823 ( \6955 , \6030 , \213 );
nor \U$6824 ( \6956 , \6954 , \6955 );
xnor \U$6825 ( \6957 , \6956 , \222 );
xor \U$6826 ( \6958 , \6953 , \6957 );
xor \U$6827 ( \6959 , \6943 , \6958 );
and \U$6828 ( \6960 , \5156 , \230 );
and \U$6829 ( \6961 , \5469 , \228 );
nor \U$6830 ( \6962 , \6960 , \6961 );
xnor \U$6831 ( \6963 , \6962 , \237 );
and \U$6832 ( \6964 , \4749 , \245 );
and \U$6833 ( \6965 , \4922 , \243 );
nor \U$6834 ( \6966 , \6964 , \6965 );
xnor \U$6835 ( \6967 , \6966 , \252 );
xor \U$6836 ( \6968 , \6963 , \6967 );
and \U$6837 ( \6969 , \4364 , \141 );
and \U$6838 ( \6970 , \4654 , \139 );
nor \U$6839 ( \6971 , \6969 , \6970 );
xnor \U$6840 ( \6972 , \6971 , \148 );
xor \U$6841 ( \6973 , \6968 , \6972 );
xor \U$6842 ( \6974 , \6959 , \6973 );
and \U$6843 ( \6975 , \1948 , \1824 );
and \U$6844 ( \6976 , \2090 , \1739 );
nor \U$6845 ( \6977 , \6975 , \6976 );
xnor \U$6846 ( \6978 , \6977 , \1697 );
and \U$6847 ( \6979 , \1684 , \2121 );
and \U$6848 ( \6980 , \1802 , \2008 );
nor \U$6849 ( \6981 , \6979 , \6980 );
xnor \U$6850 ( \6982 , \6981 , \1961 );
xor \U$6851 ( \6983 , \6978 , \6982 );
and \U$6852 ( \6984 , \1484 , \2400 );
and \U$6853 ( \6985 , \1601 , \2246 );
nor \U$6854 ( \6986 , \6984 , \6985 );
xnor \U$6855 ( \6987 , \6986 , \2195 );
xor \U$6856 ( \6988 , \6983 , \6987 );
and \U$6857 ( \6989 , \2826 , \1086 );
and \U$6858 ( \6990 , \3037 , \508 );
nor \U$6859 ( \6991 , \6989 , \6990 );
xnor \U$6860 ( \6992 , \6991 , \487 );
and \U$6861 ( \6993 , \2521 , \1301 );
and \U$6862 ( \6994 , \2757 , \1246 );
nor \U$6863 ( \6995 , \6993 , \6994 );
xnor \U$6864 ( \6996 , \6995 , \1205 );
xor \U$6865 ( \6997 , \6992 , \6996 );
and \U$6866 ( \6998 , \2182 , \1578 );
and \U$6867 ( \6999 , \2366 , \1431 );
nor \U$6868 ( \7000 , \6998 , \6999 );
xnor \U$6869 ( \7001 , \7000 , \1436 );
xor \U$6870 ( \7002 , \6997 , \7001 );
xor \U$6871 ( \7003 , \6988 , \7002 );
and \U$6872 ( \7004 , \1192 , \2669 );
and \U$6873 ( \7005 , \1333 , \2538 );
nor \U$6874 ( \7006 , \7004 , \7005 );
xnor \U$6875 ( \7007 , \7006 , \2534 );
and \U$6876 ( \7008 , \474 , \3103 );
and \U$6877 ( \7009 , \1147 , \2934 );
nor \U$6878 ( \7010 , \7008 , \7009 );
xnor \U$6879 ( \7011 , \7010 , \2839 );
xor \U$6880 ( \7012 , \7007 , \7011 );
and \U$6881 ( \7013 , \307 , \3357 );
and \U$6882 ( \7014 , \412 , \3255 );
nor \U$6883 ( \7015 , \7013 , \7014 );
xnor \U$6884 ( \7016 , \7015 , \3156 );
xor \U$6885 ( \7017 , \7012 , \7016 );
xor \U$6886 ( \7018 , \7003 , \7017 );
xor \U$6887 ( \7019 , \6974 , \7018 );
and \U$6888 ( \7020 , \232 , \5011 );
and \U$6889 ( \7021 , \209 , \4878 );
nor \U$6890 ( \7022 , \7020 , \7021 );
xnor \U$6891 ( \7023 , \7022 , \4762 );
and \U$6892 ( \7024 , \247 , \5485 );
and \U$6893 ( \7025 , \224 , \5275 );
nor \U$6894 ( \7026 , \7024 , \7025 );
xnor \U$6895 ( \7027 , \7026 , \5169 );
xor \U$6896 ( \7028 , \7023 , \7027 );
and \U$6897 ( \7029 , \143 , \5996 );
and \U$6898 ( \7030 , \240 , \5695 );
nor \U$6899 ( \7031 , \7029 , \7030 );
xnor \U$6900 ( \7032 , \7031 , \5687 );
xor \U$6901 ( \7033 , \7028 , \7032 );
and \U$6902 ( \7034 , \185 , \3813 );
and \U$6903 ( \7035 , \261 , \3557 );
nor \U$6904 ( \7036 , \7034 , \7035 );
xnor \U$6905 ( \7037 , \7036 , \3562 );
and \U$6906 ( \7038 , \197 , \4132 );
and \U$6907 ( \7039 , \178 , \4012 );
nor \U$6908 ( \7040 , \7038 , \7039 );
xnor \U$6909 ( \7041 , \7040 , \3925 );
xor \U$6910 ( \7042 , \7037 , \7041 );
and \U$6911 ( \7043 , \217 , \4581 );
and \U$6912 ( \7044 , \189 , \4424 );
nor \U$6913 ( \7045 , \7043 , \7044 );
xnor \U$6914 ( \7046 , \7045 , \4377 );
xor \U$6915 ( \7047 , \7042 , \7046 );
xor \U$6916 ( \7048 , \7033 , \7047 );
and \U$6917 ( \7049 , \158 , \6401 );
and \U$6918 ( \7050 , \134 , \6143 );
nor \U$6919 ( \7051 , \7049 , \7050 );
xnor \U$6920 ( \7052 , \7051 , \6148 );
xor \U$6921 ( \7053 , \6677 , \6674 );
not \U$6922 ( \7054 , \6675 );
and \U$6923 ( \7055 , \7053 , \7054 );
and \U$6924 ( \7056 , \166 , \7055 );
and \U$6925 ( \7057 , \150 , \6675 );
nor \U$6926 ( \7058 , \7056 , \7057 );
xnor \U$6927 ( \7059 , \7058 , \6680 );
xor \U$6928 ( \7060 , \7052 , \7059 );
xor \U$6929 ( \7061 , \7048 , \7060 );
xor \U$6930 ( \7062 , \7019 , \7061 );
xor \U$6931 ( \7063 , \6929 , \7062 );
xor \U$6932 ( \7064 , \6880 , \7063 );
xor \U$6933 ( \7065 , \6851 , \7064 );
xor \U$6934 ( \7066 , \6842 , \7065 );
and \U$6935 ( \7067 , \6562 , \6583 );
and \U$6936 ( \7068 , \6583 , \6804 );
and \U$6937 ( \7069 , \6562 , \6804 );
or \U$6938 ( \7070 , \7067 , \7068 , \7069 );
xor \U$6939 ( \7071 , \7066 , \7070 );
and \U$6940 ( \7072 , \6805 , \6809 );
and \U$6941 ( \7073 , \6810 , \6813 );
or \U$6942 ( \7074 , \7072 , \7073 );
xor \U$6943 ( \7075 , \7071 , \7074 );
buf \U$6944 ( \7076 , \7075 );
buf \U$6945 ( \7077 , \7076 );
and \U$6946 ( \7078 , \6846 , \6850 );
and \U$6947 ( \7079 , \6850 , \7064 );
and \U$6948 ( \7080 , \6846 , \7064 );
or \U$6949 ( \7081 , \7078 , \7079 , \7080 );
and \U$6950 ( \7082 , \6824 , \6828 );
and \U$6951 ( \7083 , \6828 , \6840 );
and \U$6952 ( \7084 , \6824 , \6840 );
or \U$6953 ( \7085 , \7082 , \7083 , \7084 );
and \U$6954 ( \7086 , \6865 , \6879 );
and \U$6955 ( \7087 , \6879 , \7063 );
and \U$6956 ( \7088 , \6865 , \7063 );
or \U$6957 ( \7089 , \7086 , \7087 , \7088 );
xor \U$6958 ( \7090 , \7085 , \7089 );
and \U$6959 ( \7091 , \6898 , \6912 );
and \U$6960 ( \7092 , \6912 , \6927 );
and \U$6961 ( \7093 , \6898 , \6927 );
or \U$6962 ( \7094 , \7091 , \7092 , \7093 );
and \U$6963 ( \7095 , \6933 , \6937 );
and \U$6964 ( \7096 , \6937 , \6942 );
and \U$6965 ( \7097 , \6933 , \6942 );
or \U$6966 ( \7098 , \7095 , \7096 , \7097 );
and \U$6967 ( \7099 , \6948 , \6952 );
and \U$6968 ( \7100 , \6952 , \6957 );
and \U$6969 ( \7101 , \6948 , \6957 );
or \U$6970 ( \7102 , \7099 , \7100 , \7101 );
xor \U$6971 ( \7103 , \7098 , \7102 );
and \U$6972 ( \7104 , \6963 , \6967 );
and \U$6973 ( \7105 , \6967 , \6972 );
and \U$6974 ( \7106 , \6963 , \6972 );
or \U$6975 ( \7107 , \7104 , \7105 , \7106 );
xor \U$6976 ( \7108 , \7103 , \7107 );
xor \U$6977 ( \7109 , \7094 , \7108 );
and \U$6978 ( \7110 , \6978 , \6982 );
and \U$6979 ( \7111 , \6982 , \6987 );
and \U$6980 ( \7112 , \6978 , \6987 );
or \U$6981 ( \7113 , \7110 , \7111 , \7112 );
and \U$6982 ( \7114 , \6992 , \6996 );
and \U$6983 ( \7115 , \6996 , \7001 );
and \U$6984 ( \7116 , \6992 , \7001 );
or \U$6985 ( \7117 , \7114 , \7115 , \7116 );
xor \U$6986 ( \7118 , \7113 , \7117 );
and \U$6987 ( \7119 , \7007 , \7011 );
and \U$6988 ( \7120 , \7011 , \7016 );
and \U$6989 ( \7121 , \7007 , \7016 );
or \U$6990 ( \7122 , \7119 , \7120 , \7121 );
xor \U$6991 ( \7123 , \7118 , \7122 );
and \U$6992 ( \7124 , \7023 , \7027 );
and \U$6993 ( \7125 , \7027 , \7032 );
and \U$6994 ( \7126 , \7023 , \7032 );
or \U$6995 ( \7127 , \7124 , \7125 , \7126 );
and \U$6996 ( \7128 , \7037 , \7041 );
and \U$6997 ( \7129 , \7041 , \7046 );
and \U$6998 ( \7130 , \7037 , \7046 );
or \U$6999 ( \7131 , \7128 , \7129 , \7130 );
xor \U$7000 ( \7132 , \7127 , \7131 );
and \U$7001 ( \7133 , \7052 , \7059 );
xor \U$7002 ( \7134 , \7132 , \7133 );
xor \U$7003 ( \7135 , \7123 , \7134 );
buf \U$7004 ( \7136 , RIb560a98_12);
xor \U$7005 ( \7137 , \7136 , \6677 );
nand \U$7006 ( \7138 , \166 , \7137 );
buf \U$7007 ( \7139 , RIb560b10_11);
and \U$7008 ( \7140 , \7136 , \6677 );
not \U$7009 ( \7141 , \7140 );
and \U$7010 ( \7142 , \7139 , \7141 );
xnor \U$7011 ( \7143 , \7138 , \7142 );
and \U$7012 ( \7144 , \240 , \5996 );
and \U$7013 ( \7145 , \247 , \5695 );
nor \U$7014 ( \7146 , \7144 , \7145 );
xnor \U$7015 ( \7147 , \7146 , \5687 );
and \U$7016 ( \7148 , \134 , \6401 );
and \U$7017 ( \7149 , \143 , \6143 );
nor \U$7018 ( \7150 , \7148 , \7149 );
xnor \U$7019 ( \7151 , \7150 , \6148 );
xor \U$7020 ( \7152 , \7147 , \7151 );
and \U$7021 ( \7153 , \150 , \7055 );
and \U$7022 ( \7154 , \158 , \6675 );
nor \U$7023 ( \7155 , \7153 , \7154 );
xnor \U$7024 ( \7156 , \7155 , \6680 );
xor \U$7025 ( \7157 , \7152 , \7156 );
xor \U$7026 ( \7158 , \7143 , \7157 );
and \U$7027 ( \7159 , \189 , \4581 );
and \U$7028 ( \7160 , \197 , \4424 );
nor \U$7029 ( \7161 , \7159 , \7160 );
xnor \U$7030 ( \7162 , \7161 , \4377 );
and \U$7031 ( \7163 , \209 , \5011 );
and \U$7032 ( \7164 , \217 , \4878 );
nor \U$7033 ( \7165 , \7163 , \7164 );
xnor \U$7034 ( \7166 , \7165 , \4762 );
xor \U$7035 ( \7167 , \7162 , \7166 );
and \U$7036 ( \7168 , \224 , \5485 );
and \U$7037 ( \7169 , \232 , \5275 );
nor \U$7038 ( \7170 , \7168 , \7169 );
xnor \U$7039 ( \7171 , \7170 , \5169 );
xor \U$7040 ( \7172 , \7167 , \7171 );
xor \U$7041 ( \7173 , \7158 , \7172 );
xor \U$7042 ( \7174 , \7135 , \7173 );
xor \U$7043 ( \7175 , \7109 , \7174 );
xor \U$7044 ( \7176 , \7090 , \7175 );
xor \U$7045 ( \7177 , \7081 , \7176 );
and \U$7046 ( \7178 , \6855 , \6859 );
and \U$7047 ( \7179 , \6859 , \6864 );
and \U$7048 ( \7180 , \6855 , \6864 );
or \U$7049 ( \7181 , \7178 , \7179 , \7180 );
and \U$7050 ( \7182 , \6833 , \6837 );
and \U$7051 ( \7183 , \6837 , \6839 );
and \U$7052 ( \7184 , \6833 , \6839 );
or \U$7053 ( \7185 , \7182 , \7183 , \7184 );
xor \U$7054 ( \7186 , \7181 , \7185 );
and \U$7055 ( \7187 , \6974 , \7018 );
and \U$7056 ( \7188 , \7018 , \7061 );
and \U$7057 ( \7189 , \6974 , \7061 );
or \U$7058 ( \7190 , \7187 , \7188 , \7189 );
xor \U$7059 ( \7191 , \7186 , \7190 );
and \U$7060 ( \7192 , \6869 , \6873 );
and \U$7061 ( \7193 , \6873 , \6878 );
and \U$7062 ( \7194 , \6869 , \6878 );
or \U$7063 ( \7195 , \7192 , \7193 , \7194 );
and \U$7064 ( \7196 , \6884 , \6928 );
and \U$7065 ( \7197 , \6928 , \7062 );
and \U$7066 ( \7198 , \6884 , \7062 );
or \U$7067 ( \7199 , \7196 , \7197 , \7198 );
xor \U$7068 ( \7200 , \7195 , \7199 );
and \U$7069 ( \7201 , \6888 , \6892 );
and \U$7070 ( \7202 , \6892 , \6897 );
and \U$7071 ( \7203 , \6888 , \6897 );
or \U$7072 ( \7204 , \7201 , \7202 , \7203 );
and \U$7073 ( \7205 , \6902 , \6906 );
and \U$7074 ( \7206 , \6906 , \6911 );
and \U$7075 ( \7207 , \6902 , \6911 );
or \U$7076 ( \7208 , \7205 , \7206 , \7207 );
xor \U$7077 ( \7209 , \7204 , \7208 );
and \U$7078 ( \7210 , \6917 , \6921 );
and \U$7079 ( \7211 , \6921 , \6926 );
and \U$7080 ( \7212 , \6917 , \6926 );
or \U$7081 ( \7213 , \7210 , \7211 , \7212 );
xor \U$7082 ( \7214 , \7209 , \7213 );
and \U$7083 ( \7215 , \6943 , \6958 );
and \U$7084 ( \7216 , \6958 , \6973 );
and \U$7085 ( \7217 , \6943 , \6973 );
or \U$7086 ( \7218 , \7215 , \7216 , \7217 );
and \U$7087 ( \7219 , \6988 , \7002 );
and \U$7088 ( \7220 , \7002 , \7017 );
and \U$7089 ( \7221 , \6988 , \7017 );
or \U$7090 ( \7222 , \7219 , \7220 , \7221 );
xor \U$7091 ( \7223 , \7218 , \7222 );
and \U$7092 ( \7224 , \7033 , \7047 );
and \U$7093 ( \7225 , \7047 , \7060 );
and \U$7094 ( \7226 , \7033 , \7060 );
or \U$7095 ( \7227 , \7224 , \7225 , \7226 );
xor \U$7096 ( \7228 , \7223 , \7227 );
xor \U$7097 ( \7229 , \7214 , \7228 );
and \U$7098 ( \7230 , \6945 , \183 );
buf \U$7099 ( \7231 , RIb55ec98_76);
and \U$7100 ( \7232 , \7231 , \180 );
nor \U$7101 ( \7233 , \7230 , \7232 );
xnor \U$7102 ( \7234 , \7233 , \179 );
and \U$7103 ( \7235 , \6514 , \195 );
and \U$7104 ( \7236 , \6790 , \193 );
nor \U$7105 ( \7237 , \7235 , \7236 );
xnor \U$7106 ( \7238 , \7237 , \202 );
xor \U$7107 ( \7239 , \7234 , \7238 );
xor \U$7108 ( \7240 , \7239 , \7142 );
and \U$7109 ( \7241 , \6030 , \215 );
and \U$7110 ( \7242 , \6281 , \213 );
nor \U$7111 ( \7243 , \7241 , \7242 );
xnor \U$7112 ( \7244 , \7243 , \222 );
and \U$7113 ( \7245 , \5469 , \230 );
and \U$7114 ( \7246 , \5674 , \228 );
nor \U$7115 ( \7247 , \7245 , \7246 );
xnor \U$7116 ( \7248 , \7247 , \237 );
xor \U$7117 ( \7249 , \7244 , \7248 );
and \U$7118 ( \7250 , \4922 , \245 );
and \U$7119 ( \7251 , \5156 , \243 );
nor \U$7120 ( \7252 , \7250 , \7251 );
xnor \U$7121 ( \7253 , \7252 , \252 );
xor \U$7122 ( \7254 , \7249 , \7253 );
and \U$7123 ( \7255 , \4654 , \141 );
and \U$7124 ( \7256 , \4749 , \139 );
nor \U$7125 ( \7257 , \7255 , \7256 );
xnor \U$7126 ( \7258 , \7257 , \148 );
and \U$7127 ( \7259 , \4160 , \156 );
and \U$7128 ( \7260 , \4364 , \154 );
nor \U$7129 ( \7261 , \7259 , \7260 );
xnor \U$7130 ( \7262 , \7261 , \163 );
xor \U$7131 ( \7263 , \7258 , \7262 );
and \U$7132 ( \7264 , \3736 , \296 );
and \U$7133 ( \7265 , \3912 , \168 );
nor \U$7134 ( \7266 , \7264 , \7265 );
xnor \U$7135 ( \7267 , \7266 , \173 );
xor \U$7136 ( \7268 , \7263 , \7267 );
xor \U$7137 ( \7269 , \7254 , \7268 );
and \U$7138 ( \7270 , \3395 , \438 );
and \U$7139 ( \7271 , \3646 , \336 );
nor \U$7140 ( \7272 , \7270 , \7271 );
xnor \U$7141 ( \7273 , \7272 , \320 );
and \U$7142 ( \7274 , \3037 , \1086 );
and \U$7143 ( \7275 , \3143 , \508 );
nor \U$7144 ( \7276 , \7274 , \7275 );
xnor \U$7145 ( \7277 , \7276 , \487 );
xor \U$7146 ( \7278 , \7273 , \7277 );
and \U$7147 ( \7279 , \2757 , \1301 );
and \U$7148 ( \7280 , \2826 , \1246 );
nor \U$7149 ( \7281 , \7279 , \7280 );
xnor \U$7150 ( \7282 , \7281 , \1205 );
xor \U$7151 ( \7283 , \7278 , \7282 );
xor \U$7152 ( \7284 , \7269 , \7283 );
xor \U$7153 ( \7285 , \7240 , \7284 );
and \U$7154 ( \7286 , \412 , \3357 );
and \U$7155 ( \7287 , \474 , \3255 );
nor \U$7156 ( \7288 , \7286 , \7287 );
xnor \U$7157 ( \7289 , \7288 , \3156 );
and \U$7158 ( \7290 , \261 , \3813 );
and \U$7159 ( \7291 , \307 , \3557 );
nor \U$7160 ( \7292 , \7290 , \7291 );
xnor \U$7161 ( \7293 , \7292 , \3562 );
xor \U$7162 ( \7294 , \7289 , \7293 );
and \U$7163 ( \7295 , \178 , \4132 );
and \U$7164 ( \7296 , \185 , \4012 );
nor \U$7165 ( \7297 , \7295 , \7296 );
xnor \U$7166 ( \7298 , \7297 , \3925 );
xor \U$7167 ( \7299 , \7294 , \7298 );
and \U$7168 ( \7300 , \1601 , \2400 );
and \U$7169 ( \7301 , \1684 , \2246 );
nor \U$7170 ( \7302 , \7300 , \7301 );
xnor \U$7171 ( \7303 , \7302 , \2195 );
and \U$7172 ( \7304 , \1333 , \2669 );
and \U$7173 ( \7305 , \1484 , \2538 );
nor \U$7174 ( \7306 , \7304 , \7305 );
xnor \U$7175 ( \7307 , \7306 , \2534 );
xor \U$7176 ( \7308 , \7303 , \7307 );
and \U$7177 ( \7309 , \1147 , \3103 );
and \U$7178 ( \7310 , \1192 , \2934 );
nor \U$7179 ( \7311 , \7309 , \7310 );
xnor \U$7180 ( \7312 , \7311 , \2839 );
xor \U$7181 ( \7313 , \7308 , \7312 );
xor \U$7182 ( \7314 , \7299 , \7313 );
and \U$7183 ( \7315 , \2366 , \1578 );
and \U$7184 ( \7316 , \2521 , \1431 );
nor \U$7185 ( \7317 , \7315 , \7316 );
xnor \U$7186 ( \7318 , \7317 , \1436 );
and \U$7187 ( \7319 , \2090 , \1824 );
and \U$7188 ( \7320 , \2182 , \1739 );
nor \U$7189 ( \7321 , \7319 , \7320 );
xnor \U$7190 ( \7322 , \7321 , \1697 );
xor \U$7191 ( \7323 , \7318 , \7322 );
and \U$7192 ( \7324 , \1802 , \2121 );
and \U$7193 ( \7325 , \1948 , \2008 );
nor \U$7194 ( \7326 , \7324 , \7325 );
xnor \U$7195 ( \7327 , \7326 , \1961 );
xor \U$7196 ( \7328 , \7323 , \7327 );
xor \U$7197 ( \7329 , \7314 , \7328 );
xor \U$7198 ( \7330 , \7285 , \7329 );
xor \U$7199 ( \7331 , \7229 , \7330 );
xor \U$7200 ( \7332 , \7200 , \7331 );
xor \U$7201 ( \7333 , \7191 , \7332 );
xor \U$7202 ( \7334 , \7177 , \7333 );
and \U$7203 ( \7335 , \6820 , \6841 );
and \U$7204 ( \7336 , \6841 , \7065 );
and \U$7205 ( \7337 , \6820 , \7065 );
or \U$7206 ( \7338 , \7335 , \7336 , \7337 );
xor \U$7207 ( \7339 , \7334 , \7338 );
and \U$7208 ( \7340 , \7066 , \7070 );
and \U$7209 ( \7341 , \7071 , \7074 );
or \U$7210 ( \7342 , \7340 , \7341 );
xor \U$7211 ( \7343 , \7339 , \7342 );
buf \U$7212 ( \7344 , \7343 );
buf \U$7213 ( \7345 , \7344 );
and \U$7214 ( \7346 , \7085 , \7089 );
and \U$7215 ( \7347 , \7089 , \7175 );
and \U$7216 ( \7348 , \7085 , \7175 );
or \U$7217 ( \7349 , \7346 , \7347 , \7348 );
and \U$7218 ( \7350 , \7191 , \7332 );
xor \U$7219 ( \7351 , \7349 , \7350 );
and \U$7220 ( \7352 , \7195 , \7199 );
and \U$7221 ( \7353 , \7199 , \7331 );
and \U$7222 ( \7354 , \7195 , \7331 );
or \U$7223 ( \7355 , \7352 , \7353 , \7354 );
and \U$7224 ( \7356 , \7181 , \7185 );
and \U$7225 ( \7357 , \7185 , \7190 );
and \U$7226 ( \7358 , \7181 , \7190 );
or \U$7227 ( \7359 , \7356 , \7357 , \7358 );
and \U$7228 ( \7360 , \7094 , \7108 );
and \U$7229 ( \7361 , \7108 , \7174 );
and \U$7230 ( \7362 , \7094 , \7174 );
or \U$7231 ( \7363 , \7360 , \7361 , \7362 );
xor \U$7232 ( \7364 , \7359 , \7363 );
and \U$7233 ( \7365 , \7214 , \7228 );
and \U$7234 ( \7366 , \7228 , \7330 );
and \U$7235 ( \7367 , \7214 , \7330 );
or \U$7236 ( \7368 , \7365 , \7366 , \7367 );
xor \U$7237 ( \7369 , \7364 , \7368 );
xor \U$7238 ( \7370 , \7355 , \7369 );
and \U$7239 ( \7371 , \7204 , \7208 );
and \U$7240 ( \7372 , \7208 , \7213 );
and \U$7241 ( \7373 , \7204 , \7213 );
or \U$7242 ( \7374 , \7371 , \7372 , \7373 );
and \U$7243 ( \7375 , \7218 , \7222 );
and \U$7244 ( \7376 , \7222 , \7227 );
and \U$7245 ( \7377 , \7218 , \7227 );
or \U$7246 ( \7378 , \7375 , \7376 , \7377 );
xor \U$7247 ( \7379 , \7374 , \7378 );
and \U$7248 ( \7380 , \7240 , \7284 );
and \U$7249 ( \7381 , \7284 , \7329 );
and \U$7250 ( \7382 , \7240 , \7329 );
or \U$7251 ( \7383 , \7380 , \7381 , \7382 );
xor \U$7252 ( \7384 , \7379 , \7383 );
and \U$7253 ( \7385 , \7123 , \7134 );
and \U$7254 ( \7386 , \7134 , \7173 );
and \U$7255 ( \7387 , \7123 , \7173 );
or \U$7256 ( \7388 , \7385 , \7386 , \7387 );
and \U$7257 ( \7389 , \7303 , \7307 );
and \U$7258 ( \7390 , \7307 , \7312 );
and \U$7259 ( \7391 , \7303 , \7312 );
or \U$7260 ( \7392 , \7389 , \7390 , \7391 );
and \U$7261 ( \7393 , \7273 , \7277 );
and \U$7262 ( \7394 , \7277 , \7282 );
and \U$7263 ( \7395 , \7273 , \7282 );
or \U$7264 ( \7396 , \7393 , \7394 , \7395 );
xor \U$7265 ( \7397 , \7392 , \7396 );
and \U$7266 ( \7398 , \7318 , \7322 );
and \U$7267 ( \7399 , \7322 , \7327 );
and \U$7268 ( \7400 , \7318 , \7327 );
or \U$7269 ( \7401 , \7398 , \7399 , \7400 );
xor \U$7270 ( \7402 , \7397 , \7401 );
and \U$7271 ( \7403 , \7244 , \7248 );
and \U$7272 ( \7404 , \7248 , \7253 );
and \U$7273 ( \7405 , \7244 , \7253 );
or \U$7274 ( \7406 , \7403 , \7404 , \7405 );
and \U$7275 ( \7407 , \7234 , \7238 );
and \U$7276 ( \7408 , \7238 , \7142 );
and \U$7277 ( \7409 , \7234 , \7142 );
or \U$7278 ( \7410 , \7407 , \7408 , \7409 );
xor \U$7279 ( \7411 , \7406 , \7410 );
and \U$7280 ( \7412 , \7258 , \7262 );
and \U$7281 ( \7413 , \7262 , \7267 );
and \U$7282 ( \7414 , \7258 , \7267 );
or \U$7283 ( \7415 , \7412 , \7413 , \7414 );
xor \U$7284 ( \7416 , \7411 , \7415 );
xor \U$7285 ( \7417 , \7402 , \7416 );
and \U$7286 ( \7418 , \7147 , \7151 );
and \U$7287 ( \7419 , \7151 , \7156 );
and \U$7288 ( \7420 , \7147 , \7156 );
or \U$7289 ( \7421 , \7418 , \7419 , \7420 );
and \U$7290 ( \7422 , \7289 , \7293 );
and \U$7291 ( \7423 , \7293 , \7298 );
and \U$7292 ( \7424 , \7289 , \7298 );
or \U$7293 ( \7425 , \7422 , \7423 , \7424 );
xor \U$7294 ( \7426 , \7421 , \7425 );
and \U$7295 ( \7427 , \7162 , \7166 );
and \U$7296 ( \7428 , \7166 , \7171 );
and \U$7297 ( \7429 , \7162 , \7171 );
or \U$7298 ( \7430 , \7427 , \7428 , \7429 );
xor \U$7299 ( \7431 , \7426 , \7430 );
xor \U$7300 ( \7432 , \7417 , \7431 );
xor \U$7301 ( \7433 , \7388 , \7432 );
and \U$7302 ( \7434 , \1484 , \2669 );
and \U$7303 ( \7435 , \1601 , \2538 );
nor \U$7304 ( \7436 , \7434 , \7435 );
xnor \U$7305 ( \7437 , \7436 , \2534 );
and \U$7306 ( \7438 , \1192 , \3103 );
and \U$7307 ( \7439 , \1333 , \2934 );
nor \U$7308 ( \7440 , \7438 , \7439 );
xnor \U$7309 ( \7441 , \7440 , \2839 );
xor \U$7310 ( \7442 , \7437 , \7441 );
and \U$7311 ( \7443 , \474 , \3357 );
and \U$7312 ( \7444 , \1147 , \3255 );
nor \U$7313 ( \7445 , \7443 , \7444 );
xnor \U$7314 ( \7446 , \7445 , \3156 );
xor \U$7315 ( \7447 , \7442 , \7446 );
and \U$7316 ( \7448 , \2182 , \1824 );
and \U$7317 ( \7449 , \2366 , \1739 );
nor \U$7318 ( \7450 , \7448 , \7449 );
xnor \U$7319 ( \7451 , \7450 , \1697 );
and \U$7320 ( \7452 , \1948 , \2121 );
and \U$7321 ( \7453 , \2090 , \2008 );
nor \U$7322 ( \7454 , \7452 , \7453 );
xnor \U$7323 ( \7455 , \7454 , \1961 );
xor \U$7324 ( \7456 , \7451 , \7455 );
and \U$7325 ( \7457 , \1684 , \2400 );
and \U$7326 ( \7458 , \1802 , \2246 );
nor \U$7327 ( \7459 , \7457 , \7458 );
xnor \U$7328 ( \7460 , \7459 , \2195 );
xor \U$7329 ( \7461 , \7456 , \7460 );
xor \U$7330 ( \7462 , \7447 , \7461 );
and \U$7331 ( \7463 , \3143 , \1086 );
and \U$7332 ( \7464 , \3395 , \508 );
nor \U$7333 ( \7465 , \7463 , \7464 );
xnor \U$7334 ( \7466 , \7465 , \487 );
and \U$7335 ( \7467 , \2826 , \1301 );
and \U$7336 ( \7468 , \3037 , \1246 );
nor \U$7337 ( \7469 , \7467 , \7468 );
xnor \U$7338 ( \7470 , \7469 , \1205 );
xor \U$7339 ( \7471 , \7466 , \7470 );
and \U$7340 ( \7472 , \2521 , \1578 );
and \U$7341 ( \7473 , \2757 , \1431 );
nor \U$7342 ( \7474 , \7472 , \7473 );
xnor \U$7343 ( \7475 , \7474 , \1436 );
xor \U$7344 ( \7476 , \7471 , \7475 );
xor \U$7345 ( \7477 , \7462 , \7476 );
and \U$7346 ( \7478 , \143 , \6401 );
and \U$7347 ( \7479 , \240 , \6143 );
nor \U$7348 ( \7480 , \7478 , \7479 );
xnor \U$7349 ( \7481 , \7480 , \6148 );
and \U$7350 ( \7482 , \158 , \7055 );
and \U$7351 ( \7483 , \134 , \6675 );
nor \U$7352 ( \7484 , \7482 , \7483 );
xnor \U$7353 ( \7485 , \7484 , \6680 );
xor \U$7354 ( \7486 , \7481 , \7485 );
xor \U$7355 ( \7487 , \7139 , \7136 );
not \U$7356 ( \7488 , \7137 );
and \U$7357 ( \7489 , \7487 , \7488 );
and \U$7358 ( \7490 , \166 , \7489 );
and \U$7359 ( \7491 , \150 , \7137 );
nor \U$7360 ( \7492 , \7490 , \7491 );
xnor \U$7361 ( \7493 , \7492 , \7142 );
xor \U$7362 ( \7494 , \7486 , \7493 );
and \U$7363 ( \7495 , \307 , \3813 );
and \U$7364 ( \7496 , \412 , \3557 );
nor \U$7365 ( \7497 , \7495 , \7496 );
xnor \U$7366 ( \7498 , \7497 , \3562 );
and \U$7367 ( \7499 , \185 , \4132 );
and \U$7368 ( \7500 , \261 , \4012 );
nor \U$7369 ( \7501 , \7499 , \7500 );
xnor \U$7370 ( \7502 , \7501 , \3925 );
xor \U$7371 ( \7503 , \7498 , \7502 );
and \U$7372 ( \7504 , \197 , \4581 );
and \U$7373 ( \7505 , \178 , \4424 );
nor \U$7374 ( \7506 , \7504 , \7505 );
xnor \U$7375 ( \7507 , \7506 , \4377 );
xor \U$7376 ( \7508 , \7503 , \7507 );
xor \U$7377 ( \7509 , \7494 , \7508 );
and \U$7378 ( \7510 , \217 , \5011 );
and \U$7379 ( \7511 , \189 , \4878 );
nor \U$7380 ( \7512 , \7510 , \7511 );
xnor \U$7381 ( \7513 , \7512 , \4762 );
and \U$7382 ( \7514 , \232 , \5485 );
and \U$7383 ( \7515 , \209 , \5275 );
nor \U$7384 ( \7516 , \7514 , \7515 );
xnor \U$7385 ( \7517 , \7516 , \5169 );
xor \U$7386 ( \7518 , \7513 , \7517 );
and \U$7387 ( \7519 , \247 , \5996 );
and \U$7388 ( \7520 , \224 , \5695 );
nor \U$7389 ( \7521 , \7519 , \7520 );
xnor \U$7390 ( \7522 , \7521 , \5687 );
xor \U$7391 ( \7523 , \7518 , \7522 );
xor \U$7392 ( \7524 , \7509 , \7523 );
xor \U$7393 ( \7525 , \7477 , \7524 );
and \U$7394 ( \7526 , \5674 , \230 );
and \U$7395 ( \7527 , \6030 , \228 );
nor \U$7396 ( \7528 , \7526 , \7527 );
xnor \U$7397 ( \7529 , \7528 , \237 );
and \U$7398 ( \7530 , \5156 , \245 );
and \U$7399 ( \7531 , \5469 , \243 );
nor \U$7400 ( \7532 , \7530 , \7531 );
xnor \U$7401 ( \7533 , \7532 , \252 );
xor \U$7402 ( \7534 , \7529 , \7533 );
and \U$7403 ( \7535 , \4749 , \141 );
and \U$7404 ( \7536 , \4922 , \139 );
nor \U$7405 ( \7537 , \7535 , \7536 );
xnor \U$7406 ( \7538 , \7537 , \148 );
xor \U$7407 ( \7539 , \7534 , \7538 );
and \U$7408 ( \7540 , \4364 , \156 );
and \U$7409 ( \7541 , \4654 , \154 );
nor \U$7410 ( \7542 , \7540 , \7541 );
xnor \U$7411 ( \7543 , \7542 , \163 );
and \U$7412 ( \7544 , \3912 , \296 );
and \U$7413 ( \7545 , \4160 , \168 );
nor \U$7414 ( \7546 , \7544 , \7545 );
xnor \U$7415 ( \7547 , \7546 , \173 );
xor \U$7416 ( \7548 , \7543 , \7547 );
and \U$7417 ( \7549 , \3646 , \438 );
and \U$7418 ( \7550 , \3736 , \336 );
nor \U$7419 ( \7551 , \7549 , \7550 );
xnor \U$7420 ( \7552 , \7551 , \320 );
xor \U$7421 ( \7553 , \7548 , \7552 );
xor \U$7422 ( \7554 , \7539 , \7553 );
and \U$7423 ( \7555 , \7231 , \183 );
buf \U$7424 ( \7556 , RIb55ed10_75);
and \U$7425 ( \7557 , \7556 , \180 );
nor \U$7426 ( \7558 , \7555 , \7557 );
xnor \U$7427 ( \7559 , \7558 , \179 );
and \U$7428 ( \7560 , \6790 , \195 );
and \U$7429 ( \7561 , \6945 , \193 );
nor \U$7430 ( \7562 , \7560 , \7561 );
xnor \U$7431 ( \7563 , \7562 , \202 );
xor \U$7432 ( \7564 , \7559 , \7563 );
and \U$7433 ( \7565 , \6281 , \215 );
and \U$7434 ( \7566 , \6514 , \213 );
nor \U$7435 ( \7567 , \7565 , \7566 );
xnor \U$7436 ( \7568 , \7567 , \222 );
xor \U$7437 ( \7569 , \7564 , \7568 );
xor \U$7438 ( \7570 , \7554 , \7569 );
xor \U$7439 ( \7571 , \7525 , \7570 );
xor \U$7440 ( \7572 , \7433 , \7571 );
xor \U$7441 ( \7573 , \7384 , \7572 );
and \U$7442 ( \7574 , \7113 , \7117 );
and \U$7443 ( \7575 , \7117 , \7122 );
and \U$7444 ( \7576 , \7113 , \7122 );
or \U$7445 ( \7577 , \7574 , \7575 , \7576 );
and \U$7446 ( \7578 , \7127 , \7131 );
and \U$7447 ( \7579 , \7131 , \7133 );
and \U$7448 ( \7580 , \7127 , \7133 );
or \U$7449 ( \7581 , \7578 , \7579 , \7580 );
xor \U$7450 ( \7582 , \7577 , \7581 );
and \U$7451 ( \7583 , \7098 , \7102 );
and \U$7452 ( \7584 , \7102 , \7107 );
and \U$7453 ( \7585 , \7098 , \7107 );
or \U$7454 ( \7586 , \7583 , \7584 , \7585 );
xor \U$7455 ( \7587 , \7582 , \7586 );
and \U$7456 ( \7588 , \7254 , \7268 );
and \U$7457 ( \7589 , \7268 , \7283 );
and \U$7458 ( \7590 , \7254 , \7283 );
or \U$7459 ( \7591 , \7588 , \7589 , \7590 );
and \U$7460 ( \7592 , \7143 , \7157 );
and \U$7461 ( \7593 , \7157 , \7172 );
and \U$7462 ( \7594 , \7143 , \7172 );
or \U$7463 ( \7595 , \7592 , \7593 , \7594 );
xor \U$7464 ( \7596 , \7591 , \7595 );
and \U$7465 ( \7597 , \7299 , \7313 );
and \U$7466 ( \7598 , \7313 , \7328 );
and \U$7467 ( \7599 , \7299 , \7328 );
or \U$7468 ( \7600 , \7597 , \7598 , \7599 );
xor \U$7469 ( \7601 , \7596 , \7600 );
xor \U$7470 ( \7602 , \7587 , \7601 );
xor \U$7471 ( \7603 , \7573 , \7602 );
xor \U$7472 ( \7604 , \7370 , \7603 );
xor \U$7473 ( \7605 , \7351 , \7604 );
and \U$7474 ( \7606 , \7081 , \7176 );
and \U$7475 ( \7607 , \7176 , \7333 );
and \U$7476 ( \7608 , \7081 , \7333 );
or \U$7477 ( \7609 , \7606 , \7607 , \7608 );
xor \U$7478 ( \7610 , \7605 , \7609 );
and \U$7479 ( \7611 , \7334 , \7338 );
and \U$7480 ( \7612 , \7339 , \7342 );
or \U$7481 ( \7613 , \7611 , \7612 );
xor \U$7482 ( \7614 , \7610 , \7613 );
buf \U$7483 ( \7615 , \7614 );
buf \U$7484 ( \7616 , \7615 );
and \U$7485 ( \7617 , \7355 , \7369 );
and \U$7486 ( \7618 , \7369 , \7603 );
and \U$7487 ( \7619 , \7355 , \7603 );
or \U$7488 ( \7620 , \7617 , \7618 , \7619 );
and \U$7489 ( \7621 , \7374 , \7378 );
and \U$7490 ( \7622 , \7378 , \7383 );
and \U$7491 ( \7623 , \7374 , \7383 );
or \U$7492 ( \7624 , \7621 , \7622 , \7623 );
and \U$7493 ( \7625 , \7388 , \7432 );
and \U$7494 ( \7626 , \7432 , \7571 );
and \U$7495 ( \7627 , \7388 , \7571 );
or \U$7496 ( \7628 , \7625 , \7626 , \7627 );
xor \U$7497 ( \7629 , \7624 , \7628 );
and \U$7498 ( \7630 , \7587 , \7601 );
xor \U$7499 ( \7631 , \7629 , \7630 );
xor \U$7500 ( \7632 , \7620 , \7631 );
and \U$7501 ( \7633 , \7359 , \7363 );
and \U$7502 ( \7634 , \7363 , \7368 );
and \U$7503 ( \7635 , \7359 , \7368 );
or \U$7504 ( \7636 , \7633 , \7634 , \7635 );
and \U$7505 ( \7637 , \7384 , \7572 );
and \U$7506 ( \7638 , \7572 , \7602 );
and \U$7507 ( \7639 , \7384 , \7602 );
or \U$7508 ( \7640 , \7637 , \7638 , \7639 );
xor \U$7509 ( \7641 , \7636 , \7640 );
and \U$7510 ( \7642 , \7577 , \7581 );
and \U$7511 ( \7643 , \7581 , \7586 );
and \U$7512 ( \7644 , \7577 , \7586 );
or \U$7513 ( \7645 , \7642 , \7643 , \7644 );
and \U$7514 ( \7646 , \7591 , \7595 );
and \U$7515 ( \7647 , \7595 , \7600 );
and \U$7516 ( \7648 , \7591 , \7600 );
or \U$7517 ( \7649 , \7646 , \7647 , \7648 );
xor \U$7518 ( \7650 , \7645 , \7649 );
and \U$7519 ( \7651 , \7477 , \7524 );
and \U$7520 ( \7652 , \7524 , \7570 );
and \U$7521 ( \7653 , \7477 , \7570 );
or \U$7522 ( \7654 , \7651 , \7652 , \7653 );
xor \U$7523 ( \7655 , \7650 , \7654 );
and \U$7524 ( \7656 , \7447 , \7461 );
and \U$7525 ( \7657 , \7461 , \7476 );
and \U$7526 ( \7658 , \7447 , \7476 );
or \U$7527 ( \7659 , \7656 , \7657 , \7658 );
and \U$7528 ( \7660 , \7494 , \7508 );
and \U$7529 ( \7661 , \7508 , \7523 );
and \U$7530 ( \7662 , \7494 , \7523 );
or \U$7531 ( \7663 , \7660 , \7661 , \7662 );
xor \U$7532 ( \7664 , \7659 , \7663 );
and \U$7533 ( \7665 , \7539 , \7553 );
and \U$7534 ( \7666 , \7553 , \7569 );
and \U$7535 ( \7667 , \7539 , \7569 );
or \U$7536 ( \7668 , \7665 , \7666 , \7667 );
xor \U$7537 ( \7669 , \7664 , \7668 );
and \U$7538 ( \7670 , \7392 , \7396 );
and \U$7539 ( \7671 , \7396 , \7401 );
and \U$7540 ( \7672 , \7392 , \7401 );
or \U$7541 ( \7673 , \7670 , \7671 , \7672 );
and \U$7542 ( \7674 , \7406 , \7410 );
and \U$7543 ( \7675 , \7410 , \7415 );
and \U$7544 ( \7676 , \7406 , \7415 );
or \U$7545 ( \7677 , \7674 , \7675 , \7676 );
xor \U$7546 ( \7678 , \7673 , \7677 );
and \U$7547 ( \7679 , \7421 , \7425 );
and \U$7548 ( \7680 , \7425 , \7430 );
and \U$7549 ( \7681 , \7421 , \7430 );
or \U$7550 ( \7682 , \7679 , \7680 , \7681 );
xor \U$7551 ( \7683 , \7678 , \7682 );
xor \U$7552 ( \7684 , \7669 , \7683 );
and \U$7553 ( \7685 , \6514 , \215 );
and \U$7554 ( \7686 , \6790 , \213 );
nor \U$7555 ( \7687 , \7685 , \7686 );
xnor \U$7556 ( \7688 , \7687 , \222 );
and \U$7557 ( \7689 , \6030 , \230 );
and \U$7558 ( \7690 , \6281 , \228 );
nor \U$7559 ( \7691 , \7689 , \7690 );
xnor \U$7560 ( \7692 , \7691 , \237 );
xor \U$7561 ( \7693 , \7688 , \7692 );
and \U$7562 ( \7694 , \5469 , \245 );
and \U$7563 ( \7695 , \5674 , \243 );
nor \U$7564 ( \7696 , \7694 , \7695 );
xnor \U$7565 ( \7697 , \7696 , \252 );
xor \U$7566 ( \7698 , \7693 , \7697 );
and \U$7567 ( \7699 , \7556 , \183 );
buf \U$7568 ( \7700 , RIb55ed88_74);
and \U$7569 ( \7701 , \7700 , \180 );
nor \U$7570 ( \7702 , \7699 , \7701 );
xnor \U$7571 ( \7703 , \7702 , \179 );
and \U$7572 ( \7704 , \6945 , \195 );
and \U$7573 ( \7705 , \7231 , \193 );
nor \U$7574 ( \7706 , \7704 , \7705 );
xnor \U$7575 ( \7707 , \7706 , \202 );
xor \U$7576 ( \7708 , \7703 , \7707 );
buf \U$7577 ( \7709 , RIb560c00_9);
buf \U$7578 ( \7710 , RIb560b88_10);
and \U$7579 ( \7711 , \7710 , \7139 );
not \U$7580 ( \7712 , \7711 );
and \U$7581 ( \7713 , \7709 , \7712 );
xor \U$7582 ( \7714 , \7708 , \7713 );
xor \U$7583 ( \7715 , \7698 , \7714 );
and \U$7584 ( \7716 , \4922 , \141 );
and \U$7585 ( \7717 , \5156 , \139 );
nor \U$7586 ( \7718 , \7716 , \7717 );
xnor \U$7587 ( \7719 , \7718 , \148 );
and \U$7588 ( \7720 , \4654 , \156 );
and \U$7589 ( \7721 , \4749 , \154 );
nor \U$7590 ( \7722 , \7720 , \7721 );
xnor \U$7591 ( \7723 , \7722 , \163 );
xor \U$7592 ( \7724 , \7719 , \7723 );
and \U$7593 ( \7725 , \4160 , \296 );
and \U$7594 ( \7726 , \4364 , \168 );
nor \U$7595 ( \7727 , \7725 , \7726 );
xnor \U$7596 ( \7728 , \7727 , \173 );
xor \U$7597 ( \7729 , \7724 , \7728 );
and \U$7598 ( \7730 , \2757 , \1578 );
and \U$7599 ( \7731 , \2826 , \1431 );
nor \U$7600 ( \7732 , \7730 , \7731 );
xnor \U$7601 ( \7733 , \7732 , \1436 );
and \U$7602 ( \7734 , \2366 , \1824 );
and \U$7603 ( \7735 , \2521 , \1739 );
nor \U$7604 ( \7736 , \7734 , \7735 );
xnor \U$7605 ( \7737 , \7736 , \1697 );
xor \U$7606 ( \7738 , \7733 , \7737 );
and \U$7607 ( \7739 , \2090 , \2121 );
and \U$7608 ( \7740 , \2182 , \2008 );
nor \U$7609 ( \7741 , \7739 , \7740 );
xnor \U$7610 ( \7742 , \7741 , \1961 );
xor \U$7611 ( \7743 , \7738 , \7742 );
xor \U$7612 ( \7744 , \7729 , \7743 );
and \U$7613 ( \7745 , \3736 , \438 );
and \U$7614 ( \7746 , \3912 , \336 );
nor \U$7615 ( \7747 , \7745 , \7746 );
xnor \U$7616 ( \7748 , \7747 , \320 );
and \U$7617 ( \7749 , \3395 , \1086 );
and \U$7618 ( \7750 , \3646 , \508 );
nor \U$7619 ( \7751 , \7749 , \7750 );
xnor \U$7620 ( \7752 , \7751 , \487 );
xor \U$7621 ( \7753 , \7748 , \7752 );
and \U$7622 ( \7754 , \3037 , \1301 );
and \U$7623 ( \7755 , \3143 , \1246 );
nor \U$7624 ( \7756 , \7754 , \7755 );
xnor \U$7625 ( \7757 , \7756 , \1205 );
xor \U$7626 ( \7758 , \7753 , \7757 );
xor \U$7627 ( \7759 , \7744 , \7758 );
xor \U$7628 ( \7760 , \7715 , \7759 );
xor \U$7629 ( \7761 , \7684 , \7760 );
xor \U$7630 ( \7762 , \7655 , \7761 );
and \U$7631 ( \7763 , \7402 , \7416 );
and \U$7632 ( \7764 , \7416 , \7431 );
and \U$7633 ( \7765 , \7402 , \7431 );
or \U$7634 ( \7766 , \7763 , \7764 , \7765 );
and \U$7635 ( \7767 , \7481 , \7485 );
and \U$7636 ( \7768 , \7485 , \7493 );
and \U$7637 ( \7769 , \7481 , \7493 );
or \U$7638 ( \7770 , \7767 , \7768 , \7769 );
and \U$7639 ( \7771 , \7498 , \7502 );
and \U$7640 ( \7772 , \7502 , \7507 );
and \U$7641 ( \7773 , \7498 , \7507 );
or \U$7642 ( \7774 , \7771 , \7772 , \7773 );
xor \U$7643 ( \7775 , \7770 , \7774 );
and \U$7644 ( \7776 , \7513 , \7517 );
and \U$7645 ( \7777 , \7517 , \7522 );
and \U$7646 ( \7778 , \7513 , \7522 );
or \U$7647 ( \7779 , \7776 , \7777 , \7778 );
xor \U$7648 ( \7780 , \7775 , \7779 );
and \U$7649 ( \7781 , \1802 , \2400 );
and \U$7650 ( \7782 , \1948 , \2246 );
nor \U$7651 ( \7783 , \7781 , \7782 );
xnor \U$7652 ( \7784 , \7783 , \2195 );
and \U$7653 ( \7785 , \1601 , \2669 );
and \U$7654 ( \7786 , \1684 , \2538 );
nor \U$7655 ( \7787 , \7785 , \7786 );
xnor \U$7656 ( \7788 , \7787 , \2534 );
xor \U$7657 ( \7789 , \7784 , \7788 );
and \U$7658 ( \7790 , \1333 , \3103 );
and \U$7659 ( \7791 , \1484 , \2934 );
nor \U$7660 ( \7792 , \7790 , \7791 );
xnor \U$7661 ( \7793 , \7792 , \2839 );
xor \U$7662 ( \7794 , \7789 , \7793 );
and \U$7663 ( \7795 , \1147 , \3357 );
and \U$7664 ( \7796 , \1192 , \3255 );
nor \U$7665 ( \7797 , \7795 , \7796 );
xnor \U$7666 ( \7798 , \7797 , \3156 );
and \U$7667 ( \7799 , \412 , \3813 );
and \U$7668 ( \7800 , \474 , \3557 );
nor \U$7669 ( \7801 , \7799 , \7800 );
xnor \U$7670 ( \7802 , \7801 , \3562 );
xor \U$7671 ( \7803 , \7798 , \7802 );
and \U$7672 ( \7804 , \261 , \4132 );
and \U$7673 ( \7805 , \307 , \4012 );
nor \U$7674 ( \7806 , \7804 , \7805 );
xnor \U$7675 ( \7807 , \7806 , \3925 );
xor \U$7676 ( \7808 , \7803 , \7807 );
xor \U$7677 ( \7809 , \7794 , \7808 );
and \U$7678 ( \7810 , \178 , \4581 );
and \U$7679 ( \7811 , \185 , \4424 );
nor \U$7680 ( \7812 , \7810 , \7811 );
xnor \U$7681 ( \7813 , \7812 , \4377 );
and \U$7682 ( \7814 , \189 , \5011 );
and \U$7683 ( \7815 , \197 , \4878 );
nor \U$7684 ( \7816 , \7814 , \7815 );
xnor \U$7685 ( \7817 , \7816 , \4762 );
xor \U$7686 ( \7818 , \7813 , \7817 );
and \U$7687 ( \7819 , \209 , \5485 );
and \U$7688 ( \7820 , \217 , \5275 );
nor \U$7689 ( \7821 , \7819 , \7820 );
xnor \U$7690 ( \7822 , \7821 , \5169 );
xor \U$7691 ( \7823 , \7818 , \7822 );
xor \U$7692 ( \7824 , \7809 , \7823 );
xor \U$7693 ( \7825 , \7780 , \7824 );
and \U$7694 ( \7826 , \150 , \7489 );
and \U$7695 ( \7827 , \158 , \7137 );
nor \U$7696 ( \7828 , \7826 , \7827 );
xnor \U$7697 ( \7829 , \7828 , \7142 );
xor \U$7698 ( \7830 , \7710 , \7139 );
nand \U$7699 ( \7831 , \166 , \7830 );
xnor \U$7700 ( \7832 , \7831 , \7713 );
xor \U$7701 ( \7833 , \7829 , \7832 );
and \U$7702 ( \7834 , \224 , \5996 );
and \U$7703 ( \7835 , \232 , \5695 );
nor \U$7704 ( \7836 , \7834 , \7835 );
xnor \U$7705 ( \7837 , \7836 , \5687 );
and \U$7706 ( \7838 , \240 , \6401 );
and \U$7707 ( \7839 , \247 , \6143 );
nor \U$7708 ( \7840 , \7838 , \7839 );
xnor \U$7709 ( \7841 , \7840 , \6148 );
xor \U$7710 ( \7842 , \7837 , \7841 );
and \U$7711 ( \7843 , \134 , \7055 );
and \U$7712 ( \7844 , \143 , \6675 );
nor \U$7713 ( \7845 , \7843 , \7844 );
xnor \U$7714 ( \7846 , \7845 , \6680 );
xor \U$7715 ( \7847 , \7842 , \7846 );
xor \U$7716 ( \7848 , \7833 , \7847 );
xor \U$7717 ( \7849 , \7825 , \7848 );
xor \U$7718 ( \7850 , \7766 , \7849 );
and \U$7719 ( \7851 , \7529 , \7533 );
and \U$7720 ( \7852 , \7533 , \7538 );
and \U$7721 ( \7853 , \7529 , \7538 );
or \U$7722 ( \7854 , \7851 , \7852 , \7853 );
and \U$7723 ( \7855 , \7543 , \7547 );
and \U$7724 ( \7856 , \7547 , \7552 );
and \U$7725 ( \7857 , \7543 , \7552 );
or \U$7726 ( \7858 , \7855 , \7856 , \7857 );
xor \U$7727 ( \7859 , \7854 , \7858 );
and \U$7728 ( \7860 , \7559 , \7563 );
and \U$7729 ( \7861 , \7563 , \7568 );
and \U$7730 ( \7862 , \7559 , \7568 );
or \U$7731 ( \7863 , \7860 , \7861 , \7862 );
xor \U$7732 ( \7864 , \7859 , \7863 );
and \U$7733 ( \7865 , \7437 , \7441 );
and \U$7734 ( \7866 , \7441 , \7446 );
and \U$7735 ( \7867 , \7437 , \7446 );
or \U$7736 ( \7868 , \7865 , \7866 , \7867 );
and \U$7737 ( \7869 , \7451 , \7455 );
and \U$7738 ( \7870 , \7455 , \7460 );
and \U$7739 ( \7871 , \7451 , \7460 );
or \U$7740 ( \7872 , \7869 , \7870 , \7871 );
xor \U$7741 ( \7873 , \7868 , \7872 );
and \U$7742 ( \7874 , \7466 , \7470 );
and \U$7743 ( \7875 , \7470 , \7475 );
and \U$7744 ( \7876 , \7466 , \7475 );
or \U$7745 ( \7877 , \7874 , \7875 , \7876 );
xor \U$7746 ( \7878 , \7873 , \7877 );
xor \U$7747 ( \7879 , \7864 , \7878 );
xor \U$7748 ( \7880 , \7850 , \7879 );
xor \U$7749 ( \7881 , \7762 , \7880 );
xor \U$7750 ( \7882 , \7641 , \7881 );
xor \U$7751 ( \7883 , \7632 , \7882 );
and \U$7752 ( \7884 , \7349 , \7350 );
and \U$7753 ( \7885 , \7350 , \7604 );
and \U$7754 ( \7886 , \7349 , \7604 );
or \U$7755 ( \7887 , \7884 , \7885 , \7886 );
xor \U$7756 ( \7888 , \7883 , \7887 );
and \U$7757 ( \7889 , \7605 , \7609 );
and \U$7758 ( \7890 , \7610 , \7613 );
or \U$7759 ( \7891 , \7889 , \7890 );
xor \U$7760 ( \7892 , \7888 , \7891 );
buf \U$7761 ( \7893 , \7892 );
buf \U$7762 ( \7894 , \7893 );
and \U$7763 ( \7895 , \7636 , \7640 );
and \U$7764 ( \7896 , \7640 , \7881 );
and \U$7765 ( \7897 , \7636 , \7881 );
or \U$7766 ( \7898 , \7895 , \7896 , \7897 );
and \U$7767 ( \7899 , \7624 , \7628 );
and \U$7768 ( \7900 , \7628 , \7630 );
and \U$7769 ( \7901 , \7624 , \7630 );
or \U$7770 ( \7902 , \7899 , \7900 , \7901 );
and \U$7771 ( \7903 , \7655 , \7761 );
and \U$7772 ( \7904 , \7761 , \7880 );
and \U$7773 ( \7905 , \7655 , \7880 );
or \U$7774 ( \7906 , \7903 , \7904 , \7905 );
xor \U$7775 ( \7907 , \7902 , \7906 );
and \U$7776 ( \7908 , \7659 , \7663 );
and \U$7777 ( \7909 , \7663 , \7668 );
and \U$7778 ( \7910 , \7659 , \7668 );
or \U$7779 ( \7911 , \7908 , \7909 , \7910 );
and \U$7780 ( \7912 , \7673 , \7677 );
and \U$7781 ( \7913 , \7677 , \7682 );
and \U$7782 ( \7914 , \7673 , \7682 );
or \U$7783 ( \7915 , \7912 , \7913 , \7914 );
xor \U$7784 ( \7916 , \7911 , \7915 );
and \U$7785 ( \7917 , \7698 , \7714 );
and \U$7786 ( \7918 , \7714 , \7759 );
and \U$7787 ( \7919 , \7698 , \7759 );
or \U$7788 ( \7920 , \7917 , \7918 , \7919 );
xor \U$7789 ( \7921 , \7916 , \7920 );
xor \U$7790 ( \7922 , \7907 , \7921 );
xor \U$7791 ( \7923 , \7898 , \7922 );
and \U$7792 ( \7924 , \7645 , \7649 );
and \U$7793 ( \7925 , \7649 , \7654 );
and \U$7794 ( \7926 , \7645 , \7654 );
or \U$7795 ( \7927 , \7924 , \7925 , \7926 );
and \U$7796 ( \7928 , \7669 , \7683 );
and \U$7797 ( \7929 , \7683 , \7760 );
and \U$7798 ( \7930 , \7669 , \7760 );
or \U$7799 ( \7931 , \7928 , \7929 , \7930 );
xor \U$7800 ( \7932 , \7927 , \7931 );
and \U$7801 ( \7933 , \7766 , \7849 );
and \U$7802 ( \7934 , \7849 , \7879 );
and \U$7803 ( \7935 , \7766 , \7879 );
or \U$7804 ( \7936 , \7933 , \7934 , \7935 );
xor \U$7805 ( \7937 , \7932 , \7936 );
and \U$7806 ( \7938 , \7770 , \7774 );
and \U$7807 ( \7939 , \7774 , \7779 );
and \U$7808 ( \7940 , \7770 , \7779 );
or \U$7809 ( \7941 , \7938 , \7939 , \7940 );
and \U$7810 ( \7942 , \7854 , \7858 );
and \U$7811 ( \7943 , \7858 , \7863 );
and \U$7812 ( \7944 , \7854 , \7863 );
or \U$7813 ( \7945 , \7942 , \7943 , \7944 );
xor \U$7814 ( \7946 , \7941 , \7945 );
and \U$7815 ( \7947 , \7868 , \7872 );
and \U$7816 ( \7948 , \7872 , \7877 );
and \U$7817 ( \7949 , \7868 , \7877 );
or \U$7818 ( \7950 , \7947 , \7948 , \7949 );
xor \U$7819 ( \7951 , \7946 , \7950 );
and \U$7820 ( \7952 , \7780 , \7824 );
and \U$7821 ( \7953 , \7824 , \7848 );
and \U$7822 ( \7954 , \7780 , \7848 );
or \U$7823 ( \7955 , \7952 , \7953 , \7954 );
and \U$7824 ( \7956 , \7864 , \7878 );
xor \U$7825 ( \7957 , \7955 , \7956 );
and \U$7826 ( \7958 , \7719 , \7723 );
and \U$7827 ( \7959 , \7723 , \7728 );
and \U$7828 ( \7960 , \7719 , \7728 );
or \U$7829 ( \7961 , \7958 , \7959 , \7960 );
and \U$7830 ( \7962 , \7688 , \7692 );
and \U$7831 ( \7963 , \7692 , \7697 );
and \U$7832 ( \7964 , \7688 , \7697 );
or \U$7833 ( \7965 , \7962 , \7963 , \7964 );
xor \U$7834 ( \7966 , \7961 , \7965 );
and \U$7835 ( \7967 , \7703 , \7707 );
and \U$7836 ( \7968 , \7707 , \7713 );
and \U$7837 ( \7969 , \7703 , \7713 );
or \U$7838 ( \7970 , \7967 , \7968 , \7969 );
xor \U$7839 ( \7971 , \7966 , \7970 );
xor \U$7840 ( \7972 , \7957 , \7971 );
xor \U$7841 ( \7973 , \7951 , \7972 );
and \U$7842 ( \7974 , \7794 , \7808 );
and \U$7843 ( \7975 , \7808 , \7823 );
and \U$7844 ( \7976 , \7794 , \7823 );
or \U$7845 ( \7977 , \7974 , \7975 , \7976 );
and \U$7846 ( \7978 , \7829 , \7832 );
and \U$7847 ( \7979 , \7832 , \7847 );
and \U$7848 ( \7980 , \7829 , \7847 );
or \U$7849 ( \7981 , \7978 , \7979 , \7980 );
xor \U$7850 ( \7982 , \7977 , \7981 );
and \U$7851 ( \7983 , \7729 , \7743 );
and \U$7852 ( \7984 , \7743 , \7758 );
and \U$7853 ( \7985 , \7729 , \7758 );
or \U$7854 ( \7986 , \7983 , \7984 , \7985 );
xor \U$7855 ( \7987 , \7982 , \7986 );
and \U$7856 ( \7988 , \7837 , \7841 );
and \U$7857 ( \7989 , \7841 , \7846 );
and \U$7858 ( \7990 , \7837 , \7846 );
or \U$7859 ( \7991 , \7988 , \7989 , \7990 );
and \U$7860 ( \7992 , \7798 , \7802 );
and \U$7861 ( \7993 , \7802 , \7807 );
and \U$7862 ( \7994 , \7798 , \7807 );
or \U$7863 ( \7995 , \7992 , \7993 , \7994 );
xor \U$7864 ( \7996 , \7991 , \7995 );
and \U$7865 ( \7997 , \7813 , \7817 );
and \U$7866 ( \7998 , \7817 , \7822 );
and \U$7867 ( \7999 , \7813 , \7822 );
or \U$7868 ( \8000 , \7997 , \7998 , \7999 );
xor \U$7869 ( \8001 , \7996 , \8000 );
and \U$7870 ( \8002 , \7784 , \7788 );
and \U$7871 ( \8003 , \7788 , \7793 );
and \U$7872 ( \8004 , \7784 , \7793 );
or \U$7873 ( \8005 , \8002 , \8003 , \8004 );
and \U$7874 ( \8006 , \7733 , \7737 );
and \U$7875 ( \8007 , \7737 , \7742 );
and \U$7876 ( \8008 , \7733 , \7742 );
or \U$7877 ( \8009 , \8006 , \8007 , \8008 );
xor \U$7878 ( \8010 , \8005 , \8009 );
and \U$7879 ( \8011 , \7748 , \7752 );
and \U$7880 ( \8012 , \7752 , \7757 );
and \U$7881 ( \8013 , \7748 , \7757 );
or \U$7882 ( \8014 , \8011 , \8012 , \8013 );
xor \U$7883 ( \8015 , \8010 , \8014 );
xor \U$7884 ( \8016 , \8001 , \8015 );
xor \U$7885 ( \8017 , \7709 , \7710 );
not \U$7886 ( \8018 , \7830 );
and \U$7887 ( \8019 , \8017 , \8018 );
and \U$7888 ( \8020 , \166 , \8019 );
and \U$7889 ( \8021 , \150 , \7830 );
nor \U$7890 ( \8022 , \8020 , \8021 );
xnor \U$7891 ( \8023 , \8022 , \7713 );
and \U$7892 ( \8024 , \247 , \6401 );
and \U$7893 ( \8025 , \224 , \6143 );
nor \U$7894 ( \8026 , \8024 , \8025 );
xnor \U$7895 ( \8027 , \8026 , \6148 );
and \U$7896 ( \8028 , \143 , \7055 );
and \U$7897 ( \8029 , \240 , \6675 );
nor \U$7898 ( \8030 , \8028 , \8029 );
xnor \U$7899 ( \8031 , \8030 , \6680 );
xor \U$7900 ( \8032 , \8027 , \8031 );
and \U$7901 ( \8033 , \158 , \7489 );
and \U$7902 ( \8034 , \134 , \7137 );
nor \U$7903 ( \8035 , \8033 , \8034 );
xnor \U$7904 ( \8036 , \8035 , \7142 );
xor \U$7905 ( \8037 , \8032 , \8036 );
xor \U$7906 ( \8038 , \8023 , \8037 );
and \U$7907 ( \8039 , \197 , \5011 );
and \U$7908 ( \8040 , \178 , \4878 );
nor \U$7909 ( \8041 , \8039 , \8040 );
xnor \U$7910 ( \8042 , \8041 , \4762 );
and \U$7911 ( \8043 , \217 , \5485 );
and \U$7912 ( \8044 , \189 , \5275 );
nor \U$7913 ( \8045 , \8043 , \8044 );
xnor \U$7914 ( \8046 , \8045 , \5169 );
xor \U$7915 ( \8047 , \8042 , \8046 );
and \U$7916 ( \8048 , \232 , \5996 );
and \U$7917 ( \8049 , \209 , \5695 );
nor \U$7918 ( \8050 , \8048 , \8049 );
xnor \U$7919 ( \8051 , \8050 , \5687 );
xor \U$7920 ( \8052 , \8047 , \8051 );
xor \U$7921 ( \8053 , \8038 , \8052 );
xor \U$7922 ( \8054 , \8016 , \8053 );
xor \U$7923 ( \8055 , \7987 , \8054 );
and \U$7924 ( \8056 , \7700 , \183 );
buf \U$7925 ( \8057 , RIb55ee00_73);
and \U$7926 ( \8058 , \8057 , \180 );
nor \U$7927 ( \8059 , \8056 , \8058 );
xnor \U$7928 ( \8060 , \8059 , \179 );
and \U$7929 ( \8061 , \7231 , \195 );
and \U$7930 ( \8062 , \7556 , \193 );
nor \U$7931 ( \8063 , \8061 , \8062 );
xnor \U$7932 ( \8064 , \8063 , \202 );
xor \U$7933 ( \8065 , \8060 , \8064 );
and \U$7934 ( \8066 , \6790 , \215 );
and \U$7935 ( \8067 , \6945 , \213 );
nor \U$7936 ( \8068 , \8066 , \8067 );
xnor \U$7937 ( \8069 , \8068 , \222 );
xor \U$7938 ( \8070 , \8065 , \8069 );
and \U$7939 ( \8071 , \1684 , \2669 );
and \U$7940 ( \8072 , \1802 , \2538 );
nor \U$7941 ( \8073 , \8071 , \8072 );
xnor \U$7942 ( \8074 , \8073 , \2534 );
and \U$7943 ( \8075 , \1484 , \3103 );
and \U$7944 ( \8076 , \1601 , \2934 );
nor \U$7945 ( \8077 , \8075 , \8076 );
xnor \U$7946 ( \8078 , \8077 , \2839 );
xor \U$7947 ( \8079 , \8074 , \8078 );
and \U$7948 ( \8080 , \1192 , \3357 );
and \U$7949 ( \8081 , \1333 , \3255 );
nor \U$7950 ( \8082 , \8080 , \8081 );
xnor \U$7951 ( \8083 , \8082 , \3156 );
xor \U$7952 ( \8084 , \8079 , \8083 );
and \U$7953 ( \8085 , \2521 , \1824 );
and \U$7954 ( \8086 , \2757 , \1739 );
nor \U$7955 ( \8087 , \8085 , \8086 );
xnor \U$7956 ( \8088 , \8087 , \1697 );
and \U$7957 ( \8089 , \2182 , \2121 );
and \U$7958 ( \8090 , \2366 , \2008 );
nor \U$7959 ( \8091 , \8089 , \8090 );
xnor \U$7960 ( \8092 , \8091 , \1961 );
xor \U$7961 ( \8093 , \8088 , \8092 );
and \U$7962 ( \8094 , \1948 , \2400 );
and \U$7963 ( \8095 , \2090 , \2246 );
nor \U$7964 ( \8096 , \8094 , \8095 );
xnor \U$7965 ( \8097 , \8096 , \2195 );
xor \U$7966 ( \8098 , \8093 , \8097 );
xor \U$7967 ( \8099 , \8084 , \8098 );
and \U$7968 ( \8100 , \474 , \3813 );
and \U$7969 ( \8101 , \1147 , \3557 );
nor \U$7970 ( \8102 , \8100 , \8101 );
xnor \U$7971 ( \8103 , \8102 , \3562 );
and \U$7972 ( \8104 , \307 , \4132 );
and \U$7973 ( \8105 , \412 , \4012 );
nor \U$7974 ( \8106 , \8104 , \8105 );
xnor \U$7975 ( \8107 , \8106 , \3925 );
xor \U$7976 ( \8108 , \8103 , \8107 );
and \U$7977 ( \8109 , \185 , \4581 );
and \U$7978 ( \8110 , \261 , \4424 );
nor \U$7979 ( \8111 , \8109 , \8110 );
xnor \U$7980 ( \8112 , \8111 , \4377 );
xor \U$7981 ( \8113 , \8108 , \8112 );
xor \U$7982 ( \8114 , \8099 , \8113 );
xor \U$7983 ( \8115 , \8070 , \8114 );
and \U$7984 ( \8116 , \3646 , \1086 );
and \U$7985 ( \8117 , \3736 , \508 );
nor \U$7986 ( \8118 , \8116 , \8117 );
xnor \U$7987 ( \8119 , \8118 , \487 );
and \U$7988 ( \8120 , \3143 , \1301 );
and \U$7989 ( \8121 , \3395 , \1246 );
nor \U$7990 ( \8122 , \8120 , \8121 );
xnor \U$7991 ( \8123 , \8122 , \1205 );
xor \U$7992 ( \8124 , \8119 , \8123 );
and \U$7993 ( \8125 , \2826 , \1578 );
and \U$7994 ( \8126 , \3037 , \1431 );
nor \U$7995 ( \8127 , \8125 , \8126 );
xnor \U$7996 ( \8128 , \8127 , \1436 );
xor \U$7997 ( \8129 , \8124 , \8128 );
and \U$7998 ( \8130 , \4749 , \156 );
and \U$7999 ( \8131 , \4922 , \154 );
nor \U$8000 ( \8132 , \8130 , \8131 );
xnor \U$8001 ( \8133 , \8132 , \163 );
and \U$8002 ( \8134 , \4364 , \296 );
and \U$8003 ( \8135 , \4654 , \168 );
nor \U$8004 ( \8136 , \8134 , \8135 );
xnor \U$8005 ( \8137 , \8136 , \173 );
xor \U$8006 ( \8138 , \8133 , \8137 );
and \U$8007 ( \8139 , \3912 , \438 );
and \U$8008 ( \8140 , \4160 , \336 );
nor \U$8009 ( \8141 , \8139 , \8140 );
xnor \U$8010 ( \8142 , \8141 , \320 );
xor \U$8011 ( \8143 , \8138 , \8142 );
xor \U$8012 ( \8144 , \8129 , \8143 );
and \U$8013 ( \8145 , \6281 , \230 );
and \U$8014 ( \8146 , \6514 , \228 );
nor \U$8015 ( \8147 , \8145 , \8146 );
xnor \U$8016 ( \8148 , \8147 , \237 );
and \U$8017 ( \8149 , \5674 , \245 );
and \U$8018 ( \8150 , \6030 , \243 );
nor \U$8019 ( \8151 , \8149 , \8150 );
xnor \U$8020 ( \8152 , \8151 , \252 );
xor \U$8021 ( \8153 , \8148 , \8152 );
and \U$8022 ( \8154 , \5156 , \141 );
and \U$8023 ( \8155 , \5469 , \139 );
nor \U$8024 ( \8156 , \8154 , \8155 );
xnor \U$8025 ( \8157 , \8156 , \148 );
xor \U$8026 ( \8158 , \8153 , \8157 );
xor \U$8027 ( \8159 , \8144 , \8158 );
xor \U$8028 ( \8160 , \8115 , \8159 );
xor \U$8029 ( \8161 , \8055 , \8160 );
xor \U$8030 ( \8162 , \7973 , \8161 );
xor \U$8031 ( \8163 , \7937 , \8162 );
xor \U$8032 ( \8164 , \7923 , \8163 );
and \U$8033 ( \8165 , \7620 , \7631 );
and \U$8034 ( \8166 , \7631 , \7882 );
and \U$8035 ( \8167 , \7620 , \7882 );
or \U$8036 ( \8168 , \8165 , \8166 , \8167 );
xor \U$8037 ( \8169 , \8164 , \8168 );
and \U$8038 ( \8170 , \7883 , \7887 );
and \U$8039 ( \8171 , \7888 , \7891 );
or \U$8040 ( \8172 , \8170 , \8171 );
xor \U$8041 ( \8173 , \8169 , \8172 );
buf \U$8042 ( \8174 , \8173 );
buf \U$8043 ( \8175 , \8174 );
and \U$8044 ( \8176 , \7902 , \7906 );
and \U$8045 ( \8177 , \7906 , \7921 );
and \U$8046 ( \8178 , \7902 , \7921 );
or \U$8047 ( \8179 , \8176 , \8177 , \8178 );
and \U$8048 ( \8180 , \7937 , \8162 );
xor \U$8049 ( \8181 , \8179 , \8180 );
and \U$8050 ( \8182 , \7911 , \7915 );
and \U$8051 ( \8183 , \7915 , \7920 );
and \U$8052 ( \8184 , \7911 , \7920 );
or \U$8053 ( \8185 , \8182 , \8183 , \8184 );
and \U$8054 ( \8186 , \7955 , \7956 );
and \U$8055 ( \8187 , \7956 , \7971 );
and \U$8056 ( \8188 , \7955 , \7971 );
or \U$8057 ( \8189 , \8186 , \8187 , \8188 );
xor \U$8058 ( \8190 , \8185 , \8189 );
and \U$8059 ( \8191 , \7987 , \8054 );
and \U$8060 ( \8192 , \8054 , \8160 );
and \U$8061 ( \8193 , \7987 , \8160 );
or \U$8062 ( \8194 , \8191 , \8192 , \8193 );
xor \U$8063 ( \8195 , \8190 , \8194 );
xor \U$8064 ( \8196 , \8181 , \8195 );
and \U$8065 ( \8197 , \7927 , \7931 );
and \U$8066 ( \8198 , \7931 , \7936 );
and \U$8067 ( \8199 , \7927 , \7936 );
or \U$8068 ( \8200 , \8197 , \8198 , \8199 );
and \U$8069 ( \8201 , \7951 , \7972 );
and \U$8070 ( \8202 , \7972 , \8161 );
and \U$8071 ( \8203 , \7951 , \8161 );
or \U$8072 ( \8204 , \8201 , \8202 , \8203 );
xor \U$8073 ( \8205 , \8200 , \8204 );
and \U$8074 ( \8206 , \7977 , \7981 );
and \U$8075 ( \8207 , \7981 , \7986 );
and \U$8076 ( \8208 , \7977 , \7986 );
or \U$8077 ( \8209 , \8206 , \8207 , \8208 );
and \U$8078 ( \8210 , \7941 , \7945 );
and \U$8079 ( \8211 , \7945 , \7950 );
and \U$8080 ( \8212 , \7941 , \7950 );
or \U$8081 ( \8213 , \8210 , \8211 , \8212 );
xor \U$8082 ( \8214 , \8209 , \8213 );
and \U$8083 ( \8215 , \8070 , \8114 );
and \U$8084 ( \8216 , \8114 , \8159 );
and \U$8085 ( \8217 , \8070 , \8159 );
or \U$8086 ( \8218 , \8215 , \8216 , \8217 );
xor \U$8087 ( \8219 , \8214 , \8218 );
and \U$8088 ( \8220 , \8001 , \8015 );
and \U$8089 ( \8221 , \8015 , \8053 );
and \U$8090 ( \8222 , \8001 , \8053 );
or \U$8091 ( \8223 , \8220 , \8221 , \8222 );
and \U$8092 ( \8224 , \8133 , \8137 );
and \U$8093 ( \8225 , \8137 , \8142 );
and \U$8094 ( \8226 , \8133 , \8142 );
or \U$8095 ( \8227 , \8224 , \8225 , \8226 );
and \U$8096 ( \8228 , \8060 , \8064 );
and \U$8097 ( \8229 , \8064 , \8069 );
and \U$8098 ( \8230 , \8060 , \8069 );
or \U$8099 ( \8231 , \8228 , \8229 , \8230 );
xor \U$8100 ( \8232 , \8227 , \8231 );
and \U$8101 ( \8233 , \8148 , \8152 );
and \U$8102 ( \8234 , \8152 , \8157 );
and \U$8103 ( \8235 , \8148 , \8157 );
or \U$8104 ( \8236 , \8233 , \8234 , \8235 );
xor \U$8105 ( \8237 , \8232 , \8236 );
xor \U$8106 ( \8238 , \8223 , \8237 );
and \U$8107 ( \8239 , \8119 , \8123 );
and \U$8108 ( \8240 , \8123 , \8128 );
and \U$8109 ( \8241 , \8119 , \8128 );
or \U$8110 ( \8242 , \8239 , \8240 , \8241 );
and \U$8111 ( \8243 , \8074 , \8078 );
and \U$8112 ( \8244 , \8078 , \8083 );
and \U$8113 ( \8245 , \8074 , \8083 );
or \U$8114 ( \8246 , \8243 , \8244 , \8245 );
xor \U$8115 ( \8247 , \8242 , \8246 );
and \U$8116 ( \8248 , \8088 , \8092 );
and \U$8117 ( \8249 , \8092 , \8097 );
and \U$8118 ( \8250 , \8088 , \8097 );
or \U$8119 ( \8251 , \8248 , \8249 , \8250 );
xor \U$8120 ( \8252 , \8247 , \8251 );
and \U$8121 ( \8253 , \8027 , \8031 );
and \U$8122 ( \8254 , \8031 , \8036 );
and \U$8123 ( \8255 , \8027 , \8036 );
or \U$8124 ( \8256 , \8253 , \8254 , \8255 );
and \U$8125 ( \8257 , \8042 , \8046 );
and \U$8126 ( \8258 , \8046 , \8051 );
and \U$8127 ( \8259 , \8042 , \8051 );
or \U$8128 ( \8260 , \8257 , \8258 , \8259 );
xor \U$8129 ( \8261 , \8256 , \8260 );
and \U$8130 ( \8262 , \8103 , \8107 );
and \U$8131 ( \8263 , \8107 , \8112 );
and \U$8132 ( \8264 , \8103 , \8112 );
or \U$8133 ( \8265 , \8262 , \8263 , \8264 );
xor \U$8134 ( \8266 , \8261 , \8265 );
xor \U$8135 ( \8267 , \8252 , \8266 );
and \U$8136 ( \8268 , \261 , \4581 );
and \U$8137 ( \8269 , \307 , \4424 );
nor \U$8138 ( \8270 , \8268 , \8269 );
xnor \U$8139 ( \8271 , \8270 , \4377 );
and \U$8140 ( \8272 , \178 , \5011 );
and \U$8141 ( \8273 , \185 , \4878 );
nor \U$8142 ( \8274 , \8272 , \8273 );
xnor \U$8143 ( \8275 , \8274 , \4762 );
xor \U$8144 ( \8276 , \8271 , \8275 );
and \U$8145 ( \8277 , \189 , \5485 );
and \U$8146 ( \8278 , \197 , \5275 );
nor \U$8147 ( \8279 , \8277 , \8278 );
xnor \U$8148 ( \8280 , \8279 , \5169 );
xor \U$8149 ( \8281 , \8276 , \8280 );
and \U$8150 ( \8282 , \134 , \7489 );
and \U$8151 ( \8283 , \143 , \7137 );
nor \U$8152 ( \8284 , \8282 , \8283 );
xnor \U$8153 ( \8285 , \8284 , \7142 );
and \U$8154 ( \8286 , \150 , \8019 );
and \U$8155 ( \8287 , \158 , \7830 );
nor \U$8156 ( \8288 , \8286 , \8287 );
xnor \U$8157 ( \8289 , \8288 , \7713 );
xor \U$8158 ( \8290 , \8285 , \8289 );
buf \U$8159 ( \8291 , RIb560c78_8);
xor \U$8160 ( \8292 , \8291 , \7709 );
nand \U$8161 ( \8293 , \166 , \8292 );
buf \U$8162 ( \8294 , RIb560cf0_7);
and \U$8163 ( \8295 , \8291 , \7709 );
not \U$8164 ( \8296 , \8295 );
and \U$8165 ( \8297 , \8294 , \8296 );
xnor \U$8166 ( \8298 , \8293 , \8297 );
xor \U$8167 ( \8299 , \8290 , \8298 );
xor \U$8168 ( \8300 , \8281 , \8299 );
and \U$8169 ( \8301 , \209 , \5996 );
and \U$8170 ( \8302 , \217 , \5695 );
nor \U$8171 ( \8303 , \8301 , \8302 );
xnor \U$8172 ( \8304 , \8303 , \5687 );
and \U$8173 ( \8305 , \224 , \6401 );
and \U$8174 ( \8306 , \232 , \6143 );
nor \U$8175 ( \8307 , \8305 , \8306 );
xnor \U$8176 ( \8308 , \8307 , \6148 );
xor \U$8177 ( \8309 , \8304 , \8308 );
and \U$8178 ( \8310 , \240 , \7055 );
and \U$8179 ( \8311 , \247 , \6675 );
nor \U$8180 ( \8312 , \8310 , \8311 );
xnor \U$8181 ( \8313 , \8312 , \6680 );
xor \U$8182 ( \8314 , \8309 , \8313 );
xor \U$8183 ( \8315 , \8300 , \8314 );
xor \U$8184 ( \8316 , \8267 , \8315 );
xor \U$8185 ( \8317 , \8238 , \8316 );
xor \U$8186 ( \8318 , \8219 , \8317 );
and \U$8187 ( \8319 , \8084 , \8098 );
and \U$8188 ( \8320 , \8098 , \8113 );
and \U$8189 ( \8321 , \8084 , \8113 );
or \U$8190 ( \8322 , \8319 , \8320 , \8321 );
and \U$8191 ( \8323 , \8129 , \8143 );
and \U$8192 ( \8324 , \8143 , \8158 );
and \U$8193 ( \8325 , \8129 , \8158 );
or \U$8194 ( \8326 , \8323 , \8324 , \8325 );
xor \U$8195 ( \8327 , \8322 , \8326 );
and \U$8196 ( \8328 , \8023 , \8037 );
and \U$8197 ( \8329 , \8037 , \8052 );
and \U$8198 ( \8330 , \8023 , \8052 );
or \U$8199 ( \8331 , \8328 , \8329 , \8330 );
xor \U$8200 ( \8332 , \8327 , \8331 );
and \U$8201 ( \8333 , \7961 , \7965 );
and \U$8202 ( \8334 , \7965 , \7970 );
and \U$8203 ( \8335 , \7961 , \7970 );
or \U$8204 ( \8336 , \8333 , \8334 , \8335 );
and \U$8205 ( \8337 , \7991 , \7995 );
and \U$8206 ( \8338 , \7995 , \8000 );
and \U$8207 ( \8339 , \7991 , \8000 );
or \U$8208 ( \8340 , \8337 , \8338 , \8339 );
xor \U$8209 ( \8341 , \8336 , \8340 );
and \U$8210 ( \8342 , \8005 , \8009 );
and \U$8211 ( \8343 , \8009 , \8014 );
and \U$8212 ( \8344 , \8005 , \8014 );
or \U$8213 ( \8345 , \8342 , \8343 , \8344 );
xor \U$8214 ( \8346 , \8341 , \8345 );
xor \U$8215 ( \8347 , \8332 , \8346 );
and \U$8216 ( \8348 , \8057 , \183 );
buf \U$8217 ( \8349 , RIb55ee78_72);
and \U$8218 ( \8350 , \8349 , \180 );
nor \U$8219 ( \8351 , \8348 , \8350 );
xnor \U$8220 ( \8352 , \8351 , \179 );
and \U$8221 ( \8353 , \7556 , \195 );
and \U$8222 ( \8354 , \7700 , \193 );
nor \U$8223 ( \8355 , \8353 , \8354 );
xnor \U$8224 ( \8356 , \8355 , \202 );
xor \U$8225 ( \8357 , \8352 , \8356 );
xor \U$8226 ( \8358 , \8357 , \8297 );
and \U$8227 ( \8359 , \6945 , \215 );
and \U$8228 ( \8360 , \7231 , \213 );
nor \U$8229 ( \8361 , \8359 , \8360 );
xnor \U$8230 ( \8362 , \8361 , \222 );
and \U$8231 ( \8363 , \6514 , \230 );
and \U$8232 ( \8364 , \6790 , \228 );
nor \U$8233 ( \8365 , \8363 , \8364 );
xnor \U$8234 ( \8366 , \8365 , \237 );
xor \U$8235 ( \8367 , \8362 , \8366 );
and \U$8236 ( \8368 , \6030 , \245 );
and \U$8237 ( \8369 , \6281 , \243 );
nor \U$8238 ( \8370 , \8368 , \8369 );
xnor \U$8239 ( \8371 , \8370 , \252 );
xor \U$8240 ( \8372 , \8367 , \8371 );
and \U$8241 ( \8373 , \5469 , \141 );
and \U$8242 ( \8374 , \5674 , \139 );
nor \U$8243 ( \8375 , \8373 , \8374 );
xnor \U$8244 ( \8376 , \8375 , \148 );
and \U$8245 ( \8377 , \4922 , \156 );
and \U$8246 ( \8378 , \5156 , \154 );
nor \U$8247 ( \8379 , \8377 , \8378 );
xnor \U$8248 ( \8380 , \8379 , \163 );
xor \U$8249 ( \8381 , \8376 , \8380 );
and \U$8250 ( \8382 , \4654 , \296 );
and \U$8251 ( \8383 , \4749 , \168 );
nor \U$8252 ( \8384 , \8382 , \8383 );
xnor \U$8253 ( \8385 , \8384 , \173 );
xor \U$8254 ( \8386 , \8381 , \8385 );
xor \U$8255 ( \8387 , \8372 , \8386 );
and \U$8256 ( \8388 , \4160 , \438 );
and \U$8257 ( \8389 , \4364 , \336 );
nor \U$8258 ( \8390 , \8388 , \8389 );
xnor \U$8259 ( \8391 , \8390 , \320 );
and \U$8260 ( \8392 , \3736 , \1086 );
and \U$8261 ( \8393 , \3912 , \508 );
nor \U$8262 ( \8394 , \8392 , \8393 );
xnor \U$8263 ( \8395 , \8394 , \487 );
xor \U$8264 ( \8396 , \8391 , \8395 );
and \U$8265 ( \8397 , \3395 , \1301 );
and \U$8266 ( \8398 , \3646 , \1246 );
nor \U$8267 ( \8399 , \8397 , \8398 );
xnor \U$8268 ( \8400 , \8399 , \1205 );
xor \U$8269 ( \8401 , \8396 , \8400 );
xor \U$8270 ( \8402 , \8387 , \8401 );
xor \U$8271 ( \8403 , \8358 , \8402 );
and \U$8272 ( \8404 , \2090 , \2400 );
and \U$8273 ( \8405 , \2182 , \2246 );
nor \U$8274 ( \8406 , \8404 , \8405 );
xnor \U$8275 ( \8407 , \8406 , \2195 );
and \U$8276 ( \8408 , \1802 , \2669 );
and \U$8277 ( \8409 , \1948 , \2538 );
nor \U$8278 ( \8410 , \8408 , \8409 );
xnor \U$8279 ( \8411 , \8410 , \2534 );
xor \U$8280 ( \8412 , \8407 , \8411 );
and \U$8281 ( \8413 , \1601 , \3103 );
and \U$8282 ( \8414 , \1684 , \2934 );
nor \U$8283 ( \8415 , \8413 , \8414 );
xnor \U$8284 ( \8416 , \8415 , \2839 );
xor \U$8285 ( \8417 , \8412 , \8416 );
and \U$8286 ( \8418 , \3037 , \1578 );
and \U$8287 ( \8419 , \3143 , \1431 );
nor \U$8288 ( \8420 , \8418 , \8419 );
xnor \U$8289 ( \8421 , \8420 , \1436 );
and \U$8290 ( \8422 , \2757 , \1824 );
and \U$8291 ( \8423 , \2826 , \1739 );
nor \U$8292 ( \8424 , \8422 , \8423 );
xnor \U$8293 ( \8425 , \8424 , \1697 );
xor \U$8294 ( \8426 , \8421 , \8425 );
and \U$8295 ( \8427 , \2366 , \2121 );
and \U$8296 ( \8428 , \2521 , \2008 );
nor \U$8297 ( \8429 , \8427 , \8428 );
xnor \U$8298 ( \8430 , \8429 , \1961 );
xor \U$8299 ( \8431 , \8426 , \8430 );
xor \U$8300 ( \8432 , \8417 , \8431 );
and \U$8301 ( \8433 , \1333 , \3357 );
and \U$8302 ( \8434 , \1484 , \3255 );
nor \U$8303 ( \8435 , \8433 , \8434 );
xnor \U$8304 ( \8436 , \8435 , \3156 );
and \U$8305 ( \8437 , \1147 , \3813 );
and \U$8306 ( \8438 , \1192 , \3557 );
nor \U$8307 ( \8439 , \8437 , \8438 );
xnor \U$8308 ( \8440 , \8439 , \3562 );
xor \U$8309 ( \8441 , \8436 , \8440 );
and \U$8310 ( \8442 , \412 , \4132 );
and \U$8311 ( \8443 , \474 , \4012 );
nor \U$8312 ( \8444 , \8442 , \8443 );
xnor \U$8313 ( \8445 , \8444 , \3925 );
xor \U$8314 ( \8446 , \8441 , \8445 );
xor \U$8315 ( \8447 , \8432 , \8446 );
xor \U$8316 ( \8448 , \8403 , \8447 );
xor \U$8317 ( \8449 , \8347 , \8448 );
xor \U$8318 ( \8450 , \8318 , \8449 );
xor \U$8319 ( \8451 , \8205 , \8450 );
xor \U$8320 ( \8452 , \8196 , \8451 );
and \U$8321 ( \8453 , \7898 , \7922 );
and \U$8322 ( \8454 , \7922 , \8163 );
and \U$8323 ( \8455 , \7898 , \8163 );
or \U$8324 ( \8456 , \8453 , \8454 , \8455 );
xor \U$8325 ( \8457 , \8452 , \8456 );
and \U$8326 ( \8458 , \8164 , \8168 );
and \U$8327 ( \8459 , \8169 , \8172 );
or \U$8328 ( \8460 , \8458 , \8459 );
xor \U$8329 ( \8461 , \8457 , \8460 );
buf \U$8330 ( \8462 , \8461 );
buf \U$8331 ( \8463 , \8462 );
and \U$8332 ( \8464 , \8179 , \8180 );
and \U$8333 ( \8465 , \8180 , \8195 );
and \U$8334 ( \8466 , \8179 , \8195 );
or \U$8335 ( \8467 , \8464 , \8465 , \8466 );
and \U$8336 ( \8468 , \8200 , \8204 );
and \U$8337 ( \8469 , \8204 , \8450 );
and \U$8338 ( \8470 , \8200 , \8450 );
or \U$8339 ( \8471 , \8468 , \8469 , \8470 );
and \U$8340 ( \8472 , \8209 , \8213 );
and \U$8341 ( \8473 , \8213 , \8218 );
and \U$8342 ( \8474 , \8209 , \8218 );
or \U$8343 ( \8475 , \8472 , \8473 , \8474 );
and \U$8344 ( \8476 , \8223 , \8237 );
and \U$8345 ( \8477 , \8237 , \8316 );
and \U$8346 ( \8478 , \8223 , \8316 );
or \U$8347 ( \8479 , \8476 , \8477 , \8478 );
xor \U$8348 ( \8480 , \8475 , \8479 );
and \U$8349 ( \8481 , \8332 , \8346 );
and \U$8350 ( \8482 , \8346 , \8448 );
and \U$8351 ( \8483 , \8332 , \8448 );
or \U$8352 ( \8484 , \8481 , \8482 , \8483 );
xor \U$8353 ( \8485 , \8480 , \8484 );
xor \U$8354 ( \8486 , \8471 , \8485 );
and \U$8355 ( \8487 , \8185 , \8189 );
and \U$8356 ( \8488 , \8189 , \8194 );
and \U$8357 ( \8489 , \8185 , \8194 );
or \U$8358 ( \8490 , \8487 , \8488 , \8489 );
and \U$8359 ( \8491 , \8219 , \8317 );
and \U$8360 ( \8492 , \8317 , \8449 );
and \U$8361 ( \8493 , \8219 , \8449 );
or \U$8362 ( \8494 , \8491 , \8492 , \8493 );
xor \U$8363 ( \8495 , \8490 , \8494 );
and \U$8364 ( \8496 , \8322 , \8326 );
and \U$8365 ( \8497 , \8326 , \8331 );
and \U$8366 ( \8498 , \8322 , \8331 );
or \U$8367 ( \8499 , \8496 , \8497 , \8498 );
and \U$8368 ( \8500 , \8336 , \8340 );
and \U$8369 ( \8501 , \8340 , \8345 );
and \U$8370 ( \8502 , \8336 , \8345 );
or \U$8371 ( \8503 , \8500 , \8501 , \8502 );
xor \U$8372 ( \8504 , \8499 , \8503 );
and \U$8373 ( \8505 , \8358 , \8402 );
and \U$8374 ( \8506 , \8402 , \8447 );
and \U$8375 ( \8507 , \8358 , \8447 );
or \U$8376 ( \8508 , \8505 , \8506 , \8507 );
xor \U$8377 ( \8509 , \8504 , \8508 );
and \U$8378 ( \8510 , \8252 , \8266 );
and \U$8379 ( \8511 , \8266 , \8315 );
and \U$8380 ( \8512 , \8252 , \8315 );
or \U$8381 ( \8513 , \8510 , \8511 , \8512 );
and \U$8382 ( \8514 , \8362 , \8366 );
and \U$8383 ( \8515 , \8366 , \8371 );
and \U$8384 ( \8516 , \8362 , \8371 );
or \U$8385 ( \8517 , \8514 , \8515 , \8516 );
and \U$8386 ( \8518 , \8376 , \8380 );
and \U$8387 ( \8519 , \8380 , \8385 );
and \U$8388 ( \8520 , \8376 , \8385 );
or \U$8389 ( \8521 , \8518 , \8519 , \8520 );
xor \U$8390 ( \8522 , \8517 , \8521 );
and \U$8391 ( \8523 , \8352 , \8356 );
and \U$8392 ( \8524 , \8356 , \8297 );
and \U$8393 ( \8525 , \8352 , \8297 );
or \U$8394 ( \8526 , \8523 , \8524 , \8525 );
xor \U$8395 ( \8527 , \8522 , \8526 );
xor \U$8396 ( \8528 , \8513 , \8527 );
and \U$8397 ( \8529 , \8285 , \8289 );
and \U$8398 ( \8530 , \8289 , \8298 );
and \U$8399 ( \8531 , \8285 , \8298 );
or \U$8400 ( \8532 , \8529 , \8530 , \8531 );
and \U$8401 ( \8533 , \158 , \8019 );
and \U$8402 ( \8534 , \134 , \7830 );
nor \U$8403 ( \8535 , \8533 , \8534 );
xnor \U$8404 ( \8536 , \8535 , \7713 );
xor \U$8405 ( \8537 , \8532 , \8536 );
xor \U$8406 ( \8538 , \8294 , \8291 );
not \U$8407 ( \8539 , \8292 );
and \U$8408 ( \8540 , \8538 , \8539 );
and \U$8409 ( \8541 , \166 , \8540 );
and \U$8410 ( \8542 , \150 , \8292 );
nor \U$8411 ( \8543 , \8541 , \8542 );
xnor \U$8412 ( \8544 , \8543 , \8297 );
xor \U$8413 ( \8545 , \8537 , \8544 );
and \U$8414 ( \8546 , \8407 , \8411 );
and \U$8415 ( \8547 , \8411 , \8416 );
and \U$8416 ( \8548 , \8407 , \8416 );
or \U$8417 ( \8549 , \8546 , \8547 , \8548 );
and \U$8418 ( \8550 , \8391 , \8395 );
and \U$8419 ( \8551 , \8395 , \8400 );
and \U$8420 ( \8552 , \8391 , \8400 );
or \U$8421 ( \8553 , \8550 , \8551 , \8552 );
xor \U$8422 ( \8554 , \8549 , \8553 );
and \U$8423 ( \8555 , \8421 , \8425 );
and \U$8424 ( \8556 , \8425 , \8430 );
and \U$8425 ( \8557 , \8421 , \8430 );
or \U$8426 ( \8558 , \8555 , \8556 , \8557 );
xor \U$8427 ( \8559 , \8554 , \8558 );
xor \U$8428 ( \8560 , \8545 , \8559 );
and \U$8429 ( \8561 , \8271 , \8275 );
and \U$8430 ( \8562 , \8275 , \8280 );
and \U$8431 ( \8563 , \8271 , \8280 );
or \U$8432 ( \8564 , \8561 , \8562 , \8563 );
and \U$8433 ( \8565 , \8304 , \8308 );
and \U$8434 ( \8566 , \8308 , \8313 );
and \U$8435 ( \8567 , \8304 , \8313 );
or \U$8436 ( \8568 , \8565 , \8566 , \8567 );
xor \U$8437 ( \8569 , \8564 , \8568 );
and \U$8438 ( \8570 , \8436 , \8440 );
and \U$8439 ( \8571 , \8440 , \8445 );
and \U$8440 ( \8572 , \8436 , \8445 );
or \U$8441 ( \8573 , \8570 , \8571 , \8572 );
xor \U$8442 ( \8574 , \8569 , \8573 );
xor \U$8443 ( \8575 , \8560 , \8574 );
xor \U$8444 ( \8576 , \8528 , \8575 );
xor \U$8445 ( \8577 , \8509 , \8576 );
and \U$8446 ( \8578 , \8372 , \8386 );
and \U$8447 ( \8579 , \8386 , \8401 );
and \U$8448 ( \8580 , \8372 , \8401 );
or \U$8449 ( \8581 , \8578 , \8579 , \8580 );
and \U$8450 ( \8582 , \8417 , \8431 );
and \U$8451 ( \8583 , \8431 , \8446 );
and \U$8452 ( \8584 , \8417 , \8446 );
or \U$8453 ( \8585 , \8582 , \8583 , \8584 );
xor \U$8454 ( \8586 , \8581 , \8585 );
and \U$8455 ( \8587 , \8281 , \8299 );
and \U$8456 ( \8588 , \8299 , \8314 );
and \U$8457 ( \8589 , \8281 , \8314 );
or \U$8458 ( \8590 , \8587 , \8588 , \8589 );
xor \U$8459 ( \8591 , \8586 , \8590 );
and \U$8460 ( \8592 , \8242 , \8246 );
and \U$8461 ( \8593 , \8246 , \8251 );
and \U$8462 ( \8594 , \8242 , \8251 );
or \U$8463 ( \8595 , \8592 , \8593 , \8594 );
and \U$8464 ( \8596 , \8256 , \8260 );
and \U$8465 ( \8597 , \8260 , \8265 );
and \U$8466 ( \8598 , \8256 , \8265 );
or \U$8467 ( \8599 , \8596 , \8597 , \8598 );
xor \U$8468 ( \8600 , \8595 , \8599 );
and \U$8469 ( \8601 , \8227 , \8231 );
and \U$8470 ( \8602 , \8231 , \8236 );
and \U$8471 ( \8603 , \8227 , \8236 );
or \U$8472 ( \8604 , \8601 , \8602 , \8603 );
xor \U$8473 ( \8605 , \8600 , \8604 );
xor \U$8474 ( \8606 , \8591 , \8605 );
and \U$8475 ( \8607 , \185 , \5011 );
and \U$8476 ( \8608 , \261 , \4878 );
nor \U$8477 ( \8609 , \8607 , \8608 );
xnor \U$8478 ( \8610 , \8609 , \4762 );
and \U$8479 ( \8611 , \197 , \5485 );
and \U$8480 ( \8612 , \178 , \5275 );
nor \U$8481 ( \8613 , \8611 , \8612 );
xnor \U$8482 ( \8614 , \8613 , \5169 );
xor \U$8483 ( \8615 , \8610 , \8614 );
and \U$8484 ( \8616 , \217 , \5996 );
and \U$8485 ( \8617 , \189 , \5695 );
nor \U$8486 ( \8618 , \8616 , \8617 );
xnor \U$8487 ( \8619 , \8618 , \5687 );
xor \U$8488 ( \8620 , \8615 , \8619 );
and \U$8489 ( \8621 , \232 , \6401 );
and \U$8490 ( \8622 , \209 , \6143 );
nor \U$8491 ( \8623 , \8621 , \8622 );
xnor \U$8492 ( \8624 , \8623 , \6148 );
and \U$8493 ( \8625 , \247 , \7055 );
and \U$8494 ( \8626 , \224 , \6675 );
nor \U$8495 ( \8627 , \8625 , \8626 );
xnor \U$8496 ( \8628 , \8627 , \6680 );
xor \U$8497 ( \8629 , \8624 , \8628 );
and \U$8498 ( \8630 , \143 , \7489 );
and \U$8499 ( \8631 , \240 , \7137 );
nor \U$8500 ( \8632 , \8630 , \8631 );
xnor \U$8501 ( \8633 , \8632 , \7142 );
xor \U$8502 ( \8634 , \8629 , \8633 );
xor \U$8503 ( \8635 , \8620 , \8634 );
and \U$8504 ( \8636 , \1192 , \3813 );
and \U$8505 ( \8637 , \1333 , \3557 );
nor \U$8506 ( \8638 , \8636 , \8637 );
xnor \U$8507 ( \8639 , \8638 , \3562 );
and \U$8508 ( \8640 , \474 , \4132 );
and \U$8509 ( \8641 , \1147 , \4012 );
nor \U$8510 ( \8642 , \8640 , \8641 );
xnor \U$8511 ( \8643 , \8642 , \3925 );
xor \U$8512 ( \8644 , \8639 , \8643 );
and \U$8513 ( \8645 , \307 , \4581 );
and \U$8514 ( \8646 , \412 , \4424 );
nor \U$8515 ( \8647 , \8645 , \8646 );
xnor \U$8516 ( \8648 , \8647 , \4377 );
xor \U$8517 ( \8649 , \8644 , \8648 );
xor \U$8518 ( \8650 , \8635 , \8649 );
and \U$8519 ( \8651 , \8349 , \183 );
buf \U$8520 ( \8652 , RIb55eef0_71);
and \U$8521 ( \8653 , \8652 , \180 );
nor \U$8522 ( \8654 , \8651 , \8653 );
xnor \U$8523 ( \8655 , \8654 , \179 );
and \U$8524 ( \8656 , \7700 , \195 );
and \U$8525 ( \8657 , \8057 , \193 );
nor \U$8526 ( \8658 , \8656 , \8657 );
xnor \U$8527 ( \8659 , \8658 , \202 );
xor \U$8528 ( \8660 , \8655 , \8659 );
and \U$8529 ( \8661 , \7231 , \215 );
and \U$8530 ( \8662 , \7556 , \213 );
nor \U$8531 ( \8663 , \8661 , \8662 );
xnor \U$8532 ( \8664 , \8663 , \222 );
xor \U$8533 ( \8665 , \8660 , \8664 );
and \U$8534 ( \8666 , \6790 , \230 );
and \U$8535 ( \8667 , \6945 , \228 );
nor \U$8536 ( \8668 , \8666 , \8667 );
xnor \U$8537 ( \8669 , \8668 , \237 );
and \U$8538 ( \8670 , \6281 , \245 );
and \U$8539 ( \8671 , \6514 , \243 );
nor \U$8540 ( \8672 , \8670 , \8671 );
xnor \U$8541 ( \8673 , \8672 , \252 );
xor \U$8542 ( \8674 , \8669 , \8673 );
and \U$8543 ( \8675 , \5674 , \141 );
and \U$8544 ( \8676 , \6030 , \139 );
nor \U$8545 ( \8677 , \8675 , \8676 );
xnor \U$8546 ( \8678 , \8677 , \148 );
xor \U$8547 ( \8679 , \8674 , \8678 );
xor \U$8548 ( \8680 , \8665 , \8679 );
and \U$8549 ( \8681 , \5156 , \156 );
and \U$8550 ( \8682 , \5469 , \154 );
nor \U$8551 ( \8683 , \8681 , \8682 );
xnor \U$8552 ( \8684 , \8683 , \163 );
and \U$8553 ( \8685 , \4749 , \296 );
and \U$8554 ( \8686 , \4922 , \168 );
nor \U$8555 ( \8687 , \8685 , \8686 );
xnor \U$8556 ( \8688 , \8687 , \173 );
xor \U$8557 ( \8689 , \8684 , \8688 );
and \U$8558 ( \8690 , \4364 , \438 );
and \U$8559 ( \8691 , \4654 , \336 );
nor \U$8560 ( \8692 , \8690 , \8691 );
xnor \U$8561 ( \8693 , \8692 , \320 );
xor \U$8562 ( \8694 , \8689 , \8693 );
xor \U$8563 ( \8695 , \8680 , \8694 );
xor \U$8564 ( \8696 , \8650 , \8695 );
and \U$8565 ( \8697 , \2826 , \1824 );
and \U$8566 ( \8698 , \3037 , \1739 );
nor \U$8567 ( \8699 , \8697 , \8698 );
xnor \U$8568 ( \8700 , \8699 , \1697 );
and \U$8569 ( \8701 , \2521 , \2121 );
and \U$8570 ( \8702 , \2757 , \2008 );
nor \U$8571 ( \8703 , \8701 , \8702 );
xnor \U$8572 ( \8704 , \8703 , \1961 );
xor \U$8573 ( \8705 , \8700 , \8704 );
and \U$8574 ( \8706 , \2182 , \2400 );
and \U$8575 ( \8707 , \2366 , \2246 );
nor \U$8576 ( \8708 , \8706 , \8707 );
xnor \U$8577 ( \8709 , \8708 , \2195 );
xor \U$8578 ( \8710 , \8705 , \8709 );
and \U$8579 ( \8711 , \1948 , \2669 );
and \U$8580 ( \8712 , \2090 , \2538 );
nor \U$8581 ( \8713 , \8711 , \8712 );
xnor \U$8582 ( \8714 , \8713 , \2534 );
and \U$8583 ( \8715 , \1684 , \3103 );
and \U$8584 ( \8716 , \1802 , \2934 );
nor \U$8585 ( \8717 , \8715 , \8716 );
xnor \U$8586 ( \8718 , \8717 , \2839 );
xor \U$8587 ( \8719 , \8714 , \8718 );
and \U$8588 ( \8720 , \1484 , \3357 );
and \U$8589 ( \8721 , \1601 , \3255 );
nor \U$8590 ( \8722 , \8720 , \8721 );
xnor \U$8591 ( \8723 , \8722 , \3156 );
xor \U$8592 ( \8724 , \8719 , \8723 );
xor \U$8593 ( \8725 , \8710 , \8724 );
and \U$8594 ( \8726 , \3912 , \1086 );
and \U$8595 ( \8727 , \4160 , \508 );
nor \U$8596 ( \8728 , \8726 , \8727 );
xnor \U$8597 ( \8729 , \8728 , \487 );
and \U$8598 ( \8730 , \3646 , \1301 );
and \U$8599 ( \8731 , \3736 , \1246 );
nor \U$8600 ( \8732 , \8730 , \8731 );
xnor \U$8601 ( \8733 , \8732 , \1205 );
xor \U$8602 ( \8734 , \8729 , \8733 );
and \U$8603 ( \8735 , \3143 , \1578 );
and \U$8604 ( \8736 , \3395 , \1431 );
nor \U$8605 ( \8737 , \8735 , \8736 );
xnor \U$8606 ( \8738 , \8737 , \1436 );
xor \U$8607 ( \8739 , \8734 , \8738 );
xor \U$8608 ( \8740 , \8725 , \8739 );
xor \U$8609 ( \8741 , \8696 , \8740 );
xor \U$8610 ( \8742 , \8606 , \8741 );
xor \U$8611 ( \8743 , \8577 , \8742 );
xor \U$8612 ( \8744 , \8495 , \8743 );
xor \U$8613 ( \8745 , \8486 , \8744 );
xor \U$8614 ( \8746 , \8467 , \8745 );
and \U$8615 ( \8747 , \8196 , \8451 );
xor \U$8616 ( \8748 , \8746 , \8747 );
and \U$8617 ( \8749 , \8452 , \8456 );
and \U$8618 ( \8750 , \8457 , \8460 );
or \U$8619 ( \8751 , \8749 , \8750 );
xor \U$8620 ( \8752 , \8748 , \8751 );
buf \U$8621 ( \8753 , \8752 );
buf \U$8622 ( \8754 , \8753 );
and \U$8623 ( \8755 , \8471 , \8485 );
and \U$8624 ( \8756 , \8485 , \8744 );
and \U$8625 ( \8757 , \8471 , \8744 );
or \U$8626 ( \8758 , \8755 , \8756 , \8757 );
and \U$8627 ( \8759 , \8490 , \8494 );
and \U$8628 ( \8760 , \8494 , \8743 );
and \U$8629 ( \8761 , \8490 , \8743 );
or \U$8630 ( \8762 , \8759 , \8760 , \8761 );
and \U$8631 ( \8763 , \8499 , \8503 );
and \U$8632 ( \8764 , \8503 , \8508 );
and \U$8633 ( \8765 , \8499 , \8508 );
or \U$8634 ( \8766 , \8763 , \8764 , \8765 );
and \U$8635 ( \8767 , \8513 , \8527 );
and \U$8636 ( \8768 , \8527 , \8575 );
and \U$8637 ( \8769 , \8513 , \8575 );
or \U$8638 ( \8770 , \8767 , \8768 , \8769 );
xor \U$8639 ( \8771 , \8766 , \8770 );
and \U$8640 ( \8772 , \8591 , \8605 );
and \U$8641 ( \8773 , \8605 , \8741 );
and \U$8642 ( \8774 , \8591 , \8741 );
or \U$8643 ( \8775 , \8772 , \8773 , \8774 );
xor \U$8644 ( \8776 , \8771 , \8775 );
xor \U$8645 ( \8777 , \8762 , \8776 );
and \U$8646 ( \8778 , \8475 , \8479 );
and \U$8647 ( \8779 , \8479 , \8484 );
and \U$8648 ( \8780 , \8475 , \8484 );
or \U$8649 ( \8781 , \8778 , \8779 , \8780 );
and \U$8650 ( \8782 , \8509 , \8576 );
and \U$8651 ( \8783 , \8576 , \8742 );
and \U$8652 ( \8784 , \8509 , \8742 );
or \U$8653 ( \8785 , \8782 , \8783 , \8784 );
xor \U$8654 ( \8786 , \8781 , \8785 );
and \U$8655 ( \8787 , \8581 , \8585 );
and \U$8656 ( \8788 , \8585 , \8590 );
and \U$8657 ( \8789 , \8581 , \8590 );
or \U$8658 ( \8790 , \8787 , \8788 , \8789 );
and \U$8659 ( \8791 , \8595 , \8599 );
and \U$8660 ( \8792 , \8599 , \8604 );
and \U$8661 ( \8793 , \8595 , \8604 );
or \U$8662 ( \8794 , \8791 , \8792 , \8793 );
xor \U$8663 ( \8795 , \8790 , \8794 );
and \U$8664 ( \8796 , \8650 , \8695 );
and \U$8665 ( \8797 , \8695 , \8740 );
and \U$8666 ( \8798 , \8650 , \8740 );
or \U$8667 ( \8799 , \8796 , \8797 , \8798 );
xor \U$8668 ( \8800 , \8795 , \8799 );
and \U$8669 ( \8801 , \8532 , \8536 );
and \U$8670 ( \8802 , \8536 , \8544 );
and \U$8671 ( \8803 , \8532 , \8544 );
or \U$8672 ( \8804 , \8801 , \8802 , \8803 );
and \U$8673 ( \8805 , \8620 , \8634 );
and \U$8674 ( \8806 , \8634 , \8649 );
and \U$8675 ( \8807 , \8620 , \8649 );
or \U$8676 ( \8808 , \8805 , \8806 , \8807 );
xor \U$8677 ( \8809 , \8804 , \8808 );
and \U$8678 ( \8810 , \8710 , \8724 );
and \U$8679 ( \8811 , \8724 , \8739 );
and \U$8680 ( \8812 , \8710 , \8739 );
or \U$8681 ( \8813 , \8810 , \8811 , \8812 );
xor \U$8682 ( \8814 , \8809 , \8813 );
and \U$8683 ( \8815 , \8517 , \8521 );
and \U$8684 ( \8816 , \8521 , \8526 );
and \U$8685 ( \8817 , \8517 , \8526 );
or \U$8686 ( \8818 , \8815 , \8816 , \8817 );
and \U$8687 ( \8819 , \8549 , \8553 );
and \U$8688 ( \8820 , \8553 , \8558 );
and \U$8689 ( \8821 , \8549 , \8558 );
or \U$8690 ( \8822 , \8819 , \8820 , \8821 );
xor \U$8691 ( \8823 , \8818 , \8822 );
and \U$8692 ( \8824 , \8564 , \8568 );
and \U$8693 ( \8825 , \8568 , \8573 );
and \U$8694 ( \8826 , \8564 , \8573 );
or \U$8695 ( \8827 , \8824 , \8825 , \8826 );
xor \U$8696 ( \8828 , \8823 , \8827 );
xor \U$8697 ( \8829 , \8814 , \8828 );
and \U$8698 ( \8830 , \8665 , \8679 );
and \U$8699 ( \8831 , \8679 , \8694 );
and \U$8700 ( \8832 , \8665 , \8694 );
or \U$8701 ( \8833 , \8830 , \8831 , \8832 );
and \U$8702 ( \8834 , \8652 , \183 );
buf \U$8703 ( \8835 , RIb55ef68_70);
and \U$8704 ( \8836 , \8835 , \180 );
nor \U$8705 ( \8837 , \8834 , \8836 );
xnor \U$8706 ( \8838 , \8837 , \179 );
and \U$8707 ( \8839 , \8057 , \195 );
and \U$8708 ( \8840 , \8349 , \193 );
nor \U$8709 ( \8841 , \8839 , \8840 );
xnor \U$8710 ( \8842 , \8841 , \202 );
xor \U$8711 ( \8843 , \8838 , \8842 );
buf \U$8712 ( \8844 , RIb560de0_5);
buf \U$8713 ( \8845 , RIb560d68_6);
and \U$8714 ( \8846 , \8845 , \8294 );
not \U$8715 ( \8847 , \8846 );
and \U$8716 ( \8848 , \8844 , \8847 );
xor \U$8717 ( \8849 , \8843 , \8848 );
xor \U$8718 ( \8850 , \8833 , \8849 );
and \U$8719 ( \8851 , \7556 , \215 );
and \U$8720 ( \8852 , \7700 , \213 );
nor \U$8721 ( \8853 , \8851 , \8852 );
xnor \U$8722 ( \8854 , \8853 , \222 );
and \U$8723 ( \8855 , \6945 , \230 );
and \U$8724 ( \8856 , \7231 , \228 );
nor \U$8725 ( \8857 , \8855 , \8856 );
xnor \U$8726 ( \8858 , \8857 , \237 );
xor \U$8727 ( \8859 , \8854 , \8858 );
and \U$8728 ( \8860 , \6514 , \245 );
and \U$8729 ( \8861 , \6790 , \243 );
nor \U$8730 ( \8862 , \8860 , \8861 );
xnor \U$8731 ( \8863 , \8862 , \252 );
xor \U$8732 ( \8864 , \8859 , \8863 );
xor \U$8733 ( \8865 , \8850 , \8864 );
xor \U$8734 ( \8866 , \8829 , \8865 );
xor \U$8735 ( \8867 , \8800 , \8866 );
and \U$8736 ( \8868 , \8545 , \8559 );
and \U$8737 ( \8869 , \8559 , \8574 );
and \U$8738 ( \8870 , \8545 , \8574 );
or \U$8739 ( \8871 , \8868 , \8869 , \8870 );
and \U$8740 ( \8872 , \8700 , \8704 );
and \U$8741 ( \8873 , \8704 , \8709 );
and \U$8742 ( \8874 , \8700 , \8709 );
or \U$8743 ( \8875 , \8872 , \8873 , \8874 );
and \U$8744 ( \8876 , \8714 , \8718 );
and \U$8745 ( \8877 , \8718 , \8723 );
and \U$8746 ( \8878 , \8714 , \8723 );
or \U$8747 ( \8879 , \8876 , \8877 , \8878 );
xor \U$8748 ( \8880 , \8875 , \8879 );
and \U$8749 ( \8881 , \8729 , \8733 );
and \U$8750 ( \8882 , \8733 , \8738 );
and \U$8751 ( \8883 , \8729 , \8738 );
or \U$8752 ( \8884 , \8881 , \8882 , \8883 );
xor \U$8753 ( \8885 , \8880 , \8884 );
and \U$8754 ( \8886 , \8610 , \8614 );
and \U$8755 ( \8887 , \8614 , \8619 );
and \U$8756 ( \8888 , \8610 , \8619 );
or \U$8757 ( \8889 , \8886 , \8887 , \8888 );
and \U$8758 ( \8890 , \8624 , \8628 );
and \U$8759 ( \8891 , \8628 , \8633 );
and \U$8760 ( \8892 , \8624 , \8633 );
or \U$8761 ( \8893 , \8890 , \8891 , \8892 );
xor \U$8762 ( \8894 , \8889 , \8893 );
and \U$8763 ( \8895 , \8639 , \8643 );
and \U$8764 ( \8896 , \8643 , \8648 );
and \U$8765 ( \8897 , \8639 , \8648 );
or \U$8766 ( \8898 , \8895 , \8896 , \8897 );
xor \U$8767 ( \8899 , \8894 , \8898 );
xor \U$8768 ( \8900 , \8885 , \8899 );
and \U$8769 ( \8901 , \8655 , \8659 );
and \U$8770 ( \8902 , \8659 , \8664 );
and \U$8771 ( \8903 , \8655 , \8664 );
or \U$8772 ( \8904 , \8901 , \8902 , \8903 );
and \U$8773 ( \8905 , \8669 , \8673 );
and \U$8774 ( \8906 , \8673 , \8678 );
and \U$8775 ( \8907 , \8669 , \8678 );
or \U$8776 ( \8908 , \8905 , \8906 , \8907 );
xor \U$8777 ( \8909 , \8904 , \8908 );
and \U$8778 ( \8910 , \8684 , \8688 );
and \U$8779 ( \8911 , \8688 , \8693 );
and \U$8780 ( \8912 , \8684 , \8693 );
or \U$8781 ( \8913 , \8910 , \8911 , \8912 );
xor \U$8782 ( \8914 , \8909 , \8913 );
xor \U$8783 ( \8915 , \8900 , \8914 );
xor \U$8784 ( \8916 , \8871 , \8915 );
and \U$8785 ( \8917 , \6030 , \141 );
and \U$8786 ( \8918 , \6281 , \139 );
nor \U$8787 ( \8919 , \8917 , \8918 );
xnor \U$8788 ( \8920 , \8919 , \148 );
and \U$8789 ( \8921 , \5469 , \156 );
and \U$8790 ( \8922 , \5674 , \154 );
nor \U$8791 ( \8923 , \8921 , \8922 );
xnor \U$8792 ( \8924 , \8923 , \163 );
xor \U$8793 ( \8925 , \8920 , \8924 );
and \U$8794 ( \8926 , \4922 , \296 );
and \U$8795 ( \8927 , \5156 , \168 );
nor \U$8796 ( \8928 , \8926 , \8927 );
xnor \U$8797 ( \8929 , \8928 , \173 );
xor \U$8798 ( \8930 , \8925 , \8929 );
and \U$8799 ( \8931 , \3395 , \1578 );
and \U$8800 ( \8932 , \3646 , \1431 );
nor \U$8801 ( \8933 , \8931 , \8932 );
xnor \U$8802 ( \8934 , \8933 , \1436 );
and \U$8803 ( \8935 , \3037 , \1824 );
and \U$8804 ( \8936 , \3143 , \1739 );
nor \U$8805 ( \8937 , \8935 , \8936 );
xnor \U$8806 ( \8938 , \8937 , \1697 );
xor \U$8807 ( \8939 , \8934 , \8938 );
and \U$8808 ( \8940 , \2757 , \2121 );
and \U$8809 ( \8941 , \2826 , \2008 );
nor \U$8810 ( \8942 , \8940 , \8941 );
xnor \U$8811 ( \8943 , \8942 , \1961 );
xor \U$8812 ( \8944 , \8939 , \8943 );
xor \U$8813 ( \8945 , \8930 , \8944 );
and \U$8814 ( \8946 , \4654 , \438 );
and \U$8815 ( \8947 , \4749 , \336 );
nor \U$8816 ( \8948 , \8946 , \8947 );
xnor \U$8817 ( \8949 , \8948 , \320 );
and \U$8818 ( \8950 , \4160 , \1086 );
and \U$8819 ( \8951 , \4364 , \508 );
nor \U$8820 ( \8952 , \8950 , \8951 );
xnor \U$8821 ( \8953 , \8952 , \487 );
xor \U$8822 ( \8954 , \8949 , \8953 );
and \U$8823 ( \8955 , \3736 , \1301 );
and \U$8824 ( \8956 , \3912 , \1246 );
nor \U$8825 ( \8957 , \8955 , \8956 );
xnor \U$8826 ( \8958 , \8957 , \1205 );
xor \U$8827 ( \8959 , \8954 , \8958 );
xor \U$8828 ( \8960 , \8945 , \8959 );
and \U$8829 ( \8961 , \2366 , \2400 );
and \U$8830 ( \8962 , \2521 , \2246 );
nor \U$8831 ( \8963 , \8961 , \8962 );
xnor \U$8832 ( \8964 , \8963 , \2195 );
and \U$8833 ( \8965 , \2090 , \2669 );
and \U$8834 ( \8966 , \2182 , \2538 );
nor \U$8835 ( \8967 , \8965 , \8966 );
xnor \U$8836 ( \8968 , \8967 , \2534 );
xor \U$8837 ( \8969 , \8964 , \8968 );
and \U$8838 ( \8970 , \1802 , \3103 );
and \U$8839 ( \8971 , \1948 , \2934 );
nor \U$8840 ( \8972 , \8970 , \8971 );
xnor \U$8841 ( \8973 , \8972 , \2839 );
xor \U$8842 ( \8974 , \8969 , \8973 );
and \U$8843 ( \8975 , \1601 , \3357 );
and \U$8844 ( \8976 , \1684 , \3255 );
nor \U$8845 ( \8977 , \8975 , \8976 );
xnor \U$8846 ( \8978 , \8977 , \3156 );
and \U$8847 ( \8979 , \1333 , \3813 );
and \U$8848 ( \8980 , \1484 , \3557 );
nor \U$8849 ( \8981 , \8979 , \8980 );
xnor \U$8850 ( \8982 , \8981 , \3562 );
xor \U$8851 ( \8983 , \8978 , \8982 );
and \U$8852 ( \8984 , \1147 , \4132 );
and \U$8853 ( \8985 , \1192 , \4012 );
nor \U$8854 ( \8986 , \8984 , \8985 );
xnor \U$8855 ( \8987 , \8986 , \3925 );
xor \U$8856 ( \8988 , \8983 , \8987 );
xor \U$8857 ( \8989 , \8974 , \8988 );
and \U$8858 ( \8990 , \412 , \4581 );
and \U$8859 ( \8991 , \474 , \4424 );
nor \U$8860 ( \8992 , \8990 , \8991 );
xnor \U$8861 ( \8993 , \8992 , \4377 );
and \U$8862 ( \8994 , \261 , \5011 );
and \U$8863 ( \8995 , \307 , \4878 );
nor \U$8864 ( \8996 , \8994 , \8995 );
xnor \U$8865 ( \8997 , \8996 , \4762 );
xor \U$8866 ( \8998 , \8993 , \8997 );
and \U$8867 ( \8999 , \178 , \5485 );
and \U$8868 ( \9000 , \185 , \5275 );
nor \U$8869 ( \9001 , \8999 , \9000 );
xnor \U$8870 ( \9002 , \9001 , \5169 );
xor \U$8871 ( \9003 , \8998 , \9002 );
xor \U$8872 ( \9004 , \8989 , \9003 );
xor \U$8873 ( \9005 , \8960 , \9004 );
xor \U$8874 ( \9006 , \8845 , \8294 );
nand \U$8875 ( \9007 , \166 , \9006 );
xnor \U$8876 ( \9008 , \9007 , \8848 );
and \U$8877 ( \9009 , \189 , \5996 );
and \U$8878 ( \9010 , \197 , \5695 );
nor \U$8879 ( \9011 , \9009 , \9010 );
xnor \U$8880 ( \9012 , \9011 , \5687 );
and \U$8881 ( \9013 , \209 , \6401 );
and \U$8882 ( \9014 , \217 , \6143 );
nor \U$8883 ( \9015 , \9013 , \9014 );
xnor \U$8884 ( \9016 , \9015 , \6148 );
xor \U$8885 ( \9017 , \9012 , \9016 );
and \U$8886 ( \9018 , \224 , \7055 );
and \U$8887 ( \9019 , \232 , \6675 );
nor \U$8888 ( \9020 , \9018 , \9019 );
xnor \U$8889 ( \9021 , \9020 , \6680 );
xor \U$8890 ( \9022 , \9017 , \9021 );
xor \U$8891 ( \9023 , \9008 , \9022 );
and \U$8892 ( \9024 , \240 , \7489 );
and \U$8893 ( \9025 , \247 , \7137 );
nor \U$8894 ( \9026 , \9024 , \9025 );
xnor \U$8895 ( \9027 , \9026 , \7142 );
and \U$8896 ( \9028 , \134 , \8019 );
and \U$8897 ( \9029 , \143 , \7830 );
nor \U$8898 ( \9030 , \9028 , \9029 );
xnor \U$8899 ( \9031 , \9030 , \7713 );
xor \U$8900 ( \9032 , \9027 , \9031 );
and \U$8901 ( \9033 , \150 , \8540 );
and \U$8902 ( \9034 , \158 , \8292 );
nor \U$8903 ( \9035 , \9033 , \9034 );
xnor \U$8904 ( \9036 , \9035 , \8297 );
xor \U$8905 ( \9037 , \9032 , \9036 );
xor \U$8906 ( \9038 , \9023 , \9037 );
xor \U$8907 ( \9039 , \9005 , \9038 );
xor \U$8908 ( \9040 , \8916 , \9039 );
xor \U$8909 ( \9041 , \8867 , \9040 );
xor \U$8910 ( \9042 , \8786 , \9041 );
xor \U$8911 ( \9043 , \8777 , \9042 );
xor \U$8912 ( \9044 , \8758 , \9043 );
and \U$8913 ( \9045 , \8467 , \8745 );
xor \U$8914 ( \9046 , \9044 , \9045 );
and \U$8915 ( \9047 , \8746 , \8747 );
and \U$8916 ( \9048 , \8748 , \8751 );
or \U$8917 ( \9049 , \9047 , \9048 );
xor \U$8918 ( \9050 , \9046 , \9049 );
buf \U$8919 ( \9051 , \9050 );
buf \U$8920 ( \9052 , \9051 );
and \U$8921 ( \9053 , \8762 , \8776 );
and \U$8922 ( \9054 , \8776 , \9042 );
and \U$8923 ( \9055 , \8762 , \9042 );
or \U$8924 ( \9056 , \9053 , \9054 , \9055 );
and \U$8925 ( \9057 , \8781 , \8785 );
and \U$8926 ( \9058 , \8785 , \9041 );
and \U$8927 ( \9059 , \8781 , \9041 );
or \U$8928 ( \9060 , \9057 , \9058 , \9059 );
and \U$8929 ( \9061 , \8766 , \8770 );
and \U$8930 ( \9062 , \8770 , \8775 );
and \U$8931 ( \9063 , \8766 , \8775 );
or \U$8932 ( \9064 , \9061 , \9062 , \9063 );
and \U$8933 ( \9065 , \8800 , \8866 );
and \U$8934 ( \9066 , \8866 , \9040 );
and \U$8935 ( \9067 , \8800 , \9040 );
or \U$8936 ( \9068 , \9065 , \9066 , \9067 );
xor \U$8937 ( \9069 , \9064 , \9068 );
and \U$8938 ( \9070 , \8885 , \8899 );
and \U$8939 ( \9071 , \8899 , \8914 );
and \U$8940 ( \9072 , \8885 , \8914 );
or \U$8941 ( \9073 , \9070 , \9071 , \9072 );
and \U$8942 ( \9074 , \8960 , \9004 );
and \U$8943 ( \9075 , \9004 , \9038 );
and \U$8944 ( \9076 , \8960 , \9038 );
or \U$8945 ( \9077 , \9074 , \9075 , \9076 );
xor \U$8946 ( \9078 , \9073 , \9077 );
and \U$8947 ( \9079 , \8964 , \8968 );
and \U$8948 ( \9080 , \8968 , \8973 );
and \U$8949 ( \9081 , \8964 , \8973 );
or \U$8950 ( \9082 , \9079 , \9080 , \9081 );
and \U$8951 ( \9083 , \8934 , \8938 );
and \U$8952 ( \9084 , \8938 , \8943 );
and \U$8953 ( \9085 , \8934 , \8943 );
or \U$8954 ( \9086 , \9083 , \9084 , \9085 );
xor \U$8955 ( \9087 , \9082 , \9086 );
and \U$8956 ( \9088 , \8949 , \8953 );
and \U$8957 ( \9089 , \8953 , \8958 );
and \U$8958 ( \9090 , \8949 , \8958 );
or \U$8959 ( \9091 , \9088 , \9089 , \9090 );
xor \U$8960 ( \9092 , \9087 , \9091 );
xor \U$8961 ( \9093 , \9078 , \9092 );
xor \U$8962 ( \9094 , \9069 , \9093 );
xor \U$8963 ( \9095 , \9060 , \9094 );
and \U$8964 ( \9096 , \8804 , \8808 );
and \U$8965 ( \9097 , \8808 , \8813 );
and \U$8966 ( \9098 , \8804 , \8813 );
or \U$8967 ( \9099 , \9096 , \9097 , \9098 );
and \U$8968 ( \9100 , \8818 , \8822 );
and \U$8969 ( \9101 , \8822 , \8827 );
and \U$8970 ( \9102 , \8818 , \8827 );
or \U$8971 ( \9103 , \9100 , \9101 , \9102 );
xor \U$8972 ( \9104 , \9099 , \9103 );
and \U$8973 ( \9105 , \8833 , \8849 );
and \U$8974 ( \9106 , \8849 , \8864 );
and \U$8975 ( \9107 , \8833 , \8864 );
or \U$8976 ( \9108 , \9105 , \9106 , \9107 );
xor \U$8977 ( \9109 , \9104 , \9108 );
and \U$8978 ( \9110 , \8790 , \8794 );
and \U$8979 ( \9111 , \8794 , \8799 );
and \U$8980 ( \9112 , \8790 , \8799 );
or \U$8981 ( \9113 , \9110 , \9111 , \9112 );
and \U$8982 ( \9114 , \8814 , \8828 );
and \U$8983 ( \9115 , \8828 , \8865 );
and \U$8984 ( \9116 , \8814 , \8865 );
or \U$8985 ( \9117 , \9114 , \9115 , \9116 );
xor \U$8986 ( \9118 , \9113 , \9117 );
and \U$8987 ( \9119 , \8871 , \8915 );
and \U$8988 ( \9120 , \8915 , \9039 );
and \U$8989 ( \9121 , \8871 , \9039 );
or \U$8990 ( \9122 , \9119 , \9120 , \9121 );
xor \U$8991 ( \9123 , \9118 , \9122 );
xor \U$8992 ( \9124 , \9109 , \9123 );
and \U$8993 ( \9125 , \8875 , \8879 );
and \U$8994 ( \9126 , \8879 , \8884 );
and \U$8995 ( \9127 , \8875 , \8884 );
or \U$8996 ( \9128 , \9125 , \9126 , \9127 );
and \U$8997 ( \9129 , \8889 , \8893 );
and \U$8998 ( \9130 , \8893 , \8898 );
and \U$8999 ( \9131 , \8889 , \8898 );
or \U$9000 ( \9132 , \9129 , \9130 , \9131 );
xor \U$9001 ( \9133 , \9128 , \9132 );
and \U$9002 ( \9134 , \8904 , \8908 );
and \U$9003 ( \9135 , \8908 , \8913 );
and \U$9004 ( \9136 , \8904 , \8913 );
or \U$9005 ( \9137 , \9134 , \9135 , \9136 );
xor \U$9006 ( \9138 , \9133 , \9137 );
and \U$9007 ( \9139 , \8930 , \8944 );
and \U$9008 ( \9140 , \8944 , \8959 );
and \U$9009 ( \9141 , \8930 , \8959 );
or \U$9010 ( \9142 , \9139 , \9140 , \9141 );
and \U$9011 ( \9143 , \8974 , \8988 );
and \U$9012 ( \9144 , \8988 , \9003 );
and \U$9013 ( \9145 , \8974 , \9003 );
or \U$9014 ( \9146 , \9143 , \9144 , \9145 );
xor \U$9015 ( \9147 , \9142 , \9146 );
and \U$9016 ( \9148 , \9008 , \9022 );
and \U$9017 ( \9149 , \9022 , \9037 );
and \U$9018 ( \9150 , \9008 , \9037 );
or \U$9019 ( \9151 , \9148 , \9149 , \9150 );
xor \U$9020 ( \9152 , \9147 , \9151 );
xor \U$9021 ( \9153 , \9138 , \9152 );
and \U$9022 ( \9154 , \8920 , \8924 );
and \U$9023 ( \9155 , \8924 , \8929 );
and \U$9024 ( \9156 , \8920 , \8929 );
or \U$9025 ( \9157 , \9154 , \9155 , \9156 );
and \U$9026 ( \9158 , \8838 , \8842 );
and \U$9027 ( \9159 , \8842 , \8848 );
and \U$9028 ( \9160 , \8838 , \8848 );
or \U$9029 ( \9161 , \9158 , \9159 , \9160 );
xor \U$9030 ( \9162 , \9157 , \9161 );
and \U$9031 ( \9163 , \8854 , \8858 );
and \U$9032 ( \9164 , \8858 , \8863 );
and \U$9033 ( \9165 , \8854 , \8863 );
or \U$9034 ( \9166 , \9163 , \9164 , \9165 );
xor \U$9035 ( \9167 , \9162 , \9166 );
and \U$9036 ( \9168 , \8835 , \183 );
buf \U$9037 ( \9169 , RIb55efe0_69);
and \U$9038 ( \9170 , \9169 , \180 );
nor \U$9039 ( \9171 , \9168 , \9170 );
xnor \U$9040 ( \9172 , \9171 , \179 );
and \U$9041 ( \9173 , \8349 , \195 );
and \U$9042 ( \9174 , \8652 , \193 );
nor \U$9043 ( \9175 , \9173 , \9174 );
xnor \U$9044 ( \9176 , \9175 , \202 );
xor \U$9045 ( \9177 , \9172 , \9176 );
and \U$9046 ( \9178 , \7700 , \215 );
and \U$9047 ( \9179 , \8057 , \213 );
nor \U$9048 ( \9180 , \9178 , \9179 );
xnor \U$9049 ( \9181 , \9180 , \222 );
xor \U$9050 ( \9182 , \9177 , \9181 );
and \U$9051 ( \9183 , \7231 , \230 );
and \U$9052 ( \9184 , \7556 , \228 );
nor \U$9053 ( \9185 , \9183 , \9184 );
xnor \U$9054 ( \9186 , \9185 , \237 );
and \U$9055 ( \9187 , \6790 , \245 );
and \U$9056 ( \9188 , \6945 , \243 );
nor \U$9057 ( \9189 , \9187 , \9188 );
xnor \U$9058 ( \9190 , \9189 , \252 );
xor \U$9059 ( \9191 , \9186 , \9190 );
and \U$9060 ( \9192 , \6281 , \141 );
and \U$9061 ( \9193 , \6514 , \139 );
nor \U$9062 ( \9194 , \9192 , \9193 );
xnor \U$9063 ( \9195 , \9194 , \148 );
xor \U$9064 ( \9196 , \9191 , \9195 );
xor \U$9065 ( \9197 , \9182 , \9196 );
and \U$9066 ( \9198 , \5674 , \156 );
and \U$9067 ( \9199 , \6030 , \154 );
nor \U$9068 ( \9200 , \9198 , \9199 );
xnor \U$9069 ( \9201 , \9200 , \163 );
and \U$9070 ( \9202 , \5156 , \296 );
and \U$9071 ( \9203 , \5469 , \168 );
nor \U$9072 ( \9204 , \9202 , \9203 );
xnor \U$9073 ( \9205 , \9204 , \173 );
xor \U$9074 ( \9206 , \9201 , \9205 );
and \U$9075 ( \9207 , \4749 , \438 );
and \U$9076 ( \9208 , \4922 , \336 );
nor \U$9077 ( \9209 , \9207 , \9208 );
xnor \U$9078 ( \9210 , \9209 , \320 );
xor \U$9079 ( \9211 , \9206 , \9210 );
and \U$9080 ( \9212 , \4364 , \1086 );
and \U$9081 ( \9213 , \4654 , \508 );
nor \U$9082 ( \9214 , \9212 , \9213 );
xnor \U$9083 ( \9215 , \9214 , \487 );
and \U$9084 ( \9216 , \3912 , \1301 );
and \U$9085 ( \9217 , \4160 , \1246 );
nor \U$9086 ( \9218 , \9216 , \9217 );
xnor \U$9087 ( \9219 , \9218 , \1205 );
xor \U$9088 ( \9220 , \9215 , \9219 );
and \U$9089 ( \9221 , \3646 , \1578 );
and \U$9090 ( \9222 , \3736 , \1431 );
nor \U$9091 ( \9223 , \9221 , \9222 );
xnor \U$9092 ( \9224 , \9223 , \1436 );
xor \U$9093 ( \9225 , \9220 , \9224 );
xor \U$9094 ( \9226 , \9211 , \9225 );
and \U$9095 ( \9227 , \3143 , \1824 );
and \U$9096 ( \9228 , \3395 , \1739 );
nor \U$9097 ( \9229 , \9227 , \9228 );
xnor \U$9098 ( \9230 , \9229 , \1697 );
and \U$9099 ( \9231 , \2826 , \2121 );
and \U$9100 ( \9232 , \3037 , \2008 );
nor \U$9101 ( \9233 , \9231 , \9232 );
xnor \U$9102 ( \9234 , \9233 , \1961 );
xor \U$9103 ( \9235 , \9230 , \9234 );
and \U$9104 ( \9236 , \2521 , \2400 );
and \U$9105 ( \9237 , \2757 , \2246 );
nor \U$9106 ( \9238 , \9236 , \9237 );
xnor \U$9107 ( \9239 , \9238 , \2195 );
xor \U$9108 ( \9240 , \9235 , \9239 );
xor \U$9109 ( \9241 , \9226 , \9240 );
xor \U$9110 ( \9242 , \9197 , \9241 );
xor \U$9111 ( \9243 , \9167 , \9242 );
and \U$9112 ( \9244 , \8978 , \8982 );
and \U$9113 ( \9245 , \8982 , \8987 );
and \U$9114 ( \9246 , \8978 , \8987 );
or \U$9115 ( \9247 , \9244 , \9245 , \9246 );
and \U$9116 ( \9248 , \8993 , \8997 );
and \U$9117 ( \9249 , \8997 , \9002 );
and \U$9118 ( \9250 , \8993 , \9002 );
or \U$9119 ( \9251 , \9248 , \9249 , \9250 );
xor \U$9120 ( \9252 , \9247 , \9251 );
and \U$9121 ( \9253 , \9012 , \9016 );
and \U$9122 ( \9254 , \9016 , \9021 );
and \U$9123 ( \9255 , \9012 , \9021 );
or \U$9124 ( \9256 , \9253 , \9254 , \9255 );
xor \U$9125 ( \9257 , \9252 , \9256 );
and \U$9126 ( \9258 , \2182 , \2669 );
and \U$9127 ( \9259 , \2366 , \2538 );
nor \U$9128 ( \9260 , \9258 , \9259 );
xnor \U$9129 ( \9261 , \9260 , \2534 );
and \U$9130 ( \9262 , \1948 , \3103 );
and \U$9131 ( \9263 , \2090 , \2934 );
nor \U$9132 ( \9264 , \9262 , \9263 );
xnor \U$9133 ( \9265 , \9264 , \2839 );
xor \U$9134 ( \9266 , \9261 , \9265 );
and \U$9135 ( \9267 , \1684 , \3357 );
and \U$9136 ( \9268 , \1802 , \3255 );
nor \U$9137 ( \9269 , \9267 , \9268 );
xnor \U$9138 ( \9270 , \9269 , \3156 );
xor \U$9139 ( \9271 , \9266 , \9270 );
and \U$9140 ( \9272 , \1484 , \3813 );
and \U$9141 ( \9273 , \1601 , \3557 );
nor \U$9142 ( \9274 , \9272 , \9273 );
xnor \U$9143 ( \9275 , \9274 , \3562 );
and \U$9144 ( \9276 , \1192 , \4132 );
and \U$9145 ( \9277 , \1333 , \4012 );
nor \U$9146 ( \9278 , \9276 , \9277 );
xnor \U$9147 ( \9279 , \9278 , \3925 );
xor \U$9148 ( \9280 , \9275 , \9279 );
and \U$9149 ( \9281 , \474 , \4581 );
and \U$9150 ( \9282 , \1147 , \4424 );
nor \U$9151 ( \9283 , \9281 , \9282 );
xnor \U$9152 ( \9284 , \9283 , \4377 );
xor \U$9153 ( \9285 , \9280 , \9284 );
xor \U$9154 ( \9286 , \9271 , \9285 );
and \U$9155 ( \9287 , \307 , \5011 );
and \U$9156 ( \9288 , \412 , \4878 );
nor \U$9157 ( \9289 , \9287 , \9288 );
xnor \U$9158 ( \9290 , \9289 , \4762 );
and \U$9159 ( \9291 , \185 , \5485 );
and \U$9160 ( \9292 , \261 , \5275 );
nor \U$9161 ( \9293 , \9291 , \9292 );
xnor \U$9162 ( \9294 , \9293 , \5169 );
xor \U$9163 ( \9295 , \9290 , \9294 );
and \U$9164 ( \9296 , \197 , \5996 );
and \U$9165 ( \9297 , \178 , \5695 );
nor \U$9166 ( \9298 , \9296 , \9297 );
xnor \U$9167 ( \9299 , \9298 , \5687 );
xor \U$9168 ( \9300 , \9295 , \9299 );
xor \U$9169 ( \9301 , \9286 , \9300 );
xor \U$9170 ( \9302 , \9257 , \9301 );
and \U$9171 ( \9303 , \9027 , \9031 );
and \U$9172 ( \9304 , \9031 , \9036 );
and \U$9173 ( \9305 , \9027 , \9036 );
or \U$9174 ( \9306 , \9303 , \9304 , \9305 );
and \U$9175 ( \9307 , \217 , \6401 );
and \U$9176 ( \9308 , \189 , \6143 );
nor \U$9177 ( \9309 , \9307 , \9308 );
xnor \U$9178 ( \9310 , \9309 , \6148 );
and \U$9179 ( \9311 , \232 , \7055 );
and \U$9180 ( \9312 , \209 , \6675 );
nor \U$9181 ( \9313 , \9311 , \9312 );
xnor \U$9182 ( \9314 , \9313 , \6680 );
xor \U$9183 ( \9315 , \9310 , \9314 );
and \U$9184 ( \9316 , \247 , \7489 );
and \U$9185 ( \9317 , \224 , \7137 );
nor \U$9186 ( \9318 , \9316 , \9317 );
xnor \U$9187 ( \9319 , \9318 , \7142 );
xor \U$9188 ( \9320 , \9315 , \9319 );
xor \U$9189 ( \9321 , \9306 , \9320 );
and \U$9190 ( \9322 , \143 , \8019 );
and \U$9191 ( \9323 , \240 , \7830 );
nor \U$9192 ( \9324 , \9322 , \9323 );
xnor \U$9193 ( \9325 , \9324 , \7713 );
and \U$9194 ( \9326 , \158 , \8540 );
and \U$9195 ( \9327 , \134 , \8292 );
nor \U$9196 ( \9328 , \9326 , \9327 );
xnor \U$9197 ( \9329 , \9328 , \8297 );
xor \U$9198 ( \9330 , \9325 , \9329 );
xor \U$9199 ( \9331 , \8844 , \8845 );
not \U$9200 ( \9332 , \9006 );
and \U$9201 ( \9333 , \9331 , \9332 );
and \U$9202 ( \9334 , \166 , \9333 );
and \U$9203 ( \9335 , \150 , \9006 );
nor \U$9204 ( \9336 , \9334 , \9335 );
xnor \U$9205 ( \9337 , \9336 , \8848 );
xor \U$9206 ( \9338 , \9330 , \9337 );
xor \U$9207 ( \9339 , \9321 , \9338 );
xor \U$9208 ( \9340 , \9302 , \9339 );
xor \U$9209 ( \9341 , \9243 , \9340 );
xor \U$9210 ( \9342 , \9153 , \9341 );
xor \U$9211 ( \9343 , \9124 , \9342 );
xor \U$9212 ( \9344 , \9095 , \9343 );
xor \U$9213 ( \9345 , \9056 , \9344 );
and \U$9214 ( \9346 , \8758 , \9043 );
xor \U$9215 ( \9347 , \9345 , \9346 );
and \U$9216 ( \9348 , \9044 , \9045 );
and \U$9217 ( \9349 , \9046 , \9049 );
or \U$9218 ( \9350 , \9348 , \9349 );
xor \U$9219 ( \9351 , \9347 , \9350 );
buf \U$9220 ( \9352 , \9351 );
buf \U$9221 ( \9353 , \9352 );
and \U$9222 ( \9354 , \9060 , \9094 );
and \U$9223 ( \9355 , \9094 , \9343 );
and \U$9224 ( \9356 , \9060 , \9343 );
or \U$9225 ( \9357 , \9354 , \9355 , \9356 );
and \U$9226 ( \9358 , \9064 , \9068 );
and \U$9227 ( \9359 , \9068 , \9093 );
and \U$9228 ( \9360 , \9064 , \9093 );
or \U$9229 ( \9361 , \9358 , \9359 , \9360 );
and \U$9230 ( \9362 , \9109 , \9123 );
and \U$9231 ( \9363 , \9123 , \9342 );
and \U$9232 ( \9364 , \9109 , \9342 );
or \U$9233 ( \9365 , \9362 , \9363 , \9364 );
xor \U$9234 ( \9366 , \9361 , \9365 );
and \U$9235 ( \9367 , \9099 , \9103 );
and \U$9236 ( \9368 , \9103 , \9108 );
and \U$9237 ( \9369 , \9099 , \9108 );
or \U$9238 ( \9370 , \9367 , \9368 , \9369 );
and \U$9239 ( \9371 , \9073 , \9077 );
and \U$9240 ( \9372 , \9077 , \9092 );
and \U$9241 ( \9373 , \9073 , \9092 );
or \U$9242 ( \9374 , \9371 , \9372 , \9373 );
xor \U$9243 ( \9375 , \9370 , \9374 );
and \U$9244 ( \9376 , \9167 , \9242 );
and \U$9245 ( \9377 , \9242 , \9340 );
and \U$9246 ( \9378 , \9167 , \9340 );
or \U$9247 ( \9379 , \9376 , \9377 , \9378 );
xor \U$9248 ( \9380 , \9375 , \9379 );
xor \U$9249 ( \9381 , \9366 , \9380 );
xor \U$9250 ( \9382 , \9357 , \9381 );
and \U$9251 ( \9383 , \9113 , \9117 );
and \U$9252 ( \9384 , \9117 , \9122 );
and \U$9253 ( \9385 , \9113 , \9122 );
or \U$9254 ( \9386 , \9383 , \9384 , \9385 );
and \U$9255 ( \9387 , \9138 , \9152 );
and \U$9256 ( \9388 , \9152 , \9341 );
and \U$9257 ( \9389 , \9138 , \9341 );
or \U$9258 ( \9390 , \9387 , \9388 , \9389 );
xor \U$9259 ( \9391 , \9386 , \9390 );
and \U$9260 ( \9392 , \9128 , \9132 );
and \U$9261 ( \9393 , \9132 , \9137 );
and \U$9262 ( \9394 , \9128 , \9137 );
or \U$9263 ( \9395 , \9392 , \9393 , \9394 );
and \U$9264 ( \9396 , \9142 , \9146 );
and \U$9265 ( \9397 , \9146 , \9151 );
and \U$9266 ( \9398 , \9142 , \9151 );
or \U$9267 ( \9399 , \9396 , \9397 , \9398 );
xor \U$9268 ( \9400 , \9395 , \9399 );
and \U$9269 ( \9401 , \9182 , \9196 );
and \U$9270 ( \9402 , \9196 , \9241 );
and \U$9271 ( \9403 , \9182 , \9241 );
or \U$9272 ( \9404 , \9401 , \9402 , \9403 );
xor \U$9273 ( \9405 , \9400 , \9404 );
and \U$9274 ( \9406 , \9271 , \9285 );
and \U$9275 ( \9407 , \9285 , \9300 );
and \U$9276 ( \9408 , \9271 , \9300 );
or \U$9277 ( \9409 , \9406 , \9407 , \9408 );
and \U$9278 ( \9410 , \9306 , \9320 );
and \U$9279 ( \9411 , \9320 , \9338 );
and \U$9280 ( \9412 , \9306 , \9338 );
or \U$9281 ( \9413 , \9410 , \9411 , \9412 );
xor \U$9282 ( \9414 , \9409 , \9413 );
and \U$9283 ( \9415 , \9211 , \9225 );
and \U$9284 ( \9416 , \9225 , \9240 );
and \U$9285 ( \9417 , \9211 , \9240 );
or \U$9286 ( \9418 , \9415 , \9416 , \9417 );
xor \U$9287 ( \9419 , \9414 , \9418 );
and \U$9288 ( \9420 , \9157 , \9161 );
and \U$9289 ( \9421 , \9161 , \9166 );
and \U$9290 ( \9422 , \9157 , \9166 );
or \U$9291 ( \9423 , \9420 , \9421 , \9422 );
and \U$9292 ( \9424 , \9082 , \9086 );
and \U$9293 ( \9425 , \9086 , \9091 );
and \U$9294 ( \9426 , \9082 , \9091 );
or \U$9295 ( \9427 , \9424 , \9425 , \9426 );
xor \U$9296 ( \9428 , \9423 , \9427 );
and \U$9297 ( \9429 , \9247 , \9251 );
and \U$9298 ( \9430 , \9251 , \9256 );
and \U$9299 ( \9431 , \9247 , \9256 );
or \U$9300 ( \9432 , \9429 , \9430 , \9431 );
xor \U$9301 ( \9433 , \9428 , \9432 );
xor \U$9302 ( \9434 , \9419 , \9433 );
and \U$9303 ( \9435 , \6514 , \141 );
and \U$9304 ( \9436 , \6790 , \139 );
nor \U$9305 ( \9437 , \9435 , \9436 );
xnor \U$9306 ( \9438 , \9437 , \148 );
and \U$9307 ( \9439 , \6030 , \156 );
and \U$9308 ( \9440 , \6281 , \154 );
nor \U$9309 ( \9441 , \9439 , \9440 );
xnor \U$9310 ( \9442 , \9441 , \163 );
xor \U$9311 ( \9443 , \9438 , \9442 );
and \U$9312 ( \9444 , \5469 , \296 );
and \U$9313 ( \9445 , \5674 , \168 );
nor \U$9314 ( \9446 , \9444 , \9445 );
xnor \U$9315 ( \9447 , \9446 , \173 );
xor \U$9316 ( \9448 , \9443 , \9447 );
and \U$9317 ( \9449 , \8057 , \215 );
and \U$9318 ( \9450 , \8349 , \213 );
nor \U$9319 ( \9451 , \9449 , \9450 );
xnor \U$9320 ( \9452 , \9451 , \222 );
and \U$9321 ( \9453 , \7556 , \230 );
and \U$9322 ( \9454 , \7700 , \228 );
nor \U$9323 ( \9455 , \9453 , \9454 );
xnor \U$9324 ( \9456 , \9455 , \237 );
xor \U$9325 ( \9457 , \9452 , \9456 );
and \U$9326 ( \9458 , \6945 , \245 );
and \U$9327 ( \9459 , \7231 , \243 );
nor \U$9328 ( \9460 , \9458 , \9459 );
xnor \U$9329 ( \9461 , \9460 , \252 );
xor \U$9330 ( \9462 , \9457 , \9461 );
xor \U$9331 ( \9463 , \9448 , \9462 );
and \U$9332 ( \9464 , \9169 , \183 );
buf \U$9333 ( \9465 , RIb55f058_68);
and \U$9334 ( \9466 , \9465 , \180 );
nor \U$9335 ( \9467 , \9464 , \9466 );
xnor \U$9336 ( \9468 , \9467 , \179 );
and \U$9337 ( \9469 , \8652 , \195 );
and \U$9338 ( \9470 , \8835 , \193 );
nor \U$9339 ( \9471 , \9469 , \9470 );
xnor \U$9340 ( \9472 , \9471 , \202 );
xor \U$9341 ( \9473 , \9468 , \9472 );
buf \U$9342 ( \9474 , RIb560ed0_3);
buf \U$9343 ( \9475 , RIb560e58_4);
and \U$9344 ( \9476 , \9475 , \8844 );
not \U$9345 ( \9477 , \9476 );
and \U$9346 ( \9478 , \9474 , \9477 );
xor \U$9347 ( \9479 , \9473 , \9478 );
xor \U$9348 ( \9480 , \9463 , \9479 );
and \U$9349 ( \9481 , \178 , \5996 );
and \U$9350 ( \9482 , \185 , \5695 );
nor \U$9351 ( \9483 , \9481 , \9482 );
xnor \U$9352 ( \9484 , \9483 , \5687 );
and \U$9353 ( \9485 , \189 , \6401 );
and \U$9354 ( \9486 , \197 , \6143 );
nor \U$9355 ( \9487 , \9485 , \9486 );
xnor \U$9356 ( \9488 , \9487 , \6148 );
xor \U$9357 ( \9489 , \9484 , \9488 );
and \U$9358 ( \9490 , \209 , \7055 );
and \U$9359 ( \9491 , \217 , \6675 );
nor \U$9360 ( \9492 , \9490 , \9491 );
xnor \U$9361 ( \9493 , \9492 , \6680 );
xor \U$9362 ( \9494 , \9489 , \9493 );
and \U$9363 ( \9495 , \1802 , \3357 );
and \U$9364 ( \9496 , \1948 , \3255 );
nor \U$9365 ( \9497 , \9495 , \9496 );
xnor \U$9366 ( \9498 , \9497 , \3156 );
and \U$9367 ( \9499 , \1601 , \3813 );
and \U$9368 ( \9500 , \1684 , \3557 );
nor \U$9369 ( \9501 , \9499 , \9500 );
xnor \U$9370 ( \9502 , \9501 , \3562 );
xor \U$9371 ( \9503 , \9498 , \9502 );
and \U$9372 ( \9504 , \1333 , \4132 );
and \U$9373 ( \9505 , \1484 , \4012 );
nor \U$9374 ( \9506 , \9504 , \9505 );
xnor \U$9375 ( \9507 , \9506 , \3925 );
xor \U$9376 ( \9508 , \9503 , \9507 );
xor \U$9377 ( \9509 , \9494 , \9508 );
and \U$9378 ( \9510 , \1147 , \4581 );
and \U$9379 ( \9511 , \1192 , \4424 );
nor \U$9380 ( \9512 , \9510 , \9511 );
xnor \U$9381 ( \9513 , \9512 , \4377 );
and \U$9382 ( \9514 , \412 , \5011 );
and \U$9383 ( \9515 , \474 , \4878 );
nor \U$9384 ( \9516 , \9514 , \9515 );
xnor \U$9385 ( \9517 , \9516 , \4762 );
xor \U$9386 ( \9518 , \9513 , \9517 );
and \U$9387 ( \9519 , \261 , \5485 );
and \U$9388 ( \9520 , \307 , \5275 );
nor \U$9389 ( \9521 , \9519 , \9520 );
xnor \U$9390 ( \9522 , \9521 , \5169 );
xor \U$9391 ( \9523 , \9518 , \9522 );
xor \U$9392 ( \9524 , \9509 , \9523 );
xor \U$9393 ( \9525 , \9480 , \9524 );
and \U$9394 ( \9526 , \4922 , \438 );
and \U$9395 ( \9527 , \5156 , \336 );
nor \U$9396 ( \9528 , \9526 , \9527 );
xnor \U$9397 ( \9529 , \9528 , \320 );
and \U$9398 ( \9530 , \4654 , \1086 );
and \U$9399 ( \9531 , \4749 , \508 );
nor \U$9400 ( \9532 , \9530 , \9531 );
xnor \U$9401 ( \9533 , \9532 , \487 );
xor \U$9402 ( \9534 , \9529 , \9533 );
and \U$9403 ( \9535 , \4160 , \1301 );
and \U$9404 ( \9536 , \4364 , \1246 );
nor \U$9405 ( \9537 , \9535 , \9536 );
xnor \U$9406 ( \9538 , \9537 , \1205 );
xor \U$9407 ( \9539 , \9534 , \9538 );
and \U$9408 ( \9540 , \3736 , \1578 );
and \U$9409 ( \9541 , \3912 , \1431 );
nor \U$9410 ( \9542 , \9540 , \9541 );
xnor \U$9411 ( \9543 , \9542 , \1436 );
and \U$9412 ( \9544 , \3395 , \1824 );
and \U$9413 ( \9545 , \3646 , \1739 );
nor \U$9414 ( \9546 , \9544 , \9545 );
xnor \U$9415 ( \9547 , \9546 , \1697 );
xor \U$9416 ( \9548 , \9543 , \9547 );
and \U$9417 ( \9549 , \3037 , \2121 );
and \U$9418 ( \9550 , \3143 , \2008 );
nor \U$9419 ( \9551 , \9549 , \9550 );
xnor \U$9420 ( \9552 , \9551 , \1961 );
xor \U$9421 ( \9553 , \9548 , \9552 );
xor \U$9422 ( \9554 , \9539 , \9553 );
and \U$9423 ( \9555 , \2757 , \2400 );
and \U$9424 ( \9556 , \2826 , \2246 );
nor \U$9425 ( \9557 , \9555 , \9556 );
xnor \U$9426 ( \9558 , \9557 , \2195 );
and \U$9427 ( \9559 , \2366 , \2669 );
and \U$9428 ( \9560 , \2521 , \2538 );
nor \U$9429 ( \9561 , \9559 , \9560 );
xnor \U$9430 ( \9562 , \9561 , \2534 );
xor \U$9431 ( \9563 , \9558 , \9562 );
and \U$9432 ( \9564 , \2090 , \3103 );
and \U$9433 ( \9565 , \2182 , \2934 );
nor \U$9434 ( \9566 , \9564 , \9565 );
xnor \U$9435 ( \9567 , \9566 , \2839 );
xor \U$9436 ( \9568 , \9563 , \9567 );
xor \U$9437 ( \9569 , \9554 , \9568 );
xor \U$9438 ( \9570 , \9525 , \9569 );
xor \U$9439 ( \9571 , \9434 , \9570 );
xor \U$9440 ( \9572 , \9405 , \9571 );
and \U$9441 ( \9573 , \9257 , \9301 );
and \U$9442 ( \9574 , \9301 , \9339 );
and \U$9443 ( \9575 , \9257 , \9339 );
or \U$9444 ( \9576 , \9573 , \9574 , \9575 );
and \U$9445 ( \9577 , \9201 , \9205 );
and \U$9446 ( \9578 , \9205 , \9210 );
and \U$9447 ( \9579 , \9201 , \9210 );
or \U$9448 ( \9580 , \9577 , \9578 , \9579 );
and \U$9449 ( \9581 , \9172 , \9176 );
and \U$9450 ( \9582 , \9176 , \9181 );
and \U$9451 ( \9583 , \9172 , \9181 );
or \U$9452 ( \9584 , \9581 , \9582 , \9583 );
xor \U$9453 ( \9585 , \9580 , \9584 );
and \U$9454 ( \9586 , \9186 , \9190 );
and \U$9455 ( \9587 , \9190 , \9195 );
and \U$9456 ( \9588 , \9186 , \9195 );
or \U$9457 ( \9589 , \9586 , \9587 , \9588 );
xor \U$9458 ( \9590 , \9585 , \9589 );
xor \U$9459 ( \9591 , \9576 , \9590 );
and \U$9460 ( \9592 , \9261 , \9265 );
and \U$9461 ( \9593 , \9265 , \9270 );
and \U$9462 ( \9594 , \9261 , \9270 );
or \U$9463 ( \9595 , \9592 , \9593 , \9594 );
and \U$9464 ( \9596 , \9215 , \9219 );
and \U$9465 ( \9597 , \9219 , \9224 );
and \U$9466 ( \9598 , \9215 , \9224 );
or \U$9467 ( \9599 , \9596 , \9597 , \9598 );
xor \U$9468 ( \9600 , \9595 , \9599 );
and \U$9469 ( \9601 , \9230 , \9234 );
and \U$9470 ( \9602 , \9234 , \9239 );
and \U$9471 ( \9603 , \9230 , \9239 );
or \U$9472 ( \9604 , \9601 , \9602 , \9603 );
xor \U$9473 ( \9605 , \9600 , \9604 );
and \U$9474 ( \9606 , \9275 , \9279 );
and \U$9475 ( \9607 , \9279 , \9284 );
and \U$9476 ( \9608 , \9275 , \9284 );
or \U$9477 ( \9609 , \9606 , \9607 , \9608 );
and \U$9478 ( \9610 , \9310 , \9314 );
and \U$9479 ( \9611 , \9314 , \9319 );
and \U$9480 ( \9612 , \9310 , \9319 );
or \U$9481 ( \9613 , \9610 , \9611 , \9612 );
xor \U$9482 ( \9614 , \9609 , \9613 );
and \U$9483 ( \9615 , \9290 , \9294 );
and \U$9484 ( \9616 , \9294 , \9299 );
and \U$9485 ( \9617 , \9290 , \9299 );
or \U$9486 ( \9618 , \9615 , \9616 , \9617 );
xor \U$9487 ( \9619 , \9614 , \9618 );
xor \U$9488 ( \9620 , \9605 , \9619 );
and \U$9489 ( \9621 , \9325 , \9329 );
and \U$9490 ( \9622 , \9329 , \9337 );
and \U$9491 ( \9623 , \9325 , \9337 );
or \U$9492 ( \9624 , \9621 , \9622 , \9623 );
and \U$9493 ( \9625 , \224 , \7489 );
and \U$9494 ( \9626 , \232 , \7137 );
nor \U$9495 ( \9627 , \9625 , \9626 );
xnor \U$9496 ( \9628 , \9627 , \7142 );
and \U$9497 ( \9629 , \240 , \8019 );
and \U$9498 ( \9630 , \247 , \7830 );
nor \U$9499 ( \9631 , \9629 , \9630 );
xnor \U$9500 ( \9632 , \9631 , \7713 );
xor \U$9501 ( \9633 , \9628 , \9632 );
and \U$9502 ( \9634 , \134 , \8540 );
and \U$9503 ( \9635 , \143 , \8292 );
nor \U$9504 ( \9636 , \9634 , \9635 );
xnor \U$9505 ( \9637 , \9636 , \8297 );
xor \U$9506 ( \9638 , \9633 , \9637 );
xor \U$9507 ( \9639 , \9624 , \9638 );
and \U$9508 ( \9640 , \150 , \9333 );
and \U$9509 ( \9641 , \158 , \9006 );
nor \U$9510 ( \9642 , \9640 , \9641 );
xnor \U$9511 ( \9643 , \9642 , \8848 );
xor \U$9512 ( \9644 , \9475 , \8844 );
nand \U$9513 ( \9645 , \166 , \9644 );
xnor \U$9514 ( \9646 , \9645 , \9478 );
xor \U$9515 ( \9647 , \9643 , \9646 );
xor \U$9516 ( \9648 , \9639 , \9647 );
xor \U$9517 ( \9649 , \9620 , \9648 );
xor \U$9518 ( \9650 , \9591 , \9649 );
xor \U$9519 ( \9651 , \9572 , \9650 );
xor \U$9520 ( \9652 , \9391 , \9651 );
xor \U$9521 ( \9653 , \9382 , \9652 );
and \U$9522 ( \9654 , \9056 , \9344 );
xor \U$9523 ( \9655 , \9653 , \9654 );
and \U$9524 ( \9656 , \9345 , \9346 );
and \U$9525 ( \9657 , \9347 , \9350 );
or \U$9526 ( \9658 , \9656 , \9657 );
xor \U$9527 ( \9659 , \9655 , \9658 );
buf \U$9528 ( \9660 , \9659 );
buf \U$9529 ( \9661 , \9660 );
and \U$9530 ( \9662 , \9361 , \9365 );
and \U$9531 ( \9663 , \9365 , \9380 );
and \U$9532 ( \9664 , \9361 , \9380 );
or \U$9533 ( \9665 , \9662 , \9663 , \9664 );
and \U$9534 ( \9666 , \9386 , \9390 );
and \U$9535 ( \9667 , \9390 , \9651 );
and \U$9536 ( \9668 , \9386 , \9651 );
or \U$9537 ( \9669 , \9666 , \9667 , \9668 );
and \U$9538 ( \9670 , \9395 , \9399 );
and \U$9539 ( \9671 , \9399 , \9404 );
and \U$9540 ( \9672 , \9395 , \9404 );
or \U$9541 ( \9673 , \9670 , \9671 , \9672 );
and \U$9542 ( \9674 , \9419 , \9433 );
and \U$9543 ( \9675 , \9433 , \9570 );
and \U$9544 ( \9676 , \9419 , \9570 );
or \U$9545 ( \9677 , \9674 , \9675 , \9676 );
xor \U$9546 ( \9678 , \9673 , \9677 );
and \U$9547 ( \9679 , \9576 , \9590 );
and \U$9548 ( \9680 , \9590 , \9649 );
and \U$9549 ( \9681 , \9576 , \9649 );
or \U$9550 ( \9682 , \9679 , \9680 , \9681 );
xor \U$9551 ( \9683 , \9678 , \9682 );
xor \U$9552 ( \9684 , \9669 , \9683 );
and \U$9553 ( \9685 , \9370 , \9374 );
and \U$9554 ( \9686 , \9374 , \9379 );
and \U$9555 ( \9687 , \9370 , \9379 );
or \U$9556 ( \9688 , \9685 , \9686 , \9687 );
and \U$9557 ( \9689 , \9405 , \9571 );
and \U$9558 ( \9690 , \9571 , \9650 );
and \U$9559 ( \9691 , \9405 , \9650 );
or \U$9560 ( \9692 , \9689 , \9690 , \9691 );
xor \U$9561 ( \9693 , \9688 , \9692 );
and \U$9562 ( \9694 , \9409 , \9413 );
and \U$9563 ( \9695 , \9413 , \9418 );
and \U$9564 ( \9696 , \9409 , \9418 );
or \U$9565 ( \9697 , \9694 , \9695 , \9696 );
and \U$9566 ( \9698 , \9423 , \9427 );
and \U$9567 ( \9699 , \9427 , \9432 );
and \U$9568 ( \9700 , \9423 , \9432 );
or \U$9569 ( \9701 , \9698 , \9699 , \9700 );
xor \U$9570 ( \9702 , \9697 , \9701 );
and \U$9571 ( \9703 , \9480 , \9524 );
and \U$9572 ( \9704 , \9524 , \9569 );
and \U$9573 ( \9705 , \9480 , \9569 );
or \U$9574 ( \9706 , \9703 , \9704 , \9705 );
xor \U$9575 ( \9707 , \9702 , \9706 );
and \U$9576 ( \9708 , \9605 , \9619 );
and \U$9577 ( \9709 , \9619 , \9648 );
and \U$9578 ( \9710 , \9605 , \9648 );
or \U$9579 ( \9711 , \9708 , \9709 , \9710 );
and \U$9580 ( \9712 , \9484 , \9488 );
and \U$9581 ( \9713 , \9488 , \9493 );
and \U$9582 ( \9714 , \9484 , \9493 );
or \U$9583 ( \9715 , \9712 , \9713 , \9714 );
and \U$9584 ( \9716 , \9498 , \9502 );
and \U$9585 ( \9717 , \9502 , \9507 );
and \U$9586 ( \9718 , \9498 , \9507 );
or \U$9587 ( \9719 , \9716 , \9717 , \9718 );
xor \U$9588 ( \9720 , \9715 , \9719 );
and \U$9589 ( \9721 , \9513 , \9517 );
and \U$9590 ( \9722 , \9517 , \9522 );
and \U$9591 ( \9723 , \9513 , \9522 );
or \U$9592 ( \9724 , \9721 , \9722 , \9723 );
xor \U$9593 ( \9725 , \9720 , \9724 );
and \U$9594 ( \9726 , \9438 , \9442 );
and \U$9595 ( \9727 , \9442 , \9447 );
and \U$9596 ( \9728 , \9438 , \9447 );
or \U$9597 ( \9729 , \9726 , \9727 , \9728 );
and \U$9598 ( \9730 , \9452 , \9456 );
and \U$9599 ( \9731 , \9456 , \9461 );
and \U$9600 ( \9732 , \9452 , \9461 );
or \U$9601 ( \9733 , \9730 , \9731 , \9732 );
xor \U$9602 ( \9734 , \9729 , \9733 );
and \U$9603 ( \9735 , \9468 , \9472 );
and \U$9604 ( \9736 , \9472 , \9478 );
and \U$9605 ( \9737 , \9468 , \9478 );
or \U$9606 ( \9738 , \9735 , \9736 , \9737 );
xor \U$9607 ( \9739 , \9734 , \9738 );
xor \U$9608 ( \9740 , \9725 , \9739 );
and \U$9609 ( \9741 , \9529 , \9533 );
and \U$9610 ( \9742 , \9533 , \9538 );
and \U$9611 ( \9743 , \9529 , \9538 );
or \U$9612 ( \9744 , \9741 , \9742 , \9743 );
and \U$9613 ( \9745 , \9543 , \9547 );
and \U$9614 ( \9746 , \9547 , \9552 );
and \U$9615 ( \9747 , \9543 , \9552 );
or \U$9616 ( \9748 , \9745 , \9746 , \9747 );
xor \U$9617 ( \9749 , \9744 , \9748 );
and \U$9618 ( \9750 , \9558 , \9562 );
and \U$9619 ( \9751 , \9562 , \9567 );
and \U$9620 ( \9752 , \9558 , \9567 );
or \U$9621 ( \9753 , \9750 , \9751 , \9752 );
xor \U$9622 ( \9754 , \9749 , \9753 );
xor \U$9623 ( \9755 , \9740 , \9754 );
xor \U$9624 ( \9756 , \9711 , \9755 );
and \U$9625 ( \9757 , \9628 , \9632 );
and \U$9626 ( \9758 , \9632 , \9637 );
and \U$9627 ( \9759 , \9628 , \9637 );
or \U$9628 ( \9760 , \9757 , \9758 , \9759 );
and \U$9629 ( \9761 , \9643 , \9646 );
xor \U$9630 ( \9762 , \9760 , \9761 );
xor \U$9631 ( \9763 , \9474 , \9475 );
not \U$9632 ( \9764 , \9644 );
and \U$9633 ( \9765 , \9763 , \9764 );
and \U$9634 ( \9766 , \166 , \9765 );
and \U$9635 ( \9767 , \150 , \9644 );
nor \U$9636 ( \9768 , \9766 , \9767 );
xnor \U$9637 ( \9769 , \9768 , \9478 );
xor \U$9638 ( \9770 , \9762 , \9769 );
and \U$9639 ( \9771 , \1684 , \3813 );
and \U$9640 ( \9772 , \1802 , \3557 );
nor \U$9641 ( \9773 , \9771 , \9772 );
xnor \U$9642 ( \9774 , \9773 , \3562 );
and \U$9643 ( \9775 , \1484 , \4132 );
and \U$9644 ( \9776 , \1601 , \4012 );
nor \U$9645 ( \9777 , \9775 , \9776 );
xnor \U$9646 ( \9778 , \9777 , \3925 );
xor \U$9647 ( \9779 , \9774 , \9778 );
and \U$9648 ( \9780 , \1192 , \4581 );
and \U$9649 ( \9781 , \1333 , \4424 );
nor \U$9650 ( \9782 , \9780 , \9781 );
xnor \U$9651 ( \9783 , \9782 , \4377 );
xor \U$9652 ( \9784 , \9779 , \9783 );
and \U$9653 ( \9785 , \2521 , \2669 );
and \U$9654 ( \9786 , \2757 , \2538 );
nor \U$9655 ( \9787 , \9785 , \9786 );
xnor \U$9656 ( \9788 , \9787 , \2534 );
and \U$9657 ( \9789 , \2182 , \3103 );
and \U$9658 ( \9790 , \2366 , \2934 );
nor \U$9659 ( \9791 , \9789 , \9790 );
xnor \U$9660 ( \9792 , \9791 , \2839 );
xor \U$9661 ( \9793 , \9788 , \9792 );
and \U$9662 ( \9794 , \1948 , \3357 );
and \U$9663 ( \9795 , \2090 , \3255 );
nor \U$9664 ( \9796 , \9794 , \9795 );
xnor \U$9665 ( \9797 , \9796 , \3156 );
xor \U$9666 ( \9798 , \9793 , \9797 );
xor \U$9667 ( \9799 , \9784 , \9798 );
and \U$9668 ( \9800 , \3646 , \1824 );
and \U$9669 ( \9801 , \3736 , \1739 );
nor \U$9670 ( \9802 , \9800 , \9801 );
xnor \U$9671 ( \9803 , \9802 , \1697 );
and \U$9672 ( \9804 , \3143 , \2121 );
and \U$9673 ( \9805 , \3395 , \2008 );
nor \U$9674 ( \9806 , \9804 , \9805 );
xnor \U$9675 ( \9807 , \9806 , \1961 );
xor \U$9676 ( \9808 , \9803 , \9807 );
and \U$9677 ( \9809 , \2826 , \2400 );
and \U$9678 ( \9810 , \3037 , \2246 );
nor \U$9679 ( \9811 , \9809 , \9810 );
xnor \U$9680 ( \9812 , \9811 , \2195 );
xor \U$9681 ( \9813 , \9808 , \9812 );
xor \U$9682 ( \9814 , \9799 , \9813 );
xor \U$9683 ( \9815 , \9770 , \9814 );
and \U$9684 ( \9816 , \474 , \5011 );
and \U$9685 ( \9817 , \1147 , \4878 );
nor \U$9686 ( \9818 , \9816 , \9817 );
xnor \U$9687 ( \9819 , \9818 , \4762 );
and \U$9688 ( \9820 , \307 , \5485 );
and \U$9689 ( \9821 , \412 , \5275 );
nor \U$9690 ( \9822 , \9820 , \9821 );
xnor \U$9691 ( \9823 , \9822 , \5169 );
xor \U$9692 ( \9824 , \9819 , \9823 );
and \U$9693 ( \9825 , \185 , \5996 );
and \U$9694 ( \9826 , \261 , \5695 );
nor \U$9695 ( \9827 , \9825 , \9826 );
xnor \U$9696 ( \9828 , \9827 , \5687 );
xor \U$9697 ( \9829 , \9824 , \9828 );
and \U$9698 ( \9830 , \197 , \6401 );
and \U$9699 ( \9831 , \178 , \6143 );
nor \U$9700 ( \9832 , \9830 , \9831 );
xnor \U$9701 ( \9833 , \9832 , \6148 );
and \U$9702 ( \9834 , \217 , \7055 );
and \U$9703 ( \9835 , \189 , \6675 );
nor \U$9704 ( \9836 , \9834 , \9835 );
xnor \U$9705 ( \9837 , \9836 , \6680 );
xor \U$9706 ( \9838 , \9833 , \9837 );
and \U$9707 ( \9839 , \232 , \7489 );
and \U$9708 ( \9840 , \209 , \7137 );
nor \U$9709 ( \9841 , \9839 , \9840 );
xnor \U$9710 ( \9842 , \9841 , \7142 );
xor \U$9711 ( \9843 , \9838 , \9842 );
xor \U$9712 ( \9844 , \9829 , \9843 );
and \U$9713 ( \9845 , \247 , \8019 );
and \U$9714 ( \9846 , \224 , \7830 );
nor \U$9715 ( \9847 , \9845 , \9846 );
xnor \U$9716 ( \9848 , \9847 , \7713 );
and \U$9717 ( \9849 , \143 , \8540 );
and \U$9718 ( \9850 , \240 , \8292 );
nor \U$9719 ( \9851 , \9849 , \9850 );
xnor \U$9720 ( \9852 , \9851 , \8297 );
xor \U$9721 ( \9853 , \9848 , \9852 );
and \U$9722 ( \9854 , \158 , \9333 );
and \U$9723 ( \9855 , \134 , \9006 );
nor \U$9724 ( \9856 , \9854 , \9855 );
xnor \U$9725 ( \9857 , \9856 , \8848 );
xor \U$9726 ( \9858 , \9853 , \9857 );
xor \U$9727 ( \9859 , \9844 , \9858 );
xor \U$9728 ( \9860 , \9815 , \9859 );
xor \U$9729 ( \9861 , \9756 , \9860 );
xor \U$9730 ( \9862 , \9707 , \9861 );
and \U$9731 ( \9863 , \9494 , \9508 );
and \U$9732 ( \9864 , \9508 , \9523 );
and \U$9733 ( \9865 , \9494 , \9523 );
or \U$9734 ( \9866 , \9863 , \9864 , \9865 );
and \U$9735 ( \9867 , \9539 , \9553 );
and \U$9736 ( \9868 , \9553 , \9568 );
and \U$9737 ( \9869 , \9539 , \9568 );
or \U$9738 ( \9870 , \9867 , \9868 , \9869 );
xor \U$9739 ( \9871 , \9866 , \9870 );
and \U$9740 ( \9872 , \9624 , \9638 );
and \U$9741 ( \9873 , \9638 , \9647 );
and \U$9742 ( \9874 , \9624 , \9647 );
or \U$9743 ( \9875 , \9872 , \9873 , \9874 );
xor \U$9744 ( \9876 , \9871 , \9875 );
and \U$9745 ( \9877 , \9595 , \9599 );
and \U$9746 ( \9878 , \9599 , \9604 );
and \U$9747 ( \9879 , \9595 , \9604 );
or \U$9748 ( \9880 , \9877 , \9878 , \9879 );
and \U$9749 ( \9881 , \9580 , \9584 );
and \U$9750 ( \9882 , \9584 , \9589 );
and \U$9751 ( \9883 , \9580 , \9589 );
or \U$9752 ( \9884 , \9881 , \9882 , \9883 );
xor \U$9753 ( \9885 , \9880 , \9884 );
and \U$9754 ( \9886 , \9609 , \9613 );
and \U$9755 ( \9887 , \9613 , \9618 );
and \U$9756 ( \9888 , \9609 , \9618 );
or \U$9757 ( \9889 , \9886 , \9887 , \9888 );
xor \U$9758 ( \9890 , \9885 , \9889 );
xor \U$9759 ( \9891 , \9876 , \9890 );
and \U$9760 ( \9892 , \9448 , \9462 );
and \U$9761 ( \9893 , \9462 , \9479 );
and \U$9762 ( \9894 , \9448 , \9479 );
or \U$9763 ( \9895 , \9892 , \9893 , \9894 );
and \U$9764 ( \9896 , \9465 , \183 );
buf \U$9765 ( \9897 , RIb55f0d0_67);
and \U$9766 ( \9898 , \9897 , \180 );
nor \U$9767 ( \9899 , \9896 , \9898 );
xnor \U$9768 ( \9900 , \9899 , \179 );
and \U$9769 ( \9901 , \8835 , \195 );
and \U$9770 ( \9902 , \9169 , \193 );
nor \U$9771 ( \9903 , \9901 , \9902 );
xnor \U$9772 ( \9904 , \9903 , \202 );
xor \U$9773 ( \9905 , \9900 , \9904 );
and \U$9774 ( \9906 , \8349 , \215 );
and \U$9775 ( \9907 , \8652 , \213 );
nor \U$9776 ( \9908 , \9906 , \9907 );
xnor \U$9777 ( \9909 , \9908 , \222 );
xor \U$9778 ( \9910 , \9905 , \9909 );
xor \U$9779 ( \9911 , \9895 , \9910 );
and \U$9780 ( \9912 , \7700 , \230 );
and \U$9781 ( \9913 , \8057 , \228 );
nor \U$9782 ( \9914 , \9912 , \9913 );
xnor \U$9783 ( \9915 , \9914 , \237 );
and \U$9784 ( \9916 , \7231 , \245 );
and \U$9785 ( \9917 , \7556 , \243 );
nor \U$9786 ( \9918 , \9916 , \9917 );
xnor \U$9787 ( \9919 , \9918 , \252 );
xor \U$9788 ( \9920 , \9915 , \9919 );
and \U$9789 ( \9921 , \6790 , \141 );
and \U$9790 ( \9922 , \6945 , \139 );
nor \U$9791 ( \9923 , \9921 , \9922 );
xnor \U$9792 ( \9924 , \9923 , \148 );
xor \U$9793 ( \9925 , \9920 , \9924 );
and \U$9794 ( \9926 , \4749 , \1086 );
and \U$9795 ( \9927 , \4922 , \508 );
nor \U$9796 ( \9928 , \9926 , \9927 );
xnor \U$9797 ( \9929 , \9928 , \487 );
and \U$9798 ( \9930 , \4364 , \1301 );
and \U$9799 ( \9931 , \4654 , \1246 );
nor \U$9800 ( \9932 , \9930 , \9931 );
xnor \U$9801 ( \9933 , \9932 , \1205 );
xor \U$9802 ( \9934 , \9929 , \9933 );
and \U$9803 ( \9935 , \3912 , \1578 );
and \U$9804 ( \9936 , \4160 , \1431 );
nor \U$9805 ( \9937 , \9935 , \9936 );
xnor \U$9806 ( \9938 , \9937 , \1436 );
xor \U$9807 ( \9939 , \9934 , \9938 );
xor \U$9808 ( \9940 , \9925 , \9939 );
and \U$9809 ( \9941 , \6281 , \156 );
and \U$9810 ( \9942 , \6514 , \154 );
nor \U$9811 ( \9943 , \9941 , \9942 );
xnor \U$9812 ( \9944 , \9943 , \163 );
and \U$9813 ( \9945 , \5674 , \296 );
and \U$9814 ( \9946 , \6030 , \168 );
nor \U$9815 ( \9947 , \9945 , \9946 );
xnor \U$9816 ( \9948 , \9947 , \173 );
xor \U$9817 ( \9949 , \9944 , \9948 );
and \U$9818 ( \9950 , \5156 , \438 );
and \U$9819 ( \9951 , \5469 , \336 );
nor \U$9820 ( \9952 , \9950 , \9951 );
xnor \U$9821 ( \9953 , \9952 , \320 );
xor \U$9822 ( \9954 , \9949 , \9953 );
xor \U$9823 ( \9955 , \9940 , \9954 );
xor \U$9824 ( \9956 , \9911 , \9955 );
xor \U$9825 ( \9957 , \9891 , \9956 );
xor \U$9826 ( \9958 , \9862 , \9957 );
xor \U$9827 ( \9959 , \9693 , \9958 );
xor \U$9828 ( \9960 , \9684 , \9959 );
xor \U$9829 ( \9961 , \9665 , \9960 );
and \U$9830 ( \9962 , \9357 , \9381 );
and \U$9831 ( \9963 , \9381 , \9652 );
and \U$9832 ( \9964 , \9357 , \9652 );
or \U$9833 ( \9965 , \9962 , \9963 , \9964 );
xor \U$9834 ( \9966 , \9961 , \9965 );
and \U$9835 ( \9967 , \9653 , \9654 );
and \U$9836 ( \9968 , \9655 , \9658 );
or \U$9837 ( \9969 , \9967 , \9968 );
xor \U$9838 ( \9970 , \9966 , \9969 );
buf \U$9839 ( \9971 , \9970 );
buf \U$9840 ( \9972 , \9971 );
and \U$9841 ( \9973 , \9669 , \9683 );
and \U$9842 ( \9974 , \9683 , \9959 );
and \U$9843 ( \9975 , \9669 , \9959 );
or \U$9844 ( \9976 , \9973 , \9974 , \9975 );
and \U$9845 ( \9977 , \9688 , \9692 );
and \U$9846 ( \9978 , \9692 , \9958 );
and \U$9847 ( \9979 , \9688 , \9958 );
or \U$9848 ( \9980 , \9977 , \9978 , \9979 );
and \U$9849 ( \9981 , \9673 , \9677 );
and \U$9850 ( \9982 , \9677 , \9682 );
and \U$9851 ( \9983 , \9673 , \9682 );
or \U$9852 ( \9984 , \9981 , \9982 , \9983 );
and \U$9853 ( \9985 , \9707 , \9861 );
and \U$9854 ( \9986 , \9861 , \9957 );
and \U$9855 ( \9987 , \9707 , \9957 );
or \U$9856 ( \9988 , \9985 , \9986 , \9987 );
xor \U$9857 ( \9989 , \9984 , \9988 );
and \U$9858 ( \9990 , \9725 , \9739 );
and \U$9859 ( \9991 , \9739 , \9754 );
and \U$9860 ( \9992 , \9725 , \9754 );
or \U$9861 ( \9993 , \9990 , \9991 , \9992 );
and \U$9862 ( \9994 , \9770 , \9814 );
and \U$9863 ( \9995 , \9814 , \9859 );
and \U$9864 ( \9996 , \9770 , \9859 );
or \U$9865 ( \9997 , \9994 , \9995 , \9996 );
xor \U$9866 ( \9998 , \9993 , \9997 );
and \U$9867 ( \9999 , \9929 , \9933 );
and \U$9868 ( \10000 , \9933 , \9938 );
and \U$9869 ( \10001 , \9929 , \9938 );
or \U$9870 ( \10002 , \9999 , \10000 , \10001 );
and \U$9871 ( \10003 , \9788 , \9792 );
and \U$9872 ( \10004 , \9792 , \9797 );
and \U$9873 ( \10005 , \9788 , \9797 );
or \U$9874 ( \10006 , \10003 , \10004 , \10005 );
xor \U$9875 ( \10007 , \10002 , \10006 );
and \U$9876 ( \10008 , \9803 , \9807 );
and \U$9877 ( \10009 , \9807 , \9812 );
and \U$9878 ( \10010 , \9803 , \9812 );
or \U$9879 ( \10011 , \10008 , \10009 , \10010 );
xor \U$9880 ( \10012 , \10007 , \10011 );
xor \U$9881 ( \10013 , \9998 , \10012 );
xor \U$9882 ( \10014 , \9989 , \10013 );
xor \U$9883 ( \10015 , \9980 , \10014 );
and \U$9884 ( \10016 , \9866 , \9870 );
and \U$9885 ( \10017 , \9870 , \9875 );
and \U$9886 ( \10018 , \9866 , \9875 );
or \U$9887 ( \10019 , \10016 , \10017 , \10018 );
and \U$9888 ( \10020 , \9880 , \9884 );
and \U$9889 ( \10021 , \9884 , \9889 );
and \U$9890 ( \10022 , \9880 , \9889 );
or \U$9891 ( \10023 , \10020 , \10021 , \10022 );
xor \U$9892 ( \10024 , \10019 , \10023 );
and \U$9893 ( \10025 , \9895 , \9910 );
and \U$9894 ( \10026 , \9910 , \9955 );
and \U$9895 ( \10027 , \9895 , \9955 );
or \U$9896 ( \10028 , \10025 , \10026 , \10027 );
xor \U$9897 ( \10029 , \10024 , \10028 );
and \U$9898 ( \10030 , \9697 , \9701 );
and \U$9899 ( \10031 , \9701 , \9706 );
and \U$9900 ( \10032 , \9697 , \9706 );
or \U$9901 ( \10033 , \10030 , \10031 , \10032 );
and \U$9902 ( \10034 , \9711 , \9755 );
and \U$9903 ( \10035 , \9755 , \9860 );
and \U$9904 ( \10036 , \9711 , \9860 );
or \U$9905 ( \10037 , \10034 , \10035 , \10036 );
xor \U$9906 ( \10038 , \10033 , \10037 );
and \U$9907 ( \10039 , \9876 , \9890 );
and \U$9908 ( \10040 , \9890 , \9956 );
and \U$9909 ( \10041 , \9876 , \9956 );
or \U$9910 ( \10042 , \10039 , \10040 , \10041 );
xor \U$9911 ( \10043 , \10038 , \10042 );
xor \U$9912 ( \10044 , \10029 , \10043 );
and \U$9913 ( \10045 , \9715 , \9719 );
and \U$9914 ( \10046 , \9719 , \9724 );
and \U$9915 ( \10047 , \9715 , \9724 );
or \U$9916 ( \10048 , \10045 , \10046 , \10047 );
and \U$9917 ( \10049 , \9729 , \9733 );
and \U$9918 ( \10050 , \9733 , \9738 );
and \U$9919 ( \10051 , \9729 , \9738 );
or \U$9920 ( \10052 , \10049 , \10050 , \10051 );
xor \U$9921 ( \10053 , \10048 , \10052 );
and \U$9922 ( \10054 , \9744 , \9748 );
and \U$9923 ( \10055 , \9748 , \9753 );
and \U$9924 ( \10056 , \9744 , \9753 );
or \U$9925 ( \10057 , \10054 , \10055 , \10056 );
xor \U$9926 ( \10058 , \10053 , \10057 );
and \U$9927 ( \10059 , \9760 , \9761 );
and \U$9928 ( \10060 , \9761 , \9769 );
and \U$9929 ( \10061 , \9760 , \9769 );
or \U$9930 ( \10062 , \10059 , \10060 , \10061 );
and \U$9931 ( \10063 , \9784 , \9798 );
and \U$9932 ( \10064 , \9798 , \9813 );
and \U$9933 ( \10065 , \9784 , \9813 );
or \U$9934 ( \10066 , \10063 , \10064 , \10065 );
xor \U$9935 ( \10067 , \10062 , \10066 );
and \U$9936 ( \10068 , \9829 , \9843 );
and \U$9937 ( \10069 , \9843 , \9858 );
and \U$9938 ( \10070 , \9829 , \9858 );
or \U$9939 ( \10071 , \10068 , \10069 , \10070 );
xor \U$9940 ( \10072 , \10067 , \10071 );
xor \U$9941 ( \10073 , \10058 , \10072 );
and \U$9942 ( \10074 , \9915 , \9919 );
and \U$9943 ( \10075 , \9919 , \9924 );
and \U$9944 ( \10076 , \9915 , \9924 );
or \U$9945 ( \10077 , \10074 , \10075 , \10076 );
and \U$9946 ( \10078 , \9900 , \9904 );
and \U$9947 ( \10079 , \9904 , \9909 );
and \U$9948 ( \10080 , \9900 , \9909 );
or \U$9949 ( \10081 , \10078 , \10079 , \10080 );
xor \U$9950 ( \10082 , \10077 , \10081 );
and \U$9951 ( \10083 , \9944 , \9948 );
and \U$9952 ( \10084 , \9948 , \9953 );
and \U$9953 ( \10085 , \9944 , \9953 );
or \U$9954 ( \10086 , \10083 , \10084 , \10085 );
xor \U$9955 ( \10087 , \10082 , \10086 );
and \U$9956 ( \10088 , \9819 , \9823 );
and \U$9957 ( \10089 , \9823 , \9828 );
and \U$9958 ( \10090 , \9819 , \9828 );
or \U$9959 ( \10091 , \10088 , \10089 , \10090 );
and \U$9960 ( \10092 , \9833 , \9837 );
and \U$9961 ( \10093 , \9837 , \9842 );
and \U$9962 ( \10094 , \9833 , \9842 );
or \U$9963 ( \10095 , \10092 , \10093 , \10094 );
xor \U$9964 ( \10096 , \10091 , \10095 );
and \U$9965 ( \10097 , \9774 , \9778 );
and \U$9966 ( \10098 , \9778 , \9783 );
and \U$9967 ( \10099 , \9774 , \9783 );
or \U$9968 ( \10100 , \10097 , \10098 , \10099 );
xor \U$9969 ( \10101 , \10096 , \10100 );
and \U$9970 ( \10102 , \9848 , \9852 );
and \U$9971 ( \10103 , \9852 , \9857 );
and \U$9972 ( \10104 , \9848 , \9857 );
or \U$9973 ( \10105 , \10102 , \10103 , \10104 );
and \U$9974 ( \10106 , \134 , \9333 );
and \U$9975 ( \10107 , \143 , \9006 );
nor \U$9976 ( \10108 , \10106 , \10107 );
xnor \U$9977 ( \10109 , \10108 , \8848 );
and \U$9978 ( \10110 , \150 , \9765 );
and \U$9979 ( \10111 , \158 , \9644 );
nor \U$9980 ( \10112 , \10110 , \10111 );
xnor \U$9981 ( \10113 , \10112 , \9478 );
xor \U$9982 ( \10114 , \10109 , \10113 );
buf \U$9983 ( \10115 , RIb560f48_2);
xor \U$9984 ( \10116 , \10115 , \9474 );
nand \U$9985 ( \10117 , \166 , \10116 );
buf \U$9986 ( \10118 , RIb560fc0_1);
and \U$9987 ( \10119 , \10115 , \9474 );
not \U$9988 ( \10120 , \10119 );
and \U$9989 ( \10121 , \10118 , \10120 );
xnor \U$9990 ( \10122 , \10117 , \10121 );
xor \U$9991 ( \10123 , \10114 , \10122 );
xor \U$9992 ( \10124 , \10105 , \10123 );
and \U$9993 ( \10125 , \209 , \7489 );
and \U$9994 ( \10126 , \217 , \7137 );
nor \U$9995 ( \10127 , \10125 , \10126 );
xnor \U$9996 ( \10128 , \10127 , \7142 );
and \U$9997 ( \10129 , \224 , \8019 );
and \U$9998 ( \10130 , \232 , \7830 );
nor \U$9999 ( \10131 , \10129 , \10130 );
xnor \U$10000 ( \10132 , \10131 , \7713 );
xor \U$10001 ( \10133 , \10128 , \10132 );
and \U$10002 ( \10134 , \240 , \8540 );
and \U$10003 ( \10135 , \247 , \8292 );
nor \U$10004 ( \10136 , \10134 , \10135 );
xnor \U$10005 ( \10137 , \10136 , \8297 );
xor \U$10006 ( \10138 , \10133 , \10137 );
xor \U$10007 ( \10139 , \10124 , \10138 );
xor \U$10008 ( \10140 , \10101 , \10139 );
and \U$10009 ( \10141 , \1333 , \4581 );
and \U$10010 ( \10142 , \1484 , \4424 );
nor \U$10011 ( \10143 , \10141 , \10142 );
xnor \U$10012 ( \10144 , \10143 , \4377 );
and \U$10013 ( \10145 , \1147 , \5011 );
and \U$10014 ( \10146 , \1192 , \4878 );
nor \U$10015 ( \10147 , \10145 , \10146 );
xnor \U$10016 ( \10148 , \10147 , \4762 );
xor \U$10017 ( \10149 , \10144 , \10148 );
and \U$10018 ( \10150 , \412 , \5485 );
and \U$10019 ( \10151 , \474 , \5275 );
nor \U$10020 ( \10152 , \10150 , \10151 );
xnor \U$10021 ( \10153 , \10152 , \5169 );
xor \U$10022 ( \10154 , \10149 , \10153 );
and \U$10023 ( \10155 , \2090 , \3357 );
and \U$10024 ( \10156 , \2182 , \3255 );
nor \U$10025 ( \10157 , \10155 , \10156 );
xnor \U$10026 ( \10158 , \10157 , \3156 );
and \U$10027 ( \10159 , \1802 , \3813 );
and \U$10028 ( \10160 , \1948 , \3557 );
nor \U$10029 ( \10161 , \10159 , \10160 );
xnor \U$10030 ( \10162 , \10161 , \3562 );
xor \U$10031 ( \10163 , \10158 , \10162 );
and \U$10032 ( \10164 , \1601 , \4132 );
and \U$10033 ( \10165 , \1684 , \4012 );
nor \U$10034 ( \10166 , \10164 , \10165 );
xnor \U$10035 ( \10167 , \10166 , \3925 );
xor \U$10036 ( \10168 , \10163 , \10167 );
xor \U$10037 ( \10169 , \10154 , \10168 );
and \U$10038 ( \10170 , \261 , \5996 );
and \U$10039 ( \10171 , \307 , \5695 );
nor \U$10040 ( \10172 , \10170 , \10171 );
xnor \U$10041 ( \10173 , \10172 , \5687 );
and \U$10042 ( \10174 , \178 , \6401 );
and \U$10043 ( \10175 , \185 , \6143 );
nor \U$10044 ( \10176 , \10174 , \10175 );
xnor \U$10045 ( \10177 , \10176 , \6148 );
xor \U$10046 ( \10178 , \10173 , \10177 );
and \U$10047 ( \10179 , \189 , \7055 );
and \U$10048 ( \10180 , \197 , \6675 );
nor \U$10049 ( \10181 , \10179 , \10180 );
xnor \U$10050 ( \10182 , \10181 , \6680 );
xor \U$10051 ( \10183 , \10178 , \10182 );
xor \U$10052 ( \10184 , \10169 , \10183 );
xor \U$10053 ( \10185 , \10140 , \10184 );
xor \U$10054 ( \10186 , \10087 , \10185 );
and \U$10055 ( \10187 , \9925 , \9939 );
and \U$10056 ( \10188 , \9939 , \9954 );
and \U$10057 ( \10189 , \9925 , \9954 );
or \U$10058 ( \10190 , \10187 , \10188 , \10189 );
and \U$10059 ( \10191 , \6945 , \141 );
and \U$10060 ( \10192 , \7231 , \139 );
nor \U$10061 ( \10193 , \10191 , \10192 );
xnor \U$10062 ( \10194 , \10193 , \148 );
and \U$10063 ( \10195 , \6514 , \156 );
and \U$10064 ( \10196 , \6790 , \154 );
nor \U$10065 ( \10197 , \10195 , \10196 );
xnor \U$10066 ( \10198 , \10197 , \163 );
xor \U$10067 ( \10199 , \10194 , \10198 );
and \U$10068 ( \10200 , \6030 , \296 );
and \U$10069 ( \10201 , \6281 , \168 );
nor \U$10070 ( \10202 , \10200 , \10201 );
xnor \U$10071 ( \10203 , \10202 , \173 );
xor \U$10072 ( \10204 , \10199 , \10203 );
and \U$10073 ( \10205 , \9897 , \183 );
buf \U$10074 ( \10206 , RIb55f148_66);
and \U$10075 ( \10207 , \10206 , \180 );
nor \U$10076 ( \10208 , \10205 , \10207 );
xnor \U$10077 ( \10209 , \10208 , \179 );
and \U$10078 ( \10210 , \9169 , \195 );
and \U$10079 ( \10211 , \9465 , \193 );
nor \U$10080 ( \10212 , \10210 , \10211 );
xnor \U$10081 ( \10213 , \10212 , \202 );
xor \U$10082 ( \10214 , \10209 , \10213 );
xor \U$10083 ( \10215 , \10214 , \10121 );
xor \U$10084 ( \10216 , \10204 , \10215 );
and \U$10085 ( \10217 , \8652 , \215 );
and \U$10086 ( \10218 , \8835 , \213 );
nor \U$10087 ( \10219 , \10217 , \10218 );
xnor \U$10088 ( \10220 , \10219 , \222 );
and \U$10089 ( \10221 , \8057 , \230 );
and \U$10090 ( \10222 , \8349 , \228 );
nor \U$10091 ( \10223 , \10221 , \10222 );
xnor \U$10092 ( \10224 , \10223 , \237 );
xor \U$10093 ( \10225 , \10220 , \10224 );
and \U$10094 ( \10226 , \7556 , \245 );
and \U$10095 ( \10227 , \7700 , \243 );
nor \U$10096 ( \10228 , \10226 , \10227 );
xnor \U$10097 ( \10229 , \10228 , \252 );
xor \U$10098 ( \10230 , \10225 , \10229 );
xor \U$10099 ( \10231 , \10216 , \10230 );
xor \U$10100 ( \10232 , \10190 , \10231 );
and \U$10101 ( \10233 , \4160 , \1578 );
and \U$10102 ( \10234 , \4364 , \1431 );
nor \U$10103 ( \10235 , \10233 , \10234 );
xnor \U$10104 ( \10236 , \10235 , \1436 );
and \U$10105 ( \10237 , \3736 , \1824 );
and \U$10106 ( \10238 , \3912 , \1739 );
nor \U$10107 ( \10239 , \10237 , \10238 );
xnor \U$10108 ( \10240 , \10239 , \1697 );
xor \U$10109 ( \10241 , \10236 , \10240 );
and \U$10110 ( \10242 , \3395 , \2121 );
and \U$10111 ( \10243 , \3646 , \2008 );
nor \U$10112 ( \10244 , \10242 , \10243 );
xnor \U$10113 ( \10245 , \10244 , \1961 );
xor \U$10114 ( \10246 , \10241 , \10245 );
and \U$10115 ( \10247 , \5469 , \438 );
and \U$10116 ( \10248 , \5674 , \336 );
nor \U$10117 ( \10249 , \10247 , \10248 );
xnor \U$10118 ( \10250 , \10249 , \320 );
and \U$10119 ( \10251 , \4922 , \1086 );
and \U$10120 ( \10252 , \5156 , \508 );
nor \U$10121 ( \10253 , \10251 , \10252 );
xnor \U$10122 ( \10254 , \10253 , \487 );
xor \U$10123 ( \10255 , \10250 , \10254 );
and \U$10124 ( \10256 , \4654 , \1301 );
and \U$10125 ( \10257 , \4749 , \1246 );
nor \U$10126 ( \10258 , \10256 , \10257 );
xnor \U$10127 ( \10259 , \10258 , \1205 );
xor \U$10128 ( \10260 , \10255 , \10259 );
xor \U$10129 ( \10261 , \10246 , \10260 );
and \U$10130 ( \10262 , \3037 , \2400 );
and \U$10131 ( \10263 , \3143 , \2246 );
nor \U$10132 ( \10264 , \10262 , \10263 );
xnor \U$10133 ( \10265 , \10264 , \2195 );
and \U$10134 ( \10266 , \2757 , \2669 );
and \U$10135 ( \10267 , \2826 , \2538 );
nor \U$10136 ( \10268 , \10266 , \10267 );
xnor \U$10137 ( \10269 , \10268 , \2534 );
xor \U$10138 ( \10270 , \10265 , \10269 );
and \U$10139 ( \10271 , \2366 , \3103 );
and \U$10140 ( \10272 , \2521 , \2934 );
nor \U$10141 ( \10273 , \10271 , \10272 );
xnor \U$10142 ( \10274 , \10273 , \2839 );
xor \U$10143 ( \10275 , \10270 , \10274 );
xor \U$10144 ( \10276 , \10261 , \10275 );
xor \U$10145 ( \10277 , \10232 , \10276 );
xor \U$10146 ( \10278 , \10186 , \10277 );
xor \U$10147 ( \10279 , \10073 , \10278 );
xor \U$10148 ( \10280 , \10044 , \10279 );
xor \U$10149 ( \10281 , \10015 , \10280 );
xor \U$10150 ( \10282 , \9976 , \10281 );
and \U$10151 ( \10283 , \9665 , \9960 );
xor \U$10152 ( \10284 , \10282 , \10283 );
and \U$10153 ( \10285 , \9961 , \9965 );
and \U$10154 ( \10286 , \9966 , \9969 );
or \U$10155 ( \10287 , \10285 , \10286 );
xor \U$10156 ( \10288 , \10284 , \10287 );
buf \U$10157 ( \10289 , \10288 );
buf \U$10158 ( \10290 , \10289 );
and \U$10159 ( \10291 , \9980 , \10014 );
and \U$10160 ( \10292 , \10014 , \10280 );
and \U$10161 ( \10293 , \9980 , \10280 );
or \U$10162 ( \10294 , \10291 , \10292 , \10293 );
and \U$10163 ( \10295 , \9984 , \9988 );
and \U$10164 ( \10296 , \9988 , \10013 );
and \U$10165 ( \10297 , \9984 , \10013 );
or \U$10166 ( \10298 , \10295 , \10296 , \10297 );
and \U$10167 ( \10299 , \10029 , \10043 );
and \U$10168 ( \10300 , \10043 , \10279 );
and \U$10169 ( \10301 , \10029 , \10279 );
or \U$10170 ( \10302 , \10299 , \10300 , \10301 );
xor \U$10171 ( \10303 , \10298 , \10302 );
and \U$10172 ( \10304 , \10019 , \10023 );
and \U$10173 ( \10305 , \10023 , \10028 );
and \U$10174 ( \10306 , \10019 , \10028 );
or \U$10175 ( \10307 , \10304 , \10305 , \10306 );
and \U$10176 ( \10308 , \9993 , \9997 );
and \U$10177 ( \10309 , \9997 , \10012 );
and \U$10178 ( \10310 , \9993 , \10012 );
or \U$10179 ( \10311 , \10308 , \10309 , \10310 );
xor \U$10180 ( \10312 , \10307 , \10311 );
and \U$10181 ( \10313 , \10087 , \10185 );
and \U$10182 ( \10314 , \10185 , \10277 );
and \U$10183 ( \10315 , \10087 , \10277 );
or \U$10184 ( \10316 , \10313 , \10314 , \10315 );
xor \U$10185 ( \10317 , \10312 , \10316 );
xor \U$10186 ( \10318 , \10303 , \10317 );
xor \U$10187 ( \10319 , \10294 , \10318 );
and \U$10188 ( \10320 , \10033 , \10037 );
and \U$10189 ( \10321 , \10037 , \10042 );
and \U$10190 ( \10322 , \10033 , \10042 );
or \U$10191 ( \10323 , \10320 , \10321 , \10322 );
and \U$10192 ( \10324 , \10058 , \10072 );
and \U$10193 ( \10325 , \10072 , \10278 );
and \U$10194 ( \10326 , \10058 , \10278 );
or \U$10195 ( \10327 , \10324 , \10325 , \10326 );
xor \U$10196 ( \10328 , \10323 , \10327 );
and \U$10197 ( \10329 , \10048 , \10052 );
and \U$10198 ( \10330 , \10052 , \10057 );
and \U$10199 ( \10331 , \10048 , \10057 );
or \U$10200 ( \10332 , \10329 , \10330 , \10331 );
and \U$10201 ( \10333 , \10062 , \10066 );
and \U$10202 ( \10334 , \10066 , \10071 );
and \U$10203 ( \10335 , \10062 , \10071 );
or \U$10204 ( \10336 , \10333 , \10334 , \10335 );
xor \U$10205 ( \10337 , \10332 , \10336 );
and \U$10206 ( \10338 , \10190 , \10231 );
and \U$10207 ( \10339 , \10231 , \10276 );
and \U$10208 ( \10340 , \10190 , \10276 );
or \U$10209 ( \10341 , \10338 , \10339 , \10340 );
xor \U$10210 ( \10342 , \10337 , \10341 );
and \U$10211 ( \10343 , \10101 , \10139 );
and \U$10212 ( \10344 , \10139 , \10184 );
and \U$10213 ( \10345 , \10101 , \10184 );
or \U$10214 ( \10346 , \10343 , \10344 , \10345 );
and \U$10215 ( \10347 , \10144 , \10148 );
and \U$10216 ( \10348 , \10148 , \10153 );
and \U$10217 ( \10349 , \10144 , \10153 );
or \U$10218 ( \10350 , \10347 , \10348 , \10349 );
and \U$10219 ( \10351 , \10158 , \10162 );
and \U$10220 ( \10352 , \10162 , \10167 );
and \U$10221 ( \10353 , \10158 , \10167 );
or \U$10222 ( \10354 , \10351 , \10352 , \10353 );
xor \U$10223 ( \10355 , \10350 , \10354 );
and \U$10224 ( \10356 , \10173 , \10177 );
and \U$10225 ( \10357 , \10177 , \10182 );
and \U$10226 ( \10358 , \10173 , \10182 );
or \U$10227 ( \10359 , \10356 , \10357 , \10358 );
xor \U$10228 ( \10360 , \10355 , \10359 );
and \U$10229 ( \10361 , \10194 , \10198 );
and \U$10230 ( \10362 , \10198 , \10203 );
and \U$10231 ( \10363 , \10194 , \10203 );
or \U$10232 ( \10364 , \10361 , \10362 , \10363 );
and \U$10233 ( \10365 , \10209 , \10213 );
and \U$10234 ( \10366 , \10213 , \10121 );
and \U$10235 ( \10367 , \10209 , \10121 );
or \U$10236 ( \10368 , \10365 , \10366 , \10367 );
xor \U$10237 ( \10369 , \10364 , \10368 );
and \U$10238 ( \10370 , \10220 , \10224 );
and \U$10239 ( \10371 , \10224 , \10229 );
and \U$10240 ( \10372 , \10220 , \10229 );
or \U$10241 ( \10373 , \10370 , \10371 , \10372 );
xor \U$10242 ( \10374 , \10369 , \10373 );
xor \U$10243 ( \10375 , \10360 , \10374 );
and \U$10244 ( \10376 , \10236 , \10240 );
and \U$10245 ( \10377 , \10240 , \10245 );
and \U$10246 ( \10378 , \10236 , \10245 );
or \U$10247 ( \10379 , \10376 , \10377 , \10378 );
and \U$10248 ( \10380 , \10250 , \10254 );
and \U$10249 ( \10381 , \10254 , \10259 );
and \U$10250 ( \10382 , \10250 , \10259 );
or \U$10251 ( \10383 , \10380 , \10381 , \10382 );
xor \U$10252 ( \10384 , \10379 , \10383 );
and \U$10253 ( \10385 , \10265 , \10269 );
and \U$10254 ( \10386 , \10269 , \10274 );
and \U$10255 ( \10387 , \10265 , \10274 );
or \U$10256 ( \10388 , \10385 , \10386 , \10387 );
xor \U$10257 ( \10389 , \10384 , \10388 );
xor \U$10258 ( \10390 , \10375 , \10389 );
xor \U$10259 ( \10391 , \10346 , \10390 );
and \U$10260 ( \10392 , \10109 , \10113 );
and \U$10261 ( \10393 , \10113 , \10122 );
and \U$10262 ( \10394 , \10109 , \10122 );
or \U$10263 ( \10395 , \10392 , \10393 , \10394 );
and \U$10264 ( \10396 , \10128 , \10132 );
and \U$10265 ( \10397 , \10132 , \10137 );
and \U$10266 ( \10398 , \10128 , \10137 );
or \U$10267 ( \10399 , \10396 , \10397 , \10398 );
xor \U$10268 ( \10400 , \10395 , \10399 );
and \U$10269 ( \10401 , \158 , \9765 );
and \U$10270 ( \10402 , \134 , \9644 );
nor \U$10271 ( \10403 , \10401 , \10402 );
xnor \U$10272 ( \10404 , \10403 , \9478 );
xor \U$10273 ( \10405 , \10400 , \10404 );
xor \U$10274 ( \10406 , \10118 , \10115 );
not \U$10275 ( \10407 , \10116 );
and \U$10276 ( \10408 , \10406 , \10407 );
and \U$10277 ( \10409 , \166 , \10408 );
and \U$10278 ( \10410 , \150 , \10116 );
nor \U$10279 ( \10411 , \10409 , \10410 );
xnor \U$10280 ( \10412 , \10411 , \10121 );
and \U$10281 ( \10413 , \185 , \6401 );
and \U$10282 ( \10414 , \261 , \6143 );
nor \U$10283 ( \10415 , \10413 , \10414 );
xnor \U$10284 ( \10416 , \10415 , \6148 );
and \U$10285 ( \10417 , \197 , \7055 );
and \U$10286 ( \10418 , \178 , \6675 );
nor \U$10287 ( \10419 , \10417 , \10418 );
xnor \U$10288 ( \10420 , \10419 , \6680 );
xor \U$10289 ( \10421 , \10416 , \10420 );
and \U$10290 ( \10422 , \217 , \7489 );
and \U$10291 ( \10423 , \189 , \7137 );
nor \U$10292 ( \10424 , \10422 , \10423 );
xnor \U$10293 ( \10425 , \10424 , \7142 );
xor \U$10294 ( \10426 , \10421 , \10425 );
xor \U$10295 ( \10427 , \10412 , \10426 );
and \U$10296 ( \10428 , \232 , \8019 );
and \U$10297 ( \10429 , \209 , \7830 );
nor \U$10298 ( \10430 , \10428 , \10429 );
xnor \U$10299 ( \10431 , \10430 , \7713 );
and \U$10300 ( \10432 , \247 , \8540 );
and \U$10301 ( \10433 , \224 , \8292 );
nor \U$10302 ( \10434 , \10432 , \10433 );
xnor \U$10303 ( \10435 , \10434 , \8297 );
xor \U$10304 ( \10436 , \10431 , \10435 );
and \U$10305 ( \10437 , \143 , \9333 );
and \U$10306 ( \10438 , \240 , \9006 );
nor \U$10307 ( \10439 , \10437 , \10438 );
xnor \U$10308 ( \10440 , \10439 , \8848 );
xor \U$10309 ( \10441 , \10436 , \10440 );
xor \U$10310 ( \10442 , \10427 , \10441 );
xor \U$10311 ( \10443 , \10405 , \10442 );
and \U$10312 ( \10444 , \1192 , \5011 );
and \U$10313 ( \10445 , \1333 , \4878 );
nor \U$10314 ( \10446 , \10444 , \10445 );
xnor \U$10315 ( \10447 , \10446 , \4762 );
and \U$10316 ( \10448 , \474 , \5485 );
and \U$10317 ( \10449 , \1147 , \5275 );
nor \U$10318 ( \10450 , \10448 , \10449 );
xnor \U$10319 ( \10451 , \10450 , \5169 );
xor \U$10320 ( \10452 , \10447 , \10451 );
and \U$10321 ( \10453 , \307 , \5996 );
and \U$10322 ( \10454 , \412 , \5695 );
nor \U$10323 ( \10455 , \10453 , \10454 );
xnor \U$10324 ( \10456 , \10455 , \5687 );
xor \U$10325 ( \10457 , \10452 , \10456 );
and \U$10326 ( \10458 , \1948 , \3813 );
and \U$10327 ( \10459 , \2090 , \3557 );
nor \U$10328 ( \10460 , \10458 , \10459 );
xnor \U$10329 ( \10461 , \10460 , \3562 );
and \U$10330 ( \10462 , \1684 , \4132 );
and \U$10331 ( \10463 , \1802 , \4012 );
nor \U$10332 ( \10464 , \10462 , \10463 );
xnor \U$10333 ( \10465 , \10464 , \3925 );
xor \U$10334 ( \10466 , \10461 , \10465 );
and \U$10335 ( \10467 , \1484 , \4581 );
and \U$10336 ( \10468 , \1601 , \4424 );
nor \U$10337 ( \10469 , \10467 , \10468 );
xnor \U$10338 ( \10470 , \10469 , \4377 );
xor \U$10339 ( \10471 , \10466 , \10470 );
xor \U$10340 ( \10472 , \10457 , \10471 );
and \U$10341 ( \10473 , \2826 , \2669 );
and \U$10342 ( \10474 , \3037 , \2538 );
nor \U$10343 ( \10475 , \10473 , \10474 );
xnor \U$10344 ( \10476 , \10475 , \2534 );
and \U$10345 ( \10477 , \2521 , \3103 );
and \U$10346 ( \10478 , \2757 , \2934 );
nor \U$10347 ( \10479 , \10477 , \10478 );
xnor \U$10348 ( \10480 , \10479 , \2839 );
xor \U$10349 ( \10481 , \10476 , \10480 );
and \U$10350 ( \10482 , \2182 , \3357 );
and \U$10351 ( \10483 , \2366 , \3255 );
nor \U$10352 ( \10484 , \10482 , \10483 );
xnor \U$10353 ( \10485 , \10484 , \3156 );
xor \U$10354 ( \10486 , \10481 , \10485 );
xor \U$10355 ( \10487 , \10472 , \10486 );
xor \U$10356 ( \10488 , \10443 , \10487 );
xor \U$10357 ( \10489 , \10391 , \10488 );
xor \U$10358 ( \10490 , \10342 , \10489 );
and \U$10359 ( \10491 , \10077 , \10081 );
and \U$10360 ( \10492 , \10081 , \10086 );
and \U$10361 ( \10493 , \10077 , \10086 );
or \U$10362 ( \10494 , \10491 , \10492 , \10493 );
and \U$10363 ( \10495 , \10091 , \10095 );
and \U$10364 ( \10496 , \10095 , \10100 );
and \U$10365 ( \10497 , \10091 , \10100 );
or \U$10366 ( \10498 , \10495 , \10496 , \10497 );
xor \U$10367 ( \10499 , \10494 , \10498 );
and \U$10368 ( \10500 , \10002 , \10006 );
and \U$10369 ( \10501 , \10006 , \10011 );
and \U$10370 ( \10502 , \10002 , \10011 );
or \U$10371 ( \10503 , \10500 , \10501 , \10502 );
xor \U$10372 ( \10504 , \10499 , \10503 );
and \U$10373 ( \10505 , \10246 , \10260 );
and \U$10374 ( \10506 , \10260 , \10275 );
and \U$10375 ( \10507 , \10246 , \10275 );
or \U$10376 ( \10508 , \10505 , \10506 , \10507 );
and \U$10377 ( \10509 , \10105 , \10123 );
and \U$10378 ( \10510 , \10123 , \10138 );
and \U$10379 ( \10511 , \10105 , \10138 );
or \U$10380 ( \10512 , \10509 , \10510 , \10511 );
xor \U$10381 ( \10513 , \10508 , \10512 );
and \U$10382 ( \10514 , \10154 , \10168 );
and \U$10383 ( \10515 , \10168 , \10183 );
and \U$10384 ( \10516 , \10154 , \10183 );
or \U$10385 ( \10517 , \10514 , \10515 , \10516 );
xor \U$10386 ( \10518 , \10513 , \10517 );
xor \U$10387 ( \10519 , \10504 , \10518 );
and \U$10388 ( \10520 , \10204 , \10215 );
and \U$10389 ( \10521 , \10215 , \10230 );
and \U$10390 ( \10522 , \10204 , \10230 );
or \U$10391 ( \10523 , \10520 , \10521 , \10522 );
and \U$10392 ( \10524 , \3912 , \1824 );
and \U$10393 ( \10525 , \4160 , \1739 );
nor \U$10394 ( \10526 , \10524 , \10525 );
xnor \U$10395 ( \10527 , \10526 , \1697 );
and \U$10396 ( \10528 , \3646 , \2121 );
and \U$10397 ( \10529 , \3736 , \2008 );
nor \U$10398 ( \10530 , \10528 , \10529 );
xnor \U$10399 ( \10531 , \10530 , \1961 );
xor \U$10400 ( \10532 , \10527 , \10531 );
and \U$10401 ( \10533 , \3143 , \2400 );
and \U$10402 ( \10534 , \3395 , \2246 );
nor \U$10403 ( \10535 , \10533 , \10534 );
xnor \U$10404 ( \10536 , \10535 , \2195 );
xor \U$10405 ( \10537 , \10532 , \10536 );
and \U$10406 ( \10538 , \5156 , \1086 );
and \U$10407 ( \10539 , \5469 , \508 );
nor \U$10408 ( \10540 , \10538 , \10539 );
xnor \U$10409 ( \10541 , \10540 , \487 );
and \U$10410 ( \10542 , \4749 , \1301 );
and \U$10411 ( \10543 , \4922 , \1246 );
nor \U$10412 ( \10544 , \10542 , \10543 );
xnor \U$10413 ( \10545 , \10544 , \1205 );
xor \U$10414 ( \10546 , \10541 , \10545 );
and \U$10415 ( \10547 , \4364 , \1578 );
and \U$10416 ( \10548 , \4654 , \1431 );
nor \U$10417 ( \10549 , \10547 , \10548 );
xnor \U$10418 ( \10550 , \10549 , \1436 );
xor \U$10419 ( \10551 , \10546 , \10550 );
xor \U$10420 ( \10552 , \10537 , \10551 );
and \U$10421 ( \10553 , \6790 , \156 );
and \U$10422 ( \10554 , \6945 , \154 );
nor \U$10423 ( \10555 , \10553 , \10554 );
xnor \U$10424 ( \10556 , \10555 , \163 );
and \U$10425 ( \10557 , \6281 , \296 );
and \U$10426 ( \10558 , \6514 , \168 );
nor \U$10427 ( \10559 , \10557 , \10558 );
xnor \U$10428 ( \10560 , \10559 , \173 );
xor \U$10429 ( \10561 , \10556 , \10560 );
and \U$10430 ( \10562 , \5674 , \438 );
and \U$10431 ( \10563 , \6030 , \336 );
nor \U$10432 ( \10564 , \10562 , \10563 );
xnor \U$10433 ( \10565 , \10564 , \320 );
xor \U$10434 ( \10566 , \10561 , \10565 );
xor \U$10435 ( \10567 , \10552 , \10566 );
xor \U$10436 ( \10568 , \10523 , \10567 );
and \U$10437 ( \10569 , \8349 , \230 );
and \U$10438 ( \10570 , \8652 , \228 );
nor \U$10439 ( \10571 , \10569 , \10570 );
xnor \U$10440 ( \10572 , \10571 , \237 );
and \U$10441 ( \10573 , \7700 , \245 );
and \U$10442 ( \10574 , \8057 , \243 );
nor \U$10443 ( \10575 , \10573 , \10574 );
xnor \U$10444 ( \10576 , \10575 , \252 );
xor \U$10445 ( \10577 , \10572 , \10576 );
and \U$10446 ( \10578 , \7231 , \141 );
and \U$10447 ( \10579 , \7556 , \139 );
nor \U$10448 ( \10580 , \10578 , \10579 );
xnor \U$10449 ( \10581 , \10580 , \148 );
xor \U$10450 ( \10582 , \10577 , \10581 );
and \U$10451 ( \10583 , \10206 , \183 );
buf \U$10452 ( \10584 , RIb55f1c0_65);
and \U$10453 ( \10585 , \10584 , \180 );
nor \U$10454 ( \10586 , \10583 , \10585 );
xnor \U$10455 ( \10587 , \10586 , \179 );
and \U$10456 ( \10588 , \9465 , \195 );
and \U$10457 ( \10589 , \9897 , \193 );
nor \U$10458 ( \10590 , \10588 , \10589 );
xnor \U$10459 ( \10591 , \10590 , \202 );
xor \U$10460 ( \10592 , \10587 , \10591 );
and \U$10461 ( \10593 , \8835 , \215 );
and \U$10462 ( \10594 , \9169 , \213 );
nor \U$10463 ( \10595 , \10593 , \10594 );
xnor \U$10464 ( \10596 , \10595 , \222 );
xor \U$10465 ( \10597 , \10592 , \10596 );
xor \U$10466 ( \10598 , \10582 , \10597 );
xor \U$10467 ( \10599 , \10568 , \10598 );
xor \U$10468 ( \10600 , \10519 , \10599 );
xor \U$10469 ( \10601 , \10490 , \10600 );
xor \U$10470 ( \10602 , \10328 , \10601 );
xor \U$10471 ( \10603 , \10319 , \10602 );
and \U$10472 ( \10604 , \9976 , \10281 );
xor \U$10473 ( \10605 , \10603 , \10604 );
and \U$10474 ( \10606 , \10282 , \10283 );
and \U$10475 ( \10607 , \10284 , \10287 );
or \U$10476 ( \10608 , \10606 , \10607 );
xor \U$10477 ( \10609 , \10605 , \10608 );
buf \U$10478 ( \10610 , \10609 );
buf \U$10479 ( \10611 , \10610 );
and \U$10480 ( \10612 , \10298 , \10302 );
and \U$10481 ( \10613 , \10302 , \10317 );
and \U$10482 ( \10614 , \10298 , \10317 );
or \U$10483 ( \10615 , \10612 , \10613 , \10614 );
and \U$10484 ( \10616 , \10323 , \10327 );
and \U$10485 ( \10617 , \10327 , \10601 );
and \U$10486 ( \10618 , \10323 , \10601 );
or \U$10487 ( \10619 , \10616 , \10617 , \10618 );
and \U$10488 ( \10620 , \10307 , \10311 );
and \U$10489 ( \10621 , \10311 , \10316 );
and \U$10490 ( \10622 , \10307 , \10316 );
or \U$10491 ( \10623 , \10620 , \10621 , \10622 );
and \U$10492 ( \10624 , \10342 , \10489 );
and \U$10493 ( \10625 , \10489 , \10600 );
and \U$10494 ( \10626 , \10342 , \10600 );
or \U$10495 ( \10627 , \10624 , \10625 , \10626 );
xor \U$10496 ( \10628 , \10623 , \10627 );
and \U$10497 ( \10629 , \10360 , \10374 );
and \U$10498 ( \10630 , \10374 , \10389 );
and \U$10499 ( \10631 , \10360 , \10389 );
or \U$10500 ( \10632 , \10629 , \10630 , \10631 );
and \U$10501 ( \10633 , \10405 , \10442 );
and \U$10502 ( \10634 , \10442 , \10487 );
and \U$10503 ( \10635 , \10405 , \10487 );
or \U$10504 ( \10636 , \10633 , \10634 , \10635 );
xor \U$10505 ( \10637 , \10632 , \10636 );
and \U$10506 ( \10638 , \10556 , \10560 );
and \U$10507 ( \10639 , \10560 , \10565 );
and \U$10508 ( \10640 , \10556 , \10565 );
or \U$10509 ( \10641 , \10638 , \10639 , \10640 );
and \U$10510 ( \10642 , \10572 , \10576 );
and \U$10511 ( \10643 , \10576 , \10581 );
and \U$10512 ( \10644 , \10572 , \10581 );
or \U$10513 ( \10645 , \10642 , \10643 , \10644 );
xor \U$10514 ( \10646 , \10641 , \10645 );
and \U$10515 ( \10647 , \10587 , \10591 );
and \U$10516 ( \10648 , \10591 , \10596 );
and \U$10517 ( \10649 , \10587 , \10596 );
or \U$10518 ( \10650 , \10647 , \10648 , \10649 );
xor \U$10519 ( \10651 , \10646 , \10650 );
xor \U$10520 ( \10652 , \10637 , \10651 );
xor \U$10521 ( \10653 , \10628 , \10652 );
xor \U$10522 ( \10654 , \10619 , \10653 );
and \U$10523 ( \10655 , \10494 , \10498 );
and \U$10524 ( \10656 , \10498 , \10503 );
and \U$10525 ( \10657 , \10494 , \10503 );
or \U$10526 ( \10658 , \10655 , \10656 , \10657 );
and \U$10527 ( \10659 , \10508 , \10512 );
and \U$10528 ( \10660 , \10512 , \10517 );
and \U$10529 ( \10661 , \10508 , \10517 );
or \U$10530 ( \10662 , \10659 , \10660 , \10661 );
xor \U$10531 ( \10663 , \10658 , \10662 );
and \U$10532 ( \10664 , \10523 , \10567 );
and \U$10533 ( \10665 , \10567 , \10598 );
and \U$10534 ( \10666 , \10523 , \10598 );
or \U$10535 ( \10667 , \10664 , \10665 , \10666 );
xor \U$10536 ( \10668 , \10663 , \10667 );
and \U$10537 ( \10669 , \10332 , \10336 );
and \U$10538 ( \10670 , \10336 , \10341 );
and \U$10539 ( \10671 , \10332 , \10341 );
or \U$10540 ( \10672 , \10669 , \10670 , \10671 );
and \U$10541 ( \10673 , \10346 , \10390 );
and \U$10542 ( \10674 , \10390 , \10488 );
and \U$10543 ( \10675 , \10346 , \10488 );
or \U$10544 ( \10676 , \10673 , \10674 , \10675 );
xor \U$10545 ( \10677 , \10672 , \10676 );
and \U$10546 ( \10678 , \10504 , \10518 );
and \U$10547 ( \10679 , \10518 , \10599 );
and \U$10548 ( \10680 , \10504 , \10599 );
or \U$10549 ( \10681 , \10678 , \10679 , \10680 );
xor \U$10550 ( \10682 , \10677 , \10681 );
xor \U$10551 ( \10683 , \10668 , \10682 );
and \U$10552 ( \10684 , \10395 , \10399 );
and \U$10553 ( \10685 , \10399 , \10404 );
and \U$10554 ( \10686 , \10395 , \10404 );
or \U$10555 ( \10687 , \10684 , \10685 , \10686 );
and \U$10556 ( \10688 , \10412 , \10426 );
and \U$10557 ( \10689 , \10426 , \10441 );
and \U$10558 ( \10690 , \10412 , \10441 );
or \U$10559 ( \10691 , \10688 , \10689 , \10690 );
xor \U$10560 ( \10692 , \10687 , \10691 );
and \U$10561 ( \10693 , \10457 , \10471 );
and \U$10562 ( \10694 , \10471 , \10486 );
and \U$10563 ( \10695 , \10457 , \10486 );
or \U$10564 ( \10696 , \10693 , \10694 , \10695 );
xor \U$10565 ( \10697 , \10692 , \10696 );
and \U$10566 ( \10698 , \10350 , \10354 );
and \U$10567 ( \10699 , \10354 , \10359 );
and \U$10568 ( \10700 , \10350 , \10359 );
or \U$10569 ( \10701 , \10698 , \10699 , \10700 );
and \U$10570 ( \10702 , \10364 , \10368 );
and \U$10571 ( \10703 , \10368 , \10373 );
and \U$10572 ( \10704 , \10364 , \10373 );
or \U$10573 ( \10705 , \10702 , \10703 , \10704 );
xor \U$10574 ( \10706 , \10701 , \10705 );
and \U$10575 ( \10707 , \10379 , \10383 );
and \U$10576 ( \10708 , \10383 , \10388 );
and \U$10577 ( \10709 , \10379 , \10388 );
or \U$10578 ( \10710 , \10707 , \10708 , \10709 );
xor \U$10579 ( \10711 , \10706 , \10710 );
xor \U$10580 ( \10712 , \10697 , \10711 );
and \U$10581 ( \10713 , \10527 , \10531 );
and \U$10582 ( \10714 , \10531 , \10536 );
and \U$10583 ( \10715 , \10527 , \10536 );
or \U$10584 ( \10716 , \10713 , \10714 , \10715 );
and \U$10585 ( \10717 , \10541 , \10545 );
and \U$10586 ( \10718 , \10545 , \10550 );
and \U$10587 ( \10719 , \10541 , \10550 );
or \U$10588 ( \10720 , \10717 , \10718 , \10719 );
xor \U$10589 ( \10721 , \10716 , \10720 );
and \U$10590 ( \10722 , \10476 , \10480 );
and \U$10591 ( \10723 , \10480 , \10485 );
and \U$10592 ( \10724 , \10476 , \10485 );
or \U$10593 ( \10725 , \10722 , \10723 , \10724 );
xor \U$10594 ( \10726 , \10721 , \10725 );
and \U$10595 ( \10727 , \10447 , \10451 );
and \U$10596 ( \10728 , \10451 , \10456 );
and \U$10597 ( \10729 , \10447 , \10456 );
or \U$10598 ( \10730 , \10727 , \10728 , \10729 );
and \U$10599 ( \10731 , \10461 , \10465 );
and \U$10600 ( \10732 , \10465 , \10470 );
and \U$10601 ( \10733 , \10461 , \10470 );
or \U$10602 ( \10734 , \10731 , \10732 , \10733 );
xor \U$10603 ( \10735 , \10730 , \10734 );
and \U$10604 ( \10736 , \10416 , \10420 );
and \U$10605 ( \10737 , \10420 , \10425 );
and \U$10606 ( \10738 , \10416 , \10425 );
or \U$10607 ( \10739 , \10736 , \10737 , \10738 );
xor \U$10608 ( \10740 , \10735 , \10739 );
xor \U$10609 ( \10741 , \10726 , \10740 );
and \U$10610 ( \10742 , \10431 , \10435 );
and \U$10611 ( \10743 , \10435 , \10440 );
and \U$10612 ( \10744 , \10431 , \10440 );
or \U$10613 ( \10745 , \10742 , \10743 , \10744 );
nand \U$10614 ( \10746 , \166 , \10118 );
not \U$10615 ( \10747 , \10746 );
xor \U$10616 ( \10748 , \10745 , \10747 );
and \U$10617 ( \10749 , \240 , \9333 );
and \U$10618 ( \10750 , \247 , \9006 );
nor \U$10619 ( \10751 , \10749 , \10750 );
xnor \U$10620 ( \10752 , \10751 , \8848 );
and \U$10621 ( \10753 , \134 , \9765 );
and \U$10622 ( \10754 , \143 , \9644 );
nor \U$10623 ( \10755 , \10753 , \10754 );
xnor \U$10624 ( \10756 , \10755 , \9478 );
xor \U$10625 ( \10757 , \10752 , \10756 );
and \U$10626 ( \10758 , \150 , \10408 );
and \U$10627 ( \10759 , \158 , \10116 );
nor \U$10628 ( \10760 , \10758 , \10759 );
xnor \U$10629 ( \10761 , \10760 , \10121 );
xor \U$10630 ( \10762 , \10757 , \10761 );
xor \U$10631 ( \10763 , \10748 , \10762 );
xor \U$10632 ( \10764 , \10741 , \10763 );
and \U$10633 ( \10765 , \9169 , \215 );
and \U$10634 ( \10766 , \9465 , \213 );
nor \U$10635 ( \10767 , \10765 , \10766 );
xnor \U$10636 ( \10768 , \10767 , \222 );
and \U$10637 ( \10769 , \8652 , \230 );
and \U$10638 ( \10770 , \8835 , \228 );
nor \U$10639 ( \10771 , \10769 , \10770 );
xnor \U$10640 ( \10772 , \10771 , \237 );
xor \U$10641 ( \10773 , \10768 , \10772 );
and \U$10642 ( \10774 , \8057 , \245 );
and \U$10643 ( \10775 , \8349 , \243 );
nor \U$10644 ( \10776 , \10774 , \10775 );
xnor \U$10645 ( \10777 , \10776 , \252 );
xor \U$10646 ( \10778 , \10773 , \10777 );
and \U$10647 ( \10779 , \7556 , \141 );
and \U$10648 ( \10780 , \7700 , \139 );
nor \U$10649 ( \10781 , \10779 , \10780 );
xnor \U$10650 ( \10782 , \10781 , \148 );
and \U$10651 ( \10783 , \6945 , \156 );
and \U$10652 ( \10784 , \7231 , \154 );
nor \U$10653 ( \10785 , \10783 , \10784 );
xnor \U$10654 ( \10786 , \10785 , \163 );
xor \U$10655 ( \10787 , \10782 , \10786 );
and \U$10656 ( \10788 , \6514 , \296 );
and \U$10657 ( \10789 , \6790 , \168 );
nor \U$10658 ( \10790 , \10788 , \10789 );
xnor \U$10659 ( \10791 , \10790 , \173 );
xor \U$10660 ( \10792 , \10787 , \10791 );
xor \U$10661 ( \10793 , \10778 , \10792 );
and \U$10662 ( \10794 , \6030 , \438 );
and \U$10663 ( \10795 , \6281 , \336 );
nor \U$10664 ( \10796 , \10794 , \10795 );
xnor \U$10665 ( \10797 , \10796 , \320 );
and \U$10666 ( \10798 , \5469 , \1086 );
and \U$10667 ( \10799 , \5674 , \508 );
nor \U$10668 ( \10800 , \10798 , \10799 );
xnor \U$10669 ( \10801 , \10800 , \487 );
xor \U$10670 ( \10802 , \10797 , \10801 );
and \U$10671 ( \10803 , \4922 , \1301 );
and \U$10672 ( \10804 , \5156 , \1246 );
nor \U$10673 ( \10805 , \10803 , \10804 );
xnor \U$10674 ( \10806 , \10805 , \1205 );
xor \U$10675 ( \10807 , \10802 , \10806 );
xor \U$10676 ( \10808 , \10793 , \10807 );
and \U$10677 ( \10809 , \1601 , \4581 );
and \U$10678 ( \10810 , \1684 , \4424 );
nor \U$10679 ( \10811 , \10809 , \10810 );
xnor \U$10680 ( \10812 , \10811 , \4377 );
and \U$10681 ( \10813 , \1333 , \5011 );
and \U$10682 ( \10814 , \1484 , \4878 );
nor \U$10683 ( \10815 , \10813 , \10814 );
xnor \U$10684 ( \10816 , \10815 , \4762 );
xor \U$10685 ( \10817 , \10812 , \10816 );
and \U$10686 ( \10818 , \1147 , \5485 );
and \U$10687 ( \10819 , \1192 , \5275 );
nor \U$10688 ( \10820 , \10818 , \10819 );
xnor \U$10689 ( \10821 , \10820 , \5169 );
xor \U$10690 ( \10822 , \10817 , \10821 );
and \U$10691 ( \10823 , \189 , \7489 );
and \U$10692 ( \10824 , \197 , \7137 );
nor \U$10693 ( \10825 , \10823 , \10824 );
xnor \U$10694 ( \10826 , \10825 , \7142 );
and \U$10695 ( \10827 , \209 , \8019 );
and \U$10696 ( \10828 , \217 , \7830 );
nor \U$10697 ( \10829 , \10827 , \10828 );
xnor \U$10698 ( \10830 , \10829 , \7713 );
xor \U$10699 ( \10831 , \10826 , \10830 );
and \U$10700 ( \10832 , \224 , \8540 );
and \U$10701 ( \10833 , \232 , \8292 );
nor \U$10702 ( \10834 , \10832 , \10833 );
xnor \U$10703 ( \10835 , \10834 , \8297 );
xor \U$10704 ( \10836 , \10831 , \10835 );
xor \U$10705 ( \10837 , \10822 , \10836 );
and \U$10706 ( \10838 , \412 , \5996 );
and \U$10707 ( \10839 , \474 , \5695 );
nor \U$10708 ( \10840 , \10838 , \10839 );
xnor \U$10709 ( \10841 , \10840 , \5687 );
and \U$10710 ( \10842 , \261 , \6401 );
and \U$10711 ( \10843 , \307 , \6143 );
nor \U$10712 ( \10844 , \10842 , \10843 );
xnor \U$10713 ( \10845 , \10844 , \6148 );
xor \U$10714 ( \10846 , \10841 , \10845 );
and \U$10715 ( \10847 , \178 , \7055 );
and \U$10716 ( \10848 , \185 , \6675 );
nor \U$10717 ( \10849 , \10847 , \10848 );
xnor \U$10718 ( \10850 , \10849 , \6680 );
xor \U$10719 ( \10851 , \10846 , \10850 );
xor \U$10720 ( \10852 , \10837 , \10851 );
xor \U$10721 ( \10853 , \10808 , \10852 );
and \U$10722 ( \10854 , \4654 , \1578 );
and \U$10723 ( \10855 , \4749 , \1431 );
nor \U$10724 ( \10856 , \10854 , \10855 );
xnor \U$10725 ( \10857 , \10856 , \1436 );
and \U$10726 ( \10858 , \4160 , \1824 );
and \U$10727 ( \10859 , \4364 , \1739 );
nor \U$10728 ( \10860 , \10858 , \10859 );
xnor \U$10729 ( \10861 , \10860 , \1697 );
xor \U$10730 ( \10862 , \10857 , \10861 );
and \U$10731 ( \10863 , \3736 , \2121 );
and \U$10732 ( \10864 , \3912 , \2008 );
nor \U$10733 ( \10865 , \10863 , \10864 );
xnor \U$10734 ( \10866 , \10865 , \1961 );
xor \U$10735 ( \10867 , \10862 , \10866 );
and \U$10736 ( \10868 , \3395 , \2400 );
and \U$10737 ( \10869 , \3646 , \2246 );
nor \U$10738 ( \10870 , \10868 , \10869 );
xnor \U$10739 ( \10871 , \10870 , \2195 );
and \U$10740 ( \10872 , \3037 , \2669 );
and \U$10741 ( \10873 , \3143 , \2538 );
nor \U$10742 ( \10874 , \10872 , \10873 );
xnor \U$10743 ( \10875 , \10874 , \2534 );
xor \U$10744 ( \10876 , \10871 , \10875 );
and \U$10745 ( \10877 , \2757 , \3103 );
and \U$10746 ( \10878 , \2826 , \2934 );
nor \U$10747 ( \10879 , \10877 , \10878 );
xnor \U$10748 ( \10880 , \10879 , \2839 );
xor \U$10749 ( \10881 , \10876 , \10880 );
xor \U$10750 ( \10882 , \10867 , \10881 );
and \U$10751 ( \10883 , \2366 , \3357 );
and \U$10752 ( \10884 , \2521 , \3255 );
nor \U$10753 ( \10885 , \10883 , \10884 );
xnor \U$10754 ( \10886 , \10885 , \3156 );
and \U$10755 ( \10887 , \2090 , \3813 );
and \U$10756 ( \10888 , \2182 , \3557 );
nor \U$10757 ( \10889 , \10887 , \10888 );
xnor \U$10758 ( \10890 , \10889 , \3562 );
xor \U$10759 ( \10891 , \10886 , \10890 );
and \U$10760 ( \10892 , \1802 , \4132 );
and \U$10761 ( \10893 , \1948 , \4012 );
nor \U$10762 ( \10894 , \10892 , \10893 );
xnor \U$10763 ( \10895 , \10894 , \3925 );
xor \U$10764 ( \10896 , \10891 , \10895 );
xor \U$10765 ( \10897 , \10882 , \10896 );
xor \U$10766 ( \10898 , \10853 , \10897 );
xor \U$10767 ( \10899 , \10764 , \10898 );
and \U$10768 ( \10900 , \10537 , \10551 );
and \U$10769 ( \10901 , \10551 , \10566 );
and \U$10770 ( \10902 , \10537 , \10566 );
or \U$10771 ( \10903 , \10900 , \10901 , \10902 );
and \U$10772 ( \10904 , \10582 , \10597 );
xor \U$10773 ( \10905 , \10903 , \10904 );
and \U$10774 ( \10906 , \10584 , \183 );
not \U$10775 ( \10907 , \10906 );
xnor \U$10776 ( \10908 , \10907 , \179 );
and \U$10777 ( \10909 , \9897 , \195 );
and \U$10778 ( \10910 , \10206 , \193 );
nor \U$10779 ( \10911 , \10909 , \10910 );
xnor \U$10780 ( \10912 , \10911 , \202 );
xor \U$10781 ( \10913 , \10908 , \10912 );
xor \U$10782 ( \10914 , \10905 , \10913 );
xor \U$10783 ( \10915 , \10899 , \10914 );
xor \U$10784 ( \10916 , \10712 , \10915 );
xor \U$10785 ( \10917 , \10683 , \10916 );
xor \U$10786 ( \10918 , \10654 , \10917 );
xor \U$10787 ( \10919 , \10615 , \10918 );
and \U$10788 ( \10920 , \10294 , \10318 );
and \U$10789 ( \10921 , \10318 , \10602 );
and \U$10790 ( \10922 , \10294 , \10602 );
or \U$10791 ( \10923 , \10920 , \10921 , \10922 );
xor \U$10792 ( \10924 , \10919 , \10923 );
and \U$10793 ( \10925 , \10603 , \10604 );
and \U$10794 ( \10926 , \10605 , \10608 );
or \U$10795 ( \10927 , \10925 , \10926 );
xor \U$10796 ( \10928 , \10924 , \10927 );
buf \U$10797 ( \10929 , \10928 );
buf \U$10798 ( \10930 , \10929 );
and \U$10799 ( \10931 , \10619 , \10653 );
and \U$10800 ( \10932 , \10653 , \10917 );
and \U$10801 ( \10933 , \10619 , \10917 );
or \U$10802 ( \10934 , \10931 , \10932 , \10933 );
and \U$10803 ( \10935 , \10623 , \10627 );
and \U$10804 ( \10936 , \10627 , \10652 );
and \U$10805 ( \10937 , \10623 , \10652 );
or \U$10806 ( \10938 , \10935 , \10936 , \10937 );
and \U$10807 ( \10939 , \10668 , \10682 );
and \U$10808 ( \10940 , \10682 , \10916 );
and \U$10809 ( \10941 , \10668 , \10916 );
or \U$10810 ( \10942 , \10939 , \10940 , \10941 );
xor \U$10811 ( \10943 , \10938 , \10942 );
and \U$10812 ( \10944 , \10716 , \10720 );
and \U$10813 ( \10945 , \10720 , \10725 );
and \U$10814 ( \10946 , \10716 , \10725 );
or \U$10815 ( \10947 , \10944 , \10945 , \10946 );
and \U$10816 ( \10948 , \10641 , \10645 );
and \U$10817 ( \10949 , \10645 , \10650 );
and \U$10818 ( \10950 , \10641 , \10650 );
or \U$10819 ( \10951 , \10948 , \10949 , \10950 );
xor \U$10820 ( \10952 , \10947 , \10951 );
and \U$10821 ( \10953 , \10730 , \10734 );
and \U$10822 ( \10954 , \10734 , \10739 );
and \U$10823 ( \10955 , \10730 , \10739 );
or \U$10824 ( \10956 , \10953 , \10954 , \10955 );
xor \U$10825 ( \10957 , \10952 , \10956 );
and \U$10826 ( \10958 , \10726 , \10740 );
and \U$10827 ( \10959 , \10740 , \10763 );
and \U$10828 ( \10960 , \10726 , \10763 );
or \U$10829 ( \10961 , \10958 , \10959 , \10960 );
and \U$10830 ( \10962 , \10808 , \10852 );
and \U$10831 ( \10963 , \10852 , \10897 );
and \U$10832 ( \10964 , \10808 , \10897 );
or \U$10833 ( \10965 , \10962 , \10963 , \10964 );
xor \U$10834 ( \10966 , \10961 , \10965 );
and \U$10835 ( \10967 , \10812 , \10816 );
and \U$10836 ( \10968 , \10816 , \10821 );
and \U$10837 ( \10969 , \10812 , \10821 );
or \U$10838 ( \10970 , \10967 , \10968 , \10969 );
and \U$10839 ( \10971 , \10841 , \10845 );
and \U$10840 ( \10972 , \10845 , \10850 );
and \U$10841 ( \10973 , \10841 , \10850 );
or \U$10842 ( \10974 , \10971 , \10972 , \10973 );
xor \U$10843 ( \10975 , \10970 , \10974 );
and \U$10844 ( \10976 , \10886 , \10890 );
and \U$10845 ( \10977 , \10890 , \10895 );
and \U$10846 ( \10978 , \10886 , \10895 );
or \U$10847 ( \10979 , \10976 , \10977 , \10978 );
xor \U$10848 ( \10980 , \10975 , \10979 );
and \U$10849 ( \10981 , \10857 , \10861 );
and \U$10850 ( \10982 , \10861 , \10866 );
and \U$10851 ( \10983 , \10857 , \10866 );
or \U$10852 ( \10984 , \10981 , \10982 , \10983 );
and \U$10853 ( \10985 , \10871 , \10875 );
and \U$10854 ( \10986 , \10875 , \10880 );
and \U$10855 ( \10987 , \10871 , \10880 );
or \U$10856 ( \10988 , \10985 , \10986 , \10987 );
xor \U$10857 ( \10989 , \10984 , \10988 );
and \U$10858 ( \10990 , \10797 , \10801 );
and \U$10859 ( \10991 , \10801 , \10806 );
and \U$10860 ( \10992 , \10797 , \10806 );
or \U$10861 ( \10993 , \10990 , \10991 , \10992 );
xor \U$10862 ( \10994 , \10989 , \10993 );
xor \U$10863 ( \10995 , \10980 , \10994 );
and \U$10864 ( \10996 , \10768 , \10772 );
and \U$10865 ( \10997 , \10772 , \10777 );
and \U$10866 ( \10998 , \10768 , \10777 );
or \U$10867 ( \10999 , \10996 , \10997 , \10998 );
and \U$10868 ( \11000 , \10782 , \10786 );
and \U$10869 ( \11001 , \10786 , \10791 );
and \U$10870 ( \11002 , \10782 , \10791 );
or \U$10871 ( \11003 , \11000 , \11001 , \11002 );
xor \U$10872 ( \11004 , \10999 , \11003 );
and \U$10873 ( \11005 , \10908 , \10912 );
xor \U$10874 ( \11006 , \11004 , \11005 );
xor \U$10875 ( \11007 , \10995 , \11006 );
xor \U$10876 ( \11008 , \10966 , \11007 );
xor \U$10877 ( \11009 , \10957 , \11008 );
and \U$10878 ( \11010 , \10822 , \10836 );
and \U$10879 ( \11011 , \10836 , \10851 );
and \U$10880 ( \11012 , \10822 , \10851 );
or \U$10881 ( \11013 , \11010 , \11011 , \11012 );
and \U$10882 ( \11014 , \10867 , \10881 );
and \U$10883 ( \11015 , \10881 , \10896 );
and \U$10884 ( \11016 , \10867 , \10896 );
or \U$10885 ( \11017 , \11014 , \11015 , \11016 );
xor \U$10886 ( \11018 , \11013 , \11017 );
and \U$10887 ( \11019 , \10745 , \10747 );
and \U$10888 ( \11020 , \10747 , \10762 );
and \U$10889 ( \11021 , \10745 , \10762 );
or \U$10890 ( \11022 , \11019 , \11020 , \11021 );
xor \U$10891 ( \11023 , \11018 , \11022 );
and \U$10892 ( \11024 , \1484 , \5011 );
and \U$10893 ( \11025 , \1601 , \4878 );
nor \U$10894 ( \11026 , \11024 , \11025 );
xnor \U$10895 ( \11027 , \11026 , \4762 );
and \U$10896 ( \11028 , \1192 , \5485 );
and \U$10897 ( \11029 , \1333 , \5275 );
nor \U$10898 ( \11030 , \11028 , \11029 );
xnor \U$10899 ( \11031 , \11030 , \5169 );
xor \U$10900 ( \11032 , \11027 , \11031 );
and \U$10901 ( \11033 , \474 , \5996 );
and \U$10902 ( \11034 , \1147 , \5695 );
nor \U$10903 ( \11035 , \11033 , \11034 );
xnor \U$10904 ( \11036 , \11035 , \5687 );
xor \U$10905 ( \11037 , \11032 , \11036 );
and \U$10906 ( \11038 , \2182 , \3813 );
and \U$10907 ( \11039 , \2366 , \3557 );
nor \U$10908 ( \11040 , \11038 , \11039 );
xnor \U$10909 ( \11041 , \11040 , \3562 );
and \U$10910 ( \11042 , \1948 , \4132 );
and \U$10911 ( \11043 , \2090 , \4012 );
nor \U$10912 ( \11044 , \11042 , \11043 );
xnor \U$10913 ( \11045 , \11044 , \3925 );
xor \U$10914 ( \11046 , \11041 , \11045 );
and \U$10915 ( \11047 , \1684 , \4581 );
and \U$10916 ( \11048 , \1802 , \4424 );
nor \U$10917 ( \11049 , \11047 , \11048 );
xnor \U$10918 ( \11050 , \11049 , \4377 );
xor \U$10919 ( \11051 , \11046 , \11050 );
xor \U$10920 ( \11052 , \11037 , \11051 );
and \U$10921 ( \11053 , \3143 , \2669 );
and \U$10922 ( \11054 , \3395 , \2538 );
nor \U$10923 ( \11055 , \11053 , \11054 );
xnor \U$10924 ( \11056 , \11055 , \2534 );
and \U$10925 ( \11057 , \2826 , \3103 );
and \U$10926 ( \11058 , \3037 , \2934 );
nor \U$10927 ( \11059 , \11057 , \11058 );
xnor \U$10928 ( \11060 , \11059 , \2839 );
xor \U$10929 ( \11061 , \11056 , \11060 );
and \U$10930 ( \11062 , \2521 , \3357 );
and \U$10931 ( \11063 , \2757 , \3255 );
nor \U$10932 ( \11064 , \11062 , \11063 );
xnor \U$10933 ( \11065 , \11064 , \3156 );
xor \U$10934 ( \11066 , \11061 , \11065 );
xor \U$10935 ( \11067 , \11052 , \11066 );
and \U$10936 ( \11068 , \217 , \8019 );
and \U$10937 ( \11069 , \189 , \7830 );
nor \U$10938 ( \11070 , \11068 , \11069 );
xnor \U$10939 ( \11071 , \11070 , \7713 );
and \U$10940 ( \11072 , \232 , \8540 );
and \U$10941 ( \11073 , \209 , \8292 );
nor \U$10942 ( \11074 , \11072 , \11073 );
xnor \U$10943 ( \11075 , \11074 , \8297 );
xor \U$10944 ( \11076 , \11071 , \11075 );
and \U$10945 ( \11077 , \247 , \9333 );
and \U$10946 ( \11078 , \224 , \9006 );
nor \U$10947 ( \11079 , \11077 , \11078 );
xnor \U$10948 ( \11080 , \11079 , \8848 );
xor \U$10949 ( \11081 , \11076 , \11080 );
and \U$10950 ( \11082 , \143 , \9765 );
and \U$10951 ( \11083 , \240 , \9644 );
nor \U$10952 ( \11084 , \11082 , \11083 );
xnor \U$10953 ( \11085 , \11084 , \9478 );
and \U$10954 ( \11086 , \158 , \10408 );
and \U$10955 ( \11087 , \134 , \10116 );
nor \U$10956 ( \11088 , \11086 , \11087 );
xnor \U$10957 ( \11089 , \11088 , \10121 );
xor \U$10958 ( \11090 , \11085 , \11089 );
and \U$10959 ( \11091 , \150 , \10118 );
xor \U$10960 ( \11092 , \11090 , \11091 );
xor \U$10961 ( \11093 , \11081 , \11092 );
and \U$10962 ( \11094 , \307 , \6401 );
and \U$10963 ( \11095 , \412 , \6143 );
nor \U$10964 ( \11096 , \11094 , \11095 );
xnor \U$10965 ( \11097 , \11096 , \6148 );
and \U$10966 ( \11098 , \185 , \7055 );
and \U$10967 ( \11099 , \261 , \6675 );
nor \U$10968 ( \11100 , \11098 , \11099 );
xnor \U$10969 ( \11101 , \11100 , \6680 );
xor \U$10970 ( \11102 , \11097 , \11101 );
and \U$10971 ( \11103 , \197 , \7489 );
and \U$10972 ( \11104 , \178 , \7137 );
nor \U$10973 ( \11105 , \11103 , \11104 );
xnor \U$10974 ( \11106 , \11105 , \7142 );
xor \U$10975 ( \11107 , \11102 , \11106 );
xor \U$10976 ( \11108 , \11093 , \11107 );
xor \U$10977 ( \11109 , \11067 , \11108 );
and \U$10978 ( \11110 , \10826 , \10830 );
and \U$10979 ( \11111 , \10830 , \10835 );
and \U$10980 ( \11112 , \10826 , \10835 );
or \U$10981 ( \11113 , \11110 , \11111 , \11112 );
and \U$10982 ( \11114 , \10752 , \10756 );
and \U$10983 ( \11115 , \10756 , \10761 );
and \U$10984 ( \11116 , \10752 , \10761 );
or \U$10985 ( \11117 , \11114 , \11115 , \11116 );
xnor \U$10986 ( \11118 , \11113 , \11117 );
xor \U$10987 ( \11119 , \11109 , \11118 );
xor \U$10988 ( \11120 , \11023 , \11119 );
and \U$10989 ( \11121 , \10778 , \10792 );
and \U$10990 ( \11122 , \10792 , \10807 );
and \U$10991 ( \11123 , \10778 , \10807 );
or \U$10992 ( \11124 , \11121 , \11122 , \11123 );
and \U$10993 ( \11125 , \4364 , \1824 );
and \U$10994 ( \11126 , \4654 , \1739 );
nor \U$10995 ( \11127 , \11125 , \11126 );
xnor \U$10996 ( \11128 , \11127 , \1697 );
and \U$10997 ( \11129 , \3912 , \2121 );
and \U$10998 ( \11130 , \4160 , \2008 );
nor \U$10999 ( \11131 , \11129 , \11130 );
xnor \U$11000 ( \11132 , \11131 , \1961 );
xor \U$11001 ( \11133 , \11128 , \11132 );
and \U$11002 ( \11134 , \3646 , \2400 );
and \U$11003 ( \11135 , \3736 , \2246 );
nor \U$11004 ( \11136 , \11134 , \11135 );
xnor \U$11005 ( \11137 , \11136 , \2195 );
xor \U$11006 ( \11138 , \11133 , \11137 );
and \U$11007 ( \11139 , \7231 , \156 );
and \U$11008 ( \11140 , \7556 , \154 );
nor \U$11009 ( \11141 , \11139 , \11140 );
xnor \U$11010 ( \11142 , \11141 , \163 );
and \U$11011 ( \11143 , \6790 , \296 );
and \U$11012 ( \11144 , \6945 , \168 );
nor \U$11013 ( \11145 , \11143 , \11144 );
xnor \U$11014 ( \11146 , \11145 , \173 );
xor \U$11015 ( \11147 , \11142 , \11146 );
and \U$11016 ( \11148 , \6281 , \438 );
and \U$11017 ( \11149 , \6514 , \336 );
nor \U$11018 ( \11150 , \11148 , \11149 );
xnor \U$11019 ( \11151 , \11150 , \320 );
xor \U$11020 ( \11152 , \11147 , \11151 );
xor \U$11021 ( \11153 , \11138 , \11152 );
and \U$11022 ( \11154 , \5674 , \1086 );
and \U$11023 ( \11155 , \6030 , \508 );
nor \U$11024 ( \11156 , \11154 , \11155 );
xnor \U$11025 ( \11157 , \11156 , \487 );
and \U$11026 ( \11158 , \5156 , \1301 );
and \U$11027 ( \11159 , \5469 , \1246 );
nor \U$11028 ( \11160 , \11158 , \11159 );
xnor \U$11029 ( \11161 , \11160 , \1205 );
xor \U$11030 ( \11162 , \11157 , \11161 );
and \U$11031 ( \11163 , \4749 , \1578 );
and \U$11032 ( \11164 , \4922 , \1431 );
nor \U$11033 ( \11165 , \11163 , \11164 );
xnor \U$11034 ( \11166 , \11165 , \1436 );
xor \U$11035 ( \11167 , \11162 , \11166 );
xor \U$11036 ( \11168 , \11153 , \11167 );
xor \U$11037 ( \11169 , \11124 , \11168 );
not \U$11038 ( \11170 , \179 );
and \U$11039 ( \11171 , \10206 , \195 );
and \U$11040 ( \11172 , \10584 , \193 );
nor \U$11041 ( \11173 , \11171 , \11172 );
xnor \U$11042 ( \11174 , \11173 , \202 );
xor \U$11043 ( \11175 , \11170 , \11174 );
and \U$11044 ( \11176 , \9465 , \215 );
and \U$11045 ( \11177 , \9897 , \213 );
nor \U$11046 ( \11178 , \11176 , \11177 );
xnor \U$11047 ( \11179 , \11178 , \222 );
xor \U$11048 ( \11180 , \11175 , \11179 );
and \U$11049 ( \11181 , \8835 , \230 );
and \U$11050 ( \11182 , \9169 , \228 );
nor \U$11051 ( \11183 , \11181 , \11182 );
xnor \U$11052 ( \11184 , \11183 , \237 );
and \U$11053 ( \11185 , \8349 , \245 );
and \U$11054 ( \11186 , \8652 , \243 );
nor \U$11055 ( \11187 , \11185 , \11186 );
xnor \U$11056 ( \11188 , \11187 , \252 );
xor \U$11057 ( \11189 , \11184 , \11188 );
and \U$11058 ( \11190 , \7700 , \141 );
and \U$11059 ( \11191 , \8057 , \139 );
nor \U$11060 ( \11192 , \11190 , \11191 );
xnor \U$11061 ( \11193 , \11192 , \148 );
xor \U$11062 ( \11194 , \11189 , \11193 );
xor \U$11063 ( \11195 , \11180 , \11194 );
xor \U$11064 ( \11196 , \11169 , \11195 );
xor \U$11065 ( \11197 , \11120 , \11196 );
xor \U$11066 ( \11198 , \11009 , \11197 );
xor \U$11067 ( \11199 , \10943 , \11198 );
xor \U$11068 ( \11200 , \10934 , \11199 );
and \U$11069 ( \11201 , \10658 , \10662 );
and \U$11070 ( \11202 , \10662 , \10667 );
and \U$11071 ( \11203 , \10658 , \10667 );
or \U$11072 ( \11204 , \11201 , \11202 , \11203 );
and \U$11073 ( \11205 , \10632 , \10636 );
and \U$11074 ( \11206 , \10636 , \10651 );
and \U$11075 ( \11207 , \10632 , \10651 );
or \U$11076 ( \11208 , \11205 , \11206 , \11207 );
xor \U$11077 ( \11209 , \11204 , \11208 );
and \U$11078 ( \11210 , \10764 , \10898 );
and \U$11079 ( \11211 , \10898 , \10914 );
and \U$11080 ( \11212 , \10764 , \10914 );
or \U$11081 ( \11213 , \11210 , \11211 , \11212 );
xor \U$11082 ( \11214 , \11209 , \11213 );
and \U$11083 ( \11215 , \10672 , \10676 );
and \U$11084 ( \11216 , \10676 , \10681 );
and \U$11085 ( \11217 , \10672 , \10681 );
or \U$11086 ( \11218 , \11215 , \11216 , \11217 );
and \U$11087 ( \11219 , \10697 , \10711 );
and \U$11088 ( \11220 , \10711 , \10915 );
and \U$11089 ( \11221 , \10697 , \10915 );
or \U$11090 ( \11222 , \11219 , \11220 , \11221 );
xor \U$11091 ( \11223 , \11218 , \11222 );
and \U$11092 ( \11224 , \10687 , \10691 );
and \U$11093 ( \11225 , \10691 , \10696 );
and \U$11094 ( \11226 , \10687 , \10696 );
or \U$11095 ( \11227 , \11224 , \11225 , \11226 );
and \U$11096 ( \11228 , \10701 , \10705 );
and \U$11097 ( \11229 , \10705 , \10710 );
and \U$11098 ( \11230 , \10701 , \10710 );
or \U$11099 ( \11231 , \11228 , \11229 , \11230 );
xor \U$11100 ( \11232 , \11227 , \11231 );
and \U$11101 ( \11233 , \10903 , \10904 );
and \U$11102 ( \11234 , \10904 , \10913 );
and \U$11103 ( \11235 , \10903 , \10913 );
or \U$11104 ( \11236 , \11233 , \11234 , \11235 );
xor \U$11105 ( \11237 , \11232 , \11236 );
xor \U$11106 ( \11238 , \11223 , \11237 );
xor \U$11107 ( \11239 , \11214 , \11238 );
xor \U$11108 ( \11240 , \11200 , \11239 );
and \U$11109 ( \11241 , \10615 , \10918 );
xor \U$11110 ( \11242 , \11240 , \11241 );
and \U$11111 ( \11243 , \10919 , \10923 );
and \U$11112 ( \11244 , \10924 , \10927 );
or \U$11113 ( \11245 , \11243 , \11244 );
xor \U$11114 ( \11246 , \11242 , \11245 );
buf \U$11115 ( \11247 , \11246 );
buf \U$11116 ( \11248 , \11247 );
and \U$11117 ( \11249 , \10938 , \10942 );
and \U$11118 ( \11250 , \10942 , \11198 );
and \U$11119 ( \11251 , \10938 , \11198 );
or \U$11120 ( \11252 , \11249 , \11250 , \11251 );
and \U$11121 ( \11253 , \11214 , \11238 );
xor \U$11122 ( \11254 , \11252 , \11253 );
and \U$11123 ( \11255 , \11218 , \11222 );
and \U$11124 ( \11256 , \11222 , \11237 );
and \U$11125 ( \11257 , \11218 , \11237 );
or \U$11126 ( \11258 , \11255 , \11256 , \11257 );
and \U$11127 ( \11259 , \11204 , \11208 );
and \U$11128 ( \11260 , \11208 , \11213 );
and \U$11129 ( \11261 , \11204 , \11213 );
or \U$11130 ( \11262 , \11259 , \11260 , \11261 );
and \U$11131 ( \11263 , \10957 , \11008 );
and \U$11132 ( \11264 , \11008 , \11197 );
and \U$11133 ( \11265 , \10957 , \11197 );
or \U$11134 ( \11266 , \11263 , \11264 , \11265 );
xor \U$11135 ( \11267 , \11262 , \11266 );
and \U$11136 ( \11268 , \10980 , \10994 );
and \U$11137 ( \11269 , \10994 , \11006 );
and \U$11138 ( \11270 , \10980 , \11006 );
or \U$11139 ( \11271 , \11268 , \11269 , \11270 );
and \U$11140 ( \11272 , \11067 , \11108 );
and \U$11141 ( \11273 , \11108 , \11118 );
and \U$11142 ( \11274 , \11067 , \11118 );
or \U$11143 ( \11275 , \11272 , \11273 , \11274 );
xor \U$11144 ( \11276 , \11271 , \11275 );
and \U$11145 ( \11277 , \11170 , \11174 );
and \U$11146 ( \11278 , \11174 , \11179 );
and \U$11147 ( \11279 , \11170 , \11179 );
or \U$11148 ( \11280 , \11277 , \11278 , \11279 );
and \U$11149 ( \11281 , \11184 , \11188 );
and \U$11150 ( \11282 , \11188 , \11193 );
and \U$11151 ( \11283 , \11184 , \11193 );
or \U$11152 ( \11284 , \11281 , \11282 , \11283 );
xor \U$11153 ( \11285 , \11280 , \11284 );
and \U$11154 ( \11286 , \11142 , \11146 );
and \U$11155 ( \11287 , \11146 , \11151 );
and \U$11156 ( \11288 , \11142 , \11151 );
or \U$11157 ( \11289 , \11286 , \11287 , \11288 );
xor \U$11158 ( \11290 , \11285 , \11289 );
xor \U$11159 ( \11291 , \11276 , \11290 );
xor \U$11160 ( \11292 , \11267 , \11291 );
xor \U$11161 ( \11293 , \11258 , \11292 );
and \U$11162 ( \11294 , \11013 , \11017 );
and \U$11163 ( \11295 , \11017 , \11022 );
and \U$11164 ( \11296 , \11013 , \11022 );
or \U$11165 ( \11297 , \11294 , \11295 , \11296 );
and \U$11166 ( \11298 , \10947 , \10951 );
and \U$11167 ( \11299 , \10951 , \10956 );
and \U$11168 ( \11300 , \10947 , \10956 );
or \U$11169 ( \11301 , \11298 , \11299 , \11300 );
xor \U$11170 ( \11302 , \11297 , \11301 );
and \U$11171 ( \11303 , \11124 , \11168 );
and \U$11172 ( \11304 , \11168 , \11195 );
and \U$11173 ( \11305 , \11124 , \11195 );
or \U$11174 ( \11306 , \11303 , \11304 , \11305 );
xor \U$11175 ( \11307 , \11302 , \11306 );
and \U$11176 ( \11308 , \11227 , \11231 );
and \U$11177 ( \11309 , \11231 , \11236 );
and \U$11178 ( \11310 , \11227 , \11236 );
or \U$11179 ( \11311 , \11308 , \11309 , \11310 );
and \U$11180 ( \11312 , \10961 , \10965 );
and \U$11181 ( \11313 , \10965 , \11007 );
and \U$11182 ( \11314 , \10961 , \11007 );
or \U$11183 ( \11315 , \11312 , \11313 , \11314 );
xor \U$11184 ( \11316 , \11311 , \11315 );
and \U$11185 ( \11317 , \11023 , \11119 );
and \U$11186 ( \11318 , \11119 , \11196 );
and \U$11187 ( \11319 , \11023 , \11196 );
or \U$11188 ( \11320 , \11317 , \11318 , \11319 );
xor \U$11189 ( \11321 , \11316 , \11320 );
xor \U$11190 ( \11322 , \11307 , \11321 );
and \U$11191 ( \11323 , \11037 , \11051 );
and \U$11192 ( \11324 , \11051 , \11066 );
and \U$11193 ( \11325 , \11037 , \11066 );
or \U$11194 ( \11326 , \11323 , \11324 , \11325 );
and \U$11195 ( \11327 , \11081 , \11092 );
and \U$11196 ( \11328 , \11092 , \11107 );
and \U$11197 ( \11329 , \11081 , \11107 );
or \U$11198 ( \11330 , \11327 , \11328 , \11329 );
xor \U$11199 ( \11331 , \11326 , \11330 );
or \U$11200 ( \11332 , \11113 , \11117 );
xor \U$11201 ( \11333 , \11331 , \11332 );
and \U$11202 ( \11334 , \10970 , \10974 );
and \U$11203 ( \11335 , \10974 , \10979 );
and \U$11204 ( \11336 , \10970 , \10979 );
or \U$11205 ( \11337 , \11334 , \11335 , \11336 );
and \U$11206 ( \11338 , \10984 , \10988 );
and \U$11207 ( \11339 , \10988 , \10993 );
and \U$11208 ( \11340 , \10984 , \10993 );
or \U$11209 ( \11341 , \11338 , \11339 , \11340 );
xor \U$11210 ( \11342 , \11337 , \11341 );
and \U$11211 ( \11343 , \10999 , \11003 );
and \U$11212 ( \11344 , \11003 , \11005 );
and \U$11213 ( \11345 , \10999 , \11005 );
or \U$11214 ( \11346 , \11343 , \11344 , \11345 );
xor \U$11215 ( \11347 , \11342 , \11346 );
xor \U$11216 ( \11348 , \11333 , \11347 );
and \U$11217 ( \11349 , \11138 , \11152 );
and \U$11218 ( \11350 , \11152 , \11167 );
and \U$11219 ( \11351 , \11138 , \11167 );
or \U$11220 ( \11352 , \11349 , \11350 , \11351 );
and \U$11221 ( \11353 , \11180 , \11194 );
xor \U$11222 ( \11354 , \11352 , \11353 );
and \U$11223 ( \11355 , \10584 , \195 );
not \U$11224 ( \11356 , \11355 );
xnor \U$11225 ( \11357 , \11356 , \202 );
and \U$11226 ( \11358 , \9897 , \215 );
and \U$11227 ( \11359 , \10206 , \213 );
nor \U$11228 ( \11360 , \11358 , \11359 );
xnor \U$11229 ( \11361 , \11360 , \222 );
xor \U$11230 ( \11362 , \11357 , \11361 );
and \U$11231 ( \11363 , \9169 , \230 );
and \U$11232 ( \11364 , \9465 , \228 );
nor \U$11233 ( \11365 , \11363 , \11364 );
xnor \U$11234 ( \11366 , \11365 , \237 );
xor \U$11235 ( \11367 , \11362 , \11366 );
xor \U$11236 ( \11368 , \11354 , \11367 );
and \U$11237 ( \11369 , \5469 , \1301 );
and \U$11238 ( \11370 , \5674 , \1246 );
nor \U$11239 ( \11371 , \11369 , \11370 );
xnor \U$11240 ( \11372 , \11371 , \1205 );
and \U$11241 ( \11373 , \4922 , \1578 );
and \U$11242 ( \11374 , \5156 , \1431 );
nor \U$11243 ( \11375 , \11373 , \11374 );
xnor \U$11244 ( \11376 , \11375 , \1436 );
xor \U$11245 ( \11377 , \11372 , \11376 );
and \U$11246 ( \11378 , \4654 , \1824 );
and \U$11247 ( \11379 , \4749 , \1739 );
nor \U$11248 ( \11380 , \11378 , \11379 );
xnor \U$11249 ( \11381 , \11380 , \1697 );
xor \U$11250 ( \11382 , \11377 , \11381 );
and \U$11251 ( \11383 , \6945 , \296 );
and \U$11252 ( \11384 , \7231 , \168 );
nor \U$11253 ( \11385 , \11383 , \11384 );
xnor \U$11254 ( \11386 , \11385 , \173 );
and \U$11255 ( \11387 , \6514 , \438 );
and \U$11256 ( \11388 , \6790 , \336 );
nor \U$11257 ( \11389 , \11387 , \11388 );
xnor \U$11258 ( \11390 , \11389 , \320 );
xor \U$11259 ( \11391 , \11386 , \11390 );
and \U$11260 ( \11392 , \6030 , \1086 );
and \U$11261 ( \11393 , \6281 , \508 );
nor \U$11262 ( \11394 , \11392 , \11393 );
xnor \U$11263 ( \11395 , \11394 , \487 );
xor \U$11264 ( \11396 , \11391 , \11395 );
xor \U$11265 ( \11397 , \11382 , \11396 );
and \U$11266 ( \11398 , \8652 , \245 );
and \U$11267 ( \11399 , \8835 , \243 );
nor \U$11268 ( \11400 , \11398 , \11399 );
xnor \U$11269 ( \11401 , \11400 , \252 );
and \U$11270 ( \11402 , \8057 , \141 );
and \U$11271 ( \11403 , \8349 , \139 );
nor \U$11272 ( \11404 , \11402 , \11403 );
xnor \U$11273 ( \11405 , \11404 , \148 );
xor \U$11274 ( \11406 , \11401 , \11405 );
and \U$11275 ( \11407 , \7556 , \156 );
and \U$11276 ( \11408 , \7700 , \154 );
nor \U$11277 ( \11409 , \11407 , \11408 );
xnor \U$11278 ( \11410 , \11409 , \163 );
xor \U$11279 ( \11411 , \11406 , \11410 );
xor \U$11280 ( \11412 , \11397 , \11411 );
and \U$11281 ( \11413 , \3037 , \3103 );
and \U$11282 ( \11414 , \3143 , \2934 );
nor \U$11283 ( \11415 , \11413 , \11414 );
xnor \U$11284 ( \11416 , \11415 , \2839 );
and \U$11285 ( \11417 , \2757 , \3357 );
and \U$11286 ( \11418 , \2826 , \3255 );
nor \U$11287 ( \11419 , \11417 , \11418 );
xnor \U$11288 ( \11420 , \11419 , \3156 );
xor \U$11289 ( \11421 , \11416 , \11420 );
and \U$11290 ( \11422 , \2366 , \3813 );
and \U$11291 ( \11423 , \2521 , \3557 );
nor \U$11292 ( \11424 , \11422 , \11423 );
xnor \U$11293 ( \11425 , \11424 , \3562 );
xor \U$11294 ( \11426 , \11421 , \11425 );
and \U$11295 ( \11427 , \4160 , \2121 );
and \U$11296 ( \11428 , \4364 , \2008 );
nor \U$11297 ( \11429 , \11427 , \11428 );
xnor \U$11298 ( \11430 , \11429 , \1961 );
and \U$11299 ( \11431 , \3736 , \2400 );
and \U$11300 ( \11432 , \3912 , \2246 );
nor \U$11301 ( \11433 , \11431 , \11432 );
xnor \U$11302 ( \11434 , \11433 , \2195 );
xor \U$11303 ( \11435 , \11430 , \11434 );
and \U$11304 ( \11436 , \3395 , \2669 );
and \U$11305 ( \11437 , \3646 , \2538 );
nor \U$11306 ( \11438 , \11436 , \11437 );
xnor \U$11307 ( \11439 , \11438 , \2534 );
xor \U$11308 ( \11440 , \11435 , \11439 );
xor \U$11309 ( \11441 , \11426 , \11440 );
and \U$11310 ( \11442 , \2090 , \4132 );
and \U$11311 ( \11443 , \2182 , \4012 );
nor \U$11312 ( \11444 , \11442 , \11443 );
xnor \U$11313 ( \11445 , \11444 , \3925 );
and \U$11314 ( \11446 , \1802 , \4581 );
and \U$11315 ( \11447 , \1948 , \4424 );
nor \U$11316 ( \11448 , \11446 , \11447 );
xnor \U$11317 ( \11449 , \11448 , \4377 );
xor \U$11318 ( \11450 , \11445 , \11449 );
and \U$11319 ( \11451 , \1601 , \5011 );
and \U$11320 ( \11452 , \1684 , \4878 );
nor \U$11321 ( \11453 , \11451 , \11452 );
xnor \U$11322 ( \11454 , \11453 , \4762 );
xor \U$11323 ( \11455 , \11450 , \11454 );
xor \U$11324 ( \11456 , \11441 , \11455 );
xor \U$11325 ( \11457 , \11412 , \11456 );
and \U$11326 ( \11458 , \261 , \7055 );
and \U$11327 ( \11459 , \307 , \6675 );
nor \U$11328 ( \11460 , \11458 , \11459 );
xnor \U$11329 ( \11461 , \11460 , \6680 );
and \U$11330 ( \11462 , \178 , \7489 );
and \U$11331 ( \11463 , \185 , \7137 );
nor \U$11332 ( \11464 , \11462 , \11463 );
xnor \U$11333 ( \11465 , \11464 , \7142 );
xor \U$11334 ( \11466 , \11461 , \11465 );
and \U$11335 ( \11467 , \189 , \8019 );
and \U$11336 ( \11468 , \197 , \7830 );
nor \U$11337 ( \11469 , \11467 , \11468 );
xnor \U$11338 ( \11470 , \11469 , \7713 );
xor \U$11339 ( \11471 , \11466 , \11470 );
and \U$11340 ( \11472 , \209 , \8540 );
and \U$11341 ( \11473 , \217 , \8292 );
nor \U$11342 ( \11474 , \11472 , \11473 );
xnor \U$11343 ( \11475 , \11474 , \8297 );
and \U$11344 ( \11476 , \224 , \9333 );
and \U$11345 ( \11477 , \232 , \9006 );
nor \U$11346 ( \11478 , \11476 , \11477 );
xnor \U$11347 ( \11479 , \11478 , \8848 );
xor \U$11348 ( \11480 , \11475 , \11479 );
and \U$11349 ( \11481 , \240 , \9765 );
and \U$11350 ( \11482 , \247 , \9644 );
nor \U$11351 ( \11483 , \11481 , \11482 );
xnor \U$11352 ( \11484 , \11483 , \9478 );
xor \U$11353 ( \11485 , \11480 , \11484 );
xor \U$11354 ( \11486 , \11471 , \11485 );
and \U$11355 ( \11487 , \1333 , \5485 );
and \U$11356 ( \11488 , \1484 , \5275 );
nor \U$11357 ( \11489 , \11487 , \11488 );
xnor \U$11358 ( \11490 , \11489 , \5169 );
and \U$11359 ( \11491 , \1147 , \5996 );
and \U$11360 ( \11492 , \1192 , \5695 );
nor \U$11361 ( \11493 , \11491 , \11492 );
xnor \U$11362 ( \11494 , \11493 , \5687 );
xor \U$11363 ( \11495 , \11490 , \11494 );
and \U$11364 ( \11496 , \412 , \6401 );
and \U$11365 ( \11497 , \474 , \6143 );
nor \U$11366 ( \11498 , \11496 , \11497 );
xnor \U$11367 ( \11499 , \11498 , \6148 );
xor \U$11368 ( \11500 , \11495 , \11499 );
xor \U$11369 ( \11501 , \11486 , \11500 );
xor \U$11370 ( \11502 , \11457 , \11501 );
xor \U$11371 ( \11503 , \11368 , \11502 );
and \U$11372 ( \11504 , \11027 , \11031 );
and \U$11373 ( \11505 , \11031 , \11036 );
and \U$11374 ( \11506 , \11027 , \11036 );
or \U$11375 ( \11507 , \11504 , \11505 , \11506 );
and \U$11376 ( \11508 , \11041 , \11045 );
and \U$11377 ( \11509 , \11045 , \11050 );
and \U$11378 ( \11510 , \11041 , \11050 );
or \U$11379 ( \11511 , \11508 , \11509 , \11510 );
xor \U$11380 ( \11512 , \11507 , \11511 );
and \U$11381 ( \11513 , \11097 , \11101 );
and \U$11382 ( \11514 , \11101 , \11106 );
and \U$11383 ( \11515 , \11097 , \11106 );
or \U$11384 ( \11516 , \11513 , \11514 , \11515 );
xor \U$11385 ( \11517 , \11512 , \11516 );
and \U$11386 ( \11518 , \11128 , \11132 );
and \U$11387 ( \11519 , \11132 , \11137 );
and \U$11388 ( \11520 , \11128 , \11137 );
or \U$11389 ( \11521 , \11518 , \11519 , \11520 );
and \U$11390 ( \11522 , \11056 , \11060 );
and \U$11391 ( \11523 , \11060 , \11065 );
and \U$11392 ( \11524 , \11056 , \11065 );
or \U$11393 ( \11525 , \11522 , \11523 , \11524 );
xor \U$11394 ( \11526 , \11521 , \11525 );
and \U$11395 ( \11527 , \11157 , \11161 );
and \U$11396 ( \11528 , \11161 , \11166 );
and \U$11397 ( \11529 , \11157 , \11166 );
or \U$11398 ( \11530 , \11527 , \11528 , \11529 );
xor \U$11399 ( \11531 , \11526 , \11530 );
xor \U$11400 ( \11532 , \11517 , \11531 );
and \U$11401 ( \11533 , \11071 , \11075 );
and \U$11402 ( \11534 , \11075 , \11080 );
and \U$11403 ( \11535 , \11071 , \11080 );
or \U$11404 ( \11536 , \11533 , \11534 , \11535 );
and \U$11405 ( \11537 , \11085 , \11089 );
and \U$11406 ( \11538 , \11089 , \11091 );
and \U$11407 ( \11539 , \11085 , \11091 );
or \U$11408 ( \11540 , \11537 , \11538 , \11539 );
xor \U$11409 ( \11541 , \11536 , \11540 );
and \U$11410 ( \11542 , \134 , \10408 );
and \U$11411 ( \11543 , \143 , \10116 );
nor \U$11412 ( \11544 , \11542 , \11543 );
xnor \U$11413 ( \11545 , \11544 , \10121 );
and \U$11414 ( \11546 , \158 , \10118 );
xnor \U$11415 ( \11547 , \11545 , \11546 );
xor \U$11416 ( \11548 , \11541 , \11547 );
xor \U$11417 ( \11549 , \11532 , \11548 );
xor \U$11418 ( \11550 , \11503 , \11549 );
xor \U$11419 ( \11551 , \11348 , \11550 );
xor \U$11420 ( \11552 , \11322 , \11551 );
xor \U$11421 ( \11553 , \11293 , \11552 );
xor \U$11422 ( \11554 , \11254 , \11553 );
and \U$11423 ( \11555 , \10934 , \11199 );
and \U$11424 ( \11556 , \11199 , \11239 );
and \U$11425 ( \11557 , \10934 , \11239 );
or \U$11426 ( \11558 , \11555 , \11556 , \11557 );
xor \U$11427 ( \11559 , \11554 , \11558 );
and \U$11428 ( \11560 , \11240 , \11241 );
and \U$11429 ( \11561 , \11242 , \11245 );
or \U$11430 ( \11562 , \11560 , \11561 );
xor \U$11431 ( \11563 , \11559 , \11562 );
buf \U$11432 ( \11564 , \11563 );
buf \U$11433 ( \11565 , \11564 );
and \U$11434 ( \11566 , \11258 , \11292 );
and \U$11435 ( \11567 , \11292 , \11552 );
and \U$11436 ( \11568 , \11258 , \11552 );
or \U$11437 ( \11569 , \11566 , \11567 , \11568 );
and \U$11438 ( \11570 , \11262 , \11266 );
and \U$11439 ( \11571 , \11266 , \11291 );
and \U$11440 ( \11572 , \11262 , \11291 );
or \U$11441 ( \11573 , \11570 , \11571 , \11572 );
and \U$11442 ( \11574 , \11307 , \11321 );
and \U$11443 ( \11575 , \11321 , \11551 );
and \U$11444 ( \11576 , \11307 , \11551 );
or \U$11445 ( \11577 , \11574 , \11575 , \11576 );
xor \U$11446 ( \11578 , \11573 , \11577 );
and \U$11447 ( \11579 , \11280 , \11284 );
and \U$11448 ( \11580 , \11284 , \11289 );
and \U$11449 ( \11581 , \11280 , \11289 );
or \U$11450 ( \11582 , \11579 , \11580 , \11581 );
and \U$11451 ( \11583 , \11507 , \11511 );
and \U$11452 ( \11584 , \11511 , \11516 );
and \U$11453 ( \11585 , \11507 , \11516 );
or \U$11454 ( \11586 , \11583 , \11584 , \11585 );
xor \U$11455 ( \11587 , \11582 , \11586 );
and \U$11456 ( \11588 , \11521 , \11525 );
and \U$11457 ( \11589 , \11525 , \11530 );
and \U$11458 ( \11590 , \11521 , \11530 );
or \U$11459 ( \11591 , \11588 , \11589 , \11590 );
xor \U$11460 ( \11592 , \11587 , \11591 );
and \U$11461 ( \11593 , \11412 , \11456 );
and \U$11462 ( \11594 , \11456 , \11501 );
and \U$11463 ( \11595 , \11412 , \11501 );
or \U$11464 ( \11596 , \11593 , \11594 , \11595 );
and \U$11465 ( \11597 , \11517 , \11531 );
and \U$11466 ( \11598 , \11531 , \11548 );
and \U$11467 ( \11599 , \11517 , \11548 );
or \U$11468 ( \11600 , \11597 , \11598 , \11599 );
xor \U$11469 ( \11601 , \11596 , \11600 );
and \U$11470 ( \11602 , \11386 , \11390 );
and \U$11471 ( \11603 , \11390 , \11395 );
and \U$11472 ( \11604 , \11386 , \11395 );
or \U$11473 ( \11605 , \11602 , \11603 , \11604 );
and \U$11474 ( \11606 , \11357 , \11361 );
and \U$11475 ( \11607 , \11361 , \11366 );
and \U$11476 ( \11608 , \11357 , \11366 );
or \U$11477 ( \11609 , \11606 , \11607 , \11608 );
xor \U$11478 ( \11610 , \11605 , \11609 );
and \U$11479 ( \11611 , \11401 , \11405 );
and \U$11480 ( \11612 , \11405 , \11410 );
and \U$11481 ( \11613 , \11401 , \11410 );
or \U$11482 ( \11614 , \11611 , \11612 , \11613 );
xor \U$11483 ( \11615 , \11610 , \11614 );
and \U$11484 ( \11616 , \11461 , \11465 );
and \U$11485 ( \11617 , \11465 , \11470 );
and \U$11486 ( \11618 , \11461 , \11470 );
or \U$11487 ( \11619 , \11616 , \11617 , \11618 );
and \U$11488 ( \11620 , \11445 , \11449 );
and \U$11489 ( \11621 , \11449 , \11454 );
and \U$11490 ( \11622 , \11445 , \11454 );
or \U$11491 ( \11623 , \11620 , \11621 , \11622 );
xor \U$11492 ( \11624 , \11619 , \11623 );
and \U$11493 ( \11625 , \11490 , \11494 );
and \U$11494 ( \11626 , \11494 , \11499 );
and \U$11495 ( \11627 , \11490 , \11499 );
or \U$11496 ( \11628 , \11625 , \11626 , \11627 );
xor \U$11497 ( \11629 , \11624 , \11628 );
xor \U$11498 ( \11630 , \11615 , \11629 );
and \U$11499 ( \11631 , \11372 , \11376 );
and \U$11500 ( \11632 , \11376 , \11381 );
and \U$11501 ( \11633 , \11372 , \11381 );
or \U$11502 ( \11634 , \11631 , \11632 , \11633 );
and \U$11503 ( \11635 , \11416 , \11420 );
and \U$11504 ( \11636 , \11420 , \11425 );
and \U$11505 ( \11637 , \11416 , \11425 );
or \U$11506 ( \11638 , \11635 , \11636 , \11637 );
xor \U$11507 ( \11639 , \11634 , \11638 );
and \U$11508 ( \11640 , \11430 , \11434 );
and \U$11509 ( \11641 , \11434 , \11439 );
and \U$11510 ( \11642 , \11430 , \11439 );
or \U$11511 ( \11643 , \11640 , \11641 , \11642 );
xor \U$11512 ( \11644 , \11639 , \11643 );
xor \U$11513 ( \11645 , \11630 , \11644 );
xor \U$11514 ( \11646 , \11601 , \11645 );
xor \U$11515 ( \11647 , \11592 , \11646 );
and \U$11516 ( \11648 , \11426 , \11440 );
and \U$11517 ( \11649 , \11440 , \11455 );
and \U$11518 ( \11650 , \11426 , \11455 );
or \U$11519 ( \11651 , \11648 , \11649 , \11650 );
and \U$11520 ( \11652 , \11471 , \11485 );
and \U$11521 ( \11653 , \11485 , \11500 );
and \U$11522 ( \11654 , \11471 , \11500 );
or \U$11523 ( \11655 , \11652 , \11653 , \11654 );
xor \U$11524 ( \11656 , \11651 , \11655 );
and \U$11525 ( \11657 , \11536 , \11540 );
and \U$11526 ( \11658 , \11540 , \11547 );
and \U$11527 ( \11659 , \11536 , \11547 );
or \U$11528 ( \11660 , \11657 , \11658 , \11659 );
xor \U$11529 ( \11661 , \11656 , \11660 );
and \U$11530 ( \11662 , \11475 , \11479 );
and \U$11531 ( \11663 , \11479 , \11484 );
and \U$11532 ( \11664 , \11475 , \11484 );
or \U$11533 ( \11665 , \11662 , \11663 , \11664 );
or \U$11534 ( \11666 , \11545 , \11546 );
xor \U$11535 ( \11667 , \11665 , \11666 );
and \U$11536 ( \11668 , \143 , \10408 );
and \U$11537 ( \11669 , \240 , \10116 );
nor \U$11538 ( \11670 , \11668 , \11669 );
xnor \U$11539 ( \11671 , \11670 , \10121 );
xor \U$11540 ( \11672 , \11667 , \11671 );
and \U$11541 ( \11673 , \134 , \10118 );
and \U$11542 ( \11674 , \307 , \7055 );
and \U$11543 ( \11675 , \412 , \6675 );
nor \U$11544 ( \11676 , \11674 , \11675 );
xnor \U$11545 ( \11677 , \11676 , \6680 );
and \U$11546 ( \11678 , \185 , \7489 );
and \U$11547 ( \11679 , \261 , \7137 );
nor \U$11548 ( \11680 , \11678 , \11679 );
xnor \U$11549 ( \11681 , \11680 , \7142 );
xor \U$11550 ( \11682 , \11677 , \11681 );
and \U$11551 ( \11683 , \197 , \8019 );
and \U$11552 ( \11684 , \178 , \7830 );
nor \U$11553 ( \11685 , \11683 , \11684 );
xnor \U$11554 ( \11686 , \11685 , \7713 );
xor \U$11555 ( \11687 , \11682 , \11686 );
xor \U$11556 ( \11688 , \11673 , \11687 );
and \U$11557 ( \11689 , \217 , \8540 );
and \U$11558 ( \11690 , \189 , \8292 );
nor \U$11559 ( \11691 , \11689 , \11690 );
xnor \U$11560 ( \11692 , \11691 , \8297 );
and \U$11561 ( \11693 , \232 , \9333 );
and \U$11562 ( \11694 , \209 , \9006 );
nor \U$11563 ( \11695 , \11693 , \11694 );
xnor \U$11564 ( \11696 , \11695 , \8848 );
xor \U$11565 ( \11697 , \11692 , \11696 );
and \U$11566 ( \11698 , \247 , \9765 );
and \U$11567 ( \11699 , \224 , \9644 );
nor \U$11568 ( \11700 , \11698 , \11699 );
xnor \U$11569 ( \11701 , \11700 , \9478 );
xor \U$11570 ( \11702 , \11697 , \11701 );
xor \U$11571 ( \11703 , \11688 , \11702 );
xor \U$11572 ( \11704 , \11672 , \11703 );
and \U$11573 ( \11705 , \3143 , \3103 );
and \U$11574 ( \11706 , \3395 , \2934 );
nor \U$11575 ( \11707 , \11705 , \11706 );
xnor \U$11576 ( \11708 , \11707 , \2839 );
and \U$11577 ( \11709 , \2826 , \3357 );
and \U$11578 ( \11710 , \3037 , \3255 );
nor \U$11579 ( \11711 , \11709 , \11710 );
xnor \U$11580 ( \11712 , \11711 , \3156 );
xor \U$11581 ( \11713 , \11708 , \11712 );
and \U$11582 ( \11714 , \2521 , \3813 );
and \U$11583 ( \11715 , \2757 , \3557 );
nor \U$11584 ( \11716 , \11714 , \11715 );
xnor \U$11585 ( \11717 , \11716 , \3562 );
xor \U$11586 ( \11718 , \11713 , \11717 );
and \U$11587 ( \11719 , \1484 , \5485 );
and \U$11588 ( \11720 , \1601 , \5275 );
nor \U$11589 ( \11721 , \11719 , \11720 );
xnor \U$11590 ( \11722 , \11721 , \5169 );
and \U$11591 ( \11723 , \1192 , \5996 );
and \U$11592 ( \11724 , \1333 , \5695 );
nor \U$11593 ( \11725 , \11723 , \11724 );
xnor \U$11594 ( \11726 , \11725 , \5687 );
xor \U$11595 ( \11727 , \11722 , \11726 );
and \U$11596 ( \11728 , \474 , \6401 );
and \U$11597 ( \11729 , \1147 , \6143 );
nor \U$11598 ( \11730 , \11728 , \11729 );
xnor \U$11599 ( \11731 , \11730 , \6148 );
xor \U$11600 ( \11732 , \11727 , \11731 );
xor \U$11601 ( \11733 , \11718 , \11732 );
and \U$11602 ( \11734 , \2182 , \4132 );
and \U$11603 ( \11735 , \2366 , \4012 );
nor \U$11604 ( \11736 , \11734 , \11735 );
xnor \U$11605 ( \11737 , \11736 , \3925 );
and \U$11606 ( \11738 , \1948 , \4581 );
and \U$11607 ( \11739 , \2090 , \4424 );
nor \U$11608 ( \11740 , \11738 , \11739 );
xnor \U$11609 ( \11741 , \11740 , \4377 );
xor \U$11610 ( \11742 , \11737 , \11741 );
and \U$11611 ( \11743 , \1684 , \5011 );
and \U$11612 ( \11744 , \1802 , \4878 );
nor \U$11613 ( \11745 , \11743 , \11744 );
xnor \U$11614 ( \11746 , \11745 , \4762 );
xor \U$11615 ( \11747 , \11742 , \11746 );
xor \U$11616 ( \11748 , \11733 , \11747 );
xor \U$11617 ( \11749 , \11704 , \11748 );
xor \U$11618 ( \11750 , \11661 , \11749 );
and \U$11619 ( \11751 , \11382 , \11396 );
and \U$11620 ( \11752 , \11396 , \11411 );
and \U$11621 ( \11753 , \11382 , \11411 );
or \U$11622 ( \11754 , \11751 , \11752 , \11753 );
and \U$11623 ( \11755 , \7231 , \296 );
and \U$11624 ( \11756 , \7556 , \168 );
nor \U$11625 ( \11757 , \11755 , \11756 );
xnor \U$11626 ( \11758 , \11757 , \173 );
and \U$11627 ( \11759 , \6790 , \438 );
and \U$11628 ( \11760 , \6945 , \336 );
nor \U$11629 ( \11761 , \11759 , \11760 );
xnor \U$11630 ( \11762 , \11761 , \320 );
xor \U$11631 ( \11763 , \11758 , \11762 );
and \U$11632 ( \11764 , \6281 , \1086 );
and \U$11633 ( \11765 , \6514 , \508 );
nor \U$11634 ( \11766 , \11764 , \11765 );
xnor \U$11635 ( \11767 , \11766 , \487 );
xor \U$11636 ( \11768 , \11763 , \11767 );
and \U$11637 ( \11769 , \4364 , \2121 );
and \U$11638 ( \11770 , \4654 , \2008 );
nor \U$11639 ( \11771 , \11769 , \11770 );
xnor \U$11640 ( \11772 , \11771 , \1961 );
and \U$11641 ( \11773 , \3912 , \2400 );
and \U$11642 ( \11774 , \4160 , \2246 );
nor \U$11643 ( \11775 , \11773 , \11774 );
xnor \U$11644 ( \11776 , \11775 , \2195 );
xor \U$11645 ( \11777 , \11772 , \11776 );
and \U$11646 ( \11778 , \3646 , \2669 );
and \U$11647 ( \11779 , \3736 , \2538 );
nor \U$11648 ( \11780 , \11778 , \11779 );
xnor \U$11649 ( \11781 , \11780 , \2534 );
xor \U$11650 ( \11782 , \11777 , \11781 );
xor \U$11651 ( \11783 , \11768 , \11782 );
and \U$11652 ( \11784 , \5674 , \1301 );
and \U$11653 ( \11785 , \6030 , \1246 );
nor \U$11654 ( \11786 , \11784 , \11785 );
xnor \U$11655 ( \11787 , \11786 , \1205 );
and \U$11656 ( \11788 , \5156 , \1578 );
and \U$11657 ( \11789 , \5469 , \1431 );
nor \U$11658 ( \11790 , \11788 , \11789 );
xnor \U$11659 ( \11791 , \11790 , \1436 );
xor \U$11660 ( \11792 , \11787 , \11791 );
and \U$11661 ( \11793 , \4749 , \1824 );
and \U$11662 ( \11794 , \4922 , \1739 );
nor \U$11663 ( \11795 , \11793 , \11794 );
xnor \U$11664 ( \11796 , \11795 , \1697 );
xor \U$11665 ( \11797 , \11792 , \11796 );
xor \U$11666 ( \11798 , \11783 , \11797 );
xor \U$11667 ( \11799 , \11754 , \11798 );
and \U$11668 ( \11800 , \8835 , \245 );
and \U$11669 ( \11801 , \9169 , \243 );
nor \U$11670 ( \11802 , \11800 , \11801 );
xnor \U$11671 ( \11803 , \11802 , \252 );
and \U$11672 ( \11804 , \8349 , \141 );
and \U$11673 ( \11805 , \8652 , \139 );
nor \U$11674 ( \11806 , \11804 , \11805 );
xnor \U$11675 ( \11807 , \11806 , \148 );
xor \U$11676 ( \11808 , \11803 , \11807 );
and \U$11677 ( \11809 , \7700 , \156 );
and \U$11678 ( \11810 , \8057 , \154 );
nor \U$11679 ( \11811 , \11809 , \11810 );
xnor \U$11680 ( \11812 , \11811 , \163 );
xor \U$11681 ( \11813 , \11808 , \11812 );
not \U$11682 ( \11814 , \202 );
and \U$11683 ( \11815 , \10206 , \215 );
and \U$11684 ( \11816 , \10584 , \213 );
nor \U$11685 ( \11817 , \11815 , \11816 );
xnor \U$11686 ( \11818 , \11817 , \222 );
xor \U$11687 ( \11819 , \11814 , \11818 );
and \U$11688 ( \11820 , \9465 , \230 );
and \U$11689 ( \11821 , \9897 , \228 );
nor \U$11690 ( \11822 , \11820 , \11821 );
xnor \U$11691 ( \11823 , \11822 , \237 );
xor \U$11692 ( \11824 , \11819 , \11823 );
xor \U$11693 ( \11825 , \11813 , \11824 );
xor \U$11694 ( \11826 , \11799 , \11825 );
xor \U$11695 ( \11827 , \11750 , \11826 );
xor \U$11696 ( \11828 , \11647 , \11827 );
xor \U$11697 ( \11829 , \11578 , \11828 );
xor \U$11698 ( \11830 , \11569 , \11829 );
and \U$11699 ( \11831 , \11297 , \11301 );
and \U$11700 ( \11832 , \11301 , \11306 );
and \U$11701 ( \11833 , \11297 , \11306 );
or \U$11702 ( \11834 , \11831 , \11832 , \11833 );
and \U$11703 ( \11835 , \11271 , \11275 );
and \U$11704 ( \11836 , \11275 , \11290 );
and \U$11705 ( \11837 , \11271 , \11290 );
or \U$11706 ( \11838 , \11835 , \11836 , \11837 );
xor \U$11707 ( \11839 , \11834 , \11838 );
and \U$11708 ( \11840 , \11368 , \11502 );
and \U$11709 ( \11841 , \11502 , \11549 );
and \U$11710 ( \11842 , \11368 , \11549 );
or \U$11711 ( \11843 , \11840 , \11841 , \11842 );
xor \U$11712 ( \11844 , \11839 , \11843 );
and \U$11713 ( \11845 , \11311 , \11315 );
and \U$11714 ( \11846 , \11315 , \11320 );
and \U$11715 ( \11847 , \11311 , \11320 );
or \U$11716 ( \11848 , \11845 , \11846 , \11847 );
and \U$11717 ( \11849 , \11333 , \11347 );
and \U$11718 ( \11850 , \11347 , \11550 );
and \U$11719 ( \11851 , \11333 , \11550 );
or \U$11720 ( \11852 , \11849 , \11850 , \11851 );
xor \U$11721 ( \11853 , \11848 , \11852 );
and \U$11722 ( \11854 , \11326 , \11330 );
and \U$11723 ( \11855 , \11330 , \11332 );
and \U$11724 ( \11856 , \11326 , \11332 );
or \U$11725 ( \11857 , \11854 , \11855 , \11856 );
and \U$11726 ( \11858 , \11337 , \11341 );
and \U$11727 ( \11859 , \11341 , \11346 );
and \U$11728 ( \11860 , \11337 , \11346 );
or \U$11729 ( \11861 , \11858 , \11859 , \11860 );
xor \U$11730 ( \11862 , \11857 , \11861 );
and \U$11731 ( \11863 , \11352 , \11353 );
and \U$11732 ( \11864 , \11353 , \11367 );
and \U$11733 ( \11865 , \11352 , \11367 );
or \U$11734 ( \11866 , \11863 , \11864 , \11865 );
xor \U$11735 ( \11867 , \11862 , \11866 );
xor \U$11736 ( \11868 , \11853 , \11867 );
xor \U$11737 ( \11869 , \11844 , \11868 );
xor \U$11738 ( \11870 , \11830 , \11869 );
and \U$11739 ( \11871 , \11252 , \11253 );
and \U$11740 ( \11872 , \11253 , \11553 );
and \U$11741 ( \11873 , \11252 , \11553 );
or \U$11742 ( \11874 , \11871 , \11872 , \11873 );
xor \U$11743 ( \11875 , \11870 , \11874 );
and \U$11744 ( \11876 , \11554 , \11558 );
and \U$11745 ( \11877 , \11559 , \11562 );
or \U$11746 ( \11878 , \11876 , \11877 );
xor \U$11747 ( \11879 , \11875 , \11878 );
buf \U$11748 ( \11880 , \11879 );
buf \U$11749 ( \11881 , \11880 );
and \U$11750 ( \11882 , \11573 , \11577 );
and \U$11751 ( \11883 , \11577 , \11828 );
and \U$11752 ( \11884 , \11573 , \11828 );
or \U$11753 ( \11885 , \11882 , \11883 , \11884 );
and \U$11754 ( \11886 , \11844 , \11868 );
xor \U$11755 ( \11887 , \11885 , \11886 );
and \U$11756 ( \11888 , \11848 , \11852 );
and \U$11757 ( \11889 , \11852 , \11867 );
and \U$11758 ( \11890 , \11848 , \11867 );
or \U$11759 ( \11891 , \11888 , \11889 , \11890 );
and \U$11760 ( \11892 , \11834 , \11838 );
and \U$11761 ( \11893 , \11838 , \11843 );
and \U$11762 ( \11894 , \11834 , \11843 );
or \U$11763 ( \11895 , \11892 , \11893 , \11894 );
and \U$11764 ( \11896 , \11592 , \11646 );
and \U$11765 ( \11897 , \11646 , \11827 );
and \U$11766 ( \11898 , \11592 , \11827 );
or \U$11767 ( \11899 , \11896 , \11897 , \11898 );
xor \U$11768 ( \11900 , \11895 , \11899 );
and \U$11769 ( \11901 , \11651 , \11655 );
and \U$11770 ( \11902 , \11655 , \11660 );
and \U$11771 ( \11903 , \11651 , \11660 );
or \U$11772 ( \11904 , \11901 , \11902 , \11903 );
and \U$11773 ( \11905 , \11582 , \11586 );
and \U$11774 ( \11906 , \11586 , \11591 );
and \U$11775 ( \11907 , \11582 , \11591 );
or \U$11776 ( \11908 , \11905 , \11906 , \11907 );
xor \U$11777 ( \11909 , \11904 , \11908 );
and \U$11778 ( \11910 , \11754 , \11798 );
and \U$11779 ( \11911 , \11798 , \11825 );
and \U$11780 ( \11912 , \11754 , \11825 );
or \U$11781 ( \11913 , \11910 , \11911 , \11912 );
xor \U$11782 ( \11914 , \11909 , \11913 );
xor \U$11783 ( \11915 , \11900 , \11914 );
xor \U$11784 ( \11916 , \11891 , \11915 );
and \U$11785 ( \11917 , \11857 , \11861 );
and \U$11786 ( \11918 , \11861 , \11866 );
and \U$11787 ( \11919 , \11857 , \11866 );
or \U$11788 ( \11920 , \11917 , \11918 , \11919 );
and \U$11789 ( \11921 , \11596 , \11600 );
and \U$11790 ( \11922 , \11600 , \11645 );
and \U$11791 ( \11923 , \11596 , \11645 );
or \U$11792 ( \11924 , \11921 , \11922 , \11923 );
xor \U$11793 ( \11925 , \11920 , \11924 );
and \U$11794 ( \11926 , \11661 , \11749 );
and \U$11795 ( \11927 , \11749 , \11826 );
and \U$11796 ( \11928 , \11661 , \11826 );
or \U$11797 ( \11929 , \11926 , \11927 , \11928 );
xor \U$11798 ( \11930 , \11925 , \11929 );
and \U$11799 ( \11931 , \11605 , \11609 );
and \U$11800 ( \11932 , \11609 , \11614 );
and \U$11801 ( \11933 , \11605 , \11614 );
or \U$11802 ( \11934 , \11931 , \11932 , \11933 );
and \U$11803 ( \11935 , \11619 , \11623 );
and \U$11804 ( \11936 , \11623 , \11628 );
and \U$11805 ( \11937 , \11619 , \11628 );
or \U$11806 ( \11938 , \11935 , \11936 , \11937 );
xor \U$11807 ( \11939 , \11934 , \11938 );
and \U$11808 ( \11940 , \11634 , \11638 );
and \U$11809 ( \11941 , \11638 , \11643 );
and \U$11810 ( \11942 , \11634 , \11643 );
or \U$11811 ( \11943 , \11940 , \11941 , \11942 );
xor \U$11812 ( \11944 , \11939 , \11943 );
and \U$11813 ( \11945 , \11615 , \11629 );
and \U$11814 ( \11946 , \11629 , \11644 );
and \U$11815 ( \11947 , \11615 , \11644 );
or \U$11816 ( \11948 , \11945 , \11946 , \11947 );
and \U$11817 ( \11949 , \11672 , \11703 );
and \U$11818 ( \11950 , \11703 , \11748 );
and \U$11819 ( \11951 , \11672 , \11748 );
or \U$11820 ( \11952 , \11949 , \11950 , \11951 );
xor \U$11821 ( \11953 , \11948 , \11952 );
and \U$11822 ( \11954 , \11708 , \11712 );
and \U$11823 ( \11955 , \11712 , \11717 );
and \U$11824 ( \11956 , \11708 , \11717 );
or \U$11825 ( \11957 , \11954 , \11955 , \11956 );
and \U$11826 ( \11958 , \11772 , \11776 );
and \U$11827 ( \11959 , \11776 , \11781 );
and \U$11828 ( \11960 , \11772 , \11781 );
or \U$11829 ( \11961 , \11958 , \11959 , \11960 );
xor \U$11830 ( \11962 , \11957 , \11961 );
and \U$11831 ( \11963 , \11787 , \11791 );
and \U$11832 ( \11964 , \11791 , \11796 );
and \U$11833 ( \11965 , \11787 , \11796 );
or \U$11834 ( \11966 , \11963 , \11964 , \11965 );
xor \U$11835 ( \11967 , \11962 , \11966 );
and \U$11836 ( \11968 , \11758 , \11762 );
and \U$11837 ( \11969 , \11762 , \11767 );
and \U$11838 ( \11970 , \11758 , \11767 );
or \U$11839 ( \11971 , \11968 , \11969 , \11970 );
and \U$11840 ( \11972 , \11803 , \11807 );
and \U$11841 ( \11973 , \11807 , \11812 );
and \U$11842 ( \11974 , \11803 , \11812 );
or \U$11843 ( \11975 , \11972 , \11973 , \11974 );
xor \U$11844 ( \11976 , \11971 , \11975 );
and \U$11845 ( \11977 , \11814 , \11818 );
and \U$11846 ( \11978 , \11818 , \11823 );
and \U$11847 ( \11979 , \11814 , \11823 );
or \U$11848 ( \11980 , \11977 , \11978 , \11979 );
xor \U$11849 ( \11981 , \11976 , \11980 );
xor \U$11850 ( \11982 , \11967 , \11981 );
and \U$11851 ( \11983 , \11677 , \11681 );
and \U$11852 ( \11984 , \11681 , \11686 );
and \U$11853 ( \11985 , \11677 , \11686 );
or \U$11854 ( \11986 , \11983 , \11984 , \11985 );
and \U$11855 ( \11987 , \11722 , \11726 );
and \U$11856 ( \11988 , \11726 , \11731 );
and \U$11857 ( \11989 , \11722 , \11731 );
or \U$11858 ( \11990 , \11987 , \11988 , \11989 );
xor \U$11859 ( \11991 , \11986 , \11990 );
and \U$11860 ( \11992 , \11737 , \11741 );
and \U$11861 ( \11993 , \11741 , \11746 );
and \U$11862 ( \11994 , \11737 , \11746 );
or \U$11863 ( \11995 , \11992 , \11993 , \11994 );
xor \U$11864 ( \11996 , \11991 , \11995 );
xor \U$11865 ( \11997 , \11982 , \11996 );
xor \U$11866 ( \11998 , \11953 , \11997 );
xor \U$11867 ( \11999 , \11944 , \11998 );
and \U$11868 ( \12000 , \11665 , \11666 );
and \U$11869 ( \12001 , \11666 , \11671 );
and \U$11870 ( \12002 , \11665 , \11671 );
or \U$11871 ( \12003 , \12000 , \12001 , \12002 );
and \U$11872 ( \12004 , \11673 , \11687 );
and \U$11873 ( \12005 , \11687 , \11702 );
and \U$11874 ( \12006 , \11673 , \11702 );
or \U$11875 ( \12007 , \12004 , \12005 , \12006 );
xor \U$11876 ( \12008 , \12003 , \12007 );
and \U$11877 ( \12009 , \11718 , \11732 );
and \U$11878 ( \12010 , \11732 , \11747 );
and \U$11879 ( \12011 , \11718 , \11747 );
or \U$11880 ( \12012 , \12009 , \12010 , \12011 );
xor \U$11881 ( \12013 , \12008 , \12012 );
and \U$11882 ( \12014 , \11768 , \11782 );
and \U$11883 ( \12015 , \11782 , \11797 );
and \U$11884 ( \12016 , \11768 , \11797 );
or \U$11885 ( \12017 , \12014 , \12015 , \12016 );
and \U$11886 ( \12018 , \11813 , \11824 );
xor \U$11887 ( \12019 , \12017 , \12018 );
and \U$11888 ( \12020 , \10584 , \215 );
not \U$11889 ( \12021 , \12020 );
xnor \U$11890 ( \12022 , \12021 , \222 );
and \U$11891 ( \12023 , \9897 , \230 );
and \U$11892 ( \12024 , \10206 , \228 );
nor \U$11893 ( \12025 , \12023 , \12024 );
xnor \U$11894 ( \12026 , \12025 , \237 );
xor \U$11895 ( \12027 , \12022 , \12026 );
and \U$11896 ( \12028 , \9169 , \245 );
and \U$11897 ( \12029 , \9465 , \243 );
nor \U$11898 ( \12030 , \12028 , \12029 );
xnor \U$11899 ( \12031 , \12030 , \252 );
xor \U$11900 ( \12032 , \12027 , \12031 );
and \U$11901 ( \12033 , \6945 , \438 );
and \U$11902 ( \12034 , \7231 , \336 );
nor \U$11903 ( \12035 , \12033 , \12034 );
xnor \U$11904 ( \12036 , \12035 , \320 );
and \U$11905 ( \12037 , \6514 , \1086 );
and \U$11906 ( \12038 , \6790 , \508 );
nor \U$11907 ( \12039 , \12037 , \12038 );
xnor \U$11908 ( \12040 , \12039 , \487 );
xor \U$11909 ( \12041 , \12036 , \12040 );
and \U$11910 ( \12042 , \6030 , \1301 );
and \U$11911 ( \12043 , \6281 , \1246 );
nor \U$11912 ( \12044 , \12042 , \12043 );
xnor \U$11913 ( \12045 , \12044 , \1205 );
xor \U$11914 ( \12046 , \12041 , \12045 );
xor \U$11915 ( \12047 , \12032 , \12046 );
and \U$11916 ( \12048 , \8652 , \141 );
and \U$11917 ( \12049 , \8835 , \139 );
nor \U$11918 ( \12050 , \12048 , \12049 );
xnor \U$11919 ( \12051 , \12050 , \148 );
and \U$11920 ( \12052 , \8057 , \156 );
and \U$11921 ( \12053 , \8349 , \154 );
nor \U$11922 ( \12054 , \12052 , \12053 );
xnor \U$11923 ( \12055 , \12054 , \163 );
xor \U$11924 ( \12056 , \12051 , \12055 );
and \U$11925 ( \12057 , \7556 , \296 );
and \U$11926 ( \12058 , \7700 , \168 );
nor \U$11927 ( \12059 , \12057 , \12058 );
xnor \U$11928 ( \12060 , \12059 , \173 );
xor \U$11929 ( \12061 , \12056 , \12060 );
xor \U$11930 ( \12062 , \12047 , \12061 );
xor \U$11931 ( \12063 , \12019 , \12062 );
xor \U$11932 ( \12064 , \12013 , \12063 );
and \U$11933 ( \12065 , \5469 , \1578 );
and \U$11934 ( \12066 , \5674 , \1431 );
nor \U$11935 ( \12067 , \12065 , \12066 );
xnor \U$11936 ( \12068 , \12067 , \1436 );
and \U$11937 ( \12069 , \4922 , \1824 );
and \U$11938 ( \12070 , \5156 , \1739 );
nor \U$11939 ( \12071 , \12069 , \12070 );
xnor \U$11940 ( \12072 , \12071 , \1697 );
xor \U$11941 ( \12073 , \12068 , \12072 );
and \U$11942 ( \12074 , \4654 , \2121 );
and \U$11943 ( \12075 , \4749 , \2008 );
nor \U$11944 ( \12076 , \12074 , \12075 );
xnor \U$11945 ( \12077 , \12076 , \1961 );
xor \U$11946 ( \12078 , \12073 , \12077 );
and \U$11947 ( \12079 , \3037 , \3357 );
and \U$11948 ( \12080 , \3143 , \3255 );
nor \U$11949 ( \12081 , \12079 , \12080 );
xnor \U$11950 ( \12082 , \12081 , \3156 );
and \U$11951 ( \12083 , \2757 , \3813 );
and \U$11952 ( \12084 , \2826 , \3557 );
nor \U$11953 ( \12085 , \12083 , \12084 );
xnor \U$11954 ( \12086 , \12085 , \3562 );
xor \U$11955 ( \12087 , \12082 , \12086 );
and \U$11956 ( \12088 , \2366 , \4132 );
and \U$11957 ( \12089 , \2521 , \4012 );
nor \U$11958 ( \12090 , \12088 , \12089 );
xnor \U$11959 ( \12091 , \12090 , \3925 );
xor \U$11960 ( \12092 , \12087 , \12091 );
xor \U$11961 ( \12093 , \12078 , \12092 );
and \U$11962 ( \12094 , \4160 , \2400 );
and \U$11963 ( \12095 , \4364 , \2246 );
nor \U$11964 ( \12096 , \12094 , \12095 );
xnor \U$11965 ( \12097 , \12096 , \2195 );
and \U$11966 ( \12098 , \3736 , \2669 );
and \U$11967 ( \12099 , \3912 , \2538 );
nor \U$11968 ( \12100 , \12098 , \12099 );
xnor \U$11969 ( \12101 , \12100 , \2534 );
xor \U$11970 ( \12102 , \12097 , \12101 );
and \U$11971 ( \12103 , \3395 , \3103 );
and \U$11972 ( \12104 , \3646 , \2934 );
nor \U$11973 ( \12105 , \12103 , \12104 );
xnor \U$11974 ( \12106 , \12105 , \2839 );
xor \U$11975 ( \12107 , \12102 , \12106 );
xor \U$11976 ( \12108 , \12093 , \12107 );
and \U$11977 ( \12109 , \1333 , \5996 );
and \U$11978 ( \12110 , \1484 , \5695 );
nor \U$11979 ( \12111 , \12109 , \12110 );
xnor \U$11980 ( \12112 , \12111 , \5687 );
and \U$11981 ( \12113 , \1147 , \6401 );
and \U$11982 ( \12114 , \1192 , \6143 );
nor \U$11983 ( \12115 , \12113 , \12114 );
xnor \U$11984 ( \12116 , \12115 , \6148 );
xor \U$11985 ( \12117 , \12112 , \12116 );
and \U$11986 ( \12118 , \412 , \7055 );
and \U$11987 ( \12119 , \474 , \6675 );
nor \U$11988 ( \12120 , \12118 , \12119 );
xnor \U$11989 ( \12121 , \12120 , \6680 );
xor \U$11990 ( \12122 , \12117 , \12121 );
and \U$11991 ( \12123 , \2090 , \4581 );
and \U$11992 ( \12124 , \2182 , \4424 );
nor \U$11993 ( \12125 , \12123 , \12124 );
xnor \U$11994 ( \12126 , \12125 , \4377 );
and \U$11995 ( \12127 , \1802 , \5011 );
and \U$11996 ( \12128 , \1948 , \4878 );
nor \U$11997 ( \12129 , \12127 , \12128 );
xnor \U$11998 ( \12130 , \12129 , \4762 );
xor \U$11999 ( \12131 , \12126 , \12130 );
and \U$12000 ( \12132 , \1601 , \5485 );
and \U$12001 ( \12133 , \1684 , \5275 );
nor \U$12002 ( \12134 , \12132 , \12133 );
xnor \U$12003 ( \12135 , \12134 , \5169 );
xor \U$12004 ( \12136 , \12131 , \12135 );
xor \U$12005 ( \12137 , \12122 , \12136 );
and \U$12006 ( \12138 , \261 , \7489 );
and \U$12007 ( \12139 , \307 , \7137 );
nor \U$12008 ( \12140 , \12138 , \12139 );
xnor \U$12009 ( \12141 , \12140 , \7142 );
and \U$12010 ( \12142 , \178 , \8019 );
and \U$12011 ( \12143 , \185 , \7830 );
nor \U$12012 ( \12144 , \12142 , \12143 );
xnor \U$12013 ( \12145 , \12144 , \7713 );
xor \U$12014 ( \12146 , \12141 , \12145 );
and \U$12015 ( \12147 , \189 , \8540 );
and \U$12016 ( \12148 , \197 , \8292 );
nor \U$12017 ( \12149 , \12147 , \12148 );
xnor \U$12018 ( \12150 , \12149 , \8297 );
xor \U$12019 ( \12151 , \12146 , \12150 );
xor \U$12020 ( \12152 , \12137 , \12151 );
xor \U$12021 ( \12153 , \12108 , \12152 );
and \U$12022 ( \12154 , \11692 , \11696 );
and \U$12023 ( \12155 , \11696 , \11701 );
and \U$12024 ( \12156 , \11692 , \11701 );
or \U$12025 ( \12157 , \12154 , \12155 , \12156 );
and \U$12026 ( \12158 , \209 , \9333 );
and \U$12027 ( \12159 , \217 , \9006 );
nor \U$12028 ( \12160 , \12158 , \12159 );
xnor \U$12029 ( \12161 , \12160 , \8848 );
and \U$12030 ( \12162 , \224 , \9765 );
and \U$12031 ( \12163 , \232 , \9644 );
nor \U$12032 ( \12164 , \12162 , \12163 );
xnor \U$12033 ( \12165 , \12164 , \9478 );
xor \U$12034 ( \12166 , \12161 , \12165 );
and \U$12035 ( \12167 , \240 , \10408 );
and \U$12036 ( \12168 , \247 , \10116 );
nor \U$12037 ( \12169 , \12167 , \12168 );
xnor \U$12038 ( \12170 , \12169 , \10121 );
xor \U$12039 ( \12171 , \12166 , \12170 );
xor \U$12040 ( \12172 , \12157 , \12171 );
and \U$12041 ( \12173 , \143 , \10118 );
not \U$12042 ( \12174 , \12173 );
xor \U$12043 ( \12175 , \12172 , \12174 );
xor \U$12044 ( \12176 , \12153 , \12175 );
xor \U$12045 ( \12177 , \12064 , \12176 );
xor \U$12046 ( \12178 , \11999 , \12177 );
xor \U$12047 ( \12179 , \11930 , \12178 );
xor \U$12048 ( \12180 , \11916 , \12179 );
xor \U$12049 ( \12181 , \11887 , \12180 );
and \U$12050 ( \12182 , \11569 , \11829 );
and \U$12051 ( \12183 , \11829 , \11869 );
and \U$12052 ( \12184 , \11569 , \11869 );
or \U$12053 ( \12185 , \12182 , \12183 , \12184 );
xor \U$12054 ( \12186 , \12181 , \12185 );
and \U$12055 ( \12187 , \11870 , \11874 );
and \U$12056 ( \12188 , \11875 , \11878 );
or \U$12057 ( \12189 , \12187 , \12188 );
xor \U$12058 ( \12190 , \12186 , \12189 );
buf \U$12059 ( \12191 , \12190 );
buf \U$12060 ( \12192 , \12191 );
and \U$12061 ( \12193 , \11891 , \11915 );
and \U$12062 ( \12194 , \11915 , \12179 );
and \U$12063 ( \12195 , \11891 , \12179 );
or \U$12064 ( \12196 , \12193 , \12194 , \12195 );
and \U$12065 ( \12197 , \11895 , \11899 );
and \U$12066 ( \12198 , \11899 , \11914 );
and \U$12067 ( \12199 , \11895 , \11914 );
or \U$12068 ( \12200 , \12197 , \12198 , \12199 );
and \U$12069 ( \12201 , \11930 , \12178 );
xor \U$12070 ( \12202 , \12200 , \12201 );
and \U$12071 ( \12203 , \11957 , \11961 );
and \U$12072 ( \12204 , \11961 , \11966 );
and \U$12073 ( \12205 , \11957 , \11966 );
or \U$12074 ( \12206 , \12203 , \12204 , \12205 );
and \U$12075 ( \12207 , \11971 , \11975 );
and \U$12076 ( \12208 , \11975 , \11980 );
and \U$12077 ( \12209 , \11971 , \11980 );
or \U$12078 ( \12210 , \12207 , \12208 , \12209 );
xor \U$12079 ( \12211 , \12206 , \12210 );
and \U$12080 ( \12212 , \11986 , \11990 );
and \U$12081 ( \12213 , \11990 , \11995 );
and \U$12082 ( \12214 , \11986 , \11995 );
or \U$12083 ( \12215 , \12212 , \12213 , \12214 );
xor \U$12084 ( \12216 , \12211 , \12215 );
and \U$12085 ( \12217 , \11967 , \11981 );
and \U$12086 ( \12218 , \11981 , \11996 );
and \U$12087 ( \12219 , \11967 , \11996 );
or \U$12088 ( \12220 , \12217 , \12218 , \12219 );
and \U$12089 ( \12221 , \12108 , \12152 );
and \U$12090 ( \12222 , \12152 , \12175 );
and \U$12091 ( \12223 , \12108 , \12175 );
or \U$12092 ( \12224 , \12221 , \12222 , \12223 );
xor \U$12093 ( \12225 , \12220 , \12224 );
and \U$12094 ( \12226 , \12112 , \12116 );
and \U$12095 ( \12227 , \12116 , \12121 );
and \U$12096 ( \12228 , \12112 , \12121 );
or \U$12097 ( \12229 , \12226 , \12227 , \12228 );
and \U$12098 ( \12230 , \12126 , \12130 );
and \U$12099 ( \12231 , \12130 , \12135 );
and \U$12100 ( \12232 , \12126 , \12135 );
or \U$12101 ( \12233 , \12230 , \12231 , \12232 );
xor \U$12102 ( \12234 , \12229 , \12233 );
and \U$12103 ( \12235 , \12141 , \12145 );
and \U$12104 ( \12236 , \12145 , \12150 );
and \U$12105 ( \12237 , \12141 , \12150 );
or \U$12106 ( \12238 , \12235 , \12236 , \12237 );
xor \U$12107 ( \12239 , \12234 , \12238 );
and \U$12108 ( \12240 , \12022 , \12026 );
and \U$12109 ( \12241 , \12026 , \12031 );
and \U$12110 ( \12242 , \12022 , \12031 );
or \U$12111 ( \12243 , \12240 , \12241 , \12242 );
and \U$12112 ( \12244 , \12036 , \12040 );
and \U$12113 ( \12245 , \12040 , \12045 );
and \U$12114 ( \12246 , \12036 , \12045 );
or \U$12115 ( \12247 , \12244 , \12245 , \12246 );
xor \U$12116 ( \12248 , \12243 , \12247 );
and \U$12117 ( \12249 , \12051 , \12055 );
and \U$12118 ( \12250 , \12055 , \12060 );
and \U$12119 ( \12251 , \12051 , \12060 );
or \U$12120 ( \12252 , \12249 , \12250 , \12251 );
xor \U$12121 ( \12253 , \12248 , \12252 );
xor \U$12122 ( \12254 , \12239 , \12253 );
and \U$12123 ( \12255 , \12068 , \12072 );
and \U$12124 ( \12256 , \12072 , \12077 );
and \U$12125 ( \12257 , \12068 , \12077 );
or \U$12126 ( \12258 , \12255 , \12256 , \12257 );
and \U$12127 ( \12259 , \12082 , \12086 );
and \U$12128 ( \12260 , \12086 , \12091 );
and \U$12129 ( \12261 , \12082 , \12091 );
or \U$12130 ( \12262 , \12259 , \12260 , \12261 );
xor \U$12131 ( \12263 , \12258 , \12262 );
and \U$12132 ( \12264 , \12097 , \12101 );
and \U$12133 ( \12265 , \12101 , \12106 );
and \U$12134 ( \12266 , \12097 , \12106 );
or \U$12135 ( \12267 , \12264 , \12265 , \12266 );
xor \U$12136 ( \12268 , \12263 , \12267 );
xor \U$12137 ( \12269 , \12254 , \12268 );
xor \U$12138 ( \12270 , \12225 , \12269 );
xor \U$12139 ( \12271 , \12216 , \12270 );
and \U$12140 ( \12272 , \12078 , \12092 );
and \U$12141 ( \12273 , \12092 , \12107 );
and \U$12142 ( \12274 , \12078 , \12107 );
or \U$12143 ( \12275 , \12272 , \12273 , \12274 );
and \U$12144 ( \12276 , \12122 , \12136 );
and \U$12145 ( \12277 , \12136 , \12151 );
and \U$12146 ( \12278 , \12122 , \12151 );
or \U$12147 ( \12279 , \12276 , \12277 , \12278 );
xor \U$12148 ( \12280 , \12275 , \12279 );
and \U$12149 ( \12281 , \12157 , \12171 );
and \U$12150 ( \12282 , \12171 , \12174 );
and \U$12151 ( \12283 , \12157 , \12174 );
or \U$12152 ( \12284 , \12281 , \12282 , \12283 );
xor \U$12153 ( \12285 , \12280 , \12284 );
and \U$12154 ( \12286 , \12161 , \12165 );
and \U$12155 ( \12287 , \12165 , \12170 );
and \U$12156 ( \12288 , \12161 , \12170 );
or \U$12157 ( \12289 , \12286 , \12287 , \12288 );
buf \U$12158 ( \12290 , \12173 );
xor \U$12159 ( \12291 , \12289 , \12290 );
and \U$12160 ( \12292 , \240 , \10118 );
xor \U$12161 ( \12293 , \12291 , \12292 );
and \U$12162 ( \12294 , \217 , \9333 );
and \U$12163 ( \12295 , \189 , \9006 );
nor \U$12164 ( \12296 , \12294 , \12295 );
xnor \U$12165 ( \12297 , \12296 , \8848 );
and \U$12166 ( \12298 , \232 , \9765 );
and \U$12167 ( \12299 , \209 , \9644 );
nor \U$12168 ( \12300 , \12298 , \12299 );
xnor \U$12169 ( \12301 , \12300 , \9478 );
xor \U$12170 ( \12302 , \12297 , \12301 );
and \U$12171 ( \12303 , \247 , \10408 );
and \U$12172 ( \12304 , \224 , \10116 );
nor \U$12173 ( \12305 , \12303 , \12304 );
xnor \U$12174 ( \12306 , \12305 , \10121 );
xor \U$12175 ( \12307 , \12302 , \12306 );
and \U$12176 ( \12308 , \307 , \7489 );
and \U$12177 ( \12309 , \412 , \7137 );
nor \U$12178 ( \12310 , \12308 , \12309 );
xnor \U$12179 ( \12311 , \12310 , \7142 );
and \U$12180 ( \12312 , \185 , \8019 );
and \U$12181 ( \12313 , \261 , \7830 );
nor \U$12182 ( \12314 , \12312 , \12313 );
xnor \U$12183 ( \12315 , \12314 , \7713 );
xor \U$12184 ( \12316 , \12311 , \12315 );
and \U$12185 ( \12317 , \197 , \8540 );
and \U$12186 ( \12318 , \178 , \8292 );
nor \U$12187 ( \12319 , \12317 , \12318 );
xnor \U$12188 ( \12320 , \12319 , \8297 );
xor \U$12189 ( \12321 , \12316 , \12320 );
xor \U$12190 ( \12322 , \12307 , \12321 );
and \U$12191 ( \12323 , \1484 , \5996 );
and \U$12192 ( \12324 , \1601 , \5695 );
nor \U$12193 ( \12325 , \12323 , \12324 );
xnor \U$12194 ( \12326 , \12325 , \5687 );
and \U$12195 ( \12327 , \1192 , \6401 );
and \U$12196 ( \12328 , \1333 , \6143 );
nor \U$12197 ( \12329 , \12327 , \12328 );
xnor \U$12198 ( \12330 , \12329 , \6148 );
xor \U$12199 ( \12331 , \12326 , \12330 );
and \U$12200 ( \12332 , \474 , \7055 );
and \U$12201 ( \12333 , \1147 , \6675 );
nor \U$12202 ( \12334 , \12332 , \12333 );
xnor \U$12203 ( \12335 , \12334 , \6680 );
xor \U$12204 ( \12336 , \12331 , \12335 );
xor \U$12205 ( \12337 , \12322 , \12336 );
xor \U$12206 ( \12338 , \12293 , \12337 );
and \U$12207 ( \12339 , \2182 , \4581 );
and \U$12208 ( \12340 , \2366 , \4424 );
nor \U$12209 ( \12341 , \12339 , \12340 );
xnor \U$12210 ( \12342 , \12341 , \4377 );
and \U$12211 ( \12343 , \1948 , \5011 );
and \U$12212 ( \12344 , \2090 , \4878 );
nor \U$12213 ( \12345 , \12343 , \12344 );
xnor \U$12214 ( \12346 , \12345 , \4762 );
xor \U$12215 ( \12347 , \12342 , \12346 );
and \U$12216 ( \12348 , \1684 , \5485 );
and \U$12217 ( \12349 , \1802 , \5275 );
nor \U$12218 ( \12350 , \12348 , \12349 );
xnor \U$12219 ( \12351 , \12350 , \5169 );
xor \U$12220 ( \12352 , \12347 , \12351 );
and \U$12221 ( \12353 , \4364 , \2400 );
and \U$12222 ( \12354 , \4654 , \2246 );
nor \U$12223 ( \12355 , \12353 , \12354 );
xnor \U$12224 ( \12356 , \12355 , \2195 );
and \U$12225 ( \12357 , \3912 , \2669 );
and \U$12226 ( \12358 , \4160 , \2538 );
nor \U$12227 ( \12359 , \12357 , \12358 );
xnor \U$12228 ( \12360 , \12359 , \2534 );
xor \U$12229 ( \12361 , \12356 , \12360 );
and \U$12230 ( \12362 , \3646 , \3103 );
and \U$12231 ( \12363 , \3736 , \2934 );
nor \U$12232 ( \12364 , \12362 , \12363 );
xnor \U$12233 ( \12365 , \12364 , \2839 );
xor \U$12234 ( \12366 , \12361 , \12365 );
xor \U$12235 ( \12367 , \12352 , \12366 );
and \U$12236 ( \12368 , \3143 , \3357 );
and \U$12237 ( \12369 , \3395 , \3255 );
nor \U$12238 ( \12370 , \12368 , \12369 );
xnor \U$12239 ( \12371 , \12370 , \3156 );
and \U$12240 ( \12372 , \2826 , \3813 );
and \U$12241 ( \12373 , \3037 , \3557 );
nor \U$12242 ( \12374 , \12372 , \12373 );
xnor \U$12243 ( \12375 , \12374 , \3562 );
xor \U$12244 ( \12376 , \12371 , \12375 );
and \U$12245 ( \12377 , \2521 , \4132 );
and \U$12246 ( \12378 , \2757 , \4012 );
nor \U$12247 ( \12379 , \12377 , \12378 );
xnor \U$12248 ( \12380 , \12379 , \3925 );
xor \U$12249 ( \12381 , \12376 , \12380 );
xor \U$12250 ( \12382 , \12367 , \12381 );
xor \U$12251 ( \12383 , \12338 , \12382 );
xor \U$12252 ( \12384 , \12285 , \12383 );
and \U$12253 ( \12385 , \12032 , \12046 );
and \U$12254 ( \12386 , \12046 , \12061 );
and \U$12255 ( \12387 , \12032 , \12061 );
or \U$12256 ( \12388 , \12385 , \12386 , \12387 );
not \U$12257 ( \12389 , \222 );
and \U$12258 ( \12390 , \10206 , \230 );
and \U$12259 ( \12391 , \10584 , \228 );
nor \U$12260 ( \12392 , \12390 , \12391 );
xnor \U$12261 ( \12393 , \12392 , \237 );
xor \U$12262 ( \12394 , \12389 , \12393 );
and \U$12263 ( \12395 , \9465 , \245 );
and \U$12264 ( \12396 , \9897 , \243 );
nor \U$12265 ( \12397 , \12395 , \12396 );
xnor \U$12266 ( \12398 , \12397 , \252 );
xor \U$12267 ( \12399 , \12394 , \12398 );
xor \U$12268 ( \12400 , \12388 , \12399 );
and \U$12269 ( \12401 , \7231 , \438 );
and \U$12270 ( \12402 , \7556 , \336 );
nor \U$12271 ( \12403 , \12401 , \12402 );
xnor \U$12272 ( \12404 , \12403 , \320 );
and \U$12273 ( \12405 , \6790 , \1086 );
and \U$12274 ( \12406 , \6945 , \508 );
nor \U$12275 ( \12407 , \12405 , \12406 );
xnor \U$12276 ( \12408 , \12407 , \487 );
xor \U$12277 ( \12409 , \12404 , \12408 );
and \U$12278 ( \12410 , \6281 , \1301 );
and \U$12279 ( \12411 , \6514 , \1246 );
nor \U$12280 ( \12412 , \12410 , \12411 );
xnor \U$12281 ( \12413 , \12412 , \1205 );
xor \U$12282 ( \12414 , \12409 , \12413 );
and \U$12283 ( \12415 , \8835 , \141 );
and \U$12284 ( \12416 , \9169 , \139 );
nor \U$12285 ( \12417 , \12415 , \12416 );
xnor \U$12286 ( \12418 , \12417 , \148 );
and \U$12287 ( \12419 , \8349 , \156 );
and \U$12288 ( \12420 , \8652 , \154 );
nor \U$12289 ( \12421 , \12419 , \12420 );
xnor \U$12290 ( \12422 , \12421 , \163 );
xor \U$12291 ( \12423 , \12418 , \12422 );
and \U$12292 ( \12424 , \7700 , \296 );
and \U$12293 ( \12425 , \8057 , \168 );
nor \U$12294 ( \12426 , \12424 , \12425 );
xnor \U$12295 ( \12427 , \12426 , \173 );
xor \U$12296 ( \12428 , \12423 , \12427 );
xor \U$12297 ( \12429 , \12414 , \12428 );
and \U$12298 ( \12430 , \5674 , \1578 );
and \U$12299 ( \12431 , \6030 , \1431 );
nor \U$12300 ( \12432 , \12430 , \12431 );
xnor \U$12301 ( \12433 , \12432 , \1436 );
and \U$12302 ( \12434 , \5156 , \1824 );
and \U$12303 ( \12435 , \5469 , \1739 );
nor \U$12304 ( \12436 , \12434 , \12435 );
xnor \U$12305 ( \12437 , \12436 , \1697 );
xor \U$12306 ( \12438 , \12433 , \12437 );
and \U$12307 ( \12439 , \4749 , \2121 );
and \U$12308 ( \12440 , \4922 , \2008 );
nor \U$12309 ( \12441 , \12439 , \12440 );
xnor \U$12310 ( \12442 , \12441 , \1961 );
xor \U$12311 ( \12443 , \12438 , \12442 );
xor \U$12312 ( \12444 , \12429 , \12443 );
xor \U$12313 ( \12445 , \12400 , \12444 );
xor \U$12314 ( \12446 , \12384 , \12445 );
xor \U$12315 ( \12447 , \12271 , \12446 );
xor \U$12316 ( \12448 , \12202 , \12447 );
xor \U$12317 ( \12449 , \12196 , \12448 );
and \U$12318 ( \12450 , \11904 , \11908 );
and \U$12319 ( \12451 , \11908 , \11913 );
and \U$12320 ( \12452 , \11904 , \11913 );
or \U$12321 ( \12453 , \12450 , \12451 , \12452 );
and \U$12322 ( \12454 , \11948 , \11952 );
and \U$12323 ( \12455 , \11952 , \11997 );
and \U$12324 ( \12456 , \11948 , \11997 );
or \U$12325 ( \12457 , \12454 , \12455 , \12456 );
xor \U$12326 ( \12458 , \12453 , \12457 );
and \U$12327 ( \12459 , \12013 , \12063 );
and \U$12328 ( \12460 , \12063 , \12176 );
and \U$12329 ( \12461 , \12013 , \12176 );
or \U$12330 ( \12462 , \12459 , \12460 , \12461 );
xor \U$12331 ( \12463 , \12458 , \12462 );
and \U$12332 ( \12464 , \11920 , \11924 );
and \U$12333 ( \12465 , \11924 , \11929 );
and \U$12334 ( \12466 , \11920 , \11929 );
or \U$12335 ( \12467 , \12464 , \12465 , \12466 );
and \U$12336 ( \12468 , \11944 , \11998 );
and \U$12337 ( \12469 , \11998 , \12177 );
and \U$12338 ( \12470 , \11944 , \12177 );
or \U$12339 ( \12471 , \12468 , \12469 , \12470 );
xor \U$12340 ( \12472 , \12467 , \12471 );
and \U$12341 ( \12473 , \11934 , \11938 );
and \U$12342 ( \12474 , \11938 , \11943 );
and \U$12343 ( \12475 , \11934 , \11943 );
or \U$12344 ( \12476 , \12473 , \12474 , \12475 );
and \U$12345 ( \12477 , \12003 , \12007 );
and \U$12346 ( \12478 , \12007 , \12012 );
and \U$12347 ( \12479 , \12003 , \12012 );
or \U$12348 ( \12480 , \12477 , \12478 , \12479 );
xor \U$12349 ( \12481 , \12476 , \12480 );
and \U$12350 ( \12482 , \12017 , \12018 );
and \U$12351 ( \12483 , \12018 , \12062 );
and \U$12352 ( \12484 , \12017 , \12062 );
or \U$12353 ( \12485 , \12482 , \12483 , \12484 );
xor \U$12354 ( \12486 , \12481 , \12485 );
xor \U$12355 ( \12487 , \12472 , \12486 );
xor \U$12356 ( \12488 , \12463 , \12487 );
xor \U$12357 ( \12489 , \12449 , \12488 );
and \U$12358 ( \12490 , \11885 , \11886 );
and \U$12359 ( \12491 , \11886 , \12180 );
and \U$12360 ( \12492 , \11885 , \12180 );
or \U$12361 ( \12493 , \12490 , \12491 , \12492 );
xor \U$12362 ( \12494 , \12489 , \12493 );
and \U$12363 ( \12495 , \12181 , \12185 );
and \U$12364 ( \12496 , \12186 , \12189 );
or \U$12365 ( \12497 , \12495 , \12496 );
xor \U$12366 ( \12498 , \12494 , \12497 );
buf \U$12367 ( \12499 , \12498 );
buf \U$12368 ( \12500 , \12499 );
and \U$12369 ( \12501 , \12200 , \12201 );
and \U$12370 ( \12502 , \12201 , \12447 );
and \U$12371 ( \12503 , \12200 , \12447 );
or \U$12372 ( \12504 , \12501 , \12502 , \12503 );
and \U$12373 ( \12505 , \12463 , \12487 );
xor \U$12374 ( \12506 , \12504 , \12505 );
and \U$12375 ( \12507 , \12467 , \12471 );
and \U$12376 ( \12508 , \12471 , \12486 );
and \U$12377 ( \12509 , \12467 , \12486 );
or \U$12378 ( \12510 , \12507 , \12508 , \12509 );
and \U$12379 ( \12511 , \12453 , \12457 );
and \U$12380 ( \12512 , \12457 , \12462 );
and \U$12381 ( \12513 , \12453 , \12462 );
or \U$12382 ( \12514 , \12511 , \12512 , \12513 );
and \U$12383 ( \12515 , \12216 , \12270 );
and \U$12384 ( \12516 , \12270 , \12446 );
and \U$12385 ( \12517 , \12216 , \12446 );
or \U$12386 ( \12518 , \12515 , \12516 , \12517 );
xor \U$12387 ( \12519 , \12514 , \12518 );
and \U$12388 ( \12520 , \12239 , \12253 );
and \U$12389 ( \12521 , \12253 , \12268 );
and \U$12390 ( \12522 , \12239 , \12268 );
or \U$12391 ( \12523 , \12520 , \12521 , \12522 );
and \U$12392 ( \12524 , \12293 , \12337 );
and \U$12393 ( \12525 , \12337 , \12382 );
and \U$12394 ( \12526 , \12293 , \12382 );
or \U$12395 ( \12527 , \12524 , \12525 , \12526 );
xor \U$12396 ( \12528 , \12523 , \12527 );
and \U$12397 ( \12529 , \12356 , \12360 );
and \U$12398 ( \12530 , \12360 , \12365 );
and \U$12399 ( \12531 , \12356 , \12365 );
or \U$12400 ( \12532 , \12529 , \12530 , \12531 );
and \U$12401 ( \12533 , \12371 , \12375 );
and \U$12402 ( \12534 , \12375 , \12380 );
and \U$12403 ( \12535 , \12371 , \12380 );
or \U$12404 ( \12536 , \12533 , \12534 , \12535 );
xor \U$12405 ( \12537 , \12532 , \12536 );
and \U$12406 ( \12538 , \12433 , \12437 );
and \U$12407 ( \12539 , \12437 , \12442 );
and \U$12408 ( \12540 , \12433 , \12442 );
or \U$12409 ( \12541 , \12538 , \12539 , \12540 );
xor \U$12410 ( \12542 , \12537 , \12541 );
xor \U$12411 ( \12543 , \12528 , \12542 );
xor \U$12412 ( \12544 , \12519 , \12543 );
xor \U$12413 ( \12545 , \12510 , \12544 );
and \U$12414 ( \12546 , \12206 , \12210 );
and \U$12415 ( \12547 , \12210 , \12215 );
and \U$12416 ( \12548 , \12206 , \12215 );
or \U$12417 ( \12549 , \12546 , \12547 , \12548 );
and \U$12418 ( \12550 , \12275 , \12279 );
and \U$12419 ( \12551 , \12279 , \12284 );
and \U$12420 ( \12552 , \12275 , \12284 );
or \U$12421 ( \12553 , \12550 , \12551 , \12552 );
xor \U$12422 ( \12554 , \12549 , \12553 );
and \U$12423 ( \12555 , \12388 , \12399 );
and \U$12424 ( \12556 , \12399 , \12444 );
and \U$12425 ( \12557 , \12388 , \12444 );
or \U$12426 ( \12558 , \12555 , \12556 , \12557 );
xor \U$12427 ( \12559 , \12554 , \12558 );
and \U$12428 ( \12560 , \12476 , \12480 );
and \U$12429 ( \12561 , \12480 , \12485 );
and \U$12430 ( \12562 , \12476 , \12485 );
or \U$12431 ( \12563 , \12560 , \12561 , \12562 );
and \U$12432 ( \12564 , \12220 , \12224 );
and \U$12433 ( \12565 , \12224 , \12269 );
and \U$12434 ( \12566 , \12220 , \12269 );
or \U$12435 ( \12567 , \12564 , \12565 , \12566 );
xor \U$12436 ( \12568 , \12563 , \12567 );
and \U$12437 ( \12569 , \12285 , \12383 );
and \U$12438 ( \12570 , \12383 , \12445 );
and \U$12439 ( \12571 , \12285 , \12445 );
or \U$12440 ( \12572 , \12569 , \12570 , \12571 );
xor \U$12441 ( \12573 , \12568 , \12572 );
xor \U$12442 ( \12574 , \12559 , \12573 );
and \U$12443 ( \12575 , \12229 , \12233 );
and \U$12444 ( \12576 , \12233 , \12238 );
and \U$12445 ( \12577 , \12229 , \12238 );
or \U$12446 ( \12578 , \12575 , \12576 , \12577 );
and \U$12447 ( \12579 , \12243 , \12247 );
and \U$12448 ( \12580 , \12247 , \12252 );
and \U$12449 ( \12581 , \12243 , \12252 );
or \U$12450 ( \12582 , \12579 , \12580 , \12581 );
xor \U$12451 ( \12583 , \12578 , \12582 );
and \U$12452 ( \12584 , \12258 , \12262 );
and \U$12453 ( \12585 , \12262 , \12267 );
and \U$12454 ( \12586 , \12258 , \12267 );
or \U$12455 ( \12587 , \12584 , \12585 , \12586 );
xor \U$12456 ( \12588 , \12583 , \12587 );
and \U$12457 ( \12589 , \12289 , \12290 );
and \U$12458 ( \12590 , \12290 , \12292 );
and \U$12459 ( \12591 , \12289 , \12292 );
or \U$12460 ( \12592 , \12589 , \12590 , \12591 );
and \U$12461 ( \12593 , \12307 , \12321 );
and \U$12462 ( \12594 , \12321 , \12336 );
and \U$12463 ( \12595 , \12307 , \12336 );
or \U$12464 ( \12596 , \12593 , \12594 , \12595 );
xor \U$12465 ( \12597 , \12592 , \12596 );
and \U$12466 ( \12598 , \12352 , \12366 );
and \U$12467 ( \12599 , \12366 , \12381 );
and \U$12468 ( \12600 , \12352 , \12381 );
or \U$12469 ( \12601 , \12598 , \12599 , \12600 );
xor \U$12470 ( \12602 , \12597 , \12601 );
xor \U$12471 ( \12603 , \12588 , \12602 );
and \U$12472 ( \12604 , \12389 , \12393 );
and \U$12473 ( \12605 , \12393 , \12398 );
and \U$12474 ( \12606 , \12389 , \12398 );
or \U$12475 ( \12607 , \12604 , \12605 , \12606 );
and \U$12476 ( \12608 , \12404 , \12408 );
and \U$12477 ( \12609 , \12408 , \12413 );
and \U$12478 ( \12610 , \12404 , \12413 );
or \U$12479 ( \12611 , \12608 , \12609 , \12610 );
xor \U$12480 ( \12612 , \12607 , \12611 );
and \U$12481 ( \12613 , \12418 , \12422 );
and \U$12482 ( \12614 , \12422 , \12427 );
and \U$12483 ( \12615 , \12418 , \12427 );
or \U$12484 ( \12616 , \12613 , \12614 , \12615 );
xor \U$12485 ( \12617 , \12612 , \12616 );
and \U$12486 ( \12618 , \12414 , \12428 );
and \U$12487 ( \12619 , \12428 , \12443 );
and \U$12488 ( \12620 , \12414 , \12443 );
or \U$12489 ( \12621 , \12618 , \12619 , \12620 );
and \U$12490 ( \12622 , \10584 , \230 );
not \U$12491 ( \12623 , \12622 );
xnor \U$12492 ( \12624 , \12623 , \237 );
and \U$12493 ( \12625 , \9897 , \245 );
and \U$12494 ( \12626 , \10206 , \243 );
nor \U$12495 ( \12627 , \12625 , \12626 );
xnor \U$12496 ( \12628 , \12627 , \252 );
xor \U$12497 ( \12629 , \12624 , \12628 );
and \U$12498 ( \12630 , \9169 , \141 );
and \U$12499 ( \12631 , \9465 , \139 );
nor \U$12500 ( \12632 , \12630 , \12631 );
xnor \U$12501 ( \12633 , \12632 , \148 );
xor \U$12502 ( \12634 , \12629 , \12633 );
and \U$12503 ( \12635 , \6945 , \1086 );
and \U$12504 ( \12636 , \7231 , \508 );
nor \U$12505 ( \12637 , \12635 , \12636 );
xnor \U$12506 ( \12638 , \12637 , \487 );
and \U$12507 ( \12639 , \6514 , \1301 );
and \U$12508 ( \12640 , \6790 , \1246 );
nor \U$12509 ( \12641 , \12639 , \12640 );
xnor \U$12510 ( \12642 , \12641 , \1205 );
xor \U$12511 ( \12643 , \12638 , \12642 );
and \U$12512 ( \12644 , \6030 , \1578 );
and \U$12513 ( \12645 , \6281 , \1431 );
nor \U$12514 ( \12646 , \12644 , \12645 );
xnor \U$12515 ( \12647 , \12646 , \1436 );
xor \U$12516 ( \12648 , \12643 , \12647 );
xor \U$12517 ( \12649 , \12634 , \12648 );
and \U$12518 ( \12650 , \8652 , \156 );
and \U$12519 ( \12651 , \8835 , \154 );
nor \U$12520 ( \12652 , \12650 , \12651 );
xnor \U$12521 ( \12653 , \12652 , \163 );
and \U$12522 ( \12654 , \8057 , \296 );
and \U$12523 ( \12655 , \8349 , \168 );
nor \U$12524 ( \12656 , \12654 , \12655 );
xnor \U$12525 ( \12657 , \12656 , \173 );
xor \U$12526 ( \12658 , \12653 , \12657 );
and \U$12527 ( \12659 , \7556 , \438 );
and \U$12528 ( \12660 , \7700 , \336 );
nor \U$12529 ( \12661 , \12659 , \12660 );
xnor \U$12530 ( \12662 , \12661 , \320 );
xor \U$12531 ( \12663 , \12658 , \12662 );
xor \U$12532 ( \12664 , \12649 , \12663 );
xor \U$12533 ( \12665 , \12621 , \12664 );
and \U$12534 ( \12666 , \3037 , \3813 );
and \U$12535 ( \12667 , \3143 , \3557 );
nor \U$12536 ( \12668 , \12666 , \12667 );
xnor \U$12537 ( \12669 , \12668 , \3562 );
and \U$12538 ( \12670 , \2757 , \4132 );
and \U$12539 ( \12671 , \2826 , \4012 );
nor \U$12540 ( \12672 , \12670 , \12671 );
xnor \U$12541 ( \12673 , \12672 , \3925 );
xor \U$12542 ( \12674 , \12669 , \12673 );
and \U$12543 ( \12675 , \2366 , \4581 );
and \U$12544 ( \12676 , \2521 , \4424 );
nor \U$12545 ( \12677 , \12675 , \12676 );
xnor \U$12546 ( \12678 , \12677 , \4377 );
xor \U$12547 ( \12679 , \12674 , \12678 );
and \U$12548 ( \12680 , \5469 , \1824 );
and \U$12549 ( \12681 , \5674 , \1739 );
nor \U$12550 ( \12682 , \12680 , \12681 );
xnor \U$12551 ( \12683 , \12682 , \1697 );
and \U$12552 ( \12684 , \4922 , \2121 );
and \U$12553 ( \12685 , \5156 , \2008 );
nor \U$12554 ( \12686 , \12684 , \12685 );
xnor \U$12555 ( \12687 , \12686 , \1961 );
xor \U$12556 ( \12688 , \12683 , \12687 );
and \U$12557 ( \12689 , \4654 , \2400 );
and \U$12558 ( \12690 , \4749 , \2246 );
nor \U$12559 ( \12691 , \12689 , \12690 );
xnor \U$12560 ( \12692 , \12691 , \2195 );
xor \U$12561 ( \12693 , \12688 , \12692 );
xor \U$12562 ( \12694 , \12679 , \12693 );
and \U$12563 ( \12695 , \4160 , \2669 );
and \U$12564 ( \12696 , \4364 , \2538 );
nor \U$12565 ( \12697 , \12695 , \12696 );
xnor \U$12566 ( \12698 , \12697 , \2534 );
and \U$12567 ( \12699 , \3736 , \3103 );
and \U$12568 ( \12700 , \3912 , \2934 );
nor \U$12569 ( \12701 , \12699 , \12700 );
xnor \U$12570 ( \12702 , \12701 , \2839 );
xor \U$12571 ( \12703 , \12698 , \12702 );
and \U$12572 ( \12704 , \3395 , \3357 );
and \U$12573 ( \12705 , \3646 , \3255 );
nor \U$12574 ( \12706 , \12704 , \12705 );
xnor \U$12575 ( \12707 , \12706 , \3156 );
xor \U$12576 ( \12708 , \12703 , \12707 );
xor \U$12577 ( \12709 , \12694 , \12708 );
xor \U$12578 ( \12710 , \12665 , \12709 );
xor \U$12579 ( \12711 , \12617 , \12710 );
and \U$12580 ( \12712 , \12311 , \12315 );
and \U$12581 ( \12713 , \12315 , \12320 );
and \U$12582 ( \12714 , \12311 , \12320 );
or \U$12583 ( \12715 , \12712 , \12713 , \12714 );
and \U$12584 ( \12716 , \12326 , \12330 );
and \U$12585 ( \12717 , \12330 , \12335 );
and \U$12586 ( \12718 , \12326 , \12335 );
or \U$12587 ( \12719 , \12716 , \12717 , \12718 );
xor \U$12588 ( \12720 , \12715 , \12719 );
and \U$12589 ( \12721 , \12342 , \12346 );
and \U$12590 ( \12722 , \12346 , \12351 );
and \U$12591 ( \12723 , \12342 , \12351 );
or \U$12592 ( \12724 , \12721 , \12722 , \12723 );
xor \U$12593 ( \12725 , \12720 , \12724 );
and \U$12594 ( \12726 , \261 , \8019 );
and \U$12595 ( \12727 , \307 , \7830 );
nor \U$12596 ( \12728 , \12726 , \12727 );
xnor \U$12597 ( \12729 , \12728 , \7713 );
and \U$12598 ( \12730 , \178 , \8540 );
and \U$12599 ( \12731 , \185 , \8292 );
nor \U$12600 ( \12732 , \12730 , \12731 );
xnor \U$12601 ( \12733 , \12732 , \8297 );
xor \U$12602 ( \12734 , \12729 , \12733 );
and \U$12603 ( \12735 , \189 , \9333 );
and \U$12604 ( \12736 , \197 , \9006 );
nor \U$12605 ( \12737 , \12735 , \12736 );
xnor \U$12606 ( \12738 , \12737 , \8848 );
xor \U$12607 ( \12739 , \12734 , \12738 );
and \U$12608 ( \12740 , \1333 , \6401 );
and \U$12609 ( \12741 , \1484 , \6143 );
nor \U$12610 ( \12742 , \12740 , \12741 );
xnor \U$12611 ( \12743 , \12742 , \6148 );
and \U$12612 ( \12744 , \1147 , \7055 );
and \U$12613 ( \12745 , \1192 , \6675 );
nor \U$12614 ( \12746 , \12744 , \12745 );
xnor \U$12615 ( \12747 , \12746 , \6680 );
xor \U$12616 ( \12748 , \12743 , \12747 );
and \U$12617 ( \12749 , \412 , \7489 );
and \U$12618 ( \12750 , \474 , \7137 );
nor \U$12619 ( \12751 , \12749 , \12750 );
xnor \U$12620 ( \12752 , \12751 , \7142 );
xor \U$12621 ( \12753 , \12748 , \12752 );
xor \U$12622 ( \12754 , \12739 , \12753 );
and \U$12623 ( \12755 , \2090 , \5011 );
and \U$12624 ( \12756 , \2182 , \4878 );
nor \U$12625 ( \12757 , \12755 , \12756 );
xnor \U$12626 ( \12758 , \12757 , \4762 );
and \U$12627 ( \12759 , \1802 , \5485 );
and \U$12628 ( \12760 , \1948 , \5275 );
nor \U$12629 ( \12761 , \12759 , \12760 );
xnor \U$12630 ( \12762 , \12761 , \5169 );
xor \U$12631 ( \12763 , \12758 , \12762 );
and \U$12632 ( \12764 , \1601 , \5996 );
and \U$12633 ( \12765 , \1684 , \5695 );
nor \U$12634 ( \12766 , \12764 , \12765 );
xnor \U$12635 ( \12767 , \12766 , \5687 );
xor \U$12636 ( \12768 , \12763 , \12767 );
xor \U$12637 ( \12769 , \12754 , \12768 );
xor \U$12638 ( \12770 , \12725 , \12769 );
and \U$12639 ( \12771 , \12297 , \12301 );
and \U$12640 ( \12772 , \12301 , \12306 );
and \U$12641 ( \12773 , \12297 , \12306 );
or \U$12642 ( \12774 , \12771 , \12772 , \12773 );
and \U$12643 ( \12775 , \209 , \9765 );
and \U$12644 ( \12776 , \217 , \9644 );
nor \U$12645 ( \12777 , \12775 , \12776 );
xnor \U$12646 ( \12778 , \12777 , \9478 );
and \U$12647 ( \12779 , \224 , \10408 );
and \U$12648 ( \12780 , \232 , \10116 );
nor \U$12649 ( \12781 , \12779 , \12780 );
xnor \U$12650 ( \12782 , \12781 , \10121 );
xor \U$12651 ( \12783 , \12778 , \12782 );
and \U$12652 ( \12784 , \247 , \10118 );
xor \U$12653 ( \12785 , \12783 , \12784 );
xnor \U$12654 ( \12786 , \12774 , \12785 );
xor \U$12655 ( \12787 , \12770 , \12786 );
xor \U$12656 ( \12788 , \12711 , \12787 );
xor \U$12657 ( \12789 , \12603 , \12788 );
xor \U$12658 ( \12790 , \12574 , \12789 );
xor \U$12659 ( \12791 , \12545 , \12790 );
xor \U$12660 ( \12792 , \12506 , \12791 );
and \U$12661 ( \12793 , \12196 , \12448 );
and \U$12662 ( \12794 , \12448 , \12488 );
and \U$12663 ( \12795 , \12196 , \12488 );
or \U$12664 ( \12796 , \12793 , \12794 , \12795 );
xor \U$12665 ( \12797 , \12792 , \12796 );
and \U$12666 ( \12798 , \12489 , \12493 );
and \U$12667 ( \12799 , \12494 , \12497 );
or \U$12668 ( \12800 , \12798 , \12799 );
xor \U$12669 ( \12801 , \12797 , \12800 );
buf \U$12670 ( \12802 , \12801 );
buf \U$12671 ( \12803 , \12802 );
and \U$12672 ( \12804 , \12510 , \12544 );
and \U$12673 ( \12805 , \12544 , \12790 );
and \U$12674 ( \12806 , \12510 , \12790 );
or \U$12675 ( \12807 , \12804 , \12805 , \12806 );
and \U$12676 ( \12808 , \12514 , \12518 );
and \U$12677 ( \12809 , \12518 , \12543 );
and \U$12678 ( \12810 , \12514 , \12543 );
or \U$12679 ( \12811 , \12808 , \12809 , \12810 );
and \U$12680 ( \12812 , \12559 , \12573 );
and \U$12681 ( \12813 , \12573 , \12789 );
and \U$12682 ( \12814 , \12559 , \12789 );
or \U$12683 ( \12815 , \12812 , \12813 , \12814 );
xor \U$12684 ( \12816 , \12811 , \12815 );
and \U$12685 ( \12817 , \12549 , \12553 );
and \U$12686 ( \12818 , \12553 , \12558 );
and \U$12687 ( \12819 , \12549 , \12558 );
or \U$12688 ( \12820 , \12817 , \12818 , \12819 );
and \U$12689 ( \12821 , \12523 , \12527 );
and \U$12690 ( \12822 , \12527 , \12542 );
and \U$12691 ( \12823 , \12523 , \12542 );
or \U$12692 ( \12824 , \12821 , \12822 , \12823 );
xor \U$12693 ( \12825 , \12820 , \12824 );
and \U$12694 ( \12826 , \12617 , \12710 );
and \U$12695 ( \12827 , \12710 , \12787 );
and \U$12696 ( \12828 , \12617 , \12787 );
or \U$12697 ( \12829 , \12826 , \12827 , \12828 );
xor \U$12698 ( \12830 , \12825 , \12829 );
xor \U$12699 ( \12831 , \12816 , \12830 );
xor \U$12700 ( \12832 , \12807 , \12831 );
and \U$12701 ( \12833 , \12563 , \12567 );
and \U$12702 ( \12834 , \12567 , \12572 );
and \U$12703 ( \12835 , \12563 , \12572 );
or \U$12704 ( \12836 , \12833 , \12834 , \12835 );
and \U$12705 ( \12837 , \12588 , \12602 );
and \U$12706 ( \12838 , \12602 , \12788 );
and \U$12707 ( \12839 , \12588 , \12788 );
or \U$12708 ( \12840 , \12837 , \12838 , \12839 );
xor \U$12709 ( \12841 , \12836 , \12840 );
and \U$12710 ( \12842 , \12578 , \12582 );
and \U$12711 ( \12843 , \12582 , \12587 );
and \U$12712 ( \12844 , \12578 , \12587 );
or \U$12713 ( \12845 , \12842 , \12843 , \12844 );
and \U$12714 ( \12846 , \12592 , \12596 );
and \U$12715 ( \12847 , \12596 , \12601 );
and \U$12716 ( \12848 , \12592 , \12601 );
or \U$12717 ( \12849 , \12846 , \12847 , \12848 );
xor \U$12718 ( \12850 , \12845 , \12849 );
and \U$12719 ( \12851 , \12621 , \12664 );
and \U$12720 ( \12852 , \12664 , \12709 );
and \U$12721 ( \12853 , \12621 , \12709 );
or \U$12722 ( \12854 , \12851 , \12852 , \12853 );
xor \U$12723 ( \12855 , \12850 , \12854 );
and \U$12724 ( \12856 , \12739 , \12753 );
and \U$12725 ( \12857 , \12753 , \12768 );
and \U$12726 ( \12858 , \12739 , \12768 );
or \U$12727 ( \12859 , \12856 , \12857 , \12858 );
and \U$12728 ( \12860 , \12679 , \12693 );
and \U$12729 ( \12861 , \12693 , \12708 );
and \U$12730 ( \12862 , \12679 , \12708 );
or \U$12731 ( \12863 , \12860 , \12861 , \12862 );
xor \U$12732 ( \12864 , \12859 , \12863 );
or \U$12733 ( \12865 , \12774 , \12785 );
xor \U$12734 ( \12866 , \12864 , \12865 );
and \U$12735 ( \12867 , \12607 , \12611 );
and \U$12736 ( \12868 , \12611 , \12616 );
and \U$12737 ( \12869 , \12607 , \12616 );
or \U$12738 ( \12870 , \12867 , \12868 , \12869 );
and \U$12739 ( \12871 , \12532 , \12536 );
and \U$12740 ( \12872 , \12536 , \12541 );
and \U$12741 ( \12873 , \12532 , \12541 );
or \U$12742 ( \12874 , \12871 , \12872 , \12873 );
xor \U$12743 ( \12875 , \12870 , \12874 );
and \U$12744 ( \12876 , \12715 , \12719 );
and \U$12745 ( \12877 , \12719 , \12724 );
and \U$12746 ( \12878 , \12715 , \12724 );
or \U$12747 ( \12879 , \12876 , \12877 , \12878 );
xor \U$12748 ( \12880 , \12875 , \12879 );
xor \U$12749 ( \12881 , \12866 , \12880 );
and \U$12750 ( \12882 , \12634 , \12648 );
and \U$12751 ( \12883 , \12648 , \12663 );
and \U$12752 ( \12884 , \12634 , \12663 );
or \U$12753 ( \12885 , \12882 , \12883 , \12884 );
and \U$12754 ( \12886 , \8835 , \156 );
and \U$12755 ( \12887 , \9169 , \154 );
nor \U$12756 ( \12888 , \12886 , \12887 );
xnor \U$12757 ( \12889 , \12888 , \163 );
and \U$12758 ( \12890 , \8349 , \296 );
and \U$12759 ( \12891 , \8652 , \168 );
nor \U$12760 ( \12892 , \12890 , \12891 );
xnor \U$12761 ( \12893 , \12892 , \173 );
xor \U$12762 ( \12894 , \12889 , \12893 );
and \U$12763 ( \12895 , \7700 , \438 );
and \U$12764 ( \12896 , \8057 , \336 );
nor \U$12765 ( \12897 , \12895 , \12896 );
xnor \U$12766 ( \12898 , \12897 , \320 );
xor \U$12767 ( \12899 , \12894 , \12898 );
xor \U$12768 ( \12900 , \12885 , \12899 );
not \U$12769 ( \12901 , \237 );
and \U$12770 ( \12902 , \10206 , \245 );
and \U$12771 ( \12903 , \10584 , \243 );
nor \U$12772 ( \12904 , \12902 , \12903 );
xnor \U$12773 ( \12905 , \12904 , \252 );
xor \U$12774 ( \12906 , \12901 , \12905 );
and \U$12775 ( \12907 , \9465 , \141 );
and \U$12776 ( \12908 , \9897 , \139 );
nor \U$12777 ( \12909 , \12907 , \12908 );
xnor \U$12778 ( \12910 , \12909 , \148 );
xor \U$12779 ( \12911 , \12906 , \12910 );
xor \U$12780 ( \12912 , \12900 , \12911 );
xor \U$12781 ( \12913 , \12881 , \12912 );
xor \U$12782 ( \12914 , \12855 , \12913 );
and \U$12783 ( \12915 , \12725 , \12769 );
and \U$12784 ( \12916 , \12769 , \12786 );
and \U$12785 ( \12917 , \12725 , \12786 );
or \U$12786 ( \12918 , \12915 , \12916 , \12917 );
and \U$12787 ( \12919 , \12669 , \12673 );
and \U$12788 ( \12920 , \12673 , \12678 );
and \U$12789 ( \12921 , \12669 , \12678 );
or \U$12790 ( \12922 , \12919 , \12920 , \12921 );
and \U$12791 ( \12923 , \12683 , \12687 );
and \U$12792 ( \12924 , \12687 , \12692 );
and \U$12793 ( \12925 , \12683 , \12692 );
or \U$12794 ( \12926 , \12923 , \12924 , \12925 );
xor \U$12795 ( \12927 , \12922 , \12926 );
and \U$12796 ( \12928 , \12698 , \12702 );
and \U$12797 ( \12929 , \12702 , \12707 );
and \U$12798 ( \12930 , \12698 , \12707 );
or \U$12799 ( \12931 , \12928 , \12929 , \12930 );
xor \U$12800 ( \12932 , \12927 , \12931 );
and \U$12801 ( \12933 , \12729 , \12733 );
and \U$12802 ( \12934 , \12733 , \12738 );
and \U$12803 ( \12935 , \12729 , \12738 );
or \U$12804 ( \12936 , \12933 , \12934 , \12935 );
and \U$12805 ( \12937 , \12743 , \12747 );
and \U$12806 ( \12938 , \12747 , \12752 );
and \U$12807 ( \12939 , \12743 , \12752 );
or \U$12808 ( \12940 , \12937 , \12938 , \12939 );
xor \U$12809 ( \12941 , \12936 , \12940 );
and \U$12810 ( \12942 , \12758 , \12762 );
and \U$12811 ( \12943 , \12762 , \12767 );
and \U$12812 ( \12944 , \12758 , \12767 );
or \U$12813 ( \12945 , \12942 , \12943 , \12944 );
xor \U$12814 ( \12946 , \12941 , \12945 );
xor \U$12815 ( \12947 , \12932 , \12946 );
and \U$12816 ( \12948 , \12624 , \12628 );
and \U$12817 ( \12949 , \12628 , \12633 );
and \U$12818 ( \12950 , \12624 , \12633 );
or \U$12819 ( \12951 , \12948 , \12949 , \12950 );
and \U$12820 ( \12952 , \12638 , \12642 );
and \U$12821 ( \12953 , \12642 , \12647 );
and \U$12822 ( \12954 , \12638 , \12647 );
or \U$12823 ( \12955 , \12952 , \12953 , \12954 );
xor \U$12824 ( \12956 , \12951 , \12955 );
and \U$12825 ( \12957 , \12653 , \12657 );
and \U$12826 ( \12958 , \12657 , \12662 );
and \U$12827 ( \12959 , \12653 , \12662 );
or \U$12828 ( \12960 , \12957 , \12958 , \12959 );
xor \U$12829 ( \12961 , \12956 , \12960 );
xor \U$12830 ( \12962 , \12947 , \12961 );
xor \U$12831 ( \12963 , \12918 , \12962 );
and \U$12832 ( \12964 , \7231 , \1086 );
and \U$12833 ( \12965 , \7556 , \508 );
nor \U$12834 ( \12966 , \12964 , \12965 );
xnor \U$12835 ( \12967 , \12966 , \487 );
and \U$12836 ( \12968 , \6790 , \1301 );
and \U$12837 ( \12969 , \6945 , \1246 );
nor \U$12838 ( \12970 , \12968 , \12969 );
xnor \U$12839 ( \12971 , \12970 , \1205 );
xor \U$12840 ( \12972 , \12967 , \12971 );
and \U$12841 ( \12973 , \6281 , \1578 );
and \U$12842 ( \12974 , \6514 , \1431 );
nor \U$12843 ( \12975 , \12973 , \12974 );
xnor \U$12844 ( \12976 , \12975 , \1436 );
xor \U$12845 ( \12977 , \12972 , \12976 );
and \U$12846 ( \12978 , \4364 , \2669 );
and \U$12847 ( \12979 , \4654 , \2538 );
nor \U$12848 ( \12980 , \12978 , \12979 );
xnor \U$12849 ( \12981 , \12980 , \2534 );
and \U$12850 ( \12982 , \3912 , \3103 );
and \U$12851 ( \12983 , \4160 , \2934 );
nor \U$12852 ( \12984 , \12982 , \12983 );
xnor \U$12853 ( \12985 , \12984 , \2839 );
xor \U$12854 ( \12986 , \12981 , \12985 );
and \U$12855 ( \12987 , \3646 , \3357 );
and \U$12856 ( \12988 , \3736 , \3255 );
nor \U$12857 ( \12989 , \12987 , \12988 );
xnor \U$12858 ( \12990 , \12989 , \3156 );
xor \U$12859 ( \12991 , \12986 , \12990 );
xor \U$12860 ( \12992 , \12977 , \12991 );
and \U$12861 ( \12993 , \5674 , \1824 );
and \U$12862 ( \12994 , \6030 , \1739 );
nor \U$12863 ( \12995 , \12993 , \12994 );
xnor \U$12864 ( \12996 , \12995 , \1697 );
and \U$12865 ( \12997 , \5156 , \2121 );
and \U$12866 ( \12998 , \5469 , \2008 );
nor \U$12867 ( \12999 , \12997 , \12998 );
xnor \U$12868 ( \13000 , \12999 , \1961 );
xor \U$12869 ( \13001 , \12996 , \13000 );
and \U$12870 ( \13002 , \4749 , \2400 );
and \U$12871 ( \13003 , \4922 , \2246 );
nor \U$12872 ( \13004 , \13002 , \13003 );
xnor \U$12873 ( \13005 , \13004 , \2195 );
xor \U$12874 ( \13006 , \13001 , \13005 );
xor \U$12875 ( \13007 , \12992 , \13006 );
and \U$12876 ( \13008 , \3143 , \3813 );
and \U$12877 ( \13009 , \3395 , \3557 );
nor \U$12878 ( \13010 , \13008 , \13009 );
xnor \U$12879 ( \13011 , \13010 , \3562 );
and \U$12880 ( \13012 , \2826 , \4132 );
and \U$12881 ( \13013 , \3037 , \4012 );
nor \U$12882 ( \13014 , \13012 , \13013 );
xnor \U$12883 ( \13015 , \13014 , \3925 );
xor \U$12884 ( \13016 , \13011 , \13015 );
and \U$12885 ( \13017 , \2521 , \4581 );
and \U$12886 ( \13018 , \2757 , \4424 );
nor \U$12887 ( \13019 , \13017 , \13018 );
xnor \U$12888 ( \13020 , \13019 , \4377 );
xor \U$12889 ( \13021 , \13016 , \13020 );
and \U$12890 ( \13022 , \1484 , \6401 );
and \U$12891 ( \13023 , \1601 , \6143 );
nor \U$12892 ( \13024 , \13022 , \13023 );
xnor \U$12893 ( \13025 , \13024 , \6148 );
and \U$12894 ( \13026 , \1192 , \7055 );
and \U$12895 ( \13027 , \1333 , \6675 );
nor \U$12896 ( \13028 , \13026 , \13027 );
xnor \U$12897 ( \13029 , \13028 , \6680 );
xor \U$12898 ( \13030 , \13025 , \13029 );
and \U$12899 ( \13031 , \474 , \7489 );
and \U$12900 ( \13032 , \1147 , \7137 );
nor \U$12901 ( \13033 , \13031 , \13032 );
xnor \U$12902 ( \13034 , \13033 , \7142 );
xor \U$12903 ( \13035 , \13030 , \13034 );
xor \U$12904 ( \13036 , \13021 , \13035 );
and \U$12905 ( \13037 , \2182 , \5011 );
and \U$12906 ( \13038 , \2366 , \4878 );
nor \U$12907 ( \13039 , \13037 , \13038 );
xnor \U$12908 ( \13040 , \13039 , \4762 );
and \U$12909 ( \13041 , \1948 , \5485 );
and \U$12910 ( \13042 , \2090 , \5275 );
nor \U$12911 ( \13043 , \13041 , \13042 );
xnor \U$12912 ( \13044 , \13043 , \5169 );
xor \U$12913 ( \13045 , \13040 , \13044 );
and \U$12914 ( \13046 , \1684 , \5996 );
and \U$12915 ( \13047 , \1802 , \5695 );
nor \U$12916 ( \13048 , \13046 , \13047 );
xnor \U$12917 ( \13049 , \13048 , \5687 );
xor \U$12918 ( \13050 , \13045 , \13049 );
xor \U$12919 ( \13051 , \13036 , \13050 );
xor \U$12920 ( \13052 , \13007 , \13051 );
and \U$12921 ( \13053 , \12778 , \12782 );
and \U$12922 ( \13054 , \12782 , \12784 );
and \U$12923 ( \13055 , \12778 , \12784 );
or \U$12924 ( \13056 , \13053 , \13054 , \13055 );
and \U$12925 ( \13057 , \217 , \9765 );
and \U$12926 ( \13058 , \189 , \9644 );
nor \U$12927 ( \13059 , \13057 , \13058 );
xnor \U$12928 ( \13060 , \13059 , \9478 );
and \U$12929 ( \13061 , \232 , \10408 );
and \U$12930 ( \13062 , \209 , \10116 );
nor \U$12931 ( \13063 , \13061 , \13062 );
xnor \U$12932 ( \13064 , \13063 , \10121 );
xor \U$12933 ( \13065 , \13060 , \13064 );
and \U$12934 ( \13066 , \224 , \10118 );
xor \U$12935 ( \13067 , \13065 , \13066 );
xor \U$12936 ( \13068 , \13056 , \13067 );
and \U$12937 ( \13069 , \307 , \8019 );
and \U$12938 ( \13070 , \412 , \7830 );
nor \U$12939 ( \13071 , \13069 , \13070 );
xnor \U$12940 ( \13072 , \13071 , \7713 );
and \U$12941 ( \13073 , \185 , \8540 );
and \U$12942 ( \13074 , \261 , \8292 );
nor \U$12943 ( \13075 , \13073 , \13074 );
xnor \U$12944 ( \13076 , \13075 , \8297 );
xor \U$12945 ( \13077 , \13072 , \13076 );
and \U$12946 ( \13078 , \197 , \9333 );
and \U$12947 ( \13079 , \178 , \9006 );
nor \U$12948 ( \13080 , \13078 , \13079 );
xnor \U$12949 ( \13081 , \13080 , \8848 );
xor \U$12950 ( \13082 , \13077 , \13081 );
xor \U$12951 ( \13083 , \13068 , \13082 );
xor \U$12952 ( \13084 , \13052 , \13083 );
xor \U$12953 ( \13085 , \12963 , \13084 );
xor \U$12954 ( \13086 , \12914 , \13085 );
xor \U$12955 ( \13087 , \12841 , \13086 );
xor \U$12956 ( \13088 , \12832 , \13087 );
and \U$12957 ( \13089 , \12504 , \12505 );
and \U$12958 ( \13090 , \12505 , \12791 );
and \U$12959 ( \13091 , \12504 , \12791 );
or \U$12960 ( \13092 , \13089 , \13090 , \13091 );
xor \U$12961 ( \13093 , \13088 , \13092 );
and \U$12962 ( \13094 , \12792 , \12796 );
and \U$12963 ( \13095 , \12797 , \12800 );
or \U$12964 ( \13096 , \13094 , \13095 );
xor \U$12965 ( \13097 , \13093 , \13096 );
buf \U$12966 ( \13098 , \13097 );
buf \U$12967 ( \13099 , \13098 );
and \U$12968 ( \13100 , \12811 , \12815 );
and \U$12969 ( \13101 , \12815 , \12830 );
and \U$12970 ( \13102 , \12811 , \12830 );
or \U$12971 ( \13103 , \13100 , \13101 , \13102 );
and \U$12972 ( \13104 , \12836 , \12840 );
and \U$12973 ( \13105 , \12840 , \13086 );
and \U$12974 ( \13106 , \12836 , \13086 );
or \U$12975 ( \13107 , \13104 , \13105 , \13106 );
and \U$12976 ( \13108 , \12820 , \12824 );
and \U$12977 ( \13109 , \12824 , \12829 );
and \U$12978 ( \13110 , \12820 , \12829 );
or \U$12979 ( \13111 , \13108 , \13109 , \13110 );
and \U$12980 ( \13112 , \12855 , \12913 );
and \U$12981 ( \13113 , \12913 , \13085 );
and \U$12982 ( \13114 , \12855 , \13085 );
or \U$12983 ( \13115 , \13112 , \13113 , \13114 );
xor \U$12984 ( \13116 , \13111 , \13115 );
and \U$12985 ( \13117 , \12932 , \12946 );
and \U$12986 ( \13118 , \12946 , \12961 );
and \U$12987 ( \13119 , \12932 , \12961 );
or \U$12988 ( \13120 , \13117 , \13118 , \13119 );
and \U$12989 ( \13121 , \13007 , \13051 );
and \U$12990 ( \13122 , \13051 , \13083 );
and \U$12991 ( \13123 , \13007 , \13083 );
or \U$12992 ( \13124 , \13121 , \13122 , \13123 );
xor \U$12993 ( \13125 , \13120 , \13124 );
and \U$12994 ( \13126 , \13011 , \13015 );
and \U$12995 ( \13127 , \13015 , \13020 );
and \U$12996 ( \13128 , \13011 , \13020 );
or \U$12997 ( \13129 , \13126 , \13127 , \13128 );
and \U$12998 ( \13130 , \12981 , \12985 );
and \U$12999 ( \13131 , \12985 , \12990 );
and \U$13000 ( \13132 , \12981 , \12990 );
or \U$13001 ( \13133 , \13130 , \13131 , \13132 );
xor \U$13002 ( \13134 , \13129 , \13133 );
and \U$13003 ( \13135 , \12996 , \13000 );
and \U$13004 ( \13136 , \13000 , \13005 );
and \U$13005 ( \13137 , \12996 , \13005 );
or \U$13006 ( \13138 , \13135 , \13136 , \13137 );
xor \U$13007 ( \13139 , \13134 , \13138 );
xor \U$13008 ( \13140 , \13125 , \13139 );
xor \U$13009 ( \13141 , \13116 , \13140 );
xor \U$13010 ( \13142 , \13107 , \13141 );
and \U$13011 ( \13143 , \12859 , \12863 );
and \U$13012 ( \13144 , \12863 , \12865 );
and \U$13013 ( \13145 , \12859 , \12865 );
or \U$13014 ( \13146 , \13143 , \13144 , \13145 );
and \U$13015 ( \13147 , \12870 , \12874 );
and \U$13016 ( \13148 , \12874 , \12879 );
and \U$13017 ( \13149 , \12870 , \12879 );
or \U$13018 ( \13150 , \13147 , \13148 , \13149 );
xor \U$13019 ( \13151 , \13146 , \13150 );
and \U$13020 ( \13152 , \12885 , \12899 );
and \U$13021 ( \13153 , \12899 , \12911 );
and \U$13022 ( \13154 , \12885 , \12911 );
or \U$13023 ( \13155 , \13152 , \13153 , \13154 );
xor \U$13024 ( \13156 , \13151 , \13155 );
and \U$13025 ( \13157 , \12845 , \12849 );
and \U$13026 ( \13158 , \12849 , \12854 );
and \U$13027 ( \13159 , \12845 , \12854 );
or \U$13028 ( \13160 , \13157 , \13158 , \13159 );
and \U$13029 ( \13161 , \12866 , \12880 );
and \U$13030 ( \13162 , \12880 , \12912 );
and \U$13031 ( \13163 , \12866 , \12912 );
or \U$13032 ( \13164 , \13161 , \13162 , \13163 );
xor \U$13033 ( \13165 , \13160 , \13164 );
and \U$13034 ( \13166 , \12918 , \12962 );
and \U$13035 ( \13167 , \12962 , \13084 );
and \U$13036 ( \13168 , \12918 , \13084 );
or \U$13037 ( \13169 , \13166 , \13167 , \13168 );
xor \U$13038 ( \13170 , \13165 , \13169 );
xor \U$13039 ( \13171 , \13156 , \13170 );
and \U$13040 ( \13172 , \12922 , \12926 );
and \U$13041 ( \13173 , \12926 , \12931 );
and \U$13042 ( \13174 , \12922 , \12931 );
or \U$13043 ( \13175 , \13172 , \13173 , \13174 );
and \U$13044 ( \13176 , \12936 , \12940 );
and \U$13045 ( \13177 , \12940 , \12945 );
and \U$13046 ( \13178 , \12936 , \12945 );
or \U$13047 ( \13179 , \13176 , \13177 , \13178 );
xor \U$13048 ( \13180 , \13175 , \13179 );
and \U$13049 ( \13181 , \12951 , \12955 );
and \U$13050 ( \13182 , \12955 , \12960 );
and \U$13051 ( \13183 , \12951 , \12960 );
or \U$13052 ( \13184 , \13181 , \13182 , \13183 );
xor \U$13053 ( \13185 , \13180 , \13184 );
and \U$13054 ( \13186 , \12977 , \12991 );
and \U$13055 ( \13187 , \12991 , \13006 );
and \U$13056 ( \13188 , \12977 , \13006 );
or \U$13057 ( \13189 , \13186 , \13187 , \13188 );
and \U$13058 ( \13190 , \13021 , \13035 );
and \U$13059 ( \13191 , \13035 , \13050 );
and \U$13060 ( \13192 , \13021 , \13050 );
or \U$13061 ( \13193 , \13190 , \13191 , \13192 );
xor \U$13062 ( \13194 , \13189 , \13193 );
and \U$13063 ( \13195 , \13056 , \13067 );
and \U$13064 ( \13196 , \13067 , \13082 );
and \U$13065 ( \13197 , \13056 , \13082 );
or \U$13066 ( \13198 , \13195 , \13196 , \13197 );
xor \U$13067 ( \13199 , \13194 , \13198 );
xor \U$13068 ( \13200 , \13185 , \13199 );
and \U$13069 ( \13201 , \12889 , \12893 );
and \U$13070 ( \13202 , \12893 , \12898 );
and \U$13071 ( \13203 , \12889 , \12898 );
or \U$13072 ( \13204 , \13201 , \13202 , \13203 );
and \U$13073 ( \13205 , \12901 , \12905 );
and \U$13074 ( \13206 , \12905 , \12910 );
and \U$13075 ( \13207 , \12901 , \12910 );
or \U$13076 ( \13208 , \13205 , \13206 , \13207 );
xor \U$13077 ( \13209 , \13204 , \13208 );
and \U$13078 ( \13210 , \12967 , \12971 );
and \U$13079 ( \13211 , \12971 , \12976 );
and \U$13080 ( \13212 , \12967 , \12976 );
or \U$13081 ( \13213 , \13210 , \13211 , \13212 );
xor \U$13082 ( \13214 , \13209 , \13213 );
and \U$13083 ( \13215 , \10584 , \245 );
not \U$13084 ( \13216 , \13215 );
xnor \U$13085 ( \13217 , \13216 , \252 );
and \U$13086 ( \13218 , \9897 , \141 );
and \U$13087 ( \13219 , \10206 , \139 );
nor \U$13088 ( \13220 , \13218 , \13219 );
xnor \U$13089 ( \13221 , \13220 , \148 );
xor \U$13090 ( \13222 , \13217 , \13221 );
and \U$13091 ( \13223 , \9169 , \156 );
and \U$13092 ( \13224 , \9465 , \154 );
nor \U$13093 ( \13225 , \13223 , \13224 );
xnor \U$13094 ( \13226 , \13225 , \163 );
xor \U$13095 ( \13227 , \13222 , \13226 );
and \U$13096 ( \13228 , \8652 , \296 );
and \U$13097 ( \13229 , \8835 , \168 );
nor \U$13098 ( \13230 , \13228 , \13229 );
xnor \U$13099 ( \13231 , \13230 , \173 );
and \U$13100 ( \13232 , \8057 , \438 );
and \U$13101 ( \13233 , \8349 , \336 );
nor \U$13102 ( \13234 , \13232 , \13233 );
xnor \U$13103 ( \13235 , \13234 , \320 );
xor \U$13104 ( \13236 , \13231 , \13235 );
and \U$13105 ( \13237 , \7556 , \1086 );
and \U$13106 ( \13238 , \7700 , \508 );
nor \U$13107 ( \13239 , \13237 , \13238 );
xnor \U$13108 ( \13240 , \13239 , \487 );
xor \U$13109 ( \13241 , \13236 , \13240 );
xor \U$13110 ( \13242 , \13227 , \13241 );
and \U$13111 ( \13243 , \4160 , \3103 );
and \U$13112 ( \13244 , \4364 , \2934 );
nor \U$13113 ( \13245 , \13243 , \13244 );
xnor \U$13114 ( \13246 , \13245 , \2839 );
and \U$13115 ( \13247 , \3736 , \3357 );
and \U$13116 ( \13248 , \3912 , \3255 );
nor \U$13117 ( \13249 , \13247 , \13248 );
xnor \U$13118 ( \13250 , \13249 , \3156 );
xor \U$13119 ( \13251 , \13246 , \13250 );
and \U$13120 ( \13252 , \3395 , \3813 );
and \U$13121 ( \13253 , \3646 , \3557 );
nor \U$13122 ( \13254 , \13252 , \13253 );
xnor \U$13123 ( \13255 , \13254 , \3562 );
xor \U$13124 ( \13256 , \13251 , \13255 );
and \U$13125 ( \13257 , \6945 , \1301 );
and \U$13126 ( \13258 , \7231 , \1246 );
nor \U$13127 ( \13259 , \13257 , \13258 );
xnor \U$13128 ( \13260 , \13259 , \1205 );
and \U$13129 ( \13261 , \6514 , \1578 );
and \U$13130 ( \13262 , \6790 , \1431 );
nor \U$13131 ( \13263 , \13261 , \13262 );
xnor \U$13132 ( \13264 , \13263 , \1436 );
xor \U$13133 ( \13265 , \13260 , \13264 );
and \U$13134 ( \13266 , \6030 , \1824 );
and \U$13135 ( \13267 , \6281 , \1739 );
nor \U$13136 ( \13268 , \13266 , \13267 );
xnor \U$13137 ( \13269 , \13268 , \1697 );
xor \U$13138 ( \13270 , \13265 , \13269 );
xor \U$13139 ( \13271 , \13256 , \13270 );
and \U$13140 ( \13272 , \5469 , \2121 );
and \U$13141 ( \13273 , \5674 , \2008 );
nor \U$13142 ( \13274 , \13272 , \13273 );
xnor \U$13143 ( \13275 , \13274 , \1961 );
and \U$13144 ( \13276 , \4922 , \2400 );
and \U$13145 ( \13277 , \5156 , \2246 );
nor \U$13146 ( \13278 , \13276 , \13277 );
xnor \U$13147 ( \13279 , \13278 , \2195 );
xor \U$13148 ( \13280 , \13275 , \13279 );
and \U$13149 ( \13281 , \4654 , \2669 );
and \U$13150 ( \13282 , \4749 , \2538 );
nor \U$13151 ( \13283 , \13281 , \13282 );
xnor \U$13152 ( \13284 , \13283 , \2534 );
xor \U$13153 ( \13285 , \13280 , \13284 );
xor \U$13154 ( \13286 , \13271 , \13285 );
xor \U$13155 ( \13287 , \13242 , \13286 );
xor \U$13156 ( \13288 , \13214 , \13287 );
and \U$13157 ( \13289 , \13025 , \13029 );
and \U$13158 ( \13290 , \13029 , \13034 );
and \U$13159 ( \13291 , \13025 , \13034 );
or \U$13160 ( \13292 , \13289 , \13290 , \13291 );
and \U$13161 ( \13293 , \13040 , \13044 );
and \U$13162 ( \13294 , \13044 , \13049 );
and \U$13163 ( \13295 , \13040 , \13049 );
or \U$13164 ( \13296 , \13293 , \13294 , \13295 );
xor \U$13165 ( \13297 , \13292 , \13296 );
and \U$13166 ( \13298 , \13072 , \13076 );
and \U$13167 ( \13299 , \13076 , \13081 );
and \U$13168 ( \13300 , \13072 , \13081 );
or \U$13169 ( \13301 , \13298 , \13299 , \13300 );
xor \U$13170 ( \13302 , \13297 , \13301 );
and \U$13171 ( \13303 , \3037 , \4132 );
and \U$13172 ( \13304 , \3143 , \4012 );
nor \U$13173 ( \13305 , \13303 , \13304 );
xnor \U$13174 ( \13306 , \13305 , \3925 );
and \U$13175 ( \13307 , \2757 , \4581 );
and \U$13176 ( \13308 , \2826 , \4424 );
nor \U$13177 ( \13309 , \13307 , \13308 );
xnor \U$13178 ( \13310 , \13309 , \4377 );
xor \U$13179 ( \13311 , \13306 , \13310 );
and \U$13180 ( \13312 , \2366 , \5011 );
and \U$13181 ( \13313 , \2521 , \4878 );
nor \U$13182 ( \13314 , \13312 , \13313 );
xnor \U$13183 ( \13315 , \13314 , \4762 );
xor \U$13184 ( \13316 , \13311 , \13315 );
and \U$13185 ( \13317 , \1333 , \7055 );
and \U$13186 ( \13318 , \1484 , \6675 );
nor \U$13187 ( \13319 , \13317 , \13318 );
xnor \U$13188 ( \13320 , \13319 , \6680 );
and \U$13189 ( \13321 , \1147 , \7489 );
and \U$13190 ( \13322 , \1192 , \7137 );
nor \U$13191 ( \13323 , \13321 , \13322 );
xnor \U$13192 ( \13324 , \13323 , \7142 );
xor \U$13193 ( \13325 , \13320 , \13324 );
and \U$13194 ( \13326 , \412 , \8019 );
and \U$13195 ( \13327 , \474 , \7830 );
nor \U$13196 ( \13328 , \13326 , \13327 );
xnor \U$13197 ( \13329 , \13328 , \7713 );
xor \U$13198 ( \13330 , \13325 , \13329 );
xor \U$13199 ( \13331 , \13316 , \13330 );
and \U$13200 ( \13332 , \2090 , \5485 );
and \U$13201 ( \13333 , \2182 , \5275 );
nor \U$13202 ( \13334 , \13332 , \13333 );
xnor \U$13203 ( \13335 , \13334 , \5169 );
and \U$13204 ( \13336 , \1802 , \5996 );
and \U$13205 ( \13337 , \1948 , \5695 );
nor \U$13206 ( \13338 , \13336 , \13337 );
xnor \U$13207 ( \13339 , \13338 , \5687 );
xor \U$13208 ( \13340 , \13335 , \13339 );
and \U$13209 ( \13341 , \1601 , \6401 );
and \U$13210 ( \13342 , \1684 , \6143 );
nor \U$13211 ( \13343 , \13341 , \13342 );
xnor \U$13212 ( \13344 , \13343 , \6148 );
xor \U$13213 ( \13345 , \13340 , \13344 );
xor \U$13214 ( \13346 , \13331 , \13345 );
xor \U$13215 ( \13347 , \13302 , \13346 );
and \U$13216 ( \13348 , \13060 , \13064 );
and \U$13217 ( \13349 , \13064 , \13066 );
and \U$13218 ( \13350 , \13060 , \13066 );
or \U$13219 ( \13351 , \13348 , \13349 , \13350 );
and \U$13220 ( \13352 , \261 , \8540 );
and \U$13221 ( \13353 , \307 , \8292 );
nor \U$13222 ( \13354 , \13352 , \13353 );
xnor \U$13223 ( \13355 , \13354 , \8297 );
and \U$13224 ( \13356 , \178 , \9333 );
and \U$13225 ( \13357 , \185 , \9006 );
nor \U$13226 ( \13358 , \13356 , \13357 );
xnor \U$13227 ( \13359 , \13358 , \8848 );
xor \U$13228 ( \13360 , \13355 , \13359 );
and \U$13229 ( \13361 , \189 , \9765 );
and \U$13230 ( \13362 , \197 , \9644 );
nor \U$13231 ( \13363 , \13361 , \13362 );
xnor \U$13232 ( \13364 , \13363 , \9478 );
xor \U$13233 ( \13365 , \13360 , \13364 );
xor \U$13234 ( \13366 , \13351 , \13365 );
and \U$13235 ( \13367 , \209 , \10408 );
and \U$13236 ( \13368 , \217 , \10116 );
nor \U$13237 ( \13369 , \13367 , \13368 );
xnor \U$13238 ( \13370 , \13369 , \10121 );
and \U$13239 ( \13371 , \232 , \10118 );
xnor \U$13240 ( \13372 , \13370 , \13371 );
xor \U$13241 ( \13373 , \13366 , \13372 );
xor \U$13242 ( \13374 , \13347 , \13373 );
xor \U$13243 ( \13375 , \13288 , \13374 );
xor \U$13244 ( \13376 , \13200 , \13375 );
xor \U$13245 ( \13377 , \13171 , \13376 );
xor \U$13246 ( \13378 , \13142 , \13377 );
xor \U$13247 ( \13379 , \13103 , \13378 );
and \U$13248 ( \13380 , \12807 , \12831 );
and \U$13249 ( \13381 , \12831 , \13087 );
and \U$13250 ( \13382 , \12807 , \13087 );
or \U$13251 ( \13383 , \13380 , \13381 , \13382 );
xor \U$13252 ( \13384 , \13379 , \13383 );
and \U$13253 ( \13385 , \13088 , \13092 );
and \U$13254 ( \13386 , \13093 , \13096 );
or \U$13255 ( \13387 , \13385 , \13386 );
xor \U$13256 ( \13388 , \13384 , \13387 );
buf \U$13257 ( \13389 , \13388 );
buf \U$13258 ( \13390 , \13389 );
and \U$13259 ( \13391 , \13107 , \13141 );
and \U$13260 ( \13392 , \13141 , \13377 );
and \U$13261 ( \13393 , \13107 , \13377 );
or \U$13262 ( \13394 , \13391 , \13392 , \13393 );
and \U$13263 ( \13395 , \13111 , \13115 );
and \U$13264 ( \13396 , \13115 , \13140 );
and \U$13265 ( \13397 , \13111 , \13140 );
or \U$13266 ( \13398 , \13395 , \13396 , \13397 );
and \U$13267 ( \13399 , \13156 , \13170 );
and \U$13268 ( \13400 , \13170 , \13376 );
and \U$13269 ( \13401 , \13156 , \13376 );
or \U$13270 ( \13402 , \13399 , \13400 , \13401 );
xor \U$13271 ( \13403 , \13398 , \13402 );
and \U$13272 ( \13404 , \13146 , \13150 );
and \U$13273 ( \13405 , \13150 , \13155 );
and \U$13274 ( \13406 , \13146 , \13155 );
or \U$13275 ( \13407 , \13404 , \13405 , \13406 );
and \U$13276 ( \13408 , \13120 , \13124 );
and \U$13277 ( \13409 , \13124 , \13139 );
and \U$13278 ( \13410 , \13120 , \13139 );
or \U$13279 ( \13411 , \13408 , \13409 , \13410 );
xor \U$13280 ( \13412 , \13407 , \13411 );
and \U$13281 ( \13413 , \13214 , \13287 );
and \U$13282 ( \13414 , \13287 , \13374 );
and \U$13283 ( \13415 , \13214 , \13374 );
or \U$13284 ( \13416 , \13413 , \13414 , \13415 );
xor \U$13285 ( \13417 , \13412 , \13416 );
xor \U$13286 ( \13418 , \13403 , \13417 );
xor \U$13287 ( \13419 , \13394 , \13418 );
and \U$13288 ( \13420 , \13160 , \13164 );
and \U$13289 ( \13421 , \13164 , \13169 );
and \U$13290 ( \13422 , \13160 , \13169 );
or \U$13291 ( \13423 , \13420 , \13421 , \13422 );
and \U$13292 ( \13424 , \13185 , \13199 );
and \U$13293 ( \13425 , \13199 , \13375 );
and \U$13294 ( \13426 , \13185 , \13375 );
or \U$13295 ( \13427 , \13424 , \13425 , \13426 );
xor \U$13296 ( \13428 , \13423 , \13427 );
and \U$13297 ( \13429 , \13175 , \13179 );
and \U$13298 ( \13430 , \13179 , \13184 );
and \U$13299 ( \13431 , \13175 , \13184 );
or \U$13300 ( \13432 , \13429 , \13430 , \13431 );
and \U$13301 ( \13433 , \13189 , \13193 );
and \U$13302 ( \13434 , \13193 , \13198 );
and \U$13303 ( \13435 , \13189 , \13198 );
or \U$13304 ( \13436 , \13433 , \13434 , \13435 );
xor \U$13305 ( \13437 , \13432 , \13436 );
and \U$13306 ( \13438 , \13227 , \13241 );
and \U$13307 ( \13439 , \13241 , \13286 );
and \U$13308 ( \13440 , \13227 , \13286 );
or \U$13309 ( \13441 , \13438 , \13439 , \13440 );
xor \U$13310 ( \13442 , \13437 , \13441 );
and \U$13311 ( \13443 , \13302 , \13346 );
and \U$13312 ( \13444 , \13346 , \13373 );
and \U$13313 ( \13445 , \13302 , \13373 );
or \U$13314 ( \13446 , \13443 , \13444 , \13445 );
and \U$13315 ( \13447 , \13260 , \13264 );
and \U$13316 ( \13448 , \13264 , \13269 );
and \U$13317 ( \13449 , \13260 , \13269 );
or \U$13318 ( \13450 , \13447 , \13448 , \13449 );
and \U$13319 ( \13451 , \13217 , \13221 );
and \U$13320 ( \13452 , \13221 , \13226 );
and \U$13321 ( \13453 , \13217 , \13226 );
or \U$13322 ( \13454 , \13451 , \13452 , \13453 );
xor \U$13323 ( \13455 , \13450 , \13454 );
and \U$13324 ( \13456 , \13231 , \13235 );
and \U$13325 ( \13457 , \13235 , \13240 );
and \U$13326 ( \13458 , \13231 , \13240 );
or \U$13327 ( \13459 , \13456 , \13457 , \13458 );
xor \U$13328 ( \13460 , \13455 , \13459 );
xor \U$13329 ( \13461 , \13446 , \13460 );
and \U$13330 ( \13462 , \13246 , \13250 );
and \U$13331 ( \13463 , \13250 , \13255 );
and \U$13332 ( \13464 , \13246 , \13255 );
or \U$13333 ( \13465 , \13462 , \13463 , \13464 );
and \U$13334 ( \13466 , \13306 , \13310 );
and \U$13335 ( \13467 , \13310 , \13315 );
and \U$13336 ( \13468 , \13306 , \13315 );
or \U$13337 ( \13469 , \13466 , \13467 , \13468 );
xor \U$13338 ( \13470 , \13465 , \13469 );
and \U$13339 ( \13471 , \13275 , \13279 );
and \U$13340 ( \13472 , \13279 , \13284 );
and \U$13341 ( \13473 , \13275 , \13284 );
or \U$13342 ( \13474 , \13471 , \13472 , \13473 );
xor \U$13343 ( \13475 , \13470 , \13474 );
and \U$13344 ( \13476 , \13320 , \13324 );
and \U$13345 ( \13477 , \13324 , \13329 );
and \U$13346 ( \13478 , \13320 , \13329 );
or \U$13347 ( \13479 , \13476 , \13477 , \13478 );
and \U$13348 ( \13480 , \13335 , \13339 );
and \U$13349 ( \13481 , \13339 , \13344 );
and \U$13350 ( \13482 , \13335 , \13344 );
or \U$13351 ( \13483 , \13480 , \13481 , \13482 );
xor \U$13352 ( \13484 , \13479 , \13483 );
and \U$13353 ( \13485 , \13355 , \13359 );
and \U$13354 ( \13486 , \13359 , \13364 );
and \U$13355 ( \13487 , \13355 , \13364 );
or \U$13356 ( \13488 , \13485 , \13486 , \13487 );
xor \U$13357 ( \13489 , \13484 , \13488 );
xor \U$13358 ( \13490 , \13475 , \13489 );
or \U$13359 ( \13491 , \13370 , \13371 );
and \U$13360 ( \13492 , \217 , \10408 );
and \U$13361 ( \13493 , \189 , \10116 );
nor \U$13362 ( \13494 , \13492 , \13493 );
xnor \U$13363 ( \13495 , \13494 , \10121 );
xor \U$13364 ( \13496 , \13491 , \13495 );
and \U$13365 ( \13497 , \209 , \10118 );
xor \U$13366 ( \13498 , \13496 , \13497 );
xor \U$13367 ( \13499 , \13490 , \13498 );
xor \U$13368 ( \13500 , \13461 , \13499 );
xor \U$13369 ( \13501 , \13442 , \13500 );
and \U$13370 ( \13502 , \13204 , \13208 );
and \U$13371 ( \13503 , \13208 , \13213 );
and \U$13372 ( \13504 , \13204 , \13213 );
or \U$13373 ( \13505 , \13502 , \13503 , \13504 );
and \U$13374 ( \13506 , \13129 , \13133 );
and \U$13375 ( \13507 , \13133 , \13138 );
and \U$13376 ( \13508 , \13129 , \13138 );
or \U$13377 ( \13509 , \13506 , \13507 , \13508 );
xor \U$13378 ( \13510 , \13505 , \13509 );
and \U$13379 ( \13511 , \13292 , \13296 );
and \U$13380 ( \13512 , \13296 , \13301 );
and \U$13381 ( \13513 , \13292 , \13301 );
or \U$13382 ( \13514 , \13511 , \13512 , \13513 );
xor \U$13383 ( \13515 , \13510 , \13514 );
and \U$13384 ( \13516 , \13256 , \13270 );
and \U$13385 ( \13517 , \13270 , \13285 );
and \U$13386 ( \13518 , \13256 , \13285 );
or \U$13387 ( \13519 , \13516 , \13517 , \13518 );
and \U$13388 ( \13520 , \13316 , \13330 );
and \U$13389 ( \13521 , \13330 , \13345 );
and \U$13390 ( \13522 , \13316 , \13345 );
or \U$13391 ( \13523 , \13520 , \13521 , \13522 );
xor \U$13392 ( \13524 , \13519 , \13523 );
and \U$13393 ( \13525 , \13351 , \13365 );
and \U$13394 ( \13526 , \13365 , \13372 );
and \U$13395 ( \13527 , \13351 , \13372 );
or \U$13396 ( \13528 , \13525 , \13526 , \13527 );
xor \U$13397 ( \13529 , \13524 , \13528 );
xor \U$13398 ( \13530 , \13515 , \13529 );
and \U$13399 ( \13531 , \1484 , \7055 );
and \U$13400 ( \13532 , \1601 , \6675 );
nor \U$13401 ( \13533 , \13531 , \13532 );
xnor \U$13402 ( \13534 , \13533 , \6680 );
and \U$13403 ( \13535 , \1192 , \7489 );
and \U$13404 ( \13536 , \1333 , \7137 );
nor \U$13405 ( \13537 , \13535 , \13536 );
xnor \U$13406 ( \13538 , \13537 , \7142 );
xor \U$13407 ( \13539 , \13534 , \13538 );
and \U$13408 ( \13540 , \474 , \8019 );
and \U$13409 ( \13541 , \1147 , \7830 );
nor \U$13410 ( \13542 , \13540 , \13541 );
xnor \U$13411 ( \13543 , \13542 , \7713 );
xor \U$13412 ( \13544 , \13539 , \13543 );
and \U$13413 ( \13545 , \307 , \8540 );
and \U$13414 ( \13546 , \412 , \8292 );
nor \U$13415 ( \13547 , \13545 , \13546 );
xnor \U$13416 ( \13548 , \13547 , \8297 );
and \U$13417 ( \13549 , \185 , \9333 );
and \U$13418 ( \13550 , \261 , \9006 );
nor \U$13419 ( \13551 , \13549 , \13550 );
xnor \U$13420 ( \13552 , \13551 , \8848 );
xor \U$13421 ( \13553 , \13548 , \13552 );
and \U$13422 ( \13554 , \197 , \9765 );
and \U$13423 ( \13555 , \178 , \9644 );
nor \U$13424 ( \13556 , \13554 , \13555 );
xnor \U$13425 ( \13557 , \13556 , \9478 );
xor \U$13426 ( \13558 , \13553 , \13557 );
xor \U$13427 ( \13559 , \13544 , \13558 );
and \U$13428 ( \13560 , \2182 , \5485 );
and \U$13429 ( \13561 , \2366 , \5275 );
nor \U$13430 ( \13562 , \13560 , \13561 );
xnor \U$13431 ( \13563 , \13562 , \5169 );
and \U$13432 ( \13564 , \1948 , \5996 );
and \U$13433 ( \13565 , \2090 , \5695 );
nor \U$13434 ( \13566 , \13564 , \13565 );
xnor \U$13435 ( \13567 , \13566 , \5687 );
xor \U$13436 ( \13568 , \13563 , \13567 );
and \U$13437 ( \13569 , \1684 , \6401 );
and \U$13438 ( \13570 , \1802 , \6143 );
nor \U$13439 ( \13571 , \13569 , \13570 );
xnor \U$13440 ( \13572 , \13571 , \6148 );
xor \U$13441 ( \13573 , \13568 , \13572 );
xor \U$13442 ( \13574 , \13559 , \13573 );
and \U$13443 ( \13575 , \3143 , \4132 );
and \U$13444 ( \13576 , \3395 , \4012 );
nor \U$13445 ( \13577 , \13575 , \13576 );
xnor \U$13446 ( \13578 , \13577 , \3925 );
and \U$13447 ( \13579 , \2826 , \4581 );
and \U$13448 ( \13580 , \3037 , \4424 );
nor \U$13449 ( \13581 , \13579 , \13580 );
xnor \U$13450 ( \13582 , \13581 , \4377 );
xor \U$13451 ( \13583 , \13578 , \13582 );
and \U$13452 ( \13584 , \2521 , \5011 );
and \U$13453 ( \13585 , \2757 , \4878 );
nor \U$13454 ( \13586 , \13584 , \13585 );
xnor \U$13455 ( \13587 , \13586 , \4762 );
xor \U$13456 ( \13588 , \13583 , \13587 );
and \U$13457 ( \13589 , \5674 , \2121 );
and \U$13458 ( \13590 , \6030 , \2008 );
nor \U$13459 ( \13591 , \13589 , \13590 );
xnor \U$13460 ( \13592 , \13591 , \1961 );
and \U$13461 ( \13593 , \5156 , \2400 );
and \U$13462 ( \13594 , \5469 , \2246 );
nor \U$13463 ( \13595 , \13593 , \13594 );
xnor \U$13464 ( \13596 , \13595 , \2195 );
xor \U$13465 ( \13597 , \13592 , \13596 );
and \U$13466 ( \13598 , \4749 , \2669 );
and \U$13467 ( \13599 , \4922 , \2538 );
nor \U$13468 ( \13600 , \13598 , \13599 );
xnor \U$13469 ( \13601 , \13600 , \2534 );
xor \U$13470 ( \13602 , \13597 , \13601 );
xor \U$13471 ( \13603 , \13588 , \13602 );
and \U$13472 ( \13604 , \4364 , \3103 );
and \U$13473 ( \13605 , \4654 , \2934 );
nor \U$13474 ( \13606 , \13604 , \13605 );
xnor \U$13475 ( \13607 , \13606 , \2839 );
and \U$13476 ( \13608 , \3912 , \3357 );
and \U$13477 ( \13609 , \4160 , \3255 );
nor \U$13478 ( \13610 , \13608 , \13609 );
xnor \U$13479 ( \13611 , \13610 , \3156 );
xor \U$13480 ( \13612 , \13607 , \13611 );
and \U$13481 ( \13613 , \3646 , \3813 );
and \U$13482 ( \13614 , \3736 , \3557 );
nor \U$13483 ( \13615 , \13613 , \13614 );
xnor \U$13484 ( \13616 , \13615 , \3562 );
xor \U$13485 ( \13617 , \13612 , \13616 );
xor \U$13486 ( \13618 , \13603 , \13617 );
xor \U$13487 ( \13619 , \13574 , \13618 );
and \U$13488 ( \13620 , \7231 , \1301 );
and \U$13489 ( \13621 , \7556 , \1246 );
nor \U$13490 ( \13622 , \13620 , \13621 );
xnor \U$13491 ( \13623 , \13622 , \1205 );
and \U$13492 ( \13624 , \6790 , \1578 );
and \U$13493 ( \13625 , \6945 , \1431 );
nor \U$13494 ( \13626 , \13624 , \13625 );
xnor \U$13495 ( \13627 , \13626 , \1436 );
xor \U$13496 ( \13628 , \13623 , \13627 );
and \U$13497 ( \13629 , \6281 , \1824 );
and \U$13498 ( \13630 , \6514 , \1739 );
nor \U$13499 ( \13631 , \13629 , \13630 );
xnor \U$13500 ( \13632 , \13631 , \1697 );
xor \U$13501 ( \13633 , \13628 , \13632 );
not \U$13502 ( \13634 , \252 );
and \U$13503 ( \13635 , \10206 , \141 );
and \U$13504 ( \13636 , \10584 , \139 );
nor \U$13505 ( \13637 , \13635 , \13636 );
xnor \U$13506 ( \13638 , \13637 , \148 );
xor \U$13507 ( \13639 , \13634 , \13638 );
and \U$13508 ( \13640 , \9465 , \156 );
and \U$13509 ( \13641 , \9897 , \154 );
nor \U$13510 ( \13642 , \13640 , \13641 );
xnor \U$13511 ( \13643 , \13642 , \163 );
xor \U$13512 ( \13644 , \13639 , \13643 );
xor \U$13513 ( \13645 , \13633 , \13644 );
and \U$13514 ( \13646 , \8835 , \296 );
and \U$13515 ( \13647 , \9169 , \168 );
nor \U$13516 ( \13648 , \13646 , \13647 );
xnor \U$13517 ( \13649 , \13648 , \173 );
and \U$13518 ( \13650 , \8349 , \438 );
and \U$13519 ( \13651 , \8652 , \336 );
nor \U$13520 ( \13652 , \13650 , \13651 );
xnor \U$13521 ( \13653 , \13652 , \320 );
xor \U$13522 ( \13654 , \13649 , \13653 );
and \U$13523 ( \13655 , \7700 , \1086 );
and \U$13524 ( \13656 , \8057 , \508 );
nor \U$13525 ( \13657 , \13655 , \13656 );
xnor \U$13526 ( \13658 , \13657 , \487 );
xor \U$13527 ( \13659 , \13654 , \13658 );
xor \U$13528 ( \13660 , \13645 , \13659 );
xor \U$13529 ( \13661 , \13619 , \13660 );
xor \U$13530 ( \13662 , \13530 , \13661 );
xor \U$13531 ( \13663 , \13501 , \13662 );
xor \U$13532 ( \13664 , \13428 , \13663 );
xor \U$13533 ( \13665 , \13419 , \13664 );
and \U$13534 ( \13666 , \13103 , \13378 );
xor \U$13535 ( \13667 , \13665 , \13666 );
and \U$13536 ( \13668 , \13379 , \13383 );
and \U$13537 ( \13669 , \13384 , \13387 );
or \U$13538 ( \13670 , \13668 , \13669 );
xor \U$13539 ( \13671 , \13667 , \13670 );
buf \U$13540 ( \13672 , \13671 );
buf \U$13541 ( \13673 , \13672 );
and \U$13542 ( \13674 , \13398 , \13402 );
and \U$13543 ( \13675 , \13402 , \13417 );
and \U$13544 ( \13676 , \13398 , \13417 );
or \U$13545 ( \13677 , \13674 , \13675 , \13676 );
and \U$13546 ( \13678 , \13423 , \13427 );
and \U$13547 ( \13679 , \13427 , \13663 );
and \U$13548 ( \13680 , \13423 , \13663 );
or \U$13549 ( \13681 , \13678 , \13679 , \13680 );
and \U$13550 ( \13682 , \13432 , \13436 );
and \U$13551 ( \13683 , \13436 , \13441 );
and \U$13552 ( \13684 , \13432 , \13441 );
or \U$13553 ( \13685 , \13682 , \13683 , \13684 );
and \U$13554 ( \13686 , \13446 , \13460 );
and \U$13555 ( \13687 , \13460 , \13499 );
and \U$13556 ( \13688 , \13446 , \13499 );
or \U$13557 ( \13689 , \13686 , \13687 , \13688 );
xor \U$13558 ( \13690 , \13685 , \13689 );
and \U$13559 ( \13691 , \13515 , \13529 );
and \U$13560 ( \13692 , \13529 , \13661 );
and \U$13561 ( \13693 , \13515 , \13661 );
or \U$13562 ( \13694 , \13691 , \13692 , \13693 );
xor \U$13563 ( \13695 , \13690 , \13694 );
xor \U$13564 ( \13696 , \13681 , \13695 );
and \U$13565 ( \13697 , \13407 , \13411 );
and \U$13566 ( \13698 , \13411 , \13416 );
and \U$13567 ( \13699 , \13407 , \13416 );
or \U$13568 ( \13700 , \13697 , \13698 , \13699 );
and \U$13569 ( \13701 , \13442 , \13500 );
and \U$13570 ( \13702 , \13500 , \13662 );
and \U$13571 ( \13703 , \13442 , \13662 );
or \U$13572 ( \13704 , \13701 , \13702 , \13703 );
xor \U$13573 ( \13705 , \13700 , \13704 );
and \U$13574 ( \13706 , \13505 , \13509 );
and \U$13575 ( \13707 , \13509 , \13514 );
and \U$13576 ( \13708 , \13505 , \13514 );
or \U$13577 ( \13709 , \13706 , \13707 , \13708 );
and \U$13578 ( \13710 , \13519 , \13523 );
and \U$13579 ( \13711 , \13523 , \13528 );
and \U$13580 ( \13712 , \13519 , \13528 );
or \U$13581 ( \13713 , \13710 , \13711 , \13712 );
xor \U$13582 ( \13714 , \13709 , \13713 );
and \U$13583 ( \13715 , \13574 , \13618 );
and \U$13584 ( \13716 , \13618 , \13660 );
and \U$13585 ( \13717 , \13574 , \13660 );
or \U$13586 ( \13718 , \13715 , \13716 , \13717 );
xor \U$13587 ( \13719 , \13714 , \13718 );
and \U$13588 ( \13720 , \13465 , \13469 );
and \U$13589 ( \13721 , \13469 , \13474 );
and \U$13590 ( \13722 , \13465 , \13474 );
or \U$13591 ( \13723 , \13720 , \13721 , \13722 );
and \U$13592 ( \13724 , \13479 , \13483 );
and \U$13593 ( \13725 , \13483 , \13488 );
and \U$13594 ( \13726 , \13479 , \13488 );
or \U$13595 ( \13727 , \13724 , \13725 , \13726 );
xor \U$13596 ( \13728 , \13723 , \13727 );
and \U$13597 ( \13729 , \13450 , \13454 );
and \U$13598 ( \13730 , \13454 , \13459 );
and \U$13599 ( \13731 , \13450 , \13459 );
or \U$13600 ( \13732 , \13729 , \13730 , \13731 );
xor \U$13601 ( \13733 , \13728 , \13732 );
and \U$13602 ( \13734 , \13491 , \13495 );
and \U$13603 ( \13735 , \13495 , \13497 );
and \U$13604 ( \13736 , \13491 , \13497 );
or \U$13605 ( \13737 , \13734 , \13735 , \13736 );
and \U$13606 ( \13738 , \13544 , \13558 );
and \U$13607 ( \13739 , \13558 , \13573 );
and \U$13608 ( \13740 , \13544 , \13573 );
or \U$13609 ( \13741 , \13738 , \13739 , \13740 );
xor \U$13610 ( \13742 , \13737 , \13741 );
and \U$13611 ( \13743 , \13588 , \13602 );
and \U$13612 ( \13744 , \13602 , \13617 );
and \U$13613 ( \13745 , \13588 , \13617 );
or \U$13614 ( \13746 , \13743 , \13744 , \13745 );
xor \U$13615 ( \13747 , \13742 , \13746 );
xor \U$13616 ( \13748 , \13733 , \13747 );
and \U$13617 ( \13749 , \13633 , \13644 );
and \U$13618 ( \13750 , \13644 , \13659 );
and \U$13619 ( \13751 , \13633 , \13659 );
or \U$13620 ( \13752 , \13749 , \13750 , \13751 );
and \U$13621 ( \13753 , \8652 , \438 );
and \U$13622 ( \13754 , \8835 , \336 );
nor \U$13623 ( \13755 , \13753 , \13754 );
xnor \U$13624 ( \13756 , \13755 , \320 );
and \U$13625 ( \13757 , \8057 , \1086 );
and \U$13626 ( \13758 , \8349 , \508 );
nor \U$13627 ( \13759 , \13757 , \13758 );
xnor \U$13628 ( \13760 , \13759 , \487 );
xor \U$13629 ( \13761 , \13756 , \13760 );
and \U$13630 ( \13762 , \7556 , \1301 );
and \U$13631 ( \13763 , \7700 , \1246 );
nor \U$13632 ( \13764 , \13762 , \13763 );
xnor \U$13633 ( \13765 , \13764 , \1205 );
xor \U$13634 ( \13766 , \13761 , \13765 );
xor \U$13635 ( \13767 , \13752 , \13766 );
and \U$13636 ( \13768 , \10584 , \141 );
not \U$13637 ( \13769 , \13768 );
xnor \U$13638 ( \13770 , \13769 , \148 );
and \U$13639 ( \13771 , \9897 , \156 );
and \U$13640 ( \13772 , \10206 , \154 );
nor \U$13641 ( \13773 , \13771 , \13772 );
xnor \U$13642 ( \13774 , \13773 , \163 );
xor \U$13643 ( \13775 , \13770 , \13774 );
and \U$13644 ( \13776 , \9169 , \296 );
and \U$13645 ( \13777 , \9465 , \168 );
nor \U$13646 ( \13778 , \13776 , \13777 );
xnor \U$13647 ( \13779 , \13778 , \173 );
xor \U$13648 ( \13780 , \13775 , \13779 );
xor \U$13649 ( \13781 , \13767 , \13780 );
xor \U$13650 ( \13782 , \13748 , \13781 );
xor \U$13651 ( \13783 , \13719 , \13782 );
and \U$13652 ( \13784 , \13475 , \13489 );
and \U$13653 ( \13785 , \13489 , \13498 );
and \U$13654 ( \13786 , \13475 , \13498 );
or \U$13655 ( \13787 , \13784 , \13785 , \13786 );
and \U$13656 ( \13788 , \13578 , \13582 );
and \U$13657 ( \13789 , \13582 , \13587 );
and \U$13658 ( \13790 , \13578 , \13587 );
or \U$13659 ( \13791 , \13788 , \13789 , \13790 );
and \U$13660 ( \13792 , \13592 , \13596 );
and \U$13661 ( \13793 , \13596 , \13601 );
and \U$13662 ( \13794 , \13592 , \13601 );
or \U$13663 ( \13795 , \13792 , \13793 , \13794 );
xor \U$13664 ( \13796 , \13791 , \13795 );
and \U$13665 ( \13797 , \13607 , \13611 );
and \U$13666 ( \13798 , \13611 , \13616 );
and \U$13667 ( \13799 , \13607 , \13616 );
or \U$13668 ( \13800 , \13797 , \13798 , \13799 );
xor \U$13669 ( \13801 , \13796 , \13800 );
and \U$13670 ( \13802 , \13623 , \13627 );
and \U$13671 ( \13803 , \13627 , \13632 );
and \U$13672 ( \13804 , \13623 , \13632 );
or \U$13673 ( \13805 , \13802 , \13803 , \13804 );
and \U$13674 ( \13806 , \13634 , \13638 );
and \U$13675 ( \13807 , \13638 , \13643 );
and \U$13676 ( \13808 , \13634 , \13643 );
or \U$13677 ( \13809 , \13806 , \13807 , \13808 );
xor \U$13678 ( \13810 , \13805 , \13809 );
and \U$13679 ( \13811 , \13649 , \13653 );
and \U$13680 ( \13812 , \13653 , \13658 );
and \U$13681 ( \13813 , \13649 , \13658 );
or \U$13682 ( \13814 , \13811 , \13812 , \13813 );
xor \U$13683 ( \13815 , \13810 , \13814 );
xor \U$13684 ( \13816 , \13801 , \13815 );
and \U$13685 ( \13817 , \13534 , \13538 );
and \U$13686 ( \13818 , \13538 , \13543 );
and \U$13687 ( \13819 , \13534 , \13543 );
or \U$13688 ( \13820 , \13817 , \13818 , \13819 );
and \U$13689 ( \13821 , \13548 , \13552 );
and \U$13690 ( \13822 , \13552 , \13557 );
and \U$13691 ( \13823 , \13548 , \13557 );
or \U$13692 ( \13824 , \13821 , \13822 , \13823 );
xor \U$13693 ( \13825 , \13820 , \13824 );
and \U$13694 ( \13826 , \13563 , \13567 );
and \U$13695 ( \13827 , \13567 , \13572 );
and \U$13696 ( \13828 , \13563 , \13572 );
or \U$13697 ( \13829 , \13826 , \13827 , \13828 );
xor \U$13698 ( \13830 , \13825 , \13829 );
xor \U$13699 ( \13831 , \13816 , \13830 );
xor \U$13700 ( \13832 , \13787 , \13831 );
and \U$13701 ( \13833 , \2090 , \5996 );
and \U$13702 ( \13834 , \2182 , \5695 );
nor \U$13703 ( \13835 , \13833 , \13834 );
xnor \U$13704 ( \13836 , \13835 , \5687 );
and \U$13705 ( \13837 , \1802 , \6401 );
and \U$13706 ( \13838 , \1948 , \6143 );
nor \U$13707 ( \13839 , \13837 , \13838 );
xnor \U$13708 ( \13840 , \13839 , \6148 );
xor \U$13709 ( \13841 , \13836 , \13840 );
and \U$13710 ( \13842 , \1601 , \7055 );
and \U$13711 ( \13843 , \1684 , \6675 );
nor \U$13712 ( \13844 , \13842 , \13843 );
xnor \U$13713 ( \13845 , \13844 , \6680 );
xor \U$13714 ( \13846 , \13841 , \13845 );
and \U$13715 ( \13847 , \3037 , \4581 );
and \U$13716 ( \13848 , \3143 , \4424 );
nor \U$13717 ( \13849 , \13847 , \13848 );
xnor \U$13718 ( \13850 , \13849 , \4377 );
and \U$13719 ( \13851 , \2757 , \5011 );
and \U$13720 ( \13852 , \2826 , \4878 );
nor \U$13721 ( \13853 , \13851 , \13852 );
xnor \U$13722 ( \13854 , \13853 , \4762 );
xor \U$13723 ( \13855 , \13850 , \13854 );
and \U$13724 ( \13856 , \2366 , \5485 );
and \U$13725 ( \13857 , \2521 , \5275 );
nor \U$13726 ( \13858 , \13856 , \13857 );
xnor \U$13727 ( \13859 , \13858 , \5169 );
xor \U$13728 ( \13860 , \13855 , \13859 );
xor \U$13729 ( \13861 , \13846 , \13860 );
and \U$13730 ( \13862 , \1333 , \7489 );
and \U$13731 ( \13863 , \1484 , \7137 );
nor \U$13732 ( \13864 , \13862 , \13863 );
xnor \U$13733 ( \13865 , \13864 , \7142 );
and \U$13734 ( \13866 , \1147 , \8019 );
and \U$13735 ( \13867 , \1192 , \7830 );
nor \U$13736 ( \13868 , \13866 , \13867 );
xnor \U$13737 ( \13869 , \13868 , \7713 );
xor \U$13738 ( \13870 , \13865 , \13869 );
and \U$13739 ( \13871 , \412 , \8540 );
and \U$13740 ( \13872 , \474 , \8292 );
nor \U$13741 ( \13873 , \13871 , \13872 );
xnor \U$13742 ( \13874 , \13873 , \8297 );
xor \U$13743 ( \13875 , \13870 , \13874 );
xor \U$13744 ( \13876 , \13861 , \13875 );
and \U$13745 ( \13877 , \6945 , \1578 );
and \U$13746 ( \13878 , \7231 , \1431 );
nor \U$13747 ( \13879 , \13877 , \13878 );
xnor \U$13748 ( \13880 , \13879 , \1436 );
and \U$13749 ( \13881 , \6514 , \1824 );
and \U$13750 ( \13882 , \6790 , \1739 );
nor \U$13751 ( \13883 , \13881 , \13882 );
xnor \U$13752 ( \13884 , \13883 , \1697 );
xor \U$13753 ( \13885 , \13880 , \13884 );
and \U$13754 ( \13886 , \6030 , \2121 );
and \U$13755 ( \13887 , \6281 , \2008 );
nor \U$13756 ( \13888 , \13886 , \13887 );
xnor \U$13757 ( \13889 , \13888 , \1961 );
xor \U$13758 ( \13890 , \13885 , \13889 );
and \U$13759 ( \13891 , \5469 , \2400 );
and \U$13760 ( \13892 , \5674 , \2246 );
nor \U$13761 ( \13893 , \13891 , \13892 );
xnor \U$13762 ( \13894 , \13893 , \2195 );
and \U$13763 ( \13895 , \4922 , \2669 );
and \U$13764 ( \13896 , \5156 , \2538 );
nor \U$13765 ( \13897 , \13895 , \13896 );
xnor \U$13766 ( \13898 , \13897 , \2534 );
xor \U$13767 ( \13899 , \13894 , \13898 );
and \U$13768 ( \13900 , \4654 , \3103 );
and \U$13769 ( \13901 , \4749 , \2934 );
nor \U$13770 ( \13902 , \13900 , \13901 );
xnor \U$13771 ( \13903 , \13902 , \2839 );
xor \U$13772 ( \13904 , \13899 , \13903 );
xor \U$13773 ( \13905 , \13890 , \13904 );
and \U$13774 ( \13906 , \4160 , \3357 );
and \U$13775 ( \13907 , \4364 , \3255 );
nor \U$13776 ( \13908 , \13906 , \13907 );
xnor \U$13777 ( \13909 , \13908 , \3156 );
and \U$13778 ( \13910 , \3736 , \3813 );
and \U$13779 ( \13911 , \3912 , \3557 );
nor \U$13780 ( \13912 , \13910 , \13911 );
xnor \U$13781 ( \13913 , \13912 , \3562 );
xor \U$13782 ( \13914 , \13909 , \13913 );
and \U$13783 ( \13915 , \3395 , \4132 );
and \U$13784 ( \13916 , \3646 , \4012 );
nor \U$13785 ( \13917 , \13915 , \13916 );
xnor \U$13786 ( \13918 , \13917 , \3925 );
xor \U$13787 ( \13919 , \13914 , \13918 );
xor \U$13788 ( \13920 , \13905 , \13919 );
xor \U$13789 ( \13921 , \13876 , \13920 );
and \U$13790 ( \13922 , \217 , \10118 );
and \U$13791 ( \13923 , \261 , \9333 );
and \U$13792 ( \13924 , \307 , \9006 );
nor \U$13793 ( \13925 , \13923 , \13924 );
xnor \U$13794 ( \13926 , \13925 , \8848 );
and \U$13795 ( \13927 , \178 , \9765 );
and \U$13796 ( \13928 , \185 , \9644 );
nor \U$13797 ( \13929 , \13927 , \13928 );
xnor \U$13798 ( \13930 , \13929 , \9478 );
xor \U$13799 ( \13931 , \13926 , \13930 );
and \U$13800 ( \13932 , \189 , \10408 );
and \U$13801 ( \13933 , \197 , \10116 );
nor \U$13802 ( \13934 , \13932 , \13933 );
xnor \U$13803 ( \13935 , \13934 , \10121 );
xor \U$13804 ( \13936 , \13931 , \13935 );
xnor \U$13805 ( \13937 , \13922 , \13936 );
xor \U$13806 ( \13938 , \13921 , \13937 );
xor \U$13807 ( \13939 , \13832 , \13938 );
xor \U$13808 ( \13940 , \13783 , \13939 );
xor \U$13809 ( \13941 , \13705 , \13940 );
xor \U$13810 ( \13942 , \13696 , \13941 );
xor \U$13811 ( \13943 , \13677 , \13942 );
and \U$13812 ( \13944 , \13394 , \13418 );
and \U$13813 ( \13945 , \13418 , \13664 );
and \U$13814 ( \13946 , \13394 , \13664 );
or \U$13815 ( \13947 , \13944 , \13945 , \13946 );
xor \U$13816 ( \13948 , \13943 , \13947 );
and \U$13817 ( \13949 , \13665 , \13666 );
and \U$13818 ( \13950 , \13667 , \13670 );
or \U$13819 ( \13951 , \13949 , \13950 );
xor \U$13820 ( \13952 , \13948 , \13951 );
buf \U$13821 ( \13953 , \13952 );
buf \U$13822 ( \13954 , \13953 );
and \U$13823 ( \13955 , \13681 , \13695 );
and \U$13824 ( \13956 , \13695 , \13941 );
and \U$13825 ( \13957 , \13681 , \13941 );
or \U$13826 ( \13958 , \13955 , \13956 , \13957 );
and \U$13827 ( \13959 , \13700 , \13704 );
and \U$13828 ( \13960 , \13704 , \13940 );
and \U$13829 ( \13961 , \13700 , \13940 );
or \U$13830 ( \13962 , \13959 , \13960 , \13961 );
and \U$13831 ( \13963 , \13685 , \13689 );
and \U$13832 ( \13964 , \13689 , \13694 );
and \U$13833 ( \13965 , \13685 , \13694 );
or \U$13834 ( \13966 , \13963 , \13964 , \13965 );
and \U$13835 ( \13967 , \13719 , \13782 );
and \U$13836 ( \13968 , \13782 , \13939 );
and \U$13837 ( \13969 , \13719 , \13939 );
or \U$13838 ( \13970 , \13967 , \13968 , \13969 );
xor \U$13839 ( \13971 , \13966 , \13970 );
and \U$13840 ( \13972 , \13723 , \13727 );
and \U$13841 ( \13973 , \13727 , \13732 );
and \U$13842 ( \13974 , \13723 , \13732 );
or \U$13843 ( \13975 , \13972 , \13973 , \13974 );
and \U$13844 ( \13976 , \13737 , \13741 );
and \U$13845 ( \13977 , \13741 , \13746 );
and \U$13846 ( \13978 , \13737 , \13746 );
or \U$13847 ( \13979 , \13976 , \13977 , \13978 );
xor \U$13848 ( \13980 , \13975 , \13979 );
and \U$13849 ( \13981 , \13752 , \13766 );
and \U$13850 ( \13982 , \13766 , \13780 );
and \U$13851 ( \13983 , \13752 , \13780 );
or \U$13852 ( \13984 , \13981 , \13982 , \13983 );
xor \U$13853 ( \13985 , \13980 , \13984 );
xor \U$13854 ( \13986 , \13971 , \13985 );
xor \U$13855 ( \13987 , \13962 , \13986 );
and \U$13856 ( \13988 , \13709 , \13713 );
and \U$13857 ( \13989 , \13713 , \13718 );
and \U$13858 ( \13990 , \13709 , \13718 );
or \U$13859 ( \13991 , \13988 , \13989 , \13990 );
and \U$13860 ( \13992 , \13733 , \13747 );
and \U$13861 ( \13993 , \13747 , \13781 );
and \U$13862 ( \13994 , \13733 , \13781 );
or \U$13863 ( \13995 , \13992 , \13993 , \13994 );
xor \U$13864 ( \13996 , \13991 , \13995 );
and \U$13865 ( \13997 , \13787 , \13831 );
and \U$13866 ( \13998 , \13831 , \13938 );
and \U$13867 ( \13999 , \13787 , \13938 );
or \U$13868 ( \14000 , \13997 , \13998 , \13999 );
xor \U$13869 ( \14001 , \13996 , \14000 );
and \U$13870 ( \14002 , \13791 , \13795 );
and \U$13871 ( \14003 , \13795 , \13800 );
and \U$13872 ( \14004 , \13791 , \13800 );
or \U$13873 ( \14005 , \14002 , \14003 , \14004 );
and \U$13874 ( \14006 , \13805 , \13809 );
and \U$13875 ( \14007 , \13809 , \13814 );
and \U$13876 ( \14008 , \13805 , \13814 );
or \U$13877 ( \14009 , \14006 , \14007 , \14008 );
xor \U$13878 ( \14010 , \14005 , \14009 );
and \U$13879 ( \14011 , \13820 , \13824 );
and \U$13880 ( \14012 , \13824 , \13829 );
and \U$13881 ( \14013 , \13820 , \13829 );
or \U$13882 ( \14014 , \14011 , \14012 , \14013 );
xor \U$13883 ( \14015 , \14010 , \14014 );
and \U$13884 ( \14016 , \13801 , \13815 );
and \U$13885 ( \14017 , \13815 , \13830 );
and \U$13886 ( \14018 , \13801 , \13830 );
or \U$13887 ( \14019 , \14016 , \14017 , \14018 );
and \U$13888 ( \14020 , \13876 , \13920 );
and \U$13889 ( \14021 , \13920 , \13937 );
and \U$13890 ( \14022 , \13876 , \13937 );
or \U$13891 ( \14023 , \14020 , \14021 , \14022 );
xor \U$13892 ( \14024 , \14019 , \14023 );
and \U$13893 ( \14025 , \13756 , \13760 );
and \U$13894 ( \14026 , \13760 , \13765 );
and \U$13895 ( \14027 , \13756 , \13765 );
or \U$13896 ( \14028 , \14025 , \14026 , \14027 );
and \U$13897 ( \14029 , \13880 , \13884 );
and \U$13898 ( \14030 , \13884 , \13889 );
and \U$13899 ( \14031 , \13880 , \13889 );
or \U$13900 ( \14032 , \14029 , \14030 , \14031 );
xor \U$13901 ( \14033 , \14028 , \14032 );
and \U$13902 ( \14034 , \13770 , \13774 );
and \U$13903 ( \14035 , \13774 , \13779 );
and \U$13904 ( \14036 , \13770 , \13779 );
or \U$13905 ( \14037 , \14034 , \14035 , \14036 );
xor \U$13906 ( \14038 , \14033 , \14037 );
xor \U$13907 ( \14039 , \14024 , \14038 );
xor \U$13908 ( \14040 , \14015 , \14039 );
and \U$13909 ( \14041 , \13846 , \13860 );
and \U$13910 ( \14042 , \13860 , \13875 );
and \U$13911 ( \14043 , \13846 , \13875 );
or \U$13912 ( \14044 , \14041 , \14042 , \14043 );
and \U$13913 ( \14045 , \13890 , \13904 );
and \U$13914 ( \14046 , \13904 , \13919 );
and \U$13915 ( \14047 , \13890 , \13919 );
or \U$13916 ( \14048 , \14045 , \14046 , \14047 );
xor \U$13917 ( \14049 , \14044 , \14048 );
or \U$13918 ( \14050 , \13922 , \13936 );
xor \U$13919 ( \14051 , \14049 , \14050 );
and \U$13920 ( \14052 , \13836 , \13840 );
and \U$13921 ( \14053 , \13840 , \13845 );
and \U$13922 ( \14054 , \13836 , \13845 );
or \U$13923 ( \14055 , \14052 , \14053 , \14054 );
and \U$13924 ( \14056 , \13926 , \13930 );
and \U$13925 ( \14057 , \13930 , \13935 );
and \U$13926 ( \14058 , \13926 , \13935 );
or \U$13927 ( \14059 , \14056 , \14057 , \14058 );
xor \U$13928 ( \14060 , \14055 , \14059 );
and \U$13929 ( \14061 , \13865 , \13869 );
and \U$13930 ( \14062 , \13869 , \13874 );
and \U$13931 ( \14063 , \13865 , \13874 );
or \U$13932 ( \14064 , \14061 , \14062 , \14063 );
xor \U$13933 ( \14065 , \14060 , \14064 );
and \U$13934 ( \14066 , \13850 , \13854 );
and \U$13935 ( \14067 , \13854 , \13859 );
and \U$13936 ( \14068 , \13850 , \13859 );
or \U$13937 ( \14069 , \14066 , \14067 , \14068 );
and \U$13938 ( \14070 , \13894 , \13898 );
and \U$13939 ( \14071 , \13898 , \13903 );
and \U$13940 ( \14072 , \13894 , \13903 );
or \U$13941 ( \14073 , \14070 , \14071 , \14072 );
xor \U$13942 ( \14074 , \14069 , \14073 );
and \U$13943 ( \14075 , \13909 , \13913 );
and \U$13944 ( \14076 , \13913 , \13918 );
and \U$13945 ( \14077 , \13909 , \13918 );
or \U$13946 ( \14078 , \14075 , \14076 , \14077 );
xor \U$13947 ( \14079 , \14074 , \14078 );
xor \U$13948 ( \14080 , \14065 , \14079 );
and \U$13949 ( \14081 , \189 , \10118 );
and \U$13950 ( \14082 , \1484 , \7489 );
and \U$13951 ( \14083 , \1601 , \7137 );
nor \U$13952 ( \14084 , \14082 , \14083 );
xnor \U$13953 ( \14085 , \14084 , \7142 );
and \U$13954 ( \14086 , \1192 , \8019 );
and \U$13955 ( \14087 , \1333 , \7830 );
nor \U$13956 ( \14088 , \14086 , \14087 );
xnor \U$13957 ( \14089 , \14088 , \7713 );
xor \U$13958 ( \14090 , \14085 , \14089 );
and \U$13959 ( \14091 , \474 , \8540 );
and \U$13960 ( \14092 , \1147 , \8292 );
nor \U$13961 ( \14093 , \14091 , \14092 );
xnor \U$13962 ( \14094 , \14093 , \8297 );
xor \U$13963 ( \14095 , \14090 , \14094 );
xor \U$13964 ( \14096 , \14081 , \14095 );
and \U$13965 ( \14097 , \307 , \9333 );
and \U$13966 ( \14098 , \412 , \9006 );
nor \U$13967 ( \14099 , \14097 , \14098 );
xnor \U$13968 ( \14100 , \14099 , \8848 );
and \U$13969 ( \14101 , \185 , \9765 );
and \U$13970 ( \14102 , \261 , \9644 );
nor \U$13971 ( \14103 , \14101 , \14102 );
xnor \U$13972 ( \14104 , \14103 , \9478 );
xor \U$13973 ( \14105 , \14100 , \14104 );
and \U$13974 ( \14106 , \197 , \10408 );
and \U$13975 ( \14107 , \178 , \10116 );
nor \U$13976 ( \14108 , \14106 , \14107 );
xnor \U$13977 ( \14109 , \14108 , \10121 );
xor \U$13978 ( \14110 , \14105 , \14109 );
xor \U$13979 ( \14111 , \14096 , \14110 );
xor \U$13980 ( \14112 , \14080 , \14111 );
xor \U$13981 ( \14113 , \14051 , \14112 );
not \U$13982 ( \14114 , \148 );
and \U$13983 ( \14115 , \10206 , \156 );
and \U$13984 ( \14116 , \10584 , \154 );
nor \U$13985 ( \14117 , \14115 , \14116 );
xnor \U$13986 ( \14118 , \14117 , \163 );
xor \U$13987 ( \14119 , \14114 , \14118 );
and \U$13988 ( \14120 , \9465 , \296 );
and \U$13989 ( \14121 , \9897 , \168 );
nor \U$13990 ( \14122 , \14120 , \14121 );
xnor \U$13991 ( \14123 , \14122 , \173 );
xor \U$13992 ( \14124 , \14119 , \14123 );
and \U$13993 ( \14125 , \8835 , \438 );
and \U$13994 ( \14126 , \9169 , \336 );
nor \U$13995 ( \14127 , \14125 , \14126 );
xnor \U$13996 ( \14128 , \14127 , \320 );
and \U$13997 ( \14129 , \8349 , \1086 );
and \U$13998 ( \14130 , \8652 , \508 );
nor \U$13999 ( \14131 , \14129 , \14130 );
xnor \U$14000 ( \14132 , \14131 , \487 );
xor \U$14001 ( \14133 , \14128 , \14132 );
and \U$14002 ( \14134 , \7700 , \1301 );
and \U$14003 ( \14135 , \8057 , \1246 );
nor \U$14004 ( \14136 , \14134 , \14135 );
xnor \U$14005 ( \14137 , \14136 , \1205 );
xor \U$14006 ( \14138 , \14133 , \14137 );
and \U$14007 ( \14139 , \5674 , \2400 );
and \U$14008 ( \14140 , \6030 , \2246 );
nor \U$14009 ( \14141 , \14139 , \14140 );
xnor \U$14010 ( \14142 , \14141 , \2195 );
and \U$14011 ( \14143 , \5156 , \2669 );
and \U$14012 ( \14144 , \5469 , \2538 );
nor \U$14013 ( \14145 , \14143 , \14144 );
xnor \U$14014 ( \14146 , \14145 , \2534 );
xor \U$14015 ( \14147 , \14142 , \14146 );
and \U$14016 ( \14148 , \4749 , \3103 );
and \U$14017 ( \14149 , \4922 , \2934 );
nor \U$14018 ( \14150 , \14148 , \14149 );
xnor \U$14019 ( \14151 , \14150 , \2839 );
xor \U$14020 ( \14152 , \14147 , \14151 );
xor \U$14021 ( \14153 , \14138 , \14152 );
and \U$14022 ( \14154 , \7231 , \1578 );
and \U$14023 ( \14155 , \7556 , \1431 );
nor \U$14024 ( \14156 , \14154 , \14155 );
xnor \U$14025 ( \14157 , \14156 , \1436 );
and \U$14026 ( \14158 , \6790 , \1824 );
and \U$14027 ( \14159 , \6945 , \1739 );
nor \U$14028 ( \14160 , \14158 , \14159 );
xnor \U$14029 ( \14161 , \14160 , \1697 );
xor \U$14030 ( \14162 , \14157 , \14161 );
and \U$14031 ( \14163 , \6281 , \2121 );
and \U$14032 ( \14164 , \6514 , \2008 );
nor \U$14033 ( \14165 , \14163 , \14164 );
xnor \U$14034 ( \14166 , \14165 , \1961 );
xor \U$14035 ( \14167 , \14162 , \14166 );
xor \U$14036 ( \14168 , \14153 , \14167 );
xor \U$14037 ( \14169 , \14124 , \14168 );
and \U$14038 ( \14170 , \2182 , \5996 );
and \U$14039 ( \14171 , \2366 , \5695 );
nor \U$14040 ( \14172 , \14170 , \14171 );
xnor \U$14041 ( \14173 , \14172 , \5687 );
and \U$14042 ( \14174 , \1948 , \6401 );
and \U$14043 ( \14175 , \2090 , \6143 );
nor \U$14044 ( \14176 , \14174 , \14175 );
xnor \U$14045 ( \14177 , \14176 , \6148 );
xor \U$14046 ( \14178 , \14173 , \14177 );
and \U$14047 ( \14179 , \1684 , \7055 );
and \U$14048 ( \14180 , \1802 , \6675 );
nor \U$14049 ( \14181 , \14179 , \14180 );
xnor \U$14050 ( \14182 , \14181 , \6680 );
xor \U$14051 ( \14183 , \14178 , \14182 );
and \U$14052 ( \14184 , \4364 , \3357 );
and \U$14053 ( \14185 , \4654 , \3255 );
nor \U$14054 ( \14186 , \14184 , \14185 );
xnor \U$14055 ( \14187 , \14186 , \3156 );
and \U$14056 ( \14188 , \3912 , \3813 );
and \U$14057 ( \14189 , \4160 , \3557 );
nor \U$14058 ( \14190 , \14188 , \14189 );
xnor \U$14059 ( \14191 , \14190 , \3562 );
xor \U$14060 ( \14192 , \14187 , \14191 );
and \U$14061 ( \14193 , \3646 , \4132 );
and \U$14062 ( \14194 , \3736 , \4012 );
nor \U$14063 ( \14195 , \14193 , \14194 );
xnor \U$14064 ( \14196 , \14195 , \3925 );
xor \U$14065 ( \14197 , \14192 , \14196 );
xor \U$14066 ( \14198 , \14183 , \14197 );
and \U$14067 ( \14199 , \3143 , \4581 );
and \U$14068 ( \14200 , \3395 , \4424 );
nor \U$14069 ( \14201 , \14199 , \14200 );
xnor \U$14070 ( \14202 , \14201 , \4377 );
and \U$14071 ( \14203 , \2826 , \5011 );
and \U$14072 ( \14204 , \3037 , \4878 );
nor \U$14073 ( \14205 , \14203 , \14204 );
xnor \U$14074 ( \14206 , \14205 , \4762 );
xor \U$14075 ( \14207 , \14202 , \14206 );
and \U$14076 ( \14208 , \2521 , \5485 );
and \U$14077 ( \14209 , \2757 , \5275 );
nor \U$14078 ( \14210 , \14208 , \14209 );
xnor \U$14079 ( \14211 , \14210 , \5169 );
xor \U$14080 ( \14212 , \14207 , \14211 );
xor \U$14081 ( \14213 , \14198 , \14212 );
xor \U$14082 ( \14214 , \14169 , \14213 );
xor \U$14083 ( \14215 , \14113 , \14214 );
xor \U$14084 ( \14216 , \14040 , \14215 );
xor \U$14085 ( \14217 , \14001 , \14216 );
xor \U$14086 ( \14218 , \13987 , \14217 );
xor \U$14087 ( \14219 , \13958 , \14218 );
and \U$14088 ( \14220 , \13677 , \13942 );
xor \U$14089 ( \14221 , \14219 , \14220 );
and \U$14090 ( \14222 , \13943 , \13947 );
and \U$14091 ( \14223 , \13948 , \13951 );
or \U$14092 ( \14224 , \14222 , \14223 );
xor \U$14093 ( \14225 , \14221 , \14224 );
buf \U$14094 ( \14226 , \14225 );
buf \U$14095 ( \14227 , \14226 );
and \U$14096 ( \14228 , \13962 , \13986 );
and \U$14097 ( \14229 , \13986 , \14217 );
and \U$14098 ( \14230 , \13962 , \14217 );
or \U$14099 ( \14231 , \14228 , \14229 , \14230 );
and \U$14100 ( \14232 , \13966 , \13970 );
and \U$14101 ( \14233 , \13970 , \13985 );
and \U$14102 ( \14234 , \13966 , \13985 );
or \U$14103 ( \14235 , \14232 , \14233 , \14234 );
and \U$14104 ( \14236 , \14001 , \14216 );
xor \U$14105 ( \14237 , \14235 , \14236 );
and \U$14106 ( \14238 , \13975 , \13979 );
and \U$14107 ( \14239 , \13979 , \13984 );
and \U$14108 ( \14240 , \13975 , \13984 );
or \U$14109 ( \14241 , \14238 , \14239 , \14240 );
and \U$14110 ( \14242 , \14019 , \14023 );
and \U$14111 ( \14243 , \14023 , \14038 );
and \U$14112 ( \14244 , \14019 , \14038 );
or \U$14113 ( \14245 , \14242 , \14243 , \14244 );
xor \U$14114 ( \14246 , \14241 , \14245 );
and \U$14115 ( \14247 , \14051 , \14112 );
and \U$14116 ( \14248 , \14112 , \14214 );
and \U$14117 ( \14249 , \14051 , \14214 );
or \U$14118 ( \14250 , \14247 , \14248 , \14249 );
xor \U$14119 ( \14251 , \14246 , \14250 );
xor \U$14120 ( \14252 , \14237 , \14251 );
xor \U$14121 ( \14253 , \14231 , \14252 );
and \U$14122 ( \14254 , \13991 , \13995 );
and \U$14123 ( \14255 , \13995 , \14000 );
and \U$14124 ( \14256 , \13991 , \14000 );
or \U$14125 ( \14257 , \14254 , \14255 , \14256 );
and \U$14126 ( \14258 , \14015 , \14039 );
and \U$14127 ( \14259 , \14039 , \14215 );
and \U$14128 ( \14260 , \14015 , \14215 );
or \U$14129 ( \14261 , \14258 , \14259 , \14260 );
xor \U$14130 ( \14262 , \14257 , \14261 );
and \U$14131 ( \14263 , \14005 , \14009 );
and \U$14132 ( \14264 , \14009 , \14014 );
and \U$14133 ( \14265 , \14005 , \14014 );
or \U$14134 ( \14266 , \14263 , \14264 , \14265 );
and \U$14135 ( \14267 , \14044 , \14048 );
and \U$14136 ( \14268 , \14048 , \14050 );
and \U$14137 ( \14269 , \14044 , \14050 );
or \U$14138 ( \14270 , \14267 , \14268 , \14269 );
xor \U$14139 ( \14271 , \14266 , \14270 );
and \U$14140 ( \14272 , \14124 , \14168 );
and \U$14141 ( \14273 , \14168 , \14213 );
and \U$14142 ( \14274 , \14124 , \14213 );
or \U$14143 ( \14275 , \14272 , \14273 , \14274 );
xor \U$14144 ( \14276 , \14271 , \14275 );
and \U$14145 ( \14277 , \14055 , \14059 );
and \U$14146 ( \14278 , \14059 , \14064 );
and \U$14147 ( \14279 , \14055 , \14064 );
or \U$14148 ( \14280 , \14277 , \14278 , \14279 );
and \U$14149 ( \14281 , \14028 , \14032 );
and \U$14150 ( \14282 , \14032 , \14037 );
and \U$14151 ( \14283 , \14028 , \14037 );
or \U$14152 ( \14284 , \14281 , \14282 , \14283 );
xor \U$14153 ( \14285 , \14280 , \14284 );
and \U$14154 ( \14286 , \14069 , \14073 );
and \U$14155 ( \14287 , \14073 , \14078 );
and \U$14156 ( \14288 , \14069 , \14078 );
or \U$14157 ( \14289 , \14286 , \14287 , \14288 );
xor \U$14158 ( \14290 , \14285 , \14289 );
and \U$14159 ( \14291 , \14138 , \14152 );
and \U$14160 ( \14292 , \14152 , \14167 );
and \U$14161 ( \14293 , \14138 , \14167 );
or \U$14162 ( \14294 , \14291 , \14292 , \14293 );
and \U$14163 ( \14295 , \14081 , \14095 );
and \U$14164 ( \14296 , \14095 , \14110 );
and \U$14165 ( \14297 , \14081 , \14110 );
or \U$14166 ( \14298 , \14295 , \14296 , \14297 );
xor \U$14167 ( \14299 , \14294 , \14298 );
and \U$14168 ( \14300 , \14183 , \14197 );
and \U$14169 ( \14301 , \14197 , \14212 );
and \U$14170 ( \14302 , \14183 , \14212 );
or \U$14171 ( \14303 , \14300 , \14301 , \14302 );
xor \U$14172 ( \14304 , \14299 , \14303 );
xor \U$14173 ( \14305 , \14290 , \14304 );
and \U$14174 ( \14306 , \10584 , \156 );
not \U$14175 ( \14307 , \14306 );
xnor \U$14176 ( \14308 , \14307 , \163 );
and \U$14177 ( \14309 , \9897 , \296 );
and \U$14178 ( \14310 , \10206 , \168 );
nor \U$14179 ( \14311 , \14309 , \14310 );
xnor \U$14180 ( \14312 , \14311 , \173 );
xor \U$14181 ( \14313 , \14308 , \14312 );
and \U$14182 ( \14314 , \9169 , \438 );
and \U$14183 ( \14315 , \9465 , \336 );
nor \U$14184 ( \14316 , \14314 , \14315 );
xnor \U$14185 ( \14317 , \14316 , \320 );
xor \U$14186 ( \14318 , \14313 , \14317 );
and \U$14187 ( \14319 , \8652 , \1086 );
and \U$14188 ( \14320 , \8835 , \508 );
nor \U$14189 ( \14321 , \14319 , \14320 );
xnor \U$14190 ( \14322 , \14321 , \487 );
and \U$14191 ( \14323 , \8057 , \1301 );
and \U$14192 ( \14324 , \8349 , \1246 );
nor \U$14193 ( \14325 , \14323 , \14324 );
xnor \U$14194 ( \14326 , \14325 , \1205 );
xor \U$14195 ( \14327 , \14322 , \14326 );
and \U$14196 ( \14328 , \7556 , \1578 );
and \U$14197 ( \14329 , \7700 , \1431 );
nor \U$14198 ( \14330 , \14328 , \14329 );
xnor \U$14199 ( \14331 , \14330 , \1436 );
xor \U$14200 ( \14332 , \14327 , \14331 );
and \U$14201 ( \14333 , \5469 , \2669 );
and \U$14202 ( \14334 , \5674 , \2538 );
nor \U$14203 ( \14335 , \14333 , \14334 );
xnor \U$14204 ( \14336 , \14335 , \2534 );
and \U$14205 ( \14337 , \4922 , \3103 );
and \U$14206 ( \14338 , \5156 , \2934 );
nor \U$14207 ( \14339 , \14337 , \14338 );
xnor \U$14208 ( \14340 , \14339 , \2839 );
xor \U$14209 ( \14341 , \14336 , \14340 );
and \U$14210 ( \14342 , \4654 , \3357 );
and \U$14211 ( \14343 , \4749 , \3255 );
nor \U$14212 ( \14344 , \14342 , \14343 );
xnor \U$14213 ( \14345 , \14344 , \3156 );
xor \U$14214 ( \14346 , \14341 , \14345 );
xor \U$14215 ( \14347 , \14332 , \14346 );
and \U$14216 ( \14348 , \6945 , \1824 );
and \U$14217 ( \14349 , \7231 , \1739 );
nor \U$14218 ( \14350 , \14348 , \14349 );
xnor \U$14219 ( \14351 , \14350 , \1697 );
and \U$14220 ( \14352 , \6514 , \2121 );
and \U$14221 ( \14353 , \6790 , \2008 );
nor \U$14222 ( \14354 , \14352 , \14353 );
xnor \U$14223 ( \14355 , \14354 , \1961 );
xor \U$14224 ( \14356 , \14351 , \14355 );
and \U$14225 ( \14357 , \6030 , \2400 );
and \U$14226 ( \14358 , \6281 , \2246 );
nor \U$14227 ( \14359 , \14357 , \14358 );
xnor \U$14228 ( \14360 , \14359 , \2195 );
xor \U$14229 ( \14361 , \14356 , \14360 );
xor \U$14230 ( \14362 , \14347 , \14361 );
xor \U$14231 ( \14363 , \14318 , \14362 );
and \U$14232 ( \14364 , \4160 , \3813 );
and \U$14233 ( \14365 , \4364 , \3557 );
nor \U$14234 ( \14366 , \14364 , \14365 );
xnor \U$14235 ( \14367 , \14366 , \3562 );
and \U$14236 ( \14368 , \3736 , \4132 );
and \U$14237 ( \14369 , \3912 , \4012 );
nor \U$14238 ( \14370 , \14368 , \14369 );
xnor \U$14239 ( \14371 , \14370 , \3925 );
xor \U$14240 ( \14372 , \14367 , \14371 );
and \U$14241 ( \14373 , \3395 , \4581 );
and \U$14242 ( \14374 , \3646 , \4424 );
nor \U$14243 ( \14375 , \14373 , \14374 );
xnor \U$14244 ( \14376 , \14375 , \4377 );
xor \U$14245 ( \14377 , \14372 , \14376 );
and \U$14246 ( \14378 , \2090 , \6401 );
and \U$14247 ( \14379 , \2182 , \6143 );
nor \U$14248 ( \14380 , \14378 , \14379 );
xnor \U$14249 ( \14381 , \14380 , \6148 );
and \U$14250 ( \14382 , \1802 , \7055 );
and \U$14251 ( \14383 , \1948 , \6675 );
nor \U$14252 ( \14384 , \14382 , \14383 );
xnor \U$14253 ( \14385 , \14384 , \6680 );
xor \U$14254 ( \14386 , \14381 , \14385 );
and \U$14255 ( \14387 , \1601 , \7489 );
and \U$14256 ( \14388 , \1684 , \7137 );
nor \U$14257 ( \14389 , \14387 , \14388 );
xnor \U$14258 ( \14390 , \14389 , \7142 );
xor \U$14259 ( \14391 , \14386 , \14390 );
xor \U$14260 ( \14392 , \14377 , \14391 );
and \U$14261 ( \14393 , \3037 , \5011 );
and \U$14262 ( \14394 , \3143 , \4878 );
nor \U$14263 ( \14395 , \14393 , \14394 );
xnor \U$14264 ( \14396 , \14395 , \4762 );
and \U$14265 ( \14397 , \2757 , \5485 );
and \U$14266 ( \14398 , \2826 , \5275 );
nor \U$14267 ( \14399 , \14397 , \14398 );
xnor \U$14268 ( \14400 , \14399 , \5169 );
xor \U$14269 ( \14401 , \14396 , \14400 );
and \U$14270 ( \14402 , \2366 , \5996 );
and \U$14271 ( \14403 , \2521 , \5695 );
nor \U$14272 ( \14404 , \14402 , \14403 );
xnor \U$14273 ( \14405 , \14404 , \5687 );
xor \U$14274 ( \14406 , \14401 , \14405 );
xor \U$14275 ( \14407 , \14392 , \14406 );
xor \U$14276 ( \14408 , \14363 , \14407 );
xor \U$14277 ( \14409 , \14305 , \14408 );
xor \U$14278 ( \14410 , \14276 , \14409 );
and \U$14279 ( \14411 , \14065 , \14079 );
and \U$14280 ( \14412 , \14079 , \14111 );
and \U$14281 ( \14413 , \14065 , \14111 );
or \U$14282 ( \14414 , \14411 , \14412 , \14413 );
and \U$14283 ( \14415 , \14128 , \14132 );
and \U$14284 ( \14416 , \14132 , \14137 );
and \U$14285 ( \14417 , \14128 , \14137 );
or \U$14286 ( \14418 , \14415 , \14416 , \14417 );
and \U$14287 ( \14419 , \14114 , \14118 );
and \U$14288 ( \14420 , \14118 , \14123 );
and \U$14289 ( \14421 , \14114 , \14123 );
or \U$14290 ( \14422 , \14419 , \14420 , \14421 );
xor \U$14291 ( \14423 , \14418 , \14422 );
and \U$14292 ( \14424 , \14157 , \14161 );
and \U$14293 ( \14425 , \14161 , \14166 );
and \U$14294 ( \14426 , \14157 , \14166 );
or \U$14295 ( \14427 , \14424 , \14425 , \14426 );
xor \U$14296 ( \14428 , \14423 , \14427 );
xor \U$14297 ( \14429 , \14414 , \14428 );
and \U$14298 ( \14430 , \14187 , \14191 );
and \U$14299 ( \14431 , \14191 , \14196 );
and \U$14300 ( \14432 , \14187 , \14196 );
or \U$14301 ( \14433 , \14430 , \14431 , \14432 );
and \U$14302 ( \14434 , \14142 , \14146 );
and \U$14303 ( \14435 , \14146 , \14151 );
and \U$14304 ( \14436 , \14142 , \14151 );
or \U$14305 ( \14437 , \14434 , \14435 , \14436 );
xor \U$14306 ( \14438 , \14433 , \14437 );
and \U$14307 ( \14439 , \14202 , \14206 );
and \U$14308 ( \14440 , \14206 , \14211 );
and \U$14309 ( \14441 , \14202 , \14211 );
or \U$14310 ( \14442 , \14439 , \14440 , \14441 );
xor \U$14311 ( \14443 , \14438 , \14442 );
and \U$14312 ( \14444 , \14173 , \14177 );
and \U$14313 ( \14445 , \14177 , \14182 );
and \U$14314 ( \14446 , \14173 , \14182 );
or \U$14315 ( \14447 , \14444 , \14445 , \14446 );
and \U$14316 ( \14448 , \14085 , \14089 );
and \U$14317 ( \14449 , \14089 , \14094 );
and \U$14318 ( \14450 , \14085 , \14094 );
or \U$14319 ( \14451 , \14448 , \14449 , \14450 );
xor \U$14320 ( \14452 , \14447 , \14451 );
and \U$14321 ( \14453 , \14100 , \14104 );
and \U$14322 ( \14454 , \14104 , \14109 );
and \U$14323 ( \14455 , \14100 , \14109 );
or \U$14324 ( \14456 , \14453 , \14454 , \14455 );
xor \U$14325 ( \14457 , \14452 , \14456 );
xor \U$14326 ( \14458 , \14443 , \14457 );
and \U$14327 ( \14459 , \261 , \9765 );
and \U$14328 ( \14460 , \307 , \9644 );
nor \U$14329 ( \14461 , \14459 , \14460 );
xnor \U$14330 ( \14462 , \14461 , \9478 );
and \U$14331 ( \14463 , \178 , \10408 );
and \U$14332 ( \14464 , \185 , \10116 );
nor \U$14333 ( \14465 , \14463 , \14464 );
xnor \U$14334 ( \14466 , \14465 , \10121 );
xor \U$14335 ( \14467 , \14462 , \14466 );
and \U$14336 ( \14468 , \197 , \10118 );
xor \U$14337 ( \14469 , \14467 , \14468 );
and \U$14338 ( \14470 , \1333 , \8019 );
and \U$14339 ( \14471 , \1484 , \7830 );
nor \U$14340 ( \14472 , \14470 , \14471 );
xnor \U$14341 ( \14473 , \14472 , \7713 );
and \U$14342 ( \14474 , \1147 , \8540 );
and \U$14343 ( \14475 , \1192 , \8292 );
nor \U$14344 ( \14476 , \14474 , \14475 );
xnor \U$14345 ( \14477 , \14476 , \8297 );
xor \U$14346 ( \14478 , \14473 , \14477 );
and \U$14347 ( \14479 , \412 , \9333 );
and \U$14348 ( \14480 , \474 , \9006 );
nor \U$14349 ( \14481 , \14479 , \14480 );
xnor \U$14350 ( \14482 , \14481 , \8848 );
xor \U$14351 ( \14483 , \14478 , \14482 );
xnor \U$14352 ( \14484 , \14469 , \14483 );
xor \U$14353 ( \14485 , \14458 , \14484 );
xor \U$14354 ( \14486 , \14429 , \14485 );
xor \U$14355 ( \14487 , \14410 , \14486 );
xor \U$14356 ( \14488 , \14262 , \14487 );
xor \U$14357 ( \14489 , \14253 , \14488 );
and \U$14358 ( \14490 , \13958 , \14218 );
xor \U$14359 ( \14491 , \14489 , \14490 );
and \U$14360 ( \14492 , \14219 , \14220 );
and \U$14361 ( \14493 , \14221 , \14224 );
or \U$14362 ( \14494 , \14492 , \14493 );
xor \U$14363 ( \14495 , \14491 , \14494 );
buf \U$14364 ( \14496 , \14495 );
buf \U$14365 ( \14497 , \14496 );
and \U$14366 ( \14498 , \14235 , \14236 );
and \U$14367 ( \14499 , \14236 , \14251 );
and \U$14368 ( \14500 , \14235 , \14251 );
or \U$14369 ( \14501 , \14498 , \14499 , \14500 );
and \U$14370 ( \14502 , \14257 , \14261 );
and \U$14371 ( \14503 , \14261 , \14487 );
and \U$14372 ( \14504 , \14257 , \14487 );
or \U$14373 ( \14505 , \14502 , \14503 , \14504 );
and \U$14374 ( \14506 , \14266 , \14270 );
and \U$14375 ( \14507 , \14270 , \14275 );
and \U$14376 ( \14508 , \14266 , \14275 );
or \U$14377 ( \14509 , \14506 , \14507 , \14508 );
and \U$14378 ( \14510 , \14290 , \14304 );
and \U$14379 ( \14511 , \14304 , \14408 );
and \U$14380 ( \14512 , \14290 , \14408 );
or \U$14381 ( \14513 , \14510 , \14511 , \14512 );
xor \U$14382 ( \14514 , \14509 , \14513 );
and \U$14383 ( \14515 , \14414 , \14428 );
and \U$14384 ( \14516 , \14428 , \14485 );
and \U$14385 ( \14517 , \14414 , \14485 );
or \U$14386 ( \14518 , \14515 , \14516 , \14517 );
xor \U$14387 ( \14519 , \14514 , \14518 );
xor \U$14388 ( \14520 , \14505 , \14519 );
and \U$14389 ( \14521 , \14241 , \14245 );
and \U$14390 ( \14522 , \14245 , \14250 );
and \U$14391 ( \14523 , \14241 , \14250 );
or \U$14392 ( \14524 , \14521 , \14522 , \14523 );
and \U$14393 ( \14525 , \14276 , \14409 );
and \U$14394 ( \14526 , \14409 , \14486 );
and \U$14395 ( \14527 , \14276 , \14486 );
or \U$14396 ( \14528 , \14525 , \14526 , \14527 );
xor \U$14397 ( \14529 , \14524 , \14528 );
and \U$14398 ( \14530 , \14280 , \14284 );
and \U$14399 ( \14531 , \14284 , \14289 );
and \U$14400 ( \14532 , \14280 , \14289 );
or \U$14401 ( \14533 , \14530 , \14531 , \14532 );
and \U$14402 ( \14534 , \14294 , \14298 );
and \U$14403 ( \14535 , \14298 , \14303 );
and \U$14404 ( \14536 , \14294 , \14303 );
or \U$14405 ( \14537 , \14534 , \14535 , \14536 );
xor \U$14406 ( \14538 , \14533 , \14537 );
and \U$14407 ( \14539 , \14318 , \14362 );
and \U$14408 ( \14540 , \14362 , \14407 );
and \U$14409 ( \14541 , \14318 , \14407 );
or \U$14410 ( \14542 , \14539 , \14540 , \14541 );
xor \U$14411 ( \14543 , \14538 , \14542 );
and \U$14412 ( \14544 , \14443 , \14457 );
and \U$14413 ( \14545 , \14457 , \14484 );
and \U$14414 ( \14546 , \14443 , \14484 );
or \U$14415 ( \14547 , \14544 , \14545 , \14546 );
and \U$14416 ( \14548 , \14381 , \14385 );
and \U$14417 ( \14549 , \14385 , \14390 );
and \U$14418 ( \14550 , \14381 , \14390 );
or \U$14419 ( \14551 , \14548 , \14549 , \14550 );
and \U$14420 ( \14552 , \14462 , \14466 );
and \U$14421 ( \14553 , \14466 , \14468 );
and \U$14422 ( \14554 , \14462 , \14468 );
or \U$14423 ( \14555 , \14552 , \14553 , \14554 );
xor \U$14424 ( \14556 , \14551 , \14555 );
and \U$14425 ( \14557 , \14473 , \14477 );
and \U$14426 ( \14558 , \14477 , \14482 );
and \U$14427 ( \14559 , \14473 , \14482 );
or \U$14428 ( \14560 , \14557 , \14558 , \14559 );
xor \U$14429 ( \14561 , \14556 , \14560 );
and \U$14430 ( \14562 , \14322 , \14326 );
and \U$14431 ( \14563 , \14326 , \14331 );
and \U$14432 ( \14564 , \14322 , \14331 );
or \U$14433 ( \14565 , \14562 , \14563 , \14564 );
and \U$14434 ( \14566 , \14351 , \14355 );
and \U$14435 ( \14567 , \14355 , \14360 );
and \U$14436 ( \14568 , \14351 , \14360 );
or \U$14437 ( \14569 , \14566 , \14567 , \14568 );
xor \U$14438 ( \14570 , \14565 , \14569 );
and \U$14439 ( \14571 , \14308 , \14312 );
and \U$14440 ( \14572 , \14312 , \14317 );
and \U$14441 ( \14573 , \14308 , \14317 );
or \U$14442 ( \14574 , \14571 , \14572 , \14573 );
xor \U$14443 ( \14575 , \14570 , \14574 );
xor \U$14444 ( \14576 , \14561 , \14575 );
and \U$14445 ( \14577 , \14336 , \14340 );
and \U$14446 ( \14578 , \14340 , \14345 );
and \U$14447 ( \14579 , \14336 , \14345 );
or \U$14448 ( \14580 , \14577 , \14578 , \14579 );
and \U$14449 ( \14581 , \14367 , \14371 );
and \U$14450 ( \14582 , \14371 , \14376 );
and \U$14451 ( \14583 , \14367 , \14376 );
or \U$14452 ( \14584 , \14581 , \14582 , \14583 );
xor \U$14453 ( \14585 , \14580 , \14584 );
and \U$14454 ( \14586 , \14396 , \14400 );
and \U$14455 ( \14587 , \14400 , \14405 );
and \U$14456 ( \14588 , \14396 , \14405 );
or \U$14457 ( \14589 , \14586 , \14587 , \14588 );
xor \U$14458 ( \14590 , \14585 , \14589 );
xor \U$14459 ( \14591 , \14576 , \14590 );
xor \U$14460 ( \14592 , \14547 , \14591 );
and \U$14461 ( \14593 , \307 , \9765 );
and \U$14462 ( \14594 , \412 , \9644 );
nor \U$14463 ( \14595 , \14593 , \14594 );
xnor \U$14464 ( \14596 , \14595 , \9478 );
and \U$14465 ( \14597 , \185 , \10408 );
and \U$14466 ( \14598 , \261 , \10116 );
nor \U$14467 ( \14599 , \14597 , \14598 );
xnor \U$14468 ( \14600 , \14599 , \10121 );
xor \U$14469 ( \14601 , \14596 , \14600 );
and \U$14470 ( \14602 , \178 , \10118 );
xor \U$14471 ( \14603 , \14601 , \14602 );
and \U$14472 ( \14604 , \2182 , \6401 );
and \U$14473 ( \14605 , \2366 , \6143 );
nor \U$14474 ( \14606 , \14604 , \14605 );
xnor \U$14475 ( \14607 , \14606 , \6148 );
and \U$14476 ( \14608 , \1948 , \7055 );
and \U$14477 ( \14609 , \2090 , \6675 );
nor \U$14478 ( \14610 , \14608 , \14609 );
xnor \U$14479 ( \14611 , \14610 , \6680 );
xor \U$14480 ( \14612 , \14607 , \14611 );
and \U$14481 ( \14613 , \1684 , \7489 );
and \U$14482 ( \14614 , \1802 , \7137 );
nor \U$14483 ( \14615 , \14613 , \14614 );
xnor \U$14484 ( \14616 , \14615 , \7142 );
xor \U$14485 ( \14617 , \14612 , \14616 );
xor \U$14486 ( \14618 , \14603 , \14617 );
and \U$14487 ( \14619 , \1484 , \8019 );
and \U$14488 ( \14620 , \1601 , \7830 );
nor \U$14489 ( \14621 , \14619 , \14620 );
xnor \U$14490 ( \14622 , \14621 , \7713 );
and \U$14491 ( \14623 , \1192 , \8540 );
and \U$14492 ( \14624 , \1333 , \8292 );
nor \U$14493 ( \14625 , \14623 , \14624 );
xnor \U$14494 ( \14626 , \14625 , \8297 );
xor \U$14495 ( \14627 , \14622 , \14626 );
and \U$14496 ( \14628 , \474 , \9333 );
and \U$14497 ( \14629 , \1147 , \9006 );
nor \U$14498 ( \14630 , \14628 , \14629 );
xnor \U$14499 ( \14631 , \14630 , \8848 );
xor \U$14500 ( \14632 , \14627 , \14631 );
xor \U$14501 ( \14633 , \14618 , \14632 );
and \U$14502 ( \14634 , \5674 , \2669 );
and \U$14503 ( \14635 , \6030 , \2538 );
nor \U$14504 ( \14636 , \14634 , \14635 );
xnor \U$14505 ( \14637 , \14636 , \2534 );
and \U$14506 ( \14638 , \5156 , \3103 );
and \U$14507 ( \14639 , \5469 , \2934 );
nor \U$14508 ( \14640 , \14638 , \14639 );
xnor \U$14509 ( \14641 , \14640 , \2839 );
xor \U$14510 ( \14642 , \14637 , \14641 );
and \U$14511 ( \14643 , \4749 , \3357 );
and \U$14512 ( \14644 , \4922 , \3255 );
nor \U$14513 ( \14645 , \14643 , \14644 );
xnor \U$14514 ( \14646 , \14645 , \3156 );
xor \U$14515 ( \14647 , \14642 , \14646 );
and \U$14516 ( \14648 , \4364 , \3813 );
and \U$14517 ( \14649 , \4654 , \3557 );
nor \U$14518 ( \14650 , \14648 , \14649 );
xnor \U$14519 ( \14651 , \14650 , \3562 );
and \U$14520 ( \14652 , \3912 , \4132 );
and \U$14521 ( \14653 , \4160 , \4012 );
nor \U$14522 ( \14654 , \14652 , \14653 );
xnor \U$14523 ( \14655 , \14654 , \3925 );
xor \U$14524 ( \14656 , \14651 , \14655 );
and \U$14525 ( \14657 , \3646 , \4581 );
and \U$14526 ( \14658 , \3736 , \4424 );
nor \U$14527 ( \14659 , \14657 , \14658 );
xnor \U$14528 ( \14660 , \14659 , \4377 );
xor \U$14529 ( \14661 , \14656 , \14660 );
xor \U$14530 ( \14662 , \14647 , \14661 );
and \U$14531 ( \14663 , \3143 , \5011 );
and \U$14532 ( \14664 , \3395 , \4878 );
nor \U$14533 ( \14665 , \14663 , \14664 );
xnor \U$14534 ( \14666 , \14665 , \4762 );
and \U$14535 ( \14667 , \2826 , \5485 );
and \U$14536 ( \14668 , \3037 , \5275 );
nor \U$14537 ( \14669 , \14667 , \14668 );
xnor \U$14538 ( \14670 , \14669 , \5169 );
xor \U$14539 ( \14671 , \14666 , \14670 );
and \U$14540 ( \14672 , \2521 , \5996 );
and \U$14541 ( \14673 , \2757 , \5695 );
nor \U$14542 ( \14674 , \14672 , \14673 );
xnor \U$14543 ( \14675 , \14674 , \5687 );
xor \U$14544 ( \14676 , \14671 , \14675 );
xor \U$14545 ( \14677 , \14662 , \14676 );
xor \U$14546 ( \14678 , \14633 , \14677 );
and \U$14547 ( \14679 , \8835 , \1086 );
and \U$14548 ( \14680 , \9169 , \508 );
nor \U$14549 ( \14681 , \14679 , \14680 );
xnor \U$14550 ( \14682 , \14681 , \487 );
and \U$14551 ( \14683 , \8349 , \1301 );
and \U$14552 ( \14684 , \8652 , \1246 );
nor \U$14553 ( \14685 , \14683 , \14684 );
xnor \U$14554 ( \14686 , \14685 , \1205 );
xor \U$14555 ( \14687 , \14682 , \14686 );
and \U$14556 ( \14688 , \7700 , \1578 );
and \U$14557 ( \14689 , \8057 , \1431 );
nor \U$14558 ( \14690 , \14688 , \14689 );
xnor \U$14559 ( \14691 , \14690 , \1436 );
xor \U$14560 ( \14692 , \14687 , \14691 );
and \U$14561 ( \14693 , \7231 , \1824 );
and \U$14562 ( \14694 , \7556 , \1739 );
nor \U$14563 ( \14695 , \14693 , \14694 );
xnor \U$14564 ( \14696 , \14695 , \1697 );
and \U$14565 ( \14697 , \6790 , \2121 );
and \U$14566 ( \14698 , \6945 , \2008 );
nor \U$14567 ( \14699 , \14697 , \14698 );
xnor \U$14568 ( \14700 , \14699 , \1961 );
xor \U$14569 ( \14701 , \14696 , \14700 );
and \U$14570 ( \14702 , \6281 , \2400 );
and \U$14571 ( \14703 , \6514 , \2246 );
nor \U$14572 ( \14704 , \14702 , \14703 );
xnor \U$14573 ( \14705 , \14704 , \2195 );
xor \U$14574 ( \14706 , \14701 , \14705 );
xor \U$14575 ( \14707 , \14692 , \14706 );
not \U$14576 ( \14708 , \163 );
and \U$14577 ( \14709 , \10206 , \296 );
and \U$14578 ( \14710 , \10584 , \168 );
nor \U$14579 ( \14711 , \14709 , \14710 );
xnor \U$14580 ( \14712 , \14711 , \173 );
xor \U$14581 ( \14713 , \14708 , \14712 );
and \U$14582 ( \14714 , \9465 , \438 );
and \U$14583 ( \14715 , \9897 , \336 );
nor \U$14584 ( \14716 , \14714 , \14715 );
xnor \U$14585 ( \14717 , \14716 , \320 );
xor \U$14586 ( \14718 , \14713 , \14717 );
xor \U$14587 ( \14719 , \14707 , \14718 );
xor \U$14588 ( \14720 , \14678 , \14719 );
xor \U$14589 ( \14721 , \14592 , \14720 );
xor \U$14590 ( \14722 , \14543 , \14721 );
and \U$14591 ( \14723 , \14332 , \14346 );
and \U$14592 ( \14724 , \14346 , \14361 );
and \U$14593 ( \14725 , \14332 , \14361 );
or \U$14594 ( \14726 , \14723 , \14724 , \14725 );
and \U$14595 ( \14727 , \14377 , \14391 );
and \U$14596 ( \14728 , \14391 , \14406 );
and \U$14597 ( \14729 , \14377 , \14406 );
or \U$14598 ( \14730 , \14727 , \14728 , \14729 );
xor \U$14599 ( \14731 , \14726 , \14730 );
or \U$14600 ( \14732 , \14469 , \14483 );
xor \U$14601 ( \14733 , \14731 , \14732 );
and \U$14602 ( \14734 , \14433 , \14437 );
and \U$14603 ( \14735 , \14437 , \14442 );
and \U$14604 ( \14736 , \14433 , \14442 );
or \U$14605 ( \14737 , \14734 , \14735 , \14736 );
and \U$14606 ( \14738 , \14418 , \14422 );
and \U$14607 ( \14739 , \14422 , \14427 );
and \U$14608 ( \14740 , \14418 , \14427 );
or \U$14609 ( \14741 , \14738 , \14739 , \14740 );
xor \U$14610 ( \14742 , \14737 , \14741 );
and \U$14611 ( \14743 , \14447 , \14451 );
and \U$14612 ( \14744 , \14451 , \14456 );
and \U$14613 ( \14745 , \14447 , \14456 );
or \U$14614 ( \14746 , \14743 , \14744 , \14745 );
xor \U$14615 ( \14747 , \14742 , \14746 );
xor \U$14616 ( \14748 , \14733 , \14747 );
xor \U$14617 ( \14749 , \14722 , \14748 );
xor \U$14618 ( \14750 , \14529 , \14749 );
xor \U$14619 ( \14751 , \14520 , \14750 );
xor \U$14620 ( \14752 , \14501 , \14751 );
and \U$14621 ( \14753 , \14231 , \14252 );
and \U$14622 ( \14754 , \14252 , \14488 );
and \U$14623 ( \14755 , \14231 , \14488 );
or \U$14624 ( \14756 , \14753 , \14754 , \14755 );
xor \U$14625 ( \14757 , \14752 , \14756 );
and \U$14626 ( \14758 , \14489 , \14490 );
and \U$14627 ( \14759 , \14491 , \14494 );
or \U$14628 ( \14760 , \14758 , \14759 );
xor \U$14629 ( \14761 , \14757 , \14760 );
buf \U$14630 ( \14762 , \14761 );
buf \U$14631 ( \14763 , \14762 );
and \U$14632 ( \14764 , \14505 , \14519 );
and \U$14633 ( \14765 , \14519 , \14750 );
and \U$14634 ( \14766 , \14505 , \14750 );
or \U$14635 ( \14767 , \14764 , \14765 , \14766 );
and \U$14636 ( \14768 , \14524 , \14528 );
and \U$14637 ( \14769 , \14528 , \14749 );
and \U$14638 ( \14770 , \14524 , \14749 );
or \U$14639 ( \14771 , \14768 , \14769 , \14770 );
and \U$14640 ( \14772 , \14533 , \14537 );
and \U$14641 ( \14773 , \14537 , \14542 );
and \U$14642 ( \14774 , \14533 , \14542 );
or \U$14643 ( \14775 , \14772 , \14773 , \14774 );
and \U$14644 ( \14776 , \14547 , \14591 );
and \U$14645 ( \14777 , \14591 , \14720 );
and \U$14646 ( \14778 , \14547 , \14720 );
or \U$14647 ( \14779 , \14776 , \14777 , \14778 );
xor \U$14648 ( \14780 , \14775 , \14779 );
and \U$14649 ( \14781 , \14733 , \14747 );
xor \U$14650 ( \14782 , \14780 , \14781 );
xor \U$14651 ( \14783 , \14771 , \14782 );
and \U$14652 ( \14784 , \14509 , \14513 );
and \U$14653 ( \14785 , \14513 , \14518 );
and \U$14654 ( \14786 , \14509 , \14518 );
or \U$14655 ( \14787 , \14784 , \14785 , \14786 );
and \U$14656 ( \14788 , \14543 , \14721 );
and \U$14657 ( \14789 , \14721 , \14748 );
and \U$14658 ( \14790 , \14543 , \14748 );
or \U$14659 ( \14791 , \14788 , \14789 , \14790 );
xor \U$14660 ( \14792 , \14787 , \14791 );
and \U$14661 ( \14793 , \14726 , \14730 );
and \U$14662 ( \14794 , \14730 , \14732 );
and \U$14663 ( \14795 , \14726 , \14732 );
or \U$14664 ( \14796 , \14793 , \14794 , \14795 );
and \U$14665 ( \14797 , \14737 , \14741 );
and \U$14666 ( \14798 , \14741 , \14746 );
and \U$14667 ( \14799 , \14737 , \14746 );
or \U$14668 ( \14800 , \14797 , \14798 , \14799 );
xor \U$14669 ( \14801 , \14796 , \14800 );
and \U$14670 ( \14802 , \14633 , \14677 );
and \U$14671 ( \14803 , \14677 , \14719 );
and \U$14672 ( \14804 , \14633 , \14719 );
or \U$14673 ( \14805 , \14802 , \14803 , \14804 );
xor \U$14674 ( \14806 , \14801 , \14805 );
and \U$14675 ( \14807 , \14561 , \14575 );
and \U$14676 ( \14808 , \14575 , \14590 );
and \U$14677 ( \14809 , \14561 , \14590 );
or \U$14678 ( \14810 , \14807 , \14808 , \14809 );
and \U$14679 ( \14811 , \14637 , \14641 );
and \U$14680 ( \14812 , \14641 , \14646 );
and \U$14681 ( \14813 , \14637 , \14646 );
or \U$14682 ( \14814 , \14811 , \14812 , \14813 );
and \U$14683 ( \14815 , \14651 , \14655 );
and \U$14684 ( \14816 , \14655 , \14660 );
and \U$14685 ( \14817 , \14651 , \14660 );
or \U$14686 ( \14818 , \14815 , \14816 , \14817 );
xor \U$14687 ( \14819 , \14814 , \14818 );
and \U$14688 ( \14820 , \14666 , \14670 );
and \U$14689 ( \14821 , \14670 , \14675 );
and \U$14690 ( \14822 , \14666 , \14675 );
or \U$14691 ( \14823 , \14820 , \14821 , \14822 );
xor \U$14692 ( \14824 , \14819 , \14823 );
and \U$14693 ( \14825 , \14682 , \14686 );
and \U$14694 ( \14826 , \14686 , \14691 );
and \U$14695 ( \14827 , \14682 , \14691 );
or \U$14696 ( \14828 , \14825 , \14826 , \14827 );
and \U$14697 ( \14829 , \14696 , \14700 );
and \U$14698 ( \14830 , \14700 , \14705 );
and \U$14699 ( \14831 , \14696 , \14705 );
or \U$14700 ( \14832 , \14829 , \14830 , \14831 );
xor \U$14701 ( \14833 , \14828 , \14832 );
and \U$14702 ( \14834 , \14708 , \14712 );
and \U$14703 ( \14835 , \14712 , \14717 );
and \U$14704 ( \14836 , \14708 , \14717 );
or \U$14705 ( \14837 , \14834 , \14835 , \14836 );
xor \U$14706 ( \14838 , \14833 , \14837 );
xor \U$14707 ( \14839 , \14824 , \14838 );
and \U$14708 ( \14840 , \14596 , \14600 );
and \U$14709 ( \14841 , \14600 , \14602 );
and \U$14710 ( \14842 , \14596 , \14602 );
or \U$14711 ( \14843 , \14840 , \14841 , \14842 );
and \U$14712 ( \14844 , \14607 , \14611 );
and \U$14713 ( \14845 , \14611 , \14616 );
and \U$14714 ( \14846 , \14607 , \14616 );
or \U$14715 ( \14847 , \14844 , \14845 , \14846 );
xor \U$14716 ( \14848 , \14843 , \14847 );
and \U$14717 ( \14849 , \14622 , \14626 );
and \U$14718 ( \14850 , \14626 , \14631 );
and \U$14719 ( \14851 , \14622 , \14631 );
or \U$14720 ( \14852 , \14849 , \14850 , \14851 );
xor \U$14721 ( \14853 , \14848 , \14852 );
xor \U$14722 ( \14854 , \14839 , \14853 );
xor \U$14723 ( \14855 , \14810 , \14854 );
and \U$14724 ( \14856 , \4160 , \4132 );
and \U$14725 ( \14857 , \4364 , \4012 );
nor \U$14726 ( \14858 , \14856 , \14857 );
xnor \U$14727 ( \14859 , \14858 , \3925 );
and \U$14728 ( \14860 , \3736 , \4581 );
and \U$14729 ( \14861 , \3912 , \4424 );
nor \U$14730 ( \14862 , \14860 , \14861 );
xnor \U$14731 ( \14863 , \14862 , \4377 );
xor \U$14732 ( \14864 , \14859 , \14863 );
and \U$14733 ( \14865 , \3395 , \5011 );
and \U$14734 ( \14866 , \3646 , \4878 );
nor \U$14735 ( \14867 , \14865 , \14866 );
xnor \U$14736 ( \14868 , \14867 , \4762 );
xor \U$14737 ( \14869 , \14864 , \14868 );
and \U$14738 ( \14870 , \3037 , \5485 );
and \U$14739 ( \14871 , \3143 , \5275 );
nor \U$14740 ( \14872 , \14870 , \14871 );
xnor \U$14741 ( \14873 , \14872 , \5169 );
and \U$14742 ( \14874 , \2757 , \5996 );
and \U$14743 ( \14875 , \2826 , \5695 );
nor \U$14744 ( \14876 , \14874 , \14875 );
xnor \U$14745 ( \14877 , \14876 , \5687 );
xor \U$14746 ( \14878 , \14873 , \14877 );
and \U$14747 ( \14879 , \2366 , \6401 );
and \U$14748 ( \14880 , \2521 , \6143 );
nor \U$14749 ( \14881 , \14879 , \14880 );
xnor \U$14750 ( \14882 , \14881 , \6148 );
xor \U$14751 ( \14883 , \14878 , \14882 );
xor \U$14752 ( \14884 , \14869 , \14883 );
and \U$14753 ( \14885 , \5469 , \3103 );
and \U$14754 ( \14886 , \5674 , \2934 );
nor \U$14755 ( \14887 , \14885 , \14886 );
xnor \U$14756 ( \14888 , \14887 , \2839 );
and \U$14757 ( \14889 , \4922 , \3357 );
and \U$14758 ( \14890 , \5156 , \3255 );
nor \U$14759 ( \14891 , \14889 , \14890 );
xnor \U$14760 ( \14892 , \14891 , \3156 );
xor \U$14761 ( \14893 , \14888 , \14892 );
and \U$14762 ( \14894 , \4654 , \3813 );
and \U$14763 ( \14895 , \4749 , \3557 );
nor \U$14764 ( \14896 , \14894 , \14895 );
xnor \U$14765 ( \14897 , \14896 , \3562 );
xor \U$14766 ( \14898 , \14893 , \14897 );
xor \U$14767 ( \14899 , \14884 , \14898 );
and \U$14768 ( \14900 , \6945 , \2121 );
and \U$14769 ( \14901 , \7231 , \2008 );
nor \U$14770 ( \14902 , \14900 , \14901 );
xnor \U$14771 ( \14903 , \14902 , \1961 );
and \U$14772 ( \14904 , \6514 , \2400 );
and \U$14773 ( \14905 , \6790 , \2246 );
nor \U$14774 ( \14906 , \14904 , \14905 );
xnor \U$14775 ( \14907 , \14906 , \2195 );
xor \U$14776 ( \14908 , \14903 , \14907 );
and \U$14777 ( \14909 , \6030 , \2669 );
and \U$14778 ( \14910 , \6281 , \2538 );
nor \U$14779 ( \14911 , \14909 , \14910 );
xnor \U$14780 ( \14912 , \14911 , \2534 );
xor \U$14781 ( \14913 , \14908 , \14912 );
and \U$14782 ( \14914 , \8652 , \1301 );
and \U$14783 ( \14915 , \8835 , \1246 );
nor \U$14784 ( \14916 , \14914 , \14915 );
xnor \U$14785 ( \14917 , \14916 , \1205 );
and \U$14786 ( \14918 , \8057 , \1578 );
and \U$14787 ( \14919 , \8349 , \1431 );
nor \U$14788 ( \14920 , \14918 , \14919 );
xnor \U$14789 ( \14921 , \14920 , \1436 );
xor \U$14790 ( \14922 , \14917 , \14921 );
and \U$14791 ( \14923 , \7556 , \1824 );
and \U$14792 ( \14924 , \7700 , \1739 );
nor \U$14793 ( \14925 , \14923 , \14924 );
xnor \U$14794 ( \14926 , \14925 , \1697 );
xor \U$14795 ( \14927 , \14922 , \14926 );
xor \U$14796 ( \14928 , \14913 , \14927 );
and \U$14797 ( \14929 , \10584 , \296 );
not \U$14798 ( \14930 , \14929 );
xnor \U$14799 ( \14931 , \14930 , \173 );
and \U$14800 ( \14932 , \9897 , \438 );
and \U$14801 ( \14933 , \10206 , \336 );
nor \U$14802 ( \14934 , \14932 , \14933 );
xnor \U$14803 ( \14935 , \14934 , \320 );
xor \U$14804 ( \14936 , \14931 , \14935 );
and \U$14805 ( \14937 , \9169 , \1086 );
and \U$14806 ( \14938 , \9465 , \508 );
nor \U$14807 ( \14939 , \14937 , \14938 );
xnor \U$14808 ( \14940 , \14939 , \487 );
xor \U$14809 ( \14941 , \14936 , \14940 );
xor \U$14810 ( \14942 , \14928 , \14941 );
xor \U$14811 ( \14943 , \14899 , \14942 );
and \U$14812 ( \14944 , \2090 , \7055 );
and \U$14813 ( \14945 , \2182 , \6675 );
nor \U$14814 ( \14946 , \14944 , \14945 );
xnor \U$14815 ( \14947 , \14946 , \6680 );
and \U$14816 ( \14948 , \1802 , \7489 );
and \U$14817 ( \14949 , \1948 , \7137 );
nor \U$14818 ( \14950 , \14948 , \14949 );
xnor \U$14819 ( \14951 , \14950 , \7142 );
xor \U$14820 ( \14952 , \14947 , \14951 );
and \U$14821 ( \14953 , \1601 , \8019 );
and \U$14822 ( \14954 , \1684 , \7830 );
nor \U$14823 ( \14955 , \14953 , \14954 );
xnor \U$14824 ( \14956 , \14955 , \7713 );
xor \U$14825 ( \14957 , \14952 , \14956 );
and \U$14826 ( \14958 , \1333 , \8540 );
and \U$14827 ( \14959 , \1484 , \8292 );
nor \U$14828 ( \14960 , \14958 , \14959 );
xnor \U$14829 ( \14961 , \14960 , \8297 );
and \U$14830 ( \14962 , \1147 , \9333 );
and \U$14831 ( \14963 , \1192 , \9006 );
nor \U$14832 ( \14964 , \14962 , \14963 );
xnor \U$14833 ( \14965 , \14964 , \8848 );
xor \U$14834 ( \14966 , \14961 , \14965 );
and \U$14835 ( \14967 , \412 , \9765 );
and \U$14836 ( \14968 , \474 , \9644 );
nor \U$14837 ( \14969 , \14967 , \14968 );
xnor \U$14838 ( \14970 , \14969 , \9478 );
xor \U$14839 ( \14971 , \14966 , \14970 );
xor \U$14840 ( \14972 , \14957 , \14971 );
and \U$14841 ( \14973 , \261 , \10408 );
and \U$14842 ( \14974 , \307 , \10116 );
nor \U$14843 ( \14975 , \14973 , \14974 );
xnor \U$14844 ( \14976 , \14975 , \10121 );
and \U$14845 ( \14977 , \185 , \10118 );
xnor \U$14846 ( \14978 , \14976 , \14977 );
xor \U$14847 ( \14979 , \14972 , \14978 );
xor \U$14848 ( \14980 , \14943 , \14979 );
xor \U$14849 ( \14981 , \14855 , \14980 );
xor \U$14850 ( \14982 , \14806 , \14981 );
and \U$14851 ( \14983 , \14551 , \14555 );
and \U$14852 ( \14984 , \14555 , \14560 );
and \U$14853 ( \14985 , \14551 , \14560 );
or \U$14854 ( \14986 , \14983 , \14984 , \14985 );
and \U$14855 ( \14987 , \14565 , \14569 );
and \U$14856 ( \14988 , \14569 , \14574 );
and \U$14857 ( \14989 , \14565 , \14574 );
or \U$14858 ( \14990 , \14987 , \14988 , \14989 );
xor \U$14859 ( \14991 , \14986 , \14990 );
and \U$14860 ( \14992 , \14580 , \14584 );
and \U$14861 ( \14993 , \14584 , \14589 );
and \U$14862 ( \14994 , \14580 , \14589 );
or \U$14863 ( \14995 , \14992 , \14993 , \14994 );
xor \U$14864 ( \14996 , \14991 , \14995 );
and \U$14865 ( \14997 , \14603 , \14617 );
and \U$14866 ( \14998 , \14617 , \14632 );
and \U$14867 ( \14999 , \14603 , \14632 );
or \U$14868 ( \15000 , \14997 , \14998 , \14999 );
and \U$14869 ( \15001 , \14647 , \14661 );
and \U$14870 ( \15002 , \14661 , \14676 );
and \U$14871 ( \15003 , \14647 , \14676 );
or \U$14872 ( \15004 , \15001 , \15002 , \15003 );
xor \U$14873 ( \15005 , \15000 , \15004 );
and \U$14874 ( \15006 , \14692 , \14706 );
and \U$14875 ( \15007 , \14706 , \14718 );
and \U$14876 ( \15008 , \14692 , \14718 );
or \U$14877 ( \15009 , \15006 , \15007 , \15008 );
xor \U$14878 ( \15010 , \15005 , \15009 );
xor \U$14879 ( \15011 , \14996 , \15010 );
xor \U$14880 ( \15012 , \14982 , \15011 );
xor \U$14881 ( \15013 , \14792 , \15012 );
xor \U$14882 ( \15014 , \14783 , \15013 );
xor \U$14883 ( \15015 , \14767 , \15014 );
and \U$14884 ( \15016 , \14501 , \14751 );
xor \U$14885 ( \15017 , \15015 , \15016 );
and \U$14886 ( \15018 , \14752 , \14756 );
and \U$14887 ( \15019 , \14757 , \14760 );
or \U$14888 ( \15020 , \15018 , \15019 );
xor \U$14889 ( \15021 , \15017 , \15020 );
buf \U$14890 ( \15022 , \15021 );
buf \U$14891 ( \15023 , \15022 );
and \U$14892 ( \15024 , \14771 , \14782 );
and \U$14893 ( \15025 , \14782 , \15013 );
and \U$14894 ( \15026 , \14771 , \15013 );
or \U$14895 ( \15027 , \15024 , \15025 , \15026 );
and \U$14896 ( \15028 , \14787 , \14791 );
and \U$14897 ( \15029 , \14791 , \15012 );
and \U$14898 ( \15030 , \14787 , \15012 );
or \U$14899 ( \15031 , \15028 , \15029 , \15030 );
and \U$14900 ( \15032 , \14796 , \14800 );
and \U$14901 ( \15033 , \14800 , \14805 );
and \U$14902 ( \15034 , \14796 , \14805 );
or \U$14903 ( \15035 , \15032 , \15033 , \15034 );
and \U$14904 ( \15036 , \14810 , \14854 );
and \U$14905 ( \15037 , \14854 , \14980 );
and \U$14906 ( \15038 , \14810 , \14980 );
or \U$14907 ( \15039 , \15036 , \15037 , \15038 );
xor \U$14908 ( \15040 , \15035 , \15039 );
and \U$14909 ( \15041 , \14996 , \15010 );
xor \U$14910 ( \15042 , \15040 , \15041 );
xor \U$14911 ( \15043 , \15031 , \15042 );
and \U$14912 ( \15044 , \14775 , \14779 );
and \U$14913 ( \15045 , \14779 , \14781 );
and \U$14914 ( \15046 , \14775 , \14781 );
or \U$14915 ( \15047 , \15044 , \15045 , \15046 );
and \U$14916 ( \15048 , \14806 , \14981 );
and \U$14917 ( \15049 , \14981 , \15011 );
and \U$14918 ( \15050 , \14806 , \15011 );
or \U$14919 ( \15051 , \15048 , \15049 , \15050 );
xor \U$14920 ( \15052 , \15047 , \15051 );
and \U$14921 ( \15053 , \14986 , \14990 );
and \U$14922 ( \15054 , \14990 , \14995 );
and \U$14923 ( \15055 , \14986 , \14995 );
or \U$14924 ( \15056 , \15053 , \15054 , \15055 );
and \U$14925 ( \15057 , \15000 , \15004 );
and \U$14926 ( \15058 , \15004 , \15009 );
and \U$14927 ( \15059 , \15000 , \15009 );
or \U$14928 ( \15060 , \15057 , \15058 , \15059 );
xor \U$14929 ( \15061 , \15056 , \15060 );
and \U$14930 ( \15062 , \14899 , \14942 );
and \U$14931 ( \15063 , \14942 , \14979 );
and \U$14932 ( \15064 , \14899 , \14979 );
or \U$14933 ( \15065 , \15062 , \15063 , \15064 );
xor \U$14934 ( \15066 , \15061 , \15065 );
and \U$14935 ( \15067 , \14824 , \14838 );
and \U$14936 ( \15068 , \14838 , \14853 );
and \U$14937 ( \15069 , \14824 , \14853 );
or \U$14938 ( \15070 , \15067 , \15068 , \15069 );
and \U$14939 ( \15071 , \14947 , \14951 );
and \U$14940 ( \15072 , \14951 , \14956 );
and \U$14941 ( \15073 , \14947 , \14956 );
or \U$14942 ( \15074 , \15071 , \15072 , \15073 );
and \U$14943 ( \15075 , \14961 , \14965 );
and \U$14944 ( \15076 , \14965 , \14970 );
and \U$14945 ( \15077 , \14961 , \14970 );
or \U$14946 ( \15078 , \15075 , \15076 , \15077 );
xor \U$14947 ( \15079 , \15074 , \15078 );
or \U$14948 ( \15080 , \14976 , \14977 );
xor \U$14949 ( \15081 , \15079 , \15080 );
and \U$14950 ( \15082 , \14903 , \14907 );
and \U$14951 ( \15083 , \14907 , \14912 );
and \U$14952 ( \15084 , \14903 , \14912 );
or \U$14953 ( \15085 , \15082 , \15083 , \15084 );
and \U$14954 ( \15086 , \14917 , \14921 );
and \U$14955 ( \15087 , \14921 , \14926 );
and \U$14956 ( \15088 , \14917 , \14926 );
or \U$14957 ( \15089 , \15086 , \15087 , \15088 );
xor \U$14958 ( \15090 , \15085 , \15089 );
and \U$14959 ( \15091 , \14931 , \14935 );
and \U$14960 ( \15092 , \14935 , \14940 );
and \U$14961 ( \15093 , \14931 , \14940 );
or \U$14962 ( \15094 , \15091 , \15092 , \15093 );
xor \U$14963 ( \15095 , \15090 , \15094 );
xor \U$14964 ( \15096 , \15081 , \15095 );
and \U$14965 ( \15097 , \14859 , \14863 );
and \U$14966 ( \15098 , \14863 , \14868 );
and \U$14967 ( \15099 , \14859 , \14868 );
or \U$14968 ( \15100 , \15097 , \15098 , \15099 );
and \U$14969 ( \15101 , \14873 , \14877 );
and \U$14970 ( \15102 , \14877 , \14882 );
and \U$14971 ( \15103 , \14873 , \14882 );
or \U$14972 ( \15104 , \15101 , \15102 , \15103 );
xor \U$14973 ( \15105 , \15100 , \15104 );
and \U$14974 ( \15106 , \14888 , \14892 );
and \U$14975 ( \15107 , \14892 , \14897 );
and \U$14976 ( \15108 , \14888 , \14897 );
or \U$14977 ( \15109 , \15106 , \15107 , \15108 );
xor \U$14978 ( \15110 , \15105 , \15109 );
xor \U$14979 ( \15111 , \15096 , \15110 );
xor \U$14980 ( \15112 , \15070 , \15111 );
and \U$14981 ( \15113 , \5674 , \3103 );
and \U$14982 ( \15114 , \6030 , \2934 );
nor \U$14983 ( \15115 , \15113 , \15114 );
xnor \U$14984 ( \15116 , \15115 , \2839 );
and \U$14985 ( \15117 , \5156 , \3357 );
and \U$14986 ( \15118 , \5469 , \3255 );
nor \U$14987 ( \15119 , \15117 , \15118 );
xnor \U$14988 ( \15120 , \15119 , \3156 );
xor \U$14989 ( \15121 , \15116 , \15120 );
and \U$14990 ( \15122 , \4749 , \3813 );
and \U$14991 ( \15123 , \4922 , \3557 );
nor \U$14992 ( \15124 , \15122 , \15123 );
xnor \U$14993 ( \15125 , \15124 , \3562 );
xor \U$14994 ( \15126 , \15121 , \15125 );
and \U$14995 ( \15127 , \4364 , \4132 );
and \U$14996 ( \15128 , \4654 , \4012 );
nor \U$14997 ( \15129 , \15127 , \15128 );
xnor \U$14998 ( \15130 , \15129 , \3925 );
and \U$14999 ( \15131 , \3912 , \4581 );
and \U$15000 ( \15132 , \4160 , \4424 );
nor \U$15001 ( \15133 , \15131 , \15132 );
xnor \U$15002 ( \15134 , \15133 , \4377 );
xor \U$15003 ( \15135 , \15130 , \15134 );
and \U$15004 ( \15136 , \3646 , \5011 );
and \U$15005 ( \15137 , \3736 , \4878 );
nor \U$15006 ( \15138 , \15136 , \15137 );
xnor \U$15007 ( \15139 , \15138 , \4762 );
xor \U$15008 ( \15140 , \15135 , \15139 );
xor \U$15009 ( \15141 , \15126 , \15140 );
and \U$15010 ( \15142 , \3143 , \5485 );
and \U$15011 ( \15143 , \3395 , \5275 );
nor \U$15012 ( \15144 , \15142 , \15143 );
xnor \U$15013 ( \15145 , \15144 , \5169 );
and \U$15014 ( \15146 , \2826 , \5996 );
and \U$15015 ( \15147 , \3037 , \5695 );
nor \U$15016 ( \15148 , \15146 , \15147 );
xnor \U$15017 ( \15149 , \15148 , \5687 );
xor \U$15018 ( \15150 , \15145 , \15149 );
and \U$15019 ( \15151 , \2521 , \6401 );
and \U$15020 ( \15152 , \2757 , \6143 );
nor \U$15021 ( \15153 , \15151 , \15152 );
xnor \U$15022 ( \15154 , \15153 , \6148 );
xor \U$15023 ( \15155 , \15150 , \15154 );
xor \U$15024 ( \15156 , \15141 , \15155 );
and \U$15025 ( \15157 , \8835 , \1301 );
and \U$15026 ( \15158 , \9169 , \1246 );
nor \U$15027 ( \15159 , \15157 , \15158 );
xnor \U$15028 ( \15160 , \15159 , \1205 );
and \U$15029 ( \15161 , \8349 , \1578 );
and \U$15030 ( \15162 , \8652 , \1431 );
nor \U$15031 ( \15163 , \15161 , \15162 );
xnor \U$15032 ( \15164 , \15163 , \1436 );
xor \U$15033 ( \15165 , \15160 , \15164 );
and \U$15034 ( \15166 , \7700 , \1824 );
and \U$15035 ( \15167 , \8057 , \1739 );
nor \U$15036 ( \15168 , \15166 , \15167 );
xnor \U$15037 ( \15169 , \15168 , \1697 );
xor \U$15038 ( \15170 , \15165 , \15169 );
not \U$15039 ( \15171 , \173 );
and \U$15040 ( \15172 , \10206 , \438 );
and \U$15041 ( \15173 , \10584 , \336 );
nor \U$15042 ( \15174 , \15172 , \15173 );
xnor \U$15043 ( \15175 , \15174 , \320 );
xor \U$15044 ( \15176 , \15171 , \15175 );
and \U$15045 ( \15177 , \9465 , \1086 );
and \U$15046 ( \15178 , \9897 , \508 );
nor \U$15047 ( \15179 , \15177 , \15178 );
xnor \U$15048 ( \15180 , \15179 , \487 );
xor \U$15049 ( \15181 , \15176 , \15180 );
xor \U$15050 ( \15182 , \15170 , \15181 );
and \U$15051 ( \15183 , \7231 , \2121 );
and \U$15052 ( \15184 , \7556 , \2008 );
nor \U$15053 ( \15185 , \15183 , \15184 );
xnor \U$15054 ( \15186 , \15185 , \1961 );
and \U$15055 ( \15187 , \6790 , \2400 );
and \U$15056 ( \15188 , \6945 , \2246 );
nor \U$15057 ( \15189 , \15187 , \15188 );
xnor \U$15058 ( \15190 , \15189 , \2195 );
xor \U$15059 ( \15191 , \15186 , \15190 );
and \U$15060 ( \15192 , \6281 , \2669 );
and \U$15061 ( \15193 , \6514 , \2538 );
nor \U$15062 ( \15194 , \15192 , \15193 );
xnor \U$15063 ( \15195 , \15194 , \2534 );
xor \U$15064 ( \15196 , \15191 , \15195 );
xor \U$15065 ( \15197 , \15182 , \15196 );
xor \U$15066 ( \15198 , \15156 , \15197 );
and \U$15067 ( \15199 , \2182 , \7055 );
and \U$15068 ( \15200 , \2366 , \6675 );
nor \U$15069 ( \15201 , \15199 , \15200 );
xnor \U$15070 ( \15202 , \15201 , \6680 );
and \U$15071 ( \15203 , \1948 , \7489 );
and \U$15072 ( \15204 , \2090 , \7137 );
nor \U$15073 ( \15205 , \15203 , \15204 );
xnor \U$15074 ( \15206 , \15205 , \7142 );
xor \U$15075 ( \15207 , \15202 , \15206 );
and \U$15076 ( \15208 , \1684 , \8019 );
and \U$15077 ( \15209 , \1802 , \7830 );
nor \U$15078 ( \15210 , \15208 , \15209 );
xnor \U$15079 ( \15211 , \15210 , \7713 );
xor \U$15080 ( \15212 , \15207 , \15211 );
and \U$15081 ( \15213 , \1484 , \8540 );
and \U$15082 ( \15214 , \1601 , \8292 );
nor \U$15083 ( \15215 , \15213 , \15214 );
xnor \U$15084 ( \15216 , \15215 , \8297 );
and \U$15085 ( \15217 , \1192 , \9333 );
and \U$15086 ( \15218 , \1333 , \9006 );
nor \U$15087 ( \15219 , \15217 , \15218 );
xnor \U$15088 ( \15220 , \15219 , \8848 );
xor \U$15089 ( \15221 , \15216 , \15220 );
and \U$15090 ( \15222 , \474 , \9765 );
and \U$15091 ( \15223 , \1147 , \9644 );
nor \U$15092 ( \15224 , \15222 , \15223 );
xnor \U$15093 ( \15225 , \15224 , \9478 );
xor \U$15094 ( \15226 , \15221 , \15225 );
xor \U$15095 ( \15227 , \15212 , \15226 );
and \U$15096 ( \15228 , \307 , \10408 );
and \U$15097 ( \15229 , \412 , \10116 );
nor \U$15098 ( \15230 , \15228 , \15229 );
xnor \U$15099 ( \15231 , \15230 , \10121 );
and \U$15100 ( \15232 , \261 , \10118 );
xor \U$15101 ( \15233 , \15231 , \15232 );
xor \U$15102 ( \15234 , \15227 , \15233 );
xor \U$15103 ( \15235 , \15198 , \15234 );
xor \U$15104 ( \15236 , \15112 , \15235 );
xor \U$15105 ( \15237 , \15066 , \15236 );
and \U$15106 ( \15238 , \14814 , \14818 );
and \U$15107 ( \15239 , \14818 , \14823 );
and \U$15108 ( \15240 , \14814 , \14823 );
or \U$15109 ( \15241 , \15238 , \15239 , \15240 );
and \U$15110 ( \15242 , \14828 , \14832 );
and \U$15111 ( \15243 , \14832 , \14837 );
and \U$15112 ( \15244 , \14828 , \14837 );
or \U$15113 ( \15245 , \15242 , \15243 , \15244 );
xor \U$15114 ( \15246 , \15241 , \15245 );
and \U$15115 ( \15247 , \14843 , \14847 );
and \U$15116 ( \15248 , \14847 , \14852 );
and \U$15117 ( \15249 , \14843 , \14852 );
or \U$15118 ( \15250 , \15247 , \15248 , \15249 );
xor \U$15119 ( \15251 , \15246 , \15250 );
and \U$15120 ( \15252 , \14869 , \14883 );
and \U$15121 ( \15253 , \14883 , \14898 );
and \U$15122 ( \15254 , \14869 , \14898 );
or \U$15123 ( \15255 , \15252 , \15253 , \15254 );
and \U$15124 ( \15256 , \14913 , \14927 );
and \U$15125 ( \15257 , \14927 , \14941 );
and \U$15126 ( \15258 , \14913 , \14941 );
or \U$15127 ( \15259 , \15256 , \15257 , \15258 );
xor \U$15128 ( \15260 , \15255 , \15259 );
and \U$15129 ( \15261 , \14957 , \14971 );
and \U$15130 ( \15262 , \14971 , \14978 );
and \U$15131 ( \15263 , \14957 , \14978 );
or \U$15132 ( \15264 , \15261 , \15262 , \15263 );
xor \U$15133 ( \15265 , \15260 , \15264 );
xor \U$15134 ( \15266 , \15251 , \15265 );
xor \U$15135 ( \15267 , \15237 , \15266 );
xor \U$15136 ( \15268 , \15052 , \15267 );
xor \U$15137 ( \15269 , \15043 , \15268 );
xor \U$15138 ( \15270 , \15027 , \15269 );
and \U$15139 ( \15271 , \14767 , \15014 );
xor \U$15140 ( \15272 , \15270 , \15271 );
and \U$15141 ( \15273 , \15015 , \15016 );
and \U$15142 ( \15274 , \15017 , \15020 );
or \U$15143 ( \15275 , \15273 , \15274 );
xor \U$15144 ( \15276 , \15272 , \15275 );
buf \U$15145 ( \15277 , \15276 );
buf \U$15146 ( \15278 , \15277 );
and \U$15147 ( \15279 , \15031 , \15042 );
and \U$15148 ( \15280 , \15042 , \15268 );
and \U$15149 ( \15281 , \15031 , \15268 );
or \U$15150 ( \15282 , \15279 , \15280 , \15281 );
and \U$15151 ( \15283 , \15047 , \15051 );
and \U$15152 ( \15284 , \15051 , \15267 );
and \U$15153 ( \15285 , \15047 , \15267 );
or \U$15154 ( \15286 , \15283 , \15284 , \15285 );
and \U$15155 ( \15287 , \15056 , \15060 );
and \U$15156 ( \15288 , \15060 , \15065 );
and \U$15157 ( \15289 , \15056 , \15065 );
or \U$15158 ( \15290 , \15287 , \15288 , \15289 );
and \U$15159 ( \15291 , \15070 , \15111 );
and \U$15160 ( \15292 , \15111 , \15235 );
and \U$15161 ( \15293 , \15070 , \15235 );
or \U$15162 ( \15294 , \15291 , \15292 , \15293 );
xor \U$15163 ( \15295 , \15290 , \15294 );
and \U$15164 ( \15296 , \15251 , \15265 );
xor \U$15165 ( \15297 , \15295 , \15296 );
xor \U$15166 ( \15298 , \15286 , \15297 );
and \U$15167 ( \15299 , \15035 , \15039 );
and \U$15168 ( \15300 , \15039 , \15041 );
and \U$15169 ( \15301 , \15035 , \15041 );
or \U$15170 ( \15302 , \15299 , \15300 , \15301 );
and \U$15171 ( \15303 , \15066 , \15236 );
and \U$15172 ( \15304 , \15236 , \15266 );
and \U$15173 ( \15305 , \15066 , \15266 );
or \U$15174 ( \15306 , \15303 , \15304 , \15305 );
xor \U$15175 ( \15307 , \15302 , \15306 );
and \U$15176 ( \15308 , \15241 , \15245 );
and \U$15177 ( \15309 , \15245 , \15250 );
and \U$15178 ( \15310 , \15241 , \15250 );
or \U$15179 ( \15311 , \15308 , \15309 , \15310 );
and \U$15180 ( \15312 , \15255 , \15259 );
and \U$15181 ( \15313 , \15259 , \15264 );
and \U$15182 ( \15314 , \15255 , \15264 );
or \U$15183 ( \15315 , \15312 , \15313 , \15314 );
xor \U$15184 ( \15316 , \15311 , \15315 );
and \U$15185 ( \15317 , \15156 , \15197 );
and \U$15186 ( \15318 , \15197 , \15234 );
and \U$15187 ( \15319 , \15156 , \15234 );
or \U$15188 ( \15320 , \15317 , \15318 , \15319 );
xor \U$15189 ( \15321 , \15316 , \15320 );
and \U$15190 ( \15322 , \15081 , \15095 );
and \U$15191 ( \15323 , \15095 , \15110 );
and \U$15192 ( \15324 , \15081 , \15110 );
or \U$15193 ( \15325 , \15322 , \15323 , \15324 );
and \U$15194 ( \15326 , \15160 , \15164 );
and \U$15195 ( \15327 , \15164 , \15169 );
and \U$15196 ( \15328 , \15160 , \15169 );
or \U$15197 ( \15329 , \15326 , \15327 , \15328 );
and \U$15198 ( \15330 , \15171 , \15175 );
and \U$15199 ( \15331 , \15175 , \15180 );
and \U$15200 ( \15332 , \15171 , \15180 );
or \U$15201 ( \15333 , \15330 , \15331 , \15332 );
xor \U$15202 ( \15334 , \15329 , \15333 );
and \U$15203 ( \15335 , \15186 , \15190 );
and \U$15204 ( \15336 , \15190 , \15195 );
and \U$15205 ( \15337 , \15186 , \15195 );
or \U$15206 ( \15338 , \15335 , \15336 , \15337 );
xor \U$15207 ( \15339 , \15334 , \15338 );
and \U$15208 ( \15340 , \15202 , \15206 );
and \U$15209 ( \15341 , \15206 , \15211 );
and \U$15210 ( \15342 , \15202 , \15211 );
or \U$15211 ( \15343 , \15340 , \15341 , \15342 );
and \U$15212 ( \15344 , \15216 , \15220 );
and \U$15213 ( \15345 , \15220 , \15225 );
and \U$15214 ( \15346 , \15216 , \15225 );
or \U$15215 ( \15347 , \15344 , \15345 , \15346 );
xor \U$15216 ( \15348 , \15343 , \15347 );
and \U$15217 ( \15349 , \15231 , \15232 );
xor \U$15218 ( \15350 , \15348 , \15349 );
xor \U$15219 ( \15351 , \15339 , \15350 );
and \U$15220 ( \15352 , \15116 , \15120 );
and \U$15221 ( \15353 , \15120 , \15125 );
and \U$15222 ( \15354 , \15116 , \15125 );
or \U$15223 ( \15355 , \15352 , \15353 , \15354 );
and \U$15224 ( \15356 , \15130 , \15134 );
and \U$15225 ( \15357 , \15134 , \15139 );
and \U$15226 ( \15358 , \15130 , \15139 );
or \U$15227 ( \15359 , \15356 , \15357 , \15358 );
xor \U$15228 ( \15360 , \15355 , \15359 );
and \U$15229 ( \15361 , \15145 , \15149 );
and \U$15230 ( \15362 , \15149 , \15154 );
and \U$15231 ( \15363 , \15145 , \15154 );
or \U$15232 ( \15364 , \15361 , \15362 , \15363 );
xor \U$15233 ( \15365 , \15360 , \15364 );
xor \U$15234 ( \15366 , \15351 , \15365 );
xor \U$15235 ( \15367 , \15325 , \15366 );
and \U$15236 ( \15368 , \4160 , \4581 );
and \U$15237 ( \15369 , \4364 , \4424 );
nor \U$15238 ( \15370 , \15368 , \15369 );
xnor \U$15239 ( \15371 , \15370 , \4377 );
and \U$15240 ( \15372 , \3736 , \5011 );
and \U$15241 ( \15373 , \3912 , \4878 );
nor \U$15242 ( \15374 , \15372 , \15373 );
xnor \U$15243 ( \15375 , \15374 , \4762 );
xor \U$15244 ( \15376 , \15371 , \15375 );
and \U$15245 ( \15377 , \3395 , \5485 );
and \U$15246 ( \15378 , \3646 , \5275 );
nor \U$15247 ( \15379 , \15377 , \15378 );
xnor \U$15248 ( \15380 , \15379 , \5169 );
xor \U$15249 ( \15381 , \15376 , \15380 );
and \U$15250 ( \15382 , \5469 , \3357 );
and \U$15251 ( \15383 , \5674 , \3255 );
nor \U$15252 ( \15384 , \15382 , \15383 );
xnor \U$15253 ( \15385 , \15384 , \3156 );
and \U$15254 ( \15386 , \4922 , \3813 );
and \U$15255 ( \15387 , \5156 , \3557 );
nor \U$15256 ( \15388 , \15386 , \15387 );
xnor \U$15257 ( \15389 , \15388 , \3562 );
xor \U$15258 ( \15390 , \15385 , \15389 );
and \U$15259 ( \15391 , \4654 , \4132 );
and \U$15260 ( \15392 , \4749 , \4012 );
nor \U$15261 ( \15393 , \15391 , \15392 );
xnor \U$15262 ( \15394 , \15393 , \3925 );
xor \U$15263 ( \15395 , \15390 , \15394 );
xor \U$15264 ( \15396 , \15381 , \15395 );
and \U$15265 ( \15397 , \3037 , \5996 );
and \U$15266 ( \15398 , \3143 , \5695 );
nor \U$15267 ( \15399 , \15397 , \15398 );
xnor \U$15268 ( \15400 , \15399 , \5687 );
and \U$15269 ( \15401 , \2757 , \6401 );
and \U$15270 ( \15402 , \2826 , \6143 );
nor \U$15271 ( \15403 , \15401 , \15402 );
xnor \U$15272 ( \15404 , \15403 , \6148 );
xor \U$15273 ( \15405 , \15400 , \15404 );
and \U$15274 ( \15406 , \2366 , \7055 );
and \U$15275 ( \15407 , \2521 , \6675 );
nor \U$15276 ( \15408 , \15406 , \15407 );
xnor \U$15277 ( \15409 , \15408 , \6680 );
xor \U$15278 ( \15410 , \15405 , \15409 );
xor \U$15279 ( \15411 , \15396 , \15410 );
and \U$15280 ( \15412 , \8652 , \1578 );
and \U$15281 ( \15413 , \8835 , \1431 );
nor \U$15282 ( \15414 , \15412 , \15413 );
xnor \U$15283 ( \15415 , \15414 , \1436 );
and \U$15284 ( \15416 , \8057 , \1824 );
and \U$15285 ( \15417 , \8349 , \1739 );
nor \U$15286 ( \15418 , \15416 , \15417 );
xnor \U$15287 ( \15419 , \15418 , \1697 );
xor \U$15288 ( \15420 , \15415 , \15419 );
and \U$15289 ( \15421 , \7556 , \2121 );
and \U$15290 ( \15422 , \7700 , \2008 );
nor \U$15291 ( \15423 , \15421 , \15422 );
xnor \U$15292 ( \15424 , \15423 , \1961 );
xor \U$15293 ( \15425 , \15420 , \15424 );
and \U$15294 ( \15426 , \10584 , \438 );
not \U$15295 ( \15427 , \15426 );
xnor \U$15296 ( \15428 , \15427 , \320 );
and \U$15297 ( \15429 , \9897 , \1086 );
and \U$15298 ( \15430 , \10206 , \508 );
nor \U$15299 ( \15431 , \15429 , \15430 );
xnor \U$15300 ( \15432 , \15431 , \487 );
xor \U$15301 ( \15433 , \15428 , \15432 );
and \U$15302 ( \15434 , \9169 , \1301 );
and \U$15303 ( \15435 , \9465 , \1246 );
nor \U$15304 ( \15436 , \15434 , \15435 );
xnor \U$15305 ( \15437 , \15436 , \1205 );
xor \U$15306 ( \15438 , \15433 , \15437 );
xor \U$15307 ( \15439 , \15425 , \15438 );
and \U$15308 ( \15440 , \6945 , \2400 );
and \U$15309 ( \15441 , \7231 , \2246 );
nor \U$15310 ( \15442 , \15440 , \15441 );
xnor \U$15311 ( \15443 , \15442 , \2195 );
and \U$15312 ( \15444 , \6514 , \2669 );
and \U$15313 ( \15445 , \6790 , \2538 );
nor \U$15314 ( \15446 , \15444 , \15445 );
xnor \U$15315 ( \15447 , \15446 , \2534 );
xor \U$15316 ( \15448 , \15443 , \15447 );
and \U$15317 ( \15449 , \6030 , \3103 );
and \U$15318 ( \15450 , \6281 , \2934 );
nor \U$15319 ( \15451 , \15449 , \15450 );
xnor \U$15320 ( \15452 , \15451 , \2839 );
xor \U$15321 ( \15453 , \15448 , \15452 );
xor \U$15322 ( \15454 , \15439 , \15453 );
xor \U$15323 ( \15455 , \15411 , \15454 );
and \U$15324 ( \15456 , \2090 , \7489 );
and \U$15325 ( \15457 , \2182 , \7137 );
nor \U$15326 ( \15458 , \15456 , \15457 );
xnor \U$15327 ( \15459 , \15458 , \7142 );
and \U$15328 ( \15460 , \1802 , \8019 );
and \U$15329 ( \15461 , \1948 , \7830 );
nor \U$15330 ( \15462 , \15460 , \15461 );
xnor \U$15331 ( \15463 , \15462 , \7713 );
xor \U$15332 ( \15464 , \15459 , \15463 );
and \U$15333 ( \15465 , \1601 , \8540 );
and \U$15334 ( \15466 , \1684 , \8292 );
nor \U$15335 ( \15467 , \15465 , \15466 );
xnor \U$15336 ( \15468 , \15467 , \8297 );
xor \U$15337 ( \15469 , \15464 , \15468 );
and \U$15338 ( \15470 , \1333 , \9333 );
and \U$15339 ( \15471 , \1484 , \9006 );
nor \U$15340 ( \15472 , \15470 , \15471 );
xnor \U$15341 ( \15473 , \15472 , \8848 );
and \U$15342 ( \15474 , \1147 , \9765 );
and \U$15343 ( \15475 , \1192 , \9644 );
nor \U$15344 ( \15476 , \15474 , \15475 );
xnor \U$15345 ( \15477 , \15476 , \9478 );
xor \U$15346 ( \15478 , \15473 , \15477 );
and \U$15347 ( \15479 , \412 , \10408 );
and \U$15348 ( \15480 , \474 , \10116 );
nor \U$15349 ( \15481 , \15479 , \15480 );
xnor \U$15350 ( \15482 , \15481 , \10121 );
xor \U$15351 ( \15483 , \15478 , \15482 );
xor \U$15352 ( \15484 , \15469 , \15483 );
and \U$15353 ( \15485 , \307 , \10118 );
not \U$15354 ( \15486 , \15485 );
xor \U$15355 ( \15487 , \15484 , \15486 );
xor \U$15356 ( \15488 , \15455 , \15487 );
xor \U$15357 ( \15489 , \15367 , \15488 );
xor \U$15358 ( \15490 , \15321 , \15489 );
and \U$15359 ( \15491 , \15126 , \15140 );
and \U$15360 ( \15492 , \15140 , \15155 );
and \U$15361 ( \15493 , \15126 , \15155 );
or \U$15362 ( \15494 , \15491 , \15492 , \15493 );
and \U$15363 ( \15495 , \15170 , \15181 );
and \U$15364 ( \15496 , \15181 , \15196 );
and \U$15365 ( \15497 , \15170 , \15196 );
or \U$15366 ( \15498 , \15495 , \15496 , \15497 );
xor \U$15367 ( \15499 , \15494 , \15498 );
and \U$15368 ( \15500 , \15212 , \15226 );
and \U$15369 ( \15501 , \15226 , \15233 );
and \U$15370 ( \15502 , \15212 , \15233 );
or \U$15371 ( \15503 , \15500 , \15501 , \15502 );
xor \U$15372 ( \15504 , \15499 , \15503 );
and \U$15373 ( \15505 , \15074 , \15078 );
and \U$15374 ( \15506 , \15078 , \15080 );
and \U$15375 ( \15507 , \15074 , \15080 );
or \U$15376 ( \15508 , \15505 , \15506 , \15507 );
and \U$15377 ( \15509 , \15085 , \15089 );
and \U$15378 ( \15510 , \15089 , \15094 );
and \U$15379 ( \15511 , \15085 , \15094 );
or \U$15380 ( \15512 , \15509 , \15510 , \15511 );
xor \U$15381 ( \15513 , \15508 , \15512 );
and \U$15382 ( \15514 , \15100 , \15104 );
and \U$15383 ( \15515 , \15104 , \15109 );
and \U$15384 ( \15516 , \15100 , \15109 );
or \U$15385 ( \15517 , \15514 , \15515 , \15516 );
xor \U$15386 ( \15518 , \15513 , \15517 );
xor \U$15387 ( \15519 , \15504 , \15518 );
xor \U$15388 ( \15520 , \15490 , \15519 );
xor \U$15389 ( \15521 , \15307 , \15520 );
xor \U$15390 ( \15522 , \15298 , \15521 );
xor \U$15391 ( \15523 , \15282 , \15522 );
and \U$15392 ( \15524 , \15027 , \15269 );
xor \U$15393 ( \15525 , \15523 , \15524 );
and \U$15394 ( \15526 , \15270 , \15271 );
and \U$15395 ( \15527 , \15272 , \15275 );
or \U$15396 ( \15528 , \15526 , \15527 );
xor \U$15397 ( \15529 , \15525 , \15528 );
buf \U$15398 ( \15530 , \15529 );
buf \U$15399 ( \15531 , \15530 );
and \U$15400 ( \15532 , \15286 , \15297 );
and \U$15401 ( \15533 , \15297 , \15521 );
and \U$15402 ( \15534 , \15286 , \15521 );
or \U$15403 ( \15535 , \15532 , \15533 , \15534 );
and \U$15404 ( \15536 , \15302 , \15306 );
and \U$15405 ( \15537 , \15306 , \15520 );
and \U$15406 ( \15538 , \15302 , \15520 );
or \U$15407 ( \15539 , \15536 , \15537 , \15538 );
and \U$15408 ( \15540 , \15311 , \15315 );
and \U$15409 ( \15541 , \15315 , \15320 );
and \U$15410 ( \15542 , \15311 , \15320 );
or \U$15411 ( \15543 , \15540 , \15541 , \15542 );
and \U$15412 ( \15544 , \15325 , \15366 );
and \U$15413 ( \15545 , \15366 , \15488 );
and \U$15414 ( \15546 , \15325 , \15488 );
or \U$15415 ( \15547 , \15544 , \15545 , \15546 );
xor \U$15416 ( \15548 , \15543 , \15547 );
and \U$15417 ( \15549 , \15504 , \15518 );
xor \U$15418 ( \15550 , \15548 , \15549 );
xor \U$15419 ( \15551 , \15539 , \15550 );
and \U$15420 ( \15552 , \15290 , \15294 );
and \U$15421 ( \15553 , \15294 , \15296 );
and \U$15422 ( \15554 , \15290 , \15296 );
or \U$15423 ( \15555 , \15552 , \15553 , \15554 );
and \U$15424 ( \15556 , \15321 , \15489 );
and \U$15425 ( \15557 , \15489 , \15519 );
and \U$15426 ( \15558 , \15321 , \15519 );
or \U$15427 ( \15559 , \15556 , \15557 , \15558 );
xor \U$15428 ( \15560 , \15555 , \15559 );
and \U$15429 ( \15561 , \15494 , \15498 );
and \U$15430 ( \15562 , \15498 , \15503 );
and \U$15431 ( \15563 , \15494 , \15503 );
or \U$15432 ( \15564 , \15561 , \15562 , \15563 );
and \U$15433 ( \15565 , \15508 , \15512 );
and \U$15434 ( \15566 , \15512 , \15517 );
and \U$15435 ( \15567 , \15508 , \15517 );
or \U$15436 ( \15568 , \15565 , \15566 , \15567 );
xor \U$15437 ( \15569 , \15564 , \15568 );
and \U$15438 ( \15570 , \15411 , \15454 );
and \U$15439 ( \15571 , \15454 , \15487 );
and \U$15440 ( \15572 , \15411 , \15487 );
or \U$15441 ( \15573 , \15570 , \15571 , \15572 );
xor \U$15442 ( \15574 , \15569 , \15573 );
and \U$15443 ( \15575 , \15339 , \15350 );
and \U$15444 ( \15576 , \15350 , \15365 );
and \U$15445 ( \15577 , \15339 , \15365 );
or \U$15446 ( \15578 , \15575 , \15576 , \15577 );
and \U$15447 ( \15579 , \15459 , \15463 );
and \U$15448 ( \15580 , \15463 , \15468 );
and \U$15449 ( \15581 , \15459 , \15468 );
or \U$15450 ( \15582 , \15579 , \15580 , \15581 );
and \U$15451 ( \15583 , \15473 , \15477 );
and \U$15452 ( \15584 , \15477 , \15482 );
and \U$15453 ( \15585 , \15473 , \15482 );
or \U$15454 ( \15586 , \15583 , \15584 , \15585 );
xor \U$15455 ( \15587 , \15582 , \15586 );
buf \U$15456 ( \15588 , \15485 );
xor \U$15457 ( \15589 , \15587 , \15588 );
and \U$15458 ( \15590 , \15371 , \15375 );
and \U$15459 ( \15591 , \15375 , \15380 );
and \U$15460 ( \15592 , \15371 , \15380 );
or \U$15461 ( \15593 , \15590 , \15591 , \15592 );
and \U$15462 ( \15594 , \15385 , \15389 );
and \U$15463 ( \15595 , \15389 , \15394 );
and \U$15464 ( \15596 , \15385 , \15394 );
or \U$15465 ( \15597 , \15594 , \15595 , \15596 );
xor \U$15466 ( \15598 , \15593 , \15597 );
and \U$15467 ( \15599 , \15400 , \15404 );
and \U$15468 ( \15600 , \15404 , \15409 );
and \U$15469 ( \15601 , \15400 , \15409 );
or \U$15470 ( \15602 , \15599 , \15600 , \15601 );
xor \U$15471 ( \15603 , \15598 , \15602 );
xor \U$15472 ( \15604 , \15589 , \15603 );
and \U$15473 ( \15605 , \15415 , \15419 );
and \U$15474 ( \15606 , \15419 , \15424 );
and \U$15475 ( \15607 , \15415 , \15424 );
or \U$15476 ( \15608 , \15605 , \15606 , \15607 );
and \U$15477 ( \15609 , \15428 , \15432 );
and \U$15478 ( \15610 , \15432 , \15437 );
and \U$15479 ( \15611 , \15428 , \15437 );
or \U$15480 ( \15612 , \15609 , \15610 , \15611 );
xor \U$15481 ( \15613 , \15608 , \15612 );
and \U$15482 ( \15614 , \15443 , \15447 );
and \U$15483 ( \15615 , \15447 , \15452 );
and \U$15484 ( \15616 , \15443 , \15452 );
or \U$15485 ( \15617 , \15614 , \15615 , \15616 );
xor \U$15486 ( \15618 , \15613 , \15617 );
xor \U$15487 ( \15619 , \15604 , \15618 );
xor \U$15488 ( \15620 , \15578 , \15619 );
and \U$15489 ( \15621 , \8835 , \1578 );
and \U$15490 ( \15622 , \9169 , \1431 );
nor \U$15491 ( \15623 , \15621 , \15622 );
xnor \U$15492 ( \15624 , \15623 , \1436 );
and \U$15493 ( \15625 , \8349 , \1824 );
and \U$15494 ( \15626 , \8652 , \1739 );
nor \U$15495 ( \15627 , \15625 , \15626 );
xnor \U$15496 ( \15628 , \15627 , \1697 );
xor \U$15497 ( \15629 , \15624 , \15628 );
and \U$15498 ( \15630 , \7700 , \2121 );
and \U$15499 ( \15631 , \8057 , \2008 );
nor \U$15500 ( \15632 , \15630 , \15631 );
xnor \U$15501 ( \15633 , \15632 , \1961 );
xor \U$15502 ( \15634 , \15629 , \15633 );
not \U$15503 ( \15635 , \320 );
and \U$15504 ( \15636 , \10206 , \1086 );
and \U$15505 ( \15637 , \10584 , \508 );
nor \U$15506 ( \15638 , \15636 , \15637 );
xnor \U$15507 ( \15639 , \15638 , \487 );
xor \U$15508 ( \15640 , \15635 , \15639 );
and \U$15509 ( \15641 , \9465 , \1301 );
and \U$15510 ( \15642 , \9897 , \1246 );
nor \U$15511 ( \15643 , \15641 , \15642 );
xnor \U$15512 ( \15644 , \15643 , \1205 );
xor \U$15513 ( \15645 , \15640 , \15644 );
xor \U$15514 ( \15646 , \15634 , \15645 );
and \U$15515 ( \15647 , \7231 , \2400 );
and \U$15516 ( \15648 , \7556 , \2246 );
nor \U$15517 ( \15649 , \15647 , \15648 );
xnor \U$15518 ( \15650 , \15649 , \2195 );
and \U$15519 ( \15651 , \6790 , \2669 );
and \U$15520 ( \15652 , \6945 , \2538 );
nor \U$15521 ( \15653 , \15651 , \15652 );
xnor \U$15522 ( \15654 , \15653 , \2534 );
xor \U$15523 ( \15655 , \15650 , \15654 );
and \U$15524 ( \15656 , \6281 , \3103 );
and \U$15525 ( \15657 , \6514 , \2934 );
nor \U$15526 ( \15658 , \15656 , \15657 );
xnor \U$15527 ( \15659 , \15658 , \2839 );
xor \U$15528 ( \15660 , \15655 , \15659 );
xor \U$15529 ( \15661 , \15646 , \15660 );
and \U$15530 ( \15662 , \3143 , \5996 );
and \U$15531 ( \15663 , \3395 , \5695 );
nor \U$15532 ( \15664 , \15662 , \15663 );
xnor \U$15533 ( \15665 , \15664 , \5687 );
and \U$15534 ( \15666 , \2826 , \6401 );
and \U$15535 ( \15667 , \3037 , \6143 );
nor \U$15536 ( \15668 , \15666 , \15667 );
xnor \U$15537 ( \15669 , \15668 , \6148 );
xor \U$15538 ( \15670 , \15665 , \15669 );
and \U$15539 ( \15671 , \2521 , \7055 );
and \U$15540 ( \15672 , \2757 , \6675 );
nor \U$15541 ( \15673 , \15671 , \15672 );
xnor \U$15542 ( \15674 , \15673 , \6680 );
xor \U$15543 ( \15675 , \15670 , \15674 );
and \U$15544 ( \15676 , \4364 , \4581 );
and \U$15545 ( \15677 , \4654 , \4424 );
nor \U$15546 ( \15678 , \15676 , \15677 );
xnor \U$15547 ( \15679 , \15678 , \4377 );
and \U$15548 ( \15680 , \3912 , \5011 );
and \U$15549 ( \15681 , \4160 , \4878 );
nor \U$15550 ( \15682 , \15680 , \15681 );
xnor \U$15551 ( \15683 , \15682 , \4762 );
xor \U$15552 ( \15684 , \15679 , \15683 );
and \U$15553 ( \15685 , \3646 , \5485 );
and \U$15554 ( \15686 , \3736 , \5275 );
nor \U$15555 ( \15687 , \15685 , \15686 );
xnor \U$15556 ( \15688 , \15687 , \5169 );
xor \U$15557 ( \15689 , \15684 , \15688 );
xor \U$15558 ( \15690 , \15675 , \15689 );
and \U$15559 ( \15691 , \5674 , \3357 );
and \U$15560 ( \15692 , \6030 , \3255 );
nor \U$15561 ( \15693 , \15691 , \15692 );
xnor \U$15562 ( \15694 , \15693 , \3156 );
and \U$15563 ( \15695 , \5156 , \3813 );
and \U$15564 ( \15696 , \5469 , \3557 );
nor \U$15565 ( \15697 , \15695 , \15696 );
xnor \U$15566 ( \15698 , \15697 , \3562 );
xor \U$15567 ( \15699 , \15694 , \15698 );
and \U$15568 ( \15700 , \4749 , \4132 );
and \U$15569 ( \15701 , \4922 , \4012 );
nor \U$15570 ( \15702 , \15700 , \15701 );
xnor \U$15571 ( \15703 , \15702 , \3925 );
xor \U$15572 ( \15704 , \15699 , \15703 );
xor \U$15573 ( \15705 , \15690 , \15704 );
xor \U$15574 ( \15706 , \15661 , \15705 );
and \U$15575 ( \15707 , \412 , \10118 );
and \U$15576 ( \15708 , \2182 , \7489 );
and \U$15577 ( \15709 , \2366 , \7137 );
nor \U$15578 ( \15710 , \15708 , \15709 );
xnor \U$15579 ( \15711 , \15710 , \7142 );
and \U$15580 ( \15712 , \1948 , \8019 );
and \U$15581 ( \15713 , \2090 , \7830 );
nor \U$15582 ( \15714 , \15712 , \15713 );
xnor \U$15583 ( \15715 , \15714 , \7713 );
xor \U$15584 ( \15716 , \15711 , \15715 );
and \U$15585 ( \15717 , \1684 , \8540 );
and \U$15586 ( \15718 , \1802 , \8292 );
nor \U$15587 ( \15719 , \15717 , \15718 );
xnor \U$15588 ( \15720 , \15719 , \8297 );
xor \U$15589 ( \15721 , \15716 , \15720 );
xor \U$15590 ( \15722 , \15707 , \15721 );
and \U$15591 ( \15723 , \1484 , \9333 );
and \U$15592 ( \15724 , \1601 , \9006 );
nor \U$15593 ( \15725 , \15723 , \15724 );
xnor \U$15594 ( \15726 , \15725 , \8848 );
and \U$15595 ( \15727 , \1192 , \9765 );
and \U$15596 ( \15728 , \1333 , \9644 );
nor \U$15597 ( \15729 , \15727 , \15728 );
xnor \U$15598 ( \15730 , \15729 , \9478 );
xor \U$15599 ( \15731 , \15726 , \15730 );
and \U$15600 ( \15732 , \474 , \10408 );
and \U$15601 ( \15733 , \1147 , \10116 );
nor \U$15602 ( \15734 , \15732 , \15733 );
xnor \U$15603 ( \15735 , \15734 , \10121 );
xor \U$15604 ( \15736 , \15731 , \15735 );
xor \U$15605 ( \15737 , \15722 , \15736 );
xor \U$15606 ( \15738 , \15706 , \15737 );
xor \U$15607 ( \15739 , \15620 , \15738 );
xor \U$15608 ( \15740 , \15574 , \15739 );
and \U$15609 ( \15741 , \15381 , \15395 );
and \U$15610 ( \15742 , \15395 , \15410 );
and \U$15611 ( \15743 , \15381 , \15410 );
or \U$15612 ( \15744 , \15741 , \15742 , \15743 );
and \U$15613 ( \15745 , \15425 , \15438 );
and \U$15614 ( \15746 , \15438 , \15453 );
and \U$15615 ( \15747 , \15425 , \15453 );
or \U$15616 ( \15748 , \15745 , \15746 , \15747 );
xor \U$15617 ( \15749 , \15744 , \15748 );
and \U$15618 ( \15750 , \15469 , \15483 );
and \U$15619 ( \15751 , \15483 , \15486 );
and \U$15620 ( \15752 , \15469 , \15486 );
or \U$15621 ( \15753 , \15750 , \15751 , \15752 );
xor \U$15622 ( \15754 , \15749 , \15753 );
and \U$15623 ( \15755 , \15329 , \15333 );
and \U$15624 ( \15756 , \15333 , \15338 );
and \U$15625 ( \15757 , \15329 , \15338 );
or \U$15626 ( \15758 , \15755 , \15756 , \15757 );
and \U$15627 ( \15759 , \15343 , \15347 );
and \U$15628 ( \15760 , \15347 , \15349 );
and \U$15629 ( \15761 , \15343 , \15349 );
or \U$15630 ( \15762 , \15759 , \15760 , \15761 );
xor \U$15631 ( \15763 , \15758 , \15762 );
and \U$15632 ( \15764 , \15355 , \15359 );
and \U$15633 ( \15765 , \15359 , \15364 );
and \U$15634 ( \15766 , \15355 , \15364 );
or \U$15635 ( \15767 , \15764 , \15765 , \15766 );
xor \U$15636 ( \15768 , \15763 , \15767 );
xor \U$15637 ( \15769 , \15754 , \15768 );
xor \U$15638 ( \15770 , \15740 , \15769 );
xor \U$15639 ( \15771 , \15560 , \15770 );
xor \U$15640 ( \15772 , \15551 , \15771 );
xor \U$15641 ( \15773 , \15535 , \15772 );
and \U$15642 ( \15774 , \15282 , \15522 );
xor \U$15643 ( \15775 , \15773 , \15774 );
and \U$15644 ( \15776 , \15523 , \15524 );
and \U$15645 ( \15777 , \15525 , \15528 );
or \U$15646 ( \15778 , \15776 , \15777 );
xor \U$15647 ( \15779 , \15775 , \15778 );
buf \U$15648 ( \15780 , \15779 );
buf \U$15649 ( \15781 , \15780 );
or \U$15650 ( \15782 , \1070 , \1171 , \1279 , \1390 , \1508 , \1629 , \1757 , \1888 , \2026 , \2167 , \2315 , \2466 , \2624 , \2785 , \2953 , \3124 , \3302 , \3483 , \3671 , \3862 , \4060 , \4261 , \4469 , \4680 , \4898 , \5118 , \5349 , \5580 , \5818 , \6059 , \6307 , \6558 , \6816 , \7077 , \7345 , \7616 , \7894 , \8175 , \8463 , \8754 , \9052 , \9353 , \9661 , \9972 , \10290 , \10611 , \10930 , \11248 , \11565 , \11881 , \12192 , \12500 , \12803 , \13099 , \13390 , \13673 , \13954 , \14227 , \14497 , \14763 , \15023 , \15278 , \15531 , \15781 );
and \U$15651 ( \15783 , \15539 , \15550 );
and \U$15652 ( \15784 , \15550 , \15771 );
and \U$15653 ( \15785 , \15539 , \15771 );
or \U$15654 ( \15786 , \15783 , \15784 , \15785 );
and \U$15655 ( \15787 , \15555 , \15559 );
and \U$15656 ( \15788 , \15559 , \15770 );
and \U$15657 ( \15789 , \15555 , \15770 );
or \U$15658 ( \15790 , \15787 , \15788 , \15789 );
and \U$15659 ( \15791 , \15564 , \15568 );
and \U$15660 ( \15792 , \15568 , \15573 );
and \U$15661 ( \15793 , \15564 , \15573 );
or \U$15662 ( \15794 , \15791 , \15792 , \15793 );
and \U$15663 ( \15795 , \15578 , \15619 );
and \U$15664 ( \15796 , \15619 , \15738 );
and \U$15665 ( \15797 , \15578 , \15738 );
or \U$15666 ( \15798 , \15795 , \15796 , \15797 );
xor \U$15667 ( \15799 , \15794 , \15798 );
and \U$15668 ( \15800 , \15754 , \15768 );
xor \U$15669 ( \15801 , \15799 , \15800 );
xor \U$15670 ( \15802 , \15790 , \15801 );
and \U$15671 ( \15803 , \15543 , \15547 );
and \U$15672 ( \15804 , \15547 , \15549 );
and \U$15673 ( \15805 , \15543 , \15549 );
or \U$15674 ( \15806 , \15803 , \15804 , \15805 );
and \U$15675 ( \15807 , \15574 , \15739 );
and \U$15676 ( \15808 , \15739 , \15769 );
and \U$15677 ( \15809 , \15574 , \15769 );
or \U$15678 ( \15810 , \15807 , \15808 , \15809 );
xor \U$15679 ( \15811 , \15806 , \15810 );
and \U$15680 ( \15812 , \15744 , \15748 );
and \U$15681 ( \15813 , \15748 , \15753 );
and \U$15682 ( \15814 , \15744 , \15753 );
or \U$15683 ( \15815 , \15812 , \15813 , \15814 );
and \U$15684 ( \15816 , \15758 , \15762 );
and \U$15685 ( \15817 , \15762 , \15767 );
and \U$15686 ( \15818 , \15758 , \15767 );
or \U$15687 ( \15819 , \15816 , \15817 , \15818 );
xor \U$15688 ( \15820 , \15815 , \15819 );
and \U$15689 ( \15821 , \15661 , \15705 );
and \U$15690 ( \15822 , \15705 , \15737 );
and \U$15691 ( \15823 , \15661 , \15737 );
or \U$15692 ( \15824 , \15821 , \15822 , \15823 );
xor \U$15693 ( \15825 , \15820 , \15824 );
and \U$15694 ( \15826 , \15589 , \15603 );
and \U$15695 ( \15827 , \15603 , \15618 );
and \U$15696 ( \15828 , \15589 , \15618 );
or \U$15697 ( \15829 , \15826 , \15827 , \15828 );
and \U$15698 ( \15830 , \15624 , \15628 );
and \U$15699 ( \15831 , \15628 , \15633 );
and \U$15700 ( \15832 , \15624 , \15633 );
or \U$15701 ( \15833 , \15830 , \15831 , \15832 );
and \U$15702 ( \15834 , \15635 , \15639 );
and \U$15703 ( \15835 , \15639 , \15644 );
and \U$15704 ( \15836 , \15635 , \15644 );
or \U$15705 ( \15837 , \15834 , \15835 , \15836 );
xor \U$15706 ( \15838 , \15833 , \15837 );
and \U$15707 ( \15839 , \15650 , \15654 );
and \U$15708 ( \15840 , \15654 , \15659 );
and \U$15709 ( \15841 , \15650 , \15659 );
or \U$15710 ( \15842 , \15839 , \15840 , \15841 );
xor \U$15711 ( \15843 , \15838 , \15842 );
and \U$15712 ( \15844 , \15665 , \15669 );
and \U$15713 ( \15845 , \15669 , \15674 );
and \U$15714 ( \15846 , \15665 , \15674 );
or \U$15715 ( \15847 , \15844 , \15845 , \15846 );
and \U$15716 ( \15848 , \15679 , \15683 );
and \U$15717 ( \15849 , \15683 , \15688 );
and \U$15718 ( \15850 , \15679 , \15688 );
or \U$15719 ( \15851 , \15848 , \15849 , \15850 );
xor \U$15720 ( \15852 , \15847 , \15851 );
and \U$15721 ( \15853 , \15694 , \15698 );
and \U$15722 ( \15854 , \15698 , \15703 );
and \U$15723 ( \15855 , \15694 , \15703 );
or \U$15724 ( \15856 , \15853 , \15854 , \15855 );
xor \U$15725 ( \15857 , \15852 , \15856 );
xor \U$15726 ( \15858 , \15843 , \15857 );
and \U$15727 ( \15859 , \15711 , \15715 );
and \U$15728 ( \15860 , \15715 , \15720 );
and \U$15729 ( \15861 , \15711 , \15720 );
or \U$15730 ( \15862 , \15859 , \15860 , \15861 );
and \U$15731 ( \15863 , \15726 , \15730 );
and \U$15732 ( \15864 , \15730 , \15735 );
and \U$15733 ( \15865 , \15726 , \15735 );
or \U$15734 ( \15866 , \15863 , \15864 , \15865 );
xnor \U$15735 ( \15867 , \15862 , \15866 );
xor \U$15736 ( \15868 , \15858 , \15867 );
xor \U$15737 ( \15869 , \15829 , \15868 );
and \U$15738 ( \15870 , \5469 , \3813 );
and \U$15739 ( \15871 , \5674 , \3557 );
nor \U$15740 ( \15872 , \15870 , \15871 );
xnor \U$15741 ( \15873 , \15872 , \3562 );
and \U$15742 ( \15874 , \4922 , \4132 );
and \U$15743 ( \15875 , \5156 , \4012 );
nor \U$15744 ( \15876 , \15874 , \15875 );
xnor \U$15745 ( \15877 , \15876 , \3925 );
xor \U$15746 ( \15878 , \15873 , \15877 );
and \U$15747 ( \15879 , \4654 , \4581 );
and \U$15748 ( \15880 , \4749 , \4424 );
nor \U$15749 ( \15881 , \15879 , \15880 );
xnor \U$15750 ( \15882 , \15881 , \4377 );
xor \U$15751 ( \15883 , \15878 , \15882 );
and \U$15752 ( \15884 , \4160 , \5011 );
and \U$15753 ( \15885 , \4364 , \4878 );
nor \U$15754 ( \15886 , \15884 , \15885 );
xnor \U$15755 ( \15887 , \15886 , \4762 );
and \U$15756 ( \15888 , \3736 , \5485 );
and \U$15757 ( \15889 , \3912 , \5275 );
nor \U$15758 ( \15890 , \15888 , \15889 );
xnor \U$15759 ( \15891 , \15890 , \5169 );
xor \U$15760 ( \15892 , \15887 , \15891 );
and \U$15761 ( \15893 , \3395 , \5996 );
and \U$15762 ( \15894 , \3646 , \5695 );
nor \U$15763 ( \15895 , \15893 , \15894 );
xnor \U$15764 ( \15896 , \15895 , \5687 );
xor \U$15765 ( \15897 , \15892 , \15896 );
xor \U$15766 ( \15898 , \15883 , \15897 );
and \U$15767 ( \15899 , \6945 , \2669 );
and \U$15768 ( \15900 , \7231 , \2538 );
nor \U$15769 ( \15901 , \15899 , \15900 );
xnor \U$15770 ( \15902 , \15901 , \2534 );
and \U$15771 ( \15903 , \6514 , \3103 );
and \U$15772 ( \15904 , \6790 , \2934 );
nor \U$15773 ( \15905 , \15903 , \15904 );
xnor \U$15774 ( \15906 , \15905 , \2839 );
xor \U$15775 ( \15907 , \15902 , \15906 );
and \U$15776 ( \15908 , \6030 , \3357 );
and \U$15777 ( \15909 , \6281 , \3255 );
nor \U$15778 ( \15910 , \15908 , \15909 );
xnor \U$15779 ( \15911 , \15910 , \3156 );
xor \U$15780 ( \15912 , \15907 , \15911 );
xor \U$15781 ( \15913 , \15898 , \15912 );
and \U$15782 ( \15914 , \3037 , \6401 );
and \U$15783 ( \15915 , \3143 , \6143 );
nor \U$15784 ( \15916 , \15914 , \15915 );
xnor \U$15785 ( \15917 , \15916 , \6148 );
and \U$15786 ( \15918 , \2757 , \7055 );
and \U$15787 ( \15919 , \2826 , \6675 );
nor \U$15788 ( \15920 , \15918 , \15919 );
xnor \U$15789 ( \15921 , \15920 , \6680 );
xor \U$15790 ( \15922 , \15917 , \15921 );
and \U$15791 ( \15923 , \2366 , \7489 );
and \U$15792 ( \15924 , \2521 , \7137 );
nor \U$15793 ( \15925 , \15923 , \15924 );
xnor \U$15794 ( \15926 , \15925 , \7142 );
xor \U$15795 ( \15927 , \15922 , \15926 );
and \U$15796 ( \15928 , \2090 , \8019 );
and \U$15797 ( \15929 , \2182 , \7830 );
nor \U$15798 ( \15930 , \15928 , \15929 );
xnor \U$15799 ( \15931 , \15930 , \7713 );
and \U$15800 ( \15932 , \1802 , \8540 );
and \U$15801 ( \15933 , \1948 , \8292 );
nor \U$15802 ( \15934 , \15932 , \15933 );
xnor \U$15803 ( \15935 , \15934 , \8297 );
xor \U$15804 ( \15936 , \15931 , \15935 );
and \U$15805 ( \15937 , \1601 , \9333 );
and \U$15806 ( \15938 , \1684 , \9006 );
nor \U$15807 ( \15939 , \15937 , \15938 );
xnor \U$15808 ( \15940 , \15939 , \8848 );
xor \U$15809 ( \15941 , \15936 , \15940 );
xor \U$15810 ( \15942 , \15927 , \15941 );
and \U$15811 ( \15943 , \1333 , \9765 );
and \U$15812 ( \15944 , \1484 , \9644 );
nor \U$15813 ( \15945 , \15943 , \15944 );
xnor \U$15814 ( \15946 , \15945 , \9478 );
and \U$15815 ( \15947 , \1147 , \10408 );
and \U$15816 ( \15948 , \1192 , \10116 );
nor \U$15817 ( \15949 , \15947 , \15948 );
xnor \U$15818 ( \15950 , \15949 , \10121 );
xor \U$15819 ( \15951 , \15946 , \15950 );
and \U$15820 ( \15952 , \474 , \10118 );
xor \U$15821 ( \15953 , \15951 , \15952 );
xor \U$15822 ( \15954 , \15942 , \15953 );
xor \U$15823 ( \15955 , \15913 , \15954 );
and \U$15824 ( \15956 , \10584 , \1086 );
not \U$15825 ( \15957 , \15956 );
xnor \U$15826 ( \15958 , \15957 , \487 );
and \U$15827 ( \15959 , \9897 , \1301 );
and \U$15828 ( \15960 , \10206 , \1246 );
nor \U$15829 ( \15961 , \15959 , \15960 );
xnor \U$15830 ( \15962 , \15961 , \1205 );
xor \U$15831 ( \15963 , \15958 , \15962 );
and \U$15832 ( \15964 , \9169 , \1578 );
and \U$15833 ( \15965 , \9465 , \1431 );
nor \U$15834 ( \15966 , \15964 , \15965 );
xnor \U$15835 ( \15967 , \15966 , \1436 );
xor \U$15836 ( \15968 , \15963 , \15967 );
and \U$15837 ( \15969 , \8652 , \1824 );
and \U$15838 ( \15970 , \8835 , \1739 );
nor \U$15839 ( \15971 , \15969 , \15970 );
xnor \U$15840 ( \15972 , \15971 , \1697 );
and \U$15841 ( \15973 , \8057 , \2121 );
and \U$15842 ( \15974 , \8349 , \2008 );
nor \U$15843 ( \15975 , \15973 , \15974 );
xnor \U$15844 ( \15976 , \15975 , \1961 );
xor \U$15845 ( \15977 , \15972 , \15976 );
and \U$15846 ( \15978 , \7556 , \2400 );
and \U$15847 ( \15979 , \7700 , \2246 );
nor \U$15848 ( \15980 , \15978 , \15979 );
xnor \U$15849 ( \15981 , \15980 , \2195 );
xor \U$15850 ( \15982 , \15977 , \15981 );
xor \U$15851 ( \15983 , \15968 , \15982 );
xor \U$15852 ( \15984 , \15955 , \15983 );
xor \U$15853 ( \15985 , \15869 , \15984 );
xor \U$15854 ( \15986 , \15825 , \15985 );
and \U$15855 ( \15987 , \15582 , \15586 );
and \U$15856 ( \15988 , \15586 , \15588 );
and \U$15857 ( \15989 , \15582 , \15588 );
or \U$15858 ( \15990 , \15987 , \15988 , \15989 );
and \U$15859 ( \15991 , \15593 , \15597 );
and \U$15860 ( \15992 , \15597 , \15602 );
and \U$15861 ( \15993 , \15593 , \15602 );
or \U$15862 ( \15994 , \15991 , \15992 , \15993 );
xor \U$15863 ( \15995 , \15990 , \15994 );
and \U$15864 ( \15996 , \15608 , \15612 );
and \U$15865 ( \15997 , \15612 , \15617 );
and \U$15866 ( \15998 , \15608 , \15617 );
or \U$15867 ( \15999 , \15996 , \15997 , \15998 );
xor \U$15868 ( \16000 , \15995 , \15999 );
and \U$15869 ( \16001 , \15634 , \15645 );
and \U$15870 ( \16002 , \15645 , \15660 );
and \U$15871 ( \16003 , \15634 , \15660 );
or \U$15872 ( \16004 , \16001 , \16002 , \16003 );
and \U$15873 ( \16005 , \15675 , \15689 );
and \U$15874 ( \16006 , \15689 , \15704 );
and \U$15875 ( \16007 , \15675 , \15704 );
or \U$15876 ( \16008 , \16005 , \16006 , \16007 );
xor \U$15877 ( \16009 , \16004 , \16008 );
and \U$15878 ( \16010 , \15707 , \15721 );
and \U$15879 ( \16011 , \15721 , \15736 );
and \U$15880 ( \16012 , \15707 , \15736 );
or \U$15881 ( \16013 , \16010 , \16011 , \16012 );
xor \U$15882 ( \16014 , \16009 , \16013 );
xor \U$15883 ( \16015 , \16000 , \16014 );
xor \U$15884 ( \16016 , \15986 , \16015 );
xor \U$15885 ( \16017 , \15811 , \16016 );
xor \U$15886 ( \16018 , \15802 , \16017 );
xor \U$15887 ( \16019 , \15786 , \16018 );
and \U$15888 ( \16020 , \15535 , \15772 );
xor \U$15889 ( \16021 , \16019 , \16020 );
and \U$15890 ( \16022 , \15773 , \15774 );
and \U$15891 ( \16023 , \15775 , \15778 );
or \U$15892 ( \16024 , \16022 , \16023 );
xor \U$15893 ( \16025 , \16021 , \16024 );
buf \U$15894 ( \16026 , \16025 );
buf \U$15895 ( \16027 , \16026 );
and \U$15896 ( \16028 , \15790 , \15801 );
and \U$15897 ( \16029 , \15801 , \16017 );
and \U$15898 ( \16030 , \15790 , \16017 );
or \U$15899 ( \16031 , \16028 , \16029 , \16030 );
and \U$15900 ( \16032 , \15806 , \15810 );
and \U$15901 ( \16033 , \15810 , \16016 );
and \U$15902 ( \16034 , \15806 , \16016 );
or \U$15903 ( \16035 , \16032 , \16033 , \16034 );
and \U$15904 ( \16036 , \15815 , \15819 );
and \U$15905 ( \16037 , \15819 , \15824 );
and \U$15906 ( \16038 , \15815 , \15824 );
or \U$15907 ( \16039 , \16036 , \16037 , \16038 );
and \U$15908 ( \16040 , \15829 , \15868 );
and \U$15909 ( \16041 , \15868 , \15984 );
and \U$15910 ( \16042 , \15829 , \15984 );
or \U$15911 ( \16043 , \16040 , \16041 , \16042 );
xor \U$15912 ( \16044 , \16039 , \16043 );
and \U$15913 ( \16045 , \16000 , \16014 );
xor \U$15914 ( \16046 , \16044 , \16045 );
xor \U$15915 ( \16047 , \16035 , \16046 );
and \U$15916 ( \16048 , \15794 , \15798 );
and \U$15917 ( \16049 , \15798 , \15800 );
and \U$15918 ( \16050 , \15794 , \15800 );
or \U$15919 ( \16051 , \16048 , \16049 , \16050 );
and \U$15920 ( \16052 , \15825 , \15985 );
and \U$15921 ( \16053 , \15985 , \16015 );
and \U$15922 ( \16054 , \15825 , \16015 );
or \U$15923 ( \16055 , \16052 , \16053 , \16054 );
xor \U$15924 ( \16056 , \16051 , \16055 );
and \U$15925 ( \16057 , \15990 , \15994 );
and \U$15926 ( \16058 , \15994 , \15999 );
and \U$15927 ( \16059 , \15990 , \15999 );
or \U$15928 ( \16060 , \16057 , \16058 , \16059 );
and \U$15929 ( \16061 , \16004 , \16008 );
and \U$15930 ( \16062 , \16008 , \16013 );
and \U$15931 ( \16063 , \16004 , \16013 );
or \U$15932 ( \16064 , \16061 , \16062 , \16063 );
xor \U$15933 ( \16065 , \16060 , \16064 );
and \U$15934 ( \16066 , \15913 , \15954 );
and \U$15935 ( \16067 , \15954 , \15983 );
and \U$15936 ( \16068 , \15913 , \15983 );
or \U$15937 ( \16069 , \16066 , \16067 , \16068 );
xor \U$15938 ( \16070 , \16065 , \16069 );
and \U$15939 ( \16071 , \15843 , \15857 );
and \U$15940 ( \16072 , \15857 , \15867 );
and \U$15941 ( \16073 , \15843 , \15867 );
or \U$15942 ( \16074 , \16071 , \16072 , \16073 );
not \U$15943 ( \16075 , \487 );
and \U$15944 ( \16076 , \10206 , \1301 );
and \U$15945 ( \16077 , \10584 , \1246 );
nor \U$15946 ( \16078 , \16076 , \16077 );
xnor \U$15947 ( \16079 , \16078 , \1205 );
xor \U$15948 ( \16080 , \16075 , \16079 );
and \U$15949 ( \16081 , \9465 , \1578 );
and \U$15950 ( \16082 , \9897 , \1431 );
nor \U$15951 ( \16083 , \16081 , \16082 );
xnor \U$15952 ( \16084 , \16083 , \1436 );
xor \U$15953 ( \16085 , \16080 , \16084 );
and \U$15954 ( \16086 , \5674 , \3813 );
and \U$15955 ( \16087 , \6030 , \3557 );
nor \U$15956 ( \16088 , \16086 , \16087 );
xnor \U$15957 ( \16089 , \16088 , \3562 );
and \U$15958 ( \16090 , \5156 , \4132 );
and \U$15959 ( \16091 , \5469 , \4012 );
nor \U$15960 ( \16092 , \16090 , \16091 );
xnor \U$15961 ( \16093 , \16092 , \3925 );
xor \U$15962 ( \16094 , \16089 , \16093 );
and \U$15963 ( \16095 , \4749 , \4581 );
and \U$15964 ( \16096 , \4922 , \4424 );
nor \U$15965 ( \16097 , \16095 , \16096 );
xnor \U$15966 ( \16098 , \16097 , \4377 );
xor \U$15967 ( \16099 , \16094 , \16098 );
and \U$15968 ( \16100 , \8835 , \1824 );
and \U$15969 ( \16101 , \9169 , \1739 );
nor \U$15970 ( \16102 , \16100 , \16101 );
xnor \U$15971 ( \16103 , \16102 , \1697 );
and \U$15972 ( \16104 , \8349 , \2121 );
and \U$15973 ( \16105 , \8652 , \2008 );
nor \U$15974 ( \16106 , \16104 , \16105 );
xnor \U$15975 ( \16107 , \16106 , \1961 );
xor \U$15976 ( \16108 , \16103 , \16107 );
and \U$15977 ( \16109 , \7700 , \2400 );
and \U$15978 ( \16110 , \8057 , \2246 );
nor \U$15979 ( \16111 , \16109 , \16110 );
xnor \U$15980 ( \16112 , \16111 , \2195 );
xor \U$15981 ( \16113 , \16108 , \16112 );
xor \U$15982 ( \16114 , \16099 , \16113 );
and \U$15983 ( \16115 , \7231 , \2669 );
and \U$15984 ( \16116 , \7556 , \2538 );
nor \U$15985 ( \16117 , \16115 , \16116 );
xnor \U$15986 ( \16118 , \16117 , \2534 );
and \U$15987 ( \16119 , \6790 , \3103 );
and \U$15988 ( \16120 , \6945 , \2934 );
nor \U$15989 ( \16121 , \16119 , \16120 );
xnor \U$15990 ( \16122 , \16121 , \2839 );
xor \U$15991 ( \16123 , \16118 , \16122 );
and \U$15992 ( \16124 , \6281 , \3357 );
and \U$15993 ( \16125 , \6514 , \3255 );
nor \U$15994 ( \16126 , \16124 , \16125 );
xnor \U$15995 ( \16127 , \16126 , \3156 );
xor \U$15996 ( \16128 , \16123 , \16127 );
xor \U$15997 ( \16129 , \16114 , \16128 );
xor \U$15998 ( \16130 , \16085 , \16129 );
and \U$15999 ( \16131 , \4364 , \5011 );
and \U$16000 ( \16132 , \4654 , \4878 );
nor \U$16001 ( \16133 , \16131 , \16132 );
xnor \U$16002 ( \16134 , \16133 , \4762 );
and \U$16003 ( \16135 , \3912 , \5485 );
and \U$16004 ( \16136 , \4160 , \5275 );
nor \U$16005 ( \16137 , \16135 , \16136 );
xnor \U$16006 ( \16138 , \16137 , \5169 );
xor \U$16007 ( \16139 , \16134 , \16138 );
and \U$16008 ( \16140 , \3646 , \5996 );
and \U$16009 ( \16141 , \3736 , \5695 );
nor \U$16010 ( \16142 , \16140 , \16141 );
xnor \U$16011 ( \16143 , \16142 , \5687 );
xor \U$16012 ( \16144 , \16139 , \16143 );
and \U$16013 ( \16145 , \3143 , \6401 );
and \U$16014 ( \16146 , \3395 , \6143 );
nor \U$16015 ( \16147 , \16145 , \16146 );
xnor \U$16016 ( \16148 , \16147 , \6148 );
and \U$16017 ( \16149 , \2826 , \7055 );
and \U$16018 ( \16150 , \3037 , \6675 );
nor \U$16019 ( \16151 , \16149 , \16150 );
xnor \U$16020 ( \16152 , \16151 , \6680 );
xor \U$16021 ( \16153 , \16148 , \16152 );
and \U$16022 ( \16154 , \2521 , \7489 );
and \U$16023 ( \16155 , \2757 , \7137 );
nor \U$16024 ( \16156 , \16154 , \16155 );
xnor \U$16025 ( \16157 , \16156 , \7142 );
xor \U$16026 ( \16158 , \16153 , \16157 );
xor \U$16027 ( \16159 , \16144 , \16158 );
and \U$16028 ( \16160 , \2182 , \8019 );
and \U$16029 ( \16161 , \2366 , \7830 );
nor \U$16030 ( \16162 , \16160 , \16161 );
xnor \U$16031 ( \16163 , \16162 , \7713 );
and \U$16032 ( \16164 , \1948 , \8540 );
and \U$16033 ( \16165 , \2090 , \8292 );
nor \U$16034 ( \16166 , \16164 , \16165 );
xnor \U$16035 ( \16167 , \16166 , \8297 );
xor \U$16036 ( \16168 , \16163 , \16167 );
and \U$16037 ( \16169 , \1684 , \9333 );
and \U$16038 ( \16170 , \1802 , \9006 );
nor \U$16039 ( \16171 , \16169 , \16170 );
xnor \U$16040 ( \16172 , \16171 , \8848 );
xor \U$16041 ( \16173 , \16168 , \16172 );
xor \U$16042 ( \16174 , \16159 , \16173 );
xor \U$16043 ( \16175 , \16130 , \16174 );
xor \U$16044 ( \16176 , \16074 , \16175 );
and \U$16045 ( \16177 , \15958 , \15962 );
and \U$16046 ( \16178 , \15962 , \15967 );
and \U$16047 ( \16179 , \15958 , \15967 );
or \U$16048 ( \16180 , \16177 , \16178 , \16179 );
and \U$16049 ( \16181 , \15972 , \15976 );
and \U$16050 ( \16182 , \15976 , \15981 );
and \U$16051 ( \16183 , \15972 , \15981 );
or \U$16052 ( \16184 , \16181 , \16182 , \16183 );
xor \U$16053 ( \16185 , \16180 , \16184 );
and \U$16054 ( \16186 , \15902 , \15906 );
and \U$16055 ( \16187 , \15906 , \15911 );
and \U$16056 ( \16188 , \15902 , \15911 );
or \U$16057 ( \16189 , \16186 , \16187 , \16188 );
xor \U$16058 ( \16190 , \16185 , \16189 );
and \U$16059 ( \16191 , \15873 , \15877 );
and \U$16060 ( \16192 , \15877 , \15882 );
and \U$16061 ( \16193 , \15873 , \15882 );
or \U$16062 ( \16194 , \16191 , \16192 , \16193 );
and \U$16063 ( \16195 , \15887 , \15891 );
and \U$16064 ( \16196 , \15891 , \15896 );
and \U$16065 ( \16197 , \15887 , \15896 );
or \U$16066 ( \16198 , \16195 , \16196 , \16197 );
xor \U$16067 ( \16199 , \16194 , \16198 );
and \U$16068 ( \16200 , \15917 , \15921 );
and \U$16069 ( \16201 , \15921 , \15926 );
and \U$16070 ( \16202 , \15917 , \15926 );
or \U$16071 ( \16203 , \16200 , \16201 , \16202 );
xor \U$16072 ( \16204 , \16199 , \16203 );
xor \U$16073 ( \16205 , \16190 , \16204 );
and \U$16074 ( \16206 , \15931 , \15935 );
and \U$16075 ( \16207 , \15935 , \15940 );
and \U$16076 ( \16208 , \15931 , \15940 );
or \U$16077 ( \16209 , \16206 , \16207 , \16208 );
and \U$16078 ( \16210 , \15946 , \15950 );
and \U$16079 ( \16211 , \15950 , \15952 );
and \U$16080 ( \16212 , \15946 , \15952 );
or \U$16081 ( \16213 , \16210 , \16211 , \16212 );
xor \U$16082 ( \16214 , \16209 , \16213 );
and \U$16083 ( \16215 , \1484 , \9765 );
and \U$16084 ( \16216 , \1601 , \9644 );
nor \U$16085 ( \16217 , \16215 , \16216 );
xnor \U$16086 ( \16218 , \16217 , \9478 );
and \U$16087 ( \16219 , \1192 , \10408 );
and \U$16088 ( \16220 , \1333 , \10116 );
nor \U$16089 ( \16221 , \16219 , \16220 );
xnor \U$16090 ( \16222 , \16221 , \10121 );
xor \U$16091 ( \16223 , \16218 , \16222 );
and \U$16092 ( \16224 , \1147 , \10118 );
xor \U$16093 ( \16225 , \16223 , \16224 );
xor \U$16094 ( \16226 , \16214 , \16225 );
xor \U$16095 ( \16227 , \16205 , \16226 );
xor \U$16096 ( \16228 , \16176 , \16227 );
xor \U$16097 ( \16229 , \16070 , \16228 );
and \U$16098 ( \16230 , \15833 , \15837 );
and \U$16099 ( \16231 , \15837 , \15842 );
and \U$16100 ( \16232 , \15833 , \15842 );
or \U$16101 ( \16233 , \16230 , \16231 , \16232 );
and \U$16102 ( \16234 , \15847 , \15851 );
and \U$16103 ( \16235 , \15851 , \15856 );
and \U$16104 ( \16236 , \15847 , \15856 );
or \U$16105 ( \16237 , \16234 , \16235 , \16236 );
xor \U$16106 ( \16238 , \16233 , \16237 );
or \U$16107 ( \16239 , \15862 , \15866 );
xor \U$16108 ( \16240 , \16238 , \16239 );
and \U$16109 ( \16241 , \15883 , \15897 );
and \U$16110 ( \16242 , \15897 , \15912 );
and \U$16111 ( \16243 , \15883 , \15912 );
or \U$16112 ( \16244 , \16241 , \16242 , \16243 );
and \U$16113 ( \16245 , \15927 , \15941 );
and \U$16114 ( \16246 , \15941 , \15953 );
and \U$16115 ( \16247 , \15927 , \15953 );
or \U$16116 ( \16248 , \16245 , \16246 , \16247 );
xor \U$16117 ( \16249 , \16244 , \16248 );
and \U$16118 ( \16250 , \15968 , \15982 );
xor \U$16119 ( \16251 , \16249 , \16250 );
xor \U$16120 ( \16252 , \16240 , \16251 );
xor \U$16121 ( \16253 , \16229 , \16252 );
xor \U$16122 ( \16254 , \16056 , \16253 );
xor \U$16123 ( \16255 , \16047 , \16254 );
xor \U$16124 ( \16256 , \16031 , \16255 );
and \U$16125 ( \16257 , \15786 , \16018 );
xor \U$16126 ( \16258 , \16256 , \16257 );
and \U$16127 ( \16259 , \16019 , \16020 );
and \U$16128 ( \16260 , \16021 , \16024 );
or \U$16129 ( \16261 , \16259 , \16260 );
xor \U$16130 ( \16262 , \16258 , \16261 );
buf \U$16131 ( \16263 , \16262 );
buf \U$16132 ( \16264 , \16263 );
and \U$16133 ( \16265 , \16035 , \16046 );
and \U$16134 ( \16266 , \16046 , \16254 );
and \U$16135 ( \16267 , \16035 , \16254 );
or \U$16136 ( \16268 , \16265 , \16266 , \16267 );
and \U$16137 ( \16269 , \16051 , \16055 );
and \U$16138 ( \16270 , \16055 , \16253 );
and \U$16139 ( \16271 , \16051 , \16253 );
or \U$16140 ( \16272 , \16269 , \16270 , \16271 );
and \U$16141 ( \16273 , \16060 , \16064 );
and \U$16142 ( \16274 , \16064 , \16069 );
and \U$16143 ( \16275 , \16060 , \16069 );
or \U$16144 ( \16276 , \16273 , \16274 , \16275 );
and \U$16145 ( \16277 , \16074 , \16175 );
and \U$16146 ( \16278 , \16175 , \16227 );
and \U$16147 ( \16279 , \16074 , \16227 );
or \U$16148 ( \16280 , \16277 , \16278 , \16279 );
xor \U$16149 ( \16281 , \16276 , \16280 );
and \U$16150 ( \16282 , \16240 , \16251 );
xor \U$16151 ( \16283 , \16281 , \16282 );
xor \U$16152 ( \16284 , \16272 , \16283 );
and \U$16153 ( \16285 , \16039 , \16043 );
and \U$16154 ( \16286 , \16043 , \16045 );
and \U$16155 ( \16287 , \16039 , \16045 );
or \U$16156 ( \16288 , \16285 , \16286 , \16287 );
and \U$16157 ( \16289 , \16070 , \16228 );
and \U$16158 ( \16290 , \16228 , \16252 );
and \U$16159 ( \16291 , \16070 , \16252 );
or \U$16160 ( \16292 , \16289 , \16290 , \16291 );
xor \U$16161 ( \16293 , \16288 , \16292 );
and \U$16162 ( \16294 , \16233 , \16237 );
and \U$16163 ( \16295 , \16237 , \16239 );
and \U$16164 ( \16296 , \16233 , \16239 );
or \U$16165 ( \16297 , \16294 , \16295 , \16296 );
and \U$16166 ( \16298 , \16244 , \16248 );
and \U$16167 ( \16299 , \16248 , \16250 );
and \U$16168 ( \16300 , \16244 , \16250 );
or \U$16169 ( \16301 , \16298 , \16299 , \16300 );
xor \U$16170 ( \16302 , \16297 , \16301 );
and \U$16171 ( \16303 , \16085 , \16129 );
and \U$16172 ( \16304 , \16129 , \16174 );
and \U$16173 ( \16305 , \16085 , \16174 );
or \U$16174 ( \16306 , \16303 , \16304 , \16305 );
xor \U$16175 ( \16307 , \16302 , \16306 );
and \U$16176 ( \16308 , \16190 , \16204 );
and \U$16177 ( \16309 , \16204 , \16226 );
and \U$16178 ( \16310 , \16190 , \16226 );
or \U$16179 ( \16311 , \16308 , \16309 , \16310 );
and \U$16180 ( \16312 , \16075 , \16079 );
and \U$16181 ( \16313 , \16079 , \16084 );
and \U$16182 ( \16314 , \16075 , \16084 );
or \U$16183 ( \16315 , \16312 , \16313 , \16314 );
and \U$16184 ( \16316 , \16103 , \16107 );
and \U$16185 ( \16317 , \16107 , \16112 );
and \U$16186 ( \16318 , \16103 , \16112 );
or \U$16187 ( \16319 , \16316 , \16317 , \16318 );
xor \U$16188 ( \16320 , \16315 , \16319 );
and \U$16189 ( \16321 , \16118 , \16122 );
and \U$16190 ( \16322 , \16122 , \16127 );
and \U$16191 ( \16323 , \16118 , \16127 );
or \U$16192 ( \16324 , \16321 , \16322 , \16323 );
xor \U$16193 ( \16325 , \16320 , \16324 );
xor \U$16194 ( \16326 , \16311 , \16325 );
and \U$16195 ( \16327 , \16089 , \16093 );
and \U$16196 ( \16328 , \16093 , \16098 );
and \U$16197 ( \16329 , \16089 , \16098 );
or \U$16198 ( \16330 , \16327 , \16328 , \16329 );
and \U$16199 ( \16331 , \16134 , \16138 );
and \U$16200 ( \16332 , \16138 , \16143 );
and \U$16201 ( \16333 , \16134 , \16143 );
or \U$16202 ( \16334 , \16331 , \16332 , \16333 );
xor \U$16203 ( \16335 , \16330 , \16334 );
and \U$16204 ( \16336 , \16148 , \16152 );
and \U$16205 ( \16337 , \16152 , \16157 );
and \U$16206 ( \16338 , \16148 , \16157 );
or \U$16207 ( \16339 , \16336 , \16337 , \16338 );
xor \U$16208 ( \16340 , \16335 , \16339 );
xor \U$16209 ( \16341 , \16326 , \16340 );
xor \U$16210 ( \16342 , \16307 , \16341 );
and \U$16211 ( \16343 , \16180 , \16184 );
and \U$16212 ( \16344 , \16184 , \16189 );
and \U$16213 ( \16345 , \16180 , \16189 );
or \U$16214 ( \16346 , \16343 , \16344 , \16345 );
and \U$16215 ( \16347 , \16194 , \16198 );
and \U$16216 ( \16348 , \16198 , \16203 );
and \U$16217 ( \16349 , \16194 , \16203 );
or \U$16218 ( \16350 , \16347 , \16348 , \16349 );
xor \U$16219 ( \16351 , \16346 , \16350 );
and \U$16220 ( \16352 , \16209 , \16213 );
and \U$16221 ( \16353 , \16213 , \16225 );
and \U$16222 ( \16354 , \16209 , \16225 );
or \U$16223 ( \16355 , \16352 , \16353 , \16354 );
xor \U$16224 ( \16356 , \16351 , \16355 );
and \U$16225 ( \16357 , \16099 , \16113 );
and \U$16226 ( \16358 , \16113 , \16128 );
and \U$16227 ( \16359 , \16099 , \16128 );
or \U$16228 ( \16360 , \16357 , \16358 , \16359 );
and \U$16229 ( \16361 , \16144 , \16158 );
and \U$16230 ( \16362 , \16158 , \16173 );
and \U$16231 ( \16363 , \16144 , \16173 );
or \U$16232 ( \16364 , \16361 , \16362 , \16363 );
xor \U$16233 ( \16365 , \16360 , \16364 );
and \U$16234 ( \16366 , \10584 , \1301 );
not \U$16235 ( \16367 , \16366 );
xnor \U$16236 ( \16368 , \16367 , \1205 );
and \U$16237 ( \16369 , \9897 , \1578 );
and \U$16238 ( \16370 , \10206 , \1431 );
nor \U$16239 ( \16371 , \16369 , \16370 );
xnor \U$16240 ( \16372 , \16371 , \1436 );
xor \U$16241 ( \16373 , \16368 , \16372 );
and \U$16242 ( \16374 , \9169 , \1824 );
and \U$16243 ( \16375 , \9465 , \1739 );
nor \U$16244 ( \16376 , \16374 , \16375 );
xnor \U$16245 ( \16377 , \16376 , \1697 );
xor \U$16246 ( \16378 , \16373 , \16377 );
xor \U$16247 ( \16379 , \16365 , \16378 );
xor \U$16248 ( \16380 , \16356 , \16379 );
and \U$16249 ( \16381 , \2090 , \8540 );
and \U$16250 ( \16382 , \2182 , \8292 );
nor \U$16251 ( \16383 , \16381 , \16382 );
xnor \U$16252 ( \16384 , \16383 , \8297 );
and \U$16253 ( \16385 , \1802 , \9333 );
and \U$16254 ( \16386 , \1948 , \9006 );
nor \U$16255 ( \16387 , \16385 , \16386 );
xnor \U$16256 ( \16388 , \16387 , \8848 );
xor \U$16257 ( \16389 , \16384 , \16388 );
and \U$16258 ( \16390 , \1601 , \9765 );
and \U$16259 ( \16391 , \1684 , \9644 );
nor \U$16260 ( \16392 , \16390 , \16391 );
xnor \U$16261 ( \16393 , \16392 , \9478 );
xor \U$16262 ( \16394 , \16389 , \16393 );
and \U$16263 ( \16395 , \4160 , \5485 );
and \U$16264 ( \16396 , \4364 , \5275 );
nor \U$16265 ( \16397 , \16395 , \16396 );
xnor \U$16266 ( \16398 , \16397 , \5169 );
and \U$16267 ( \16399 , \3736 , \5996 );
and \U$16268 ( \16400 , \3912 , \5695 );
nor \U$16269 ( \16401 , \16399 , \16400 );
xnor \U$16270 ( \16402 , \16401 , \5687 );
xor \U$16271 ( \16403 , \16398 , \16402 );
and \U$16272 ( \16404 , \3395 , \6401 );
and \U$16273 ( \16405 , \3646 , \6143 );
nor \U$16274 ( \16406 , \16404 , \16405 );
xnor \U$16275 ( \16407 , \16406 , \6148 );
xor \U$16276 ( \16408 , \16403 , \16407 );
xor \U$16277 ( \16409 , \16394 , \16408 );
and \U$16278 ( \16410 , \3037 , \7055 );
and \U$16279 ( \16411 , \3143 , \6675 );
nor \U$16280 ( \16412 , \16410 , \16411 );
xnor \U$16281 ( \16413 , \16412 , \6680 );
and \U$16282 ( \16414 , \2757 , \7489 );
and \U$16283 ( \16415 , \2826 , \7137 );
nor \U$16284 ( \16416 , \16414 , \16415 );
xnor \U$16285 ( \16417 , \16416 , \7142 );
xor \U$16286 ( \16418 , \16413 , \16417 );
and \U$16287 ( \16419 , \2366 , \8019 );
and \U$16288 ( \16420 , \2521 , \7830 );
nor \U$16289 ( \16421 , \16419 , \16420 );
xnor \U$16290 ( \16422 , \16421 , \7713 );
xor \U$16291 ( \16423 , \16418 , \16422 );
xor \U$16292 ( \16424 , \16409 , \16423 );
and \U$16293 ( \16425 , \5469 , \4132 );
and \U$16294 ( \16426 , \5674 , \4012 );
nor \U$16295 ( \16427 , \16425 , \16426 );
xnor \U$16296 ( \16428 , \16427 , \3925 );
and \U$16297 ( \16429 , \4922 , \4581 );
and \U$16298 ( \16430 , \5156 , \4424 );
nor \U$16299 ( \16431 , \16429 , \16430 );
xnor \U$16300 ( \16432 , \16431 , \4377 );
xor \U$16301 ( \16433 , \16428 , \16432 );
and \U$16302 ( \16434 , \4654 , \5011 );
and \U$16303 ( \16435 , \4749 , \4878 );
nor \U$16304 ( \16436 , \16434 , \16435 );
xnor \U$16305 ( \16437 , \16436 , \4762 );
xor \U$16306 ( \16438 , \16433 , \16437 );
and \U$16307 ( \16439 , \6945 , \3103 );
and \U$16308 ( \16440 , \7231 , \2934 );
nor \U$16309 ( \16441 , \16439 , \16440 );
xnor \U$16310 ( \16442 , \16441 , \2839 );
and \U$16311 ( \16443 , \6514 , \3357 );
and \U$16312 ( \16444 , \6790 , \3255 );
nor \U$16313 ( \16445 , \16443 , \16444 );
xnor \U$16314 ( \16446 , \16445 , \3156 );
xor \U$16315 ( \16447 , \16442 , \16446 );
and \U$16316 ( \16448 , \6030 , \3813 );
and \U$16317 ( \16449 , \6281 , \3557 );
nor \U$16318 ( \16450 , \16448 , \16449 );
xnor \U$16319 ( \16451 , \16450 , \3562 );
xor \U$16320 ( \16452 , \16447 , \16451 );
xor \U$16321 ( \16453 , \16438 , \16452 );
and \U$16322 ( \16454 , \8652 , \2121 );
and \U$16323 ( \16455 , \8835 , \2008 );
nor \U$16324 ( \16456 , \16454 , \16455 );
xnor \U$16325 ( \16457 , \16456 , \1961 );
and \U$16326 ( \16458 , \8057 , \2400 );
and \U$16327 ( \16459 , \8349 , \2246 );
nor \U$16328 ( \16460 , \16458 , \16459 );
xnor \U$16329 ( \16461 , \16460 , \2195 );
xor \U$16330 ( \16462 , \16457 , \16461 );
and \U$16331 ( \16463 , \7556 , \2669 );
and \U$16332 ( \16464 , \7700 , \2538 );
nor \U$16333 ( \16465 , \16463 , \16464 );
xnor \U$16334 ( \16466 , \16465 , \2534 );
xor \U$16335 ( \16467 , \16462 , \16466 );
xor \U$16336 ( \16468 , \16453 , \16467 );
xor \U$16337 ( \16469 , \16424 , \16468 );
and \U$16338 ( \16470 , \16218 , \16222 );
and \U$16339 ( \16471 , \16222 , \16224 );
and \U$16340 ( \16472 , \16218 , \16224 );
or \U$16341 ( \16473 , \16470 , \16471 , \16472 );
and \U$16342 ( \16474 , \16163 , \16167 );
and \U$16343 ( \16475 , \16167 , \16172 );
and \U$16344 ( \16476 , \16163 , \16172 );
or \U$16345 ( \16477 , \16474 , \16475 , \16476 );
xor \U$16346 ( \16478 , \16473 , \16477 );
and \U$16347 ( \16479 , \1333 , \10408 );
and \U$16348 ( \16480 , \1484 , \10116 );
nor \U$16349 ( \16481 , \16479 , \16480 );
xnor \U$16350 ( \16482 , \16481 , \10121 );
and \U$16351 ( \16483 , \1192 , \10118 );
xnor \U$16352 ( \16484 , \16482 , \16483 );
xor \U$16353 ( \16485 , \16478 , \16484 );
xor \U$16354 ( \16486 , \16469 , \16485 );
xor \U$16355 ( \16487 , \16380 , \16486 );
xor \U$16356 ( \16488 , \16342 , \16487 );
xor \U$16357 ( \16489 , \16293 , \16488 );
xor \U$16358 ( \16490 , \16284 , \16489 );
xor \U$16359 ( \16491 , \16268 , \16490 );
and \U$16360 ( \16492 , \16031 , \16255 );
xor \U$16361 ( \16493 , \16491 , \16492 );
and \U$16362 ( \16494 , \16256 , \16257 );
and \U$16363 ( \16495 , \16258 , \16261 );
or \U$16364 ( \16496 , \16494 , \16495 );
xor \U$16365 ( \16497 , \16493 , \16496 );
buf \U$16366 ( \16498 , \16497 );
buf \U$16367 ( \16499 , \16498 );
and \U$16368 ( \16500 , \16272 , \16283 );
and \U$16369 ( \16501 , \16283 , \16489 );
and \U$16370 ( \16502 , \16272 , \16489 );
or \U$16371 ( \16503 , \16500 , \16501 , \16502 );
and \U$16372 ( \16504 , \16288 , \16292 );
and \U$16373 ( \16505 , \16292 , \16488 );
and \U$16374 ( \16506 , \16288 , \16488 );
or \U$16375 ( \16507 , \16504 , \16505 , \16506 );
and \U$16376 ( \16508 , \16297 , \16301 );
and \U$16377 ( \16509 , \16301 , \16306 );
and \U$16378 ( \16510 , \16297 , \16306 );
or \U$16379 ( \16511 , \16508 , \16509 , \16510 );
and \U$16380 ( \16512 , \16311 , \16325 );
and \U$16381 ( \16513 , \16325 , \16340 );
and \U$16382 ( \16514 , \16311 , \16340 );
or \U$16383 ( \16515 , \16512 , \16513 , \16514 );
xor \U$16384 ( \16516 , \16511 , \16515 );
and \U$16385 ( \16517 , \16356 , \16379 );
and \U$16386 ( \16518 , \16379 , \16486 );
and \U$16387 ( \16519 , \16356 , \16486 );
or \U$16388 ( \16520 , \16517 , \16518 , \16519 );
xor \U$16389 ( \16521 , \16516 , \16520 );
xor \U$16390 ( \16522 , \16507 , \16521 );
and \U$16391 ( \16523 , \16276 , \16280 );
and \U$16392 ( \16524 , \16280 , \16282 );
and \U$16393 ( \16525 , \16276 , \16282 );
or \U$16394 ( \16526 , \16523 , \16524 , \16525 );
and \U$16395 ( \16527 , \16307 , \16341 );
and \U$16396 ( \16528 , \16341 , \16487 );
and \U$16397 ( \16529 , \16307 , \16487 );
or \U$16398 ( \16530 , \16527 , \16528 , \16529 );
xor \U$16399 ( \16531 , \16526 , \16530 );
and \U$16400 ( \16532 , \16315 , \16319 );
and \U$16401 ( \16533 , \16319 , \16324 );
and \U$16402 ( \16534 , \16315 , \16324 );
or \U$16403 ( \16535 , \16532 , \16533 , \16534 );
and \U$16404 ( \16536 , \16330 , \16334 );
and \U$16405 ( \16537 , \16334 , \16339 );
and \U$16406 ( \16538 , \16330 , \16339 );
or \U$16407 ( \16539 , \16536 , \16537 , \16538 );
xor \U$16408 ( \16540 , \16535 , \16539 );
and \U$16409 ( \16541 , \16473 , \16477 );
and \U$16410 ( \16542 , \16477 , \16484 );
and \U$16411 ( \16543 , \16473 , \16484 );
or \U$16412 ( \16544 , \16541 , \16542 , \16543 );
xor \U$16413 ( \16545 , \16540 , \16544 );
and \U$16414 ( \16546 , \16346 , \16350 );
and \U$16415 ( \16547 , \16350 , \16355 );
and \U$16416 ( \16548 , \16346 , \16355 );
or \U$16417 ( \16549 , \16546 , \16547 , \16548 );
and \U$16418 ( \16550 , \16360 , \16364 );
and \U$16419 ( \16551 , \16364 , \16378 );
and \U$16420 ( \16552 , \16360 , \16378 );
or \U$16421 ( \16553 , \16550 , \16551 , \16552 );
xor \U$16422 ( \16554 , \16549 , \16553 );
and \U$16423 ( \16555 , \16424 , \16468 );
and \U$16424 ( \16556 , \16468 , \16485 );
and \U$16425 ( \16557 , \16424 , \16485 );
or \U$16426 ( \16558 , \16555 , \16556 , \16557 );
xor \U$16427 ( \16559 , \16554 , \16558 );
xor \U$16428 ( \16560 , \16545 , \16559 );
and \U$16429 ( \16561 , \16394 , \16408 );
and \U$16430 ( \16562 , \16408 , \16423 );
and \U$16431 ( \16563 , \16394 , \16423 );
or \U$16432 ( \16564 , \16561 , \16562 , \16563 );
and \U$16433 ( \16565 , \16438 , \16452 );
and \U$16434 ( \16566 , \16452 , \16467 );
and \U$16435 ( \16567 , \16438 , \16467 );
or \U$16436 ( \16568 , \16565 , \16566 , \16567 );
xor \U$16437 ( \16569 , \16564 , \16568 );
and \U$16438 ( \16570 , \8835 , \2121 );
and \U$16439 ( \16571 , \9169 , \2008 );
nor \U$16440 ( \16572 , \16570 , \16571 );
xnor \U$16441 ( \16573 , \16572 , \1961 );
and \U$16442 ( \16574 , \8349 , \2400 );
and \U$16443 ( \16575 , \8652 , \2246 );
nor \U$16444 ( \16576 , \16574 , \16575 );
xnor \U$16445 ( \16577 , \16576 , \2195 );
xor \U$16446 ( \16578 , \16573 , \16577 );
and \U$16447 ( \16579 , \7700 , \2669 );
and \U$16448 ( \16580 , \8057 , \2538 );
nor \U$16449 ( \16581 , \16579 , \16580 );
xnor \U$16450 ( \16582 , \16581 , \2534 );
xor \U$16451 ( \16583 , \16578 , \16582 );
xor \U$16452 ( \16584 , \16569 , \16583 );
and \U$16453 ( \16585 , \16368 , \16372 );
and \U$16454 ( \16586 , \16372 , \16377 );
and \U$16455 ( \16587 , \16368 , \16377 );
or \U$16456 ( \16588 , \16585 , \16586 , \16587 );
and \U$16457 ( \16589 , \16442 , \16446 );
and \U$16458 ( \16590 , \16446 , \16451 );
and \U$16459 ( \16591 , \16442 , \16451 );
or \U$16460 ( \16592 , \16589 , \16590 , \16591 );
xor \U$16461 ( \16593 , \16588 , \16592 );
and \U$16462 ( \16594 , \16457 , \16461 );
and \U$16463 ( \16595 , \16461 , \16466 );
and \U$16464 ( \16596 , \16457 , \16466 );
or \U$16465 ( \16597 , \16594 , \16595 , \16596 );
xor \U$16466 ( \16598 , \16593 , \16597 );
and \U$16467 ( \16599 , \16384 , \16388 );
and \U$16468 ( \16600 , \16388 , \16393 );
and \U$16469 ( \16601 , \16384 , \16393 );
or \U$16470 ( \16602 , \16599 , \16600 , \16601 );
or \U$16471 ( \16603 , \16482 , \16483 );
xor \U$16472 ( \16604 , \16602 , \16603 );
and \U$16473 ( \16605 , \1484 , \10408 );
and \U$16474 ( \16606 , \1601 , \10116 );
nor \U$16475 ( \16607 , \16605 , \16606 );
xnor \U$16476 ( \16608 , \16607 , \10121 );
xor \U$16477 ( \16609 , \16604 , \16608 );
xor \U$16478 ( \16610 , \16598 , \16609 );
and \U$16479 ( \16611 , \16428 , \16432 );
and \U$16480 ( \16612 , \16432 , \16437 );
and \U$16481 ( \16613 , \16428 , \16437 );
or \U$16482 ( \16614 , \16611 , \16612 , \16613 );
and \U$16483 ( \16615 , \16398 , \16402 );
and \U$16484 ( \16616 , \16402 , \16407 );
and \U$16485 ( \16617 , \16398 , \16407 );
or \U$16486 ( \16618 , \16615 , \16616 , \16617 );
xor \U$16487 ( \16619 , \16614 , \16618 );
and \U$16488 ( \16620 , \16413 , \16417 );
and \U$16489 ( \16621 , \16417 , \16422 );
and \U$16490 ( \16622 , \16413 , \16422 );
or \U$16491 ( \16623 , \16620 , \16621 , \16622 );
xor \U$16492 ( \16624 , \16619 , \16623 );
xor \U$16493 ( \16625 , \16610 , \16624 );
xor \U$16494 ( \16626 , \16584 , \16625 );
not \U$16495 ( \16627 , \1205 );
and \U$16496 ( \16628 , \10206 , \1578 );
and \U$16497 ( \16629 , \10584 , \1431 );
nor \U$16498 ( \16630 , \16628 , \16629 );
xnor \U$16499 ( \16631 , \16630 , \1436 );
xor \U$16500 ( \16632 , \16627 , \16631 );
and \U$16501 ( \16633 , \9465 , \1824 );
and \U$16502 ( \16634 , \9897 , \1739 );
nor \U$16503 ( \16635 , \16633 , \16634 );
xnor \U$16504 ( \16636 , \16635 , \1697 );
xor \U$16505 ( \16637 , \16632 , \16636 );
and \U$16506 ( \16638 , \1333 , \10118 );
and \U$16507 ( \16639 , \2182 , \8540 );
and \U$16508 ( \16640 , \2366 , \8292 );
nor \U$16509 ( \16641 , \16639 , \16640 );
xnor \U$16510 ( \16642 , \16641 , \8297 );
and \U$16511 ( \16643 , \1948 , \9333 );
and \U$16512 ( \16644 , \2090 , \9006 );
nor \U$16513 ( \16645 , \16643 , \16644 );
xnor \U$16514 ( \16646 , \16645 , \8848 );
xor \U$16515 ( \16647 , \16642 , \16646 );
and \U$16516 ( \16648 , \1684 , \9765 );
and \U$16517 ( \16649 , \1802 , \9644 );
nor \U$16518 ( \16650 , \16648 , \16649 );
xnor \U$16519 ( \16651 , \16650 , \9478 );
xor \U$16520 ( \16652 , \16647 , \16651 );
xor \U$16521 ( \16653 , \16638 , \16652 );
and \U$16522 ( \16654 , \3143 , \7055 );
and \U$16523 ( \16655 , \3395 , \6675 );
nor \U$16524 ( \16656 , \16654 , \16655 );
xnor \U$16525 ( \16657 , \16656 , \6680 );
and \U$16526 ( \16658 , \2826 , \7489 );
and \U$16527 ( \16659 , \3037 , \7137 );
nor \U$16528 ( \16660 , \16658 , \16659 );
xnor \U$16529 ( \16661 , \16660 , \7142 );
xor \U$16530 ( \16662 , \16657 , \16661 );
and \U$16531 ( \16663 , \2521 , \8019 );
and \U$16532 ( \16664 , \2757 , \7830 );
nor \U$16533 ( \16665 , \16663 , \16664 );
xnor \U$16534 ( \16666 , \16665 , \7713 );
xor \U$16535 ( \16667 , \16662 , \16666 );
xor \U$16536 ( \16668 , \16653 , \16667 );
xor \U$16537 ( \16669 , \16637 , \16668 );
and \U$16538 ( \16670 , \5674 , \4132 );
and \U$16539 ( \16671 , \6030 , \4012 );
nor \U$16540 ( \16672 , \16670 , \16671 );
xnor \U$16541 ( \16673 , \16672 , \3925 );
and \U$16542 ( \16674 , \5156 , \4581 );
and \U$16543 ( \16675 , \5469 , \4424 );
nor \U$16544 ( \16676 , \16674 , \16675 );
xnor \U$16545 ( \16677 , \16676 , \4377 );
xor \U$16546 ( \16678 , \16673 , \16677 );
and \U$16547 ( \16679 , \4749 , \5011 );
and \U$16548 ( \16680 , \4922 , \4878 );
nor \U$16549 ( \16681 , \16679 , \16680 );
xnor \U$16550 ( \16682 , \16681 , \4762 );
xor \U$16551 ( \16683 , \16678 , \16682 );
and \U$16552 ( \16684 , \7231 , \3103 );
and \U$16553 ( \16685 , \7556 , \2934 );
nor \U$16554 ( \16686 , \16684 , \16685 );
xnor \U$16555 ( \16687 , \16686 , \2839 );
and \U$16556 ( \16688 , \6790 , \3357 );
and \U$16557 ( \16689 , \6945 , \3255 );
nor \U$16558 ( \16690 , \16688 , \16689 );
xnor \U$16559 ( \16691 , \16690 , \3156 );
xor \U$16560 ( \16692 , \16687 , \16691 );
and \U$16561 ( \16693 , \6281 , \3813 );
and \U$16562 ( \16694 , \6514 , \3557 );
nor \U$16563 ( \16695 , \16693 , \16694 );
xnor \U$16564 ( \16696 , \16695 , \3562 );
xor \U$16565 ( \16697 , \16692 , \16696 );
xor \U$16566 ( \16698 , \16683 , \16697 );
and \U$16567 ( \16699 , \4364 , \5485 );
and \U$16568 ( \16700 , \4654 , \5275 );
nor \U$16569 ( \16701 , \16699 , \16700 );
xnor \U$16570 ( \16702 , \16701 , \5169 );
and \U$16571 ( \16703 , \3912 , \5996 );
and \U$16572 ( \16704 , \4160 , \5695 );
nor \U$16573 ( \16705 , \16703 , \16704 );
xnor \U$16574 ( \16706 , \16705 , \5687 );
xor \U$16575 ( \16707 , \16702 , \16706 );
and \U$16576 ( \16708 , \3646 , \6401 );
and \U$16577 ( \16709 , \3736 , \6143 );
nor \U$16578 ( \16710 , \16708 , \16709 );
xnor \U$16579 ( \16711 , \16710 , \6148 );
xor \U$16580 ( \16712 , \16707 , \16711 );
xor \U$16581 ( \16713 , \16698 , \16712 );
xor \U$16582 ( \16714 , \16669 , \16713 );
xor \U$16583 ( \16715 , \16626 , \16714 );
xor \U$16584 ( \16716 , \16560 , \16715 );
xor \U$16585 ( \16717 , \16531 , \16716 );
xor \U$16586 ( \16718 , \16522 , \16717 );
xor \U$16587 ( \16719 , \16503 , \16718 );
and \U$16588 ( \16720 , \16268 , \16490 );
xor \U$16589 ( \16721 , \16719 , \16720 );
and \U$16590 ( \16722 , \16491 , \16492 );
and \U$16591 ( \16723 , \16493 , \16496 );
or \U$16592 ( \16724 , \16722 , \16723 );
xor \U$16593 ( \16725 , \16721 , \16724 );
buf \U$16594 ( \16726 , \16725 );
buf \U$16595 ( \16727 , \16726 );
and \U$16596 ( \16728 , \16507 , \16521 );
and \U$16597 ( \16729 , \16521 , \16717 );
and \U$16598 ( \16730 , \16507 , \16717 );
or \U$16599 ( \16731 , \16728 , \16729 , \16730 );
and \U$16600 ( \16732 , \16526 , \16530 );
and \U$16601 ( \16733 , \16530 , \16716 );
and \U$16602 ( \16734 , \16526 , \16716 );
or \U$16603 ( \16735 , \16732 , \16733 , \16734 );
and \U$16604 ( \16736 , \16549 , \16553 );
and \U$16605 ( \16737 , \16553 , \16558 );
and \U$16606 ( \16738 , \16549 , \16558 );
or \U$16607 ( \16739 , \16736 , \16737 , \16738 );
and \U$16608 ( \16740 , \16584 , \16625 );
and \U$16609 ( \16741 , \16625 , \16714 );
and \U$16610 ( \16742 , \16584 , \16714 );
or \U$16611 ( \16743 , \16740 , \16741 , \16742 );
xor \U$16612 ( \16744 , \16739 , \16743 );
and \U$16613 ( \16745 , \16638 , \16652 );
and \U$16614 ( \16746 , \16652 , \16667 );
and \U$16615 ( \16747 , \16638 , \16667 );
or \U$16616 ( \16748 , \16745 , \16746 , \16747 );
and \U$16617 ( \16749 , \16683 , \16697 );
and \U$16618 ( \16750 , \16697 , \16712 );
and \U$16619 ( \16751 , \16683 , \16712 );
or \U$16620 ( \16752 , \16749 , \16750 , \16751 );
xor \U$16621 ( \16753 , \16748 , \16752 );
and \U$16622 ( \16754 , \6945 , \3357 );
and \U$16623 ( \16755 , \7231 , \3255 );
nor \U$16624 ( \16756 , \16754 , \16755 );
xnor \U$16625 ( \16757 , \16756 , \3156 );
and \U$16626 ( \16758 , \6514 , \3813 );
and \U$16627 ( \16759 , \6790 , \3557 );
nor \U$16628 ( \16760 , \16758 , \16759 );
xnor \U$16629 ( \16761 , \16760 , \3562 );
xor \U$16630 ( \16762 , \16757 , \16761 );
and \U$16631 ( \16763 , \6030 , \4132 );
and \U$16632 ( \16764 , \6281 , \4012 );
nor \U$16633 ( \16765 , \16763 , \16764 );
xnor \U$16634 ( \16766 , \16765 , \3925 );
xor \U$16635 ( \16767 , \16762 , \16766 );
and \U$16636 ( \16768 , \10584 , \1578 );
not \U$16637 ( \16769 , \16768 );
xnor \U$16638 ( \16770 , \16769 , \1436 );
and \U$16639 ( \16771 , \9897 , \1824 );
and \U$16640 ( \16772 , \10206 , \1739 );
nor \U$16641 ( \16773 , \16771 , \16772 );
xnor \U$16642 ( \16774 , \16773 , \1697 );
xor \U$16643 ( \16775 , \16770 , \16774 );
and \U$16644 ( \16776 , \9169 , \2121 );
and \U$16645 ( \16777 , \9465 , \2008 );
nor \U$16646 ( \16778 , \16776 , \16777 );
xnor \U$16647 ( \16779 , \16778 , \1961 );
xor \U$16648 ( \16780 , \16775 , \16779 );
xor \U$16649 ( \16781 , \16767 , \16780 );
and \U$16650 ( \16782 , \8652 , \2400 );
and \U$16651 ( \16783 , \8835 , \2246 );
nor \U$16652 ( \16784 , \16782 , \16783 );
xnor \U$16653 ( \16785 , \16784 , \2195 );
and \U$16654 ( \16786 , \8057 , \2669 );
and \U$16655 ( \16787 , \8349 , \2538 );
nor \U$16656 ( \16788 , \16786 , \16787 );
xnor \U$16657 ( \16789 , \16788 , \2534 );
xor \U$16658 ( \16790 , \16785 , \16789 );
and \U$16659 ( \16791 , \7556 , \3103 );
and \U$16660 ( \16792 , \7700 , \2934 );
nor \U$16661 ( \16793 , \16791 , \16792 );
xnor \U$16662 ( \16794 , \16793 , \2839 );
xor \U$16663 ( \16795 , \16790 , \16794 );
xor \U$16664 ( \16796 , \16781 , \16795 );
xor \U$16665 ( \16797 , \16753 , \16796 );
xor \U$16666 ( \16798 , \16744 , \16797 );
xor \U$16667 ( \16799 , \16735 , \16798 );
and \U$16668 ( \16800 , \16511 , \16515 );
and \U$16669 ( \16801 , \16515 , \16520 );
and \U$16670 ( \16802 , \16511 , \16520 );
or \U$16671 ( \16803 , \16800 , \16801 , \16802 );
and \U$16672 ( \16804 , \16545 , \16559 );
and \U$16673 ( \16805 , \16559 , \16715 );
and \U$16674 ( \16806 , \16545 , \16715 );
or \U$16675 ( \16807 , \16804 , \16805 , \16806 );
xor \U$16676 ( \16808 , \16803 , \16807 );
and \U$16677 ( \16809 , \16588 , \16592 );
and \U$16678 ( \16810 , \16592 , \16597 );
and \U$16679 ( \16811 , \16588 , \16597 );
or \U$16680 ( \16812 , \16809 , \16810 , \16811 );
and \U$16681 ( \16813 , \16602 , \16603 );
and \U$16682 ( \16814 , \16603 , \16608 );
and \U$16683 ( \16815 , \16602 , \16608 );
or \U$16684 ( \16816 , \16813 , \16814 , \16815 );
xor \U$16685 ( \16817 , \16812 , \16816 );
and \U$16686 ( \16818 , \16614 , \16618 );
and \U$16687 ( \16819 , \16618 , \16623 );
and \U$16688 ( \16820 , \16614 , \16623 );
or \U$16689 ( \16821 , \16818 , \16819 , \16820 );
xor \U$16690 ( \16822 , \16817 , \16821 );
and \U$16691 ( \16823 , \16535 , \16539 );
and \U$16692 ( \16824 , \16539 , \16544 );
and \U$16693 ( \16825 , \16535 , \16544 );
or \U$16694 ( \16826 , \16823 , \16824 , \16825 );
and \U$16695 ( \16827 , \16564 , \16568 );
and \U$16696 ( \16828 , \16568 , \16583 );
and \U$16697 ( \16829 , \16564 , \16583 );
or \U$16698 ( \16830 , \16827 , \16828 , \16829 );
xor \U$16699 ( \16831 , \16826 , \16830 );
and \U$16700 ( \16832 , \16637 , \16668 );
and \U$16701 ( \16833 , \16668 , \16713 );
and \U$16702 ( \16834 , \16637 , \16713 );
or \U$16703 ( \16835 , \16832 , \16833 , \16834 );
xor \U$16704 ( \16836 , \16831 , \16835 );
xor \U$16705 ( \16837 , \16822 , \16836 );
and \U$16706 ( \16838 , \16598 , \16609 );
and \U$16707 ( \16839 , \16609 , \16624 );
and \U$16708 ( \16840 , \16598 , \16624 );
or \U$16709 ( \16841 , \16838 , \16839 , \16840 );
and \U$16710 ( \16842 , \16687 , \16691 );
and \U$16711 ( \16843 , \16691 , \16696 );
and \U$16712 ( \16844 , \16687 , \16696 );
or \U$16713 ( \16845 , \16842 , \16843 , \16844 );
and \U$16714 ( \16846 , \16627 , \16631 );
and \U$16715 ( \16847 , \16631 , \16636 );
and \U$16716 ( \16848 , \16627 , \16636 );
or \U$16717 ( \16849 , \16846 , \16847 , \16848 );
xor \U$16718 ( \16850 , \16845 , \16849 );
and \U$16719 ( \16851 , \16573 , \16577 );
and \U$16720 ( \16852 , \16577 , \16582 );
and \U$16721 ( \16853 , \16573 , \16582 );
or \U$16722 ( \16854 , \16851 , \16852 , \16853 );
xor \U$16723 ( \16855 , \16850 , \16854 );
xor \U$16724 ( \16856 , \16841 , \16855 );
and \U$16725 ( \16857 , \16673 , \16677 );
and \U$16726 ( \16858 , \16677 , \16682 );
and \U$16727 ( \16859 , \16673 , \16682 );
or \U$16728 ( \16860 , \16857 , \16858 , \16859 );
and \U$16729 ( \16861 , \16657 , \16661 );
and \U$16730 ( \16862 , \16661 , \16666 );
and \U$16731 ( \16863 , \16657 , \16666 );
or \U$16732 ( \16864 , \16861 , \16862 , \16863 );
xor \U$16733 ( \16865 , \16860 , \16864 );
and \U$16734 ( \16866 , \16702 , \16706 );
and \U$16735 ( \16867 , \16706 , \16711 );
and \U$16736 ( \16868 , \16702 , \16711 );
or \U$16737 ( \16869 , \16866 , \16867 , \16868 );
xor \U$16738 ( \16870 , \16865 , \16869 );
and \U$16739 ( \16871 , \3037 , \7489 );
and \U$16740 ( \16872 , \3143 , \7137 );
nor \U$16741 ( \16873 , \16871 , \16872 );
xnor \U$16742 ( \16874 , \16873 , \7142 );
and \U$16743 ( \16875 , \2757 , \8019 );
and \U$16744 ( \16876 , \2826 , \7830 );
nor \U$16745 ( \16877 , \16875 , \16876 );
xnor \U$16746 ( \16878 , \16877 , \7713 );
xor \U$16747 ( \16879 , \16874 , \16878 );
and \U$16748 ( \16880 , \2366 , \8540 );
and \U$16749 ( \16881 , \2521 , \8292 );
nor \U$16750 ( \16882 , \16880 , \16881 );
xnor \U$16751 ( \16883 , \16882 , \8297 );
xor \U$16752 ( \16884 , \16879 , \16883 );
and \U$16753 ( \16885 , \4160 , \5996 );
and \U$16754 ( \16886 , \4364 , \5695 );
nor \U$16755 ( \16887 , \16885 , \16886 );
xnor \U$16756 ( \16888 , \16887 , \5687 );
and \U$16757 ( \16889 , \3736 , \6401 );
and \U$16758 ( \16890 , \3912 , \6143 );
nor \U$16759 ( \16891 , \16889 , \16890 );
xnor \U$16760 ( \16892 , \16891 , \6148 );
xor \U$16761 ( \16893 , \16888 , \16892 );
and \U$16762 ( \16894 , \3395 , \7055 );
and \U$16763 ( \16895 , \3646 , \6675 );
nor \U$16764 ( \16896 , \16894 , \16895 );
xnor \U$16765 ( \16897 , \16896 , \6680 );
xor \U$16766 ( \16898 , \16893 , \16897 );
xor \U$16767 ( \16899 , \16884 , \16898 );
and \U$16768 ( \16900 , \5469 , \4581 );
and \U$16769 ( \16901 , \5674 , \4424 );
nor \U$16770 ( \16902 , \16900 , \16901 );
xnor \U$16771 ( \16903 , \16902 , \4377 );
and \U$16772 ( \16904 , \4922 , \5011 );
and \U$16773 ( \16905 , \5156 , \4878 );
nor \U$16774 ( \16906 , \16904 , \16905 );
xnor \U$16775 ( \16907 , \16906 , \4762 );
xor \U$16776 ( \16908 , \16903 , \16907 );
and \U$16777 ( \16909 , \4654 , \5485 );
and \U$16778 ( \16910 , \4749 , \5275 );
nor \U$16779 ( \16911 , \16909 , \16910 );
xnor \U$16780 ( \16912 , \16911 , \5169 );
xor \U$16781 ( \16913 , \16908 , \16912 );
xor \U$16782 ( \16914 , \16899 , \16913 );
xor \U$16783 ( \16915 , \16870 , \16914 );
and \U$16784 ( \16916 , \16642 , \16646 );
and \U$16785 ( \16917 , \16646 , \16651 );
and \U$16786 ( \16918 , \16642 , \16651 );
or \U$16787 ( \16919 , \16916 , \16917 , \16918 );
and \U$16788 ( \16920 , \2090 , \9333 );
and \U$16789 ( \16921 , \2182 , \9006 );
nor \U$16790 ( \16922 , \16920 , \16921 );
xnor \U$16791 ( \16923 , \16922 , \8848 );
and \U$16792 ( \16924 , \1802 , \9765 );
and \U$16793 ( \16925 , \1948 , \9644 );
nor \U$16794 ( \16926 , \16924 , \16925 );
xnor \U$16795 ( \16927 , \16926 , \9478 );
xor \U$16796 ( \16928 , \16923 , \16927 );
and \U$16797 ( \16929 , \1601 , \10408 );
and \U$16798 ( \16930 , \1684 , \10116 );
nor \U$16799 ( \16931 , \16929 , \16930 );
xnor \U$16800 ( \16932 , \16931 , \10121 );
xor \U$16801 ( \16933 , \16928 , \16932 );
xor \U$16802 ( \16934 , \16919 , \16933 );
and \U$16803 ( \16935 , \1484 , \10118 );
not \U$16804 ( \16936 , \16935 );
xor \U$16805 ( \16937 , \16934 , \16936 );
xor \U$16806 ( \16938 , \16915 , \16937 );
xor \U$16807 ( \16939 , \16856 , \16938 );
xor \U$16808 ( \16940 , \16837 , \16939 );
xor \U$16809 ( \16941 , \16808 , \16940 );
xor \U$16810 ( \16942 , \16799 , \16941 );
xor \U$16811 ( \16943 , \16731 , \16942 );
and \U$16812 ( \16944 , \16503 , \16718 );
xor \U$16813 ( \16945 , \16943 , \16944 );
and \U$16814 ( \16946 , \16719 , \16720 );
and \U$16815 ( \16947 , \16721 , \16724 );
or \U$16816 ( \16948 , \16946 , \16947 );
xor \U$16817 ( \16949 , \16945 , \16948 );
buf \U$16818 ( \16950 , \16949 );
buf \U$16819 ( \16951 , \16950 );
and \U$16820 ( \16952 , \16735 , \16798 );
and \U$16821 ( \16953 , \16798 , \16941 );
and \U$16822 ( \16954 , \16735 , \16941 );
or \U$16823 ( \16955 , \16952 , \16953 , \16954 );
and \U$16824 ( \16956 , \16803 , \16807 );
and \U$16825 ( \16957 , \16807 , \16940 );
and \U$16826 ( \16958 , \16803 , \16940 );
or \U$16827 ( \16959 , \16956 , \16957 , \16958 );
and \U$16828 ( \16960 , \16826 , \16830 );
and \U$16829 ( \16961 , \16830 , \16835 );
and \U$16830 ( \16962 , \16826 , \16835 );
or \U$16831 ( \16963 , \16960 , \16961 , \16962 );
and \U$16832 ( \16964 , \16841 , \16855 );
and \U$16833 ( \16965 , \16855 , \16938 );
and \U$16834 ( \16966 , \16841 , \16938 );
or \U$16835 ( \16967 , \16964 , \16965 , \16966 );
xor \U$16836 ( \16968 , \16963 , \16967 );
and \U$16837 ( \16969 , \16884 , \16898 );
and \U$16838 ( \16970 , \16898 , \16913 );
and \U$16839 ( \16971 , \16884 , \16913 );
or \U$16840 ( \16972 , \16969 , \16970 , \16971 );
and \U$16841 ( \16973 , \16767 , \16780 );
and \U$16842 ( \16974 , \16780 , \16795 );
and \U$16843 ( \16975 , \16767 , \16795 );
or \U$16844 ( \16976 , \16973 , \16974 , \16975 );
xor \U$16845 ( \16977 , \16972 , \16976 );
not \U$16846 ( \16978 , \1436 );
and \U$16847 ( \16979 , \10206 , \1824 );
and \U$16848 ( \16980 , \10584 , \1739 );
nor \U$16849 ( \16981 , \16979 , \16980 );
xnor \U$16850 ( \16982 , \16981 , \1697 );
xor \U$16851 ( \16983 , \16978 , \16982 );
and \U$16852 ( \16984 , \9465 , \2121 );
and \U$16853 ( \16985 , \9897 , \2008 );
nor \U$16854 ( \16986 , \16984 , \16985 );
xnor \U$16855 ( \16987 , \16986 , \1961 );
xor \U$16856 ( \16988 , \16983 , \16987 );
xor \U$16857 ( \16989 , \16977 , \16988 );
xor \U$16858 ( \16990 , \16968 , \16989 );
xor \U$16859 ( \16991 , \16959 , \16990 );
and \U$16860 ( \16992 , \16739 , \16743 );
and \U$16861 ( \16993 , \16743 , \16797 );
and \U$16862 ( \16994 , \16739 , \16797 );
or \U$16863 ( \16995 , \16992 , \16993 , \16994 );
and \U$16864 ( \16996 , \16822 , \16836 );
and \U$16865 ( \16997 , \16836 , \16939 );
and \U$16866 ( \16998 , \16822 , \16939 );
or \U$16867 ( \16999 , \16996 , \16997 , \16998 );
xor \U$16868 ( \17000 , \16995 , \16999 );
and \U$16869 ( \17001 , \16845 , \16849 );
and \U$16870 ( \17002 , \16849 , \16854 );
and \U$16871 ( \17003 , \16845 , \16854 );
or \U$16872 ( \17004 , \17001 , \17002 , \17003 );
and \U$16873 ( \17005 , \16860 , \16864 );
and \U$16874 ( \17006 , \16864 , \16869 );
and \U$16875 ( \17007 , \16860 , \16869 );
or \U$16876 ( \17008 , \17005 , \17006 , \17007 );
xor \U$16877 ( \17009 , \17004 , \17008 );
and \U$16878 ( \17010 , \16919 , \16933 );
and \U$16879 ( \17011 , \16933 , \16936 );
and \U$16880 ( \17012 , \16919 , \16936 );
or \U$16881 ( \17013 , \17010 , \17011 , \17012 );
xor \U$16882 ( \17014 , \17009 , \17013 );
and \U$16883 ( \17015 , \16812 , \16816 );
and \U$16884 ( \17016 , \16816 , \16821 );
and \U$16885 ( \17017 , \16812 , \16821 );
or \U$16886 ( \17018 , \17015 , \17016 , \17017 );
and \U$16887 ( \17019 , \16748 , \16752 );
and \U$16888 ( \17020 , \16752 , \16796 );
and \U$16889 ( \17021 , \16748 , \16796 );
or \U$16890 ( \17022 , \17019 , \17020 , \17021 );
xor \U$16891 ( \17023 , \17018 , \17022 );
and \U$16892 ( \17024 , \16870 , \16914 );
and \U$16893 ( \17025 , \16914 , \16937 );
and \U$16894 ( \17026 , \16870 , \16937 );
or \U$16895 ( \17027 , \17024 , \17025 , \17026 );
xor \U$16896 ( \17028 , \17023 , \17027 );
xor \U$16897 ( \17029 , \17014 , \17028 );
and \U$16898 ( \17030 , \16757 , \16761 );
and \U$16899 ( \17031 , \16761 , \16766 );
and \U$16900 ( \17032 , \16757 , \16766 );
or \U$16901 ( \17033 , \17030 , \17031 , \17032 );
and \U$16902 ( \17034 , \16770 , \16774 );
and \U$16903 ( \17035 , \16774 , \16779 );
and \U$16904 ( \17036 , \16770 , \16779 );
or \U$16905 ( \17037 , \17034 , \17035 , \17036 );
xor \U$16906 ( \17038 , \17033 , \17037 );
and \U$16907 ( \17039 , \16785 , \16789 );
and \U$16908 ( \17040 , \16789 , \16794 );
and \U$16909 ( \17041 , \16785 , \16794 );
or \U$16910 ( \17042 , \17039 , \17040 , \17041 );
xor \U$16911 ( \17043 , \17038 , \17042 );
and \U$16912 ( \17044 , \16874 , \16878 );
and \U$16913 ( \17045 , \16878 , \16883 );
and \U$16914 ( \17046 , \16874 , \16883 );
or \U$16915 ( \17047 , \17044 , \17045 , \17046 );
and \U$16916 ( \17048 , \16888 , \16892 );
and \U$16917 ( \17049 , \16892 , \16897 );
and \U$16918 ( \17050 , \16888 , \16897 );
or \U$16919 ( \17051 , \17048 , \17049 , \17050 );
xor \U$16920 ( \17052 , \17047 , \17051 );
and \U$16921 ( \17053 , \16903 , \16907 );
and \U$16922 ( \17054 , \16907 , \16912 );
and \U$16923 ( \17055 , \16903 , \16912 );
or \U$16924 ( \17056 , \17053 , \17054 , \17055 );
xor \U$16925 ( \17057 , \17052 , \17056 );
xor \U$16926 ( \17058 , \17043 , \17057 );
and \U$16927 ( \17059 , \16923 , \16927 );
and \U$16928 ( \17060 , \16927 , \16932 );
and \U$16929 ( \17061 , \16923 , \16932 );
or \U$16930 ( \17062 , \17059 , \17060 , \17061 );
buf \U$16931 ( \17063 , \16935 );
xor \U$16932 ( \17064 , \17062 , \17063 );
and \U$16933 ( \17065 , \1601 , \10118 );
xor \U$16934 ( \17066 , \17064 , \17065 );
and \U$16935 ( \17067 , \3143 , \7489 );
and \U$16936 ( \17068 , \3395 , \7137 );
nor \U$16937 ( \17069 , \17067 , \17068 );
xnor \U$16938 ( \17070 , \17069 , \7142 );
and \U$16939 ( \17071 , \2826 , \8019 );
and \U$16940 ( \17072 , \3037 , \7830 );
nor \U$16941 ( \17073 , \17071 , \17072 );
xnor \U$16942 ( \17074 , \17073 , \7713 );
xor \U$16943 ( \17075 , \17070 , \17074 );
and \U$16944 ( \17076 , \2521 , \8540 );
and \U$16945 ( \17077 , \2757 , \8292 );
nor \U$16946 ( \17078 , \17076 , \17077 );
xnor \U$16947 ( \17079 , \17078 , \8297 );
xor \U$16948 ( \17080 , \17075 , \17079 );
and \U$16949 ( \17081 , \4364 , \5996 );
and \U$16950 ( \17082 , \4654 , \5695 );
nor \U$16951 ( \17083 , \17081 , \17082 );
xnor \U$16952 ( \17084 , \17083 , \5687 );
and \U$16953 ( \17085 , \3912 , \6401 );
and \U$16954 ( \17086 , \4160 , \6143 );
nor \U$16955 ( \17087 , \17085 , \17086 );
xnor \U$16956 ( \17088 , \17087 , \6148 );
xor \U$16957 ( \17089 , \17084 , \17088 );
and \U$16958 ( \17090 , \3646 , \7055 );
and \U$16959 ( \17091 , \3736 , \6675 );
nor \U$16960 ( \17092 , \17090 , \17091 );
xnor \U$16961 ( \17093 , \17092 , \6680 );
xor \U$16962 ( \17094 , \17089 , \17093 );
xor \U$16963 ( \17095 , \17080 , \17094 );
and \U$16964 ( \17096 , \2182 , \9333 );
and \U$16965 ( \17097 , \2366 , \9006 );
nor \U$16966 ( \17098 , \17096 , \17097 );
xnor \U$16967 ( \17099 , \17098 , \8848 );
and \U$16968 ( \17100 , \1948 , \9765 );
and \U$16969 ( \17101 , \2090 , \9644 );
nor \U$16970 ( \17102 , \17100 , \17101 );
xnor \U$16971 ( \17103 , \17102 , \9478 );
xor \U$16972 ( \17104 , \17099 , \17103 );
and \U$16973 ( \17105 , \1684 , \10408 );
and \U$16974 ( \17106 , \1802 , \10116 );
nor \U$16975 ( \17107 , \17105 , \17106 );
xnor \U$16976 ( \17108 , \17107 , \10121 );
xor \U$16977 ( \17109 , \17104 , \17108 );
xor \U$16978 ( \17110 , \17095 , \17109 );
xor \U$16979 ( \17111 , \17066 , \17110 );
and \U$16980 ( \17112 , \7231 , \3357 );
and \U$16981 ( \17113 , \7556 , \3255 );
nor \U$16982 ( \17114 , \17112 , \17113 );
xnor \U$16983 ( \17115 , \17114 , \3156 );
and \U$16984 ( \17116 , \6790 , \3813 );
and \U$16985 ( \17117 , \6945 , \3557 );
nor \U$16986 ( \17118 , \17116 , \17117 );
xnor \U$16987 ( \17119 , \17118 , \3562 );
xor \U$16988 ( \17120 , \17115 , \17119 );
and \U$16989 ( \17121 , \6281 , \4132 );
and \U$16990 ( \17122 , \6514 , \4012 );
nor \U$16991 ( \17123 , \17121 , \17122 );
xnor \U$16992 ( \17124 , \17123 , \3925 );
xor \U$16993 ( \17125 , \17120 , \17124 );
and \U$16994 ( \17126 , \5674 , \4581 );
and \U$16995 ( \17127 , \6030 , \4424 );
nor \U$16996 ( \17128 , \17126 , \17127 );
xnor \U$16997 ( \17129 , \17128 , \4377 );
and \U$16998 ( \17130 , \5156 , \5011 );
and \U$16999 ( \17131 , \5469 , \4878 );
nor \U$17000 ( \17132 , \17130 , \17131 );
xnor \U$17001 ( \17133 , \17132 , \4762 );
xor \U$17002 ( \17134 , \17129 , \17133 );
and \U$17003 ( \17135 , \4749 , \5485 );
and \U$17004 ( \17136 , \4922 , \5275 );
nor \U$17005 ( \17137 , \17135 , \17136 );
xnor \U$17006 ( \17138 , \17137 , \5169 );
xor \U$17007 ( \17139 , \17134 , \17138 );
xor \U$17008 ( \17140 , \17125 , \17139 );
and \U$17009 ( \17141 , \8835 , \2400 );
and \U$17010 ( \17142 , \9169 , \2246 );
nor \U$17011 ( \17143 , \17141 , \17142 );
xnor \U$17012 ( \17144 , \17143 , \2195 );
and \U$17013 ( \17145 , \8349 , \2669 );
and \U$17014 ( \17146 , \8652 , \2538 );
nor \U$17015 ( \17147 , \17145 , \17146 );
xnor \U$17016 ( \17148 , \17147 , \2534 );
xor \U$17017 ( \17149 , \17144 , \17148 );
and \U$17018 ( \17150 , \7700 , \3103 );
and \U$17019 ( \17151 , \8057 , \2934 );
nor \U$17020 ( \17152 , \17150 , \17151 );
xnor \U$17021 ( \17153 , \17152 , \2839 );
xor \U$17022 ( \17154 , \17149 , \17153 );
xor \U$17023 ( \17155 , \17140 , \17154 );
xor \U$17024 ( \17156 , \17111 , \17155 );
xor \U$17025 ( \17157 , \17058 , \17156 );
xor \U$17026 ( \17158 , \17029 , \17157 );
xor \U$17027 ( \17159 , \17000 , \17158 );
xor \U$17028 ( \17160 , \16991 , \17159 );
xor \U$17029 ( \17161 , \16955 , \17160 );
and \U$17030 ( \17162 , \16731 , \16942 );
xor \U$17031 ( \17163 , \17161 , \17162 );
and \U$17032 ( \17164 , \16943 , \16944 );
and \U$17033 ( \17165 , \16945 , \16948 );
or \U$17034 ( \17166 , \17164 , \17165 );
xor \U$17035 ( \17167 , \17163 , \17166 );
buf \U$17036 ( \17168 , \17167 );
buf \U$17037 ( \17169 , \17168 );
and \U$17038 ( \17170 , \16959 , \16990 );
and \U$17039 ( \17171 , \16990 , \17159 );
and \U$17040 ( \17172 , \16959 , \17159 );
or \U$17041 ( \17173 , \17170 , \17171 , \17172 );
and \U$17042 ( \17174 , \16995 , \16999 );
and \U$17043 ( \17175 , \16999 , \17158 );
and \U$17044 ( \17176 , \16995 , \17158 );
or \U$17045 ( \17177 , \17174 , \17175 , \17176 );
and \U$17046 ( \17178 , \16963 , \16967 );
and \U$17047 ( \17179 , \16967 , \16989 );
and \U$17048 ( \17180 , \16963 , \16989 );
or \U$17049 ( \17181 , \17178 , \17179 , \17180 );
and \U$17050 ( \17182 , \17014 , \17028 );
and \U$17051 ( \17183 , \17028 , \17157 );
and \U$17052 ( \17184 , \17014 , \17157 );
or \U$17053 ( \17185 , \17182 , \17183 , \17184 );
xor \U$17054 ( \17186 , \17181 , \17185 );
and \U$17055 ( \17187 , \17115 , \17119 );
and \U$17056 ( \17188 , \17119 , \17124 );
and \U$17057 ( \17189 , \17115 , \17124 );
or \U$17058 ( \17190 , \17187 , \17188 , \17189 );
and \U$17059 ( \17191 , \16978 , \16982 );
and \U$17060 ( \17192 , \16982 , \16987 );
and \U$17061 ( \17193 , \16978 , \16987 );
or \U$17062 ( \17194 , \17191 , \17192 , \17193 );
xor \U$17063 ( \17195 , \17190 , \17194 );
and \U$17064 ( \17196 , \17144 , \17148 );
and \U$17065 ( \17197 , \17148 , \17153 );
and \U$17066 ( \17198 , \17144 , \17153 );
or \U$17067 ( \17199 , \17196 , \17197 , \17198 );
xor \U$17068 ( \17200 , \17195 , \17199 );
and \U$17069 ( \17201 , \17080 , \17094 );
and \U$17070 ( \17202 , \17094 , \17109 );
and \U$17071 ( \17203 , \17080 , \17109 );
or \U$17072 ( \17204 , \17201 , \17202 , \17203 );
and \U$17073 ( \17205 , \17125 , \17139 );
and \U$17074 ( \17206 , \17139 , \17154 );
and \U$17075 ( \17207 , \17125 , \17154 );
or \U$17076 ( \17208 , \17205 , \17206 , \17207 );
xor \U$17077 ( \17209 , \17204 , \17208 );
and \U$17078 ( \17210 , \10584 , \1824 );
not \U$17079 ( \17211 , \17210 );
xnor \U$17080 ( \17212 , \17211 , \1697 );
and \U$17081 ( \17213 , \9897 , \2121 );
and \U$17082 ( \17214 , \10206 , \2008 );
nor \U$17083 ( \17215 , \17213 , \17214 );
xnor \U$17084 ( \17216 , \17215 , \1961 );
xor \U$17085 ( \17217 , \17212 , \17216 );
and \U$17086 ( \17218 , \9169 , \2400 );
and \U$17087 ( \17219 , \9465 , \2246 );
nor \U$17088 ( \17220 , \17218 , \17219 );
xnor \U$17089 ( \17221 , \17220 , \2195 );
xor \U$17090 ( \17222 , \17217 , \17221 );
and \U$17091 ( \17223 , \8652 , \2669 );
and \U$17092 ( \17224 , \8835 , \2538 );
nor \U$17093 ( \17225 , \17223 , \17224 );
xnor \U$17094 ( \17226 , \17225 , \2534 );
and \U$17095 ( \17227 , \8057 , \3103 );
and \U$17096 ( \17228 , \8349 , \2934 );
nor \U$17097 ( \17229 , \17227 , \17228 );
xnor \U$17098 ( \17230 , \17229 , \2839 );
xor \U$17099 ( \17231 , \17226 , \17230 );
and \U$17100 ( \17232 , \7556 , \3357 );
and \U$17101 ( \17233 , \7700 , \3255 );
nor \U$17102 ( \17234 , \17232 , \17233 );
xnor \U$17103 ( \17235 , \17234 , \3156 );
xor \U$17104 ( \17236 , \17231 , \17235 );
xor \U$17105 ( \17237 , \17222 , \17236 );
and \U$17106 ( \17238 , \6945 , \3813 );
and \U$17107 ( \17239 , \7231 , \3557 );
nor \U$17108 ( \17240 , \17238 , \17239 );
xnor \U$17109 ( \17241 , \17240 , \3562 );
and \U$17110 ( \17242 , \6514 , \4132 );
and \U$17111 ( \17243 , \6790 , \4012 );
nor \U$17112 ( \17244 , \17242 , \17243 );
xnor \U$17113 ( \17245 , \17244 , \3925 );
xor \U$17114 ( \17246 , \17241 , \17245 );
and \U$17115 ( \17247 , \6030 , \4581 );
and \U$17116 ( \17248 , \6281 , \4424 );
nor \U$17117 ( \17249 , \17247 , \17248 );
xnor \U$17118 ( \17250 , \17249 , \4377 );
xor \U$17119 ( \17251 , \17246 , \17250 );
xor \U$17120 ( \17252 , \17237 , \17251 );
xor \U$17121 ( \17253 , \17209 , \17252 );
xor \U$17122 ( \17254 , \17200 , \17253 );
and \U$17123 ( \17255 , \17070 , \17074 );
and \U$17124 ( \17256 , \17074 , \17079 );
and \U$17125 ( \17257 , \17070 , \17079 );
or \U$17126 ( \17258 , \17255 , \17256 , \17257 );
and \U$17127 ( \17259 , \17129 , \17133 );
and \U$17128 ( \17260 , \17133 , \17138 );
and \U$17129 ( \17261 , \17129 , \17138 );
or \U$17130 ( \17262 , \17259 , \17260 , \17261 );
xor \U$17131 ( \17263 , \17258 , \17262 );
and \U$17132 ( \17264 , \17084 , \17088 );
and \U$17133 ( \17265 , \17088 , \17093 );
and \U$17134 ( \17266 , \17084 , \17093 );
or \U$17135 ( \17267 , \17264 , \17265 , \17266 );
xor \U$17136 ( \17268 , \17263 , \17267 );
and \U$17137 ( \17269 , \3037 , \8019 );
and \U$17138 ( \17270 , \3143 , \7830 );
nor \U$17139 ( \17271 , \17269 , \17270 );
xnor \U$17140 ( \17272 , \17271 , \7713 );
and \U$17141 ( \17273 , \2757 , \8540 );
and \U$17142 ( \17274 , \2826 , \8292 );
nor \U$17143 ( \17275 , \17273 , \17274 );
xnor \U$17144 ( \17276 , \17275 , \8297 );
xor \U$17145 ( \17277 , \17272 , \17276 );
and \U$17146 ( \17278 , \2366 , \9333 );
and \U$17147 ( \17279 , \2521 , \9006 );
nor \U$17148 ( \17280 , \17278 , \17279 );
xnor \U$17149 ( \17281 , \17280 , \8848 );
xor \U$17150 ( \17282 , \17277 , \17281 );
and \U$17151 ( \17283 , \5469 , \5011 );
and \U$17152 ( \17284 , \5674 , \4878 );
nor \U$17153 ( \17285 , \17283 , \17284 );
xnor \U$17154 ( \17286 , \17285 , \4762 );
and \U$17155 ( \17287 , \4922 , \5485 );
and \U$17156 ( \17288 , \5156 , \5275 );
nor \U$17157 ( \17289 , \17287 , \17288 );
xnor \U$17158 ( \17290 , \17289 , \5169 );
xor \U$17159 ( \17291 , \17286 , \17290 );
and \U$17160 ( \17292 , \4654 , \5996 );
and \U$17161 ( \17293 , \4749 , \5695 );
nor \U$17162 ( \17294 , \17292 , \17293 );
xnor \U$17163 ( \17295 , \17294 , \5687 );
xor \U$17164 ( \17296 , \17291 , \17295 );
xor \U$17165 ( \17297 , \17282 , \17296 );
and \U$17166 ( \17298 , \4160 , \6401 );
and \U$17167 ( \17299 , \4364 , \6143 );
nor \U$17168 ( \17300 , \17298 , \17299 );
xnor \U$17169 ( \17301 , \17300 , \6148 );
and \U$17170 ( \17302 , \3736 , \7055 );
and \U$17171 ( \17303 , \3912 , \6675 );
nor \U$17172 ( \17304 , \17302 , \17303 );
xnor \U$17173 ( \17305 , \17304 , \6680 );
xor \U$17174 ( \17306 , \17301 , \17305 );
and \U$17175 ( \17307 , \3395 , \7489 );
and \U$17176 ( \17308 , \3646 , \7137 );
nor \U$17177 ( \17309 , \17307 , \17308 );
xnor \U$17178 ( \17310 , \17309 , \7142 );
xor \U$17179 ( \17311 , \17306 , \17310 );
xor \U$17180 ( \17312 , \17297 , \17311 );
xor \U$17181 ( \17313 , \17268 , \17312 );
and \U$17182 ( \17314 , \17099 , \17103 );
and \U$17183 ( \17315 , \17103 , \17108 );
and \U$17184 ( \17316 , \17099 , \17108 );
or \U$17185 ( \17317 , \17314 , \17315 , \17316 );
and \U$17186 ( \17318 , \2090 , \9765 );
and \U$17187 ( \17319 , \2182 , \9644 );
nor \U$17188 ( \17320 , \17318 , \17319 );
xnor \U$17189 ( \17321 , \17320 , \9478 );
and \U$17190 ( \17322 , \1802 , \10408 );
and \U$17191 ( \17323 , \1948 , \10116 );
nor \U$17192 ( \17324 , \17322 , \17323 );
xnor \U$17193 ( \17325 , \17324 , \10121 );
xor \U$17194 ( \17326 , \17321 , \17325 );
and \U$17195 ( \17327 , \1684 , \10118 );
xor \U$17196 ( \17328 , \17326 , \17327 );
xnor \U$17197 ( \17329 , \17317 , \17328 );
xor \U$17198 ( \17330 , \17313 , \17329 );
xor \U$17199 ( \17331 , \17254 , \17330 );
xor \U$17200 ( \17332 , \17186 , \17331 );
xor \U$17201 ( \17333 , \17177 , \17332 );
and \U$17202 ( \17334 , \17004 , \17008 );
and \U$17203 ( \17335 , \17008 , \17013 );
and \U$17204 ( \17336 , \17004 , \17013 );
or \U$17205 ( \17337 , \17334 , \17335 , \17336 );
and \U$17206 ( \17338 , \16972 , \16976 );
and \U$17207 ( \17339 , \16976 , \16988 );
and \U$17208 ( \17340 , \16972 , \16988 );
or \U$17209 ( \17341 , \17338 , \17339 , \17340 );
xor \U$17210 ( \17342 , \17337 , \17341 );
and \U$17211 ( \17343 , \17066 , \17110 );
and \U$17212 ( \17344 , \17110 , \17155 );
and \U$17213 ( \17345 , \17066 , \17155 );
or \U$17214 ( \17346 , \17343 , \17344 , \17345 );
xor \U$17215 ( \17347 , \17342 , \17346 );
and \U$17216 ( \17348 , \17018 , \17022 );
and \U$17217 ( \17349 , \17022 , \17027 );
and \U$17218 ( \17350 , \17018 , \17027 );
or \U$17219 ( \17351 , \17348 , \17349 , \17350 );
and \U$17220 ( \17352 , \17043 , \17057 );
and \U$17221 ( \17353 , \17057 , \17156 );
and \U$17222 ( \17354 , \17043 , \17156 );
or \U$17223 ( \17355 , \17352 , \17353 , \17354 );
xor \U$17224 ( \17356 , \17351 , \17355 );
and \U$17225 ( \17357 , \17062 , \17063 );
and \U$17226 ( \17358 , \17063 , \17065 );
and \U$17227 ( \17359 , \17062 , \17065 );
or \U$17228 ( \17360 , \17357 , \17358 , \17359 );
and \U$17229 ( \17361 , \17033 , \17037 );
and \U$17230 ( \17362 , \17037 , \17042 );
and \U$17231 ( \17363 , \17033 , \17042 );
or \U$17232 ( \17364 , \17361 , \17362 , \17363 );
xor \U$17233 ( \17365 , \17360 , \17364 );
and \U$17234 ( \17366 , \17047 , \17051 );
and \U$17235 ( \17367 , \17051 , \17056 );
and \U$17236 ( \17368 , \17047 , \17056 );
or \U$17237 ( \17369 , \17366 , \17367 , \17368 );
xor \U$17238 ( \17370 , \17365 , \17369 );
xor \U$17239 ( \17371 , \17356 , \17370 );
xor \U$17240 ( \17372 , \17347 , \17371 );
xor \U$17241 ( \17373 , \17333 , \17372 );
xor \U$17242 ( \17374 , \17173 , \17373 );
and \U$17243 ( \17375 , \16955 , \17160 );
xor \U$17244 ( \17376 , \17374 , \17375 );
and \U$17245 ( \17377 , \17161 , \17162 );
and \U$17246 ( \17378 , \17163 , \17166 );
or \U$17247 ( \17379 , \17377 , \17378 );
xor \U$17248 ( \17380 , \17376 , \17379 );
buf \U$17249 ( \17381 , \17380 );
buf \U$17250 ( \17382 , \17381 );
and \U$17251 ( \17383 , \17177 , \17332 );
and \U$17252 ( \17384 , \17332 , \17372 );
and \U$17253 ( \17385 , \17177 , \17372 );
or \U$17254 ( \17386 , \17383 , \17384 , \17385 );
and \U$17255 ( \17387 , \17181 , \17185 );
and \U$17256 ( \17388 , \17185 , \17331 );
and \U$17257 ( \17389 , \17181 , \17331 );
or \U$17258 ( \17390 , \17387 , \17388 , \17389 );
and \U$17259 ( \17391 , \17347 , \17371 );
xor \U$17260 ( \17392 , \17390 , \17391 );
and \U$17261 ( \17393 , \17351 , \17355 );
and \U$17262 ( \17394 , \17355 , \17370 );
and \U$17263 ( \17395 , \17351 , \17370 );
or \U$17264 ( \17396 , \17393 , \17394 , \17395 );
and \U$17265 ( \17397 , \17337 , \17341 );
and \U$17266 ( \17398 , \17341 , \17346 );
and \U$17267 ( \17399 , \17337 , \17346 );
or \U$17268 ( \17400 , \17397 , \17398 , \17399 );
and \U$17269 ( \17401 , \17200 , \17253 );
and \U$17270 ( \17402 , \17253 , \17330 );
and \U$17271 ( \17403 , \17200 , \17330 );
or \U$17272 ( \17404 , \17401 , \17402 , \17403 );
xor \U$17273 ( \17405 , \17400 , \17404 );
and \U$17274 ( \17406 , \17282 , \17296 );
and \U$17275 ( \17407 , \17296 , \17311 );
and \U$17276 ( \17408 , \17282 , \17311 );
or \U$17277 ( \17409 , \17406 , \17407 , \17408 );
and \U$17278 ( \17410 , \17222 , \17236 );
and \U$17279 ( \17411 , \17236 , \17251 );
and \U$17280 ( \17412 , \17222 , \17251 );
or \U$17281 ( \17413 , \17410 , \17411 , \17412 );
xor \U$17282 ( \17414 , \17409 , \17413 );
and \U$17283 ( \17415 , \8835 , \2669 );
and \U$17284 ( \17416 , \9169 , \2538 );
nor \U$17285 ( \17417 , \17415 , \17416 );
xnor \U$17286 ( \17418 , \17417 , \2534 );
and \U$17287 ( \17419 , \8349 , \3103 );
and \U$17288 ( \17420 , \8652 , \2934 );
nor \U$17289 ( \17421 , \17419 , \17420 );
xnor \U$17290 ( \17422 , \17421 , \2839 );
xor \U$17291 ( \17423 , \17418 , \17422 );
and \U$17292 ( \17424 , \7700 , \3357 );
and \U$17293 ( \17425 , \8057 , \3255 );
nor \U$17294 ( \17426 , \17424 , \17425 );
xnor \U$17295 ( \17427 , \17426 , \3156 );
xor \U$17296 ( \17428 , \17423 , \17427 );
xor \U$17297 ( \17429 , \17414 , \17428 );
xor \U$17298 ( \17430 , \17405 , \17429 );
xor \U$17299 ( \17431 , \17396 , \17430 );
and \U$17300 ( \17432 , \17190 , \17194 );
and \U$17301 ( \17433 , \17194 , \17199 );
and \U$17302 ( \17434 , \17190 , \17199 );
or \U$17303 ( \17435 , \17432 , \17433 , \17434 );
and \U$17304 ( \17436 , \17258 , \17262 );
and \U$17305 ( \17437 , \17262 , \17267 );
and \U$17306 ( \17438 , \17258 , \17267 );
or \U$17307 ( \17439 , \17436 , \17437 , \17438 );
xor \U$17308 ( \17440 , \17435 , \17439 );
or \U$17309 ( \17441 , \17317 , \17328 );
xor \U$17310 ( \17442 , \17440 , \17441 );
and \U$17311 ( \17443 , \17360 , \17364 );
and \U$17312 ( \17444 , \17364 , \17369 );
and \U$17313 ( \17445 , \17360 , \17369 );
or \U$17314 ( \17446 , \17443 , \17444 , \17445 );
and \U$17315 ( \17447 , \17204 , \17208 );
and \U$17316 ( \17448 , \17208 , \17252 );
and \U$17317 ( \17449 , \17204 , \17252 );
or \U$17318 ( \17450 , \17447 , \17448 , \17449 );
xor \U$17319 ( \17451 , \17446 , \17450 );
and \U$17320 ( \17452 , \17268 , \17312 );
and \U$17321 ( \17453 , \17312 , \17329 );
and \U$17322 ( \17454 , \17268 , \17329 );
or \U$17323 ( \17455 , \17452 , \17453 , \17454 );
xor \U$17324 ( \17456 , \17451 , \17455 );
xor \U$17325 ( \17457 , \17442 , \17456 );
and \U$17326 ( \17458 , \17212 , \17216 );
and \U$17327 ( \17459 , \17216 , \17221 );
and \U$17328 ( \17460 , \17212 , \17221 );
or \U$17329 ( \17461 , \17458 , \17459 , \17460 );
and \U$17330 ( \17462 , \17226 , \17230 );
and \U$17331 ( \17463 , \17230 , \17235 );
and \U$17332 ( \17464 , \17226 , \17235 );
or \U$17333 ( \17465 , \17462 , \17463 , \17464 );
xor \U$17334 ( \17466 , \17461 , \17465 );
and \U$17335 ( \17467 , \17241 , \17245 );
and \U$17336 ( \17468 , \17245 , \17250 );
and \U$17337 ( \17469 , \17241 , \17250 );
or \U$17338 ( \17470 , \17467 , \17468 , \17469 );
xor \U$17339 ( \17471 , \17466 , \17470 );
and \U$17340 ( \17472 , \17272 , \17276 );
and \U$17341 ( \17473 , \17276 , \17281 );
and \U$17342 ( \17474 , \17272 , \17281 );
or \U$17343 ( \17475 , \17472 , \17473 , \17474 );
and \U$17344 ( \17476 , \17286 , \17290 );
and \U$17345 ( \17477 , \17290 , \17295 );
and \U$17346 ( \17478 , \17286 , \17295 );
or \U$17347 ( \17479 , \17476 , \17477 , \17478 );
xor \U$17348 ( \17480 , \17475 , \17479 );
and \U$17349 ( \17481 , \17301 , \17305 );
and \U$17350 ( \17482 , \17305 , \17310 );
and \U$17351 ( \17483 , \17301 , \17310 );
or \U$17352 ( \17484 , \17481 , \17482 , \17483 );
xor \U$17353 ( \17485 , \17480 , \17484 );
xor \U$17354 ( \17486 , \17471 , \17485 );
not \U$17355 ( \17487 , \1697 );
and \U$17356 ( \17488 , \10206 , \2121 );
and \U$17357 ( \17489 , \10584 , \2008 );
nor \U$17358 ( \17490 , \17488 , \17489 );
xnor \U$17359 ( \17491 , \17490 , \1961 );
xor \U$17360 ( \17492 , \17487 , \17491 );
and \U$17361 ( \17493 , \9465 , \2400 );
and \U$17362 ( \17494 , \9897 , \2246 );
nor \U$17363 ( \17495 , \17493 , \17494 );
xnor \U$17364 ( \17496 , \17495 , \2195 );
xor \U$17365 ( \17497 , \17492 , \17496 );
and \U$17366 ( \17498 , \4364 , \6401 );
and \U$17367 ( \17499 , \4654 , \6143 );
nor \U$17368 ( \17500 , \17498 , \17499 );
xnor \U$17369 ( \17501 , \17500 , \6148 );
and \U$17370 ( \17502 , \3912 , \7055 );
and \U$17371 ( \17503 , \4160 , \6675 );
nor \U$17372 ( \17504 , \17502 , \17503 );
xnor \U$17373 ( \17505 , \17504 , \6680 );
xor \U$17374 ( \17506 , \17501 , \17505 );
and \U$17375 ( \17507 , \3646 , \7489 );
and \U$17376 ( \17508 , \3736 , \7137 );
nor \U$17377 ( \17509 , \17507 , \17508 );
xnor \U$17378 ( \17510 , \17509 , \7142 );
xor \U$17379 ( \17511 , \17506 , \17510 );
and \U$17380 ( \17512 , \5674 , \5011 );
and \U$17381 ( \17513 , \6030 , \4878 );
nor \U$17382 ( \17514 , \17512 , \17513 );
xnor \U$17383 ( \17515 , \17514 , \4762 );
and \U$17384 ( \17516 , \5156 , \5485 );
and \U$17385 ( \17517 , \5469 , \5275 );
nor \U$17386 ( \17518 , \17516 , \17517 );
xnor \U$17387 ( \17519 , \17518 , \5169 );
xor \U$17388 ( \17520 , \17515 , \17519 );
and \U$17389 ( \17521 , \4749 , \5996 );
and \U$17390 ( \17522 , \4922 , \5695 );
nor \U$17391 ( \17523 , \17521 , \17522 );
xnor \U$17392 ( \17524 , \17523 , \5687 );
xor \U$17393 ( \17525 , \17520 , \17524 );
xor \U$17394 ( \17526 , \17511 , \17525 );
and \U$17395 ( \17527 , \7231 , \3813 );
and \U$17396 ( \17528 , \7556 , \3557 );
nor \U$17397 ( \17529 , \17527 , \17528 );
xnor \U$17398 ( \17530 , \17529 , \3562 );
and \U$17399 ( \17531 , \6790 , \4132 );
and \U$17400 ( \17532 , \6945 , \4012 );
nor \U$17401 ( \17533 , \17531 , \17532 );
xnor \U$17402 ( \17534 , \17533 , \3925 );
xor \U$17403 ( \17535 , \17530 , \17534 );
and \U$17404 ( \17536 , \6281 , \4581 );
and \U$17405 ( \17537 , \6514 , \4424 );
nor \U$17406 ( \17538 , \17536 , \17537 );
xnor \U$17407 ( \17539 , \17538 , \4377 );
xor \U$17408 ( \17540 , \17535 , \17539 );
xor \U$17409 ( \17541 , \17526 , \17540 );
xor \U$17410 ( \17542 , \17497 , \17541 );
and \U$17411 ( \17543 , \17321 , \17325 );
and \U$17412 ( \17544 , \17325 , \17327 );
and \U$17413 ( \17545 , \17321 , \17327 );
or \U$17414 ( \17546 , \17543 , \17544 , \17545 );
and \U$17415 ( \17547 , \2182 , \9765 );
and \U$17416 ( \17548 , \2366 , \9644 );
nor \U$17417 ( \17549 , \17547 , \17548 );
xnor \U$17418 ( \17550 , \17549 , \9478 );
and \U$17419 ( \17551 , \1948 , \10408 );
and \U$17420 ( \17552 , \2090 , \10116 );
nor \U$17421 ( \17553 , \17551 , \17552 );
xnor \U$17422 ( \17554 , \17553 , \10121 );
xor \U$17423 ( \17555 , \17550 , \17554 );
and \U$17424 ( \17556 , \1802 , \10118 );
xor \U$17425 ( \17557 , \17555 , \17556 );
xor \U$17426 ( \17558 , \17546 , \17557 );
and \U$17427 ( \17559 , \3143 , \8019 );
and \U$17428 ( \17560 , \3395 , \7830 );
nor \U$17429 ( \17561 , \17559 , \17560 );
xnor \U$17430 ( \17562 , \17561 , \7713 );
and \U$17431 ( \17563 , \2826 , \8540 );
and \U$17432 ( \17564 , \3037 , \8292 );
nor \U$17433 ( \17565 , \17563 , \17564 );
xnor \U$17434 ( \17566 , \17565 , \8297 );
xor \U$17435 ( \17567 , \17562 , \17566 );
and \U$17436 ( \17568 , \2521 , \9333 );
and \U$17437 ( \17569 , \2757 , \9006 );
nor \U$17438 ( \17570 , \17568 , \17569 );
xnor \U$17439 ( \17571 , \17570 , \8848 );
xor \U$17440 ( \17572 , \17567 , \17571 );
xor \U$17441 ( \17573 , \17558 , \17572 );
xor \U$17442 ( \17574 , \17542 , \17573 );
xor \U$17443 ( \17575 , \17486 , \17574 );
xor \U$17444 ( \17576 , \17457 , \17575 );
xor \U$17445 ( \17577 , \17431 , \17576 );
xor \U$17446 ( \17578 , \17392 , \17577 );
xor \U$17447 ( \17579 , \17386 , \17578 );
and \U$17448 ( \17580 , \17173 , \17373 );
xor \U$17449 ( \17581 , \17579 , \17580 );
and \U$17450 ( \17582 , \17374 , \17375 );
and \U$17451 ( \17583 , \17376 , \17379 );
or \U$17452 ( \17584 , \17582 , \17583 );
xor \U$17453 ( \17585 , \17581 , \17584 );
buf \U$17454 ( \17586 , \17585 );
buf \U$17455 ( \17587 , \17586 );
and \U$17456 ( \17588 , \17390 , \17391 );
and \U$17457 ( \17589 , \17391 , \17577 );
and \U$17458 ( \17590 , \17390 , \17577 );
or \U$17459 ( \17591 , \17588 , \17589 , \17590 );
and \U$17460 ( \17592 , \17396 , \17430 );
and \U$17461 ( \17593 , \17430 , \17576 );
and \U$17462 ( \17594 , \17396 , \17576 );
or \U$17463 ( \17595 , \17592 , \17593 , \17594 );
and \U$17464 ( \17596 , \17400 , \17404 );
and \U$17465 ( \17597 , \17404 , \17429 );
and \U$17466 ( \17598 , \17400 , \17429 );
or \U$17467 ( \17599 , \17596 , \17597 , \17598 );
and \U$17468 ( \17600 , \17442 , \17456 );
and \U$17469 ( \17601 , \17456 , \17575 );
and \U$17470 ( \17602 , \17442 , \17575 );
or \U$17471 ( \17603 , \17600 , \17601 , \17602 );
xor \U$17472 ( \17604 , \17599 , \17603 );
and \U$17473 ( \17605 , \17435 , \17439 );
and \U$17474 ( \17606 , \17439 , \17441 );
and \U$17475 ( \17607 , \17435 , \17441 );
or \U$17476 ( \17608 , \17605 , \17606 , \17607 );
and \U$17477 ( \17609 , \17409 , \17413 );
and \U$17478 ( \17610 , \17413 , \17428 );
and \U$17479 ( \17611 , \17409 , \17428 );
or \U$17480 ( \17612 , \17609 , \17610 , \17611 );
xor \U$17481 ( \17613 , \17608 , \17612 );
and \U$17482 ( \17614 , \17497 , \17541 );
and \U$17483 ( \17615 , \17541 , \17573 );
and \U$17484 ( \17616 , \17497 , \17573 );
or \U$17485 ( \17617 , \17614 , \17615 , \17616 );
xor \U$17486 ( \17618 , \17613 , \17617 );
xor \U$17487 ( \17619 , \17604 , \17618 );
xor \U$17488 ( \17620 , \17595 , \17619 );
and \U$17489 ( \17621 , \17446 , \17450 );
and \U$17490 ( \17622 , \17450 , \17455 );
and \U$17491 ( \17623 , \17446 , \17455 );
or \U$17492 ( \17624 , \17621 , \17622 , \17623 );
and \U$17493 ( \17625 , \17471 , \17485 );
and \U$17494 ( \17626 , \17485 , \17574 );
and \U$17495 ( \17627 , \17471 , \17574 );
or \U$17496 ( \17628 , \17625 , \17626 , \17627 );
xor \U$17497 ( \17629 , \17624 , \17628 );
and \U$17498 ( \17630 , \17461 , \17465 );
and \U$17499 ( \17631 , \17465 , \17470 );
and \U$17500 ( \17632 , \17461 , \17470 );
or \U$17501 ( \17633 , \17630 , \17631 , \17632 );
and \U$17502 ( \17634 , \17475 , \17479 );
and \U$17503 ( \17635 , \17479 , \17484 );
and \U$17504 ( \17636 , \17475 , \17484 );
or \U$17505 ( \17637 , \17634 , \17635 , \17636 );
xor \U$17506 ( \17638 , \17633 , \17637 );
and \U$17507 ( \17639 , \17546 , \17557 );
and \U$17508 ( \17640 , \17557 , \17572 );
and \U$17509 ( \17641 , \17546 , \17572 );
or \U$17510 ( \17642 , \17639 , \17640 , \17641 );
xor \U$17511 ( \17643 , \17638 , \17642 );
and \U$17512 ( \17644 , \17501 , \17505 );
and \U$17513 ( \17645 , \17505 , \17510 );
and \U$17514 ( \17646 , \17501 , \17510 );
or \U$17515 ( \17647 , \17644 , \17645 , \17646 );
and \U$17516 ( \17648 , \17515 , \17519 );
and \U$17517 ( \17649 , \17519 , \17524 );
and \U$17518 ( \17650 , \17515 , \17524 );
or \U$17519 ( \17651 , \17648 , \17649 , \17650 );
xor \U$17520 ( \17652 , \17647 , \17651 );
and \U$17521 ( \17653 , \17562 , \17566 );
and \U$17522 ( \17654 , \17566 , \17571 );
and \U$17523 ( \17655 , \17562 , \17571 );
or \U$17524 ( \17656 , \17653 , \17654 , \17655 );
xor \U$17525 ( \17657 , \17652 , \17656 );
and \U$17526 ( \17658 , \17487 , \17491 );
and \U$17527 ( \17659 , \17491 , \17496 );
and \U$17528 ( \17660 , \17487 , \17496 );
or \U$17529 ( \17661 , \17658 , \17659 , \17660 );
and \U$17530 ( \17662 , \17418 , \17422 );
and \U$17531 ( \17663 , \17422 , \17427 );
and \U$17532 ( \17664 , \17418 , \17427 );
or \U$17533 ( \17665 , \17662 , \17663 , \17664 );
xor \U$17534 ( \17666 , \17661 , \17665 );
and \U$17535 ( \17667 , \17530 , \17534 );
and \U$17536 ( \17668 , \17534 , \17539 );
and \U$17537 ( \17669 , \17530 , \17539 );
or \U$17538 ( \17670 , \17667 , \17668 , \17669 );
xor \U$17539 ( \17671 , \17666 , \17670 );
xor \U$17540 ( \17672 , \17657 , \17671 );
and \U$17541 ( \17673 , \17550 , \17554 );
and \U$17542 ( \17674 , \17554 , \17556 );
and \U$17543 ( \17675 , \17550 , \17556 );
or \U$17544 ( \17676 , \17673 , \17674 , \17675 );
and \U$17545 ( \17677 , \3037 , \8540 );
and \U$17546 ( \17678 , \3143 , \8292 );
nor \U$17547 ( \17679 , \17677 , \17678 );
xnor \U$17548 ( \17680 , \17679 , \8297 );
and \U$17549 ( \17681 , \2757 , \9333 );
and \U$17550 ( \17682 , \2826 , \9006 );
nor \U$17551 ( \17683 , \17681 , \17682 );
xnor \U$17552 ( \17684 , \17683 , \8848 );
xor \U$17553 ( \17685 , \17680 , \17684 );
and \U$17554 ( \17686 , \2366 , \9765 );
and \U$17555 ( \17687 , \2521 , \9644 );
nor \U$17556 ( \17688 , \17686 , \17687 );
xnor \U$17557 ( \17689 , \17688 , \9478 );
xor \U$17558 ( \17690 , \17685 , \17689 );
xor \U$17559 ( \17691 , \17676 , \17690 );
and \U$17560 ( \17692 , \2090 , \10408 );
and \U$17561 ( \17693 , \2182 , \10116 );
nor \U$17562 ( \17694 , \17692 , \17693 );
xnor \U$17563 ( \17695 , \17694 , \10121 );
and \U$17564 ( \17696 , \1948 , \10118 );
xnor \U$17565 ( \17697 , \17695 , \17696 );
xor \U$17566 ( \17698 , \17691 , \17697 );
xor \U$17567 ( \17699 , \17672 , \17698 );
xor \U$17568 ( \17700 , \17643 , \17699 );
and \U$17569 ( \17701 , \17511 , \17525 );
and \U$17570 ( \17702 , \17525 , \17540 );
and \U$17571 ( \17703 , \17511 , \17540 );
or \U$17572 ( \17704 , \17701 , \17702 , \17703 );
and \U$17573 ( \17705 , \5469 , \5485 );
and \U$17574 ( \17706 , \5674 , \5275 );
nor \U$17575 ( \17707 , \17705 , \17706 );
xnor \U$17576 ( \17708 , \17707 , \5169 );
and \U$17577 ( \17709 , \4922 , \5996 );
and \U$17578 ( \17710 , \5156 , \5695 );
nor \U$17579 ( \17711 , \17709 , \17710 );
xnor \U$17580 ( \17712 , \17711 , \5687 );
xor \U$17581 ( \17713 , \17708 , \17712 );
and \U$17582 ( \17714 , \4654 , \6401 );
and \U$17583 ( \17715 , \4749 , \6143 );
nor \U$17584 ( \17716 , \17714 , \17715 );
xnor \U$17585 ( \17717 , \17716 , \6148 );
xor \U$17586 ( \17718 , \17713 , \17717 );
and \U$17587 ( \17719 , \4160 , \7055 );
and \U$17588 ( \17720 , \4364 , \6675 );
nor \U$17589 ( \17721 , \17719 , \17720 );
xnor \U$17590 ( \17722 , \17721 , \6680 );
and \U$17591 ( \17723 , \3736 , \7489 );
and \U$17592 ( \17724 , \3912 , \7137 );
nor \U$17593 ( \17725 , \17723 , \17724 );
xnor \U$17594 ( \17726 , \17725 , \7142 );
xor \U$17595 ( \17727 , \17722 , \17726 );
and \U$17596 ( \17728 , \3395 , \8019 );
and \U$17597 ( \17729 , \3646 , \7830 );
nor \U$17598 ( \17730 , \17728 , \17729 );
xnor \U$17599 ( \17731 , \17730 , \7713 );
xor \U$17600 ( \17732 , \17727 , \17731 );
xor \U$17601 ( \17733 , \17718 , \17732 );
and \U$17602 ( \17734 , \6945 , \4132 );
and \U$17603 ( \17735 , \7231 , \4012 );
nor \U$17604 ( \17736 , \17734 , \17735 );
xnor \U$17605 ( \17737 , \17736 , \3925 );
and \U$17606 ( \17738 , \6514 , \4581 );
and \U$17607 ( \17739 , \6790 , \4424 );
nor \U$17608 ( \17740 , \17738 , \17739 );
xnor \U$17609 ( \17741 , \17740 , \4377 );
xor \U$17610 ( \17742 , \17737 , \17741 );
and \U$17611 ( \17743 , \6030 , \5011 );
and \U$17612 ( \17744 , \6281 , \4878 );
nor \U$17613 ( \17745 , \17743 , \17744 );
xnor \U$17614 ( \17746 , \17745 , \4762 );
xor \U$17615 ( \17747 , \17742 , \17746 );
xor \U$17616 ( \17748 , \17733 , \17747 );
xor \U$17617 ( \17749 , \17704 , \17748 );
and \U$17618 ( \17750 , \10584 , \2121 );
not \U$17619 ( \17751 , \17750 );
xnor \U$17620 ( \17752 , \17751 , \1961 );
and \U$17621 ( \17753 , \9897 , \2400 );
and \U$17622 ( \17754 , \10206 , \2246 );
nor \U$17623 ( \17755 , \17753 , \17754 );
xnor \U$17624 ( \17756 , \17755 , \2195 );
xor \U$17625 ( \17757 , \17752 , \17756 );
and \U$17626 ( \17758 , \9169 , \2669 );
and \U$17627 ( \17759 , \9465 , \2538 );
nor \U$17628 ( \17760 , \17758 , \17759 );
xnor \U$17629 ( \17761 , \17760 , \2534 );
xor \U$17630 ( \17762 , \17757 , \17761 );
and \U$17631 ( \17763 , \8652 , \3103 );
and \U$17632 ( \17764 , \8835 , \2934 );
nor \U$17633 ( \17765 , \17763 , \17764 );
xnor \U$17634 ( \17766 , \17765 , \2839 );
and \U$17635 ( \17767 , \8057 , \3357 );
and \U$17636 ( \17768 , \8349 , \3255 );
nor \U$17637 ( \17769 , \17767 , \17768 );
xnor \U$17638 ( \17770 , \17769 , \3156 );
xor \U$17639 ( \17771 , \17766 , \17770 );
and \U$17640 ( \17772 , \7556 , \3813 );
and \U$17641 ( \17773 , \7700 , \3557 );
nor \U$17642 ( \17774 , \17772 , \17773 );
xnor \U$17643 ( \17775 , \17774 , \3562 );
xor \U$17644 ( \17776 , \17771 , \17775 );
xor \U$17645 ( \17777 , \17762 , \17776 );
xor \U$17646 ( \17778 , \17749 , \17777 );
xor \U$17647 ( \17779 , \17700 , \17778 );
xor \U$17648 ( \17780 , \17629 , \17779 );
xor \U$17649 ( \17781 , \17620 , \17780 );
xor \U$17650 ( \17782 , \17591 , \17781 );
and \U$17651 ( \17783 , \17386 , \17578 );
xor \U$17652 ( \17784 , \17782 , \17783 );
and \U$17653 ( \17785 , \17579 , \17580 );
and \U$17654 ( \17786 , \17581 , \17584 );
or \U$17655 ( \17787 , \17785 , \17786 );
xor \U$17656 ( \17788 , \17784 , \17787 );
buf \U$17657 ( \17789 , \17788 );
buf \U$17658 ( \17790 , \17789 );
and \U$17659 ( \17791 , \17599 , \17603 );
and \U$17660 ( \17792 , \17603 , \17618 );
and \U$17661 ( \17793 , \17599 , \17618 );
or \U$17662 ( \17794 , \17791 , \17792 , \17793 );
and \U$17663 ( \17795 , \17595 , \17619 );
and \U$17664 ( \17796 , \17619 , \17780 );
and \U$17665 ( \17797 , \17595 , \17780 );
or \U$17666 ( \17798 , \17795 , \17796 , \17797 );
xor \U$17667 ( \17799 , \17794 , \17798 );
and \U$17668 ( \17800 , \17624 , \17628 );
and \U$17669 ( \17801 , \17628 , \17779 );
and \U$17670 ( \17802 , \17624 , \17779 );
or \U$17671 ( \17803 , \17800 , \17801 , \17802 );
and \U$17672 ( \17804 , \17608 , \17612 );
and \U$17673 ( \17805 , \17612 , \17617 );
and \U$17674 ( \17806 , \17608 , \17617 );
or \U$17675 ( \17807 , \17804 , \17805 , \17806 );
and \U$17676 ( \17808 , \17643 , \17699 );
and \U$17677 ( \17809 , \17699 , \17778 );
and \U$17678 ( \17810 , \17643 , \17778 );
or \U$17679 ( \17811 , \17808 , \17809 , \17810 );
xor \U$17680 ( \17812 , \17807 , \17811 );
and \U$17681 ( \17813 , \17647 , \17651 );
and \U$17682 ( \17814 , \17651 , \17656 );
and \U$17683 ( \17815 , \17647 , \17656 );
or \U$17684 ( \17816 , \17813 , \17814 , \17815 );
and \U$17685 ( \17817 , \17661 , \17665 );
and \U$17686 ( \17818 , \17665 , \17670 );
and \U$17687 ( \17819 , \17661 , \17670 );
or \U$17688 ( \17820 , \17817 , \17818 , \17819 );
xor \U$17689 ( \17821 , \17816 , \17820 );
and \U$17690 ( \17822 , \17676 , \17690 );
and \U$17691 ( \17823 , \17690 , \17697 );
and \U$17692 ( \17824 , \17676 , \17697 );
or \U$17693 ( \17825 , \17822 , \17823 , \17824 );
xor \U$17694 ( \17826 , \17821 , \17825 );
xor \U$17695 ( \17827 , \17812 , \17826 );
xor \U$17696 ( \17828 , \17803 , \17827 );
and \U$17697 ( \17829 , \17633 , \17637 );
and \U$17698 ( \17830 , \17637 , \17642 );
and \U$17699 ( \17831 , \17633 , \17642 );
or \U$17700 ( \17832 , \17829 , \17830 , \17831 );
and \U$17701 ( \17833 , \17657 , \17671 );
and \U$17702 ( \17834 , \17671 , \17698 );
and \U$17703 ( \17835 , \17657 , \17698 );
or \U$17704 ( \17836 , \17833 , \17834 , \17835 );
xor \U$17705 ( \17837 , \17832 , \17836 );
and \U$17706 ( \17838 , \17704 , \17748 );
and \U$17707 ( \17839 , \17748 , \17777 );
and \U$17708 ( \17840 , \17704 , \17777 );
or \U$17709 ( \17841 , \17838 , \17839 , \17840 );
xor \U$17710 ( \17842 , \17837 , \17841 );
and \U$17711 ( \17843 , \17752 , \17756 );
and \U$17712 ( \17844 , \17756 , \17761 );
and \U$17713 ( \17845 , \17752 , \17761 );
or \U$17714 ( \17846 , \17843 , \17844 , \17845 );
and \U$17715 ( \17847 , \17766 , \17770 );
and \U$17716 ( \17848 , \17770 , \17775 );
and \U$17717 ( \17849 , \17766 , \17775 );
or \U$17718 ( \17850 , \17847 , \17848 , \17849 );
xor \U$17719 ( \17851 , \17846 , \17850 );
and \U$17720 ( \17852 , \17737 , \17741 );
and \U$17721 ( \17853 , \17741 , \17746 );
and \U$17722 ( \17854 , \17737 , \17746 );
or \U$17723 ( \17855 , \17852 , \17853 , \17854 );
xor \U$17724 ( \17856 , \17851 , \17855 );
and \U$17725 ( \17857 , \17718 , \17732 );
and \U$17726 ( \17858 , \17732 , \17747 );
and \U$17727 ( \17859 , \17718 , \17747 );
or \U$17728 ( \17860 , \17857 , \17858 , \17859 );
and \U$17729 ( \17861 , \17762 , \17776 );
xor \U$17730 ( \17862 , \17860 , \17861 );
not \U$17731 ( \17863 , \1961 );
and \U$17732 ( \17864 , \10206 , \2400 );
and \U$17733 ( \17865 , \10584 , \2246 );
nor \U$17734 ( \17866 , \17864 , \17865 );
xnor \U$17735 ( \17867 , \17866 , \2195 );
xor \U$17736 ( \17868 , \17863 , \17867 );
and \U$17737 ( \17869 , \9465 , \2669 );
and \U$17738 ( \17870 , \9897 , \2538 );
nor \U$17739 ( \17871 , \17869 , \17870 );
xnor \U$17740 ( \17872 , \17871 , \2534 );
xor \U$17741 ( \17873 , \17868 , \17872 );
and \U$17742 ( \17874 , \8835 , \3103 );
and \U$17743 ( \17875 , \9169 , \2934 );
nor \U$17744 ( \17876 , \17874 , \17875 );
xnor \U$17745 ( \17877 , \17876 , \2839 );
and \U$17746 ( \17878 , \8349 , \3357 );
and \U$17747 ( \17879 , \8652 , \3255 );
nor \U$17748 ( \17880 , \17878 , \17879 );
xnor \U$17749 ( \17881 , \17880 , \3156 );
xor \U$17750 ( \17882 , \17877 , \17881 );
and \U$17751 ( \17883 , \7700 , \3813 );
and \U$17752 ( \17884 , \8057 , \3557 );
nor \U$17753 ( \17885 , \17883 , \17884 );
xnor \U$17754 ( \17886 , \17885 , \3562 );
xor \U$17755 ( \17887 , \17882 , \17886 );
xor \U$17756 ( \17888 , \17873 , \17887 );
and \U$17757 ( \17889 , \7231 , \4132 );
and \U$17758 ( \17890 , \7556 , \4012 );
nor \U$17759 ( \17891 , \17889 , \17890 );
xnor \U$17760 ( \17892 , \17891 , \3925 );
and \U$17761 ( \17893 , \6790 , \4581 );
and \U$17762 ( \17894 , \6945 , \4424 );
nor \U$17763 ( \17895 , \17893 , \17894 );
xnor \U$17764 ( \17896 , \17895 , \4377 );
xor \U$17765 ( \17897 , \17892 , \17896 );
and \U$17766 ( \17898 , \6281 , \5011 );
and \U$17767 ( \17899 , \6514 , \4878 );
nor \U$17768 ( \17900 , \17898 , \17899 );
xnor \U$17769 ( \17901 , \17900 , \4762 );
xor \U$17770 ( \17902 , \17897 , \17901 );
xor \U$17771 ( \17903 , \17888 , \17902 );
xor \U$17772 ( \17904 , \17862 , \17903 );
xor \U$17773 ( \17905 , \17856 , \17904 );
and \U$17774 ( \17906 , \17708 , \17712 );
and \U$17775 ( \17907 , \17712 , \17717 );
and \U$17776 ( \17908 , \17708 , \17717 );
or \U$17777 ( \17909 , \17906 , \17907 , \17908 );
and \U$17778 ( \17910 , \17722 , \17726 );
and \U$17779 ( \17911 , \17726 , \17731 );
and \U$17780 ( \17912 , \17722 , \17731 );
or \U$17781 ( \17913 , \17910 , \17911 , \17912 );
xor \U$17782 ( \17914 , \17909 , \17913 );
and \U$17783 ( \17915 , \17680 , \17684 );
and \U$17784 ( \17916 , \17684 , \17689 );
and \U$17785 ( \17917 , \17680 , \17689 );
or \U$17786 ( \17918 , \17915 , \17916 , \17917 );
xor \U$17787 ( \17919 , \17914 , \17918 );
or \U$17788 ( \17920 , \17695 , \17696 );
and \U$17789 ( \17921 , \2182 , \10408 );
and \U$17790 ( \17922 , \2366 , \10116 );
nor \U$17791 ( \17923 , \17921 , \17922 );
xnor \U$17792 ( \17924 , \17923 , \10121 );
xor \U$17793 ( \17925 , \17920 , \17924 );
and \U$17794 ( \17926 , \2090 , \10118 );
xor \U$17795 ( \17927 , \17925 , \17926 );
xor \U$17796 ( \17928 , \17919 , \17927 );
and \U$17797 ( \17929 , \4364 , \7055 );
and \U$17798 ( \17930 , \4654 , \6675 );
nor \U$17799 ( \17931 , \17929 , \17930 );
xnor \U$17800 ( \17932 , \17931 , \6680 );
and \U$17801 ( \17933 , \3912 , \7489 );
and \U$17802 ( \17934 , \4160 , \7137 );
nor \U$17803 ( \17935 , \17933 , \17934 );
xnor \U$17804 ( \17936 , \17935 , \7142 );
xor \U$17805 ( \17937 , \17932 , \17936 );
and \U$17806 ( \17938 , \3646 , \8019 );
and \U$17807 ( \17939 , \3736 , \7830 );
nor \U$17808 ( \17940 , \17938 , \17939 );
xnor \U$17809 ( \17941 , \17940 , \7713 );
xor \U$17810 ( \17942 , \17937 , \17941 );
and \U$17811 ( \17943 , \5674 , \5485 );
and \U$17812 ( \17944 , \6030 , \5275 );
nor \U$17813 ( \17945 , \17943 , \17944 );
xnor \U$17814 ( \17946 , \17945 , \5169 );
and \U$17815 ( \17947 , \5156 , \5996 );
and \U$17816 ( \17948 , \5469 , \5695 );
nor \U$17817 ( \17949 , \17947 , \17948 );
xnor \U$17818 ( \17950 , \17949 , \5687 );
xor \U$17819 ( \17951 , \17946 , \17950 );
and \U$17820 ( \17952 , \4749 , \6401 );
and \U$17821 ( \17953 , \4922 , \6143 );
nor \U$17822 ( \17954 , \17952 , \17953 );
xnor \U$17823 ( \17955 , \17954 , \6148 );
xor \U$17824 ( \17956 , \17951 , \17955 );
xor \U$17825 ( \17957 , \17942 , \17956 );
and \U$17826 ( \17958 , \3143 , \8540 );
and \U$17827 ( \17959 , \3395 , \8292 );
nor \U$17828 ( \17960 , \17958 , \17959 );
xnor \U$17829 ( \17961 , \17960 , \8297 );
and \U$17830 ( \17962 , \2826 , \9333 );
and \U$17831 ( \17963 , \3037 , \9006 );
nor \U$17832 ( \17964 , \17962 , \17963 );
xnor \U$17833 ( \17965 , \17964 , \8848 );
xor \U$17834 ( \17966 , \17961 , \17965 );
and \U$17835 ( \17967 , \2521 , \9765 );
and \U$17836 ( \17968 , \2757 , \9644 );
nor \U$17837 ( \17969 , \17967 , \17968 );
xnor \U$17838 ( \17970 , \17969 , \9478 );
xor \U$17839 ( \17971 , \17966 , \17970 );
xor \U$17840 ( \17972 , \17957 , \17971 );
xor \U$17841 ( \17973 , \17928 , \17972 );
xor \U$17842 ( \17974 , \17905 , \17973 );
xor \U$17843 ( \17975 , \17842 , \17974 );
xor \U$17844 ( \17976 , \17828 , \17975 );
xor \U$17845 ( \17977 , \17799 , \17976 );
and \U$17846 ( \17978 , \17591 , \17781 );
xor \U$17847 ( \17979 , \17977 , \17978 );
and \U$17848 ( \17980 , \17782 , \17783 );
and \U$17849 ( \17981 , \17784 , \17787 );
or \U$17850 ( \17982 , \17980 , \17981 );
xor \U$17851 ( \17983 , \17979 , \17982 );
buf \U$17852 ( \17984 , \17983 );
buf \U$17853 ( \17985 , \17984 );
and \U$17854 ( \17986 , \17803 , \17827 );
and \U$17855 ( \17987 , \17827 , \17975 );
and \U$17856 ( \17988 , \17803 , \17975 );
or \U$17857 ( \17989 , \17986 , \17987 , \17988 );
and \U$17858 ( \17990 , \17832 , \17836 );
and \U$17859 ( \17991 , \17836 , \17841 );
and \U$17860 ( \17992 , \17832 , \17841 );
or \U$17861 ( \17993 , \17990 , \17991 , \17992 );
and \U$17862 ( \17994 , \17856 , \17904 );
and \U$17863 ( \17995 , \17904 , \17973 );
and \U$17864 ( \17996 , \17856 , \17973 );
or \U$17865 ( \17997 , \17994 , \17995 , \17996 );
xor \U$17866 ( \17998 , \17993 , \17997 );
and \U$17867 ( \17999 , \17942 , \17956 );
and \U$17868 ( \18000 , \17956 , \17971 );
and \U$17869 ( \18001 , \17942 , \17971 );
or \U$17870 ( \18002 , \17999 , \18000 , \18001 );
and \U$17871 ( \18003 , \17873 , \17887 );
and \U$17872 ( \18004 , \17887 , \17902 );
and \U$17873 ( \18005 , \17873 , \17902 );
or \U$17874 ( \18006 , \18003 , \18004 , \18005 );
xor \U$17875 ( \18007 , \18002 , \18006 );
and \U$17876 ( \18008 , \8652 , \3357 );
and \U$17877 ( \18009 , \8835 , \3255 );
nor \U$17878 ( \18010 , \18008 , \18009 );
xnor \U$17879 ( \18011 , \18010 , \3156 );
and \U$17880 ( \18012 , \8057 , \3813 );
and \U$17881 ( \18013 , \8349 , \3557 );
nor \U$17882 ( \18014 , \18012 , \18013 );
xnor \U$17883 ( \18015 , \18014 , \3562 );
xor \U$17884 ( \18016 , \18011 , \18015 );
and \U$17885 ( \18017 , \7556 , \4132 );
and \U$17886 ( \18018 , \7700 , \4012 );
nor \U$17887 ( \18019 , \18017 , \18018 );
xnor \U$17888 ( \18020 , \18019 , \3925 );
xor \U$17889 ( \18021 , \18016 , \18020 );
xor \U$17890 ( \18022 , \18007 , \18021 );
xor \U$17891 ( \18023 , \17998 , \18022 );
xor \U$17892 ( \18024 , \17989 , \18023 );
and \U$17893 ( \18025 , \17807 , \17811 );
and \U$17894 ( \18026 , \17811 , \17826 );
and \U$17895 ( \18027 , \17807 , \17826 );
or \U$17896 ( \18028 , \18025 , \18026 , \18027 );
and \U$17897 ( \18029 , \17842 , \17974 );
xor \U$17898 ( \18030 , \18028 , \18029 );
and \U$17899 ( \18031 , \17909 , \17913 );
and \U$17900 ( \18032 , \17913 , \17918 );
and \U$17901 ( \18033 , \17909 , \17918 );
or \U$17902 ( \18034 , \18031 , \18032 , \18033 );
and \U$17903 ( \18035 , \17920 , \17924 );
and \U$17904 ( \18036 , \17924 , \17926 );
and \U$17905 ( \18037 , \17920 , \17926 );
or \U$17906 ( \18038 , \18035 , \18036 , \18037 );
xor \U$17907 ( \18039 , \18034 , \18038 );
and \U$17908 ( \18040 , \17846 , \17850 );
and \U$17909 ( \18041 , \17850 , \17855 );
and \U$17910 ( \18042 , \17846 , \17855 );
or \U$17911 ( \18043 , \18040 , \18041 , \18042 );
xor \U$17912 ( \18044 , \18039 , \18043 );
and \U$17913 ( \18045 , \17816 , \17820 );
and \U$17914 ( \18046 , \17820 , \17825 );
and \U$17915 ( \18047 , \17816 , \17825 );
or \U$17916 ( \18048 , \18045 , \18046 , \18047 );
and \U$17917 ( \18049 , \17860 , \17861 );
and \U$17918 ( \18050 , \17861 , \17903 );
and \U$17919 ( \18051 , \17860 , \17903 );
or \U$17920 ( \18052 , \18049 , \18050 , \18051 );
xor \U$17921 ( \18053 , \18048 , \18052 );
and \U$17922 ( \18054 , \17919 , \17927 );
and \U$17923 ( \18055 , \17927 , \17972 );
and \U$17924 ( \18056 , \17919 , \17972 );
or \U$17925 ( \18057 , \18054 , \18055 , \18056 );
xor \U$17926 ( \18058 , \18053 , \18057 );
xor \U$17927 ( \18059 , \18044 , \18058 );
and \U$17928 ( \18060 , \17863 , \17867 );
and \U$17929 ( \18061 , \17867 , \17872 );
and \U$17930 ( \18062 , \17863 , \17872 );
or \U$17931 ( \18063 , \18060 , \18061 , \18062 );
and \U$17932 ( \18064 , \17877 , \17881 );
and \U$17933 ( \18065 , \17881 , \17886 );
and \U$17934 ( \18066 , \17877 , \17886 );
or \U$17935 ( \18067 , \18064 , \18065 , \18066 );
xor \U$17936 ( \18068 , \18063 , \18067 );
and \U$17937 ( \18069 , \17892 , \17896 );
and \U$17938 ( \18070 , \17896 , \17901 );
and \U$17939 ( \18071 , \17892 , \17901 );
or \U$17940 ( \18072 , \18069 , \18070 , \18071 );
xor \U$17941 ( \18073 , \18068 , \18072 );
and \U$17942 ( \18074 , \17932 , \17936 );
and \U$17943 ( \18075 , \17936 , \17941 );
and \U$17944 ( \18076 , \17932 , \17941 );
or \U$17945 ( \18077 , \18074 , \18075 , \18076 );
and \U$17946 ( \18078 , \17946 , \17950 );
and \U$17947 ( \18079 , \17950 , \17955 );
and \U$17948 ( \18080 , \17946 , \17955 );
or \U$17949 ( \18081 , \18078 , \18079 , \18080 );
xor \U$17950 ( \18082 , \18077 , \18081 );
and \U$17951 ( \18083 , \17961 , \17965 );
and \U$17952 ( \18084 , \17965 , \17970 );
and \U$17953 ( \18085 , \17961 , \17970 );
or \U$17954 ( \18086 , \18083 , \18084 , \18085 );
xor \U$17955 ( \18087 , \18082 , \18086 );
xor \U$17956 ( \18088 , \18073 , \18087 );
and \U$17957 ( \18089 , \10584 , \2400 );
not \U$17958 ( \18090 , \18089 );
xnor \U$17959 ( \18091 , \18090 , \2195 );
and \U$17960 ( \18092 , \9897 , \2669 );
and \U$17961 ( \18093 , \10206 , \2538 );
nor \U$17962 ( \18094 , \18092 , \18093 );
xnor \U$17963 ( \18095 , \18094 , \2534 );
xor \U$17964 ( \18096 , \18091 , \18095 );
and \U$17965 ( \18097 , \9169 , \3103 );
and \U$17966 ( \18098 , \9465 , \2934 );
nor \U$17967 ( \18099 , \18097 , \18098 );
xnor \U$17968 ( \18100 , \18099 , \2839 );
xor \U$17969 ( \18101 , \18096 , \18100 );
and \U$17970 ( \18102 , \6945 , \4581 );
and \U$17971 ( \18103 , \7231 , \4424 );
nor \U$17972 ( \18104 , \18102 , \18103 );
xnor \U$17973 ( \18105 , \18104 , \4377 );
and \U$17974 ( \18106 , \6514 , \5011 );
and \U$17975 ( \18107 , \6790 , \4878 );
nor \U$17976 ( \18108 , \18106 , \18107 );
xnor \U$17977 ( \18109 , \18108 , \4762 );
xor \U$17978 ( \18110 , \18105 , \18109 );
and \U$17979 ( \18111 , \6030 , \5485 );
and \U$17980 ( \18112 , \6281 , \5275 );
nor \U$17981 ( \18113 , \18111 , \18112 );
xnor \U$17982 ( \18114 , \18113 , \5169 );
xor \U$17983 ( \18115 , \18110 , \18114 );
and \U$17984 ( \18116 , \5469 , \5996 );
and \U$17985 ( \18117 , \5674 , \5695 );
nor \U$17986 ( \18118 , \18116 , \18117 );
xnor \U$17987 ( \18119 , \18118 , \5687 );
and \U$17988 ( \18120 , \4922 , \6401 );
and \U$17989 ( \18121 , \5156 , \6143 );
nor \U$17990 ( \18122 , \18120 , \18121 );
xnor \U$17991 ( \18123 , \18122 , \6148 );
xor \U$17992 ( \18124 , \18119 , \18123 );
and \U$17993 ( \18125 , \4654 , \7055 );
and \U$17994 ( \18126 , \4749 , \6675 );
nor \U$17995 ( \18127 , \18125 , \18126 );
xnor \U$17996 ( \18128 , \18127 , \6680 );
xor \U$17997 ( \18129 , \18124 , \18128 );
xor \U$17998 ( \18130 , \18115 , \18129 );
and \U$17999 ( \18131 , \4160 , \7489 );
and \U$18000 ( \18132 , \4364 , \7137 );
nor \U$18001 ( \18133 , \18131 , \18132 );
xnor \U$18002 ( \18134 , \18133 , \7142 );
and \U$18003 ( \18135 , \3736 , \8019 );
and \U$18004 ( \18136 , \3912 , \7830 );
nor \U$18005 ( \18137 , \18135 , \18136 );
xnor \U$18006 ( \18138 , \18137 , \7713 );
xor \U$18007 ( \18139 , \18134 , \18138 );
and \U$18008 ( \18140 , \3395 , \8540 );
and \U$18009 ( \18141 , \3646 , \8292 );
nor \U$18010 ( \18142 , \18140 , \18141 );
xnor \U$18011 ( \18143 , \18142 , \8297 );
xor \U$18012 ( \18144 , \18139 , \18143 );
xor \U$18013 ( \18145 , \18130 , \18144 );
xor \U$18014 ( \18146 , \18101 , \18145 );
and \U$18015 ( \18147 , \2182 , \10118 );
and \U$18016 ( \18148 , \3037 , \9333 );
and \U$18017 ( \18149 , \3143 , \9006 );
nor \U$18018 ( \18150 , \18148 , \18149 );
xnor \U$18019 ( \18151 , \18150 , \8848 );
and \U$18020 ( \18152 , \2757 , \9765 );
and \U$18021 ( \18153 , \2826 , \9644 );
nor \U$18022 ( \18154 , \18152 , \18153 );
xnor \U$18023 ( \18155 , \18154 , \9478 );
xor \U$18024 ( \18156 , \18151 , \18155 );
and \U$18025 ( \18157 , \2366 , \10408 );
and \U$18026 ( \18158 , \2521 , \10116 );
nor \U$18027 ( \18159 , \18157 , \18158 );
xnor \U$18028 ( \18160 , \18159 , \10121 );
xor \U$18029 ( \18161 , \18156 , \18160 );
xnor \U$18030 ( \18162 , \18147 , \18161 );
xor \U$18031 ( \18163 , \18146 , \18162 );
xor \U$18032 ( \18164 , \18088 , \18163 );
xor \U$18033 ( \18165 , \18059 , \18164 );
xor \U$18034 ( \18166 , \18030 , \18165 );
xor \U$18035 ( \18167 , \18024 , \18166 );
and \U$18036 ( \18168 , \17794 , \17798 );
and \U$18037 ( \18169 , \17798 , \17976 );
and \U$18038 ( \18170 , \17794 , \17976 );
or \U$18039 ( \18171 , \18168 , \18169 , \18170 );
xor \U$18040 ( \18172 , \18167 , \18171 );
and \U$18041 ( \18173 , \17977 , \17978 );
and \U$18042 ( \18174 , \17979 , \17982 );
or \U$18043 ( \18175 , \18173 , \18174 );
xor \U$18044 ( \18176 , \18172 , \18175 );
buf \U$18045 ( \18177 , \18176 );
buf \U$18046 ( \18178 , \18177 );
and \U$18047 ( \18179 , \18028 , \18029 );
and \U$18048 ( \18180 , \18029 , \18165 );
and \U$18049 ( \18181 , \18028 , \18165 );
or \U$18050 ( \18182 , \18179 , \18180 , \18181 );
and \U$18051 ( \18183 , \17993 , \17997 );
and \U$18052 ( \18184 , \17997 , \18022 );
and \U$18053 ( \18185 , \17993 , \18022 );
or \U$18054 ( \18186 , \18183 , \18184 , \18185 );
and \U$18055 ( \18187 , \18044 , \18058 );
and \U$18056 ( \18188 , \18058 , \18164 );
and \U$18057 ( \18189 , \18044 , \18164 );
or \U$18058 ( \18190 , \18187 , \18188 , \18189 );
xor \U$18059 ( \18191 , \18186 , \18190 );
and \U$18060 ( \18192 , \18034 , \18038 );
and \U$18061 ( \18193 , \18038 , \18043 );
and \U$18062 ( \18194 , \18034 , \18043 );
or \U$18063 ( \18195 , \18192 , \18193 , \18194 );
and \U$18064 ( \18196 , \18002 , \18006 );
and \U$18065 ( \18197 , \18006 , \18021 );
and \U$18066 ( \18198 , \18002 , \18021 );
or \U$18067 ( \18199 , \18196 , \18197 , \18198 );
xor \U$18068 ( \18200 , \18195 , \18199 );
and \U$18069 ( \18201 , \18101 , \18145 );
and \U$18070 ( \18202 , \18145 , \18162 );
and \U$18071 ( \18203 , \18101 , \18162 );
or \U$18072 ( \18204 , \18201 , \18202 , \18203 );
xor \U$18073 ( \18205 , \18200 , \18204 );
xor \U$18074 ( \18206 , \18191 , \18205 );
xor \U$18075 ( \18207 , \18182 , \18206 );
and \U$18076 ( \18208 , \18048 , \18052 );
and \U$18077 ( \18209 , \18052 , \18057 );
and \U$18078 ( \18210 , \18048 , \18057 );
or \U$18079 ( \18211 , \18208 , \18209 , \18210 );
and \U$18080 ( \18212 , \18073 , \18087 );
and \U$18081 ( \18213 , \18087 , \18163 );
and \U$18082 ( \18214 , \18073 , \18163 );
or \U$18083 ( \18215 , \18212 , \18213 , \18214 );
xor \U$18084 ( \18216 , \18211 , \18215 );
and \U$18085 ( \18217 , \18063 , \18067 );
and \U$18086 ( \18218 , \18067 , \18072 );
and \U$18087 ( \18219 , \18063 , \18072 );
or \U$18088 ( \18220 , \18217 , \18218 , \18219 );
and \U$18089 ( \18221 , \18077 , \18081 );
and \U$18090 ( \18222 , \18081 , \18086 );
and \U$18091 ( \18223 , \18077 , \18086 );
or \U$18092 ( \18224 , \18221 , \18222 , \18223 );
xor \U$18093 ( \18225 , \18220 , \18224 );
or \U$18094 ( \18226 , \18147 , \18161 );
xor \U$18095 ( \18227 , \18225 , \18226 );
and \U$18096 ( \18228 , \18115 , \18129 );
and \U$18097 ( \18229 , \18129 , \18144 );
and \U$18098 ( \18230 , \18115 , \18144 );
or \U$18099 ( \18231 , \18228 , \18229 , \18230 );
not \U$18100 ( \18232 , \2195 );
and \U$18101 ( \18233 , \10206 , \2669 );
and \U$18102 ( \18234 , \10584 , \2538 );
nor \U$18103 ( \18235 , \18233 , \18234 );
xnor \U$18104 ( \18236 , \18235 , \2534 );
xor \U$18105 ( \18237 , \18232 , \18236 );
and \U$18106 ( \18238 , \9465 , \3103 );
and \U$18107 ( \18239 , \9897 , \2934 );
nor \U$18108 ( \18240 , \18238 , \18239 );
xnor \U$18109 ( \18241 , \18240 , \2839 );
xor \U$18110 ( \18242 , \18237 , \18241 );
xor \U$18111 ( \18243 , \18231 , \18242 );
and \U$18112 ( \18244 , \7231 , \4581 );
and \U$18113 ( \18245 , \7556 , \4424 );
nor \U$18114 ( \18246 , \18244 , \18245 );
xnor \U$18115 ( \18247 , \18246 , \4377 );
and \U$18116 ( \18248 , \6790 , \5011 );
and \U$18117 ( \18249 , \6945 , \4878 );
nor \U$18118 ( \18250 , \18248 , \18249 );
xnor \U$18119 ( \18251 , \18250 , \4762 );
xor \U$18120 ( \18252 , \18247 , \18251 );
and \U$18121 ( \18253 , \6281 , \5485 );
and \U$18122 ( \18254 , \6514 , \5275 );
nor \U$18123 ( \18255 , \18253 , \18254 );
xnor \U$18124 ( \18256 , \18255 , \5169 );
xor \U$18125 ( \18257 , \18252 , \18256 );
and \U$18126 ( \18258 , \5674 , \5996 );
and \U$18127 ( \18259 , \6030 , \5695 );
nor \U$18128 ( \18260 , \18258 , \18259 );
xnor \U$18129 ( \18261 , \18260 , \5687 );
and \U$18130 ( \18262 , \5156 , \6401 );
and \U$18131 ( \18263 , \5469 , \6143 );
nor \U$18132 ( \18264 , \18262 , \18263 );
xnor \U$18133 ( \18265 , \18264 , \6148 );
xor \U$18134 ( \18266 , \18261 , \18265 );
and \U$18135 ( \18267 , \4749 , \7055 );
and \U$18136 ( \18268 , \4922 , \6675 );
nor \U$18137 ( \18269 , \18267 , \18268 );
xnor \U$18138 ( \18270 , \18269 , \6680 );
xor \U$18139 ( \18271 , \18266 , \18270 );
xor \U$18140 ( \18272 , \18257 , \18271 );
and \U$18141 ( \18273 , \8835 , \3357 );
and \U$18142 ( \18274 , \9169 , \3255 );
nor \U$18143 ( \18275 , \18273 , \18274 );
xnor \U$18144 ( \18276 , \18275 , \3156 );
and \U$18145 ( \18277 , \8349 , \3813 );
and \U$18146 ( \18278 , \8652 , \3557 );
nor \U$18147 ( \18279 , \18277 , \18278 );
xnor \U$18148 ( \18280 , \18279 , \3562 );
xor \U$18149 ( \18281 , \18276 , \18280 );
and \U$18150 ( \18282 , \7700 , \4132 );
and \U$18151 ( \18283 , \8057 , \4012 );
nor \U$18152 ( \18284 , \18282 , \18283 );
xnor \U$18153 ( \18285 , \18284 , \3925 );
xor \U$18154 ( \18286 , \18281 , \18285 );
xor \U$18155 ( \18287 , \18272 , \18286 );
xor \U$18156 ( \18288 , \18243 , \18287 );
xor \U$18157 ( \18289 , \18227 , \18288 );
and \U$18158 ( \18290 , \18105 , \18109 );
and \U$18159 ( \18291 , \18109 , \18114 );
and \U$18160 ( \18292 , \18105 , \18114 );
or \U$18161 ( \18293 , \18290 , \18291 , \18292 );
and \U$18162 ( \18294 , \18011 , \18015 );
and \U$18163 ( \18295 , \18015 , \18020 );
and \U$18164 ( \18296 , \18011 , \18020 );
or \U$18165 ( \18297 , \18294 , \18295 , \18296 );
xor \U$18166 ( \18298 , \18293 , \18297 );
and \U$18167 ( \18299 , \18091 , \18095 );
and \U$18168 ( \18300 , \18095 , \18100 );
and \U$18169 ( \18301 , \18091 , \18100 );
or \U$18170 ( \18302 , \18299 , \18300 , \18301 );
xor \U$18171 ( \18303 , \18298 , \18302 );
and \U$18172 ( \18304 , \18119 , \18123 );
and \U$18173 ( \18305 , \18123 , \18128 );
and \U$18174 ( \18306 , \18119 , \18128 );
or \U$18175 ( \18307 , \18304 , \18305 , \18306 );
and \U$18176 ( \18308 , \18151 , \18155 );
and \U$18177 ( \18309 , \18155 , \18160 );
and \U$18178 ( \18310 , \18151 , \18160 );
or \U$18179 ( \18311 , \18308 , \18309 , \18310 );
xor \U$18180 ( \18312 , \18307 , \18311 );
and \U$18181 ( \18313 , \18134 , \18138 );
and \U$18182 ( \18314 , \18138 , \18143 );
and \U$18183 ( \18315 , \18134 , \18143 );
or \U$18184 ( \18316 , \18313 , \18314 , \18315 );
xor \U$18185 ( \18317 , \18312 , \18316 );
xor \U$18186 ( \18318 , \18303 , \18317 );
and \U$18187 ( \18319 , \2366 , \10118 );
and \U$18188 ( \18320 , \3143 , \9333 );
and \U$18189 ( \18321 , \3395 , \9006 );
nor \U$18190 ( \18322 , \18320 , \18321 );
xnor \U$18191 ( \18323 , \18322 , \8848 );
and \U$18192 ( \18324 , \2826 , \9765 );
and \U$18193 ( \18325 , \3037 , \9644 );
nor \U$18194 ( \18326 , \18324 , \18325 );
xnor \U$18195 ( \18327 , \18326 , \9478 );
xor \U$18196 ( \18328 , \18323 , \18327 );
and \U$18197 ( \18329 , \2521 , \10408 );
and \U$18198 ( \18330 , \2757 , \10116 );
nor \U$18199 ( \18331 , \18329 , \18330 );
xnor \U$18200 ( \18332 , \18331 , \10121 );
xor \U$18201 ( \18333 , \18328 , \18332 );
xor \U$18202 ( \18334 , \18319 , \18333 );
and \U$18203 ( \18335 , \4364 , \7489 );
and \U$18204 ( \18336 , \4654 , \7137 );
nor \U$18205 ( \18337 , \18335 , \18336 );
xnor \U$18206 ( \18338 , \18337 , \7142 );
and \U$18207 ( \18339 , \3912 , \8019 );
and \U$18208 ( \18340 , \4160 , \7830 );
nor \U$18209 ( \18341 , \18339 , \18340 );
xnor \U$18210 ( \18342 , \18341 , \7713 );
xor \U$18211 ( \18343 , \18338 , \18342 );
and \U$18212 ( \18344 , \3646 , \8540 );
and \U$18213 ( \18345 , \3736 , \8292 );
nor \U$18214 ( \18346 , \18344 , \18345 );
xnor \U$18215 ( \18347 , \18346 , \8297 );
xor \U$18216 ( \18348 , \18343 , \18347 );
xor \U$18217 ( \18349 , \18334 , \18348 );
xor \U$18218 ( \18350 , \18318 , \18349 );
xor \U$18219 ( \18351 , \18289 , \18350 );
xor \U$18220 ( \18352 , \18216 , \18351 );
xor \U$18221 ( \18353 , \18207 , \18352 );
and \U$18222 ( \18354 , \17989 , \18023 );
and \U$18223 ( \18355 , \18023 , \18166 );
and \U$18224 ( \18356 , \17989 , \18166 );
or \U$18225 ( \18357 , \18354 , \18355 , \18356 );
xor \U$18226 ( \18358 , \18353 , \18357 );
and \U$18227 ( \18359 , \18167 , \18171 );
and \U$18228 ( \18360 , \18172 , \18175 );
or \U$18229 ( \18361 , \18359 , \18360 );
xor \U$18230 ( \18362 , \18358 , \18361 );
buf \U$18231 ( \18363 , \18362 );
buf \U$18232 ( \18364 , \18363 );
and \U$18233 ( \18365 , \18186 , \18190 );
and \U$18234 ( \18366 , \18190 , \18205 );
and \U$18235 ( \18367 , \18186 , \18205 );
or \U$18236 ( \18368 , \18365 , \18366 , \18367 );
and \U$18237 ( \18369 , \18211 , \18215 );
and \U$18238 ( \18370 , \18215 , \18351 );
and \U$18239 ( \18371 , \18211 , \18351 );
or \U$18240 ( \18372 , \18369 , \18370 , \18371 );
and \U$18241 ( \18373 , \18220 , \18224 );
and \U$18242 ( \18374 , \18224 , \18226 );
and \U$18243 ( \18375 , \18220 , \18226 );
or \U$18244 ( \18376 , \18373 , \18374 , \18375 );
and \U$18245 ( \18377 , \18231 , \18242 );
and \U$18246 ( \18378 , \18242 , \18287 );
and \U$18247 ( \18379 , \18231 , \18287 );
or \U$18248 ( \18380 , \18377 , \18378 , \18379 );
xor \U$18249 ( \18381 , \18376 , \18380 );
and \U$18250 ( \18382 , \18303 , \18317 );
and \U$18251 ( \18383 , \18317 , \18349 );
and \U$18252 ( \18384 , \18303 , \18349 );
or \U$18253 ( \18385 , \18382 , \18383 , \18384 );
xor \U$18254 ( \18386 , \18381 , \18385 );
xor \U$18255 ( \18387 , \18372 , \18386 );
and \U$18256 ( \18388 , \18195 , \18199 );
and \U$18257 ( \18389 , \18199 , \18204 );
and \U$18258 ( \18390 , \18195 , \18204 );
or \U$18259 ( \18391 , \18388 , \18389 , \18390 );
and \U$18260 ( \18392 , \18227 , \18288 );
and \U$18261 ( \18393 , \18288 , \18350 );
and \U$18262 ( \18394 , \18227 , \18350 );
or \U$18263 ( \18395 , \18392 , \18393 , \18394 );
xor \U$18264 ( \18396 , \18391 , \18395 );
and \U$18265 ( \18397 , \18293 , \18297 );
and \U$18266 ( \18398 , \18297 , \18302 );
and \U$18267 ( \18399 , \18293 , \18302 );
or \U$18268 ( \18400 , \18397 , \18398 , \18399 );
and \U$18269 ( \18401 , \18307 , \18311 );
and \U$18270 ( \18402 , \18311 , \18316 );
and \U$18271 ( \18403 , \18307 , \18316 );
or \U$18272 ( \18404 , \18401 , \18402 , \18403 );
xor \U$18273 ( \18405 , \18400 , \18404 );
and \U$18274 ( \18406 , \18319 , \18333 );
and \U$18275 ( \18407 , \18333 , \18348 );
and \U$18276 ( \18408 , \18319 , \18348 );
or \U$18277 ( \18409 , \18406 , \18407 , \18408 );
xor \U$18278 ( \18410 , \18405 , \18409 );
and \U$18279 ( \18411 , \18257 , \18271 );
and \U$18280 ( \18412 , \18271 , \18286 );
and \U$18281 ( \18413 , \18257 , \18286 );
or \U$18282 ( \18414 , \18411 , \18412 , \18413 );
and \U$18283 ( \18415 , \10584 , \2669 );
not \U$18284 ( \18416 , \18415 );
xnor \U$18285 ( \18417 , \18416 , \2534 );
and \U$18286 ( \18418 , \9897 , \3103 );
and \U$18287 ( \18419 , \10206 , \2934 );
nor \U$18288 ( \18420 , \18418 , \18419 );
xnor \U$18289 ( \18421 , \18420 , \2839 );
xor \U$18290 ( \18422 , \18417 , \18421 );
and \U$18291 ( \18423 , \9169 , \3357 );
and \U$18292 ( \18424 , \9465 , \3255 );
nor \U$18293 ( \18425 , \18423 , \18424 );
xnor \U$18294 ( \18426 , \18425 , \3156 );
xor \U$18295 ( \18427 , \18422 , \18426 );
xor \U$18296 ( \18428 , \18414 , \18427 );
and \U$18297 ( \18429 , \8652 , \3813 );
and \U$18298 ( \18430 , \8835 , \3557 );
nor \U$18299 ( \18431 , \18429 , \18430 );
xnor \U$18300 ( \18432 , \18431 , \3562 );
and \U$18301 ( \18433 , \8057 , \4132 );
and \U$18302 ( \18434 , \8349 , \4012 );
nor \U$18303 ( \18435 , \18433 , \18434 );
xnor \U$18304 ( \18436 , \18435 , \3925 );
xor \U$18305 ( \18437 , \18432 , \18436 );
and \U$18306 ( \18438 , \7556 , \4581 );
and \U$18307 ( \18439 , \7700 , \4424 );
nor \U$18308 ( \18440 , \18438 , \18439 );
xnor \U$18309 ( \18441 , \18440 , \4377 );
xor \U$18310 ( \18442 , \18437 , \18441 );
and \U$18311 ( \18443 , \6945 , \5011 );
and \U$18312 ( \18444 , \7231 , \4878 );
nor \U$18313 ( \18445 , \18443 , \18444 );
xnor \U$18314 ( \18446 , \18445 , \4762 );
and \U$18315 ( \18447 , \6514 , \5485 );
and \U$18316 ( \18448 , \6790 , \5275 );
nor \U$18317 ( \18449 , \18447 , \18448 );
xnor \U$18318 ( \18450 , \18449 , \5169 );
xor \U$18319 ( \18451 , \18446 , \18450 );
and \U$18320 ( \18452 , \6030 , \5996 );
and \U$18321 ( \18453 , \6281 , \5695 );
nor \U$18322 ( \18454 , \18452 , \18453 );
xnor \U$18323 ( \18455 , \18454 , \5687 );
xor \U$18324 ( \18456 , \18451 , \18455 );
xor \U$18325 ( \18457 , \18442 , \18456 );
and \U$18326 ( \18458 , \5469 , \6401 );
and \U$18327 ( \18459 , \5674 , \6143 );
nor \U$18328 ( \18460 , \18458 , \18459 );
xnor \U$18329 ( \18461 , \18460 , \6148 );
and \U$18330 ( \18462 , \4922 , \7055 );
and \U$18331 ( \18463 , \5156 , \6675 );
nor \U$18332 ( \18464 , \18462 , \18463 );
xnor \U$18333 ( \18465 , \18464 , \6680 );
xor \U$18334 ( \18466 , \18461 , \18465 );
and \U$18335 ( \18467 , \4654 , \7489 );
and \U$18336 ( \18468 , \4749 , \7137 );
nor \U$18337 ( \18469 , \18467 , \18468 );
xnor \U$18338 ( \18470 , \18469 , \7142 );
xor \U$18339 ( \18471 , \18466 , \18470 );
xor \U$18340 ( \18472 , \18457 , \18471 );
xor \U$18341 ( \18473 , \18428 , \18472 );
xor \U$18342 ( \18474 , \18410 , \18473 );
and \U$18343 ( \18475 , \18247 , \18251 );
and \U$18344 ( \18476 , \18251 , \18256 );
and \U$18345 ( \18477 , \18247 , \18256 );
or \U$18346 ( \18478 , \18475 , \18476 , \18477 );
and \U$18347 ( \18479 , \18232 , \18236 );
and \U$18348 ( \18480 , \18236 , \18241 );
and \U$18349 ( \18481 , \18232 , \18241 );
or \U$18350 ( \18482 , \18479 , \18480 , \18481 );
xor \U$18351 ( \18483 , \18478 , \18482 );
and \U$18352 ( \18484 , \18276 , \18280 );
and \U$18353 ( \18485 , \18280 , \18285 );
and \U$18354 ( \18486 , \18276 , \18285 );
or \U$18355 ( \18487 , \18484 , \18485 , \18486 );
xor \U$18356 ( \18488 , \18483 , \18487 );
and \U$18357 ( \18489 , \18323 , \18327 );
and \U$18358 ( \18490 , \18327 , \18332 );
and \U$18359 ( \18491 , \18323 , \18332 );
or \U$18360 ( \18492 , \18489 , \18490 , \18491 );
and \U$18361 ( \18493 , \18261 , \18265 );
and \U$18362 ( \18494 , \18265 , \18270 );
and \U$18363 ( \18495 , \18261 , \18270 );
or \U$18364 ( \18496 , \18493 , \18494 , \18495 );
xor \U$18365 ( \18497 , \18492 , \18496 );
and \U$18366 ( \18498 , \18338 , \18342 );
and \U$18367 ( \18499 , \18342 , \18347 );
and \U$18368 ( \18500 , \18338 , \18347 );
or \U$18369 ( \18501 , \18498 , \18499 , \18500 );
xor \U$18370 ( \18502 , \18497 , \18501 );
xor \U$18371 ( \18503 , \18488 , \18502 );
and \U$18372 ( \18504 , \3037 , \9765 );
and \U$18373 ( \18505 , \3143 , \9644 );
nor \U$18374 ( \18506 , \18504 , \18505 );
xnor \U$18375 ( \18507 , \18506 , \9478 );
and \U$18376 ( \18508 , \2757 , \10408 );
and \U$18377 ( \18509 , \2826 , \10116 );
nor \U$18378 ( \18510 , \18508 , \18509 );
xnor \U$18379 ( \18511 , \18510 , \10121 );
xor \U$18380 ( \18512 , \18507 , \18511 );
and \U$18381 ( \18513 , \2521 , \10118 );
xor \U$18382 ( \18514 , \18512 , \18513 );
and \U$18383 ( \18515 , \4160 , \8019 );
and \U$18384 ( \18516 , \4364 , \7830 );
nor \U$18385 ( \18517 , \18515 , \18516 );
xnor \U$18386 ( \18518 , \18517 , \7713 );
and \U$18387 ( \18519 , \3736 , \8540 );
and \U$18388 ( \18520 , \3912 , \8292 );
nor \U$18389 ( \18521 , \18519 , \18520 );
xnor \U$18390 ( \18522 , \18521 , \8297 );
xor \U$18391 ( \18523 , \18518 , \18522 );
and \U$18392 ( \18524 , \3395 , \9333 );
and \U$18393 ( \18525 , \3646 , \9006 );
nor \U$18394 ( \18526 , \18524 , \18525 );
xnor \U$18395 ( \18527 , \18526 , \8848 );
xor \U$18396 ( \18528 , \18523 , \18527 );
xnor \U$18397 ( \18529 , \18514 , \18528 );
xor \U$18398 ( \18530 , \18503 , \18529 );
xor \U$18399 ( \18531 , \18474 , \18530 );
xor \U$18400 ( \18532 , \18396 , \18531 );
xor \U$18401 ( \18533 , \18387 , \18532 );
xor \U$18402 ( \18534 , \18368 , \18533 );
and \U$18403 ( \18535 , \18182 , \18206 );
and \U$18404 ( \18536 , \18206 , \18352 );
and \U$18405 ( \18537 , \18182 , \18352 );
or \U$18406 ( \18538 , \18535 , \18536 , \18537 );
xor \U$18407 ( \18539 , \18534 , \18538 );
and \U$18408 ( \18540 , \18353 , \18357 );
and \U$18409 ( \18541 , \18358 , \18361 );
or \U$18410 ( \18542 , \18540 , \18541 );
xor \U$18411 ( \18543 , \18539 , \18542 );
buf \U$18412 ( \18544 , \18543 );
buf \U$18413 ( \18545 , \18544 );
and \U$18414 ( \18546 , \18372 , \18386 );
and \U$18415 ( \18547 , \18386 , \18532 );
and \U$18416 ( \18548 , \18372 , \18532 );
or \U$18417 ( \18549 , \18546 , \18547 , \18548 );
and \U$18418 ( \18550 , \18391 , \18395 );
and \U$18419 ( \18551 , \18395 , \18531 );
and \U$18420 ( \18552 , \18391 , \18531 );
or \U$18421 ( \18553 , \18550 , \18551 , \18552 );
and \U$18422 ( \18554 , \18400 , \18404 );
and \U$18423 ( \18555 , \18404 , \18409 );
and \U$18424 ( \18556 , \18400 , \18409 );
or \U$18425 ( \18557 , \18554 , \18555 , \18556 );
and \U$18426 ( \18558 , \18414 , \18427 );
and \U$18427 ( \18559 , \18427 , \18472 );
and \U$18428 ( \18560 , \18414 , \18472 );
or \U$18429 ( \18561 , \18558 , \18559 , \18560 );
xor \U$18430 ( \18562 , \18557 , \18561 );
and \U$18431 ( \18563 , \18488 , \18502 );
and \U$18432 ( \18564 , \18502 , \18529 );
and \U$18433 ( \18565 , \18488 , \18529 );
or \U$18434 ( \18566 , \18563 , \18564 , \18565 );
xor \U$18435 ( \18567 , \18562 , \18566 );
xor \U$18436 ( \18568 , \18553 , \18567 );
and \U$18437 ( \18569 , \18376 , \18380 );
and \U$18438 ( \18570 , \18380 , \18385 );
and \U$18439 ( \18571 , \18376 , \18385 );
or \U$18440 ( \18572 , \18569 , \18570 , \18571 );
and \U$18441 ( \18573 , \18410 , \18473 );
and \U$18442 ( \18574 , \18473 , \18530 );
and \U$18443 ( \18575 , \18410 , \18530 );
or \U$18444 ( \18576 , \18573 , \18574 , \18575 );
xor \U$18445 ( \18577 , \18572 , \18576 );
and \U$18446 ( \18578 , \18478 , \18482 );
and \U$18447 ( \18579 , \18482 , \18487 );
and \U$18448 ( \18580 , \18478 , \18487 );
or \U$18449 ( \18581 , \18578 , \18579 , \18580 );
and \U$18450 ( \18582 , \18492 , \18496 );
and \U$18451 ( \18583 , \18496 , \18501 );
and \U$18452 ( \18584 , \18492 , \18501 );
or \U$18453 ( \18585 , \18582 , \18583 , \18584 );
xor \U$18454 ( \18586 , \18581 , \18585 );
or \U$18455 ( \18587 , \18514 , \18528 );
xor \U$18456 ( \18588 , \18586 , \18587 );
and \U$18457 ( \18589 , \18442 , \18456 );
and \U$18458 ( \18590 , \18456 , \18471 );
and \U$18459 ( \18591 , \18442 , \18471 );
or \U$18460 ( \18592 , \18589 , \18590 , \18591 );
and \U$18461 ( \18593 , \3143 , \9765 );
and \U$18462 ( \18594 , \3395 , \9644 );
nor \U$18463 ( \18595 , \18593 , \18594 );
xnor \U$18464 ( \18596 , \18595 , \9478 );
and \U$18465 ( \18597 , \2826 , \10408 );
and \U$18466 ( \18598 , \3037 , \10116 );
nor \U$18467 ( \18599 , \18597 , \18598 );
xnor \U$18468 ( \18600 , \18599 , \10121 );
xor \U$18469 ( \18601 , \18596 , \18600 );
and \U$18470 ( \18602 , \2757 , \10118 );
xor \U$18471 ( \18603 , \18601 , \18602 );
and \U$18472 ( \18604 , \4364 , \8019 );
and \U$18473 ( \18605 , \4654 , \7830 );
nor \U$18474 ( \18606 , \18604 , \18605 );
xnor \U$18475 ( \18607 , \18606 , \7713 );
and \U$18476 ( \18608 , \3912 , \8540 );
and \U$18477 ( \18609 , \4160 , \8292 );
nor \U$18478 ( \18610 , \18608 , \18609 );
xnor \U$18479 ( \18611 , \18610 , \8297 );
xor \U$18480 ( \18612 , \18607 , \18611 );
and \U$18481 ( \18613 , \3646 , \9333 );
and \U$18482 ( \18614 , \3736 , \9006 );
nor \U$18483 ( \18615 , \18613 , \18614 );
xnor \U$18484 ( \18616 , \18615 , \8848 );
xor \U$18485 ( \18617 , \18612 , \18616 );
xor \U$18486 ( \18618 , \18603 , \18617 );
and \U$18487 ( \18619 , \5674 , \6401 );
and \U$18488 ( \18620 , \6030 , \6143 );
nor \U$18489 ( \18621 , \18619 , \18620 );
xnor \U$18490 ( \18622 , \18621 , \6148 );
and \U$18491 ( \18623 , \5156 , \7055 );
and \U$18492 ( \18624 , \5469 , \6675 );
nor \U$18493 ( \18625 , \18623 , \18624 );
xnor \U$18494 ( \18626 , \18625 , \6680 );
xor \U$18495 ( \18627 , \18622 , \18626 );
and \U$18496 ( \18628 , \4749 , \7489 );
and \U$18497 ( \18629 , \4922 , \7137 );
nor \U$18498 ( \18630 , \18628 , \18629 );
xnor \U$18499 ( \18631 , \18630 , \7142 );
xor \U$18500 ( \18632 , \18627 , \18631 );
xor \U$18501 ( \18633 , \18618 , \18632 );
xor \U$18502 ( \18634 , \18592 , \18633 );
and \U$18503 ( \18635 , \8835 , \3813 );
and \U$18504 ( \18636 , \9169 , \3557 );
nor \U$18505 ( \18637 , \18635 , \18636 );
xnor \U$18506 ( \18638 , \18637 , \3562 );
and \U$18507 ( \18639 , \8349 , \4132 );
and \U$18508 ( \18640 , \8652 , \4012 );
nor \U$18509 ( \18641 , \18639 , \18640 );
xnor \U$18510 ( \18642 , \18641 , \3925 );
xor \U$18511 ( \18643 , \18638 , \18642 );
and \U$18512 ( \18644 , \7700 , \4581 );
and \U$18513 ( \18645 , \8057 , \4424 );
nor \U$18514 ( \18646 , \18644 , \18645 );
xnor \U$18515 ( \18647 , \18646 , \4377 );
xor \U$18516 ( \18648 , \18643 , \18647 );
and \U$18517 ( \18649 , \7231 , \5011 );
and \U$18518 ( \18650 , \7556 , \4878 );
nor \U$18519 ( \18651 , \18649 , \18650 );
xnor \U$18520 ( \18652 , \18651 , \4762 );
and \U$18521 ( \18653 , \6790 , \5485 );
and \U$18522 ( \18654 , \6945 , \5275 );
nor \U$18523 ( \18655 , \18653 , \18654 );
xnor \U$18524 ( \18656 , \18655 , \5169 );
xor \U$18525 ( \18657 , \18652 , \18656 );
and \U$18526 ( \18658 , \6281 , \5996 );
and \U$18527 ( \18659 , \6514 , \5695 );
nor \U$18528 ( \18660 , \18658 , \18659 );
xnor \U$18529 ( \18661 , \18660 , \5687 );
xor \U$18530 ( \18662 , \18657 , \18661 );
xor \U$18531 ( \18663 , \18648 , \18662 );
not \U$18532 ( \18664 , \2534 );
and \U$18533 ( \18665 , \10206 , \3103 );
and \U$18534 ( \18666 , \10584 , \2934 );
nor \U$18535 ( \18667 , \18665 , \18666 );
xnor \U$18536 ( \18668 , \18667 , \2839 );
xor \U$18537 ( \18669 , \18664 , \18668 );
and \U$18538 ( \18670 , \9465 , \3357 );
and \U$18539 ( \18671 , \9897 , \3255 );
nor \U$18540 ( \18672 , \18670 , \18671 );
xnor \U$18541 ( \18673 , \18672 , \3156 );
xor \U$18542 ( \18674 , \18669 , \18673 );
xor \U$18543 ( \18675 , \18663 , \18674 );
xor \U$18544 ( \18676 , \18634 , \18675 );
xor \U$18545 ( \18677 , \18588 , \18676 );
and \U$18546 ( \18678 , \18507 , \18511 );
and \U$18547 ( \18679 , \18511 , \18513 );
and \U$18548 ( \18680 , \18507 , \18513 );
or \U$18549 ( \18681 , \18678 , \18679 , \18680 );
and \U$18550 ( \18682 , \18518 , \18522 );
and \U$18551 ( \18683 , \18522 , \18527 );
and \U$18552 ( \18684 , \18518 , \18527 );
or \U$18553 ( \18685 , \18682 , \18683 , \18684 );
xor \U$18554 ( \18686 , \18681 , \18685 );
and \U$18555 ( \18687 , \18461 , \18465 );
and \U$18556 ( \18688 , \18465 , \18470 );
and \U$18557 ( \18689 , \18461 , \18470 );
or \U$18558 ( \18690 , \18687 , \18688 , \18689 );
xor \U$18559 ( \18691 , \18686 , \18690 );
and \U$18560 ( \18692 , \18432 , \18436 );
and \U$18561 ( \18693 , \18436 , \18441 );
and \U$18562 ( \18694 , \18432 , \18441 );
or \U$18563 ( \18695 , \18692 , \18693 , \18694 );
and \U$18564 ( \18696 , \18417 , \18421 );
and \U$18565 ( \18697 , \18421 , \18426 );
and \U$18566 ( \18698 , \18417 , \18426 );
or \U$18567 ( \18699 , \18696 , \18697 , \18698 );
xor \U$18568 ( \18700 , \18695 , \18699 );
and \U$18569 ( \18701 , \18446 , \18450 );
and \U$18570 ( \18702 , \18450 , \18455 );
and \U$18571 ( \18703 , \18446 , \18455 );
or \U$18572 ( \18704 , \18701 , \18702 , \18703 );
xor \U$18573 ( \18705 , \18700 , \18704 );
xor \U$18574 ( \18706 , \18691 , \18705 );
xor \U$18575 ( \18707 , \18677 , \18706 );
xor \U$18576 ( \18708 , \18577 , \18707 );
xor \U$18577 ( \18709 , \18568 , \18708 );
xor \U$18578 ( \18710 , \18549 , \18709 );
and \U$18579 ( \18711 , \18368 , \18533 );
xor \U$18580 ( \18712 , \18710 , \18711 );
and \U$18581 ( \18713 , \18534 , \18538 );
and \U$18582 ( \18714 , \18539 , \18542 );
or \U$18583 ( \18715 , \18713 , \18714 );
xor \U$18584 ( \18716 , \18712 , \18715 );
buf \U$18585 ( \18717 , \18716 );
buf \U$18586 ( \18718 , \18717 );
and \U$18587 ( \18719 , \18553 , \18567 );
and \U$18588 ( \18720 , \18567 , \18708 );
and \U$18589 ( \18721 , \18553 , \18708 );
or \U$18590 ( \18722 , \18719 , \18720 , \18721 );
and \U$18591 ( \18723 , \18572 , \18576 );
and \U$18592 ( \18724 , \18576 , \18707 );
and \U$18593 ( \18725 , \18572 , \18707 );
or \U$18594 ( \18726 , \18723 , \18724 , \18725 );
and \U$18595 ( \18727 , \18581 , \18585 );
and \U$18596 ( \18728 , \18585 , \18587 );
and \U$18597 ( \18729 , \18581 , \18587 );
or \U$18598 ( \18730 , \18727 , \18728 , \18729 );
and \U$18599 ( \18731 , \18592 , \18633 );
and \U$18600 ( \18732 , \18633 , \18675 );
and \U$18601 ( \18733 , \18592 , \18675 );
or \U$18602 ( \18734 , \18731 , \18732 , \18733 );
xor \U$18603 ( \18735 , \18730 , \18734 );
and \U$18604 ( \18736 , \18691 , \18705 );
xor \U$18605 ( \18737 , \18735 , \18736 );
xor \U$18606 ( \18738 , \18726 , \18737 );
and \U$18607 ( \18739 , \18557 , \18561 );
and \U$18608 ( \18740 , \18561 , \18566 );
and \U$18609 ( \18741 , \18557 , \18566 );
or \U$18610 ( \18742 , \18739 , \18740 , \18741 );
and \U$18611 ( \18743 , \18588 , \18676 );
and \U$18612 ( \18744 , \18676 , \18706 );
and \U$18613 ( \18745 , \18588 , \18706 );
or \U$18614 ( \18746 , \18743 , \18744 , \18745 );
xor \U$18615 ( \18747 , \18742 , \18746 );
and \U$18616 ( \18748 , \18681 , \18685 );
and \U$18617 ( \18749 , \18685 , \18690 );
and \U$18618 ( \18750 , \18681 , \18690 );
or \U$18619 ( \18751 , \18748 , \18749 , \18750 );
and \U$18620 ( \18752 , \18695 , \18699 );
and \U$18621 ( \18753 , \18699 , \18704 );
and \U$18622 ( \18754 , \18695 , \18704 );
or \U$18623 ( \18755 , \18752 , \18753 , \18754 );
xor \U$18624 ( \18756 , \18751 , \18755 );
and \U$18625 ( \18757 , \18603 , \18617 );
and \U$18626 ( \18758 , \18617 , \18632 );
and \U$18627 ( \18759 , \18603 , \18632 );
or \U$18628 ( \18760 , \18757 , \18758 , \18759 );
xor \U$18629 ( \18761 , \18756 , \18760 );
and \U$18630 ( \18762 , \18648 , \18662 );
and \U$18631 ( \18763 , \18662 , \18674 );
and \U$18632 ( \18764 , \18648 , \18674 );
or \U$18633 ( \18765 , \18762 , \18763 , \18764 );
and \U$18634 ( \18766 , \10584 , \3103 );
not \U$18635 ( \18767 , \18766 );
xnor \U$18636 ( \18768 , \18767 , \2839 );
and \U$18637 ( \18769 , \9897 , \3357 );
and \U$18638 ( \18770 , \10206 , \3255 );
nor \U$18639 ( \18771 , \18769 , \18770 );
xnor \U$18640 ( \18772 , \18771 , \3156 );
xor \U$18641 ( \18773 , \18768 , \18772 );
and \U$18642 ( \18774 , \9169 , \3813 );
and \U$18643 ( \18775 , \9465 , \3557 );
nor \U$18644 ( \18776 , \18774 , \18775 );
xnor \U$18645 ( \18777 , \18776 , \3562 );
xor \U$18646 ( \18778 , \18773 , \18777 );
and \U$18647 ( \18779 , \6945 , \5485 );
and \U$18648 ( \18780 , \7231 , \5275 );
nor \U$18649 ( \18781 , \18779 , \18780 );
xnor \U$18650 ( \18782 , \18781 , \5169 );
and \U$18651 ( \18783 , \6514 , \5996 );
and \U$18652 ( \18784 , \6790 , \5695 );
nor \U$18653 ( \18785 , \18783 , \18784 );
xnor \U$18654 ( \18786 , \18785 , \5687 );
xor \U$18655 ( \18787 , \18782 , \18786 );
and \U$18656 ( \18788 , \6030 , \6401 );
and \U$18657 ( \18789 , \6281 , \6143 );
nor \U$18658 ( \18790 , \18788 , \18789 );
xnor \U$18659 ( \18791 , \18790 , \6148 );
xor \U$18660 ( \18792 , \18787 , \18791 );
xor \U$18661 ( \18793 , \18778 , \18792 );
and \U$18662 ( \18794 , \8652 , \4132 );
and \U$18663 ( \18795 , \8835 , \4012 );
nor \U$18664 ( \18796 , \18794 , \18795 );
xnor \U$18665 ( \18797 , \18796 , \3925 );
and \U$18666 ( \18798 , \8057 , \4581 );
and \U$18667 ( \18799 , \8349 , \4424 );
nor \U$18668 ( \18800 , \18798 , \18799 );
xnor \U$18669 ( \18801 , \18800 , \4377 );
xor \U$18670 ( \18802 , \18797 , \18801 );
and \U$18671 ( \18803 , \7556 , \5011 );
and \U$18672 ( \18804 , \7700 , \4878 );
nor \U$18673 ( \18805 , \18803 , \18804 );
xnor \U$18674 ( \18806 , \18805 , \4762 );
xor \U$18675 ( \18807 , \18802 , \18806 );
xor \U$18676 ( \18808 , \18793 , \18807 );
xor \U$18677 ( \18809 , \18765 , \18808 );
and \U$18678 ( \18810 , \4160 , \8540 );
and \U$18679 ( \18811 , \4364 , \8292 );
nor \U$18680 ( \18812 , \18810 , \18811 );
xnor \U$18681 ( \18813 , \18812 , \8297 );
and \U$18682 ( \18814 , \3736 , \9333 );
and \U$18683 ( \18815 , \3912 , \9006 );
nor \U$18684 ( \18816 , \18814 , \18815 );
xnor \U$18685 ( \18817 , \18816 , \8848 );
xor \U$18686 ( \18818 , \18813 , \18817 );
and \U$18687 ( \18819 , \3395 , \9765 );
and \U$18688 ( \18820 , \3646 , \9644 );
nor \U$18689 ( \18821 , \18819 , \18820 );
xnor \U$18690 ( \18822 , \18821 , \9478 );
xor \U$18691 ( \18823 , \18818 , \18822 );
and \U$18692 ( \18824 , \5469 , \7055 );
and \U$18693 ( \18825 , \5674 , \6675 );
nor \U$18694 ( \18826 , \18824 , \18825 );
xnor \U$18695 ( \18827 , \18826 , \6680 );
and \U$18696 ( \18828 , \4922 , \7489 );
and \U$18697 ( \18829 , \5156 , \7137 );
nor \U$18698 ( \18830 , \18828 , \18829 );
xnor \U$18699 ( \18831 , \18830 , \7142 );
xor \U$18700 ( \18832 , \18827 , \18831 );
and \U$18701 ( \18833 , \4654 , \8019 );
and \U$18702 ( \18834 , \4749 , \7830 );
nor \U$18703 ( \18835 , \18833 , \18834 );
xnor \U$18704 ( \18836 , \18835 , \7713 );
xor \U$18705 ( \18837 , \18832 , \18836 );
xor \U$18706 ( \18838 , \18823 , \18837 );
and \U$18707 ( \18839 , \3037 , \10408 );
and \U$18708 ( \18840 , \3143 , \10116 );
nor \U$18709 ( \18841 , \18839 , \18840 );
xnor \U$18710 ( \18842 , \18841 , \10121 );
and \U$18711 ( \18843 , \2826 , \10118 );
xnor \U$18712 ( \18844 , \18842 , \18843 );
xor \U$18713 ( \18845 , \18838 , \18844 );
xor \U$18714 ( \18846 , \18809 , \18845 );
xor \U$18715 ( \18847 , \18761 , \18846 );
and \U$18716 ( \18848 , \18638 , \18642 );
and \U$18717 ( \18849 , \18642 , \18647 );
and \U$18718 ( \18850 , \18638 , \18647 );
or \U$18719 ( \18851 , \18848 , \18849 , \18850 );
and \U$18720 ( \18852 , \18652 , \18656 );
and \U$18721 ( \18853 , \18656 , \18661 );
and \U$18722 ( \18854 , \18652 , \18661 );
or \U$18723 ( \18855 , \18852 , \18853 , \18854 );
xor \U$18724 ( \18856 , \18851 , \18855 );
and \U$18725 ( \18857 , \18664 , \18668 );
and \U$18726 ( \18858 , \18668 , \18673 );
and \U$18727 ( \18859 , \18664 , \18673 );
or \U$18728 ( \18860 , \18857 , \18858 , \18859 );
xor \U$18729 ( \18861 , \18856 , \18860 );
and \U$18730 ( \18862 , \18596 , \18600 );
and \U$18731 ( \18863 , \18600 , \18602 );
and \U$18732 ( \18864 , \18596 , \18602 );
or \U$18733 ( \18865 , \18862 , \18863 , \18864 );
and \U$18734 ( \18866 , \18607 , \18611 );
and \U$18735 ( \18867 , \18611 , \18616 );
and \U$18736 ( \18868 , \18607 , \18616 );
or \U$18737 ( \18869 , \18866 , \18867 , \18868 );
xor \U$18738 ( \18870 , \18865 , \18869 );
and \U$18739 ( \18871 , \18622 , \18626 );
and \U$18740 ( \18872 , \18626 , \18631 );
and \U$18741 ( \18873 , \18622 , \18631 );
or \U$18742 ( \18874 , \18871 , \18872 , \18873 );
xor \U$18743 ( \18875 , \18870 , \18874 );
xor \U$18744 ( \18876 , \18861 , \18875 );
xor \U$18745 ( \18877 , \18847 , \18876 );
xor \U$18746 ( \18878 , \18747 , \18877 );
xor \U$18747 ( \18879 , \18738 , \18878 );
xor \U$18748 ( \18880 , \18722 , \18879 );
and \U$18749 ( \18881 , \18549 , \18709 );
xor \U$18750 ( \18882 , \18880 , \18881 );
and \U$18751 ( \18883 , \18710 , \18711 );
and \U$18752 ( \18884 , \18712 , \18715 );
or \U$18753 ( \18885 , \18883 , \18884 );
xor \U$18754 ( \18886 , \18882 , \18885 );
buf \U$18755 ( \18887 , \18886 );
buf \U$18756 ( \18888 , \18887 );
and \U$18757 ( \18889 , \18726 , \18737 );
and \U$18758 ( \18890 , \18737 , \18878 );
and \U$18759 ( \18891 , \18726 , \18878 );
or \U$18760 ( \18892 , \18889 , \18890 , \18891 );
and \U$18761 ( \18893 , \18742 , \18746 );
and \U$18762 ( \18894 , \18746 , \18877 );
and \U$18763 ( \18895 , \18742 , \18877 );
or \U$18764 ( \18896 , \18893 , \18894 , \18895 );
and \U$18765 ( \18897 , \18751 , \18755 );
and \U$18766 ( \18898 , \18755 , \18760 );
and \U$18767 ( \18899 , \18751 , \18760 );
or \U$18768 ( \18900 , \18897 , \18898 , \18899 );
and \U$18769 ( \18901 , \18765 , \18808 );
and \U$18770 ( \18902 , \18808 , \18845 );
and \U$18771 ( \18903 , \18765 , \18845 );
or \U$18772 ( \18904 , \18901 , \18902 , \18903 );
xor \U$18773 ( \18905 , \18900 , \18904 );
and \U$18774 ( \18906 , \18861 , \18875 );
xor \U$18775 ( \18907 , \18905 , \18906 );
xor \U$18776 ( \18908 , \18896 , \18907 );
and \U$18777 ( \18909 , \18730 , \18734 );
and \U$18778 ( \18910 , \18734 , \18736 );
and \U$18779 ( \18911 , \18730 , \18736 );
or \U$18780 ( \18912 , \18909 , \18910 , \18911 );
and \U$18781 ( \18913 , \18761 , \18846 );
and \U$18782 ( \18914 , \18846 , \18876 );
and \U$18783 ( \18915 , \18761 , \18876 );
or \U$18784 ( \18916 , \18913 , \18914 , \18915 );
xor \U$18785 ( \18917 , \18912 , \18916 );
and \U$18786 ( \18918 , \18851 , \18855 );
and \U$18787 ( \18919 , \18855 , \18860 );
and \U$18788 ( \18920 , \18851 , \18860 );
or \U$18789 ( \18921 , \18918 , \18919 , \18920 );
and \U$18790 ( \18922 , \18865 , \18869 );
and \U$18791 ( \18923 , \18869 , \18874 );
and \U$18792 ( \18924 , \18865 , \18874 );
or \U$18793 ( \18925 , \18922 , \18923 , \18924 );
xor \U$18794 ( \18926 , \18921 , \18925 );
and \U$18795 ( \18927 , \18823 , \18837 );
and \U$18796 ( \18928 , \18837 , \18844 );
and \U$18797 ( \18929 , \18823 , \18844 );
or \U$18798 ( \18930 , \18927 , \18928 , \18929 );
xor \U$18799 ( \18931 , \18926 , \18930 );
and \U$18800 ( \18932 , \18778 , \18792 );
and \U$18801 ( \18933 , \18792 , \18807 );
and \U$18802 ( \18934 , \18778 , \18807 );
or \U$18803 ( \18935 , \18932 , \18933 , \18934 );
and \U$18804 ( \18936 , \7231 , \5485 );
and \U$18805 ( \18937 , \7556 , \5275 );
nor \U$18806 ( \18938 , \18936 , \18937 );
xnor \U$18807 ( \18939 , \18938 , \5169 );
and \U$18808 ( \18940 , \6790 , \5996 );
and \U$18809 ( \18941 , \6945 , \5695 );
nor \U$18810 ( \18942 , \18940 , \18941 );
xnor \U$18811 ( \18943 , \18942 , \5687 );
xor \U$18812 ( \18944 , \18939 , \18943 );
and \U$18813 ( \18945 , \6281 , \6401 );
and \U$18814 ( \18946 , \6514 , \6143 );
nor \U$18815 ( \18947 , \18945 , \18946 );
xnor \U$18816 ( \18948 , \18947 , \6148 );
xor \U$18817 ( \18949 , \18944 , \18948 );
not \U$18818 ( \18950 , \2839 );
and \U$18819 ( \18951 , \10206 , \3357 );
and \U$18820 ( \18952 , \10584 , \3255 );
nor \U$18821 ( \18953 , \18951 , \18952 );
xnor \U$18822 ( \18954 , \18953 , \3156 );
xor \U$18823 ( \18955 , \18950 , \18954 );
and \U$18824 ( \18956 , \9465 , \3813 );
and \U$18825 ( \18957 , \9897 , \3557 );
nor \U$18826 ( \18958 , \18956 , \18957 );
xnor \U$18827 ( \18959 , \18958 , \3562 );
xor \U$18828 ( \18960 , \18955 , \18959 );
xor \U$18829 ( \18961 , \18949 , \18960 );
and \U$18830 ( \18962 , \8835 , \4132 );
and \U$18831 ( \18963 , \9169 , \4012 );
nor \U$18832 ( \18964 , \18962 , \18963 );
xnor \U$18833 ( \18965 , \18964 , \3925 );
and \U$18834 ( \18966 , \8349 , \4581 );
and \U$18835 ( \18967 , \8652 , \4424 );
nor \U$18836 ( \18968 , \18966 , \18967 );
xnor \U$18837 ( \18969 , \18968 , \4377 );
xor \U$18838 ( \18970 , \18965 , \18969 );
and \U$18839 ( \18971 , \7700 , \5011 );
and \U$18840 ( \18972 , \8057 , \4878 );
nor \U$18841 ( \18973 , \18971 , \18972 );
xnor \U$18842 ( \18974 , \18973 , \4762 );
xor \U$18843 ( \18975 , \18970 , \18974 );
xor \U$18844 ( \18976 , \18961 , \18975 );
xor \U$18845 ( \18977 , \18935 , \18976 );
and \U$18846 ( \18978 , \4364 , \8540 );
and \U$18847 ( \18979 , \4654 , \8292 );
nor \U$18848 ( \18980 , \18978 , \18979 );
xnor \U$18849 ( \18981 , \18980 , \8297 );
and \U$18850 ( \18982 , \3912 , \9333 );
and \U$18851 ( \18983 , \4160 , \9006 );
nor \U$18852 ( \18984 , \18982 , \18983 );
xnor \U$18853 ( \18985 , \18984 , \8848 );
xor \U$18854 ( \18986 , \18981 , \18985 );
and \U$18855 ( \18987 , \3646 , \9765 );
and \U$18856 ( \18988 , \3736 , \9644 );
nor \U$18857 ( \18989 , \18987 , \18988 );
xnor \U$18858 ( \18990 , \18989 , \9478 );
xor \U$18859 ( \18991 , \18986 , \18990 );
and \U$18860 ( \18992 , \5674 , \7055 );
and \U$18861 ( \18993 , \6030 , \6675 );
nor \U$18862 ( \18994 , \18992 , \18993 );
xnor \U$18863 ( \18995 , \18994 , \6680 );
and \U$18864 ( \18996 , \5156 , \7489 );
and \U$18865 ( \18997 , \5469 , \7137 );
nor \U$18866 ( \18998 , \18996 , \18997 );
xnor \U$18867 ( \18999 , \18998 , \7142 );
xor \U$18868 ( \19000 , \18995 , \18999 );
and \U$18869 ( \19001 , \4749 , \8019 );
and \U$18870 ( \19002 , \4922 , \7830 );
nor \U$18871 ( \19003 , \19001 , \19002 );
xnor \U$18872 ( \19004 , \19003 , \7713 );
xor \U$18873 ( \19005 , \19000 , \19004 );
xor \U$18874 ( \19006 , \18991 , \19005 );
and \U$18875 ( \19007 , \3143 , \10408 );
and \U$18876 ( \19008 , \3395 , \10116 );
nor \U$18877 ( \19009 , \19007 , \19008 );
xnor \U$18878 ( \19010 , \19009 , \10121 );
and \U$18879 ( \19011 , \3037 , \10118 );
xor \U$18880 ( \19012 , \19010 , \19011 );
xor \U$18881 ( \19013 , \19006 , \19012 );
xor \U$18882 ( \19014 , \18977 , \19013 );
xor \U$18883 ( \19015 , \18931 , \19014 );
and \U$18884 ( \19016 , \18768 , \18772 );
and \U$18885 ( \19017 , \18772 , \18777 );
and \U$18886 ( \19018 , \18768 , \18777 );
or \U$18887 ( \19019 , \19016 , \19017 , \19018 );
and \U$18888 ( \19020 , \18782 , \18786 );
and \U$18889 ( \19021 , \18786 , \18791 );
and \U$18890 ( \19022 , \18782 , \18791 );
or \U$18891 ( \19023 , \19020 , \19021 , \19022 );
xor \U$18892 ( \19024 , \19019 , \19023 );
and \U$18893 ( \19025 , \18797 , \18801 );
and \U$18894 ( \19026 , \18801 , \18806 );
and \U$18895 ( \19027 , \18797 , \18806 );
or \U$18896 ( \19028 , \19025 , \19026 , \19027 );
xor \U$18897 ( \19029 , \19024 , \19028 );
and \U$18898 ( \19030 , \18813 , \18817 );
and \U$18899 ( \19031 , \18817 , \18822 );
and \U$18900 ( \19032 , \18813 , \18822 );
or \U$18901 ( \19033 , \19030 , \19031 , \19032 );
and \U$18902 ( \19034 , \18827 , \18831 );
and \U$18903 ( \19035 , \18831 , \18836 );
and \U$18904 ( \19036 , \18827 , \18836 );
or \U$18905 ( \19037 , \19034 , \19035 , \19036 );
xor \U$18906 ( \19038 , \19033 , \19037 );
or \U$18907 ( \19039 , \18842 , \18843 );
xor \U$18908 ( \19040 , \19038 , \19039 );
xor \U$18909 ( \19041 , \19029 , \19040 );
xor \U$18910 ( \19042 , \19015 , \19041 );
xor \U$18911 ( \19043 , \18917 , \19042 );
xor \U$18912 ( \19044 , \18908 , \19043 );
xor \U$18913 ( \19045 , \18892 , \19044 );
and \U$18914 ( \19046 , \18722 , \18879 );
xor \U$18915 ( \19047 , \19045 , \19046 );
and \U$18916 ( \19048 , \18880 , \18881 );
and \U$18917 ( \19049 , \18882 , \18885 );
or \U$18918 ( \19050 , \19048 , \19049 );
xor \U$18919 ( \19051 , \19047 , \19050 );
buf \U$18920 ( \19052 , \19051 );
buf \U$18921 ( \19053 , \19052 );
and \U$18922 ( \19054 , \18896 , \18907 );
and \U$18923 ( \19055 , \18907 , \19043 );
and \U$18924 ( \19056 , \18896 , \19043 );
or \U$18925 ( \19057 , \19054 , \19055 , \19056 );
and \U$18926 ( \19058 , \18912 , \18916 );
and \U$18927 ( \19059 , \18916 , \19042 );
and \U$18928 ( \19060 , \18912 , \19042 );
or \U$18929 ( \19061 , \19058 , \19059 , \19060 );
and \U$18930 ( \19062 , \18921 , \18925 );
and \U$18931 ( \19063 , \18925 , \18930 );
and \U$18932 ( \19064 , \18921 , \18930 );
or \U$18933 ( \19065 , \19062 , \19063 , \19064 );
and \U$18934 ( \19066 , \18935 , \18976 );
and \U$18935 ( \19067 , \18976 , \19013 );
and \U$18936 ( \19068 , \18935 , \19013 );
or \U$18937 ( \19069 , \19066 , \19067 , \19068 );
xor \U$18938 ( \19070 , \19065 , \19069 );
and \U$18939 ( \19071 , \19029 , \19040 );
xor \U$18940 ( \19072 , \19070 , \19071 );
xor \U$18941 ( \19073 , \19061 , \19072 );
and \U$18942 ( \19074 , \18900 , \18904 );
and \U$18943 ( \19075 , \18904 , \18906 );
and \U$18944 ( \19076 , \18900 , \18906 );
or \U$18945 ( \19077 , \19074 , \19075 , \19076 );
and \U$18946 ( \19078 , \18931 , \19014 );
and \U$18947 ( \19079 , \19014 , \19041 );
and \U$18948 ( \19080 , \18931 , \19041 );
or \U$18949 ( \19081 , \19078 , \19079 , \19080 );
xor \U$18950 ( \19082 , \19077 , \19081 );
and \U$18951 ( \19083 , \19019 , \19023 );
and \U$18952 ( \19084 , \19023 , \19028 );
and \U$18953 ( \19085 , \19019 , \19028 );
or \U$18954 ( \19086 , \19083 , \19084 , \19085 );
and \U$18955 ( \19087 , \19033 , \19037 );
and \U$18956 ( \19088 , \19037 , \19039 );
and \U$18957 ( \19089 , \19033 , \19039 );
or \U$18958 ( \19090 , \19087 , \19088 , \19089 );
xor \U$18959 ( \19091 , \19086 , \19090 );
and \U$18960 ( \19092 , \18991 , \19005 );
and \U$18961 ( \19093 , \19005 , \19012 );
and \U$18962 ( \19094 , \18991 , \19012 );
or \U$18963 ( \19095 , \19092 , \19093 , \19094 );
xor \U$18964 ( \19096 , \19091 , \19095 );
and \U$18965 ( \19097 , \18949 , \18960 );
and \U$18966 ( \19098 , \18960 , \18975 );
and \U$18967 ( \19099 , \18949 , \18975 );
or \U$18968 ( \19100 , \19097 , \19098 , \19099 );
and \U$18969 ( \19101 , \8652 , \4581 );
and \U$18970 ( \19102 , \8835 , \4424 );
nor \U$18971 ( \19103 , \19101 , \19102 );
xnor \U$18972 ( \19104 , \19103 , \4377 );
and \U$18973 ( \19105 , \8057 , \5011 );
and \U$18974 ( \19106 , \8349 , \4878 );
nor \U$18975 ( \19107 , \19105 , \19106 );
xnor \U$18976 ( \19108 , \19107 , \4762 );
xor \U$18977 ( \19109 , \19104 , \19108 );
and \U$18978 ( \19110 , \7556 , \5485 );
and \U$18979 ( \19111 , \7700 , \5275 );
nor \U$18980 ( \19112 , \19110 , \19111 );
xnor \U$18981 ( \19113 , \19112 , \5169 );
xor \U$18982 ( \19114 , \19109 , \19113 );
and \U$18983 ( \19115 , \10584 , \3357 );
not \U$18984 ( \19116 , \19115 );
xnor \U$18985 ( \19117 , \19116 , \3156 );
and \U$18986 ( \19118 , \9897 , \3813 );
and \U$18987 ( \19119 , \10206 , \3557 );
nor \U$18988 ( \19120 , \19118 , \19119 );
xnor \U$18989 ( \19121 , \19120 , \3562 );
xor \U$18990 ( \19122 , \19117 , \19121 );
and \U$18991 ( \19123 , \9169 , \4132 );
and \U$18992 ( \19124 , \9465 , \4012 );
nor \U$18993 ( \19125 , \19123 , \19124 );
xnor \U$18994 ( \19126 , \19125 , \3925 );
xor \U$18995 ( \19127 , \19122 , \19126 );
xor \U$18996 ( \19128 , \19114 , \19127 );
and \U$18997 ( \19129 , \6945 , \5996 );
and \U$18998 ( \19130 , \7231 , \5695 );
nor \U$18999 ( \19131 , \19129 , \19130 );
xnor \U$19000 ( \19132 , \19131 , \5687 );
and \U$19001 ( \19133 , \6514 , \6401 );
and \U$19002 ( \19134 , \6790 , \6143 );
nor \U$19003 ( \19135 , \19133 , \19134 );
xnor \U$19004 ( \19136 , \19135 , \6148 );
xor \U$19005 ( \19137 , \19132 , \19136 );
and \U$19006 ( \19138 , \6030 , \7055 );
and \U$19007 ( \19139 , \6281 , \6675 );
nor \U$19008 ( \19140 , \19138 , \19139 );
xnor \U$19009 ( \19141 , \19140 , \6680 );
xor \U$19010 ( \19142 , \19137 , \19141 );
xor \U$19011 ( \19143 , \19128 , \19142 );
xor \U$19012 ( \19144 , \19100 , \19143 );
and \U$19013 ( \19145 , \4160 , \9333 );
and \U$19014 ( \19146 , \4364 , \9006 );
nor \U$19015 ( \19147 , \19145 , \19146 );
xnor \U$19016 ( \19148 , \19147 , \8848 );
and \U$19017 ( \19149 , \3736 , \9765 );
and \U$19018 ( \19150 , \3912 , \9644 );
nor \U$19019 ( \19151 , \19149 , \19150 );
xnor \U$19020 ( \19152 , \19151 , \9478 );
xor \U$19021 ( \19153 , \19148 , \19152 );
and \U$19022 ( \19154 , \3395 , \10408 );
and \U$19023 ( \19155 , \3646 , \10116 );
nor \U$19024 ( \19156 , \19154 , \19155 );
xnor \U$19025 ( \19157 , \19156 , \10121 );
xor \U$19026 ( \19158 , \19153 , \19157 );
and \U$19027 ( \19159 , \5469 , \7489 );
and \U$19028 ( \19160 , \5674 , \7137 );
nor \U$19029 ( \19161 , \19159 , \19160 );
xnor \U$19030 ( \19162 , \19161 , \7142 );
and \U$19031 ( \19163 , \4922 , \8019 );
and \U$19032 ( \19164 , \5156 , \7830 );
nor \U$19033 ( \19165 , \19163 , \19164 );
xnor \U$19034 ( \19166 , \19165 , \7713 );
xor \U$19035 ( \19167 , \19162 , \19166 );
and \U$19036 ( \19168 , \4654 , \8540 );
and \U$19037 ( \19169 , \4749 , \8292 );
nor \U$19038 ( \19170 , \19168 , \19169 );
xnor \U$19039 ( \19171 , \19170 , \8297 );
xor \U$19040 ( \19172 , \19167 , \19171 );
xor \U$19041 ( \19173 , \19158 , \19172 );
and \U$19042 ( \19174 , \3143 , \10118 );
not \U$19043 ( \19175 , \19174 );
xor \U$19044 ( \19176 , \19173 , \19175 );
xor \U$19045 ( \19177 , \19144 , \19176 );
xor \U$19046 ( \19178 , \19096 , \19177 );
and \U$19047 ( \19179 , \18939 , \18943 );
and \U$19048 ( \19180 , \18943 , \18948 );
and \U$19049 ( \19181 , \18939 , \18948 );
or \U$19050 ( \19182 , \19179 , \19180 , \19181 );
and \U$19051 ( \19183 , \18950 , \18954 );
and \U$19052 ( \19184 , \18954 , \18959 );
and \U$19053 ( \19185 , \18950 , \18959 );
or \U$19054 ( \19186 , \19183 , \19184 , \19185 );
xor \U$19055 ( \19187 , \19182 , \19186 );
and \U$19056 ( \19188 , \18965 , \18969 );
and \U$19057 ( \19189 , \18969 , \18974 );
and \U$19058 ( \19190 , \18965 , \18974 );
or \U$19059 ( \19191 , \19188 , \19189 , \19190 );
xor \U$19060 ( \19192 , \19187 , \19191 );
and \U$19061 ( \19193 , \18981 , \18985 );
and \U$19062 ( \19194 , \18985 , \18990 );
and \U$19063 ( \19195 , \18981 , \18990 );
or \U$19064 ( \19196 , \19193 , \19194 , \19195 );
and \U$19065 ( \19197 , \18995 , \18999 );
and \U$19066 ( \19198 , \18999 , \19004 );
and \U$19067 ( \19199 , \18995 , \19004 );
or \U$19068 ( \19200 , \19197 , \19198 , \19199 );
xor \U$19069 ( \19201 , \19196 , \19200 );
and \U$19070 ( \19202 , \19010 , \19011 );
xor \U$19071 ( \19203 , \19201 , \19202 );
xor \U$19072 ( \19204 , \19192 , \19203 );
xor \U$19073 ( \19205 , \19178 , \19204 );
xor \U$19074 ( \19206 , \19082 , \19205 );
xor \U$19075 ( \19207 , \19073 , \19206 );
xor \U$19076 ( \19208 , \19057 , \19207 );
and \U$19077 ( \19209 , \18892 , \19044 );
xor \U$19078 ( \19210 , \19208 , \19209 );
and \U$19079 ( \19211 , \19045 , \19046 );
and \U$19080 ( \19212 , \19047 , \19050 );
or \U$19081 ( \19213 , \19211 , \19212 );
xor \U$19082 ( \19214 , \19210 , \19213 );
buf \U$19083 ( \19215 , \19214 );
buf \U$19084 ( \19216 , \19215 );
and \U$19085 ( \19217 , \19061 , \19072 );
and \U$19086 ( \19218 , \19072 , \19206 );
and \U$19087 ( \19219 , \19061 , \19206 );
or \U$19088 ( \19220 , \19217 , \19218 , \19219 );
and \U$19089 ( \19221 , \19077 , \19081 );
and \U$19090 ( \19222 , \19081 , \19205 );
and \U$19091 ( \19223 , \19077 , \19205 );
or \U$19092 ( \19224 , \19221 , \19222 , \19223 );
and \U$19093 ( \19225 , \19086 , \19090 );
and \U$19094 ( \19226 , \19090 , \19095 );
and \U$19095 ( \19227 , \19086 , \19095 );
or \U$19096 ( \19228 , \19225 , \19226 , \19227 );
and \U$19097 ( \19229 , \19100 , \19143 );
and \U$19098 ( \19230 , \19143 , \19176 );
and \U$19099 ( \19231 , \19100 , \19176 );
or \U$19100 ( \19232 , \19229 , \19230 , \19231 );
xor \U$19101 ( \19233 , \19228 , \19232 );
and \U$19102 ( \19234 , \19192 , \19203 );
xor \U$19103 ( \19235 , \19233 , \19234 );
xor \U$19104 ( \19236 , \19224 , \19235 );
and \U$19105 ( \19237 , \19065 , \19069 );
and \U$19106 ( \19238 , \19069 , \19071 );
and \U$19107 ( \19239 , \19065 , \19071 );
or \U$19108 ( \19240 , \19237 , \19238 , \19239 );
and \U$19109 ( \19241 , \19096 , \19177 );
and \U$19110 ( \19242 , \19177 , \19204 );
and \U$19111 ( \19243 , \19096 , \19204 );
or \U$19112 ( \19244 , \19241 , \19242 , \19243 );
xor \U$19113 ( \19245 , \19240 , \19244 );
and \U$19114 ( \19246 , \19182 , \19186 );
and \U$19115 ( \19247 , \19186 , \19191 );
and \U$19116 ( \19248 , \19182 , \19191 );
or \U$19117 ( \19249 , \19246 , \19247 , \19248 );
and \U$19118 ( \19250 , \19196 , \19200 );
and \U$19119 ( \19251 , \19200 , \19202 );
and \U$19120 ( \19252 , \19196 , \19202 );
or \U$19121 ( \19253 , \19250 , \19251 , \19252 );
xor \U$19122 ( \19254 , \19249 , \19253 );
and \U$19123 ( \19255 , \19158 , \19172 );
and \U$19124 ( \19256 , \19172 , \19175 );
and \U$19125 ( \19257 , \19158 , \19175 );
or \U$19126 ( \19258 , \19255 , \19256 , \19257 );
xor \U$19127 ( \19259 , \19254 , \19258 );
and \U$19128 ( \19260 , \19114 , \19127 );
and \U$19129 ( \19261 , \19127 , \19142 );
and \U$19130 ( \19262 , \19114 , \19142 );
or \U$19131 ( \19263 , \19260 , \19261 , \19262 );
and \U$19132 ( \19264 , \8835 , \4581 );
and \U$19133 ( \19265 , \9169 , \4424 );
nor \U$19134 ( \19266 , \19264 , \19265 );
xnor \U$19135 ( \19267 , \19266 , \4377 );
and \U$19136 ( \19268 , \8349 , \5011 );
and \U$19137 ( \19269 , \8652 , \4878 );
nor \U$19138 ( \19270 , \19268 , \19269 );
xnor \U$19139 ( \19271 , \19270 , \4762 );
xor \U$19140 ( \19272 , \19267 , \19271 );
and \U$19141 ( \19273 , \7700 , \5485 );
and \U$19142 ( \19274 , \8057 , \5275 );
nor \U$19143 ( \19275 , \19273 , \19274 );
xnor \U$19144 ( \19276 , \19275 , \5169 );
xor \U$19145 ( \19277 , \19272 , \19276 );
not \U$19146 ( \19278 , \3156 );
and \U$19147 ( \19279 , \10206 , \3813 );
and \U$19148 ( \19280 , \10584 , \3557 );
nor \U$19149 ( \19281 , \19279 , \19280 );
xnor \U$19150 ( \19282 , \19281 , \3562 );
xor \U$19151 ( \19283 , \19278 , \19282 );
and \U$19152 ( \19284 , \9465 , \4132 );
and \U$19153 ( \19285 , \9897 , \4012 );
nor \U$19154 ( \19286 , \19284 , \19285 );
xnor \U$19155 ( \19287 , \19286 , \3925 );
xor \U$19156 ( \19288 , \19283 , \19287 );
xor \U$19157 ( \19289 , \19277 , \19288 );
and \U$19158 ( \19290 , \7231 , \5996 );
and \U$19159 ( \19291 , \7556 , \5695 );
nor \U$19160 ( \19292 , \19290 , \19291 );
xnor \U$19161 ( \19293 , \19292 , \5687 );
and \U$19162 ( \19294 , \6790 , \6401 );
and \U$19163 ( \19295 , \6945 , \6143 );
nor \U$19164 ( \19296 , \19294 , \19295 );
xnor \U$19165 ( \19297 , \19296 , \6148 );
xor \U$19166 ( \19298 , \19293 , \19297 );
and \U$19167 ( \19299 , \6281 , \7055 );
and \U$19168 ( \19300 , \6514 , \6675 );
nor \U$19169 ( \19301 , \19299 , \19300 );
xnor \U$19170 ( \19302 , \19301 , \6680 );
xor \U$19171 ( \19303 , \19298 , \19302 );
xor \U$19172 ( \19304 , \19289 , \19303 );
xor \U$19173 ( \19305 , \19263 , \19304 );
and \U$19174 ( \19306 , \3395 , \10118 );
and \U$19175 ( \19307 , \4364 , \9333 );
and \U$19176 ( \19308 , \4654 , \9006 );
nor \U$19177 ( \19309 , \19307 , \19308 );
xnor \U$19178 ( \19310 , \19309 , \8848 );
and \U$19179 ( \19311 , \3912 , \9765 );
and \U$19180 ( \19312 , \4160 , \9644 );
nor \U$19181 ( \19313 , \19311 , \19312 );
xnor \U$19182 ( \19314 , \19313 , \9478 );
xor \U$19183 ( \19315 , \19310 , \19314 );
and \U$19184 ( \19316 , \3646 , \10408 );
and \U$19185 ( \19317 , \3736 , \10116 );
nor \U$19186 ( \19318 , \19316 , \19317 );
xnor \U$19187 ( \19319 , \19318 , \10121 );
xor \U$19188 ( \19320 , \19315 , \19319 );
xor \U$19189 ( \19321 , \19306 , \19320 );
and \U$19190 ( \19322 , \5674 , \7489 );
and \U$19191 ( \19323 , \6030 , \7137 );
nor \U$19192 ( \19324 , \19322 , \19323 );
xnor \U$19193 ( \19325 , \19324 , \7142 );
and \U$19194 ( \19326 , \5156 , \8019 );
and \U$19195 ( \19327 , \5469 , \7830 );
nor \U$19196 ( \19328 , \19326 , \19327 );
xnor \U$19197 ( \19329 , \19328 , \7713 );
xor \U$19198 ( \19330 , \19325 , \19329 );
and \U$19199 ( \19331 , \4749 , \8540 );
and \U$19200 ( \19332 , \4922 , \8292 );
nor \U$19201 ( \19333 , \19331 , \19332 );
xnor \U$19202 ( \19334 , \19333 , \8297 );
xor \U$19203 ( \19335 , \19330 , \19334 );
xor \U$19204 ( \19336 , \19321 , \19335 );
xor \U$19205 ( \19337 , \19305 , \19336 );
xor \U$19206 ( \19338 , \19259 , \19337 );
and \U$19207 ( \19339 , \19104 , \19108 );
and \U$19208 ( \19340 , \19108 , \19113 );
and \U$19209 ( \19341 , \19104 , \19113 );
or \U$19210 ( \19342 , \19339 , \19340 , \19341 );
and \U$19211 ( \19343 , \19117 , \19121 );
and \U$19212 ( \19344 , \19121 , \19126 );
and \U$19213 ( \19345 , \19117 , \19126 );
or \U$19214 ( \19346 , \19343 , \19344 , \19345 );
xor \U$19215 ( \19347 , \19342 , \19346 );
and \U$19216 ( \19348 , \19132 , \19136 );
and \U$19217 ( \19349 , \19136 , \19141 );
and \U$19218 ( \19350 , \19132 , \19141 );
or \U$19219 ( \19351 , \19348 , \19349 , \19350 );
xor \U$19220 ( \19352 , \19347 , \19351 );
and \U$19221 ( \19353 , \19148 , \19152 );
and \U$19222 ( \19354 , \19152 , \19157 );
and \U$19223 ( \19355 , \19148 , \19157 );
or \U$19224 ( \19356 , \19353 , \19354 , \19355 );
and \U$19225 ( \19357 , \19162 , \19166 );
and \U$19226 ( \19358 , \19166 , \19171 );
and \U$19227 ( \19359 , \19162 , \19171 );
or \U$19228 ( \19360 , \19357 , \19358 , \19359 );
xor \U$19229 ( \19361 , \19356 , \19360 );
buf \U$19230 ( \19362 , \19174 );
xor \U$19231 ( \19363 , \19361 , \19362 );
xor \U$19232 ( \19364 , \19352 , \19363 );
xor \U$19233 ( \19365 , \19338 , \19364 );
xor \U$19234 ( \19366 , \19245 , \19365 );
xor \U$19235 ( \19367 , \19236 , \19366 );
xor \U$19236 ( \19368 , \19220 , \19367 );
and \U$19237 ( \19369 , \19057 , \19207 );
xor \U$19238 ( \19370 , \19368 , \19369 );
and \U$19239 ( \19371 , \19208 , \19209 );
and \U$19240 ( \19372 , \19210 , \19213 );
or \U$19241 ( \19373 , \19371 , \19372 );
xor \U$19242 ( \19374 , \19370 , \19373 );
buf \U$19243 ( \19375 , \19374 );
buf \U$19244 ( \19376 , \19375 );
and \U$19245 ( \19377 , \19224 , \19235 );
and \U$19246 ( \19378 , \19235 , \19366 );
and \U$19247 ( \19379 , \19224 , \19366 );
or \U$19248 ( \19380 , \19377 , \19378 , \19379 );
and \U$19249 ( \19381 , \19240 , \19244 );
and \U$19250 ( \19382 , \19244 , \19365 );
and \U$19251 ( \19383 , \19240 , \19365 );
or \U$19252 ( \19384 , \19381 , \19382 , \19383 );
and \U$19253 ( \19385 , \19249 , \19253 );
and \U$19254 ( \19386 , \19253 , \19258 );
and \U$19255 ( \19387 , \19249 , \19258 );
or \U$19256 ( \19388 , \19385 , \19386 , \19387 );
and \U$19257 ( \19389 , \19263 , \19304 );
and \U$19258 ( \19390 , \19304 , \19336 );
and \U$19259 ( \19391 , \19263 , \19336 );
or \U$19260 ( \19392 , \19389 , \19390 , \19391 );
xor \U$19261 ( \19393 , \19388 , \19392 );
and \U$19262 ( \19394 , \19352 , \19363 );
xor \U$19263 ( \19395 , \19393 , \19394 );
xor \U$19264 ( \19396 , \19384 , \19395 );
and \U$19265 ( \19397 , \19228 , \19232 );
and \U$19266 ( \19398 , \19232 , \19234 );
and \U$19267 ( \19399 , \19228 , \19234 );
or \U$19268 ( \19400 , \19397 , \19398 , \19399 );
and \U$19269 ( \19401 , \19259 , \19337 );
and \U$19270 ( \19402 , \19337 , \19364 );
and \U$19271 ( \19403 , \19259 , \19364 );
or \U$19272 ( \19404 , \19401 , \19402 , \19403 );
xor \U$19273 ( \19405 , \19400 , \19404 );
and \U$19274 ( \19406 , \19342 , \19346 );
and \U$19275 ( \19407 , \19346 , \19351 );
and \U$19276 ( \19408 , \19342 , \19351 );
or \U$19277 ( \19409 , \19406 , \19407 , \19408 );
and \U$19278 ( \19410 , \19356 , \19360 );
and \U$19279 ( \19411 , \19360 , \19362 );
and \U$19280 ( \19412 , \19356 , \19362 );
or \U$19281 ( \19413 , \19410 , \19411 , \19412 );
xor \U$19282 ( \19414 , \19409 , \19413 );
and \U$19283 ( \19415 , \19306 , \19320 );
and \U$19284 ( \19416 , \19320 , \19335 );
and \U$19285 ( \19417 , \19306 , \19335 );
or \U$19286 ( \19418 , \19415 , \19416 , \19417 );
xor \U$19287 ( \19419 , \19414 , \19418 );
and \U$19288 ( \19420 , \19277 , \19288 );
and \U$19289 ( \19421 , \19288 , \19303 );
and \U$19290 ( \19422 , \19277 , \19303 );
or \U$19291 ( \19423 , \19420 , \19421 , \19422 );
and \U$19292 ( \19424 , \10584 , \3813 );
not \U$19293 ( \19425 , \19424 );
xnor \U$19294 ( \19426 , \19425 , \3562 );
and \U$19295 ( \19427 , \9897 , \4132 );
and \U$19296 ( \19428 , \10206 , \4012 );
nor \U$19297 ( \19429 , \19427 , \19428 );
xnor \U$19298 ( \19430 , \19429 , \3925 );
xor \U$19299 ( \19431 , \19426 , \19430 );
and \U$19300 ( \19432 , \9169 , \4581 );
and \U$19301 ( \19433 , \9465 , \4424 );
nor \U$19302 ( \19434 , \19432 , \19433 );
xnor \U$19303 ( \19435 , \19434 , \4377 );
xor \U$19304 ( \19436 , \19431 , \19435 );
xor \U$19305 ( \19437 , \19423 , \19436 );
and \U$19306 ( \19438 , \8652 , \5011 );
and \U$19307 ( \19439 , \8835 , \4878 );
nor \U$19308 ( \19440 , \19438 , \19439 );
xnor \U$19309 ( \19441 , \19440 , \4762 );
and \U$19310 ( \19442 , \8057 , \5485 );
and \U$19311 ( \19443 , \8349 , \5275 );
nor \U$19312 ( \19444 , \19442 , \19443 );
xnor \U$19313 ( \19445 , \19444 , \5169 );
xor \U$19314 ( \19446 , \19441 , \19445 );
and \U$19315 ( \19447 , \7556 , \5996 );
and \U$19316 ( \19448 , \7700 , \5695 );
nor \U$19317 ( \19449 , \19447 , \19448 );
xnor \U$19318 ( \19450 , \19449 , \5687 );
xor \U$19319 ( \19451 , \19446 , \19450 );
xor \U$19320 ( \19452 , \19437 , \19451 );
xor \U$19321 ( \19453 , \19419 , \19452 );
and \U$19322 ( \19454 , \19267 , \19271 );
and \U$19323 ( \19455 , \19271 , \19276 );
and \U$19324 ( \19456 , \19267 , \19276 );
or \U$19325 ( \19457 , \19454 , \19455 , \19456 );
and \U$19326 ( \19458 , \19278 , \19282 );
and \U$19327 ( \19459 , \19282 , \19287 );
and \U$19328 ( \19460 , \19278 , \19287 );
or \U$19329 ( \19461 , \19458 , \19459 , \19460 );
xor \U$19330 ( \19462 , \19457 , \19461 );
and \U$19331 ( \19463 , \19293 , \19297 );
and \U$19332 ( \19464 , \19297 , \19302 );
and \U$19333 ( \19465 , \19293 , \19302 );
or \U$19334 ( \19466 , \19463 , \19464 , \19465 );
xor \U$19335 ( \19467 , \19462 , \19466 );
and \U$19336 ( \19468 , \5469 , \8019 );
and \U$19337 ( \19469 , \5674 , \7830 );
nor \U$19338 ( \19470 , \19468 , \19469 );
xnor \U$19339 ( \19471 , \19470 , \7713 );
and \U$19340 ( \19472 , \4922 , \8540 );
and \U$19341 ( \19473 , \5156 , \8292 );
nor \U$19342 ( \19474 , \19472 , \19473 );
xnor \U$19343 ( \19475 , \19474 , \8297 );
xor \U$19344 ( \19476 , \19471 , \19475 );
and \U$19345 ( \19477 , \4654 , \9333 );
and \U$19346 ( \19478 , \4749 , \9006 );
nor \U$19347 ( \19479 , \19477 , \19478 );
xnor \U$19348 ( \19480 , \19479 , \8848 );
xor \U$19349 ( \19481 , \19476 , \19480 );
and \U$19350 ( \19482 , \4160 , \9765 );
and \U$19351 ( \19483 , \4364 , \9644 );
nor \U$19352 ( \19484 , \19482 , \19483 );
xnor \U$19353 ( \19485 , \19484 , \9478 );
and \U$19354 ( \19486 , \3736 , \10408 );
and \U$19355 ( \19487 , \3912 , \10116 );
nor \U$19356 ( \19488 , \19486 , \19487 );
xnor \U$19357 ( \19489 , \19488 , \10121 );
xor \U$19358 ( \19490 , \19485 , \19489 );
and \U$19359 ( \19491 , \3646 , \10118 );
xor \U$19360 ( \19492 , \19490 , \19491 );
xor \U$19361 ( \19493 , \19481 , \19492 );
and \U$19362 ( \19494 , \6945 , \6401 );
and \U$19363 ( \19495 , \7231 , \6143 );
nor \U$19364 ( \19496 , \19494 , \19495 );
xnor \U$19365 ( \19497 , \19496 , \6148 );
and \U$19366 ( \19498 , \6514 , \7055 );
and \U$19367 ( \19499 , \6790 , \6675 );
nor \U$19368 ( \19500 , \19498 , \19499 );
xnor \U$19369 ( \19501 , \19500 , \6680 );
xor \U$19370 ( \19502 , \19497 , \19501 );
and \U$19371 ( \19503 , \6030 , \7489 );
and \U$19372 ( \19504 , \6281 , \7137 );
nor \U$19373 ( \19505 , \19503 , \19504 );
xnor \U$19374 ( \19506 , \19505 , \7142 );
xor \U$19375 ( \19507 , \19502 , \19506 );
xor \U$19376 ( \19508 , \19493 , \19507 );
xor \U$19377 ( \19509 , \19467 , \19508 );
and \U$19378 ( \19510 , \19310 , \19314 );
and \U$19379 ( \19511 , \19314 , \19319 );
and \U$19380 ( \19512 , \19310 , \19319 );
or \U$19381 ( \19513 , \19510 , \19511 , \19512 );
and \U$19382 ( \19514 , \19325 , \19329 );
and \U$19383 ( \19515 , \19329 , \19334 );
and \U$19384 ( \19516 , \19325 , \19334 );
or \U$19385 ( \19517 , \19514 , \19515 , \19516 );
xnor \U$19386 ( \19518 , \19513 , \19517 );
xor \U$19387 ( \19519 , \19509 , \19518 );
xor \U$19388 ( \19520 , \19453 , \19519 );
xor \U$19389 ( \19521 , \19405 , \19520 );
xor \U$19390 ( \19522 , \19396 , \19521 );
xor \U$19391 ( \19523 , \19380 , \19522 );
and \U$19392 ( \19524 , \19220 , \19367 );
xor \U$19393 ( \19525 , \19523 , \19524 );
and \U$19394 ( \19526 , \19368 , \19369 );
and \U$19395 ( \19527 , \19370 , \19373 );
or \U$19396 ( \19528 , \19526 , \19527 );
xor \U$19397 ( \19529 , \19525 , \19528 );
buf \U$19398 ( \19530 , \19529 );
buf \U$19399 ( \19531 , \19530 );
and \U$19400 ( \19532 , \19384 , \19395 );
and \U$19401 ( \19533 , \19395 , \19521 );
and \U$19402 ( \19534 , \19384 , \19521 );
or \U$19403 ( \19535 , \19532 , \19533 , \19534 );
and \U$19404 ( \19536 , \19400 , \19404 );
and \U$19405 ( \19537 , \19404 , \19520 );
and \U$19406 ( \19538 , \19400 , \19520 );
or \U$19407 ( \19539 , \19536 , \19537 , \19538 );
and \U$19408 ( \19540 , \19409 , \19413 );
and \U$19409 ( \19541 , \19413 , \19418 );
and \U$19410 ( \19542 , \19409 , \19418 );
or \U$19411 ( \19543 , \19540 , \19541 , \19542 );
and \U$19412 ( \19544 , \19423 , \19436 );
and \U$19413 ( \19545 , \19436 , \19451 );
and \U$19414 ( \19546 , \19423 , \19451 );
or \U$19415 ( \19547 , \19544 , \19545 , \19546 );
xor \U$19416 ( \19548 , \19543 , \19547 );
and \U$19417 ( \19549 , \19467 , \19508 );
and \U$19418 ( \19550 , \19508 , \19518 );
and \U$19419 ( \19551 , \19467 , \19518 );
or \U$19420 ( \19552 , \19549 , \19550 , \19551 );
xor \U$19421 ( \19553 , \19548 , \19552 );
xor \U$19422 ( \19554 , \19539 , \19553 );
and \U$19423 ( \19555 , \19388 , \19392 );
and \U$19424 ( \19556 , \19392 , \19394 );
and \U$19425 ( \19557 , \19388 , \19394 );
or \U$19426 ( \19558 , \19555 , \19556 , \19557 );
and \U$19427 ( \19559 , \19419 , \19452 );
and \U$19428 ( \19560 , \19452 , \19519 );
and \U$19429 ( \19561 , \19419 , \19519 );
or \U$19430 ( \19562 , \19559 , \19560 , \19561 );
xor \U$19431 ( \19563 , \19558 , \19562 );
and \U$19432 ( \19564 , \19426 , \19430 );
and \U$19433 ( \19565 , \19430 , \19435 );
and \U$19434 ( \19566 , \19426 , \19435 );
or \U$19435 ( \19567 , \19564 , \19565 , \19566 );
and \U$19436 ( \19568 , \19441 , \19445 );
and \U$19437 ( \19569 , \19445 , \19450 );
and \U$19438 ( \19570 , \19441 , \19450 );
or \U$19439 ( \19571 , \19568 , \19569 , \19570 );
xor \U$19440 ( \19572 , \19567 , \19571 );
and \U$19441 ( \19573 , \19497 , \19501 );
and \U$19442 ( \19574 , \19501 , \19506 );
and \U$19443 ( \19575 , \19497 , \19506 );
or \U$19444 ( \19576 , \19573 , \19574 , \19575 );
xor \U$19445 ( \19577 , \19572 , \19576 );
and \U$19446 ( \19578 , \19457 , \19461 );
and \U$19447 ( \19579 , \19461 , \19466 );
and \U$19448 ( \19580 , \19457 , \19466 );
or \U$19449 ( \19581 , \19578 , \19579 , \19580 );
and \U$19450 ( \19582 , \19481 , \19492 );
and \U$19451 ( \19583 , \19492 , \19507 );
and \U$19452 ( \19584 , \19481 , \19507 );
or \U$19453 ( \19585 , \19582 , \19583 , \19584 );
xor \U$19454 ( \19586 , \19581 , \19585 );
or \U$19455 ( \19587 , \19513 , \19517 );
xor \U$19456 ( \19588 , \19586 , \19587 );
xor \U$19457 ( \19589 , \19577 , \19588 );
not \U$19458 ( \19590 , \3562 );
and \U$19459 ( \19591 , \10206 , \4132 );
and \U$19460 ( \19592 , \10584 , \4012 );
nor \U$19461 ( \19593 , \19591 , \19592 );
xnor \U$19462 ( \19594 , \19593 , \3925 );
xor \U$19463 ( \19595 , \19590 , \19594 );
and \U$19464 ( \19596 , \9465 , \4581 );
and \U$19465 ( \19597 , \9897 , \4424 );
nor \U$19466 ( \19598 , \19596 , \19597 );
xnor \U$19467 ( \19599 , \19598 , \4377 );
xor \U$19468 ( \19600 , \19595 , \19599 );
and \U$19469 ( \19601 , \19471 , \19475 );
and \U$19470 ( \19602 , \19475 , \19480 );
and \U$19471 ( \19603 , \19471 , \19480 );
or \U$19472 ( \19604 , \19601 , \19602 , \19603 );
and \U$19473 ( \19605 , \19485 , \19489 );
and \U$19474 ( \19606 , \19489 , \19491 );
and \U$19475 ( \19607 , \19485 , \19491 );
or \U$19476 ( \19608 , \19605 , \19606 , \19607 );
xor \U$19477 ( \19609 , \19604 , \19608 );
and \U$19478 ( \19610 , \4364 , \9765 );
and \U$19479 ( \19611 , \4654 , \9644 );
nor \U$19480 ( \19612 , \19610 , \19611 );
xnor \U$19481 ( \19613 , \19612 , \9478 );
and \U$19482 ( \19614 , \3912 , \10408 );
and \U$19483 ( \19615 , \4160 , \10116 );
nor \U$19484 ( \19616 , \19614 , \19615 );
xnor \U$19485 ( \19617 , \19616 , \10121 );
xor \U$19486 ( \19618 , \19613 , \19617 );
and \U$19487 ( \19619 , \3736 , \10118 );
xor \U$19488 ( \19620 , \19618 , \19619 );
xor \U$19489 ( \19621 , \19609 , \19620 );
xor \U$19490 ( \19622 , \19600 , \19621 );
and \U$19491 ( \19623 , \8835 , \5011 );
and \U$19492 ( \19624 , \9169 , \4878 );
nor \U$19493 ( \19625 , \19623 , \19624 );
xnor \U$19494 ( \19626 , \19625 , \4762 );
and \U$19495 ( \19627 , \8349 , \5485 );
and \U$19496 ( \19628 , \8652 , \5275 );
nor \U$19497 ( \19629 , \19627 , \19628 );
xnor \U$19498 ( \19630 , \19629 , \5169 );
xor \U$19499 ( \19631 , \19626 , \19630 );
and \U$19500 ( \19632 , \7700 , \5996 );
and \U$19501 ( \19633 , \8057 , \5695 );
nor \U$19502 ( \19634 , \19632 , \19633 );
xnor \U$19503 ( \19635 , \19634 , \5687 );
xor \U$19504 ( \19636 , \19631 , \19635 );
and \U$19505 ( \19637 , \5674 , \8019 );
and \U$19506 ( \19638 , \6030 , \7830 );
nor \U$19507 ( \19639 , \19637 , \19638 );
xnor \U$19508 ( \19640 , \19639 , \7713 );
and \U$19509 ( \19641 , \5156 , \8540 );
and \U$19510 ( \19642 , \5469 , \8292 );
nor \U$19511 ( \19643 , \19641 , \19642 );
xnor \U$19512 ( \19644 , \19643 , \8297 );
xor \U$19513 ( \19645 , \19640 , \19644 );
and \U$19514 ( \19646 , \4749 , \9333 );
and \U$19515 ( \19647 , \4922 , \9006 );
nor \U$19516 ( \19648 , \19646 , \19647 );
xnor \U$19517 ( \19649 , \19648 , \8848 );
xor \U$19518 ( \19650 , \19645 , \19649 );
xor \U$19519 ( \19651 , \19636 , \19650 );
and \U$19520 ( \19652 , \7231 , \6401 );
and \U$19521 ( \19653 , \7556 , \6143 );
nor \U$19522 ( \19654 , \19652 , \19653 );
xnor \U$19523 ( \19655 , \19654 , \6148 );
and \U$19524 ( \19656 , \6790 , \7055 );
and \U$19525 ( \19657 , \6945 , \6675 );
nor \U$19526 ( \19658 , \19656 , \19657 );
xnor \U$19527 ( \19659 , \19658 , \6680 );
xor \U$19528 ( \19660 , \19655 , \19659 );
and \U$19529 ( \19661 , \6281 , \7489 );
and \U$19530 ( \19662 , \6514 , \7137 );
nor \U$19531 ( \19663 , \19661 , \19662 );
xnor \U$19532 ( \19664 , \19663 , \7142 );
xor \U$19533 ( \19665 , \19660 , \19664 );
xor \U$19534 ( \19666 , \19651 , \19665 );
xor \U$19535 ( \19667 , \19622 , \19666 );
xor \U$19536 ( \19668 , \19589 , \19667 );
xor \U$19537 ( \19669 , \19563 , \19668 );
xor \U$19538 ( \19670 , \19554 , \19669 );
xor \U$19539 ( \19671 , \19535 , \19670 );
and \U$19540 ( \19672 , \19380 , \19522 );
xor \U$19541 ( \19673 , \19671 , \19672 );
and \U$19542 ( \19674 , \19523 , \19524 );
and \U$19543 ( \19675 , \19525 , \19528 );
or \U$19544 ( \19676 , \19674 , \19675 );
xor \U$19545 ( \19677 , \19673 , \19676 );
buf \U$19546 ( \19678 , \19677 );
buf \U$19547 ( \19679 , \19678 );
and \U$19548 ( \19680 , \19539 , \19553 );
and \U$19549 ( \19681 , \19553 , \19669 );
and \U$19550 ( \19682 , \19539 , \19669 );
or \U$19551 ( \19683 , \19680 , \19681 , \19682 );
and \U$19552 ( \19684 , \19558 , \19562 );
and \U$19553 ( \19685 , \19562 , \19668 );
and \U$19554 ( \19686 , \19558 , \19668 );
or \U$19555 ( \19687 , \19684 , \19685 , \19686 );
and \U$19556 ( \19688 , \19543 , \19547 );
and \U$19557 ( \19689 , \19547 , \19552 );
and \U$19558 ( \19690 , \19543 , \19552 );
or \U$19559 ( \19691 , \19688 , \19689 , \19690 );
and \U$19560 ( \19692 , \19577 , \19588 );
and \U$19561 ( \19693 , \19588 , \19667 );
and \U$19562 ( \19694 , \19577 , \19667 );
or \U$19563 ( \19695 , \19692 , \19693 , \19694 );
xor \U$19564 ( \19696 , \19691 , \19695 );
and \U$19565 ( \19697 , \10584 , \4132 );
not \U$19566 ( \19698 , \19697 );
xnor \U$19567 ( \19699 , \19698 , \3925 );
and \U$19568 ( \19700 , \9897 , \4581 );
and \U$19569 ( \19701 , \10206 , \4424 );
nor \U$19570 ( \19702 , \19700 , \19701 );
xnor \U$19571 ( \19703 , \19702 , \4377 );
xor \U$19572 ( \19704 , \19699 , \19703 );
and \U$19573 ( \19705 , \9169 , \5011 );
and \U$19574 ( \19706 , \9465 , \4878 );
nor \U$19575 ( \19707 , \19705 , \19706 );
xnor \U$19576 ( \19708 , \19707 , \4762 );
xor \U$19577 ( \19709 , \19704 , \19708 );
and \U$19578 ( \19710 , \6945 , \7055 );
and \U$19579 ( \19711 , \7231 , \6675 );
nor \U$19580 ( \19712 , \19710 , \19711 );
xnor \U$19581 ( \19713 , \19712 , \6680 );
and \U$19582 ( \19714 , \6514 , \7489 );
and \U$19583 ( \19715 , \6790 , \7137 );
nor \U$19584 ( \19716 , \19714 , \19715 );
xnor \U$19585 ( \19717 , \19716 , \7142 );
xor \U$19586 ( \19718 , \19713 , \19717 );
and \U$19587 ( \19719 , \6030 , \8019 );
and \U$19588 ( \19720 , \6281 , \7830 );
nor \U$19589 ( \19721 , \19719 , \19720 );
xnor \U$19590 ( \19722 , \19721 , \7713 );
xor \U$19591 ( \19723 , \19718 , \19722 );
and \U$19592 ( \19724 , \8652 , \5485 );
and \U$19593 ( \19725 , \8835 , \5275 );
nor \U$19594 ( \19726 , \19724 , \19725 );
xnor \U$19595 ( \19727 , \19726 , \5169 );
and \U$19596 ( \19728 , \8057 , \5996 );
and \U$19597 ( \19729 , \8349 , \5695 );
nor \U$19598 ( \19730 , \19728 , \19729 );
xnor \U$19599 ( \19731 , \19730 , \5687 );
xor \U$19600 ( \19732 , \19727 , \19731 );
and \U$19601 ( \19733 , \7556 , \6401 );
and \U$19602 ( \19734 , \7700 , \6143 );
nor \U$19603 ( \19735 , \19733 , \19734 );
xnor \U$19604 ( \19736 , \19735 , \6148 );
xor \U$19605 ( \19737 , \19732 , \19736 );
xor \U$19606 ( \19738 , \19723 , \19737 );
and \U$19607 ( \19739 , \5469 , \8540 );
and \U$19608 ( \19740 , \5674 , \8292 );
nor \U$19609 ( \19741 , \19739 , \19740 );
xnor \U$19610 ( \19742 , \19741 , \8297 );
and \U$19611 ( \19743 , \4922 , \9333 );
and \U$19612 ( \19744 , \5156 , \9006 );
nor \U$19613 ( \19745 , \19743 , \19744 );
xnor \U$19614 ( \19746 , \19745 , \8848 );
xor \U$19615 ( \19747 , \19742 , \19746 );
and \U$19616 ( \19748 , \4654 , \9765 );
and \U$19617 ( \19749 , \4749 , \9644 );
nor \U$19618 ( \19750 , \19748 , \19749 );
xnor \U$19619 ( \19751 , \19750 , \9478 );
xor \U$19620 ( \19752 , \19747 , \19751 );
xor \U$19621 ( \19753 , \19738 , \19752 );
xor \U$19622 ( \19754 , \19709 , \19753 );
and \U$19623 ( \19755 , \19613 , \19617 );
and \U$19624 ( \19756 , \19617 , \19619 );
and \U$19625 ( \19757 , \19613 , \19619 );
or \U$19626 ( \19758 , \19755 , \19756 , \19757 );
and \U$19627 ( \19759 , \19640 , \19644 );
and \U$19628 ( \19760 , \19644 , \19649 );
and \U$19629 ( \19761 , \19640 , \19649 );
or \U$19630 ( \19762 , \19759 , \19760 , \19761 );
xor \U$19631 ( \19763 , \19758 , \19762 );
and \U$19632 ( \19764 , \4160 , \10408 );
and \U$19633 ( \19765 , \4364 , \10116 );
nor \U$19634 ( \19766 , \19764 , \19765 );
xnor \U$19635 ( \19767 , \19766 , \10121 );
and \U$19636 ( \19768 , \3912 , \10118 );
xnor \U$19637 ( \19769 , \19767 , \19768 );
xor \U$19638 ( \19770 , \19763 , \19769 );
xor \U$19639 ( \19771 , \19754 , \19770 );
xor \U$19640 ( \19772 , \19696 , \19771 );
xor \U$19641 ( \19773 , \19687 , \19772 );
and \U$19642 ( \19774 , \19567 , \19571 );
and \U$19643 ( \19775 , \19571 , \19576 );
and \U$19644 ( \19776 , \19567 , \19576 );
or \U$19645 ( \19777 , \19774 , \19775 , \19776 );
and \U$19646 ( \19778 , \19604 , \19608 );
and \U$19647 ( \19779 , \19608 , \19620 );
and \U$19648 ( \19780 , \19604 , \19620 );
or \U$19649 ( \19781 , \19778 , \19779 , \19780 );
xor \U$19650 ( \19782 , \19777 , \19781 );
and \U$19651 ( \19783 , \19636 , \19650 );
and \U$19652 ( \19784 , \19650 , \19665 );
and \U$19653 ( \19785 , \19636 , \19665 );
or \U$19654 ( \19786 , \19783 , \19784 , \19785 );
xor \U$19655 ( \19787 , \19782 , \19786 );
and \U$19656 ( \19788 , \19581 , \19585 );
and \U$19657 ( \19789 , \19585 , \19587 );
and \U$19658 ( \19790 , \19581 , \19587 );
or \U$19659 ( \19791 , \19788 , \19789 , \19790 );
and \U$19660 ( \19792 , \19600 , \19621 );
and \U$19661 ( \19793 , \19621 , \19666 );
and \U$19662 ( \19794 , \19600 , \19666 );
or \U$19663 ( \19795 , \19792 , \19793 , \19794 );
xor \U$19664 ( \19796 , \19791 , \19795 );
and \U$19665 ( \19797 , \19590 , \19594 );
and \U$19666 ( \19798 , \19594 , \19599 );
and \U$19667 ( \19799 , \19590 , \19599 );
or \U$19668 ( \19800 , \19797 , \19798 , \19799 );
and \U$19669 ( \19801 , \19626 , \19630 );
and \U$19670 ( \19802 , \19630 , \19635 );
and \U$19671 ( \19803 , \19626 , \19635 );
or \U$19672 ( \19804 , \19801 , \19802 , \19803 );
xor \U$19673 ( \19805 , \19800 , \19804 );
and \U$19674 ( \19806 , \19655 , \19659 );
and \U$19675 ( \19807 , \19659 , \19664 );
and \U$19676 ( \19808 , \19655 , \19664 );
or \U$19677 ( \19809 , \19806 , \19807 , \19808 );
xor \U$19678 ( \19810 , \19805 , \19809 );
xor \U$19679 ( \19811 , \19796 , \19810 );
xor \U$19680 ( \19812 , \19787 , \19811 );
xor \U$19681 ( \19813 , \19773 , \19812 );
xor \U$19682 ( \19814 , \19683 , \19813 );
and \U$19683 ( \19815 , \19535 , \19670 );
xor \U$19684 ( \19816 , \19814 , \19815 );
and \U$19685 ( \19817 , \19671 , \19672 );
and \U$19686 ( \19818 , \19673 , \19676 );
or \U$19687 ( \19819 , \19817 , \19818 );
xor \U$19688 ( \19820 , \19816 , \19819 );
buf \U$19689 ( \19821 , \19820 );
buf \U$19690 ( \19822 , \19821 );
and \U$19691 ( \19823 , \19687 , \19772 );
and \U$19692 ( \19824 , \19772 , \19812 );
and \U$19693 ( \19825 , \19687 , \19812 );
or \U$19694 ( \19826 , \19823 , \19824 , \19825 );
and \U$19695 ( \19827 , \19691 , \19695 );
and \U$19696 ( \19828 , \19695 , \19771 );
and \U$19697 ( \19829 , \19691 , \19771 );
or \U$19698 ( \19830 , \19827 , \19828 , \19829 );
and \U$19699 ( \19831 , \19787 , \19811 );
xor \U$19700 ( \19832 , \19830 , \19831 );
and \U$19701 ( \19833 , \19791 , \19795 );
and \U$19702 ( \19834 , \19795 , \19810 );
and \U$19703 ( \19835 , \19791 , \19810 );
or \U$19704 ( \19836 , \19833 , \19834 , \19835 );
and \U$19705 ( \19837 , \19777 , \19781 );
and \U$19706 ( \19838 , \19781 , \19786 );
and \U$19707 ( \19839 , \19777 , \19786 );
or \U$19708 ( \19840 , \19837 , \19838 , \19839 );
and \U$19709 ( \19841 , \19709 , \19753 );
and \U$19710 ( \19842 , \19753 , \19770 );
and \U$19711 ( \19843 , \19709 , \19770 );
or \U$19712 ( \19844 , \19841 , \19842 , \19843 );
xor \U$19713 ( \19845 , \19840 , \19844 );
and \U$19714 ( \19846 , \19742 , \19746 );
and \U$19715 ( \19847 , \19746 , \19751 );
and \U$19716 ( \19848 , \19742 , \19751 );
or \U$19717 ( \19849 , \19846 , \19847 , \19848 );
or \U$19718 ( \19850 , \19767 , \19768 );
xor \U$19719 ( \19851 , \19849 , \19850 );
and \U$19720 ( \19852 , \4364 , \10408 );
and \U$19721 ( \19853 , \4654 , \10116 );
nor \U$19722 ( \19854 , \19852 , \19853 );
xnor \U$19723 ( \19855 , \19854 , \10121 );
xor \U$19724 ( \19856 , \19851 , \19855 );
xor \U$19725 ( \19857 , \19845 , \19856 );
xor \U$19726 ( \19858 , \19836 , \19857 );
and \U$19727 ( \19859 , \19713 , \19717 );
and \U$19728 ( \19860 , \19717 , \19722 );
and \U$19729 ( \19861 , \19713 , \19722 );
or \U$19730 ( \19862 , \19859 , \19860 , \19861 );
and \U$19731 ( \19863 , \19727 , \19731 );
and \U$19732 ( \19864 , \19731 , \19736 );
and \U$19733 ( \19865 , \19727 , \19736 );
or \U$19734 ( \19866 , \19863 , \19864 , \19865 );
xor \U$19735 ( \19867 , \19862 , \19866 );
and \U$19736 ( \19868 , \19699 , \19703 );
and \U$19737 ( \19869 , \19703 , \19708 );
and \U$19738 ( \19870 , \19699 , \19708 );
or \U$19739 ( \19871 , \19868 , \19869 , \19870 );
xor \U$19740 ( \19872 , \19867 , \19871 );
and \U$19741 ( \19873 , \19800 , \19804 );
and \U$19742 ( \19874 , \19804 , \19809 );
and \U$19743 ( \19875 , \19800 , \19809 );
or \U$19744 ( \19876 , \19873 , \19874 , \19875 );
and \U$19745 ( \19877 , \19723 , \19737 );
and \U$19746 ( \19878 , \19737 , \19752 );
and \U$19747 ( \19879 , \19723 , \19752 );
or \U$19748 ( \19880 , \19877 , \19878 , \19879 );
xor \U$19749 ( \19881 , \19876 , \19880 );
and \U$19750 ( \19882 , \19758 , \19762 );
and \U$19751 ( \19883 , \19762 , \19769 );
and \U$19752 ( \19884 , \19758 , \19769 );
or \U$19753 ( \19885 , \19882 , \19883 , \19884 );
xor \U$19754 ( \19886 , \19881 , \19885 );
xor \U$19755 ( \19887 , \19872 , \19886 );
and \U$19756 ( \19888 , \8835 , \5485 );
and \U$19757 ( \19889 , \9169 , \5275 );
nor \U$19758 ( \19890 , \19888 , \19889 );
xnor \U$19759 ( \19891 , \19890 , \5169 );
and \U$19760 ( \19892 , \8349 , \5996 );
and \U$19761 ( \19893 , \8652 , \5695 );
nor \U$19762 ( \19894 , \19892 , \19893 );
xnor \U$19763 ( \19895 , \19894 , \5687 );
xor \U$19764 ( \19896 , \19891 , \19895 );
and \U$19765 ( \19897 , \7700 , \6401 );
and \U$19766 ( \19898 , \8057 , \6143 );
nor \U$19767 ( \19899 , \19897 , \19898 );
xnor \U$19768 ( \19900 , \19899 , \6148 );
xor \U$19769 ( \19901 , \19896 , \19900 );
not \U$19770 ( \19902 , \3925 );
and \U$19771 ( \19903 , \10206 , \4581 );
and \U$19772 ( \19904 , \10584 , \4424 );
nor \U$19773 ( \19905 , \19903 , \19904 );
xnor \U$19774 ( \19906 , \19905 , \4377 );
xor \U$19775 ( \19907 , \19902 , \19906 );
and \U$19776 ( \19908 , \9465 , \5011 );
and \U$19777 ( \19909 , \9897 , \4878 );
nor \U$19778 ( \19910 , \19908 , \19909 );
xnor \U$19779 ( \19911 , \19910 , \4762 );
xor \U$19780 ( \19912 , \19907 , \19911 );
xor \U$19781 ( \19913 , \19901 , \19912 );
and \U$19782 ( \19914 , \4160 , \10118 );
and \U$19783 ( \19915 , \7231 , \7055 );
and \U$19784 ( \19916 , \7556 , \6675 );
nor \U$19785 ( \19917 , \19915 , \19916 );
xnor \U$19786 ( \19918 , \19917 , \6680 );
and \U$19787 ( \19919 , \6790 , \7489 );
and \U$19788 ( \19920 , \6945 , \7137 );
nor \U$19789 ( \19921 , \19919 , \19920 );
xnor \U$19790 ( \19922 , \19921 , \7142 );
xor \U$19791 ( \19923 , \19918 , \19922 );
and \U$19792 ( \19924 , \6281 , \8019 );
and \U$19793 ( \19925 , \6514 , \7830 );
nor \U$19794 ( \19926 , \19924 , \19925 );
xnor \U$19795 ( \19927 , \19926 , \7713 );
xor \U$19796 ( \19928 , \19923 , \19927 );
xor \U$19797 ( \19929 , \19914 , \19928 );
and \U$19798 ( \19930 , \5674 , \8540 );
and \U$19799 ( \19931 , \6030 , \8292 );
nor \U$19800 ( \19932 , \19930 , \19931 );
xnor \U$19801 ( \19933 , \19932 , \8297 );
and \U$19802 ( \19934 , \5156 , \9333 );
and \U$19803 ( \19935 , \5469 , \9006 );
nor \U$19804 ( \19936 , \19934 , \19935 );
xnor \U$19805 ( \19937 , \19936 , \8848 );
xor \U$19806 ( \19938 , \19933 , \19937 );
and \U$19807 ( \19939 , \4749 , \9765 );
and \U$19808 ( \19940 , \4922 , \9644 );
nor \U$19809 ( \19941 , \19939 , \19940 );
xnor \U$19810 ( \19942 , \19941 , \9478 );
xor \U$19811 ( \19943 , \19938 , \19942 );
xor \U$19812 ( \19944 , \19929 , \19943 );
xor \U$19813 ( \19945 , \19913 , \19944 );
xor \U$19814 ( \19946 , \19887 , \19945 );
xor \U$19815 ( \19947 , \19858 , \19946 );
xor \U$19816 ( \19948 , \19832 , \19947 );
xor \U$19817 ( \19949 , \19826 , \19948 );
and \U$19818 ( \19950 , \19683 , \19813 );
xor \U$19819 ( \19951 , \19949 , \19950 );
and \U$19820 ( \19952 , \19814 , \19815 );
and \U$19821 ( \19953 , \19816 , \19819 );
or \U$19822 ( \19954 , \19952 , \19953 );
xor \U$19823 ( \19955 , \19951 , \19954 );
buf \U$19824 ( \19956 , \19955 );
buf \U$19825 ( \19957 , \19956 );
and \U$19826 ( \19958 , \19830 , \19831 );
and \U$19827 ( \19959 , \19831 , \19947 );
and \U$19828 ( \19960 , \19830 , \19947 );
or \U$19829 ( \19961 , \19958 , \19959 , \19960 );
and \U$19830 ( \19962 , \19836 , \19857 );
and \U$19831 ( \19963 , \19857 , \19946 );
and \U$19832 ( \19964 , \19836 , \19946 );
or \U$19833 ( \19965 , \19962 , \19963 , \19964 );
and \U$19834 ( \19966 , \19840 , \19844 );
and \U$19835 ( \19967 , \19844 , \19856 );
and \U$19836 ( \19968 , \19840 , \19856 );
or \U$19837 ( \19969 , \19966 , \19967 , \19968 );
and \U$19838 ( \19970 , \19872 , \19886 );
and \U$19839 ( \19971 , \19886 , \19945 );
and \U$19840 ( \19972 , \19872 , \19945 );
or \U$19841 ( \19973 , \19970 , \19971 , \19972 );
xor \U$19842 ( \19974 , \19969 , \19973 );
and \U$19843 ( \19975 , \19849 , \19850 );
and \U$19844 ( \19976 , \19850 , \19855 );
and \U$19845 ( \19977 , \19849 , \19855 );
or \U$19846 ( \19978 , \19975 , \19976 , \19977 );
and \U$19847 ( \19979 , \19862 , \19866 );
and \U$19848 ( \19980 , \19866 , \19871 );
and \U$19849 ( \19981 , \19862 , \19871 );
or \U$19850 ( \19982 , \19979 , \19980 , \19981 );
xor \U$19851 ( \19983 , \19978 , \19982 );
and \U$19852 ( \19984 , \19914 , \19928 );
and \U$19853 ( \19985 , \19928 , \19943 );
and \U$19854 ( \19986 , \19914 , \19943 );
or \U$19855 ( \19987 , \19984 , \19985 , \19986 );
xor \U$19856 ( \19988 , \19983 , \19987 );
xor \U$19857 ( \19989 , \19974 , \19988 );
xor \U$19858 ( \19990 , \19965 , \19989 );
and \U$19859 ( \19991 , \19876 , \19880 );
and \U$19860 ( \19992 , \19880 , \19885 );
and \U$19861 ( \19993 , \19876 , \19885 );
or \U$19862 ( \19994 , \19991 , \19992 , \19993 );
and \U$19863 ( \19995 , \19901 , \19912 );
and \U$19864 ( \19996 , \19912 , \19944 );
and \U$19865 ( \19997 , \19901 , \19944 );
or \U$19866 ( \19998 , \19995 , \19996 , \19997 );
xor \U$19867 ( \19999 , \19994 , \19998 );
and \U$19868 ( \20000 , \19918 , \19922 );
and \U$19869 ( \20001 , \19922 , \19927 );
and \U$19870 ( \20002 , \19918 , \19927 );
or \U$19871 ( \20003 , \20000 , \20001 , \20002 );
and \U$19872 ( \20004 , \19891 , \19895 );
and \U$19873 ( \20005 , \19895 , \19900 );
and \U$19874 ( \20006 , \19891 , \19900 );
or \U$19875 ( \20007 , \20004 , \20005 , \20006 );
xor \U$19876 ( \20008 , \20003 , \20007 );
and \U$19877 ( \20009 , \19902 , \19906 );
and \U$19878 ( \20010 , \19906 , \19911 );
and \U$19879 ( \20011 , \19902 , \19911 );
or \U$19880 ( \20012 , \20009 , \20010 , \20011 );
xor \U$19881 ( \20013 , \20008 , \20012 );
and \U$19882 ( \20014 , \8652 , \5996 );
and \U$19883 ( \20015 , \8835 , \5695 );
nor \U$19884 ( \20016 , \20014 , \20015 );
xnor \U$19885 ( \20017 , \20016 , \5687 );
and \U$19886 ( \20018 , \8057 , \6401 );
and \U$19887 ( \20019 , \8349 , \6143 );
nor \U$19888 ( \20020 , \20018 , \20019 );
xnor \U$19889 ( \20021 , \20020 , \6148 );
xor \U$19890 ( \20022 , \20017 , \20021 );
and \U$19891 ( \20023 , \7556 , \7055 );
and \U$19892 ( \20024 , \7700 , \6675 );
nor \U$19893 ( \20025 , \20023 , \20024 );
xnor \U$19894 ( \20026 , \20025 , \6680 );
xor \U$19895 ( \20027 , \20022 , \20026 );
and \U$19896 ( \20028 , \10584 , \4581 );
not \U$19897 ( \20029 , \20028 );
xnor \U$19898 ( \20030 , \20029 , \4377 );
and \U$19899 ( \20031 , \9897 , \5011 );
and \U$19900 ( \20032 , \10206 , \4878 );
nor \U$19901 ( \20033 , \20031 , \20032 );
xnor \U$19902 ( \20034 , \20033 , \4762 );
xor \U$19903 ( \20035 , \20030 , \20034 );
and \U$19904 ( \20036 , \9169 , \5485 );
and \U$19905 ( \20037 , \9465 , \5275 );
nor \U$19906 ( \20038 , \20036 , \20037 );
xnor \U$19907 ( \20039 , \20038 , \5169 );
xor \U$19908 ( \20040 , \20035 , \20039 );
xor \U$19909 ( \20041 , \20027 , \20040 );
and \U$19910 ( \20042 , \6945 , \7489 );
and \U$19911 ( \20043 , \7231 , \7137 );
nor \U$19912 ( \20044 , \20042 , \20043 );
xnor \U$19913 ( \20045 , \20044 , \7142 );
and \U$19914 ( \20046 , \6514 , \8019 );
and \U$19915 ( \20047 , \6790 , \7830 );
nor \U$19916 ( \20048 , \20046 , \20047 );
xnor \U$19917 ( \20049 , \20048 , \7713 );
xor \U$19918 ( \20050 , \20045 , \20049 );
and \U$19919 ( \20051 , \6030 , \8540 );
and \U$19920 ( \20052 , \6281 , \8292 );
nor \U$19921 ( \20053 , \20051 , \20052 );
xnor \U$19922 ( \20054 , \20053 , \8297 );
xor \U$19923 ( \20055 , \20050 , \20054 );
xor \U$19924 ( \20056 , \20041 , \20055 );
xor \U$19925 ( \20057 , \20013 , \20056 );
and \U$19926 ( \20058 , \19933 , \19937 );
and \U$19927 ( \20059 , \19937 , \19942 );
and \U$19928 ( \20060 , \19933 , \19942 );
or \U$19929 ( \20061 , \20058 , \20059 , \20060 );
and \U$19930 ( \20062 , \5469 , \9333 );
and \U$19931 ( \20063 , \5674 , \9006 );
nor \U$19932 ( \20064 , \20062 , \20063 );
xnor \U$19933 ( \20065 , \20064 , \8848 );
and \U$19934 ( \20066 , \4922 , \9765 );
and \U$19935 ( \20067 , \5156 , \9644 );
nor \U$19936 ( \20068 , \20066 , \20067 );
xnor \U$19937 ( \20069 , \20068 , \9478 );
xor \U$19938 ( \20070 , \20065 , \20069 );
and \U$19939 ( \20071 , \4654 , \10408 );
and \U$19940 ( \20072 , \4749 , \10116 );
nor \U$19941 ( \20073 , \20071 , \20072 );
xnor \U$19942 ( \20074 , \20073 , \10121 );
xor \U$19943 ( \20075 , \20070 , \20074 );
xor \U$19944 ( \20076 , \20061 , \20075 );
and \U$19945 ( \20077 , \4364 , \10118 );
not \U$19946 ( \20078 , \20077 );
xor \U$19947 ( \20079 , \20076 , \20078 );
xor \U$19948 ( \20080 , \20057 , \20079 );
xor \U$19949 ( \20081 , \19999 , \20080 );
xor \U$19950 ( \20082 , \19990 , \20081 );
xor \U$19951 ( \20083 , \19961 , \20082 );
and \U$19952 ( \20084 , \19826 , \19948 );
xor \U$19953 ( \20085 , \20083 , \20084 );
and \U$19954 ( \20086 , \19949 , \19950 );
and \U$19955 ( \20087 , \19951 , \19954 );
or \U$19956 ( \20088 , \20086 , \20087 );
xor \U$19957 ( \20089 , \20085 , \20088 );
buf \U$19958 ( \20090 , \20089 );
buf \U$19959 ( \20091 , \20090 );
and \U$19960 ( \20092 , \19969 , \19973 );
and \U$19961 ( \20093 , \19973 , \19988 );
and \U$19962 ( \20094 , \19969 , \19988 );
or \U$19963 ( \20095 , \20092 , \20093 , \20094 );
and \U$19964 ( \20096 , \19965 , \19989 );
and \U$19965 ( \20097 , \19989 , \20081 );
and \U$19966 ( \20098 , \19965 , \20081 );
or \U$19967 ( \20099 , \20096 , \20097 , \20098 );
xor \U$19968 ( \20100 , \20095 , \20099 );
and \U$19969 ( \20101 , \19994 , \19998 );
and \U$19970 ( \20102 , \19998 , \20080 );
and \U$19971 ( \20103 , \19994 , \20080 );
or \U$19972 ( \20104 , \20101 , \20102 , \20103 );
and \U$19973 ( \20105 , \19978 , \19982 );
and \U$19974 ( \20106 , \19982 , \19987 );
and \U$19975 ( \20107 , \19978 , \19987 );
or \U$19976 ( \20108 , \20105 , \20106 , \20107 );
and \U$19977 ( \20109 , \20013 , \20056 );
and \U$19978 ( \20110 , \20056 , \20079 );
and \U$19979 ( \20111 , \20013 , \20079 );
or \U$19980 ( \20112 , \20109 , \20110 , \20111 );
xor \U$19981 ( \20113 , \20108 , \20112 );
and \U$19982 ( \20114 , \20017 , \20021 );
and \U$19983 ( \20115 , \20021 , \20026 );
and \U$19984 ( \20116 , \20017 , \20026 );
or \U$19985 ( \20117 , \20114 , \20115 , \20116 );
and \U$19986 ( \20118 , \20030 , \20034 );
and \U$19987 ( \20119 , \20034 , \20039 );
and \U$19988 ( \20120 , \20030 , \20039 );
or \U$19989 ( \20121 , \20118 , \20119 , \20120 );
xor \U$19990 ( \20122 , \20117 , \20121 );
and \U$19991 ( \20123 , \20045 , \20049 );
and \U$19992 ( \20124 , \20049 , \20054 );
and \U$19993 ( \20125 , \20045 , \20054 );
or \U$19994 ( \20126 , \20123 , \20124 , \20125 );
xor \U$19995 ( \20127 , \20122 , \20126 );
xor \U$19996 ( \20128 , \20113 , \20127 );
xor \U$19997 ( \20129 , \20104 , \20128 );
and \U$19998 ( \20130 , \20003 , \20007 );
and \U$19999 ( \20131 , \20007 , \20012 );
and \U$20000 ( \20132 , \20003 , \20012 );
or \U$20001 ( \20133 , \20130 , \20131 , \20132 );
and \U$20002 ( \20134 , \20027 , \20040 );
and \U$20003 ( \20135 , \20040 , \20055 );
and \U$20004 ( \20136 , \20027 , \20055 );
or \U$20005 ( \20137 , \20134 , \20135 , \20136 );
xor \U$20006 ( \20138 , \20133 , \20137 );
and \U$20007 ( \20139 , \20061 , \20075 );
and \U$20008 ( \20140 , \20075 , \20078 );
and \U$20009 ( \20141 , \20061 , \20078 );
or \U$20010 ( \20142 , \20139 , \20140 , \20141 );
xor \U$20011 ( \20143 , \20138 , \20142 );
not \U$20012 ( \20144 , \4377 );
and \U$20013 ( \20145 , \10206 , \5011 );
and \U$20014 ( \20146 , \10584 , \4878 );
nor \U$20015 ( \20147 , \20145 , \20146 );
xnor \U$20016 ( \20148 , \20147 , \4762 );
xor \U$20017 ( \20149 , \20144 , \20148 );
and \U$20018 ( \20150 , \9465 , \5485 );
and \U$20019 ( \20151 , \9897 , \5275 );
nor \U$20020 ( \20152 , \20150 , \20151 );
xnor \U$20021 ( \20153 , \20152 , \5169 );
xor \U$20022 ( \20154 , \20149 , \20153 );
and \U$20023 ( \20155 , \20065 , \20069 );
and \U$20024 ( \20156 , \20069 , \20074 );
and \U$20025 ( \20157 , \20065 , \20074 );
or \U$20026 ( \20158 , \20155 , \20156 , \20157 );
buf \U$20027 ( \20159 , \20077 );
xor \U$20028 ( \20160 , \20158 , \20159 );
and \U$20029 ( \20161 , \4654 , \10118 );
xor \U$20030 ( \20162 , \20160 , \20161 );
xor \U$20031 ( \20163 , \20154 , \20162 );
and \U$20032 ( \20164 , \8835 , \5996 );
and \U$20033 ( \20165 , \9169 , \5695 );
nor \U$20034 ( \20166 , \20164 , \20165 );
xnor \U$20035 ( \20167 , \20166 , \5687 );
and \U$20036 ( \20168 , \8349 , \6401 );
and \U$20037 ( \20169 , \8652 , \6143 );
nor \U$20038 ( \20170 , \20168 , \20169 );
xnor \U$20039 ( \20171 , \20170 , \6148 );
xor \U$20040 ( \20172 , \20167 , \20171 );
and \U$20041 ( \20173 , \7700 , \7055 );
and \U$20042 ( \20174 , \8057 , \6675 );
nor \U$20043 ( \20175 , \20173 , \20174 );
xnor \U$20044 ( \20176 , \20175 , \6680 );
xor \U$20045 ( \20177 , \20172 , \20176 );
and \U$20046 ( \20178 , \5674 , \9333 );
and \U$20047 ( \20179 , \6030 , \9006 );
nor \U$20048 ( \20180 , \20178 , \20179 );
xnor \U$20049 ( \20181 , \20180 , \8848 );
and \U$20050 ( \20182 , \5156 , \9765 );
and \U$20051 ( \20183 , \5469 , \9644 );
nor \U$20052 ( \20184 , \20182 , \20183 );
xnor \U$20053 ( \20185 , \20184 , \9478 );
xor \U$20054 ( \20186 , \20181 , \20185 );
and \U$20055 ( \20187 , \4749 , \10408 );
and \U$20056 ( \20188 , \4922 , \10116 );
nor \U$20057 ( \20189 , \20187 , \20188 );
xnor \U$20058 ( \20190 , \20189 , \10121 );
xor \U$20059 ( \20191 , \20186 , \20190 );
xor \U$20060 ( \20192 , \20177 , \20191 );
and \U$20061 ( \20193 , \7231 , \7489 );
and \U$20062 ( \20194 , \7556 , \7137 );
nor \U$20063 ( \20195 , \20193 , \20194 );
xnor \U$20064 ( \20196 , \20195 , \7142 );
and \U$20065 ( \20197 , \6790 , \8019 );
and \U$20066 ( \20198 , \6945 , \7830 );
nor \U$20067 ( \20199 , \20197 , \20198 );
xnor \U$20068 ( \20200 , \20199 , \7713 );
xor \U$20069 ( \20201 , \20196 , \20200 );
and \U$20070 ( \20202 , \6281 , \8540 );
and \U$20071 ( \20203 , \6514 , \8292 );
nor \U$20072 ( \20204 , \20202 , \20203 );
xnor \U$20073 ( \20205 , \20204 , \8297 );
xor \U$20074 ( \20206 , \20201 , \20205 );
xor \U$20075 ( \20207 , \20192 , \20206 );
xor \U$20076 ( \20208 , \20163 , \20207 );
xor \U$20077 ( \20209 , \20143 , \20208 );
xor \U$20078 ( \20210 , \20129 , \20209 );
xor \U$20079 ( \20211 , \20100 , \20210 );
and \U$20080 ( \20212 , \19961 , \20082 );
xor \U$20081 ( \20213 , \20211 , \20212 );
and \U$20082 ( \20214 , \20083 , \20084 );
and \U$20083 ( \20215 , \20085 , \20088 );
or \U$20084 ( \20216 , \20214 , \20215 );
xor \U$20085 ( \20217 , \20213 , \20216 );
buf \U$20086 ( \20218 , \20217 );
buf \U$20087 ( \20219 , \20218 );
and \U$20088 ( \20220 , \20104 , \20128 );
and \U$20089 ( \20221 , \20128 , \20209 );
and \U$20090 ( \20222 , \20104 , \20209 );
or \U$20091 ( \20223 , \20220 , \20221 , \20222 );
and \U$20092 ( \20224 , \20108 , \20112 );
and \U$20093 ( \20225 , \20112 , \20127 );
and \U$20094 ( \20226 , \20108 , \20127 );
or \U$20095 ( \20227 , \20224 , \20225 , \20226 );
and \U$20096 ( \20228 , \20143 , \20208 );
xor \U$20097 ( \20229 , \20227 , \20228 );
and \U$20098 ( \20230 , \20158 , \20159 );
and \U$20099 ( \20231 , \20159 , \20161 );
and \U$20100 ( \20232 , \20158 , \20161 );
or \U$20101 ( \20233 , \20230 , \20231 , \20232 );
and \U$20102 ( \20234 , \20117 , \20121 );
and \U$20103 ( \20235 , \20121 , \20126 );
and \U$20104 ( \20236 , \20117 , \20126 );
or \U$20105 ( \20237 , \20234 , \20235 , \20236 );
xor \U$20106 ( \20238 , \20233 , \20237 );
and \U$20107 ( \20239 , \20177 , \20191 );
and \U$20108 ( \20240 , \20191 , \20206 );
and \U$20109 ( \20241 , \20177 , \20206 );
or \U$20110 ( \20242 , \20239 , \20240 , \20241 );
xor \U$20111 ( \20243 , \20238 , \20242 );
xor \U$20112 ( \20244 , \20229 , \20243 );
xor \U$20113 ( \20245 , \20223 , \20244 );
and \U$20114 ( \20246 , \20133 , \20137 );
and \U$20115 ( \20247 , \20137 , \20142 );
and \U$20116 ( \20248 , \20133 , \20142 );
or \U$20117 ( \20249 , \20246 , \20247 , \20248 );
and \U$20118 ( \20250 , \20154 , \20162 );
and \U$20119 ( \20251 , \20162 , \20207 );
and \U$20120 ( \20252 , \20154 , \20207 );
or \U$20121 ( \20253 , \20250 , \20251 , \20252 );
xor \U$20122 ( \20254 , \20249 , \20253 );
and \U$20123 ( \20255 , \20144 , \20148 );
and \U$20124 ( \20256 , \20148 , \20153 );
and \U$20125 ( \20257 , \20144 , \20153 );
or \U$20126 ( \20258 , \20255 , \20256 , \20257 );
and \U$20127 ( \20259 , \20167 , \20171 );
and \U$20128 ( \20260 , \20171 , \20176 );
and \U$20129 ( \20261 , \20167 , \20176 );
or \U$20130 ( \20262 , \20259 , \20260 , \20261 );
xor \U$20131 ( \20263 , \20258 , \20262 );
and \U$20132 ( \20264 , \20196 , \20200 );
and \U$20133 ( \20265 , \20200 , \20205 );
and \U$20134 ( \20266 , \20196 , \20205 );
or \U$20135 ( \20267 , \20264 , \20265 , \20266 );
xor \U$20136 ( \20268 , \20263 , \20267 );
and \U$20137 ( \20269 , \10584 , \5011 );
not \U$20138 ( \20270 , \20269 );
xnor \U$20139 ( \20271 , \20270 , \4762 );
and \U$20140 ( \20272 , \9897 , \5485 );
and \U$20141 ( \20273 , \10206 , \5275 );
nor \U$20142 ( \20274 , \20272 , \20273 );
xnor \U$20143 ( \20275 , \20274 , \5169 );
xor \U$20144 ( \20276 , \20271 , \20275 );
and \U$20145 ( \20277 , \9169 , \5996 );
and \U$20146 ( \20278 , \9465 , \5695 );
nor \U$20147 ( \20279 , \20277 , \20278 );
xnor \U$20148 ( \20280 , \20279 , \5687 );
xor \U$20149 ( \20281 , \20276 , \20280 );
and \U$20150 ( \20282 , \6945 , \8019 );
and \U$20151 ( \20283 , \7231 , \7830 );
nor \U$20152 ( \20284 , \20282 , \20283 );
xnor \U$20153 ( \20285 , \20284 , \7713 );
and \U$20154 ( \20286 , \6514 , \8540 );
and \U$20155 ( \20287 , \6790 , \8292 );
nor \U$20156 ( \20288 , \20286 , \20287 );
xnor \U$20157 ( \20289 , \20288 , \8297 );
xor \U$20158 ( \20290 , \20285 , \20289 );
and \U$20159 ( \20291 , \6030 , \9333 );
and \U$20160 ( \20292 , \6281 , \9006 );
nor \U$20161 ( \20293 , \20291 , \20292 );
xnor \U$20162 ( \20294 , \20293 , \8848 );
xor \U$20163 ( \20295 , \20290 , \20294 );
xor \U$20164 ( \20296 , \20281 , \20295 );
and \U$20165 ( \20297 , \8652 , \6401 );
and \U$20166 ( \20298 , \8835 , \6143 );
nor \U$20167 ( \20299 , \20297 , \20298 );
xnor \U$20168 ( \20300 , \20299 , \6148 );
and \U$20169 ( \20301 , \8057 , \7055 );
and \U$20170 ( \20302 , \8349 , \6675 );
nor \U$20171 ( \20303 , \20301 , \20302 );
xnor \U$20172 ( \20304 , \20303 , \6680 );
xor \U$20173 ( \20305 , \20300 , \20304 );
and \U$20174 ( \20306 , \7556 , \7489 );
and \U$20175 ( \20307 , \7700 , \7137 );
nor \U$20176 ( \20308 , \20306 , \20307 );
xnor \U$20177 ( \20309 , \20308 , \7142 );
xor \U$20178 ( \20310 , \20305 , \20309 );
xor \U$20179 ( \20311 , \20296 , \20310 );
xor \U$20180 ( \20312 , \20268 , \20311 );
and \U$20181 ( \20313 , \20181 , \20185 );
and \U$20182 ( \20314 , \20185 , \20190 );
and \U$20183 ( \20315 , \20181 , \20190 );
or \U$20184 ( \20316 , \20313 , \20314 , \20315 );
and \U$20185 ( \20317 , \5469 , \9765 );
and \U$20186 ( \20318 , \5674 , \9644 );
nor \U$20187 ( \20319 , \20317 , \20318 );
xnor \U$20188 ( \20320 , \20319 , \9478 );
and \U$20189 ( \20321 , \4922 , \10408 );
and \U$20190 ( \20322 , \5156 , \10116 );
nor \U$20191 ( \20323 , \20321 , \20322 );
xnor \U$20192 ( \20324 , \20323 , \10121 );
xor \U$20193 ( \20325 , \20320 , \20324 );
and \U$20194 ( \20326 , \4749 , \10118 );
xor \U$20195 ( \20327 , \20325 , \20326 );
xnor \U$20196 ( \20328 , \20316 , \20327 );
xor \U$20197 ( \20329 , \20312 , \20328 );
xor \U$20198 ( \20330 , \20254 , \20329 );
xor \U$20199 ( \20331 , \20245 , \20330 );
and \U$20200 ( \20332 , \20095 , \20099 );
and \U$20201 ( \20333 , \20099 , \20210 );
and \U$20202 ( \20334 , \20095 , \20210 );
or \U$20203 ( \20335 , \20332 , \20333 , \20334 );
xor \U$20204 ( \20336 , \20331 , \20335 );
and \U$20205 ( \20337 , \20211 , \20212 );
and \U$20206 ( \20338 , \20213 , \20216 );
or \U$20207 ( \20339 , \20337 , \20338 );
xor \U$20208 ( \20340 , \20336 , \20339 );
buf \U$20209 ( \20341 , \20340 );
buf \U$20210 ( \20342 , \20341 );
and \U$20211 ( \20343 , \20227 , \20228 );
and \U$20212 ( \20344 , \20228 , \20243 );
and \U$20213 ( \20345 , \20227 , \20243 );
or \U$20214 ( \20346 , \20343 , \20344 , \20345 );
and \U$20215 ( \20347 , \20249 , \20253 );
and \U$20216 ( \20348 , \20253 , \20329 );
and \U$20217 ( \20349 , \20249 , \20329 );
or \U$20218 ( \20350 , \20347 , \20348 , \20349 );
and \U$20219 ( \20351 , \20258 , \20262 );
and \U$20220 ( \20352 , \20262 , \20267 );
and \U$20221 ( \20353 , \20258 , \20267 );
or \U$20222 ( \20354 , \20351 , \20352 , \20353 );
and \U$20223 ( \20355 , \20281 , \20295 );
and \U$20224 ( \20356 , \20295 , \20310 );
and \U$20225 ( \20357 , \20281 , \20310 );
or \U$20226 ( \20358 , \20355 , \20356 , \20357 );
xor \U$20227 ( \20359 , \20354 , \20358 );
or \U$20228 ( \20360 , \20316 , \20327 );
xor \U$20229 ( \20361 , \20359 , \20360 );
xor \U$20230 ( \20362 , \20350 , \20361 );
and \U$20231 ( \20363 , \20233 , \20237 );
and \U$20232 ( \20364 , \20237 , \20242 );
and \U$20233 ( \20365 , \20233 , \20242 );
or \U$20234 ( \20366 , \20363 , \20364 , \20365 );
and \U$20235 ( \20367 , \20268 , \20311 );
and \U$20236 ( \20368 , \20311 , \20328 );
and \U$20237 ( \20369 , \20268 , \20328 );
or \U$20238 ( \20370 , \20367 , \20368 , \20369 );
xor \U$20239 ( \20371 , \20366 , \20370 );
and \U$20240 ( \20372 , \20271 , \20275 );
and \U$20241 ( \20373 , \20275 , \20280 );
and \U$20242 ( \20374 , \20271 , \20280 );
or \U$20243 ( \20375 , \20372 , \20373 , \20374 );
and \U$20244 ( \20376 , \20285 , \20289 );
and \U$20245 ( \20377 , \20289 , \20294 );
and \U$20246 ( \20378 , \20285 , \20294 );
or \U$20247 ( \20379 , \20376 , \20377 , \20378 );
xor \U$20248 ( \20380 , \20375 , \20379 );
and \U$20249 ( \20381 , \20300 , \20304 );
and \U$20250 ( \20382 , \20304 , \20309 );
and \U$20251 ( \20383 , \20300 , \20309 );
or \U$20252 ( \20384 , \20381 , \20382 , \20383 );
xor \U$20253 ( \20385 , \20380 , \20384 );
and \U$20254 ( \20386 , \20320 , \20324 );
and \U$20255 ( \20387 , \20324 , \20326 );
and \U$20256 ( \20388 , \20320 , \20326 );
or \U$20257 ( \20389 , \20386 , \20387 , \20388 );
and \U$20258 ( \20390 , \5674 , \9765 );
and \U$20259 ( \20391 , \6030 , \9644 );
nor \U$20260 ( \20392 , \20390 , \20391 );
xnor \U$20261 ( \20393 , \20392 , \9478 );
and \U$20262 ( \20394 , \5156 , \10408 );
and \U$20263 ( \20395 , \5469 , \10116 );
nor \U$20264 ( \20396 , \20394 , \20395 );
xnor \U$20265 ( \20397 , \20396 , \10121 );
xor \U$20266 ( \20398 , \20393 , \20397 );
and \U$20267 ( \20399 , \4922 , \10118 );
xor \U$20268 ( \20400 , \20398 , \20399 );
xor \U$20269 ( \20401 , \20389 , \20400 );
and \U$20270 ( \20402 , \7231 , \8019 );
and \U$20271 ( \20403 , \7556 , \7830 );
nor \U$20272 ( \20404 , \20402 , \20403 );
xnor \U$20273 ( \20405 , \20404 , \7713 );
and \U$20274 ( \20406 , \6790 , \8540 );
and \U$20275 ( \20407 , \6945 , \8292 );
nor \U$20276 ( \20408 , \20406 , \20407 );
xnor \U$20277 ( \20409 , \20408 , \8297 );
xor \U$20278 ( \20410 , \20405 , \20409 );
and \U$20279 ( \20411 , \6281 , \9333 );
and \U$20280 ( \20412 , \6514 , \9006 );
nor \U$20281 ( \20413 , \20411 , \20412 );
xnor \U$20282 ( \20414 , \20413 , \8848 );
xor \U$20283 ( \20415 , \20410 , \20414 );
xor \U$20284 ( \20416 , \20401 , \20415 );
xor \U$20285 ( \20417 , \20385 , \20416 );
not \U$20286 ( \20418 , \4762 );
and \U$20287 ( \20419 , \10206 , \5485 );
and \U$20288 ( \20420 , \10584 , \5275 );
nor \U$20289 ( \20421 , \20419 , \20420 );
xnor \U$20290 ( \20422 , \20421 , \5169 );
xor \U$20291 ( \20423 , \20418 , \20422 );
and \U$20292 ( \20424 , \9465 , \5996 );
and \U$20293 ( \20425 , \9897 , \5695 );
nor \U$20294 ( \20426 , \20424 , \20425 );
xnor \U$20295 ( \20427 , \20426 , \5687 );
xor \U$20296 ( \20428 , \20423 , \20427 );
and \U$20297 ( \20429 , \8835 , \6401 );
and \U$20298 ( \20430 , \9169 , \6143 );
nor \U$20299 ( \20431 , \20429 , \20430 );
xnor \U$20300 ( \20432 , \20431 , \6148 );
and \U$20301 ( \20433 , \8349 , \7055 );
and \U$20302 ( \20434 , \8652 , \6675 );
nor \U$20303 ( \20435 , \20433 , \20434 );
xnor \U$20304 ( \20436 , \20435 , \6680 );
xor \U$20305 ( \20437 , \20432 , \20436 );
and \U$20306 ( \20438 , \7700 , \7489 );
and \U$20307 ( \20439 , \8057 , \7137 );
nor \U$20308 ( \20440 , \20438 , \20439 );
xnor \U$20309 ( \20441 , \20440 , \7142 );
xor \U$20310 ( \20442 , \20437 , \20441 );
xor \U$20311 ( \20443 , \20428 , \20442 );
xor \U$20312 ( \20444 , \20417 , \20443 );
xor \U$20313 ( \20445 , \20371 , \20444 );
xor \U$20314 ( \20446 , \20362 , \20445 );
xor \U$20315 ( \20447 , \20346 , \20446 );
and \U$20316 ( \20448 , \20223 , \20244 );
and \U$20317 ( \20449 , \20244 , \20330 );
and \U$20318 ( \20450 , \20223 , \20330 );
or \U$20319 ( \20451 , \20448 , \20449 , \20450 );
xor \U$20320 ( \20452 , \20447 , \20451 );
and \U$20321 ( \20453 , \20331 , \20335 );
and \U$20322 ( \20454 , \20336 , \20339 );
or \U$20323 ( \20455 , \20453 , \20454 );
xor \U$20324 ( \20456 , \20452 , \20455 );
buf \U$20325 ( \20457 , \20456 );
buf \U$20326 ( \20458 , \20457 );
and \U$20327 ( \20459 , \20350 , \20361 );
and \U$20328 ( \20460 , \20361 , \20445 );
and \U$20329 ( \20461 , \20350 , \20445 );
or \U$20330 ( \20462 , \20459 , \20460 , \20461 );
and \U$20331 ( \20463 , \20366 , \20370 );
and \U$20332 ( \20464 , \20370 , \20444 );
and \U$20333 ( \20465 , \20366 , \20444 );
or \U$20334 ( \20466 , \20463 , \20464 , \20465 );
and \U$20335 ( \20467 , \20375 , \20379 );
and \U$20336 ( \20468 , \20379 , \20384 );
and \U$20337 ( \20469 , \20375 , \20384 );
or \U$20338 ( \20470 , \20467 , \20468 , \20469 );
and \U$20339 ( \20471 , \20389 , \20400 );
and \U$20340 ( \20472 , \20400 , \20415 );
and \U$20341 ( \20473 , \20389 , \20415 );
or \U$20342 ( \20474 , \20471 , \20472 , \20473 );
xor \U$20343 ( \20475 , \20470 , \20474 );
and \U$20344 ( \20476 , \20428 , \20442 );
xor \U$20345 ( \20477 , \20475 , \20476 );
xor \U$20346 ( \20478 , \20466 , \20477 );
and \U$20347 ( \20479 , \20354 , \20358 );
and \U$20348 ( \20480 , \20358 , \20360 );
and \U$20349 ( \20481 , \20354 , \20360 );
or \U$20350 ( \20482 , \20479 , \20480 , \20481 );
and \U$20351 ( \20483 , \20385 , \20416 );
and \U$20352 ( \20484 , \20416 , \20443 );
and \U$20353 ( \20485 , \20385 , \20443 );
or \U$20354 ( \20486 , \20483 , \20484 , \20485 );
xor \U$20355 ( \20487 , \20482 , \20486 );
and \U$20356 ( \20488 , \20418 , \20422 );
and \U$20357 ( \20489 , \20422 , \20427 );
and \U$20358 ( \20490 , \20418 , \20427 );
or \U$20359 ( \20491 , \20488 , \20489 , \20490 );
and \U$20360 ( \20492 , \20405 , \20409 );
and \U$20361 ( \20493 , \20409 , \20414 );
and \U$20362 ( \20494 , \20405 , \20414 );
or \U$20363 ( \20495 , \20492 , \20493 , \20494 );
xor \U$20364 ( \20496 , \20491 , \20495 );
and \U$20365 ( \20497 , \20432 , \20436 );
and \U$20366 ( \20498 , \20436 , \20441 );
and \U$20367 ( \20499 , \20432 , \20441 );
or \U$20368 ( \20500 , \20497 , \20498 , \20499 );
xor \U$20369 ( \20501 , \20496 , \20500 );
and \U$20370 ( \20502 , \20393 , \20397 );
and \U$20371 ( \20503 , \20397 , \20399 );
and \U$20372 ( \20504 , \20393 , \20399 );
or \U$20373 ( \20505 , \20502 , \20503 , \20504 );
and \U$20374 ( \20506 , \6945 , \8540 );
and \U$20375 ( \20507 , \7231 , \8292 );
nor \U$20376 ( \20508 , \20506 , \20507 );
xnor \U$20377 ( \20509 , \20508 , \8297 );
and \U$20378 ( \20510 , \6514 , \9333 );
and \U$20379 ( \20511 , \6790 , \9006 );
nor \U$20380 ( \20512 , \20510 , \20511 );
xnor \U$20381 ( \20513 , \20512 , \8848 );
xor \U$20382 ( \20514 , \20509 , \20513 );
and \U$20383 ( \20515 , \6030 , \9765 );
and \U$20384 ( \20516 , \6281 , \9644 );
nor \U$20385 ( \20517 , \20515 , \20516 );
xnor \U$20386 ( \20518 , \20517 , \9478 );
xor \U$20387 ( \20519 , \20514 , \20518 );
xor \U$20388 ( \20520 , \20505 , \20519 );
and \U$20389 ( \20521 , \5469 , \10408 );
and \U$20390 ( \20522 , \5674 , \10116 );
nor \U$20391 ( \20523 , \20521 , \20522 );
xnor \U$20392 ( \20524 , \20523 , \10121 );
and \U$20393 ( \20525 , \5156 , \10118 );
xnor \U$20394 ( \20526 , \20524 , \20525 );
xor \U$20395 ( \20527 , \20520 , \20526 );
xor \U$20396 ( \20528 , \20501 , \20527 );
and \U$20397 ( \20529 , \8652 , \7055 );
and \U$20398 ( \20530 , \8835 , \6675 );
nor \U$20399 ( \20531 , \20529 , \20530 );
xnor \U$20400 ( \20532 , \20531 , \6680 );
and \U$20401 ( \20533 , \8057 , \7489 );
and \U$20402 ( \20534 , \8349 , \7137 );
nor \U$20403 ( \20535 , \20533 , \20534 );
xnor \U$20404 ( \20536 , \20535 , \7142 );
xor \U$20405 ( \20537 , \20532 , \20536 );
and \U$20406 ( \20538 , \7556 , \8019 );
and \U$20407 ( \20539 , \7700 , \7830 );
nor \U$20408 ( \20540 , \20538 , \20539 );
xnor \U$20409 ( \20541 , \20540 , \7713 );
xor \U$20410 ( \20542 , \20537 , \20541 );
and \U$20411 ( \20543 , \10584 , \5485 );
not \U$20412 ( \20544 , \20543 );
xnor \U$20413 ( \20545 , \20544 , \5169 );
and \U$20414 ( \20546 , \9897 , \5996 );
and \U$20415 ( \20547 , \10206 , \5695 );
nor \U$20416 ( \20548 , \20546 , \20547 );
xnor \U$20417 ( \20549 , \20548 , \5687 );
xor \U$20418 ( \20550 , \20545 , \20549 );
and \U$20419 ( \20551 , \9169 , \6401 );
and \U$20420 ( \20552 , \9465 , \6143 );
nor \U$20421 ( \20553 , \20551 , \20552 );
xnor \U$20422 ( \20554 , \20553 , \6148 );
xor \U$20423 ( \20555 , \20550 , \20554 );
xor \U$20424 ( \20556 , \20542 , \20555 );
xor \U$20425 ( \20557 , \20528 , \20556 );
xor \U$20426 ( \20558 , \20487 , \20557 );
xor \U$20427 ( \20559 , \20478 , \20558 );
xor \U$20428 ( \20560 , \20462 , \20559 );
and \U$20429 ( \20561 , \20346 , \20446 );
xor \U$20430 ( \20562 , \20560 , \20561 );
and \U$20431 ( \20563 , \20447 , \20451 );
and \U$20432 ( \20564 , \20452 , \20455 );
or \U$20433 ( \20565 , \20563 , \20564 );
xor \U$20434 ( \20566 , \20562 , \20565 );
buf \U$20435 ( \20567 , \20566 );
buf \U$20436 ( \20568 , \20567 );
and \U$20437 ( \20569 , \20466 , \20477 );
and \U$20438 ( \20570 , \20477 , \20558 );
and \U$20439 ( \20571 , \20466 , \20558 );
or \U$20440 ( \20572 , \20569 , \20570 , \20571 );
and \U$20441 ( \20573 , \20482 , \20486 );
and \U$20442 ( \20574 , \20486 , \20557 );
and \U$20443 ( \20575 , \20482 , \20557 );
or \U$20444 ( \20576 , \20573 , \20574 , \20575 );
and \U$20445 ( \20577 , \20491 , \20495 );
and \U$20446 ( \20578 , \20495 , \20500 );
and \U$20447 ( \20579 , \20491 , \20500 );
or \U$20448 ( \20580 , \20577 , \20578 , \20579 );
and \U$20449 ( \20581 , \20505 , \20519 );
and \U$20450 ( \20582 , \20519 , \20526 );
and \U$20451 ( \20583 , \20505 , \20526 );
or \U$20452 ( \20584 , \20581 , \20582 , \20583 );
xor \U$20453 ( \20585 , \20580 , \20584 );
and \U$20454 ( \20586 , \20542 , \20555 );
xor \U$20455 ( \20587 , \20585 , \20586 );
xor \U$20456 ( \20588 , \20576 , \20587 );
and \U$20457 ( \20589 , \20470 , \20474 );
and \U$20458 ( \20590 , \20474 , \20476 );
and \U$20459 ( \20591 , \20470 , \20476 );
or \U$20460 ( \20592 , \20589 , \20590 , \20591 );
and \U$20461 ( \20593 , \20501 , \20527 );
and \U$20462 ( \20594 , \20527 , \20556 );
and \U$20463 ( \20595 , \20501 , \20556 );
or \U$20464 ( \20596 , \20593 , \20594 , \20595 );
xor \U$20465 ( \20597 , \20592 , \20596 );
and \U$20466 ( \20598 , \20509 , \20513 );
and \U$20467 ( \20599 , \20513 , \20518 );
and \U$20468 ( \20600 , \20509 , \20518 );
or \U$20469 ( \20601 , \20598 , \20599 , \20600 );
and \U$20470 ( \20602 , \20532 , \20536 );
and \U$20471 ( \20603 , \20536 , \20541 );
and \U$20472 ( \20604 , \20532 , \20541 );
or \U$20473 ( \20605 , \20602 , \20603 , \20604 );
xor \U$20474 ( \20606 , \20601 , \20605 );
and \U$20475 ( \20607 , \20545 , \20549 );
and \U$20476 ( \20608 , \20549 , \20554 );
and \U$20477 ( \20609 , \20545 , \20554 );
or \U$20478 ( \20610 , \20607 , \20608 , \20609 );
xor \U$20479 ( \20611 , \20606 , \20610 );
or \U$20480 ( \20612 , \20524 , \20525 );
and \U$20481 ( \20613 , \5674 , \10408 );
and \U$20482 ( \20614 , \6030 , \10116 );
nor \U$20483 ( \20615 , \20613 , \20614 );
xnor \U$20484 ( \20616 , \20615 , \10121 );
xor \U$20485 ( \20617 , \20612 , \20616 );
and \U$20486 ( \20618 , \5469 , \10118 );
xor \U$20487 ( \20619 , \20617 , \20618 );
xor \U$20488 ( \20620 , \20611 , \20619 );
not \U$20489 ( \20621 , \5169 );
and \U$20490 ( \20622 , \10206 , \5996 );
and \U$20491 ( \20623 , \10584 , \5695 );
nor \U$20492 ( \20624 , \20622 , \20623 );
xnor \U$20493 ( \20625 , \20624 , \5687 );
xor \U$20494 ( \20626 , \20621 , \20625 );
and \U$20495 ( \20627 , \9465 , \6401 );
and \U$20496 ( \20628 , \9897 , \6143 );
nor \U$20497 ( \20629 , \20627 , \20628 );
xnor \U$20498 ( \20630 , \20629 , \6148 );
xor \U$20499 ( \20631 , \20626 , \20630 );
and \U$20500 ( \20632 , \8835 , \7055 );
and \U$20501 ( \20633 , \9169 , \6675 );
nor \U$20502 ( \20634 , \20632 , \20633 );
xnor \U$20503 ( \20635 , \20634 , \6680 );
and \U$20504 ( \20636 , \8349 , \7489 );
and \U$20505 ( \20637 , \8652 , \7137 );
nor \U$20506 ( \20638 , \20636 , \20637 );
xnor \U$20507 ( \20639 , \20638 , \7142 );
xor \U$20508 ( \20640 , \20635 , \20639 );
and \U$20509 ( \20641 , \7700 , \8019 );
and \U$20510 ( \20642 , \8057 , \7830 );
nor \U$20511 ( \20643 , \20641 , \20642 );
xnor \U$20512 ( \20644 , \20643 , \7713 );
xor \U$20513 ( \20645 , \20640 , \20644 );
xor \U$20514 ( \20646 , \20631 , \20645 );
and \U$20515 ( \20647 , \7231 , \8540 );
and \U$20516 ( \20648 , \7556 , \8292 );
nor \U$20517 ( \20649 , \20647 , \20648 );
xnor \U$20518 ( \20650 , \20649 , \8297 );
and \U$20519 ( \20651 , \6790 , \9333 );
and \U$20520 ( \20652 , \6945 , \9006 );
nor \U$20521 ( \20653 , \20651 , \20652 );
xnor \U$20522 ( \20654 , \20653 , \8848 );
xor \U$20523 ( \20655 , \20650 , \20654 );
and \U$20524 ( \20656 , \6281 , \9765 );
and \U$20525 ( \20657 , \6514 , \9644 );
nor \U$20526 ( \20658 , \20656 , \20657 );
xnor \U$20527 ( \20659 , \20658 , \9478 );
xor \U$20528 ( \20660 , \20655 , \20659 );
xor \U$20529 ( \20661 , \20646 , \20660 );
xor \U$20530 ( \20662 , \20620 , \20661 );
xor \U$20531 ( \20663 , \20597 , \20662 );
xor \U$20532 ( \20664 , \20588 , \20663 );
xor \U$20533 ( \20665 , \20572 , \20664 );
and \U$20534 ( \20666 , \20462 , \20559 );
xor \U$20535 ( \20667 , \20665 , \20666 );
and \U$20536 ( \20668 , \20560 , \20561 );
and \U$20537 ( \20669 , \20562 , \20565 );
or \U$20538 ( \20670 , \20668 , \20669 );
xor \U$20539 ( \20671 , \20667 , \20670 );
buf \U$20540 ( \20672 , \20671 );
buf \U$20541 ( \20673 , \20672 );
and \U$20542 ( \20674 , \20576 , \20587 );
and \U$20543 ( \20675 , \20587 , \20663 );
and \U$20544 ( \20676 , \20576 , \20663 );
or \U$20545 ( \20677 , \20674 , \20675 , \20676 );
and \U$20546 ( \20678 , \20592 , \20596 );
and \U$20547 ( \20679 , \20596 , \20662 );
and \U$20548 ( \20680 , \20592 , \20662 );
or \U$20549 ( \20681 , \20678 , \20679 , \20680 );
and \U$20550 ( \20682 , \20601 , \20605 );
and \U$20551 ( \20683 , \20605 , \20610 );
and \U$20552 ( \20684 , \20601 , \20610 );
or \U$20553 ( \20685 , \20682 , \20683 , \20684 );
and \U$20554 ( \20686 , \20612 , \20616 );
and \U$20555 ( \20687 , \20616 , \20618 );
and \U$20556 ( \20688 , \20612 , \20618 );
or \U$20557 ( \20689 , \20686 , \20687 , \20688 );
xor \U$20558 ( \20690 , \20685 , \20689 );
and \U$20559 ( \20691 , \20631 , \20645 );
and \U$20560 ( \20692 , \20645 , \20660 );
and \U$20561 ( \20693 , \20631 , \20660 );
or \U$20562 ( \20694 , \20691 , \20692 , \20693 );
xor \U$20563 ( \20695 , \20690 , \20694 );
xor \U$20564 ( \20696 , \20681 , \20695 );
and \U$20565 ( \20697 , \20580 , \20584 );
and \U$20566 ( \20698 , \20584 , \20586 );
and \U$20567 ( \20699 , \20580 , \20586 );
or \U$20568 ( \20700 , \20697 , \20698 , \20699 );
and \U$20569 ( \20701 , \20611 , \20619 );
and \U$20570 ( \20702 , \20619 , \20661 );
and \U$20571 ( \20703 , \20611 , \20661 );
or \U$20572 ( \20704 , \20701 , \20702 , \20703 );
xor \U$20573 ( \20705 , \20700 , \20704 );
and \U$20574 ( \20706 , \20621 , \20625 );
and \U$20575 ( \20707 , \20625 , \20630 );
and \U$20576 ( \20708 , \20621 , \20630 );
or \U$20577 ( \20709 , \20706 , \20707 , \20708 );
and \U$20578 ( \20710 , \20635 , \20639 );
and \U$20579 ( \20711 , \20639 , \20644 );
and \U$20580 ( \20712 , \20635 , \20644 );
or \U$20581 ( \20713 , \20710 , \20711 , \20712 );
xor \U$20582 ( \20714 , \20709 , \20713 );
and \U$20583 ( \20715 , \20650 , \20654 );
and \U$20584 ( \20716 , \20654 , \20659 );
and \U$20585 ( \20717 , \20650 , \20659 );
or \U$20586 ( \20718 , \20715 , \20716 , \20717 );
xor \U$20587 ( \20719 , \20714 , \20718 );
and \U$20588 ( \20720 , \5674 , \10118 );
and \U$20589 ( \20721 , \6945 , \9333 );
and \U$20590 ( \20722 , \7231 , \9006 );
nor \U$20591 ( \20723 , \20721 , \20722 );
xnor \U$20592 ( \20724 , \20723 , \8848 );
and \U$20593 ( \20725 , \6514 , \9765 );
and \U$20594 ( \20726 , \6790 , \9644 );
nor \U$20595 ( \20727 , \20725 , \20726 );
xnor \U$20596 ( \20728 , \20727 , \9478 );
xor \U$20597 ( \20729 , \20724 , \20728 );
and \U$20598 ( \20730 , \6030 , \10408 );
and \U$20599 ( \20731 , \6281 , \10116 );
nor \U$20600 ( \20732 , \20730 , \20731 );
xnor \U$20601 ( \20733 , \20732 , \10121 );
xor \U$20602 ( \20734 , \20729 , \20733 );
xnor \U$20603 ( \20735 , \20720 , \20734 );
xor \U$20604 ( \20736 , \20719 , \20735 );
and \U$20605 ( \20737 , \8652 , \7489 );
and \U$20606 ( \20738 , \8835 , \7137 );
nor \U$20607 ( \20739 , \20737 , \20738 );
xnor \U$20608 ( \20740 , \20739 , \7142 );
and \U$20609 ( \20741 , \8057 , \8019 );
and \U$20610 ( \20742 , \8349 , \7830 );
nor \U$20611 ( \20743 , \20741 , \20742 );
xnor \U$20612 ( \20744 , \20743 , \7713 );
xor \U$20613 ( \20745 , \20740 , \20744 );
and \U$20614 ( \20746 , \7556 , \8540 );
and \U$20615 ( \20747 , \7700 , \8292 );
nor \U$20616 ( \20748 , \20746 , \20747 );
xnor \U$20617 ( \20749 , \20748 , \8297 );
xor \U$20618 ( \20750 , \20745 , \20749 );
and \U$20619 ( \20751 , \10584 , \5996 );
not \U$20620 ( \20752 , \20751 );
xnor \U$20621 ( \20753 , \20752 , \5687 );
and \U$20622 ( \20754 , \9897 , \6401 );
and \U$20623 ( \20755 , \10206 , \6143 );
nor \U$20624 ( \20756 , \20754 , \20755 );
xnor \U$20625 ( \20757 , \20756 , \6148 );
xor \U$20626 ( \20758 , \20753 , \20757 );
and \U$20627 ( \20759 , \9169 , \7055 );
and \U$20628 ( \20760 , \9465 , \6675 );
nor \U$20629 ( \20761 , \20759 , \20760 );
xnor \U$20630 ( \20762 , \20761 , \6680 );
xor \U$20631 ( \20763 , \20758 , \20762 );
xor \U$20632 ( \20764 , \20750 , \20763 );
xor \U$20633 ( \20765 , \20736 , \20764 );
xor \U$20634 ( \20766 , \20705 , \20765 );
xor \U$20635 ( \20767 , \20696 , \20766 );
xor \U$20636 ( \20768 , \20677 , \20767 );
and \U$20637 ( \20769 , \20572 , \20664 );
xor \U$20638 ( \20770 , \20768 , \20769 );
and \U$20639 ( \20771 , \20665 , \20666 );
and \U$20640 ( \20772 , \20667 , \20670 );
or \U$20641 ( \20773 , \20771 , \20772 );
xor \U$20642 ( \20774 , \20770 , \20773 );
buf \U$20643 ( \20775 , \20774 );
buf \U$20644 ( \20776 , \20775 );
and \U$20645 ( \20777 , \20681 , \20695 );
and \U$20646 ( \20778 , \20695 , \20766 );
and \U$20647 ( \20779 , \20681 , \20766 );
or \U$20648 ( \20780 , \20777 , \20778 , \20779 );
and \U$20649 ( \20781 , \20700 , \20704 );
and \U$20650 ( \20782 , \20704 , \20765 );
and \U$20651 ( \20783 , \20700 , \20765 );
or \U$20652 ( \20784 , \20781 , \20782 , \20783 );
and \U$20653 ( \20785 , \20709 , \20713 );
and \U$20654 ( \20786 , \20713 , \20718 );
and \U$20655 ( \20787 , \20709 , \20718 );
or \U$20656 ( \20788 , \20785 , \20786 , \20787 );
or \U$20657 ( \20789 , \20720 , \20734 );
xor \U$20658 ( \20790 , \20788 , \20789 );
and \U$20659 ( \20791 , \20750 , \20763 );
xor \U$20660 ( \20792 , \20790 , \20791 );
xor \U$20661 ( \20793 , \20784 , \20792 );
and \U$20662 ( \20794 , \20685 , \20689 );
and \U$20663 ( \20795 , \20689 , \20694 );
and \U$20664 ( \20796 , \20685 , \20694 );
or \U$20665 ( \20797 , \20794 , \20795 , \20796 );
and \U$20666 ( \20798 , \20719 , \20735 );
and \U$20667 ( \20799 , \20735 , \20764 );
and \U$20668 ( \20800 , \20719 , \20764 );
or \U$20669 ( \20801 , \20798 , \20799 , \20800 );
xor \U$20670 ( \20802 , \20797 , \20801 );
not \U$20671 ( \20803 , \5687 );
and \U$20672 ( \20804 , \10206 , \6401 );
and \U$20673 ( \20805 , \10584 , \6143 );
nor \U$20674 ( \20806 , \20804 , \20805 );
xnor \U$20675 ( \20807 , \20806 , \6148 );
xor \U$20676 ( \20808 , \20803 , \20807 );
and \U$20677 ( \20809 , \9465 , \7055 );
and \U$20678 ( \20810 , \9897 , \6675 );
nor \U$20679 ( \20811 , \20809 , \20810 );
xnor \U$20680 ( \20812 , \20811 , \6680 );
xor \U$20681 ( \20813 , \20808 , \20812 );
and \U$20682 ( \20814 , \20740 , \20744 );
and \U$20683 ( \20815 , \20744 , \20749 );
and \U$20684 ( \20816 , \20740 , \20749 );
or \U$20685 ( \20817 , \20814 , \20815 , \20816 );
and \U$20686 ( \20818 , \20753 , \20757 );
and \U$20687 ( \20819 , \20757 , \20762 );
and \U$20688 ( \20820 , \20753 , \20762 );
or \U$20689 ( \20821 , \20818 , \20819 , \20820 );
xor \U$20690 ( \20822 , \20817 , \20821 );
and \U$20691 ( \20823 , \20724 , \20728 );
and \U$20692 ( \20824 , \20728 , \20733 );
and \U$20693 ( \20825 , \20724 , \20733 );
or \U$20694 ( \20826 , \20823 , \20824 , \20825 );
xor \U$20695 ( \20827 , \20822 , \20826 );
xor \U$20696 ( \20828 , \20813 , \20827 );
and \U$20697 ( \20829 , \6030 , \10118 );
and \U$20698 ( \20830 , \8835 , \7489 );
and \U$20699 ( \20831 , \9169 , \7137 );
nor \U$20700 ( \20832 , \20830 , \20831 );
xnor \U$20701 ( \20833 , \20832 , \7142 );
and \U$20702 ( \20834 , \8349 , \8019 );
and \U$20703 ( \20835 , \8652 , \7830 );
nor \U$20704 ( \20836 , \20834 , \20835 );
xnor \U$20705 ( \20837 , \20836 , \7713 );
xor \U$20706 ( \20838 , \20833 , \20837 );
and \U$20707 ( \20839 , \7700 , \8540 );
and \U$20708 ( \20840 , \8057 , \8292 );
nor \U$20709 ( \20841 , \20839 , \20840 );
xnor \U$20710 ( \20842 , \20841 , \8297 );
xor \U$20711 ( \20843 , \20838 , \20842 );
xor \U$20712 ( \20844 , \20829 , \20843 );
and \U$20713 ( \20845 , \7231 , \9333 );
and \U$20714 ( \20846 , \7556 , \9006 );
nor \U$20715 ( \20847 , \20845 , \20846 );
xnor \U$20716 ( \20848 , \20847 , \8848 );
and \U$20717 ( \20849 , \6790 , \9765 );
and \U$20718 ( \20850 , \6945 , \9644 );
nor \U$20719 ( \20851 , \20849 , \20850 );
xnor \U$20720 ( \20852 , \20851 , \9478 );
xor \U$20721 ( \20853 , \20848 , \20852 );
and \U$20722 ( \20854 , \6281 , \10408 );
and \U$20723 ( \20855 , \6514 , \10116 );
nor \U$20724 ( \20856 , \20854 , \20855 );
xnor \U$20725 ( \20857 , \20856 , \10121 );
xor \U$20726 ( \20858 , \20853 , \20857 );
xor \U$20727 ( \20859 , \20844 , \20858 );
xor \U$20728 ( \20860 , \20828 , \20859 );
xor \U$20729 ( \20861 , \20802 , \20860 );
xor \U$20730 ( \20862 , \20793 , \20861 );
xor \U$20731 ( \20863 , \20780 , \20862 );
and \U$20732 ( \20864 , \20677 , \20767 );
xor \U$20733 ( \20865 , \20863 , \20864 );
and \U$20734 ( \20866 , \20768 , \20769 );
and \U$20735 ( \20867 , \20770 , \20773 );
or \U$20736 ( \20868 , \20866 , \20867 );
xor \U$20737 ( \20869 , \20865 , \20868 );
buf \U$20738 ( \20870 , \20869 );
buf \U$20739 ( \20871 , \20870 );
and \U$20740 ( \20872 , \20784 , \20792 );
and \U$20741 ( \20873 , \20792 , \20861 );
and \U$20742 ( \20874 , \20784 , \20861 );
or \U$20743 ( \20875 , \20872 , \20873 , \20874 );
and \U$20744 ( \20876 , \20797 , \20801 );
and \U$20745 ( \20877 , \20801 , \20860 );
and \U$20746 ( \20878 , \20797 , \20860 );
or \U$20747 ( \20879 , \20876 , \20877 , \20878 );
and \U$20748 ( \20880 , \20788 , \20789 );
and \U$20749 ( \20881 , \20789 , \20791 );
and \U$20750 ( \20882 , \20788 , \20791 );
or \U$20751 ( \20883 , \20880 , \20881 , \20882 );
and \U$20752 ( \20884 , \20813 , \20827 );
and \U$20753 ( \20885 , \20827 , \20859 );
and \U$20754 ( \20886 , \20813 , \20859 );
or \U$20755 ( \20887 , \20884 , \20885 , \20886 );
xor \U$20756 ( \20888 , \20883 , \20887 );
and \U$20757 ( \20889 , \6945 , \9765 );
and \U$20758 ( \20890 , \7231 , \9644 );
nor \U$20759 ( \20891 , \20889 , \20890 );
xnor \U$20760 ( \20892 , \20891 , \9478 );
and \U$20761 ( \20893 , \6514 , \10408 );
and \U$20762 ( \20894 , \6790 , \10116 );
nor \U$20763 ( \20895 , \20893 , \20894 );
xnor \U$20764 ( \20896 , \20895 , \10121 );
xor \U$20765 ( \20897 , \20892 , \20896 );
and \U$20766 ( \20898 , \6281 , \10118 );
xor \U$20767 ( \20899 , \20897 , \20898 );
and \U$20768 ( \20900 , \8652 , \8019 );
and \U$20769 ( \20901 , \8835 , \7830 );
nor \U$20770 ( \20902 , \20900 , \20901 );
xnor \U$20771 ( \20903 , \20902 , \7713 );
and \U$20772 ( \20904 , \8057 , \8540 );
and \U$20773 ( \20905 , \8349 , \8292 );
nor \U$20774 ( \20906 , \20904 , \20905 );
xnor \U$20775 ( \20907 , \20906 , \8297 );
xor \U$20776 ( \20908 , \20903 , \20907 );
and \U$20777 ( \20909 , \7556 , \9333 );
and \U$20778 ( \20910 , \7700 , \9006 );
nor \U$20779 ( \20911 , \20909 , \20910 );
xnor \U$20780 ( \20912 , \20911 , \8848 );
xor \U$20781 ( \20913 , \20908 , \20912 );
xnor \U$20782 ( \20914 , \20899 , \20913 );
xor \U$20783 ( \20915 , \20888 , \20914 );
xor \U$20784 ( \20916 , \20879 , \20915 );
and \U$20785 ( \20917 , \20833 , \20837 );
and \U$20786 ( \20918 , \20837 , \20842 );
and \U$20787 ( \20919 , \20833 , \20842 );
or \U$20788 ( \20920 , \20917 , \20918 , \20919 );
and \U$20789 ( \20921 , \20803 , \20807 );
and \U$20790 ( \20922 , \20807 , \20812 );
and \U$20791 ( \20923 , \20803 , \20812 );
or \U$20792 ( \20924 , \20921 , \20922 , \20923 );
xor \U$20793 ( \20925 , \20920 , \20924 );
and \U$20794 ( \20926 , \20848 , \20852 );
and \U$20795 ( \20927 , \20852 , \20857 );
and \U$20796 ( \20928 , \20848 , \20857 );
or \U$20797 ( \20929 , \20926 , \20927 , \20928 );
xor \U$20798 ( \20930 , \20925 , \20929 );
and \U$20799 ( \20931 , \20817 , \20821 );
and \U$20800 ( \20932 , \20821 , \20826 );
and \U$20801 ( \20933 , \20817 , \20826 );
or \U$20802 ( \20934 , \20931 , \20932 , \20933 );
and \U$20803 ( \20935 , \20829 , \20843 );
and \U$20804 ( \20936 , \20843 , \20858 );
and \U$20805 ( \20937 , \20829 , \20858 );
or \U$20806 ( \20938 , \20935 , \20936 , \20937 );
xor \U$20807 ( \20939 , \20934 , \20938 );
and \U$20808 ( \20940 , \10584 , \6401 );
not \U$20809 ( \20941 , \20940 );
xnor \U$20810 ( \20942 , \20941 , \6148 );
and \U$20811 ( \20943 , \9897 , \7055 );
and \U$20812 ( \20944 , \10206 , \6675 );
nor \U$20813 ( \20945 , \20943 , \20944 );
xnor \U$20814 ( \20946 , \20945 , \6680 );
xor \U$20815 ( \20947 , \20942 , \20946 );
and \U$20816 ( \20948 , \9169 , \7489 );
and \U$20817 ( \20949 , \9465 , \7137 );
nor \U$20818 ( \20950 , \20948 , \20949 );
xnor \U$20819 ( \20951 , \20950 , \7142 );
xor \U$20820 ( \20952 , \20947 , \20951 );
xor \U$20821 ( \20953 , \20939 , \20952 );
xor \U$20822 ( \20954 , \20930 , \20953 );
xor \U$20823 ( \20955 , \20916 , \20954 );
xor \U$20824 ( \20956 , \20875 , \20955 );
and \U$20825 ( \20957 , \20780 , \20862 );
xor \U$20826 ( \20958 , \20956 , \20957 );
and \U$20827 ( \20959 , \20863 , \20864 );
and \U$20828 ( \20960 , \20865 , \20868 );
or \U$20829 ( \20961 , \20959 , \20960 );
xor \U$20830 ( \20962 , \20958 , \20961 );
buf \U$20831 ( \20963 , \20962 );
buf \U$20832 ( \20964 , \20963 );
and \U$20833 ( \20965 , \20879 , \20915 );
and \U$20834 ( \20966 , \20915 , \20954 );
and \U$20835 ( \20967 , \20879 , \20954 );
or \U$20836 ( \20968 , \20965 , \20966 , \20967 );
and \U$20837 ( \20969 , \20883 , \20887 );
and \U$20838 ( \20970 , \20887 , \20914 );
and \U$20839 ( \20971 , \20883 , \20914 );
or \U$20840 ( \20972 , \20969 , \20970 , \20971 );
and \U$20841 ( \20973 , \20930 , \20953 );
xor \U$20842 ( \20974 , \20972 , \20973 );
and \U$20843 ( \20975 , \20934 , \20938 );
and \U$20844 ( \20976 , \20938 , \20952 );
and \U$20845 ( \20977 , \20934 , \20952 );
or \U$20846 ( \20978 , \20975 , \20976 , \20977 );
and \U$20847 ( \20979 , \20892 , \20896 );
and \U$20848 ( \20980 , \20896 , \20898 );
and \U$20849 ( \20981 , \20892 , \20898 );
or \U$20850 ( \20982 , \20979 , \20980 , \20981 );
and \U$20851 ( \20983 , \20942 , \20946 );
and \U$20852 ( \20984 , \20946 , \20951 );
and \U$20853 ( \20985 , \20942 , \20951 );
or \U$20854 ( \20986 , \20983 , \20984 , \20985 );
xor \U$20855 ( \20987 , \20982 , \20986 );
and \U$20856 ( \20988 , \20903 , \20907 );
and \U$20857 ( \20989 , \20907 , \20912 );
and \U$20858 ( \20990 , \20903 , \20912 );
or \U$20859 ( \20991 , \20988 , \20989 , \20990 );
xor \U$20860 ( \20992 , \20987 , \20991 );
xor \U$20861 ( \20993 , \20978 , \20992 );
and \U$20862 ( \20994 , \20920 , \20924 );
and \U$20863 ( \20995 , \20924 , \20929 );
and \U$20864 ( \20996 , \20920 , \20929 );
or \U$20865 ( \20997 , \20994 , \20995 , \20996 );
or \U$20866 ( \20998 , \20899 , \20913 );
xor \U$20867 ( \20999 , \20997 , \20998 );
not \U$20868 ( \21000 , \6148 );
and \U$20869 ( \21001 , \10206 , \7055 );
and \U$20870 ( \21002 , \10584 , \6675 );
nor \U$20871 ( \21003 , \21001 , \21002 );
xnor \U$20872 ( \21004 , \21003 , \6680 );
xor \U$20873 ( \21005 , \21000 , \21004 );
and \U$20874 ( \21006 , \9465 , \7489 );
and \U$20875 ( \21007 , \9897 , \7137 );
nor \U$20876 ( \21008 , \21006 , \21007 );
xnor \U$20877 ( \21009 , \21008 , \7142 );
xor \U$20878 ( \21010 , \21005 , \21009 );
and \U$20879 ( \21011 , \7231 , \9765 );
and \U$20880 ( \21012 , \7556 , \9644 );
nor \U$20881 ( \21013 , \21011 , \21012 );
xnor \U$20882 ( \21014 , \21013 , \9478 );
and \U$20883 ( \21015 , \6790 , \10408 );
and \U$20884 ( \21016 , \6945 , \10116 );
nor \U$20885 ( \21017 , \21015 , \21016 );
xnor \U$20886 ( \21018 , \21017 , \10121 );
xor \U$20887 ( \21019 , \21014 , \21018 );
and \U$20888 ( \21020 , \6514 , \10118 );
xor \U$20889 ( \21021 , \21019 , \21020 );
xor \U$20890 ( \21022 , \21010 , \21021 );
and \U$20891 ( \21023 , \8835 , \8019 );
and \U$20892 ( \21024 , \9169 , \7830 );
nor \U$20893 ( \21025 , \21023 , \21024 );
xnor \U$20894 ( \21026 , \21025 , \7713 );
and \U$20895 ( \21027 , \8349 , \8540 );
and \U$20896 ( \21028 , \8652 , \8292 );
nor \U$20897 ( \21029 , \21027 , \21028 );
xnor \U$20898 ( \21030 , \21029 , \8297 );
xor \U$20899 ( \21031 , \21026 , \21030 );
and \U$20900 ( \21032 , \7700 , \9333 );
and \U$20901 ( \21033 , \8057 , \9006 );
nor \U$20902 ( \21034 , \21032 , \21033 );
xnor \U$20903 ( \21035 , \21034 , \8848 );
xor \U$20904 ( \21036 , \21031 , \21035 );
xor \U$20905 ( \21037 , \21022 , \21036 );
xor \U$20906 ( \21038 , \20999 , \21037 );
xor \U$20907 ( \21039 , \20993 , \21038 );
xor \U$20908 ( \21040 , \20974 , \21039 );
xor \U$20909 ( \21041 , \20968 , \21040 );
and \U$20910 ( \21042 , \20875 , \20955 );
xor \U$20911 ( \21043 , \21041 , \21042 );
and \U$20912 ( \21044 , \20956 , \20957 );
and \U$20913 ( \21045 , \20958 , \20961 );
or \U$20914 ( \21046 , \21044 , \21045 );
xor \U$20915 ( \21047 , \21043 , \21046 );
buf \U$20916 ( \21048 , \21047 );
buf \U$20917 ( \21049 , \21048 );
and \U$20918 ( \21050 , \20978 , \20992 );
and \U$20919 ( \21051 , \20992 , \21038 );
and \U$20920 ( \21052 , \20978 , \21038 );
or \U$20921 ( \21053 , \21050 , \21051 , \21052 );
and \U$20922 ( \21054 , \20972 , \20973 );
and \U$20923 ( \21055 , \20973 , \21039 );
and \U$20924 ( \21056 , \20972 , \21039 );
or \U$20925 ( \21057 , \21054 , \21055 , \21056 );
xor \U$20926 ( \21058 , \21053 , \21057 );
and \U$20927 ( \21059 , \20997 , \20998 );
and \U$20928 ( \21060 , \20998 , \21037 );
and \U$20929 ( \21061 , \20997 , \21037 );
or \U$20930 ( \21062 , \21059 , \21060 , \21061 );
and \U$20931 ( \21063 , \21000 , \21004 );
and \U$20932 ( \21064 , \21004 , \21009 );
and \U$20933 ( \21065 , \21000 , \21009 );
or \U$20934 ( \21066 , \21063 , \21064 , \21065 );
and \U$20935 ( \21067 , \21014 , \21018 );
and \U$20936 ( \21068 , \21018 , \21020 );
and \U$20937 ( \21069 , \21014 , \21020 );
or \U$20938 ( \21070 , \21067 , \21068 , \21069 );
xor \U$20939 ( \21071 , \21066 , \21070 );
and \U$20940 ( \21072 , \21026 , \21030 );
and \U$20941 ( \21073 , \21030 , \21035 );
and \U$20942 ( \21074 , \21026 , \21035 );
or \U$20943 ( \21075 , \21072 , \21073 , \21074 );
xor \U$20944 ( \21076 , \21071 , \21075 );
xor \U$20945 ( \21077 , \21062 , \21076 );
and \U$20946 ( \21078 , \20982 , \20986 );
and \U$20947 ( \21079 , \20986 , \20991 );
and \U$20948 ( \21080 , \20982 , \20991 );
or \U$20949 ( \21081 , \21078 , \21079 , \21080 );
and \U$20950 ( \21082 , \21010 , \21021 );
and \U$20951 ( \21083 , \21021 , \21036 );
and \U$20952 ( \21084 , \21010 , \21036 );
or \U$20953 ( \21085 , \21082 , \21083 , \21084 );
xor \U$20954 ( \21086 , \21081 , \21085 );
and \U$20955 ( \21087 , \10584 , \7055 );
not \U$20956 ( \21088 , \21087 );
xnor \U$20957 ( \21089 , \21088 , \6680 );
and \U$20958 ( \21090 , \9897 , \7489 );
and \U$20959 ( \21091 , \10206 , \7137 );
nor \U$20960 ( \21092 , \21090 , \21091 );
xnor \U$20961 ( \21093 , \21092 , \7142 );
xor \U$20962 ( \21094 , \21089 , \21093 );
and \U$20963 ( \21095 , \9169 , \8019 );
and \U$20964 ( \21096 , \9465 , \7830 );
nor \U$20965 ( \21097 , \21095 , \21096 );
xnor \U$20966 ( \21098 , \21097 , \7713 );
xor \U$20967 ( \21099 , \21094 , \21098 );
and \U$20968 ( \21100 , \8652 , \8540 );
and \U$20969 ( \21101 , \8835 , \8292 );
nor \U$20970 ( \21102 , \21100 , \21101 );
xnor \U$20971 ( \21103 , \21102 , \8297 );
and \U$20972 ( \21104 , \8057 , \9333 );
and \U$20973 ( \21105 , \8349 , \9006 );
nor \U$20974 ( \21106 , \21104 , \21105 );
xnor \U$20975 ( \21107 , \21106 , \8848 );
xor \U$20976 ( \21108 , \21103 , \21107 );
and \U$20977 ( \21109 , \7556 , \9765 );
and \U$20978 ( \21110 , \7700 , \9644 );
nor \U$20979 ( \21111 , \21109 , \21110 );
xnor \U$20980 ( \21112 , \21111 , \9478 );
xor \U$20981 ( \21113 , \21108 , \21112 );
xor \U$20982 ( \21114 , \21099 , \21113 );
and \U$20983 ( \21115 , \6945 , \10408 );
and \U$20984 ( \21116 , \7231 , \10116 );
nor \U$20985 ( \21117 , \21115 , \21116 );
xnor \U$20986 ( \21118 , \21117 , \10121 );
and \U$20987 ( \21119 , \6790 , \10118 );
xnor \U$20988 ( \21120 , \21118 , \21119 );
xor \U$20989 ( \21121 , \21114 , \21120 );
xor \U$20990 ( \21122 , \21086 , \21121 );
xor \U$20991 ( \21123 , \21077 , \21122 );
xor \U$20992 ( \21124 , \21058 , \21123 );
and \U$20993 ( \21125 , \20968 , \21040 );
xor \U$20994 ( \21126 , \21124 , \21125 );
and \U$20995 ( \21127 , \21041 , \21042 );
and \U$20996 ( \21128 , \21043 , \21046 );
or \U$20997 ( \21129 , \21127 , \21128 );
xor \U$20998 ( \21130 , \21126 , \21129 );
buf \U$20999 ( \21131 , \21130 );
buf \U$21000 ( \21132 , \21131 );
and \U$21001 ( \21133 , \21062 , \21076 );
and \U$21002 ( \21134 , \21076 , \21122 );
and \U$21003 ( \21135 , \21062 , \21122 );
or \U$21004 ( \21136 , \21133 , \21134 , \21135 );
and \U$21005 ( \21137 , \21081 , \21085 );
and \U$21006 ( \21138 , \21085 , \21121 );
and \U$21007 ( \21139 , \21081 , \21121 );
or \U$21008 ( \21140 , \21137 , \21138 , \21139 );
and \U$21009 ( \21141 , \21089 , \21093 );
and \U$21010 ( \21142 , \21093 , \21098 );
and \U$21011 ( \21143 , \21089 , \21098 );
or \U$21012 ( \21144 , \21141 , \21142 , \21143 );
and \U$21013 ( \21145 , \21103 , \21107 );
and \U$21014 ( \21146 , \21107 , \21112 );
and \U$21015 ( \21147 , \21103 , \21112 );
or \U$21016 ( \21148 , \21145 , \21146 , \21147 );
xor \U$21017 ( \21149 , \21144 , \21148 );
or \U$21018 ( \21150 , \21118 , \21119 );
xor \U$21019 ( \21151 , \21149 , \21150 );
xor \U$21020 ( \21152 , \21140 , \21151 );
and \U$21021 ( \21153 , \21066 , \21070 );
and \U$21022 ( \21154 , \21070 , \21075 );
and \U$21023 ( \21155 , \21066 , \21075 );
or \U$21024 ( \21156 , \21153 , \21154 , \21155 );
and \U$21025 ( \21157 , \21099 , \21113 );
and \U$21026 ( \21158 , \21113 , \21120 );
and \U$21027 ( \21159 , \21099 , \21120 );
or \U$21028 ( \21160 , \21157 , \21158 , \21159 );
xor \U$21029 ( \21161 , \21156 , \21160 );
not \U$21030 ( \21162 , \6680 );
and \U$21031 ( \21163 , \10206 , \7489 );
and \U$21032 ( \21164 , \10584 , \7137 );
nor \U$21033 ( \21165 , \21163 , \21164 );
xnor \U$21034 ( \21166 , \21165 , \7142 );
xor \U$21035 ( \21167 , \21162 , \21166 );
and \U$21036 ( \21168 , \9465 , \8019 );
and \U$21037 ( \21169 , \9897 , \7830 );
nor \U$21038 ( \21170 , \21168 , \21169 );
xnor \U$21039 ( \21171 , \21170 , \7713 );
xor \U$21040 ( \21172 , \21167 , \21171 );
and \U$21041 ( \21173 , \8835 , \8540 );
and \U$21042 ( \21174 , \9169 , \8292 );
nor \U$21043 ( \21175 , \21173 , \21174 );
xnor \U$21044 ( \21176 , \21175 , \8297 );
and \U$21045 ( \21177 , \8349 , \9333 );
and \U$21046 ( \21178 , \8652 , \9006 );
nor \U$21047 ( \21179 , \21177 , \21178 );
xnor \U$21048 ( \21180 , \21179 , \8848 );
xor \U$21049 ( \21181 , \21176 , \21180 );
and \U$21050 ( \21182 , \7700 , \9765 );
and \U$21051 ( \21183 , \8057 , \9644 );
nor \U$21052 ( \21184 , \21182 , \21183 );
xnor \U$21053 ( \21185 , \21184 , \9478 );
xor \U$21054 ( \21186 , \21181 , \21185 );
xor \U$21055 ( \21187 , \21172 , \21186 );
and \U$21056 ( \21188 , \7231 , \10408 );
and \U$21057 ( \21189 , \7556 , \10116 );
nor \U$21058 ( \21190 , \21188 , \21189 );
xnor \U$21059 ( \21191 , \21190 , \10121 );
and \U$21060 ( \21192 , \6945 , \10118 );
xor \U$21061 ( \21193 , \21191 , \21192 );
xor \U$21062 ( \21194 , \21187 , \21193 );
xor \U$21063 ( \21195 , \21161 , \21194 );
xor \U$21064 ( \21196 , \21152 , \21195 );
xor \U$21065 ( \21197 , \21136 , \21196 );
and \U$21066 ( \21198 , \21053 , \21057 );
and \U$21067 ( \21199 , \21057 , \21123 );
and \U$21068 ( \21200 , \21053 , \21123 );
or \U$21069 ( \21201 , \21198 , \21199 , \21200 );
xor \U$21070 ( \21202 , \21197 , \21201 );
and \U$21071 ( \21203 , \21124 , \21125 );
and \U$21072 ( \21204 , \21126 , \21129 );
or \U$21073 ( \21205 , \21203 , \21204 );
xor \U$21074 ( \21206 , \21202 , \21205 );
buf \U$21075 ( \21207 , \21206 );
buf \U$21076 ( \21208 , \21207 );
and \U$21077 ( \21209 , \21140 , \21151 );
and \U$21078 ( \21210 , \21151 , \21195 );
and \U$21079 ( \21211 , \21140 , \21195 );
or \U$21080 ( \21212 , \21209 , \21210 , \21211 );
and \U$21081 ( \21213 , \21156 , \21160 );
and \U$21082 ( \21214 , \21160 , \21194 );
and \U$21083 ( \21215 , \21156 , \21194 );
or \U$21084 ( \21216 , \21213 , \21214 , \21215 );
and \U$21085 ( \21217 , \21162 , \21166 );
and \U$21086 ( \21218 , \21166 , \21171 );
and \U$21087 ( \21219 , \21162 , \21171 );
or \U$21088 ( \21220 , \21217 , \21218 , \21219 );
and \U$21089 ( \21221 , \21176 , \21180 );
and \U$21090 ( \21222 , \21180 , \21185 );
and \U$21091 ( \21223 , \21176 , \21185 );
or \U$21092 ( \21224 , \21221 , \21222 , \21223 );
xor \U$21093 ( \21225 , \21220 , \21224 );
and \U$21094 ( \21226 , \21191 , \21192 );
xor \U$21095 ( \21227 , \21225 , \21226 );
xor \U$21096 ( \21228 , \21216 , \21227 );
and \U$21097 ( \21229 , \21144 , \21148 );
and \U$21098 ( \21230 , \21148 , \21150 );
and \U$21099 ( \21231 , \21144 , \21150 );
or \U$21100 ( \21232 , \21229 , \21230 , \21231 );
and \U$21101 ( \21233 , \21172 , \21186 );
and \U$21102 ( \21234 , \21186 , \21193 );
and \U$21103 ( \21235 , \21172 , \21193 );
or \U$21104 ( \21236 , \21233 , \21234 , \21235 );
xor \U$21105 ( \21237 , \21232 , \21236 );
and \U$21106 ( \21238 , \8652 , \9333 );
and \U$21107 ( \21239 , \8835 , \9006 );
nor \U$21108 ( \21240 , \21238 , \21239 );
xnor \U$21109 ( \21241 , \21240 , \8848 );
and \U$21110 ( \21242 , \8057 , \9765 );
and \U$21111 ( \21243 , \8349 , \9644 );
nor \U$21112 ( \21244 , \21242 , \21243 );
xnor \U$21113 ( \21245 , \21244 , \9478 );
xor \U$21114 ( \21246 , \21241 , \21245 );
and \U$21115 ( \21247 , \7556 , \10408 );
and \U$21116 ( \21248 , \7700 , \10116 );
nor \U$21117 ( \21249 , \21247 , \21248 );
xnor \U$21118 ( \21250 , \21249 , \10121 );
xor \U$21119 ( \21251 , \21246 , \21250 );
and \U$21120 ( \21252 , \10584 , \7489 );
not \U$21121 ( \21253 , \21252 );
xnor \U$21122 ( \21254 , \21253 , \7142 );
and \U$21123 ( \21255 , \9897 , \8019 );
and \U$21124 ( \21256 , \10206 , \7830 );
nor \U$21125 ( \21257 , \21255 , \21256 );
xnor \U$21126 ( \21258 , \21257 , \7713 );
xor \U$21127 ( \21259 , \21254 , \21258 );
and \U$21128 ( \21260 , \9169 , \8540 );
and \U$21129 ( \21261 , \9465 , \8292 );
nor \U$21130 ( \21262 , \21260 , \21261 );
xnor \U$21131 ( \21263 , \21262 , \8297 );
xor \U$21132 ( \21264 , \21259 , \21263 );
xor \U$21133 ( \21265 , \21251 , \21264 );
and \U$21134 ( \21266 , \7231 , \10118 );
not \U$21135 ( \21267 , \21266 );
xor \U$21136 ( \21268 , \21265 , \21267 );
xor \U$21137 ( \21269 , \21237 , \21268 );
xor \U$21138 ( \21270 , \21228 , \21269 );
xor \U$21139 ( \21271 , \21212 , \21270 );
and \U$21140 ( \21272 , \21136 , \21196 );
xor \U$21141 ( \21273 , \21271 , \21272 );
and \U$21142 ( \21274 , \21197 , \21201 );
and \U$21143 ( \21275 , \21202 , \21205 );
or \U$21144 ( \21276 , \21274 , \21275 );
xor \U$21145 ( \21277 , \21273 , \21276 );
buf \U$21146 ( \21278 , \21277 );
buf \U$21147 ( \21279 , \21278 );
and \U$21148 ( \21280 , \21216 , \21227 );
and \U$21149 ( \21281 , \21227 , \21269 );
and \U$21150 ( \21282 , \21216 , \21269 );
or \U$21151 ( \21283 , \21280 , \21281 , \21282 );
and \U$21152 ( \21284 , \21232 , \21236 );
and \U$21153 ( \21285 , \21236 , \21268 );
and \U$21154 ( \21286 , \21232 , \21268 );
or \U$21155 ( \21287 , \21284 , \21285 , \21286 );
and \U$21156 ( \21288 , \21241 , \21245 );
and \U$21157 ( \21289 , \21245 , \21250 );
and \U$21158 ( \21290 , \21241 , \21250 );
or \U$21159 ( \21291 , \21288 , \21289 , \21290 );
and \U$21160 ( \21292 , \21254 , \21258 );
and \U$21161 ( \21293 , \21258 , \21263 );
and \U$21162 ( \21294 , \21254 , \21263 );
or \U$21163 ( \21295 , \21292 , \21293 , \21294 );
xor \U$21164 ( \21296 , \21291 , \21295 );
buf \U$21165 ( \21297 , \21266 );
xor \U$21166 ( \21298 , \21296 , \21297 );
xor \U$21167 ( \21299 , \21287 , \21298 );
and \U$21168 ( \21300 , \21220 , \21224 );
and \U$21169 ( \21301 , \21224 , \21226 );
and \U$21170 ( \21302 , \21220 , \21226 );
or \U$21171 ( \21303 , \21300 , \21301 , \21302 );
and \U$21172 ( \21304 , \21251 , \21264 );
and \U$21173 ( \21305 , \21264 , \21267 );
and \U$21174 ( \21306 , \21251 , \21267 );
or \U$21175 ( \21307 , \21304 , \21305 , \21306 );
xor \U$21176 ( \21308 , \21303 , \21307 );
and \U$21177 ( \21309 , \7556 , \10118 );
and \U$21178 ( \21310 , \8835 , \9333 );
and \U$21179 ( \21311 , \9169 , \9006 );
nor \U$21180 ( \21312 , \21310 , \21311 );
xnor \U$21181 ( \21313 , \21312 , \8848 );
and \U$21182 ( \21314 , \8349 , \9765 );
and \U$21183 ( \21315 , \8652 , \9644 );
nor \U$21184 ( \21316 , \21314 , \21315 );
xnor \U$21185 ( \21317 , \21316 , \9478 );
xor \U$21186 ( \21318 , \21313 , \21317 );
and \U$21187 ( \21319 , \7700 , \10408 );
and \U$21188 ( \21320 , \8057 , \10116 );
nor \U$21189 ( \21321 , \21319 , \21320 );
xnor \U$21190 ( \21322 , \21321 , \10121 );
xor \U$21191 ( \21323 , \21318 , \21322 );
xor \U$21192 ( \21324 , \21309 , \21323 );
not \U$21193 ( \21325 , \7142 );
and \U$21194 ( \21326 , \10206 , \8019 );
and \U$21195 ( \21327 , \10584 , \7830 );
nor \U$21196 ( \21328 , \21326 , \21327 );
xnor \U$21197 ( \21329 , \21328 , \7713 );
xor \U$21198 ( \21330 , \21325 , \21329 );
and \U$21199 ( \21331 , \9465 , \8540 );
and \U$21200 ( \21332 , \9897 , \8292 );
nor \U$21201 ( \21333 , \21331 , \21332 );
xnor \U$21202 ( \21334 , \21333 , \8297 );
xor \U$21203 ( \21335 , \21330 , \21334 );
xor \U$21204 ( \21336 , \21324 , \21335 );
xor \U$21205 ( \21337 , \21308 , \21336 );
xor \U$21206 ( \21338 , \21299 , \21337 );
xor \U$21207 ( \21339 , \21283 , \21338 );
and \U$21208 ( \21340 , \21212 , \21270 );
xor \U$21209 ( \21341 , \21339 , \21340 );
and \U$21210 ( \21342 , \21271 , \21272 );
and \U$21211 ( \21343 , \21273 , \21276 );
or \U$21212 ( \21344 , \21342 , \21343 );
xor \U$21213 ( \21345 , \21341 , \21344 );
buf \U$21214 ( \21346 , \21345 );
buf \U$21215 ( \21347 , \21346 );
and \U$21216 ( \21348 , \21287 , \21298 );
and \U$21217 ( \21349 , \21298 , \21337 );
and \U$21218 ( \21350 , \21287 , \21337 );
or \U$21219 ( \21351 , \21348 , \21349 , \21350 );
and \U$21220 ( \21352 , \21303 , \21307 );
and \U$21221 ( \21353 , \21307 , \21336 );
and \U$21222 ( \21354 , \21303 , \21336 );
or \U$21223 ( \21355 , \21352 , \21353 , \21354 );
and \U$21224 ( \21356 , \21291 , \21295 );
and \U$21225 ( \21357 , \21295 , \21297 );
and \U$21226 ( \21358 , \21291 , \21297 );
or \U$21227 ( \21359 , \21356 , \21357 , \21358 );
and \U$21228 ( \21360 , \21309 , \21323 );
and \U$21229 ( \21361 , \21323 , \21335 );
and \U$21230 ( \21362 , \21309 , \21335 );
or \U$21231 ( \21363 , \21360 , \21361 , \21362 );
xor \U$21232 ( \21364 , \21359 , \21363 );
and \U$21233 ( \21365 , \8652 , \9765 );
and \U$21234 ( \21366 , \8835 , \9644 );
nor \U$21235 ( \21367 , \21365 , \21366 );
xnor \U$21236 ( \21368 , \21367 , \9478 );
and \U$21237 ( \21369 , \8057 , \10408 );
and \U$21238 ( \21370 , \8349 , \10116 );
nor \U$21239 ( \21371 , \21369 , \21370 );
xnor \U$21240 ( \21372 , \21371 , \10121 );
xor \U$21241 ( \21373 , \21368 , \21372 );
and \U$21242 ( \21374 , \7700 , \10118 );
xor \U$21243 ( \21375 , \21373 , \21374 );
xor \U$21244 ( \21376 , \21364 , \21375 );
xor \U$21245 ( \21377 , \21355 , \21376 );
and \U$21246 ( \21378 , \10584 , \8019 );
not \U$21247 ( \21379 , \21378 );
xnor \U$21248 ( \21380 , \21379 , \7713 );
and \U$21249 ( \21381 , \9897 , \8540 );
and \U$21250 ( \21382 , \10206 , \8292 );
nor \U$21251 ( \21383 , \21381 , \21382 );
xnor \U$21252 ( \21384 , \21383 , \8297 );
xor \U$21253 ( \21385 , \21380 , \21384 );
and \U$21254 ( \21386 , \9169 , \9333 );
and \U$21255 ( \21387 , \9465 , \9006 );
nor \U$21256 ( \21388 , \21386 , \21387 );
xnor \U$21257 ( \21389 , \21388 , \8848 );
xor \U$21258 ( \21390 , \21385 , \21389 );
and \U$21259 ( \21391 , \21313 , \21317 );
and \U$21260 ( \21392 , \21317 , \21322 );
and \U$21261 ( \21393 , \21313 , \21322 );
or \U$21262 ( \21394 , \21391 , \21392 , \21393 );
and \U$21263 ( \21395 , \21325 , \21329 );
and \U$21264 ( \21396 , \21329 , \21334 );
and \U$21265 ( \21397 , \21325 , \21334 );
or \U$21266 ( \21398 , \21395 , \21396 , \21397 );
xnor \U$21267 ( \21399 , \21394 , \21398 );
xor \U$21268 ( \21400 , \21390 , \21399 );
xor \U$21269 ( \21401 , \21377 , \21400 );
xor \U$21270 ( \21402 , \21351 , \21401 );
and \U$21271 ( \21403 , \21283 , \21338 );
xor \U$21272 ( \21404 , \21402 , \21403 );
and \U$21273 ( \21405 , \21339 , \21340 );
and \U$21274 ( \21406 , \21341 , \21344 );
or \U$21275 ( \21407 , \21405 , \21406 );
xor \U$21276 ( \21408 , \21404 , \21407 );
buf \U$21277 ( \21409 , \21408 );
buf \U$21278 ( \21410 , \21409 );
and \U$21279 ( \21411 , \21355 , \21376 );
and \U$21280 ( \21412 , \21376 , \21400 );
and \U$21281 ( \21413 , \21355 , \21400 );
or \U$21282 ( \21414 , \21411 , \21412 , \21413 );
and \U$21283 ( \21415 , \21359 , \21363 );
and \U$21284 ( \21416 , \21363 , \21375 );
and \U$21285 ( \21417 , \21359 , \21375 );
or \U$21286 ( \21418 , \21415 , \21416 , \21417 );
and \U$21287 ( \21419 , \21390 , \21399 );
xor \U$21288 ( \21420 , \21418 , \21419 );
or \U$21289 ( \21421 , \21394 , \21398 );
not \U$21290 ( \21422 , \7713 );
and \U$21291 ( \21423 , \10206 , \8540 );
and \U$21292 ( \21424 , \10584 , \8292 );
nor \U$21293 ( \21425 , \21423 , \21424 );
xnor \U$21294 ( \21426 , \21425 , \8297 );
xor \U$21295 ( \21427 , \21422 , \21426 );
and \U$21296 ( \21428 , \9465 , \9333 );
and \U$21297 ( \21429 , \9897 , \9006 );
nor \U$21298 ( \21430 , \21428 , \21429 );
xnor \U$21299 ( \21431 , \21430 , \8848 );
xor \U$21300 ( \21432 , \21427 , \21431 );
xor \U$21301 ( \21433 , \21421 , \21432 );
and \U$21302 ( \21434 , \21380 , \21384 );
and \U$21303 ( \21435 , \21384 , \21389 );
and \U$21304 ( \21436 , \21380 , \21389 );
or \U$21305 ( \21437 , \21434 , \21435 , \21436 );
and \U$21306 ( \21438 , \21368 , \21372 );
and \U$21307 ( \21439 , \21372 , \21374 );
and \U$21308 ( \21440 , \21368 , \21374 );
or \U$21309 ( \21441 , \21438 , \21439 , \21440 );
xor \U$21310 ( \21442 , \21437 , \21441 );
and \U$21311 ( \21443 , \8835 , \9765 );
and \U$21312 ( \21444 , \9169 , \9644 );
nor \U$21313 ( \21445 , \21443 , \21444 );
xnor \U$21314 ( \21446 , \21445 , \9478 );
and \U$21315 ( \21447 , \8349 , \10408 );
and \U$21316 ( \21448 , \8652 , \10116 );
nor \U$21317 ( \21449 , \21447 , \21448 );
xnor \U$21318 ( \21450 , \21449 , \10121 );
xor \U$21319 ( \21451 , \21446 , \21450 );
and \U$21320 ( \21452 , \8057 , \10118 );
xor \U$21321 ( \21453 , \21451 , \21452 );
xor \U$21322 ( \21454 , \21442 , \21453 );
xor \U$21323 ( \21455 , \21433 , \21454 );
xor \U$21324 ( \21456 , \21420 , \21455 );
xor \U$21325 ( \21457 , \21414 , \21456 );
and \U$21326 ( \21458 , \21351 , \21401 );
xor \U$21327 ( \21459 , \21457 , \21458 );
and \U$21328 ( \21460 , \21402 , \21403 );
and \U$21329 ( \21461 , \21404 , \21407 );
or \U$21330 ( \21462 , \21460 , \21461 );
xor \U$21331 ( \21463 , \21459 , \21462 );
buf \U$21332 ( \21464 , \21463 );
buf \U$21333 ( \21465 , \21464 );
and \U$21334 ( \21466 , \21421 , \21432 );
and \U$21335 ( \21467 , \21432 , \21454 );
and \U$21336 ( \21468 , \21421 , \21454 );
or \U$21337 ( \21469 , \21466 , \21467 , \21468 );
and \U$21338 ( \21470 , \21418 , \21419 );
and \U$21339 ( \21471 , \21419 , \21455 );
and \U$21340 ( \21472 , \21418 , \21455 );
or \U$21341 ( \21473 , \21470 , \21471 , \21472 );
xor \U$21342 ( \21474 , \21469 , \21473 );
and \U$21343 ( \21475 , \21437 , \21441 );
and \U$21344 ( \21476 , \21441 , \21453 );
and \U$21345 ( \21477 , \21437 , \21453 );
or \U$21346 ( \21478 , \21475 , \21476 , \21477 );
and \U$21347 ( \21479 , \10584 , \8540 );
not \U$21348 ( \21480 , \21479 );
xnor \U$21349 ( \21481 , \21480 , \8297 );
and \U$21350 ( \21482 , \9897 , \9333 );
and \U$21351 ( \21483 , \10206 , \9006 );
nor \U$21352 ( \21484 , \21482 , \21483 );
xnor \U$21353 ( \21485 , \21484 , \8848 );
xor \U$21354 ( \21486 , \21481 , \21485 );
and \U$21355 ( \21487 , \9169 , \9765 );
and \U$21356 ( \21488 , \9465 , \9644 );
nor \U$21357 ( \21489 , \21487 , \21488 );
xnor \U$21358 ( \21490 , \21489 , \9478 );
xor \U$21359 ( \21491 , \21486 , \21490 );
xor \U$21360 ( \21492 , \21478 , \21491 );
and \U$21361 ( \21493 , \21422 , \21426 );
and \U$21362 ( \21494 , \21426 , \21431 );
and \U$21363 ( \21495 , \21422 , \21431 );
or \U$21364 ( \21496 , \21493 , \21494 , \21495 );
and \U$21365 ( \21497 , \21446 , \21450 );
and \U$21366 ( \21498 , \21450 , \21452 );
and \U$21367 ( \21499 , \21446 , \21452 );
or \U$21368 ( \21500 , \21497 , \21498 , \21499 );
xor \U$21369 ( \21501 , \21496 , \21500 );
and \U$21370 ( \21502 , \8652 , \10408 );
and \U$21371 ( \21503 , \8835 , \10116 );
nor \U$21372 ( \21504 , \21502 , \21503 );
xnor \U$21373 ( \21505 , \21504 , \10121 );
and \U$21374 ( \21506 , \8349 , \10118 );
xnor \U$21375 ( \21507 , \21505 , \21506 );
xor \U$21376 ( \21508 , \21501 , \21507 );
xor \U$21377 ( \21509 , \21492 , \21508 );
xor \U$21378 ( \21510 , \21474 , \21509 );
and \U$21379 ( \21511 , \21414 , \21456 );
xor \U$21380 ( \21512 , \21510 , \21511 );
and \U$21381 ( \21513 , \21457 , \21458 );
and \U$21382 ( \21514 , \21459 , \21462 );
or \U$21383 ( \21515 , \21513 , \21514 );
xor \U$21384 ( \21516 , \21512 , \21515 );
buf \U$21385 ( \21517 , \21516 );
buf \U$21386 ( \21518 , \21517 );
and \U$21387 ( \21519 , \21478 , \21491 );
and \U$21388 ( \21520 , \21491 , \21508 );
and \U$21389 ( \21521 , \21478 , \21508 );
or \U$21390 ( \21522 , \21519 , \21520 , \21521 );
and \U$21391 ( \21523 , \21496 , \21500 );
and \U$21392 ( \21524 , \21500 , \21507 );
and \U$21393 ( \21525 , \21496 , \21507 );
or \U$21394 ( \21526 , \21523 , \21524 , \21525 );
and \U$21395 ( \21527 , \21481 , \21485 );
and \U$21396 ( \21528 , \21485 , \21490 );
and \U$21397 ( \21529 , \21481 , \21490 );
or \U$21398 ( \21530 , \21527 , \21528 , \21529 );
or \U$21399 ( \21531 , \21505 , \21506 );
xor \U$21400 ( \21532 , \21530 , \21531 );
and \U$21401 ( \21533 , \8835 , \10408 );
and \U$21402 ( \21534 , \9169 , \10116 );
nor \U$21403 ( \21535 , \21533 , \21534 );
xnor \U$21404 ( \21536 , \21535 , \10121 );
xor \U$21405 ( \21537 , \21532 , \21536 );
xor \U$21406 ( \21538 , \21526 , \21537 );
and \U$21407 ( \21539 , \8652 , \10118 );
not \U$21408 ( \21540 , \8297 );
and \U$21409 ( \21541 , \10206 , \9333 );
and \U$21410 ( \21542 , \10584 , \9006 );
nor \U$21411 ( \21543 , \21541 , \21542 );
xnor \U$21412 ( \21544 , \21543 , \8848 );
xor \U$21413 ( \21545 , \21540 , \21544 );
and \U$21414 ( \21546 , \9465 , \9765 );
and \U$21415 ( \21547 , \9897 , \9644 );
nor \U$21416 ( \21548 , \21546 , \21547 );
xnor \U$21417 ( \21549 , \21548 , \9478 );
xor \U$21418 ( \21550 , \21545 , \21549 );
xor \U$21419 ( \21551 , \21539 , \21550 );
xor \U$21420 ( \21552 , \21538 , \21551 );
xor \U$21421 ( \21553 , \21522 , \21552 );
and \U$21422 ( \21554 , \21469 , \21473 );
and \U$21423 ( \21555 , \21473 , \21509 );
and \U$21424 ( \21556 , \21469 , \21509 );
or \U$21425 ( \21557 , \21554 , \21555 , \21556 );
xor \U$21426 ( \21558 , \21553 , \21557 );
and \U$21427 ( \21559 , \21510 , \21511 );
and \U$21428 ( \21560 , \21512 , \21515 );
or \U$21429 ( \21561 , \21559 , \21560 );
xor \U$21430 ( \21562 , \21558 , \21561 );
buf \U$21431 ( \21563 , \21562 );
buf \U$21432 ( \21564 , \21563 );
and \U$21433 ( \21565 , \21526 , \21537 );
and \U$21434 ( \21566 , \21537 , \21551 );
and \U$21435 ( \21567 , \21526 , \21551 );
or \U$21436 ( \21568 , \21565 , \21566 , \21567 );
and \U$21437 ( \21569 , \21530 , \21531 );
and \U$21438 ( \21570 , \21531 , \21536 );
and \U$21439 ( \21571 , \21530 , \21536 );
or \U$21440 ( \21572 , \21569 , \21570 , \21571 );
and \U$21441 ( \21573 , \21539 , \21550 );
xor \U$21442 ( \21574 , \21572 , \21573 );
and \U$21443 ( \21575 , \21540 , \21544 );
and \U$21444 ( \21576 , \21544 , \21549 );
and \U$21445 ( \21577 , \21540 , \21549 );
or \U$21446 ( \21578 , \21575 , \21576 , \21577 );
and \U$21447 ( \21579 , \10584 , \9333 );
not \U$21448 ( \21580 , \21579 );
xnor \U$21449 ( \21581 , \21580 , \8848 );
and \U$21450 ( \21582 , \9897 , \9765 );
and \U$21451 ( \21583 , \10206 , \9644 );
nor \U$21452 ( \21584 , \21582 , \21583 );
xnor \U$21453 ( \21585 , \21584 , \9478 );
xor \U$21454 ( \21586 , \21581 , \21585 );
and \U$21455 ( \21587 , \9169 , \10408 );
and \U$21456 ( \21588 , \9465 , \10116 );
nor \U$21457 ( \21589 , \21587 , \21588 );
xnor \U$21458 ( \21590 , \21589 , \10121 );
xor \U$21459 ( \21591 , \21586 , \21590 );
xor \U$21460 ( \21592 , \21578 , \21591 );
and \U$21461 ( \21593 , \8835 , \10118 );
not \U$21462 ( \21594 , \21593 );
xor \U$21463 ( \21595 , \21592 , \21594 );
xor \U$21464 ( \21596 , \21574 , \21595 );
xor \U$21465 ( \21597 , \21568 , \21596 );
and \U$21466 ( \21598 , \21522 , \21552 );
xor \U$21467 ( \21599 , \21597 , \21598 );
and \U$21468 ( \21600 , \21553 , \21557 );
and \U$21469 ( \21601 , \21558 , \21561 );
or \U$21470 ( \21602 , \21600 , \21601 );
xor \U$21471 ( \21603 , \21599 , \21602 );
buf \U$21472 ( \21604 , \21603 );
buf \U$21473 ( \21605 , \21604 );
and \U$21474 ( \21606 , \21572 , \21573 );
and \U$21475 ( \21607 , \21573 , \21595 );
and \U$21476 ( \21608 , \21572 , \21595 );
or \U$21477 ( \21609 , \21606 , \21607 , \21608 );
and \U$21478 ( \21610 , \21578 , \21591 );
and \U$21479 ( \21611 , \21591 , \21594 );
and \U$21480 ( \21612 , \21578 , \21594 );
or \U$21481 ( \21613 , \21610 , \21611 , \21612 );
not \U$21482 ( \21614 , \8848 );
and \U$21483 ( \21615 , \10206 , \9765 );
and \U$21484 ( \21616 , \10584 , \9644 );
nor \U$21485 ( \21617 , \21615 , \21616 );
xnor \U$21486 ( \21618 , \21617 , \9478 );
xor \U$21487 ( \21619 , \21614 , \21618 );
and \U$21488 ( \21620 , \9465 , \10408 );
and \U$21489 ( \21621 , \9897 , \10116 );
nor \U$21490 ( \21622 , \21620 , \21621 );
xnor \U$21491 ( \21623 , \21622 , \10121 );
xor \U$21492 ( \21624 , \21619 , \21623 );
xor \U$21493 ( \21625 , \21613 , \21624 );
and \U$21494 ( \21626 , \21581 , \21585 );
and \U$21495 ( \21627 , \21585 , \21590 );
and \U$21496 ( \21628 , \21581 , \21590 );
or \U$21497 ( \21629 , \21626 , \21627 , \21628 );
buf \U$21498 ( \21630 , \21593 );
xor \U$21499 ( \21631 , \21629 , \21630 );
and \U$21500 ( \21632 , \9169 , \10118 );
xor \U$21501 ( \21633 , \21631 , \21632 );
xor \U$21502 ( \21634 , \21625 , \21633 );
xor \U$21503 ( \21635 , \21609 , \21634 );
and \U$21504 ( \21636 , \21568 , \21596 );
xor \U$21505 ( \21637 , \21635 , \21636 );
and \U$21506 ( \21638 , \21597 , \21598 );
and \U$21507 ( \21639 , \21599 , \21602 );
or \U$21508 ( \21640 , \21638 , \21639 );
xor \U$21509 ( \21641 , \21637 , \21640 );
buf \U$21510 ( \21642 , \21641 );
buf \U$21511 ( \21643 , \21642 );
and \U$21512 ( \21644 , \21629 , \21630 );
and \U$21513 ( \21645 , \21630 , \21632 );
and \U$21514 ( \21646 , \21629 , \21632 );
or \U$21515 ( \21647 , \21644 , \21645 , \21646 );
and \U$21516 ( \21648 , \21613 , \21624 );
and \U$21517 ( \21649 , \21624 , \21633 );
and \U$21518 ( \21650 , \21613 , \21633 );
or \U$21519 ( \21651 , \21648 , \21649 , \21650 );
xor \U$21520 ( \21652 , \21647 , \21651 );
and \U$21521 ( \21653 , \21614 , \21618 );
and \U$21522 ( \21654 , \21618 , \21623 );
and \U$21523 ( \21655 , \21614 , \21623 );
or \U$21524 ( \21656 , \21653 , \21654 , \21655 );
and \U$21525 ( \21657 , \10584 , \9765 );
not \U$21526 ( \21658 , \21657 );
xnor \U$21527 ( \21659 , \21658 , \9478 );
and \U$21528 ( \21660 , \9897 , \10408 );
and \U$21529 ( \21661 , \10206 , \10116 );
nor \U$21530 ( \21662 , \21660 , \21661 );
xnor \U$21531 ( \21663 , \21662 , \10121 );
xor \U$21532 ( \21664 , \21659 , \21663 );
and \U$21533 ( \21665 , \9465 , \10118 );
xor \U$21534 ( \21666 , \21664 , \21665 );
xnor \U$21535 ( \21667 , \21656 , \21666 );
xor \U$21536 ( \21668 , \21652 , \21667 );
and \U$21537 ( \21669 , \21609 , \21634 );
xor \U$21538 ( \21670 , \21668 , \21669 );
and \U$21539 ( \21671 , \21635 , \21636 );
and \U$21540 ( \21672 , \21637 , \21640 );
or \U$21541 ( \21673 , \21671 , \21672 );
xor \U$21542 ( \21674 , \21670 , \21673 );
buf \U$21543 ( \21675 , \21674 );
buf \U$21544 ( \21676 , \21675 );
and \U$21545 ( \21677 , \21659 , \21663 );
and \U$21546 ( \21678 , \21663 , \21665 );
and \U$21547 ( \21679 , \21659 , \21665 );
or \U$21548 ( \21680 , \21677 , \21678 , \21679 );
or \U$21549 ( \21681 , \21656 , \21666 );
xor \U$21550 ( \21682 , \21680 , \21681 );
not \U$21551 ( \21683 , \9478 );
and \U$21552 ( \21684 , \10206 , \10408 );
and \U$21553 ( \21685 , \10584 , \10116 );
nor \U$21554 ( \21686 , \21684 , \21685 );
xnor \U$21555 ( \21687 , \21686 , \10121 );
xor \U$21556 ( \21688 , \21683 , \21687 );
and \U$21557 ( \21689 , \9897 , \10118 );
xor \U$21558 ( \21690 , \21688 , \21689 );
xor \U$21559 ( \21691 , \21682 , \21690 );
and \U$21560 ( \21692 , \21647 , \21651 );
and \U$21561 ( \21693 , \21651 , \21667 );
and \U$21562 ( \21694 , \21647 , \21667 );
or \U$21563 ( \21695 , \21692 , \21693 , \21694 );
xor \U$21564 ( \21696 , \21691 , \21695 );
and \U$21565 ( \21697 , \21668 , \21669 );
and \U$21566 ( \21698 , \21670 , \21673 );
or \U$21567 ( \21699 , \21697 , \21698 );
xor \U$21568 ( \21700 , \21696 , \21699 );
buf \U$21569 ( \21701 , \21700 );
buf \U$21570 ( \21702 , \21701 );
and \U$21571 ( \21703 , \21683 , \21687 );
and \U$21572 ( \21704 , \21687 , \21689 );
and \U$21573 ( \21705 , \21683 , \21689 );
or \U$21574 ( \21706 , \21703 , \21704 , \21705 );
and \U$21575 ( \21707 , \10584 , \10408 );
not \U$21576 ( \21708 , \21707 );
xnor \U$21577 ( \21709 , \21708 , \10121 );
and \U$21578 ( \21710 , \10206 , \10118 );
xnor \U$21579 ( \21711 , \21709 , \21710 );
xor \U$21580 ( \21712 , \21706 , \21711 );
and \U$21581 ( \21713 , \21680 , \21681 );
and \U$21582 ( \21714 , \21681 , \21690 );
and \U$21583 ( \21715 , \21680 , \21690 );
or \U$21584 ( \21716 , \21713 , \21714 , \21715 );
xor \U$21585 ( \21717 , \21712 , \21716 );
and \U$21586 ( \21718 , \21691 , \21695 );
and \U$21587 ( \21719 , \21696 , \21699 );
or \U$21588 ( \21720 , \21718 , \21719 );
xor \U$21589 ( \21721 , \21717 , \21720 );
buf \U$21590 ( \21722 , \21721 );
buf \U$21591 ( \21723 , \21722 );
or \U$21592 ( \21724 , \21709 , \21710 );
not \U$21593 ( \21725 , \10121 );
xor \U$21594 ( \21726 , \21724 , \21725 );
and \U$21595 ( \21727 , \10584 , \10118 );
xor \U$21596 ( \21728 , \21726 , \21727 );
and \U$21597 ( \21729 , \21706 , \21711 );
xor \U$21598 ( \21730 , \21728 , \21729 );
and \U$21599 ( \21731 , \21712 , \21716 );
and \U$21600 ( \21732 , \21717 , \21720 );
or \U$21601 ( \21733 , \21731 , \21732 );
xor \U$21602 ( \21734 , \21730 , \21733 );
buf \U$21603 ( \21735 , \21734 );
buf \U$21604 ( \21736 , \21735 );
xor \U$21605 ( \21737 , \649 , \1063 );
buf \U$21606 ( \21738 , \21737 );
buf \U$21607 ( \21739 , \21738 );
xor \U$21608 ( \21740 , \594 , \1065 );
buf \U$21609 ( \21741 , \21740 );
buf \U$21610 ( \21742 , \21741 );
xor \U$21611 ( \21743 , \865 , \1055 );
buf \U$21612 ( \21744 , \21743 );
buf \U$21613 ( \21745 , \21744 );
xor \U$21614 ( \21746 , \812 , \1057 );
buf \U$21615 ( \21747 , \21746 );
buf \U$21616 ( \21748 , \21747 );
xor \U$21617 ( \21749 , \773 , \1059 );
buf \U$21618 ( \21750 , \21749 );
buf \U$21619 ( \21751 , \21750 );
xor \U$21620 ( \21752 , \720 , \1061 );
buf \U$21621 ( \21753 , \21752 );
buf \U$21622 ( \21754 , \21753 );
xor \U$21623 ( \21755 , \907 , \1051 );
buf \U$21624 ( \21756 , \21755 );
buf \U$21625 ( \21757 , \21756 );
xor \U$21626 ( \21758 , \873 , \1053 );
buf \U$21627 ( \21759 , \21758 );
buf \U$21628 ( \21760 , \21759 );
xor \U$21629 ( \21761 , \941 , \1049 );
buf \U$21630 ( \21762 , \21761 );
buf \U$21631 ( \21763 , \21762 );
xor \U$21632 ( \21764 , \949 , \1047 );
buf \U$21633 ( \21765 , \21764 );
buf \U$21634 ( \21766 , \21765 );
xor \U$21635 ( \21767 , \994 , \1043 );
buf \U$21636 ( \21768 , \21767 );
buf \U$21637 ( \21769 , \21768 );
xor \U$21638 ( \21770 , \975 , \1045 );
buf \U$21639 ( \21771 , \21770 );
buf \U$21640 ( \21772 , \21771 );
or \U$21641 ( \21773 , \21769 , \21772 );
and \U$21642 ( \21774 , \21766 , \21773 );
or \U$21643 ( \21775 , \21763 , \21774 );
and \U$21644 ( \21776 , \21757 , \21760 , \21775 );
or \U$21645 ( \21777 , \21745 , \21748 , \21751 , \21754 , \21776 );
and \U$21646 ( \21778 , \21739 , \21742 , \21777 );
or \U$21647 ( \21779 , \16027 , \16264 , \16499 , \16727 , \16951 , \17169 , \17382 , \17587 , \17790 , \17985 , \18178 , \18364 , \18545 , \18718 , \18888 , \19053 , \19216 , \19376 , \19531 , \19679 , \19822 , \19957 , \20091 , \20219 , \20342 , \20458 , \20568 , \20673 , \20776 , \20871 , \20964 , \21049 , \21132 , \21208 , \21279 , \21347 , \21410 , \21465 , \21518 , \21564 , \21605 , \21643 , \21676 , \21702 , \21723 , \21736 , \21778 );
or \U$21648 ( \21780 , \15782 , \21779 );
buf \U$21649 ( \21781 , \21780 );
buf \U$21650 ( \21782 , \1069 );
buf \U$21651 ( \21783 , \1170 );
buf \U$21652 ( \21784 , \1278 );
buf \U$21653 ( \21785 , \1389 );
buf \U$21654 ( \21786 , \1507 );
buf \U$21655 ( \21787 , \1628 );
buf \U$21656 ( \21788 , \1756 );
buf \U$21657 ( \21789 , \1887 );
buf \U$21658 ( \21790 , \2025 );
buf \U$21659 ( \21791 , \2166 );
buf \U$21660 ( \21792 , \2314 );
buf \U$21661 ( \21793 , \2465 );
buf \U$21662 ( \21794 , \2623 );
buf \U$21663 ( \21795 , \2784 );
buf \U$21664 ( \21796 , \2952 );
buf \U$21665 ( \21797 , \3123 );
buf \U$21666 ( \21798 , \3301 );
buf \U$21667 ( \21799 , \3482 );
buf \U$21668 ( \21800 , \3670 );
buf \U$21669 ( \21801 , \3861 );
buf \U$21670 ( \21802 , \4059 );
buf \U$21671 ( \21803 , \4260 );
buf \U$21672 ( \21804 , \4468 );
buf \U$21673 ( \21805 , \4679 );
buf \U$21674 ( \21806 , \4897 );
buf \U$21675 ( \21807 , \5117 );
buf \U$21676 ( \21808 , \5348 );
buf \U$21677 ( \21809 , \5579 );
buf \U$21678 ( \21810 , \5817 );
buf \U$21679 ( \21811 , \6058 );
buf \U$21680 ( \21812 , \6306 );
buf \U$21681 ( \21813 , \6557 );
buf \U$21682 ( \21814 , \6815 );
buf \U$21683 ( \21815 , \7076 );
buf \U$21684 ( \21816 , \7344 );
buf \U$21685 ( \21817 , \7615 );
buf \U$21686 ( \21818 , \7893 );
buf \U$21687 ( \21819 , \8174 );
buf \U$21688 ( \21820 , \8462 );
buf \U$21689 ( \21821 , \8753 );
buf \U$21690 ( \21822 , \9051 );
buf \U$21691 ( \21823 , \9352 );
buf \U$21692 ( \21824 , \9660 );
buf \U$21693 ( \21825 , \9971 );
buf \U$21694 ( \21826 , \10289 );
buf \U$21695 ( \21827 , \10610 );
buf \U$21696 ( \21828 , \10929 );
buf \U$21697 ( \21829 , \11247 );
buf \U$21698 ( \21830 , \11564 );
buf \U$21699 ( \21831 , \11880 );
buf \U$21700 ( \21832 , \12191 );
buf \U$21701 ( \21833 , \12499 );
buf \U$21702 ( \21834 , \12802 );
buf \U$21703 ( \21835 , \13098 );
buf \U$21704 ( \21836 , \13389 );
buf \U$21705 ( \21837 , \13672 );
buf \U$21706 ( \21838 , \13953 );
buf \U$21707 ( \21839 , \14226 );
buf \U$21708 ( \21840 , \14496 );
buf \U$21709 ( \21841 , \14762 );
buf \U$21710 ( \21842 , \15022 );
buf \U$21711 ( \21843 , \15277 );
buf \U$21712 ( \21844 , \15530 );
buf \U$21713 ( \21845 , \15780 );
or \U$21714 ( \21846 , \21782 , \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 );
buf \U$21715 ( \21847 , \16026 );
buf \U$21716 ( \21848 , \16263 );
buf \U$21717 ( \21849 , \16498 );
buf \U$21718 ( \21850 , \16726 );
buf \U$21719 ( \21851 , \16950 );
buf \U$21720 ( \21852 , \17168 );
buf \U$21721 ( \21853 , \17381 );
buf \U$21722 ( \21854 , \17586 );
buf \U$21723 ( \21855 , \17789 );
buf \U$21724 ( \21856 , \17984 );
buf \U$21725 ( \21857 , \18177 );
buf \U$21726 ( \21858 , \18363 );
buf \U$21727 ( \21859 , \18544 );
buf \U$21728 ( \21860 , \18717 );
buf \U$21729 ( \21861 , \18887 );
buf \U$21730 ( \21862 , \19052 );
buf \U$21731 ( \21863 , \19215 );
buf \U$21732 ( \21864 , \19375 );
buf \U$21733 ( \21865 , \19530 );
buf \U$21734 ( \21866 , \19678 );
buf \U$21735 ( \21867 , \19821 );
buf \U$21736 ( \21868 , \19956 );
buf \U$21737 ( \21869 , \20090 );
buf \U$21738 ( \21870 , \20218 );
buf \U$21739 ( \21871 , \20341 );
buf \U$21740 ( \21872 , \20457 );
buf \U$21741 ( \21873 , \20567 );
buf \U$21742 ( \21874 , \20672 );
buf \U$21743 ( \21875 , \20775 );
buf \U$21744 ( \21876 , \20870 );
buf \U$21745 ( \21877 , \20963 );
buf \U$21746 ( \21878 , \21048 );
buf \U$21747 ( \21879 , \21131 );
buf \U$21748 ( \21880 , \21207 );
buf \U$21749 ( \21881 , \21278 );
buf \U$21750 ( \21882 , \21346 );
buf \U$21751 ( \21883 , \21409 );
buf \U$21752 ( \21884 , \21464 );
buf \U$21753 ( \21885 , \21517 );
buf \U$21754 ( \21886 , \21563 );
buf \U$21755 ( \21887 , \21604 );
buf \U$21756 ( \21888 , \21642 );
buf \U$21757 ( \21889 , \21675 );
buf \U$21758 ( \21890 , \21701 );
buf \U$21759 ( \21891 , \21722 );
buf \U$21760 ( \21892 , \21735 );
buf \U$21761 ( \21893 , \21738 );
buf \U$21762 ( \21894 , \21741 );
buf \U$21763 ( \21895 , \21750 );
buf \U$21764 ( \21896 , \21753 );
buf \U$21765 ( \21897 , \21759 );
buf \U$21766 ( \21898 , \21744 );
buf \U$21767 ( \21899 , \21747 );
buf \U$21768 ( \21900 , \21765 );
buf \U$21769 ( \21901 , \21762 );
buf \U$21770 ( \21902 , \21756 );
buf \U$21771 ( \21903 , \21771 );
buf \U$21772 ( \21904 , \21768 );
xor \U$21773 ( \21905 , \1002 , \1041 );
buf \U$21774 ( \21906 , \21905 );
buf \U$21775 ( \21907 , \21906 );
xor \U$21776 ( \21908 , \1022 , \1037 );
buf \U$21777 ( \21909 , \21908 );
buf \U$21778 ( \21910 , \21909 );
xor \U$21779 ( \21911 , \1014 , \1039 );
buf \U$21780 ( \21912 , \21911 );
buf \U$21781 ( \21913 , \21912 );
xor \U$21782 ( \21914 , \1033 , \179 );
buf \U$21783 ( \21915 , \21914 );
buf \U$21784 ( \21916 , \21915 );
xor \U$21785 ( \21917 , \1031 , \1034 );
buf \U$21786 ( \21918 , \21917 );
buf \U$21787 ( \21919 , \21918 );
xor \U$21788 ( \21920 , \1027 , \1035 );
buf \U$21789 ( \21921 , \21920 );
buf \U$21790 ( \21922 , \21921 );
and \U$21791 ( \21923 , \21916 , \21919 , \21922 );
or \U$21792 ( \21924 , \21910 , \21913 , \21923 );
and \U$21793 ( \21925 , \21907 , \21924 );
or \U$21794 ( \21926 , \21904 , \21925 );
and \U$21795 ( \21927 , \21903 , \21926 );
or \U$21796 ( \21928 , \21900 , \21901 , \21902 , \21927 );
and \U$21797 ( \21929 , \21897 , \21898 , \21899 , \21928 );
or \U$21798 ( \21930 , \21895 , \21896 , \21929 );
and \U$21799 ( \21931 , \21893 , \21894 , \21930 );
or \U$21800 ( \21932 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21931 );
nor \U$21801 ( \21933 , \21846 , \21932 );
buf \U$21802 ( \21934 , \21933 );
and \U$21803 ( \21935 , \21781 , \21934 );
not \U$21804 ( \21936 , \21935 );
_DC r56af ( \21937_nR56af , 1'b0 , \21936 );
buf \U$21805 ( \21938 , \21937_nR56af );
endmodule

