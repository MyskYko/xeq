//
// Conformal-LEC Version 20.10-d132 (30-Jun-2020)
//
module top(RIde68638_3981,RIde67cd8_3982,RIde68f20_3980,RIb79b518_270,RIdbb8138_3227,RIe548ff0_6844,RIe549ef0_6842,RIe5319e0_6884,RIe549770_6843,
        RIe4f85f0_6398,RIdaea590_2835,RIe4301f0_6000,RIde3d1e0_4027,RIe00b330_4420,RIe160838_5254,RIe0d49f0_4816,RIda11c00_2446,RIe269120_5609,RId958f08_2058,
        RId888d80_1669,RIdc6ed48_3642,RIe5c2e08_6791,RId6f3a80_883,RId7bf4e0_1272,RIb7b93b0_251,RIdba4548_3251,RIe4fa198_6396,RIdaebc88_2833,RIe431ac8_5998,
        RIde3ed88_4025,RIe00ce60_4418,RIe1615d0_5253,RIe0d62c8_4814,RIda13640_2444,RIe26a7a0_5607,RId95a600_2056,RId88a478_1667,RIdc70800_3640,RIe5c4500_6789,
        RId6f5100_881,RId7c0e30_1270,RIb7b94a0_249,RIdbb7328_3228,RIe4f7a38_6399,RIdae97f8_2836,RIe42f4d0_6001,RIde3c448_4028,RIe00a598_4421,RIe172718_5244,
        RIe0d3dc0_4817,RIda10df0_2447,RIe268568_5610,RId9582d8_2059,RId888240_1670,RIdc6e280_3643,RIe5c22c8_6792,RId7064a0_859,RId7be838_1273,RIb7af720_252,
        RIdbb6518_3229,RIe4f6ef8_6400,RIdae8a60_2837,RIe42e8a0_6002,RIde3b728_4029,RIe009710_4422,RIe163e20_5250,RIe0d2e48_4818,RIda101c0_2448,RIe2679b0_5611,
        RId957720_2060,RId89b638_1645,RIdc6d740_3644,RIe5c1710_6793,RId705780_860,RId7d2338_1248,RIb7af6a8_253,RIe4faf30_6395,RIdba51f0_3250,RIe4326f8_5997,
        RIdad5d70_2860,RIde3fb20_4024,RIe00db80_4417,RIe164b40_5249,RIe0d6fe8_4813,RIda143d8_2443,RIe26b2e0_5606,RId95b1b8_2055,RId88b030_1666,RIdc71610_3639,
        RIe5c4fc8_6788,RId6f5cb8_880,RId7c1b50_1269,RIb7b9518_248,RIdba3828_3252,RIe4f9388_6397,RIdaeb0d0_2834,RIe430e20_5999,RIde3df00_4026,RIe00c0c8_4419,
        RIe163088_5251,RIe0d55a8_4815,RIda12920_2445,RIe269c60_5608,RId959a48_2057,RId889938_1668,RIdc6f9f0_3641,RIe5c3948_6790,RId6f4638_882,RId7c0110_1271,
        RIb7b9428_250,RIdba6bb8_3248,RIe4fc9e8_6393,RIdad7918_2858,RIe4340c0_5995,RIde415d8_4022,RIe00f6b0_4415,RIe162368_5252,RIe0d89b0_4811,RIda15da0_2441,
        RIe26ce10_5604,RId95c8b0_2053,RId88c728_1664,RIdd731d8_3637,RId7c3590_1267,RIe5c6738_6786,RId6f73b0_878,RIb7b9608_246,RIdba5e98_3249,RIe4fbcc8_6394,
        RIdad6b80_2859,RIe4333a0_5996,RIde408b8_4023,RIe00e918_4416,RIe1658d8_5248,RIe0d7d08_4812,RIda150f8_2442,RIe26c000_5605,RId95bcf8_2054,RId88bbe8_1665,
        RIdc72420_3638,RIe5c5bf8_6787,RId6f68e8_879,RId7c2870_1268,RIb7b9590_247,RIe5349b0_6879,RIe5341b8_6880,RIe5339c0_6881,RIe5331c8_6882,RIe5329d0_6883,
        RIeb72150_6905,RIe5359a0_6877,RIe5351a8_6878,RIeab7d00_6896,RIeab78c8_6895,RIeab6518_6891,RIeacfa18_6902,RIeab80c0_6897,RIeb352c8_6904,RIea94af8_6890,
        RIeab87c8_6898,RIe15c260_5259,RIe0f3878_4787,RIde5d760_3998,RIdfce700_4467,RIe3f7760_6049,RIe3887c0_5578,RIe5e3568_6762,RIe51acb8_6366,RId7e6f90_1232,
        RId71e398_838,RId8ac078_1630,RId97ab20_2022,RIdb01d80_2813,RIda2def0_2418,RIdbcc7f0_3208,RIdd963e0_3603,RIb7af3d8_259,RIe182a68_5243,RIe0f3008_4788,
        RIde5ad30_4003,RIdfc11b8_4469,RIe3f8a98_6047,RIe385d90_5583,RIe5e09d0_6767,RIe4af828_6445,RId7e5f28_1234,RId71bad0_843,RId8ab538_1631,RId977f88_2027,
        RIdaff2d8_2817,RIda2b970_2422,RIdbcac48_3211,RIdd93500_3608,RIb7af630_254,RIdaffda0_2816,RIda2c258_2421,RIdb62338_3285,RIdd93ed8_3607,RIde5b618_4002,
        RIdfc07e0_4470,RIe1bcc68_5184,RIe088e38_4865,RId978960_2026,RId8ae508_1629,RId71c2c8_842,RId7827c0_1310,RIe386678_5582,RIe450d88_5972,RIe519818_6368,
        RIe5e1330_6766,RIb7af5b8_255,RIdabee68_2890,RIda2cbb8_2420,RIdb8a760_3284,RIdd95288_3605,RIde5c6f8_4000,RIe02a8c0_4391,RIe1bdd48_5182,RIe0aeb60_4864,
        RId9799c8_2024,RId8aed00_1628,RId71d330_840,RId790848_1309,RIe3876e0_5580,RIe3e5628_6050,RIe51a2e0_6367,RIe5e2488_6764,RIb7af4c8_257,RIe1be5b8_5181,
        RIe0b0870_4861,RIde5dfd0_3997,RIdfcf2b8_4466,RIe451670_5971,RIe388fb8_5577,RIe588848_6840,RIe4bd310_6442,RId7a4bb8_1307,RId71ec08_837,RId86c4d8_1705,
        RId97b318_2021,RIdb02668_2812,RIda2e760_2417,RIdbcd0d8_3207,RIdd96cc8_3602,RIb7a5bf8_260,RIe15b900_5260,RIe0f4070_4786,RIde5e840_3996,RIdfcfc90_4465,
        RIe3f9470_6046,RIe3898a0_5576,RIe5e3e50_6761,RIe4b0a70_6443,RId7e7800_1231,RId71f400_836,RId8b0290_1626,RId97bc00_2020,RIdb02f50_2811,RIda2f0c0_2416,
        RIdbcd9c0_3206,RIdd97538_3601,RIb7a0c48_261,RIe3f9e48_6045,RIe387ed8_5579,RIe5e2d70_6763,RIe4bdce8_6441,RIde5cf68_3999,RIdfcdc38_4468,RIe183440_5242,
        RIe0aff10_4862,RId97a238_2023,RId8af7c8_1627,RId71dba0_839,RId7a41e0_1308,RIda2d4a0_2419,RIdb01498_2814,RIdbcbe18_3209,RIdd95b70_3604,RIb7af450_258,
        RIde5be10_4001,RIe02a050_4392,RIe1bd4d8_5183,RIe0af538_4863,RIe3f8048_6048,RIe386e70_5581,RIe5e1ba0_6765,RIe4b0200_6444,RId9791d0_2025,RId86cf28_1704,
        RId71cb38_841,RId7e6798_1233,RId9cdfc8_2495,RIdb00bb0_2815,RIdbcb530_3210,RIdd94928_3606,RIb7af540_256,RIea91330_6888,RIb7b9680_245,RIde4ec88_4006,
        RIb79b4a0_271,RIb79b338_274,RIde612e8_3992,RIde5fec0_3994,RIde60988_3993,RIde69970_3979,RIde6a2d0_3978,RIde6ad98_3977,RIde63250_3989,RIde62878_3990,
        RIde61e28_3991,RIb839848_152,RIe545dc8_6851,RIe545648_6852,RIea90778_6887,RIe546890_6849,RIe546098_6850,RIb8396e0_155,RIb839668_156,RIb79b3b0_273,
        RIde5f3f8_3995,RIde4c8e8_4009,RIb7b96f8_244,RIde4d6f8_4008,RIb7c20c8_243,RIde431f8_4020,RIb7c5728_242,RIde43f90_4019,RIb7c57a0_241,RIde44da0_4018,
        RIb7c5818_240,RIde45ac0_4017,RIb7c5890_239,RIde468d0_4016,RIb7c5908_238,RIde4fb10_4005,RIb7a09f0_266,RIde49300_4013,RIb7a0a68_265,RIde4a020_4012,
        RIb7a0ae0_264,RIde4ae30_4011,RIb7a0b58_263,RIde4bb50_4010,RIb7a0bd0_262,RIdbee210_3713,RIb839b90_145,RIe667bb0_6885,RIe667f70_6886,RIea91768_6889,
        RIeab7058_6894,RIb87eb00_69,RIb7c5980_237,RIdbecc08_3714,RIb87eb78_68,RIb7c59f8_236,RIdbebab0_3715,RIb87ebf0_67,RIb7c5a70_235,RIdbea4a8_3716,
        RIb882ca0_66,RIb7cade0_234,RIdbe9350_3717,RIb885310_65,RIb7cae58_233,RIdbe7d48_3718,RIb885388_64,RIb7caed0_232,RIdbe6bf0_3719,RIb885400_63,
        RIb7caf48_231,RIdbe5a98_3720,RIb885478_62,RIb7cafc0_230,RIdbe4490_3721,RIb8854f0_61,RIb7cb038_229,RIdbe3338_3722,RIb885568_60,RIb7cb0b0_228,
        RIdbe1d30_3723,RIb8855e0_59,RIb7cb128_227,RIdbe0bd8_3724,RIb885658_58,RIb7d00d8_226,RIdaab098_3725,RIb8856d0_57,RIb8263d8_225,RIdaaf0d0_3726,
        RIb885748_56,RIb826e28_224,RIdab2fa0_3727,RIb8857c0_55,RIb826ea0_223,RIdab8e50_3728,RIb885838_54,RIb826f18_222,RIdabcf00_3729,RIb8858b0_53,
        RIb826f90_221,RIdac3788_3730,RIb885928_52,RIb8293a8_220,RIdac8eb8_3731,RIb8859a0_51,RIb829420_219,RIdacf650_3732,RIb885a18_50,RIb829498_218,
        RIdad4fd8_3733,RIb885a90_49,RIb829510_217,RIdadaf00_3734,RIb885b08_48,RIb829588_216,RIdae2610_3735,RIb885b80_47,RIb829600_215,RIdae8268_3736,
        RIb885bf8_46,RIb829678_214,RIdaef720_3737,RIb885c70_45,RIb8296f0_213,RIdaf4e50_3738,RIb885ce8_44,RIb82dae8_212,RIdafa508_3739,RIb885d60_43,
        RIb82db60_211,RIdafe630_3740,RIb885dd8_42,RIb82dbd8_210,RIdb03b08_3741,RIb885e50_41,RIb82dc50_209,RIdb09d00_3742,RIb885ec8_40,RIb82dcc8_208,
        RIdb0e440_3743,RIb885f40_39,RIb82dd40_207,RIdb13468_3744,RIb885fb8_38,RIb82ddb8_206,RId9d7370_3745,RIb886030_37,RIb82de30_205,RId9d25a0_3746,
        RIb8860a8_36,RIb832228_204,RId9cd0c8_3747,RIb886120_35,RIb8322a0_203,RId9c86b8_3748,RIb886198_34,RIb832318_202,RIda940a0_3749,RIb886210_33,
        RIb832390_201,RIda91850_3750,RIb886288_32,RIb832408_200,RIda8dbd8_3751,RIb886300_31,RIb832480_199,RIda8a7d0_3752,RIb886378_30,RIb8324f8_198,
        RIda86978_3753,RIb8863f0_29,RIb832570_197,RIda835e8_3754,RIb886468_28,RIb8383a8_196,RIda80f00_3755,RIb8864e0_27,RIb838420_195,RIda7daf8_3756,
        RIb886558_26,RIb838498_194,RIda7a7e0_3757,RIb8865d0_25,RIb838510_193,RIda745e8_3758,RIb886648_24,RIb838588_192,RIda6e018_3759,RIb8866c0_23,
        RIb838600_191,RIda65e40_3760,RIb886738_22,RIb838678_190,RIda5f888_3761,RIb8867b0_21,RIb8386f0_189,RIda59780_3762,RIb886828_20,RIb838768_188,
        RIda510f8_3763,RIb8868a0_19,RIb8387e0_187,RIda4aff0_3764,RIb886918_18,RIb838858_186,RId927408_3765,RIb886990_17,RIb8388d0_185,RId943680_3766,
        RIb886a08_16,RIb838948_184,RId96ccd8_3767,RIb886a80_15,RIb8389c0_183,RId988b30_3768,RIb886af8_14,RIb838a38_182,RId90bb68_3769,RIb886b70_13,
        RIb838ab0_181,RId8f7438_3770,RIb886be8_12,RIb838b28_180,RId8d6dc8_3771,RIb886c60_11,RIb838ba0_179,RId6c4d70_3772,RIb886cd8_10,RIb838c18_178,
        RId6ae7c8_3773,RIb886d50_9,RIb838c90_177,RId835578_3774,RIb886dc8_8,RIb838d08_176,RId8a9d50_3775,RIb886e40_7,RIb838d80_175,RId862aa0_3776,
        RIb886eb8_6,RIb838df8_174,RId99e778_3777,RId9ac620_3778,RId9b8290_3779,RId9bdfd8_3780,RId90fe70_3781,RId918b10_3782,RIda42698_3783,RIda33a58_3784,
        RIda28b08_3785,RIda18aa0_3786,RIda0b288_3787,RId9f8d18_3788,RId9ec9a0_3789,RId9e3418_3790,RIdb156a0_3791,RIdb17f68_3792,RIdb1b640_3793,RIdb1df08_3794,
        RIdb215e0_3795,RIdb23ea8_3796,RIdb26c20_3797,RIdb29e48_3798,RIdb2cbc0_3799,RIdb2fde8_3800,RIdb32b60_3801,RIdb35d88_3802,RIdb38b00_3803,RIdb3b3c8_3804,
        RIdb3eaa0_3805,RIdb404e0_3806,RIdb422e0_3807,RIdb43ac8_3808,RIdb45850_3809,RIdb47128_3810,RIdb483e8_3811,RIdb49888_3812,RIdb4abc0_3813,RIdb4c330_3814,
        RIdb4d410_3815,RIdb4e5e0_3816,RIdb4fa08_3817,RIdb51100_3818,RIdb52c30_3819,RIdb541c0_3820,RIdb559a8_3821,RIdb56e48_3822,RIdb58900_3823,RIdb5a070_3824,
        RIdb5b588_3825,RIdb5d0b8_3826,RIdb5e3f0_3827,RIda95720_3828,RIda97598_3829,RIda99a28_3830,RIda9bd50_3831,RIda9df10_3832,RIda9f4a0_3833,RIdaa1228_3834,
        RIdaa2d58_3835,RIdaa4a68_3836,RIdaa6b38_3837,RIdaa89b0_3838,RIdbdf030_3839,RIdbdcd80_3840,RIdbdaff8_3841,RIdbd9540_3842,RIdbd6e58_3843,RIdbd4860_3844,
        RIdbd25b0_3845,RIdbd0030_3846,RIdbcdc18_3847,RIdbcb800_3848,RIdbc9730_3849,RIdbc7a20_3850,RIdbc5e78_3851,RIdbc40f0_3852,RIdbc1f30_3853,RIdbbf938_3854,
        RIdbbd4a8_3855,RIdbba910_3856,RIdbb8480_3857,RIdbb58e8_3858,RIdbb2648_3859,RIdbb0758_3860,RIdbad788_3861,RIdbaad58_3862,RIdba7d88_3863,RIdba55b0_3864,
        RIdba2ce8_3865,RIdb9fe80_3866,RIdb9d4c8_3867,RIdb9acf0_3868,RIdb98c20_3869,RIdb96178_3870,RIdb93ce8_3871,RIdb916f0_3872,RIdb8e2e8_3873,RIdb8b840_3874,
        RIdb890e0_3875,RIdb86cc8_3876,RIdb84ec8_3877,RIdb83410_3878,RIdb81700_3879,RIdb7fa68_3880,RIdb7db78_3881,RIdb7bb98_3882,RIdb79e10_3883,RIdb78268_3884,
        RIdb76828_3885,RIdb746e0_3886,RIdda9490_3887,RIdda9c88_3888,RIddaa480_3889,RIddaac78_3890,RIddab470_3891,RIddabc68_3892,RIddac460_3893,RIddacc58_3894,
        RIddad450_3895,RIddadc48_3896,RIddae440_3897,RIddaec38_3898,RIddaf430_3899,RIddafc28_3900,RIddb0420_3901,RIddb0c18_3902,RIddb1410_3903,RIddb1c08_3904,
        RIddb2400_3905,RIddb2bf8_3906,RIddb33f0_3907,RIddb3be8_3908,RIddb43e0_3909,RIddb4bd8_3910,RIddb53d0_3911,RIddb5bc8_3912,RIddb63c0_3913,RIddb6bb8_3914,
        RIddb73b0_3915,RIddb7ba8_3916,RIddb83a0_3917,RIddb8b98_3918,RIddb9390_3919,RIddb9b88_3920,RIddba380_3921,RIddbab78_3922,RIddbb370_3923,RIddbbb68_3924,
        RIddbc360_3925,RIddbcb58_3926,RIddbd350_3927,RIddbdb48_3928,RIddbe340_3929,RIddbeb38_3930,RIddbf330_3931,RIddbfb28_3932,RIddc0320_3933,RIddc0b18_3934,
        RIddc1310_3935,RIddc1b08_3936,RIddc2300_3937,RIddc2af8_3938,RIddc32f0_3939,RIddc3ae8_3940,RIddc42e0_3941,RIddc4ad8_3942,RIddc52d0_3943,RIddc5ac8_3944,
        RIddc62c0_3945,RIddc6ab8_3946,RIddc72b0_3947,RIddc7aa8_3948,RIddc82a0_3949,RIddc8a98_3950,RIddc9290_3951,RIddc9a88_3952,RIddca280_3953,RIddcaa78_3954,
        RIddcb270_3955,RIddcba68_3956,RIddcc260_3957,RIddcca58_3958,RIddcd250_3959,RIddcda48_3960,RIddce240_3961,RIddcea38_3962,RIddcf230_3963,RIddcfa28_3964,
        RIddd0220_3965,RIddd0a18_3966,RIddd1210_3967,RIddd1a08_3968,RIdc0fbb8_3681,RIb86fc68_77,RIdc0f0f0_3682,RIb86fce0_76,RIdc0e5b0_3683,RIb86fd58_75,
        RIdc0dae8_3684,RIb87e8a8_74,RIdc0cfa8_3685,RIb87e920_73,RIdc0c3f0_3686,RIb87e998_72,RIdc0b7c0_3687,RIb87ea10_71,RIdc0ac08_3688,RIb87ea88_70,
        RIdc09f60_3689,RIdc093a8_3690,RIdc08700_3691,RIdc07878_3692,RIdc06270_3693,RIdc05118_3694,RIdc03b10_3695,RIdc029b8_3696,RIdc013b0_3697,RIdc00258_3698,
        RIdbff100_3699,RIdbfdaf8_3700,RIdbfc9a0_3701,RIdbfb398_3702,RIdbfa240_3703,RIdbf8c38_3704,RIdbf7ae0_3705,RIdbf6988_3706,RIdbf5380_3707,RIdbf4228_3708,
        RIdbf2c20_3709,RIdbf1ac8_3710,RIdbf04c0_3711,RIdbef368_3712,RIb79b428_272,RIdda31a8_3581,RIdbd9c48_3186,RIe036f80_4371,RIe100460_4766,RIda3bc30_2396,
        RIde6b9c8_3976,RIdb0e968_2791,RId987e10_2001,RIe527288_6346,RIe45e528_5951,RIe395df8_5556,RIe1ca840_5161,RId72b4a8_816,RIe5efc28_6741,RId8bc950_1606,
        RId7f4028_1211,RId710748_846,RId96d278_2032,RId8aa728_1632,RId7dcb80_1235,RIdbc4870_3212,RIdd8ba30_3609,RIda25c28_2423,RIdaf5f30_2820,RIe022a30_4393,
        RIe0e8ec8_4791,RIe1ac2a0_5191,RIe444fb0_5975,RIe37f9b8_5584,RIe5d6d40_6768,RIe5117a8_6369,RIe3ac2b0_6083,RIe3aaca8_6084,RIe3a9b50_6085,RIe3a8548_6086,
        RIe3a73f0_6087,RIe3a6298_6088,RIe3a4c90_6089,RIe3a3b38_6090,RIe3a2530_6091,RIe3a13d8_6092,RIe39fdd0_6093,RIe39ec78_6094,RIe39db20_6095,RIe39c518_6096,
        RIe1694d8_6097,RIe16e398_6098,RIe173270_6099,RIe178388_6100,RIe17c780_6101,RIe1805d8_6102,RIe1877c0_6103,RIe18c9c8_6104,RIe192ff8_6105,RIe198cc8_6106,
        RIe1a05b8_6107,RIe1a6300_6108,RIe1ac318_6109,RIe1b2420_6110,RIe1b7970_6111,RIe1bce48_6112,RIe1c12b8_6113,RIe1c7960_6114,RIe1cc820_6115,RIe1d0fd8_6116,
        RIe094940_6117,RIe090368_6118,RIe08b700_6119,RIe087a10_6120,RIe14c9f0_6121,RIe1495e8_6122,RIe146348_6123,RIe143210_6124,RIe140a38_6125,RIe13d4c8_6126,
        RIe13a660_6127,RIe137168_6128,RIe133a18_6129,RIe12fda0_6130,RIe1280f0_6131,RIe121b38_6132,RIe1194b0_6133,RIe1133a8_6134,RIe10ad20_6135,RIdfd70d0_6136,
        RIdff52b0_6137,RIe01ea70_6138,RIe03a5e0_6139,RIdfb6cb8_6140,RIdfa46d0_6141,RIdf7c7e8_6142,RIdc22218_6143,RIda953d8_6144,RIddeaf80_6145,RIde58a80_6146,
        RIe03fa40_6147,RIe04e338_6148,RIe0629f0_6149,RIe06c608_6150,RIe0732e0_6151,RIe07d0d8_6152,RIe084158_6153,RIdfc61e0_6154,RIe106838_6155,RIe0f8198_6156,
        RIe0eed00_6157,RIe0e2b68_6158,RIe0d0b98_6159,RIe0c3998_6160,RIe0b0960_6161,RIe0a6988_6162,RIe099440_6163,RIe1d3c60_6164,RIe1d69d8_6165,RIe1d9c00_6166,
        RIe1dc978_6167,RIe1dfba0_6168,RIe1e2918_6169,RIe1e5b40_6170,RIe1e88b8_6171,RIe1eb180_6172,RIe1ee858_6173,RIe1f1120_6174,RIe1f47f8_6175,RIe1f70c0_6176,
        RIe1fa180_6177,RIe1fbad0_6178,RIe1fd330_6179,RIe1ff568_6180,RIe2012f0_6181,RIe203000_6182,RIe203f00_6183,RIe2053a0_6184,RIe2066d8_6185,RIe207920_6186,
        RIe208be0_6187,RIe209d38_6188,RIe20b958_6189,RIe20cf60_6190,RIe20e4f0_6191,RIe20f5d0_6192,RIe211178_6193,RIe212c30_6194,RIe214148_6195,RIe215c00_6196,
        RIe217460_6197,RIe218798_6198,RIe2199e0_6199,RIe14e868_6200,RIe151130_6201,RIe153020_6202,RIe154ad8_6203,RIe156518_6204,RIe158228_6205,RIe15a280_6206,
        RIe15c3c8_6207,RIe15ef60_6208,RIe1616c0_6209,RIe164168_6210,RIe166c10_6211,RIe39a100_6212,RIe3984e0_6213,RIe3967d0_6214,RIe3941d8_6215,RIe391c58_6216,
        RIe38f5e8_6217,RIe38d428_6218,RIe38ae30_6219,RIe389030_6220,RIe386fd8_6221,RIe384ff8_6222,RIe3832e8_6223,RIe381218_6224,RIe37f148_6225,RIe37ce20_6226,
        RIe37aeb8_6227,RIe378668_6228,RIe3755a8_6229,RIe372c68_6230,RIe2703f8_6231,RIe26d4a0_6232,RIe26aae8_6233,RIe2686d0_6234,RIe265ca0_6235,RIe264170_6236,
        RIe2616c8_6237,RIe25f238_6238,RIe25c6a0_6239,RIe259ec8_6240,RIe257240_6241,RIe254018_6242,RIe251408_6243,RIe24e8e8_6244,RIe24c110_6245,RIe248d08_6246,
        RIe246170_6247,RIe2435d8_6248,RIe2418c8_6249,RIe23fb40_6250,RIe23dcc8_6251,RIe23ba18_6252,RIe239948_6253,RIe2381d8_6254,RIe236720_6255,RIe2346c8_6256,
        RIe232a30_6257,RIe230bb8_6258,RIe465cb0_6259,RIe4664a8_6260,RIe466ca0_6261,RIe467498_6262,RIe467c90_6263,RIe468488_6264,RIe468c80_6265,RIe469478_6266,
        RIe469c70_6267,RIe46a468_6268,RIe46ac60_6269,RIe46b458_6270,RIe46bc50_6271,RIe46c448_6272,RIe46cc40_6273,RIe46d438_6274,RIe46dc30_6275,RIe46e428_6276,
        RIe46ec20_6277,RIe46f418_6278,RIe46fc10_6279,RIe470408_6280,RIe470c00_6281,RIe4713f8_6282,RIe471bf0_6283,RIe4723e8_6284,RIe472bf8_6285,RIe4733f0_6286,
        RIe473be8_6287,RIe4743e0_6288,RIe474bd8_6289,RIe4753d0_6290,RIe475bc8_6291,RIe4763c0_6292,RIe476bb8_6293,RIe4773b0_6294,RIe477ba8_6295,RIe4783a0_6296,
        RIe478b98_6297,RIe479390_6298,RIe479b88_6299,RIe47a380_6300,RIe47ab78_6301,RIe47b370_6302,RIe47bb68_6303,RIe47c360_6304,RIe47cb58_6305,RIe47d350_6306,
        RIe47db48_6307,RIe47e340_6308,RIe47eb38_6309,RIe47f330_6310,RIe47fb28_6311,RIe480320_6312,RIe480b18_6313,RIe481310_6314,RIe481b08_6315,RIe482300_6316,
        RIe482af8_6317,RIe4832f0_6318,RIe483ae8_6319,RIe4842e0_6320,RIe484ad8_6321,RIe4852d0_6322,RIe485ac8_6323,RIe4862c0_6324,RIe486ab8_6325,RIe4872b0_6326,
        RIe487aa8_6327,RIe4882a0_6328,RIe488a98_6329,RIe489290_6330,RIe489a88_6331,RIe48a280_6332,RIe48aa78_6333,RIe48b270_6334,RIe48ba68_6335,RIe48c260_6336,
        RIe48ca58_6337,RIe48d250_6338,RIe3cd190_6051,RIe3cc3f8_6052,RIe3cb750_6053,RIe3ca9b8_6054,RIe3c9e00_6055,RIe3c9248_6056,RIe3c8708_6057,RIe3c7bc8_6058,
        RIe3c7100_6059,RIe3c6638_6060,RIe3c5af8_6061,RIe3c4ec8_6062,RIe3c4130_6063,RIe3c31b8_6064,RIe3c1bb0_6065,RIe3c0a58_6066,RIe3bf900_6067,RIe3be2f8_6068,
        RIe3bd1a0_6069,RIe3bbb98_6070,RIe3baa40_6071,RIe3b9438_6072,RIe3b82e0_6073,RIe3b7188_6074,RIe3b5b80_6075,RIe3b4a28_6076,RIe3b3420_6077,RIe3b22c8_6078,
        RIe3b0cc0_6079,RIe3afb68_6080,RIe3aea10_6081,RIe3ad408_6082,RIe51b690_6365,RIe500d68_6388,RIe501998_6387,RIe5026b8_6386,RIe5032e8_6385,RIe503f90_6384,
        RIe504d28_6383,RIe505958_6382,RIe50ef58_6371,RIe50ac50_6376,RIe50b880_6375,RIe50c690_6374,RIe50d428_6373,RIe524060_6351,RIe523688_6352,RIe524948_6350,
        RIe51d5f8_6362,RIe51c158_6364,RIe51cc20_6363,RIe51f290_6359,RIe51dee0_6361,RIe51e840_6360,RIe525410_6349,RIe525d70_6348,RIe5267c0_6347,RIe1e2210_5688,
        RIe1e10b8_5689,RIe1dfab0_5690,RIe1de958_5691,RIe1dd350_5692,RIe1dc1f8_5693,RIe1dabf0_5694,RIe1d9a98_5695,RIe1d8940_5696,RIe1d7338_5697,RIe1d61e0_5698,
        RIe1d4bd8_5699,RIe1d3a80_5700,RIe1d2478_5701,RIe099530_5702,RIe09d298_5703,RIe0a2338_5704,RIe0a6fa0_5705,RIe0ac310_5706,RIe0b16f8_5707,RIe0b9240_5708,
        RIe0bf438_5709,RIe0c4730_5710,RIe0cb0a8_5711,RIe0d0df0_5712,RIe0d8aa0_5713,RIe0de608_5714,RIe0e5ca0_5715,RIe0eb358_5716,RIe0ef138_5717,RIe0f3bc0_5718,
        RIe0f8300_5719,RIe0ff380_5720,RIe103430_5721,RIdfce868_5722,RIdfc9fc0_5723,RIdfc6000_5724,RIdfc1410_5725,RIdfbcc58_5726,RIe082f10_5727,RIe0800a8_5728,
        RIe07bd28_5729,RIe078ec0_5730,RIe075ab8_5731,RIe071f18_5732,RIe06f308_5733,RIe06b0f0_5734,RIe067928_5735,RIe0608a8_5736,RIe05a2f0_5737,RIe0541e8_5738,
        RIe04bb60_5739,RIe045a58_5740,RIe03d3d0_5741,RIde1d908_5742,RIde4a200_5743,RIde62e18_5744,RIdc30d68_5745,RIdde3e10_5746,RIddce948_5747,RIdb96b50_5748,
        RIda0b300_5749,RIdc00960_5750,RIdb708e8_5751,RIdc692d0_5752,RIdf7e930_5753,RIdf8d6d8_5754,RIdf9f978_5755,RIdfa6f20_5756,RIdfaf968_5757,RIdfb74b0_5758,
        RIddf5a98_5759,RIde028d8_5760,RIe036620_5761,RIe027530_5762,RIe01deb8_5763,RIe00b3a8_5764,RIdffd938_5765,RIdfefb08_5766,RIdfe0838_5767,RIdfd6680_5768,
        RIe1084d0_5769,RIe10ad98_5770,RIe10e470_5771,RIe110d38_5772,RIe113ab0_5773,RIe116cd8_5774,RIe119a50_5775,RIe11cc78_5776,RIe11f9f0_5777,RIe122c18_5778,
        RIe125990_5779,RIe128258_5780,RIe12b930_5781,RIe12e1f8_5782,RIe1308e0_5783,RIe132398_5784,RIe134300_5785,RIe135ae8_5786,RIe137258_5787,RIe138608_5788,
        RIe139850_5789,RIe13ab88_5790,RIe13c028_5791,RIe13d5b8_5792,RIe13ead0_5793,RIe13fef8_5794,RIe141230_5795,RIe142568_5796,RIe1434e0_5797,RIe144638_5798,
        RIe145880_5799,RIe146ac8_5800,RIe1486e8_5801,RIe149f48_5802,RIe14b550_5803,RIe14c978_5804,RIe14e430_5805,RIe0865e8_5806,RIe087f38_5807,RIe089db0_5808,
        RIe08b7f0_5809,RIe08d578_5810,RIe08f120_5811,RIe091100_5812,RIe093248_5813,RIe0950c0_5814,RIe096998_5815,RIe0986a8_5816,RIe1cfd18_5817,RIe1ce080_5818,
        RIe1cc550_5819,RIe1ca048_5820,RIe1c78e8_5821,RIe1c4f30_5822,RIe1c26e0_5823,RIe1c0b38_5824,RIe1be9f0_5825,RIe1bcce0_5826,RIe1baf58_5827,RIe1b9158_5828,
        RIe1b6908_5829,RIe1b3b90_5830,RIe1b1d18_5831,RIe1aff90_5832,RIe1ae2f8_5833,RIe1ab940_5834,RIe1a8628_5835,RIe1a6030_5836,RIe1a2d90_5837,RIe1a0540_5838,
        RIe19da20_5839,RIe19a870_5840,RIe197cd8_5841,RIe195410_5842,RIe192e90_5843,RIe190460_5844,RIe18e0c0_5845,RIe18bc30_5846,RIe189098_5847,RIe186c08_5848,
        RIe1839e0_5849,RIe1817a8_5850,RIe17fb88_5851,RIe17def0_5852,RIe17c3c0_5853,RIe17a458_5854,RIe1781a8_5855,RIe176240_5856,RIe174530_5857,RIe172988_5858,
        RIe16fc70_5859,RIe16e140_5860,RIe16c1d8_5861,RIe16a5b8_5862,RIe168a88_5863,RIe167138_5864,RIe39c680_5865,RIe39ce78_5866,RIe39d670_5867,RIe39de68_5868,
        RIe39e660_5869,RIe39ee58_5870,RIe39f650_5871,RIe39fe48_5872,RIe3a0640_5873,RIe3a0e38_5874,RIe3a1630_5875,RIe3a1e28_5876,RIe3a2620_5877,RIe3a2e18_5878,
        RIe3a3610_5879,RIe3a3e08_5880,RIe3a4600_5881,RIe3a4df8_5882,RIe3a55f0_5883,RIe3a5de8_5884,RIe3a65e0_5885,RIe3a6dd8_5886,RIe3a75d0_5887,RIe3a7dc8_5888,
        RIe3a85c0_5889,RIe3a8db8_5890,RIe3a95b0_5891,RIe3a9da8_5892,RIe3aa5a0_5893,RIe3aad98_5894,RIe3ab590_5895,RIe3abd88_5896,RIe3ac580_5897,RIe3acd78_5898,
        RIe3ad570_5899,RIe3add68_5900,RIe3ae560_5901,RIe3aed58_5902,RIe3af550_5903,RIe3afd48_5904,RIe3b0540_5905,RIe3b0d38_5906,RIe3b1530_5907,RIe3b1d28_5908,
        RIe3b2520_5909,RIe3b2d18_5910,RIe3b3510_5911,RIe3b3d08_5912,RIe3b4500_5913,RIe3b4cf8_5914,RIe3b54f0_5915,RIe3b5ce8_5916,RIe3b64e0_5917,RIe3b6cd8_5918,
        RIe3b74d0_5919,RIe3b7cc8_5920,RIe3b84c0_5921,RIe3b8cb8_5922,RIe3b94b0_5923,RIe3b9ca8_5924,RIe3ba4a0_5925,RIe3bac98_5926,RIe3bb490_5927,RIe3bbc88_5928,
        RIe3bc480_5929,RIe3bcc78_5930,RIe3bd470_5931,RIe3bdc68_5932,RIe3be460_5933,RIe3bec58_5934,RIe3bf450_5935,RIe3bfc48_5936,RIe3c0440_5937,RIe3c0c38_5938,
        RIe3c1430_5939,RIe3c1c28_5940,RIe3c2420_5941,RIe3c2c18_5942,RIe3c3410_5943,RIe202f10_5656,RIe202448_5657,RIe201980_5658,RIe200e40_5659,RIe2000a8_5660,
        RIe1ff310_5661,RIe1fe668_5662,RIe1fd9c0_5663,RIe1fce80_5664,RIe1fc340_5665,RIe1fb878_5666,RIe1facc0_5667,RIe1fa090_5668,RIe1f9118_5669,RIe1f7fc0_5670,
        RIe1f69b8_5671,RIe1f5860_5672,RIe1f4258_5673,RIe1f3100_5674,RIe1f1fa8_5675,RIe1f09a0_5676,RIe1ef848_5677,RIe1ee240_5678,RIe1ed0e8_5679,RIe1ebae0_5680,
        RIe1ea988_5681,RIe1e9830_5682,RIe1e8228_5683,RIe1e70d0_5684,RIe1e5ac8_5685,RIe1e4970_5686,RIe1e3368_5687,RIe4520c0_5970,RIe438440_5990,RIe4390e8_5989,
        RIe439f70_5988,RIe43ad80_5987,RIe43ba28_5986,RIe43c7c0_5985,RIe43d5d0_5984,RIe445e38_5974,RIe441c98_5979,RIe4429b8_5978,RIe443750_5977,RIe437630_5991,
        RIe455e28_5964,RIe454988_5966,RIe4554c8_5965,RIe45c278_5954,RIe45cdb8_5953,RIe45d880_5952,RIe45aec8_5956,RIe45a478_5957,RIe45b8a0_5955,RIe4534e8_5968,
        RIe452b88_5969,RIe453fb0_5967,RIe116b70_5293,RIe115a18_5294,RIe114410_5295,RIe1132b8_5296,RIe111cb0_5297,RIe110b58_5298,RIe10f550_5299,RIe10e3f8_5300,
        RIe10d2a0_5301,RIe10bc98_5302,RIe10ab40_5303,RIe109538_5304,RIe1083e0_5305,RIe106dd8_5306,RIdfd3728_5307,RIdfd71c0_5308,RIdfdc8f0_5309,RIdfe0b80_5310,
        RIdfe6760_5311,RIdfeb788_5312,RIdff1f98_5313,RIdff7f38_5314,RIdffe400_5315,RIe005750_5316,RIe00b420_5317,RIe0132b0_5318,RIe0193b8_5319,RIe0202d0_5320,
        RIe023de0_5321,RIe027878_5322,RIe02ccd8_5323,RIe0322a0_5324,RIe038768_5325,RIe03c728_5326,RIde01258_5327,RIddfd748_5328,RIddf9788_5329,RIddf3d88_5330,
        RIdfba228_5331,RIdfb5e30_5332,RIdfb2aa0_5333,RIdfaec48_5334,RIdfabf48_5335,RIdfa97e8_5336,RIdfa5e40_5337,RIdfa2f60_5338,RIdf9e4d8_5339,RIdf99618_5340,
        RIdf90f90_5341,RIdf8ae88_5342,RIdf848d0_5343,RIdf7c248_5344,RIdf76140_5345,RIdc56298_5346,RIdd75f50_5347,RIdd9d6b8_5348,RIdb67180_5349,RIdc198c0_5350,
        RIdc008e8_5351,RIdacdc88_5352,RId8fd180_5353,RIdb353b0_5354,RIdbdbca0_5355,RIdb8b8b8_5356,RIddb1a28_5357,RIddc60e0_5358,RIddd3cb8_5359,RIdddeaa0_5360,
        RIdde50d0_5361,RIddeee50_5362,RIdc2bb60_5363,RIdc34788_5364,RIde6e7b8_5365,RIde62ad0_5366,RIde55510_5367,RIde4a188_5368,RIde36d90_5369,RIde29c80_5370,
        RIde1c210_5371,RIde0cb08_5372,RIe03d4c0_5373,RIe040b98_5374,RIe043460_5375,RIe046b38_5376,RIe049400_5377,RIe04c178_5378,RIe04f3a0_5379,RIe052118_5380,
        RIe055340_5381,RIe0580b8_5382,RIe05b2e0_5383,RIe05e058_5384,RIe060920_5385,RIe063ff8_5386,RIe0662a8_5387,RIe068288_5388,RIe069a70_5389,RIe06b870_5390,
        RIe06cf68_5391,RIe06e6d8_5392,RIe06fa10_5393,RIe070eb0_5394,RIe0721e8_5395,RIe073808_5396,RIe074960_5397,RIe0762b0_5398,RIe0779a8_5399,RIe079118_5400,
        RIe07a798_5401,RIe07bcb0_5402,RIe07d768_5403,RIe07f220_5404,RIe080cd8_5405,RIe082088_5406,RIe083078_5407,RIe0843b0_5408,RIdfbbbf0_5409,RIdfbd5b8_5410,
        RIdfbf3b8_5411,RIdfc15f0_5412,RIdfc30a8_5413,RIdfc4f20_5414,RIdfc6f00_5415,RIdfc85f8_5416,RIdfca3f8_5417,RIdfcc720_5418,RIdfce8e0_5419,RIe106478_5420,
        RIe104948_5421,RIe102b48_5422,RIe100f28_5423,RIe0fea20_5424,RIe0fcd10_5425,RIe0fa3d0_5426,RIe0f7838_5427,RIe0f5a38_5428,RIe0f3968_5429,RIe0f1b68_5430,
        RIe0f0290_5431,RIe0ee508_5432,RIe0ec690_5433,RIe0eaea8_5434,RIe0e8658_5435,RIe0e54a8_5436,RIe0e2988_5437,RIe0e0228_5438,RIe0dd7f8_5439,RIe0da828_5440,
        RIe0d7f60_5441,RIe0d4f18_5442,RIe0d3280_5443,RIe0d02b0_5444,RIe0cdad8_5445,RIe0cae50_5446,RIe0c8150_5447,RIe0c5d38_5448,RIe0c3290_5449,RIe0c0d88_5450,
        RIe0be628_5451,RIe0bbdd8_5452,RIe0b91c8_5453,RIe0b5f28_5454,RIe0b3318_5455,RIe0b02d0_5456,RIe0adeb8_5457,RIe0ac0b8_5458,RIe0aa330_5459,RIe0a83c8_5460,
        RIe0a6a00_5461,RIe0a40c0_5462,RIe0a2158_5463,RIe0a0010_5464,RIe09e378_5465,RIe09c668_5466,RIe09a8e0_5467,RIe099080_5468,RIe1d1cf8_5469,RIe1d24f0_5470,
        RIe1d2ce8_5471,RIe1d34e0_5472,RIe1d3cd8_5473,RIe1d44d0_5474,RIe1d4cc8_5475,RIe1d54c0_5476,RIe1d5cb8_5477,RIe1d64b0_5478,RIe1d6ca8_5479,RIe1d74a0_5480,
        RIe1d7c98_5481,RIe1d8490_5482,RIe1d8c88_5483,RIe1d9480_5484,RIe1d9c78_5485,RIe1da470_5486,RIe1dac68_5487,RIe1db460_5488,RIe1dbc58_5489,RIe1dc450_5490,
        RIe1dcc48_5491,RIe1dd440_5492,RIe1ddc38_5493,RIe1de430_5494,RIe1dec28_5495,RIe1df420_5496,RIe1dfc18_5497,RIe1e0410_5498,RIe1e0c08_5499,RIe1e1400_5500,
        RIe1e1bf8_5501,RIe1e23f0_5502,RIe1e2be8_5503,RIe1e33e0_5504,RIe1e3bd8_5505,RIe1e43d0_5506,RIe1e4bc8_5507,RIe1e53c0_5508,RIe1e5bb8_5509,RIe1e63b0_5510,
        RIe1e6ba8_5511,RIe1e73a0_5512,RIe1e7b98_5513,RIe1e8390_5514,RIe1e8b88_5515,RIe1e9380_5516,RIe1e9b78_5517,RIe1ea370_5518,RIe1eab68_5519,RIe1eb360_5520,
        RIe1ebb58_5521,RIe1ec350_5522,RIe1ecb48_5523,RIe1ed340_5524,RIe1edb38_5525,RIe1ee330_5526,RIe1eeb28_5527,RIe1ef320_5528,RIe1efb18_5529,RIe1f0310_5530,
        RIe1f0b08_5531,RIe1f1300_5532,RIe1f1af8_5533,RIe1f22f0_5534,RIe1f2ae8_5535,RIe1f32e0_5536,RIe1f3ad8_5537,RIe1f42d0_5538,RIe1f4ac8_5539,RIe1f52c0_5540,
        RIe1f5ab8_5541,RIe1f62b0_5542,RIe1f6aa8_5543,RIe1f72a0_5544,RIe1f7a98_5545,RIe1f8290_5546,RIe1f8a88_5547,RIe1f9280_5548,RIe137870_5261,RIe136da8_5262,
        RIe136358_5263,RIe135890_5264,RIe134d50_5265,RIe134288_5266,RIe1337c0_5267,RIe132c08_5268,RIe131fd8_5269,RIe1313a8_5270,RIe1307f0_5271,RIe12fbc0_5272,
        RIe12f080_5273,RIe12da78_5274,RIe12c920_5275,RIe12b318_5276,RIe12a1c0_5277,RIe128bb8_5278,RIe127a60_5279,RIe126908_5280,RIe125300_5281,RIe1241a8_5282,
        RIe122ba0_5283,RIe121a48_5284,RIe120440_5285,RIe11f2e8_5286,RIe11e190_5287,RIe11cb88_5288,RIe11ba30_5289,RIe11a428_5290,RIe1192d0_5291,RIe117cc8_5292,
        RIe38a110_5575,RIe378410_5590,RIe379220_5589,RIe379e50_5588,RIe26f4f8_5601,RIe270290_5600,RIe270ec0_5599,RIe271be0_5598,RIe37b908_5586,RIe375008_5594,
        RIe375da0_5593,RIe376a48_5592,RIe377768_5591,RIe392b58_5561,RIe3921f8_5562,RIe3934b8_5560,RIe38b9e8_5572,RIe38a908_5574,RIe38b1f0_5573,RIe38da40_5569,
        RIe38c4b0_5571,RIe38cf78_5570,RIe393e90_5559,RIe394868_5558,RIe3951c8_5557,RIe04cad8_4898,RIe04b980_4899,RIe04a378_4900,RIe049220_4901,RIe047c18_4902,
        RIe046ac0_4903,RIe045968_4904,RIe044360_4905,RIe043208_4906,RIe041c00_4907,RIe040aa8_4908,RIe03f4a0_4909,RIe03e348_4910,RIe03d1f0_4911,RIde08bc0_4912,
        RIde0d030_4913,RIde131b0_4914,RIde17968_4915,RIde1f528_4916,RIde24e38_4917,RIde29ed8_4918,RIde31390_4919,RIde36e08_4920,RIde3efe0_4921,RIde45070_4922,
        RIde4c9d8_4923,RIde51b68_4924,RIde553a8_4925,RIde59c50_4926,RIde5e390_4927,RIde65668_4928,RIde6a4b0_4929,RIde6f820_4930,RIdf73710_4931,RIdc38040_4932,
        RIdc32b68_4933,RIdc2ee78_4934,RIdc29bf8_4935,RIddf1628_4936,RIddee388_4937,RIddeaa58_4938,RIdde7a88_4939,RIdde35a0_4940,RIdde0cd8_4941,RIddddf60_4942,
        RIdddb710_4943,RIddd5e78_4944,RIddd2278_4945,RIddcc080_4946,RIddc39f8_4947,RIddbd8f0_4948,RIddb5268_4949,RIddaf160_4950,RIdb7c228_4951,RIdb96c40_4952,
        RIdbbbd38_4953,RIdbdcdf8_4954,RIdb5db80_4955,RIdb48190_4956,RIdb26ba8_4957,RId917aa8_4958,RId986da8_4959,RIda7eb60_4960,RIdaf90e0_4961,RIdab27a8_4962,
        RIdbf1ca8_4963,RIdc00a50_4964,RIdc0fe88_4965,RIdc16080_4966,RIdc1c098_4967,RIdc25080_4968,RIdb67810_4969,RIdda8518_4970,RIdd9d5c8_4971,RIdd8f270_4972,
        RIdd82fe8_4973,RIdd74150_4974,RIdc641b8_4975,RIdc54600_4976,RIdc46848_4977,RIdc3b970_4978,RIdf77220_4979,RIdf79f98_4980,RIdf7c860_4981,RIdf7ff38_4982,
        RIdf82800_4983,RIdf85ed8_4984,RIdf887a0_4985,RIdf8be78_4986,RIdf8e740_4987,RIdf91008_4988,RIdf946e0_4989,RIdf96fa8_4990,RIdf9a680_4991,RIdf9ccf0_4992,
        RIdf9ec58_4993,RIdfa04b8_4994,RIdfa1bb0_4995,RIdfa3b18_4996,RIdfa4dd8_4997,RIdfa6110_4998,RIdfa75b0_4999,RIdfa88e8_5000,RIdfa9d10_5001,RIdfab048_5002,
        RIdfac218_5003,RIdfad460_5004,RIdfaecc0_5005,RIdfb0610_5006,RIdfb1c90_5007,RIdfb3310_5008,RIdfb4828_5009,RIdfb5d40_5010,RIdfb77f8_5011,RIdfb92b0_5012,
        RIdfba9a8_5013,RIddf2ca8_5014,RIddf4580_5015,RIddf6308_5016,RIddf8270_5017,RIddf9e90_5018,RIddfbdf8_5019,RIddfdb08_5020,RIddff548_5021,RIde015a0_5022,
        RIde03508_5023,RIde04fc0_5024,RIe03bbe8_5025,RIe039cf8_5026,RIe038600_5027,RIe0363c8_5028,RIe033b78_5029,RIe031580_5030,RIe02ee98_5031,RIe02c4e0_5032,
        RIe02a488_5033,RIe028958_5034,RIe026b58_5035,RIe025460_5036,RIe023b88_5037,RIe021fe0_5038,RIe020168_5039,RIe01dcd8_5040,RIe01b758_5041,RIe018440_5042,
        RIe0157b8_5043,RIe012590_5044,RIe010628_5045,RIe00d298_5046,RIe00a778_5047,RIe007e38_5048,RIe004df0_5049,RIe0024b0_5050,RIdfff558_5051,RIdffcd08_5052,
        RIdffa260_5053,RIdff7b78_5054,RIdff4f68_5055,RIdff1ea8_5056,R_25610_96cc360,R_25642_95f0d48,R_25644_9598060,R_25646_95984f8,R_25614_953c348,R_25616_96251f8,
        R_25618_96ed6b0,R_2561a_95f00d0,R_2561c_95f0418,R_2561e_95f0760,R_25620_953c3f0,R_25622_953c690,R_25612_953c9d8,R_25624_95f08b0,R_25626_953ca80,R_25628_96253f0,
        R_2562a_9632be8,R_253fc_9d20ef0,R_25412_9530108,R_25428_95f75a0,R_2543e_95301b0,R_25454_95304f8,R_2546a_9533198,R_25474_95332e8,R_25476_96dee60,R_25478_95f7798,
        R_2547a_96def08,R_253fe_95f7990,R_25400_9d21190,R_25402_9d21388,R_25404_9589e90,R_25406_9d21430,R_25408_9533780,R_2540a_9533b70,R_2540c_9d216d0,R_2540e_958a5c8,
        R_25410_96defb0,R_25414_9d21778,R_25416_9d21cb8,R_25418_95f7ae0,R_2541a_9d21d60,R_2541c_96df100,R_2541e_9d221f8,R_25420_958ac58,R_25422_95f7b88,R_25424_9533c18,
        R_25426_958b630,R_2542a_9d222a0,R_2542c_9533d68,R_2542e_95f7c30,R_25430_9d22498,R_25432_9d22540,R_25434_9533f60,R_25436_96df1a8,R_25438_95f7f78,R_2543a_9534008,
        R_2543c_9534200,R_25440_95f80c8,R_25442_96df250,R_25444_9d22690,R_25446_95fa438,R_25448_95fa4e0,R_2544a_958bcc0,R_2544c_9d22738,R_2544e_9d227e0,R_25450_9d22888,
        R_25452_9d22930,R_25456_9d229d8,R_25458_95fa588,R_2545a_9534350,R_2545c_95fa828,R_2545e_9d22a80,R_25460_96df2f8,R_25462_96df3a0,R_25464_95343f8,R_25466_95fa8d0,
        R_25468_95faac8,R_2546c_958bd68,R_2546e_958be10,R_25470_95fab70,R_25472_9d22b28,R_2547c_958beb8,R_25492_9d22bd0,R_254a8_958bf60,R_254be_9d22c78,R_254d4_9d22dc8,
        R_254ea_9d22e70,R_254f4_958c0b0,R_254f6_9d22f18,R_254f8_958c158,R_254fa_9d22fc0,R_2547e_958c200,R_25480_9d23068,R_25482_9d231b8,R_25484_958c2a8,R_25486_958c350,
        R_25488_9d23458,R_2548a_958c4a0,R_2548c_9d235a8,R_2548e_9d236f8,R_25490_958c548,R_25494_958c5f0,R_25496_9d237a0,R_25498_958c698,R_2549a_958f728,R_2549c_9d23848,
        R_2549e_958f7d0,R_254a0_958f878,R_254a2_9d23998,R_254a4_9d23ae8,R_254a6_9d23c38,R_254aa_9d23d88,R_254ac_9d23e30,R_254ae_9d23f80,R_254b0_9d24028,R_254b2_9d240d0,
        R_254b4_9d24220,R_254b6_9d242c8,R_254b8_9590988,R_254ba_9590a30,R_254bc_9590cd0,R_254c0_9d24418,R_254c2_9590d78,R_254c4_9590f70,R_254c6_9591178,R_254c8_9d24568,
        R_254ca_9d24bf8,R_254cc_9d25090,R_254ce_95916b8,R_254d0_9591808,R_254d2_9d251e0,R_254d6_9d25f10,R_254d8_9d25fb8,R_254da_95918b0,R_254dc_9d265a0,R_254de_9591958,
        R_254e0_9d26990,R_254e2_9d26c30,R_254e4_9591a00,R_254e6_95347e8,R_254e8_9591b50,R_254ec_9591bf8,R_254ee_9d26d80,R_254f0_9d27368,R_254f2_9d27410,R_254fc_96df4f0,
        R_25512_9d276b0,R_25528_96df598,R_2553e_9534890,R_25554_9d27c98,R_2556a_96df640,R_25574_9d27de8,R_25576_96df6e8,R_25578_9534bd8,R_2557a_96df838,R_254fe_96dfad8,
        R_25500_9534d28,R_25502_9534dd0,R_25504_9534f20,R_25506_9d281d8,R_25508_96dfb80,R_2550a_9d28328,R_2550c_9d283d0,R_2550e_96dfc28,R_25510_9534fc8,R_25514_96dfcd0,
        R_25516_9d28520,R_25518_96dfe20,R_2551a_96dfec8,R_2551c_9535070,R_2551e_95351c0,R_25520_9535268,R_25522_96dff70,R_25524_96e0018,R_25526_96e00c0,R_2552a_9535310,
        R_2552c_96e0168,R_2552e_96e0210,R_25530_96e02b8,R_25532_96e0408,R_25534_96e0558,R_25536_96e0600,R_25538_9535658,R_2553a_9d289b8,R_2553c_96e06a8,R_25540_95358f8,
        R_25542_96e0750,R_25544_96e0b40,R_25546_96e0be8,R_25548_96e0c90,R_2554a_96e0d38,R_2554c_95359a0,R_2554e_9d28a60,R_25550_96e0e88,R_25552_9535a48,R_25556_96e0f30,
        R_25558_9535b98,R_2555a_9d28c58,R_2555c_96e0fd8,R_2555e_9d28d00,R_25560_9535c40,R_25562_95362d0,R_25564_9536810,R_25566_9536a08,R_25568_96e1080,R_2556c_96e1128,
        R_2556e_9d28ef8,R_25570_96e11d0,R_25572_96e1c50,R_2557c_9591d48,R_25592_9591df0,R_255a8_96e2e08,R_255be_9591e98,R_255d4_9591f40,R_255ea_96e3690,R_255f4_96e6918,
        R_255f6_96e69c0,R_255f8_9d29048,R_255fa_9d28718,R_2557e_9591fe8,R_25580_96e6fa8,R_25582_96e72f0,R_25584_9d287c0,R_25586_9592090,R_25588_9592138,R_2558a_96e7398,
        R_2558c_9d28868,R_2558e_9d290f0,R_25590_9d29240,R_25594_96e7cc8,R_25596_95921e0,R_25598_9592288,R_2559a_9592330,R_2559c_96e82b0,R_2559e_9d292e8,R_255a0_9d2dfb0,
        R_255a2_9592528,R_255a4_9592678,R_255a6_9d2e058,R_255aa_96e8358,R_255ac_9592918,R_255ae_96e86a0,R_255b0_9d2e988,R_255b2_9d29390,R_255b4_9d2ec28,R_255b6_9d294e0,
        R_255b8_9d2f360,R_255ba_9592a68,R_255bc_9592b10,R_255c0_9d30128,R_255c2_9592c60,R_255c4_96e8940,R_255c6_96e89e8,R_255c8_9d30278,R_255ca_96e8be0,R_255cc_9592f00,
        R_255ce_9d29588,R_255d0_9d296d8,R_255d2_9d30518,R_255d6_9d29828,R_255d8_96e9120,R_255da_96e93c0,R_255dc_96e9510,R_255de_9d307b8,R_255e0_9d29cc0,R_255e2_9592fa8,
        R_255e4_9593050,R_255e6_96e9858,R_255e8_96e9a50,R_255ec_95930f8,R_255ee_9d29eb8,R_255f0_96ea038,R_255f2_95931a0,R_253bc_96eacb0,R_253be_9593248,R_253c0_9d29f60,
        R_253c2_95932f0,R_253c4_96eae00,R_253c6_9536b58,R_253c8_9593398,R_253ca_9d2a350,R_253cc_b7dc210,R_253ce_b7dcd38,R_253d0_b7dcde0,R_253d2_9593590,R_253d4_96376b8,
        R_253d6_9d2a4a0,R_253d8_9596038,R_253da_b7dc2b8,R_253dc_96eb0a0,R_253de_9596578,R_253e0_9536f48,R_253e2_96eb298,R_253e4_9537098,R_253e6_96eb340,R_253e8_95373e0,
        R_253ea_9596a10,R_253ec_9d30860,R_253ee_9ef0090,R_253f0_9d30f98,R_253f2_9ef05d0,R_253f4_9d31040,R_253f6_9d31238,R_253f8_9d314d8,R_253fa_9d316d0,R_25666_96346d0,
        R_1a4_b821b50,R_1a3_b821aa8,R_23ca4_96329f0,R_23cba_9f596e0,R_23cd0_962b7c0,R_23ce6_955f268,R_23cfc_9f5c4d0,R_23d12_9d225e8,R_23d1c_962b910,R_23d1e_95a3470,
        R_23d20_9632c90,R_23d22_95a3710,R_23ca6_9ee76c0,R_23ca8_9ee7810,R_23caa_9ee78b8,R_23cac_9ee8140,R_23cae_962bbb0,R_23cb0_9ee8920,R_23cb2_9d22d20,R_23cb4_9ee8bc0,
        R_23cb6_9632d38,R_23cb8_9d23110,R_23cbc_962bc58,R_23cbe_9ee9ad8,R_23cc0_9d23260,R_23cc2_9632f30,R_23cc4_9eec430,R_23cc6_9d23308,R_23cc8_9eef4c0,R_23cca_9eefca0,
        R_23ccc_9d23650,R_23cce_9ef0678,R_23cd2_95a3908,R_23cd4_962bd00,R_23cd6_9632fd8,R_23cd8_962be50,R_23cda_96331d0,R_23cdc_962bef8,R_23cde_9d30ef0,R_23ce0_9d238f0,
        R_23ce2_9d23b90,R_23ce4_962bfa0,R_23ce8_962c048,R_23cea_95a3a58,R_23cec_9d23ed8,R_23cee_9ef09c0,R_23cf0_9ef4380,R_23cf2_95a3ba8,R_23cf4_9ef4a10,R_23cf6_962c0f0,
        R_23cf8_96c3060,R_23cfa_96c6d68,R_23cfe_9d310e8,R_23d00_96c72a8,R_23d02_962c390,R_23d04_96c74a0,R_23d06_962da88,R_23d08_9d24178,R_23d0a_962df20,R_23d0c_9633278,
        R_23d0e_9633320,R_23d10_95a3e48,R_23d14_95a4040,R_23d16_9d24370,R_23d18_96c7e78,R_23d1a_96333c8,R_23d24_9633470,R_23d3a_9633518,R_23d50_962dfc8,R_23d66_9629b88,
        R_23d7c_95547c8,R_23d92_96335c0,R_23d9c_96337b8,R_23d9e_9633908,R_23da0_9633a58,R_23da2_962e7a8,R_23d26_9554870,R_23d28_962a560,R_23d2a_962ee38,R_23d2c_962a8a8,
        R_23d2e_962f2d0,R_23d30_95549c0,R_23d32_9633cf8,R_23d34_962f4c8,R_23d36_9633da0,R_23d38_9633e48,R_23d3c_9633ef0,R_23d3e_962c4e0,R_23d40_9554bb8,R_23d42_9554d08,
        R_23d44_9634040,R_23d46_962f6c0,R_23d48_9554f00,R_23d4a_962c8d0,R_23d4c_9635000,R_23d4e_962fab0,R_23d52_95552f0,R_23d54_96350a8,R_23d56_96351f8,R_23d58_962fc00,
        R_23d5a_95554e8,R_23d5c_9555638,R_23d5e_9635540,R_23d60_96355e8,R_23d62_9635738,R_23d64_96359d8,R_23d68_962ca20,R_23d6a_9635f18,R_23d6c_962ff48,R_23d6e_9636068,
        R_23d70_96363b0,R_23d72_9636ae8,R_23d74_9637220,R_23d76_9637e98,R_23d78_9638b10,R_23d7a_962d4a0,R_23d7e_96305d8,R_23d80_9638bb8,R_23d82_9638fa8,R_23d84_962d548,
        R_23d86_9639398,R_23d88_95556e0,R_23d8a_9639440,R_23d8c_9d18d00,R_23d8e_9d19d68,R_23d90_9630a70,R_23d94_9d1a008,R_23d96_9d1a350,R_23d98_9d1a9e0,R_23d9a_96314f0,
        R_23da4_9634430,R_23dba_95558d8,R_23dd0_9555a28,R_23de6_9d1ac80,R_23dfc_962d9e0,R_23e12_9555b78,R_23e1c_96344d8,R_23e1e_9555e18,R_23e20_9d1b070,R_23e22_9d1b8f8,
        R_23da6_9634a18,R_23da8_9555f68,R_23daa_9635150,R_23dac_96352a0,R_23dae_9556010,R_23db0_9557078,R_23db2_96353f0,R_23db4_9d1ba48,R_23db6_962db30,R_23db8_96357e0,
        R_23dbc_9559730,R_23dbe_955bde8,R_23dc0_955dd68,R_23dc2_9d1baf0,R_23dc4_955e158,R_23dc6_9638db0,R_23dc8_9d1bb98,R_23dca_9639248,R_23dcc_9d1bce8,R_23dce_96c81c0,
        R_23dd2_955e4a0,R_23dd4_955ea88,R_23dd6_96392f0,R_23dd8_9d15d18,R_23dda_955ee78,R_23ddc_9d168e8,R_23dde_9d16ae0,R_23de0_962e310,R_23de2_9d16c30,R_23de4_9d16e28,
        R_23de8_9d170c8,R_23dea_955f1c0,R_23dec_96c87a8,R_23dee_955f310,R_23df0_9d1bee0,R_23df2_955f3b8,R_23df4_95a39b0,R_23df6_96c8af0,R_23df8_95a3b00,R_23dfa_95a40e8,
        R_23dfe_95a44d8,R_23e00_9d1bf88,R_23e02_95a4580,R_23e04_95a4c10,R_23e06_9d17218,R_23e08_95a5348,R_23e0a_962ec40,R_23e0c_9d17608,R_23e0e_95a57e0,R_23e10_95a5930,
        R_23e14_9d18910,R_23e16_9d19630,R_23e18_95a5c78,R_23e1a_95a6260,R_23e24_9d1c030,R_23e3a_95a4628,R_23e50_95a48c8,R_23e66_95a4b68,R_23e7c_95b1438,R_23e92_9d19780,
        R_23e9c_95a6d88,R_23e9e_95b1780,R_23ea0_95a7028,R_23ea2_95a70d0,R_23e26_95b1828,R_23e28_95a7220,R_23e2a_95b2bd8,R_23e2c_95b3310,R_23e2e_95818b0,R_23e30_9582138,
        R_23e32_9582288,R_23e34_95a7760,R_23e36_9582870,R_23e38_95a78b0,R_23e3c_9d1c0d8,R_23e3e_9582a68,R_23e40_9d1b118,R_23e42_9582e58,R_23e44_9582f00,R_23e46_95830f8,
        R_23e48_958cbd8,R_23e4a_958cc80,R_23e4c_95a7aa8,R_23e4e_958f5d8,R_23e52_958f920,R_23e54_9590058,R_23e56_95a7bf8,R_23e58_95a7ca0,R_23e5a_95901a8,R_23e5c_959fdb8,
        R_23e5e_95a0b80,R_23e60_9d1c4c8,R_23e62_9625b28,R_23e64_96261b8,R_23e68_9d1b268,R_23e6a_9d1c570,R_23e6c_95a7d48,R_23e6e_9626458,R_23e70_95a8090,R_23e72_9628330,
        R_23e74_9628480,R_23e76_9628528,R_23e78_95a8138,R_23e7a_96285d0,R_23e7e_9628720,R_23e80_9628bb8,R_23e82_962c198,R_23e84_9d1c618,R_23e86_95a8288,R_23e88_9634238,
        R_23e8a_9d1c6c0,R_23e8c_96342e0,R_23e8e_9634970,R_23e90_9d1c8b8,R_23e94_9639830,R_23e96_9d159d0,R_23e98_9d15e68,R_23e9a_95a83d8,R_23c64_96c9a08,R_23c66_9d1b658,
        R_23c68_96ca920,R_23c6a_9d244c0,R_23c6c_96cb4f0,R_23c6e_9d1b700,R_23c70_9d1ca08,R_23c72_96cb640,R_23c74_962f030,R_23c76_9d1cc00,R_23c78_9d1cd50,R_23c7a_9d1cdf8,
        R_23c7c_9d1b7a8,R_23c7e_9d1cf48,R_23c80_9d1d098,R_23c82_9d1d1e8,R_23c84_95a8528,R_23c86_9d1b9a0,R_23c88_95a8720,R_23c8a_9d1be38,R_23c8c_9d246b8,R_23c8e_96cb838,
        R_23c90_9d24760,R_23c92_9d1c2d0,R_23c94_9d1d3e0,R_23c96_95a87c8,R_23c98_9d19438,R_23c9a_9d1c378,R_23c9c_9d1c768,R_23c9e_9d1d488,R_23ca0_9d1c960,R_23ca2_9d1e8e0,
        R_23ebc_9667ae0,R_23ebe_965f6f8,R_23ec0_9667b88,R_23ec2_96688a8,R_23ec4_95ac230,R_23ec6_95ac428,R_23ec8_966a780,R_23eca_966a8d0,R_23eba_965f8f0,R_23ecc_95ac620,
        R_23ece_95ac770,R_23ed0_966a978,R_23ed2_966aa20,R_23eb8_966aac8,R_23eea_95b1588,R_23eec_9d1e448,R_23eee_9d1e790,R_23a0c_95b1630,R_23a22_95b1c18,R_23a38_966acc0,
        R_23a4e_95b1d68,R_23a64_966ad68,R_23a7a_95b2c80,R_23a84_9661a68,R_23a86_9d1d7d0,R_23a88_966ae10,R_23a8a_966b0b0,R_23a0e_962f420,R_23a10_966ba88,R_23a12_95b2fc8,
        R_23a14_9d1f6a8,R_23a16_952daf8,R_23a18_95b3268,R_23a1a_9581220,R_23a1c_9d1d878,R_23a1e_9663160,R_23a20_9d1e250,R_23a24_9d1fb40,R_23a26_95305a0,R_23a28_95812c8,
        R_23a2a_9530798,R_23a2c_95816b8,R_23a2e_9663550,R_23a30_9531e90,R_23a32_9531f38,R_23a34_9532130,R_23a36_9532280,R_23a3a_9532328,R_23a3c_9581760,R_23a3e_9581f40,
        R_23a40_95323d0,R_23a42_9532868,R_23a44_9582720,R_23a46_9532b08,R_23a48_9532c58,R_23a4a_9582918,R_23a4c_966a4e0,R_23a50_9532e50,R_23a52_9d24808,R_23a54_9533390,
        R_23a56_9d20668,R_23a58_9582db0,R_23a5a_9583050,R_23a5c_9533978,R_23a5e_9534158,R_23a60_9d20710,R_23a62_95349e0,R_23a66_9537290,R_23a68_9d1f750,R_23a6a_966a6d8,
        R_23a6c_966aeb8,R_23a6e_966b158,R_23a70_9537a70,R_23a72_9539f30,R_23a74_95831a0,R_23a76_9537c68,R_23a78_9d20a58,R_23a7c_9537d10,R_23a7e_9537e60,R_23a80_9538250,
        R_23a82_95382f8,R_23a8c_9d21e08,R_23aa2_9583440,R_23ab8_9d1f8a0,R_23ace_9d1ff30,R_23ae4_9d23ce0,R_23afa_95834e8,R_23b04_9583590,R_23b06_9d20860,R_23b08_9d24958,
        R_23b0a_9d24ca0,R_23a8e_95836e0,R_23a90_9583e18,R_23a92_9d25288,R_23a94_9d20908,R_23a96_9d25330,R_23a98_9d22348,R_23a9a_9d253d8,R_23a9c_9d233b0,R_23a9e_9d25528,
        R_23aa0_9d255d0,R_23aa4_9d23500,R_23aa6_9d25678,R_23aa8_9d23a40,R_23aaa_9d24610,R_23aac_9d25880,R_23aae_9d248b0,R_23ab0_9d26258,R_23ab2_9584898,R_23ab4_9d24a00,
        R_23ab6_9d26450,R_23aba_9d26648,R_23abc_9d26e28,R_23abe_9d270c8,R_23ac0_9584c88,R_23ac2_9d24aa8,R_23ac4_9d24d48,R_23ac6_9585270,R_23ac8_9585708,R_23aca_9d27bf0,
        R_23acc_9d28910,R_23ad0_9d29198,R_23ad2_9d29630,R_23ad4_9d24fe8,R_23ad6_95857b0,R_23ad8_9d2a0b0,R_23ada_9585900,R_23adc_9d2a200,R_23ade_9d2a3f8,R_23ae0_9d2a7e8,
        R_23ae2_9d25138,R_23ae6_9d2ad28,R_23ae8_95860e0,R_23aea_9d25480,R_23aec_9d25928,R_23aee_9d25bc8,R_23af0_95864d0,R_23af2_9d25e68,R_23af4_95866c8,R_23af6_9586770,
        R_23af8_9587688,R_23afc_9d26ed0,R_23afe_9587730,R_23b00_9d27aa0,R_23b02_9d2add0,R_23b0c_95877d8,R_23b22_95386e8,R_23b38_95388e0,R_23b4e_9588108,R_23b64_9538ad8,
        R_23b7a_9d2b118,R_23b84_95881b0,R_23b86_95899f8,R_23b88_9589aa0,R_23b8a_9d2b460,R_23b0e_958d268,R_23b10_95390c0,R_23b12_9539168,R_23b14_95394b0,R_23b16_95399f0,
        R_23b18_9539c90,R_23b1a_953ba18,R_23b1c_953bac0,R_23b1e_958d460,R_23b20_9d2b508,R_23b24_953bf58,R_23b26_953c0a8,R_23b28_953c1f8,R_23b2a_953c540,R_23b2c_9d2b5b0,
        R_23b2e_953c888,R_23b30_953cdc8,R_23b32_958da48,R_23b34_9d2b700,R_23b36_953cf18,R_23b3a_958de38,R_23b3c_958e180,R_23b3e_96ddca8,R_23b40_96dddf8,R_23b42_958e570,
        R_23b44_958e810,R_23b46_96de098,R_23b48_9d285c8,R_23b4a_96de3e0,R_23b4c_9d28b08,R_23b50_96de530,R_23b52_958ef48,R_23b54_9d24b50,R_23b56_9d25d18,R_23b58_958ff08,
        R_23b5a_96e6c60,R_23b5c_96e8160,R_23b5e_96ebc70,R_23b60_95903a0,R_23b62_95906e8,R_23b66_96ebdc0,R_23b68_95efb90,R_23b6a_9596d58,R_23b6c_9d2b7a8,R_23b6e_9598c30,
        R_23b70_95f0220,R_23b72_9598cd8,R_23b74_95f1918,R_23b76_9599170,R_23b78_9d28bb0,R_23b7c_95f37f0,R_23b7e_95f41c8,R_23b80_95f4318,R_23b82_95992c0,R_23b8c_9599608,
        R_23ba2_9599758,R_23bb8_9599800,R_23bce_9599950,R_23be4_962f570,R_23bfa_9599b48,R_23c04_959a088,R_23c06_959a130,R_23c08_959a1d8,R_23c0a_962f618,R_23b8e_959a5c8,
        R_23b90_959a9b8,R_23b92_959ac58,R_23b94_959aef8,R_23b96_962f8b8,R_23b98_959afa0,R_23b9a_959b048,R_23b9c_959b0f0,R_23b9e_959b198,R_23ba0_959b240,R_23ba4_959b6d8,
        R_23ba6_959b828,R_23ba8_959b8d0,R_23baa_959ba20,R_23bac_9d28da8,R_23bae_959bac8,R_23bb0_959d268,R_23bb2_959d508,R_23bb4_959dce8,R_23bb6_959e420,R_23bba_9d28fa0,
        R_23bbc_962f960,R_23bbe_9d298d0,R_23bc0_959e618,R_23bc2_959eea0,R_23bc4_959f098,R_23bc6_9d29978,R_23bc8_9d25dc0,R_23bca_959f9c8,R_23bcc_9d29a20,R_23bd0_95a0e20,
        R_23bd2_9d29b70,R_23bd4_962fb58,R_23bd6_95a0f70,R_23bd8_9d29c18,R_23bda_9619ae0,R_23bdc_9619b88,R_23bde_9619d80,R_23be0_9619e28,R_23be2_961a020,R_23be6_961a0c8,
        R_23be8_961a218,R_23bea_961a4b8,R_23bec_961a800,R_23bee_961a8a8,R_23bf0_961a950,R_23bf2_961ad40,R_23bf4_961ade8,R_23bf6_961ae90,R_23bf8_961af38,R_23bfc_9d26060,
        R_23bfe_961b088,R_23c00_9d29d68,R_23c02_961b1d8,R_239cc_95f4af8,R_239ce_962fd50,R_239d0_9558e00,R_239d2_9d261b0,R_239d4_95f52d8,R_239d6_9558ea8,R_239d8_961b670,
        R_239da_95f5620,R_239dc_961b910,R_239de_9d2b850,R_239e0_9d2b9a0,R_239e2_9d29e10,R_239e4_9d2a158,R_239e6_961bb08,R_239e8_961c978,R_239ea_961cd68,R_239ec_9d2baf0,
        R_239ee_95f5968,R_239f0_95f5ab8,R_239f2_9d2a2a8,R_239f4_961ce10,R_239f6_9634e08,R_239f8_9d2bb98,R_239fa_9d2bd90,R_239fc_962fdf8,R_239fe_962fea0,R_23a00_961d200,
        R_23a02_961d5f0,R_23a04_961d698,R_23a06_962fff0,R_23a08_961d740,R_23a0a_961d938,R_23c24_9d2a698,R_23c26_9d2c420,R_23c28_962ac98,R_23c2a_9d2c4c8,R_23c2c_9d2c570,
        R_23c2e_95f63e8,R_23c30_9d2a890,R_23c32_962ad40,R_23c22_9d2aa88,R_23c34_9d2c810,R_23c36_9d2ab30,R_23c38_9d2c8b8,R_23c3a_9d2cab0,R_23c20_9635e70,R_23c52_962b868,
        R_23c54_9d2af20,R_23c56_9d2b310,R_23774_9630098,R_2378a_962b9b8,R_237a0_9d2cd50,R_237b6_962bb08,R_237cc_9d2cff0,R_237e2_9d2d098,R_237ec_9d2d140,R_237ee_9d2d290,
        R_237f0_962c240,R_237f2_9559688,R_23776_96301e8,R_23778_9d2d7d0,R_2377a_962c2e8,R_2377c_9d2d878,R_2377e_962ce10,R_23780_9d2d920,R_23782_962d938,R_23784_962e5b0,
        R_23786_9d2d9c8,R_23788_9d2dc68,R_2378c_9d2dd10,R_2378e_9d2ddb8,R_23790_9d2e100,R_23792_9d2e1a8,R_23794_9d2f0c0,R_23796_9630290,R_23798_96303e0,R_2379a_9d2f210,
        R_2379c_9d2f7f8,R_2379e_9630728,R_237a2_96307d0,R_237a4_9d2fb40,R_237a6_9d301d0,R_237a8_9559bc8,R_237aa_9630140,R_237ac_96312f8,R_237ae_9d30710,R_237b0_9630b18,
        R_237b2_9630c68,R_237b4_9d309b0,R_237b8_9630d10,R_237ba_9630fb0,R_237bc_9631100,R_237be_9d30a58,R_237c0_9d30da0,R_237c2_96311a8,R_237c4_96313a0,R_237c6_96318e0,
        R_237c8_9631a30,R_237ca_9d30e48,R_237ce_9d31190,R_237d0_9631b80,R_237d2_9d31f58,R_237d4_9631448,R_237d6_9631790,R_237d8_9d323f0,R_237da_9631ad8,R_237dc_9d32540,
        R_237de_9632018,R_237e0_9631cd0,R_237e4_9632210,R_237e6_9d32690,R_237e8_96322b8,R_237ea_9d32888,R_237f4_9631e20,R_2380a_9d329d8,R_23820_9d32a80,R_23836_9d32f18,
        R_2384c_9d2b3b8,R_23862_9631ec8,R_2386c_9632360,R_2386e_9632a98,R_23870_9d32fc0,R_23872_9632408,R_237f6_9632600,R_237f8_9d33500,R_237fa_96326a8,R_237fc_9d33650,
        R_237fe_9d336f8,R_23800_9d33a40,R_23802_9632750,R_23804_96328a0,R_23806_9d340d0,R_23808_9632948,R_2380c_9d2b658,R_2380e_9d34418,R_23810_9d34760,R_23812_9d34fe8,
        R_23814_9632de0,R_23816_9632e88,R_23818_9d35720,R_2381a_9d2bc40,R_2381c_b805670,R_2381e_b805868,R_23822_9633080,R_23824_b8060f0,R_23826_9633128,R_23828_9633b00,
        R_2382a_9632b40,R_2382c_9634190,R_2382e_9638720,R_23830_9d2c180,R_23832_96389c0,R_23834_9638a68,R_23838_9d15880,R_2383a_b806198,R_2383c_9d2c768,R_2383e_9d16a38,
        R_23840_9d2ca08,R_23842_b806240,R_23844_9d17170,R_23846_9d17c98,R_23848_b8062e8,R_2384a_b806390,R_2384e_9d2cca8,R_23850_9d17fe0,R_23852_9d18328,R_23854_9d2d1e8,
        R_23856_9d1fd38,R_23858_b8064e0,R_2385a_9d2d3e0,R_2385c_9d220a8,R_2385e_9535d90,R_23860_b806588,R_23864_9d25720,R_23866_b8066d8,R_23868_b806780,R_2386a_9d2d530,
        R_23874_95f7840,R_2388a_95f7e28,R_238a0_9d28e50,R_238b6_95f8170,R_238cc_95fcd90,R_238e2_95fda08,R_238ec_95fdb58,R_238ee_95fdca8,R_238f0_95fdd50,R_238f2_9d2d728,
        R_23876_95ff6e8,R_23878_9535e38,R_2387a_9633668,R_2387c_9f4ddd0,R_2387e_9f51b80,R_23880_9f51e20,R_23882_9d29ac8,R_23884_9f53278,R_23886_9f53320,R_23888_9f54580,
        R_2388c_9f54778,R_2388e_9d2dbc0,R_23890_9d2e250,R_23892_9f548c8,R_23894_9f54970,R_23896_9f54c10,R_23898_9f55348,R_2389a_9f55498,R_2389c_9d2a740,R_2389e_9d2e3a0,
        R_238a2_9d2b070,R_238a4_9633710,R_238a6_9f55b28,R_238a8_9f56260,R_238aa_9f56500,R_238ac_9f5baf8,R_238ae_9ee9d78,R_238b0_9d2ba48,R_238b2_9d2bce8,R_238b4_9eea0c0,
        R_238b8_9eeb518,R_238ba_9eedf18,R_238bc_9eee6f8,R_238be_9ef2010,R_238c0_9537530,R_238c2_9ef2208,R_238c4_9ef3660,R_238c6_9ef3858,R_238c8_9633860,R_238ca_9ef3a50,
        R_238ce_9ef3af8,R_238d0_9ef3ba0,R_238d2_9ef3c48,R_238d4_9ef4620,R_238d6_9d2c2d0,R_238d8_9ef4770,R_238da_9d2cb58,R_238dc_9ef4ab8,R_238de_9ef4c08,R_238e0_9ef4ff8,
        R_238e4_9ef5148,R_238e6_9ef51f0,R_238e8_9d2cf48,R_238ea_9ef53e8,R_238f4_9d2e4f0,R_2390a_96339b0,R_23920_9633c50,R_23936_9d266f0,R_2394c_9d2e838,R_23962_9d2ecd0,
        R_2396c_9d2ed78,R_2396e_9d2f018,R_23970_9d2f168,R_23972_b8068d0,R_238f6_9d2f2b8,R_238f8_9d2f9f0,R_238fa_9d2fde0,R_238fc_9633f98,R_238fe_b806a20,R_23900_96340e8,
        R_23902_9d30320,R_23904_9634580,R_23906_9d305c0,R_23908_9634b68,R_2390c_9d30ba8,R_2390e_9d30c50,R_23910_b806ac8,R_23912_9d32000,R_23914_b806b70,R_23916_9d320a8,
        R_23918_9634c10,R_2391a_9d32150,R_2391c_9634cb8,R_2391e_9d32498,R_23922_9d32738,R_23924_9d327e0,R_23926_9d32b28,R_23928_9d32bd0,R_2392a_9635348,R_2392c_9635690,
        R_2392e_9d32c78,R_23930_9d32d20,R_23932_9635a80,R_23934_9d32dc8,R_23938_9d331b8,R_2393a_9d2d488,R_2393c_9d333b0,R_2393e_9d335a8,R_23940_9d337a0,R_23942_9635b28,
        R_23944_9d2d5d8,R_23946_9d338f0,R_23948_9635bd0,R_2394a_9d33998,R_2394e_9d33ae8,R_23950_9d33b90,R_23952_9636110,R_23954_9d33ce0,R_23956_b806c18,R_23958_9d33ed8,
        R_2395a_9d33f80,R_2395c_9636308,R_2395e_b806cc0,R_23960_9d34028,R_23964_9d34178,R_23966_9d2db18,R_23968_96365a8,R_2396a_9636848,R_23734_96368f0,R_23736_9636998,
        R_23738_9636a40,R_2373a_b7dc0c0,R_2373c_9636b90,R_2373e_9636c38,R_23740_b7dc168,R_23742_b806d68,R_23744_b806e10,R_23746_9636ed8,R_23748_b806eb8,R_2374a_9637028,
        R_2374c_b806f60,R_2374e_b8070b0,R_23750_9d33308,R_23752_b807158,R_23754_9ef5880,R_23756_9d26798,R_23758_9d342c8,R_2375a_9ef5928,R_2375c_96c2b20,R_2375e_9d31820,
        R_23760_9d31970,R_23762_9637178,R_23764_9d26840,R_23766_96372c8,R_23768_9d268e8,R_2376a_9d26a38,R_2376c_9d26ae0,R_2376e_9637370,R_23770_9d26b88,R_23772_9637418,
        R_2398c_96c2fb8,R_2398e_9559c70,R_23990_96c35a0,R_23992_96e8010,R_23994_955a300,R_23996_955a450,R_23998_9d34ca0,R_2399a_96c3840,R_2398a_9d34d48,R_2399c_96c3a38,
        R_2399e_96c3d80,R_239a0_955a840,R_239a2_96c59b8,R_23988_96eaf50,R_239ba_96ca728,R_239bc_955b8a8,R_239be_b7db6e8,R_234dc_b8085b0,R_234f2_b80b988,R_23508_b808658,
        R_2351e_b808700,R_23534_b8087a8,R_2354a_b8088f8,R_23554_b80ba30,R_23556_b80bb80,R_23558_b80bec8,R_2355a_b80bf70,R_234de_b8089a0,R_234e0_b808a48,R_234e2_b809768,
        R_234e4_b809df8,R_234e6_b80c2b8,R_234e8_b80e040,R_234ea_b80e580,R_234ec_b80c600,R_234ee_b80f0a8,R_234f0_b80fd20,R_234f4_b80c750,R_234f6_b80ffc0,R_234f8_b7ddf98,
        R_234fa_b80c7f8,R_234fc_b7de0e8,R_234fe_b7de388,R_23500_b7de430,R_23502_b80c9f0,R_23504_b7de580,R_23506_b80ca98,R_2350a_b7de820,R_2350c_b7dea18,R_2350e_b7dee08,
        R_23510_b80cc90,R_23512_b80cd38,R_23514_b7df1f8,R_23516_b80ce88,R_23518_b7df348,R_2351a_b7df540,R_2351c_b80cf30,R_23520_b7dfc78,R_23522_b80d080,R_23524_b80d278,
        R_23526_b7dff18,R_23528_b80d320,R_2352a_b7e0068,R_2352c_b80d5c0,R_2352e_b7e01b8,R_23530_b80d668,R_23532_b7e0458,R_23536_b7e05a8,R_23538_b80d7b8,R_2353a_b80de48,
        R_2353c_b7e0998,R_2353e_b7e0b90,R_23540_b7e1178,R_23542_b80e430,R_23544_b80e628,R_23546_b80e778,R_23548_b7e1568,R_2354c_b80e970,R_2354e_b7e16b8,R_23550_b80eb68,
        R_23552_b7e1808,R_2355c_b7e18b0,R_23572_b805c58,R_23588_b7e1958,R_2359e_b80ed60,R_235b4_95ad7d8,R_235ca_b806438,R_235d4_b7e1a00,R_235d6_b80f000,R_235d8_b7e1bf8,
        R_235da_b7e1ca0,R_2355e_b7e1e98,R_23560_95ad9d0,R_23562_b7e1f40,R_23564_95adb20,R_23566_b7e1fe8,R_23568_b80f3f0,R_2356a_b80f5e8,R_2356c_b806630,R_2356e_b7e2090,
        R_23570_b80f690,R_23574_b7e2138,R_23576_b7e21e0,R_23578_b7e23d8,R_2357a_b7e2720,R_2357c_b7e2870,R_2357e_b7e29c0,R_23580_b806828,R_23582_b7e2a68,R_23584_b7e2c60,
        R_23586_b7e2f00,R_2358a_b80f7e0,R_2358c_96cb8e0,R_2358e_b7e2fa8,R_23590_b7e30f8,R_23592_b806978,R_23594_b807008,R_23596_b7e32f0,R_23598_b80fb28,R_2359a_b7e3398,
        R_2359c_b807698,R_235a0_b7e34e8,R_235a2_96cbb80,R_235a4_b80fbd0,R_235a6_96cc018,R_235a8_95adf10,R_235aa_b7e36e0,R_235ac_b807890,R_235ae_b7e3788,R_235b0_b7e38d8,
        R_235b2_b7e3ad0,R_235b6_b7e3cc8,R_235b8_b7e3f68,R_235ba_b807f20,R_235bc_b807fc8,R_235be_b8101b8,R_235c0_b7e40b8,R_235c2_b7e4208,R_235c4_b8105a8,R_235c6_b810650,
        R_235c8_96cc210,R_235cc_b7e42b0,R_235ce_b7e4400,R_235d0_b7e4550,R_235d2_b7e45f8,R_235dc_b8106f8,R_235f2_b7e46a0,R_23608_b808118,R_2361e_b7e47f0,R_23634_b7e49e8,
        R_2364a_b7dd860,R_23654_95ae060,R_23656_b7dd908,R_23658_b7ddda0,R_2365a_b7dde48,R_235de_9637b50,R_235e0_95ae1b0,R_235e2_b7ddef0,R_235e4_b7de238,R_235e6_b7e4b38,
        R_235e8_9637fe8,R_235ea_b7de2e0,R_235ec_b808310,R_235ee_9638138,R_235f0_96381e0,R_235f4_b7e4d30,R_235f6_96383d8,R_235f8_b7de6d0,R_235fa_9638480,R_235fc_b7de8c8,
        R_235fe_9638528,R_23600_96385d0,R_23602_b7de970,R_23604_b7deac0,R_23606_9638678,R_2360a_96387c8);
input RIde68638_3981,RIde67cd8_3982,RIde68f20_3980,RIb79b518_270,RIdbb8138_3227,RIe548ff0_6844,RIe549ef0_6842,RIe5319e0_6884,RIe549770_6843,
        RIe4f85f0_6398,RIdaea590_2835,RIe4301f0_6000,RIde3d1e0_4027,RIe00b330_4420,RIe160838_5254,RIe0d49f0_4816,RIda11c00_2446,RIe269120_5609,RId958f08_2058,
        RId888d80_1669,RIdc6ed48_3642,RIe5c2e08_6791,RId6f3a80_883,RId7bf4e0_1272,RIb7b93b0_251,RIdba4548_3251,RIe4fa198_6396,RIdaebc88_2833,RIe431ac8_5998,
        RIde3ed88_4025,RIe00ce60_4418,RIe1615d0_5253,RIe0d62c8_4814,RIda13640_2444,RIe26a7a0_5607,RId95a600_2056,RId88a478_1667,RIdc70800_3640,RIe5c4500_6789,
        RId6f5100_881,RId7c0e30_1270,RIb7b94a0_249,RIdbb7328_3228,RIe4f7a38_6399,RIdae97f8_2836,RIe42f4d0_6001,RIde3c448_4028,RIe00a598_4421,RIe172718_5244,
        RIe0d3dc0_4817,RIda10df0_2447,RIe268568_5610,RId9582d8_2059,RId888240_1670,RIdc6e280_3643,RIe5c22c8_6792,RId7064a0_859,RId7be838_1273,RIb7af720_252,
        RIdbb6518_3229,RIe4f6ef8_6400,RIdae8a60_2837,RIe42e8a0_6002,RIde3b728_4029,RIe009710_4422,RIe163e20_5250,RIe0d2e48_4818,RIda101c0_2448,RIe2679b0_5611,
        RId957720_2060,RId89b638_1645,RIdc6d740_3644,RIe5c1710_6793,RId705780_860,RId7d2338_1248,RIb7af6a8_253,RIe4faf30_6395,RIdba51f0_3250,RIe4326f8_5997,
        RIdad5d70_2860,RIde3fb20_4024,RIe00db80_4417,RIe164b40_5249,RIe0d6fe8_4813,RIda143d8_2443,RIe26b2e0_5606,RId95b1b8_2055,RId88b030_1666,RIdc71610_3639,
        RIe5c4fc8_6788,RId6f5cb8_880,RId7c1b50_1269,RIb7b9518_248,RIdba3828_3252,RIe4f9388_6397,RIdaeb0d0_2834,RIe430e20_5999,RIde3df00_4026,RIe00c0c8_4419,
        RIe163088_5251,RIe0d55a8_4815,RIda12920_2445,RIe269c60_5608,RId959a48_2057,RId889938_1668,RIdc6f9f0_3641,RIe5c3948_6790,RId6f4638_882,RId7c0110_1271,
        RIb7b9428_250,RIdba6bb8_3248,RIe4fc9e8_6393,RIdad7918_2858,RIe4340c0_5995,RIde415d8_4022,RIe00f6b0_4415,RIe162368_5252,RIe0d89b0_4811,RIda15da0_2441,
        RIe26ce10_5604,RId95c8b0_2053,RId88c728_1664,RIdd731d8_3637,RId7c3590_1267,RIe5c6738_6786,RId6f73b0_878,RIb7b9608_246,RIdba5e98_3249,RIe4fbcc8_6394,
        RIdad6b80_2859,RIe4333a0_5996,RIde408b8_4023,RIe00e918_4416,RIe1658d8_5248,RIe0d7d08_4812,RIda150f8_2442,RIe26c000_5605,RId95bcf8_2054,RId88bbe8_1665,
        RIdc72420_3638,RIe5c5bf8_6787,RId6f68e8_879,RId7c2870_1268,RIb7b9590_247,RIe5349b0_6879,RIe5341b8_6880,RIe5339c0_6881,RIe5331c8_6882,RIe5329d0_6883,
        RIeb72150_6905,RIe5359a0_6877,RIe5351a8_6878,RIeab7d00_6896,RIeab78c8_6895,RIeab6518_6891,RIeacfa18_6902,RIeab80c0_6897,RIeb352c8_6904,RIea94af8_6890,
        RIeab87c8_6898,RIe15c260_5259,RIe0f3878_4787,RIde5d760_3998,RIdfce700_4467,RIe3f7760_6049,RIe3887c0_5578,RIe5e3568_6762,RIe51acb8_6366,RId7e6f90_1232,
        RId71e398_838,RId8ac078_1630,RId97ab20_2022,RIdb01d80_2813,RIda2def0_2418,RIdbcc7f0_3208,RIdd963e0_3603,RIb7af3d8_259,RIe182a68_5243,RIe0f3008_4788,
        RIde5ad30_4003,RIdfc11b8_4469,RIe3f8a98_6047,RIe385d90_5583,RIe5e09d0_6767,RIe4af828_6445,RId7e5f28_1234,RId71bad0_843,RId8ab538_1631,RId977f88_2027,
        RIdaff2d8_2817,RIda2b970_2422,RIdbcac48_3211,RIdd93500_3608,RIb7af630_254,RIdaffda0_2816,RIda2c258_2421,RIdb62338_3285,RIdd93ed8_3607,RIde5b618_4002,
        RIdfc07e0_4470,RIe1bcc68_5184,RIe088e38_4865,RId978960_2026,RId8ae508_1629,RId71c2c8_842,RId7827c0_1310,RIe386678_5582,RIe450d88_5972,RIe519818_6368,
        RIe5e1330_6766,RIb7af5b8_255,RIdabee68_2890,RIda2cbb8_2420,RIdb8a760_3284,RIdd95288_3605,RIde5c6f8_4000,RIe02a8c0_4391,RIe1bdd48_5182,RIe0aeb60_4864,
        RId9799c8_2024,RId8aed00_1628,RId71d330_840,RId790848_1309,RIe3876e0_5580,RIe3e5628_6050,RIe51a2e0_6367,RIe5e2488_6764,RIb7af4c8_257,RIe1be5b8_5181,
        RIe0b0870_4861,RIde5dfd0_3997,RIdfcf2b8_4466,RIe451670_5971,RIe388fb8_5577,RIe588848_6840,RIe4bd310_6442,RId7a4bb8_1307,RId71ec08_837,RId86c4d8_1705,
        RId97b318_2021,RIdb02668_2812,RIda2e760_2417,RIdbcd0d8_3207,RIdd96cc8_3602,RIb7a5bf8_260,RIe15b900_5260,RIe0f4070_4786,RIde5e840_3996,RIdfcfc90_4465,
        RIe3f9470_6046,RIe3898a0_5576,RIe5e3e50_6761,RIe4b0a70_6443,RId7e7800_1231,RId71f400_836,RId8b0290_1626,RId97bc00_2020,RIdb02f50_2811,RIda2f0c0_2416,
        RIdbcd9c0_3206,RIdd97538_3601,RIb7a0c48_261,RIe3f9e48_6045,RIe387ed8_5579,RIe5e2d70_6763,RIe4bdce8_6441,RIde5cf68_3999,RIdfcdc38_4468,RIe183440_5242,
        RIe0aff10_4862,RId97a238_2023,RId8af7c8_1627,RId71dba0_839,RId7a41e0_1308,RIda2d4a0_2419,RIdb01498_2814,RIdbcbe18_3209,RIdd95b70_3604,RIb7af450_258,
        RIde5be10_4001,RIe02a050_4392,RIe1bd4d8_5183,RIe0af538_4863,RIe3f8048_6048,RIe386e70_5581,RIe5e1ba0_6765,RIe4b0200_6444,RId9791d0_2025,RId86cf28_1704,
        RId71cb38_841,RId7e6798_1233,RId9cdfc8_2495,RIdb00bb0_2815,RIdbcb530_3210,RIdd94928_3606,RIb7af540_256,RIea91330_6888,RIb7b9680_245,RIde4ec88_4006,
        RIb79b4a0_271,RIb79b338_274,RIde612e8_3992,RIde5fec0_3994,RIde60988_3993,RIde69970_3979,RIde6a2d0_3978,RIde6ad98_3977,RIde63250_3989,RIde62878_3990,
        RIde61e28_3991,RIb839848_152,RIe545dc8_6851,RIe545648_6852,RIea90778_6887,RIe546890_6849,RIe546098_6850,RIb8396e0_155,RIb839668_156,RIb79b3b0_273,
        RIde5f3f8_3995,RIde4c8e8_4009,RIb7b96f8_244,RIde4d6f8_4008,RIb7c20c8_243,RIde431f8_4020,RIb7c5728_242,RIde43f90_4019,RIb7c57a0_241,RIde44da0_4018,
        RIb7c5818_240,RIde45ac0_4017,RIb7c5890_239,RIde468d0_4016,RIb7c5908_238,RIde4fb10_4005,RIb7a09f0_266,RIde49300_4013,RIb7a0a68_265,RIde4a020_4012,
        RIb7a0ae0_264,RIde4ae30_4011,RIb7a0b58_263,RIde4bb50_4010,RIb7a0bd0_262,RIdbee210_3713,RIb839b90_145,RIe667bb0_6885,RIe667f70_6886,RIea91768_6889,
        RIeab7058_6894,RIb87eb00_69,RIb7c5980_237,RIdbecc08_3714,RIb87eb78_68,RIb7c59f8_236,RIdbebab0_3715,RIb87ebf0_67,RIb7c5a70_235,RIdbea4a8_3716,
        RIb882ca0_66,RIb7cade0_234,RIdbe9350_3717,RIb885310_65,RIb7cae58_233,RIdbe7d48_3718,RIb885388_64,RIb7caed0_232,RIdbe6bf0_3719,RIb885400_63,
        RIb7caf48_231,RIdbe5a98_3720,RIb885478_62,RIb7cafc0_230,RIdbe4490_3721,RIb8854f0_61,RIb7cb038_229,RIdbe3338_3722,RIb885568_60,RIb7cb0b0_228,
        RIdbe1d30_3723,RIb8855e0_59,RIb7cb128_227,RIdbe0bd8_3724,RIb885658_58,RIb7d00d8_226,RIdaab098_3725,RIb8856d0_57,RIb8263d8_225,RIdaaf0d0_3726,
        RIb885748_56,RIb826e28_224,RIdab2fa0_3727,RIb8857c0_55,RIb826ea0_223,RIdab8e50_3728,RIb885838_54,RIb826f18_222,RIdabcf00_3729,RIb8858b0_53,
        RIb826f90_221,RIdac3788_3730,RIb885928_52,RIb8293a8_220,RIdac8eb8_3731,RIb8859a0_51,RIb829420_219,RIdacf650_3732,RIb885a18_50,RIb829498_218,
        RIdad4fd8_3733,RIb885a90_49,RIb829510_217,RIdadaf00_3734,RIb885b08_48,RIb829588_216,RIdae2610_3735,RIb885b80_47,RIb829600_215,RIdae8268_3736,
        RIb885bf8_46,RIb829678_214,RIdaef720_3737,RIb885c70_45,RIb8296f0_213,RIdaf4e50_3738,RIb885ce8_44,RIb82dae8_212,RIdafa508_3739,RIb885d60_43,
        RIb82db60_211,RIdafe630_3740,RIb885dd8_42,RIb82dbd8_210,RIdb03b08_3741,RIb885e50_41,RIb82dc50_209,RIdb09d00_3742,RIb885ec8_40,RIb82dcc8_208,
        RIdb0e440_3743,RIb885f40_39,RIb82dd40_207,RIdb13468_3744,RIb885fb8_38,RIb82ddb8_206,RId9d7370_3745,RIb886030_37,RIb82de30_205,RId9d25a0_3746,
        RIb8860a8_36,RIb832228_204,RId9cd0c8_3747,RIb886120_35,RIb8322a0_203,RId9c86b8_3748,RIb886198_34,RIb832318_202,RIda940a0_3749,RIb886210_33,
        RIb832390_201,RIda91850_3750,RIb886288_32,RIb832408_200,RIda8dbd8_3751,RIb886300_31,RIb832480_199,RIda8a7d0_3752,RIb886378_30,RIb8324f8_198,
        RIda86978_3753,RIb8863f0_29,RIb832570_197,RIda835e8_3754,RIb886468_28,RIb8383a8_196,RIda80f00_3755,RIb8864e0_27,RIb838420_195,RIda7daf8_3756,
        RIb886558_26,RIb838498_194,RIda7a7e0_3757,RIb8865d0_25,RIb838510_193,RIda745e8_3758,RIb886648_24,RIb838588_192,RIda6e018_3759,RIb8866c0_23,
        RIb838600_191,RIda65e40_3760,RIb886738_22,RIb838678_190,RIda5f888_3761,RIb8867b0_21,RIb8386f0_189,RIda59780_3762,RIb886828_20,RIb838768_188,
        RIda510f8_3763,RIb8868a0_19,RIb8387e0_187,RIda4aff0_3764,RIb886918_18,RIb838858_186,RId927408_3765,RIb886990_17,RIb8388d0_185,RId943680_3766,
        RIb886a08_16,RIb838948_184,RId96ccd8_3767,RIb886a80_15,RIb8389c0_183,RId988b30_3768,RIb886af8_14,RIb838a38_182,RId90bb68_3769,RIb886b70_13,
        RIb838ab0_181,RId8f7438_3770,RIb886be8_12,RIb838b28_180,RId8d6dc8_3771,RIb886c60_11,RIb838ba0_179,RId6c4d70_3772,RIb886cd8_10,RIb838c18_178,
        RId6ae7c8_3773,RIb886d50_9,RIb838c90_177,RId835578_3774,RIb886dc8_8,RIb838d08_176,RId8a9d50_3775,RIb886e40_7,RIb838d80_175,RId862aa0_3776,
        RIb886eb8_6,RIb838df8_174,RId99e778_3777,RId9ac620_3778,RId9b8290_3779,RId9bdfd8_3780,RId90fe70_3781,RId918b10_3782,RIda42698_3783,RIda33a58_3784,
        RIda28b08_3785,RIda18aa0_3786,RIda0b288_3787,RId9f8d18_3788,RId9ec9a0_3789,RId9e3418_3790,RIdb156a0_3791,RIdb17f68_3792,RIdb1b640_3793,RIdb1df08_3794,
        RIdb215e0_3795,RIdb23ea8_3796,RIdb26c20_3797,RIdb29e48_3798,RIdb2cbc0_3799,RIdb2fde8_3800,RIdb32b60_3801,RIdb35d88_3802,RIdb38b00_3803,RIdb3b3c8_3804,
        RIdb3eaa0_3805,RIdb404e0_3806,RIdb422e0_3807,RIdb43ac8_3808,RIdb45850_3809,RIdb47128_3810,RIdb483e8_3811,RIdb49888_3812,RIdb4abc0_3813,RIdb4c330_3814,
        RIdb4d410_3815,RIdb4e5e0_3816,RIdb4fa08_3817,RIdb51100_3818,RIdb52c30_3819,RIdb541c0_3820,RIdb559a8_3821,RIdb56e48_3822,RIdb58900_3823,RIdb5a070_3824,
        RIdb5b588_3825,RIdb5d0b8_3826,RIdb5e3f0_3827,RIda95720_3828,RIda97598_3829,RIda99a28_3830,RIda9bd50_3831,RIda9df10_3832,RIda9f4a0_3833,RIdaa1228_3834,
        RIdaa2d58_3835,RIdaa4a68_3836,RIdaa6b38_3837,RIdaa89b0_3838,RIdbdf030_3839,RIdbdcd80_3840,RIdbdaff8_3841,RIdbd9540_3842,RIdbd6e58_3843,RIdbd4860_3844,
        RIdbd25b0_3845,RIdbd0030_3846,RIdbcdc18_3847,RIdbcb800_3848,RIdbc9730_3849,RIdbc7a20_3850,RIdbc5e78_3851,RIdbc40f0_3852,RIdbc1f30_3853,RIdbbf938_3854,
        RIdbbd4a8_3855,RIdbba910_3856,RIdbb8480_3857,RIdbb58e8_3858,RIdbb2648_3859,RIdbb0758_3860,RIdbad788_3861,RIdbaad58_3862,RIdba7d88_3863,RIdba55b0_3864,
        RIdba2ce8_3865,RIdb9fe80_3866,RIdb9d4c8_3867,RIdb9acf0_3868,RIdb98c20_3869,RIdb96178_3870,RIdb93ce8_3871,RIdb916f0_3872,RIdb8e2e8_3873,RIdb8b840_3874,
        RIdb890e0_3875,RIdb86cc8_3876,RIdb84ec8_3877,RIdb83410_3878,RIdb81700_3879,RIdb7fa68_3880,RIdb7db78_3881,RIdb7bb98_3882,RIdb79e10_3883,RIdb78268_3884,
        RIdb76828_3885,RIdb746e0_3886,RIdda9490_3887,RIdda9c88_3888,RIddaa480_3889,RIddaac78_3890,RIddab470_3891,RIddabc68_3892,RIddac460_3893,RIddacc58_3894,
        RIddad450_3895,RIddadc48_3896,RIddae440_3897,RIddaec38_3898,RIddaf430_3899,RIddafc28_3900,RIddb0420_3901,RIddb0c18_3902,RIddb1410_3903,RIddb1c08_3904,
        RIddb2400_3905,RIddb2bf8_3906,RIddb33f0_3907,RIddb3be8_3908,RIddb43e0_3909,RIddb4bd8_3910,RIddb53d0_3911,RIddb5bc8_3912,RIddb63c0_3913,RIddb6bb8_3914,
        RIddb73b0_3915,RIddb7ba8_3916,RIddb83a0_3917,RIddb8b98_3918,RIddb9390_3919,RIddb9b88_3920,RIddba380_3921,RIddbab78_3922,RIddbb370_3923,RIddbbb68_3924,
        RIddbc360_3925,RIddbcb58_3926,RIddbd350_3927,RIddbdb48_3928,RIddbe340_3929,RIddbeb38_3930,RIddbf330_3931,RIddbfb28_3932,RIddc0320_3933,RIddc0b18_3934,
        RIddc1310_3935,RIddc1b08_3936,RIddc2300_3937,RIddc2af8_3938,RIddc32f0_3939,RIddc3ae8_3940,RIddc42e0_3941,RIddc4ad8_3942,RIddc52d0_3943,RIddc5ac8_3944,
        RIddc62c0_3945,RIddc6ab8_3946,RIddc72b0_3947,RIddc7aa8_3948,RIddc82a0_3949,RIddc8a98_3950,RIddc9290_3951,RIddc9a88_3952,RIddca280_3953,RIddcaa78_3954,
        RIddcb270_3955,RIddcba68_3956,RIddcc260_3957,RIddcca58_3958,RIddcd250_3959,RIddcda48_3960,RIddce240_3961,RIddcea38_3962,RIddcf230_3963,RIddcfa28_3964,
        RIddd0220_3965,RIddd0a18_3966,RIddd1210_3967,RIddd1a08_3968,RIdc0fbb8_3681,RIb86fc68_77,RIdc0f0f0_3682,RIb86fce0_76,RIdc0e5b0_3683,RIb86fd58_75,
        RIdc0dae8_3684,RIb87e8a8_74,RIdc0cfa8_3685,RIb87e920_73,RIdc0c3f0_3686,RIb87e998_72,RIdc0b7c0_3687,RIb87ea10_71,RIdc0ac08_3688,RIb87ea88_70,
        RIdc09f60_3689,RIdc093a8_3690,RIdc08700_3691,RIdc07878_3692,RIdc06270_3693,RIdc05118_3694,RIdc03b10_3695,RIdc029b8_3696,RIdc013b0_3697,RIdc00258_3698,
        RIdbff100_3699,RIdbfdaf8_3700,RIdbfc9a0_3701,RIdbfb398_3702,RIdbfa240_3703,RIdbf8c38_3704,RIdbf7ae0_3705,RIdbf6988_3706,RIdbf5380_3707,RIdbf4228_3708,
        RIdbf2c20_3709,RIdbf1ac8_3710,RIdbf04c0_3711,RIdbef368_3712,RIb79b428_272,RIdda31a8_3581,RIdbd9c48_3186,RIe036f80_4371,RIe100460_4766,RIda3bc30_2396,
        RIde6b9c8_3976,RIdb0e968_2791,RId987e10_2001,RIe527288_6346,RIe45e528_5951,RIe395df8_5556,RIe1ca840_5161,RId72b4a8_816,RIe5efc28_6741,RId8bc950_1606,
        RId7f4028_1211,RId710748_846,RId96d278_2032,RId8aa728_1632,RId7dcb80_1235,RIdbc4870_3212,RIdd8ba30_3609,RIda25c28_2423,RIdaf5f30_2820,RIe022a30_4393,
        RIe0e8ec8_4791,RIe1ac2a0_5191,RIe444fb0_5975,RIe37f9b8_5584,RIe5d6d40_6768,RIe5117a8_6369,RIe3ac2b0_6083,RIe3aaca8_6084,RIe3a9b50_6085,RIe3a8548_6086,
        RIe3a73f0_6087,RIe3a6298_6088,RIe3a4c90_6089,RIe3a3b38_6090,RIe3a2530_6091,RIe3a13d8_6092,RIe39fdd0_6093,RIe39ec78_6094,RIe39db20_6095,RIe39c518_6096,
        RIe1694d8_6097,RIe16e398_6098,RIe173270_6099,RIe178388_6100,RIe17c780_6101,RIe1805d8_6102,RIe1877c0_6103,RIe18c9c8_6104,RIe192ff8_6105,RIe198cc8_6106,
        RIe1a05b8_6107,RIe1a6300_6108,RIe1ac318_6109,RIe1b2420_6110,RIe1b7970_6111,RIe1bce48_6112,RIe1c12b8_6113,RIe1c7960_6114,RIe1cc820_6115,RIe1d0fd8_6116,
        RIe094940_6117,RIe090368_6118,RIe08b700_6119,RIe087a10_6120,RIe14c9f0_6121,RIe1495e8_6122,RIe146348_6123,RIe143210_6124,RIe140a38_6125,RIe13d4c8_6126,
        RIe13a660_6127,RIe137168_6128,RIe133a18_6129,RIe12fda0_6130,RIe1280f0_6131,RIe121b38_6132,RIe1194b0_6133,RIe1133a8_6134,RIe10ad20_6135,RIdfd70d0_6136,
        RIdff52b0_6137,RIe01ea70_6138,RIe03a5e0_6139,RIdfb6cb8_6140,RIdfa46d0_6141,RIdf7c7e8_6142,RIdc22218_6143,RIda953d8_6144,RIddeaf80_6145,RIde58a80_6146,
        RIe03fa40_6147,RIe04e338_6148,RIe0629f0_6149,RIe06c608_6150,RIe0732e0_6151,RIe07d0d8_6152,RIe084158_6153,RIdfc61e0_6154,RIe106838_6155,RIe0f8198_6156,
        RIe0eed00_6157,RIe0e2b68_6158,RIe0d0b98_6159,RIe0c3998_6160,RIe0b0960_6161,RIe0a6988_6162,RIe099440_6163,RIe1d3c60_6164,RIe1d69d8_6165,RIe1d9c00_6166,
        RIe1dc978_6167,RIe1dfba0_6168,RIe1e2918_6169,RIe1e5b40_6170,RIe1e88b8_6171,RIe1eb180_6172,RIe1ee858_6173,RIe1f1120_6174,RIe1f47f8_6175,RIe1f70c0_6176,
        RIe1fa180_6177,RIe1fbad0_6178,RIe1fd330_6179,RIe1ff568_6180,RIe2012f0_6181,RIe203000_6182,RIe203f00_6183,RIe2053a0_6184,RIe2066d8_6185,RIe207920_6186,
        RIe208be0_6187,RIe209d38_6188,RIe20b958_6189,RIe20cf60_6190,RIe20e4f0_6191,RIe20f5d0_6192,RIe211178_6193,RIe212c30_6194,RIe214148_6195,RIe215c00_6196,
        RIe217460_6197,RIe218798_6198,RIe2199e0_6199,RIe14e868_6200,RIe151130_6201,RIe153020_6202,RIe154ad8_6203,RIe156518_6204,RIe158228_6205,RIe15a280_6206,
        RIe15c3c8_6207,RIe15ef60_6208,RIe1616c0_6209,RIe164168_6210,RIe166c10_6211,RIe39a100_6212,RIe3984e0_6213,RIe3967d0_6214,RIe3941d8_6215,RIe391c58_6216,
        RIe38f5e8_6217,RIe38d428_6218,RIe38ae30_6219,RIe389030_6220,RIe386fd8_6221,RIe384ff8_6222,RIe3832e8_6223,RIe381218_6224,RIe37f148_6225,RIe37ce20_6226,
        RIe37aeb8_6227,RIe378668_6228,RIe3755a8_6229,RIe372c68_6230,RIe2703f8_6231,RIe26d4a0_6232,RIe26aae8_6233,RIe2686d0_6234,RIe265ca0_6235,RIe264170_6236,
        RIe2616c8_6237,RIe25f238_6238,RIe25c6a0_6239,RIe259ec8_6240,RIe257240_6241,RIe254018_6242,RIe251408_6243,RIe24e8e8_6244,RIe24c110_6245,RIe248d08_6246,
        RIe246170_6247,RIe2435d8_6248,RIe2418c8_6249,RIe23fb40_6250,RIe23dcc8_6251,RIe23ba18_6252,RIe239948_6253,RIe2381d8_6254,RIe236720_6255,RIe2346c8_6256,
        RIe232a30_6257,RIe230bb8_6258,RIe465cb0_6259,RIe4664a8_6260,RIe466ca0_6261,RIe467498_6262,RIe467c90_6263,RIe468488_6264,RIe468c80_6265,RIe469478_6266,
        RIe469c70_6267,RIe46a468_6268,RIe46ac60_6269,RIe46b458_6270,RIe46bc50_6271,RIe46c448_6272,RIe46cc40_6273,RIe46d438_6274,RIe46dc30_6275,RIe46e428_6276,
        RIe46ec20_6277,RIe46f418_6278,RIe46fc10_6279,RIe470408_6280,RIe470c00_6281,RIe4713f8_6282,RIe471bf0_6283,RIe4723e8_6284,RIe472bf8_6285,RIe4733f0_6286,
        RIe473be8_6287,RIe4743e0_6288,RIe474bd8_6289,RIe4753d0_6290,RIe475bc8_6291,RIe4763c0_6292,RIe476bb8_6293,RIe4773b0_6294,RIe477ba8_6295,RIe4783a0_6296,
        RIe478b98_6297,RIe479390_6298,RIe479b88_6299,RIe47a380_6300,RIe47ab78_6301,RIe47b370_6302,RIe47bb68_6303,RIe47c360_6304,RIe47cb58_6305,RIe47d350_6306,
        RIe47db48_6307,RIe47e340_6308,RIe47eb38_6309,RIe47f330_6310,RIe47fb28_6311,RIe480320_6312,RIe480b18_6313,RIe481310_6314,RIe481b08_6315,RIe482300_6316,
        RIe482af8_6317,RIe4832f0_6318,RIe483ae8_6319,RIe4842e0_6320,RIe484ad8_6321,RIe4852d0_6322,RIe485ac8_6323,RIe4862c0_6324,RIe486ab8_6325,RIe4872b0_6326,
        RIe487aa8_6327,RIe4882a0_6328,RIe488a98_6329,RIe489290_6330,RIe489a88_6331,RIe48a280_6332,RIe48aa78_6333,RIe48b270_6334,RIe48ba68_6335,RIe48c260_6336,
        RIe48ca58_6337,RIe48d250_6338,RIe3cd190_6051,RIe3cc3f8_6052,RIe3cb750_6053,RIe3ca9b8_6054,RIe3c9e00_6055,RIe3c9248_6056,RIe3c8708_6057,RIe3c7bc8_6058,
        RIe3c7100_6059,RIe3c6638_6060,RIe3c5af8_6061,RIe3c4ec8_6062,RIe3c4130_6063,RIe3c31b8_6064,RIe3c1bb0_6065,RIe3c0a58_6066,RIe3bf900_6067,RIe3be2f8_6068,
        RIe3bd1a0_6069,RIe3bbb98_6070,RIe3baa40_6071,RIe3b9438_6072,RIe3b82e0_6073,RIe3b7188_6074,RIe3b5b80_6075,RIe3b4a28_6076,RIe3b3420_6077,RIe3b22c8_6078,
        RIe3b0cc0_6079,RIe3afb68_6080,RIe3aea10_6081,RIe3ad408_6082,RIe51b690_6365,RIe500d68_6388,RIe501998_6387,RIe5026b8_6386,RIe5032e8_6385,RIe503f90_6384,
        RIe504d28_6383,RIe505958_6382,RIe50ef58_6371,RIe50ac50_6376,RIe50b880_6375,RIe50c690_6374,RIe50d428_6373,RIe524060_6351,RIe523688_6352,RIe524948_6350,
        RIe51d5f8_6362,RIe51c158_6364,RIe51cc20_6363,RIe51f290_6359,RIe51dee0_6361,RIe51e840_6360,RIe525410_6349,RIe525d70_6348,RIe5267c0_6347,RIe1e2210_5688,
        RIe1e10b8_5689,RIe1dfab0_5690,RIe1de958_5691,RIe1dd350_5692,RIe1dc1f8_5693,RIe1dabf0_5694,RIe1d9a98_5695,RIe1d8940_5696,RIe1d7338_5697,RIe1d61e0_5698,
        RIe1d4bd8_5699,RIe1d3a80_5700,RIe1d2478_5701,RIe099530_5702,RIe09d298_5703,RIe0a2338_5704,RIe0a6fa0_5705,RIe0ac310_5706,RIe0b16f8_5707,RIe0b9240_5708,
        RIe0bf438_5709,RIe0c4730_5710,RIe0cb0a8_5711,RIe0d0df0_5712,RIe0d8aa0_5713,RIe0de608_5714,RIe0e5ca0_5715,RIe0eb358_5716,RIe0ef138_5717,RIe0f3bc0_5718,
        RIe0f8300_5719,RIe0ff380_5720,RIe103430_5721,RIdfce868_5722,RIdfc9fc0_5723,RIdfc6000_5724,RIdfc1410_5725,RIdfbcc58_5726,RIe082f10_5727,RIe0800a8_5728,
        RIe07bd28_5729,RIe078ec0_5730,RIe075ab8_5731,RIe071f18_5732,RIe06f308_5733,RIe06b0f0_5734,RIe067928_5735,RIe0608a8_5736,RIe05a2f0_5737,RIe0541e8_5738,
        RIe04bb60_5739,RIe045a58_5740,RIe03d3d0_5741,RIde1d908_5742,RIde4a200_5743,RIde62e18_5744,RIdc30d68_5745,RIdde3e10_5746,RIddce948_5747,RIdb96b50_5748,
        RIda0b300_5749,RIdc00960_5750,RIdb708e8_5751,RIdc692d0_5752,RIdf7e930_5753,RIdf8d6d8_5754,RIdf9f978_5755,RIdfa6f20_5756,RIdfaf968_5757,RIdfb74b0_5758,
        RIddf5a98_5759,RIde028d8_5760,RIe036620_5761,RIe027530_5762,RIe01deb8_5763,RIe00b3a8_5764,RIdffd938_5765,RIdfefb08_5766,RIdfe0838_5767,RIdfd6680_5768,
        RIe1084d0_5769,RIe10ad98_5770,RIe10e470_5771,RIe110d38_5772,RIe113ab0_5773,RIe116cd8_5774,RIe119a50_5775,RIe11cc78_5776,RIe11f9f0_5777,RIe122c18_5778,
        RIe125990_5779,RIe128258_5780,RIe12b930_5781,RIe12e1f8_5782,RIe1308e0_5783,RIe132398_5784,RIe134300_5785,RIe135ae8_5786,RIe137258_5787,RIe138608_5788,
        RIe139850_5789,RIe13ab88_5790,RIe13c028_5791,RIe13d5b8_5792,RIe13ead0_5793,RIe13fef8_5794,RIe141230_5795,RIe142568_5796,RIe1434e0_5797,RIe144638_5798,
        RIe145880_5799,RIe146ac8_5800,RIe1486e8_5801,RIe149f48_5802,RIe14b550_5803,RIe14c978_5804,RIe14e430_5805,RIe0865e8_5806,RIe087f38_5807,RIe089db0_5808,
        RIe08b7f0_5809,RIe08d578_5810,RIe08f120_5811,RIe091100_5812,RIe093248_5813,RIe0950c0_5814,RIe096998_5815,RIe0986a8_5816,RIe1cfd18_5817,RIe1ce080_5818,
        RIe1cc550_5819,RIe1ca048_5820,RIe1c78e8_5821,RIe1c4f30_5822,RIe1c26e0_5823,RIe1c0b38_5824,RIe1be9f0_5825,RIe1bcce0_5826,RIe1baf58_5827,RIe1b9158_5828,
        RIe1b6908_5829,RIe1b3b90_5830,RIe1b1d18_5831,RIe1aff90_5832,RIe1ae2f8_5833,RIe1ab940_5834,RIe1a8628_5835,RIe1a6030_5836,RIe1a2d90_5837,RIe1a0540_5838,
        RIe19da20_5839,RIe19a870_5840,RIe197cd8_5841,RIe195410_5842,RIe192e90_5843,RIe190460_5844,RIe18e0c0_5845,RIe18bc30_5846,RIe189098_5847,RIe186c08_5848,
        RIe1839e0_5849,RIe1817a8_5850,RIe17fb88_5851,RIe17def0_5852,RIe17c3c0_5853,RIe17a458_5854,RIe1781a8_5855,RIe176240_5856,RIe174530_5857,RIe172988_5858,
        RIe16fc70_5859,RIe16e140_5860,RIe16c1d8_5861,RIe16a5b8_5862,RIe168a88_5863,RIe167138_5864,RIe39c680_5865,RIe39ce78_5866,RIe39d670_5867,RIe39de68_5868,
        RIe39e660_5869,RIe39ee58_5870,RIe39f650_5871,RIe39fe48_5872,RIe3a0640_5873,RIe3a0e38_5874,RIe3a1630_5875,RIe3a1e28_5876,RIe3a2620_5877,RIe3a2e18_5878,
        RIe3a3610_5879,RIe3a3e08_5880,RIe3a4600_5881,RIe3a4df8_5882,RIe3a55f0_5883,RIe3a5de8_5884,RIe3a65e0_5885,RIe3a6dd8_5886,RIe3a75d0_5887,RIe3a7dc8_5888,
        RIe3a85c0_5889,RIe3a8db8_5890,RIe3a95b0_5891,RIe3a9da8_5892,RIe3aa5a0_5893,RIe3aad98_5894,RIe3ab590_5895,RIe3abd88_5896,RIe3ac580_5897,RIe3acd78_5898,
        RIe3ad570_5899,RIe3add68_5900,RIe3ae560_5901,RIe3aed58_5902,RIe3af550_5903,RIe3afd48_5904,RIe3b0540_5905,RIe3b0d38_5906,RIe3b1530_5907,RIe3b1d28_5908,
        RIe3b2520_5909,RIe3b2d18_5910,RIe3b3510_5911,RIe3b3d08_5912,RIe3b4500_5913,RIe3b4cf8_5914,RIe3b54f0_5915,RIe3b5ce8_5916,RIe3b64e0_5917,RIe3b6cd8_5918,
        RIe3b74d0_5919,RIe3b7cc8_5920,RIe3b84c0_5921,RIe3b8cb8_5922,RIe3b94b0_5923,RIe3b9ca8_5924,RIe3ba4a0_5925,RIe3bac98_5926,RIe3bb490_5927,RIe3bbc88_5928,
        RIe3bc480_5929,RIe3bcc78_5930,RIe3bd470_5931,RIe3bdc68_5932,RIe3be460_5933,RIe3bec58_5934,RIe3bf450_5935,RIe3bfc48_5936,RIe3c0440_5937,RIe3c0c38_5938,
        RIe3c1430_5939,RIe3c1c28_5940,RIe3c2420_5941,RIe3c2c18_5942,RIe3c3410_5943,RIe202f10_5656,RIe202448_5657,RIe201980_5658,RIe200e40_5659,RIe2000a8_5660,
        RIe1ff310_5661,RIe1fe668_5662,RIe1fd9c0_5663,RIe1fce80_5664,RIe1fc340_5665,RIe1fb878_5666,RIe1facc0_5667,RIe1fa090_5668,RIe1f9118_5669,RIe1f7fc0_5670,
        RIe1f69b8_5671,RIe1f5860_5672,RIe1f4258_5673,RIe1f3100_5674,RIe1f1fa8_5675,RIe1f09a0_5676,RIe1ef848_5677,RIe1ee240_5678,RIe1ed0e8_5679,RIe1ebae0_5680,
        RIe1ea988_5681,RIe1e9830_5682,RIe1e8228_5683,RIe1e70d0_5684,RIe1e5ac8_5685,RIe1e4970_5686,RIe1e3368_5687,RIe4520c0_5970,RIe438440_5990,RIe4390e8_5989,
        RIe439f70_5988,RIe43ad80_5987,RIe43ba28_5986,RIe43c7c0_5985,RIe43d5d0_5984,RIe445e38_5974,RIe441c98_5979,RIe4429b8_5978,RIe443750_5977,RIe437630_5991,
        RIe455e28_5964,RIe454988_5966,RIe4554c8_5965,RIe45c278_5954,RIe45cdb8_5953,RIe45d880_5952,RIe45aec8_5956,RIe45a478_5957,RIe45b8a0_5955,RIe4534e8_5968,
        RIe452b88_5969,RIe453fb0_5967,RIe116b70_5293,RIe115a18_5294,RIe114410_5295,RIe1132b8_5296,RIe111cb0_5297,RIe110b58_5298,RIe10f550_5299,RIe10e3f8_5300,
        RIe10d2a0_5301,RIe10bc98_5302,RIe10ab40_5303,RIe109538_5304,RIe1083e0_5305,RIe106dd8_5306,RIdfd3728_5307,RIdfd71c0_5308,RIdfdc8f0_5309,RIdfe0b80_5310,
        RIdfe6760_5311,RIdfeb788_5312,RIdff1f98_5313,RIdff7f38_5314,RIdffe400_5315,RIe005750_5316,RIe00b420_5317,RIe0132b0_5318,RIe0193b8_5319,RIe0202d0_5320,
        RIe023de0_5321,RIe027878_5322,RIe02ccd8_5323,RIe0322a0_5324,RIe038768_5325,RIe03c728_5326,RIde01258_5327,RIddfd748_5328,RIddf9788_5329,RIddf3d88_5330,
        RIdfba228_5331,RIdfb5e30_5332,RIdfb2aa0_5333,RIdfaec48_5334,RIdfabf48_5335,RIdfa97e8_5336,RIdfa5e40_5337,RIdfa2f60_5338,RIdf9e4d8_5339,RIdf99618_5340,
        RIdf90f90_5341,RIdf8ae88_5342,RIdf848d0_5343,RIdf7c248_5344,RIdf76140_5345,RIdc56298_5346,RIdd75f50_5347,RIdd9d6b8_5348,RIdb67180_5349,RIdc198c0_5350,
        RIdc008e8_5351,RIdacdc88_5352,RId8fd180_5353,RIdb353b0_5354,RIdbdbca0_5355,RIdb8b8b8_5356,RIddb1a28_5357,RIddc60e0_5358,RIddd3cb8_5359,RIdddeaa0_5360,
        RIdde50d0_5361,RIddeee50_5362,RIdc2bb60_5363,RIdc34788_5364,RIde6e7b8_5365,RIde62ad0_5366,RIde55510_5367,RIde4a188_5368,RIde36d90_5369,RIde29c80_5370,
        RIde1c210_5371,RIde0cb08_5372,RIe03d4c0_5373,RIe040b98_5374,RIe043460_5375,RIe046b38_5376,RIe049400_5377,RIe04c178_5378,RIe04f3a0_5379,RIe052118_5380,
        RIe055340_5381,RIe0580b8_5382,RIe05b2e0_5383,RIe05e058_5384,RIe060920_5385,RIe063ff8_5386,RIe0662a8_5387,RIe068288_5388,RIe069a70_5389,RIe06b870_5390,
        RIe06cf68_5391,RIe06e6d8_5392,RIe06fa10_5393,RIe070eb0_5394,RIe0721e8_5395,RIe073808_5396,RIe074960_5397,RIe0762b0_5398,RIe0779a8_5399,RIe079118_5400,
        RIe07a798_5401,RIe07bcb0_5402,RIe07d768_5403,RIe07f220_5404,RIe080cd8_5405,RIe082088_5406,RIe083078_5407,RIe0843b0_5408,RIdfbbbf0_5409,RIdfbd5b8_5410,
        RIdfbf3b8_5411,RIdfc15f0_5412,RIdfc30a8_5413,RIdfc4f20_5414,RIdfc6f00_5415,RIdfc85f8_5416,RIdfca3f8_5417,RIdfcc720_5418,RIdfce8e0_5419,RIe106478_5420,
        RIe104948_5421,RIe102b48_5422,RIe100f28_5423,RIe0fea20_5424,RIe0fcd10_5425,RIe0fa3d0_5426,RIe0f7838_5427,RIe0f5a38_5428,RIe0f3968_5429,RIe0f1b68_5430,
        RIe0f0290_5431,RIe0ee508_5432,RIe0ec690_5433,RIe0eaea8_5434,RIe0e8658_5435,RIe0e54a8_5436,RIe0e2988_5437,RIe0e0228_5438,RIe0dd7f8_5439,RIe0da828_5440,
        RIe0d7f60_5441,RIe0d4f18_5442,RIe0d3280_5443,RIe0d02b0_5444,RIe0cdad8_5445,RIe0cae50_5446,RIe0c8150_5447,RIe0c5d38_5448,RIe0c3290_5449,RIe0c0d88_5450,
        RIe0be628_5451,RIe0bbdd8_5452,RIe0b91c8_5453,RIe0b5f28_5454,RIe0b3318_5455,RIe0b02d0_5456,RIe0adeb8_5457,RIe0ac0b8_5458,RIe0aa330_5459,RIe0a83c8_5460,
        RIe0a6a00_5461,RIe0a40c0_5462,RIe0a2158_5463,RIe0a0010_5464,RIe09e378_5465,RIe09c668_5466,RIe09a8e0_5467,RIe099080_5468,RIe1d1cf8_5469,RIe1d24f0_5470,
        RIe1d2ce8_5471,RIe1d34e0_5472,RIe1d3cd8_5473,RIe1d44d0_5474,RIe1d4cc8_5475,RIe1d54c0_5476,RIe1d5cb8_5477,RIe1d64b0_5478,RIe1d6ca8_5479,RIe1d74a0_5480,
        RIe1d7c98_5481,RIe1d8490_5482,RIe1d8c88_5483,RIe1d9480_5484,RIe1d9c78_5485,RIe1da470_5486,RIe1dac68_5487,RIe1db460_5488,RIe1dbc58_5489,RIe1dc450_5490,
        RIe1dcc48_5491,RIe1dd440_5492,RIe1ddc38_5493,RIe1de430_5494,RIe1dec28_5495,RIe1df420_5496,RIe1dfc18_5497,RIe1e0410_5498,RIe1e0c08_5499,RIe1e1400_5500,
        RIe1e1bf8_5501,RIe1e23f0_5502,RIe1e2be8_5503,RIe1e33e0_5504,RIe1e3bd8_5505,RIe1e43d0_5506,RIe1e4bc8_5507,RIe1e53c0_5508,RIe1e5bb8_5509,RIe1e63b0_5510,
        RIe1e6ba8_5511,RIe1e73a0_5512,RIe1e7b98_5513,RIe1e8390_5514,RIe1e8b88_5515,RIe1e9380_5516,RIe1e9b78_5517,RIe1ea370_5518,RIe1eab68_5519,RIe1eb360_5520,
        RIe1ebb58_5521,RIe1ec350_5522,RIe1ecb48_5523,RIe1ed340_5524,RIe1edb38_5525,RIe1ee330_5526,RIe1eeb28_5527,RIe1ef320_5528,RIe1efb18_5529,RIe1f0310_5530,
        RIe1f0b08_5531,RIe1f1300_5532,RIe1f1af8_5533,RIe1f22f0_5534,RIe1f2ae8_5535,RIe1f32e0_5536,RIe1f3ad8_5537,RIe1f42d0_5538,RIe1f4ac8_5539,RIe1f52c0_5540,
        RIe1f5ab8_5541,RIe1f62b0_5542,RIe1f6aa8_5543,RIe1f72a0_5544,RIe1f7a98_5545,RIe1f8290_5546,RIe1f8a88_5547,RIe1f9280_5548,RIe137870_5261,RIe136da8_5262,
        RIe136358_5263,RIe135890_5264,RIe134d50_5265,RIe134288_5266,RIe1337c0_5267,RIe132c08_5268,RIe131fd8_5269,RIe1313a8_5270,RIe1307f0_5271,RIe12fbc0_5272,
        RIe12f080_5273,RIe12da78_5274,RIe12c920_5275,RIe12b318_5276,RIe12a1c0_5277,RIe128bb8_5278,RIe127a60_5279,RIe126908_5280,RIe125300_5281,RIe1241a8_5282,
        RIe122ba0_5283,RIe121a48_5284,RIe120440_5285,RIe11f2e8_5286,RIe11e190_5287,RIe11cb88_5288,RIe11ba30_5289,RIe11a428_5290,RIe1192d0_5291,RIe117cc8_5292,
        RIe38a110_5575,RIe378410_5590,RIe379220_5589,RIe379e50_5588,RIe26f4f8_5601,RIe270290_5600,RIe270ec0_5599,RIe271be0_5598,RIe37b908_5586,RIe375008_5594,
        RIe375da0_5593,RIe376a48_5592,RIe377768_5591,RIe392b58_5561,RIe3921f8_5562,RIe3934b8_5560,RIe38b9e8_5572,RIe38a908_5574,RIe38b1f0_5573,RIe38da40_5569,
        RIe38c4b0_5571,RIe38cf78_5570,RIe393e90_5559,RIe394868_5558,RIe3951c8_5557,RIe04cad8_4898,RIe04b980_4899,RIe04a378_4900,RIe049220_4901,RIe047c18_4902,
        RIe046ac0_4903,RIe045968_4904,RIe044360_4905,RIe043208_4906,RIe041c00_4907,RIe040aa8_4908,RIe03f4a0_4909,RIe03e348_4910,RIe03d1f0_4911,RIde08bc0_4912,
        RIde0d030_4913,RIde131b0_4914,RIde17968_4915,RIde1f528_4916,RIde24e38_4917,RIde29ed8_4918,RIde31390_4919,RIde36e08_4920,RIde3efe0_4921,RIde45070_4922,
        RIde4c9d8_4923,RIde51b68_4924,RIde553a8_4925,RIde59c50_4926,RIde5e390_4927,RIde65668_4928,RIde6a4b0_4929,RIde6f820_4930,RIdf73710_4931,RIdc38040_4932,
        RIdc32b68_4933,RIdc2ee78_4934,RIdc29bf8_4935,RIddf1628_4936,RIddee388_4937,RIddeaa58_4938,RIdde7a88_4939,RIdde35a0_4940,RIdde0cd8_4941,RIddddf60_4942,
        RIdddb710_4943,RIddd5e78_4944,RIddd2278_4945,RIddcc080_4946,RIddc39f8_4947,RIddbd8f0_4948,RIddb5268_4949,RIddaf160_4950,RIdb7c228_4951,RIdb96c40_4952,
        RIdbbbd38_4953,RIdbdcdf8_4954,RIdb5db80_4955,RIdb48190_4956,RIdb26ba8_4957,RId917aa8_4958,RId986da8_4959,RIda7eb60_4960,RIdaf90e0_4961,RIdab27a8_4962,
        RIdbf1ca8_4963,RIdc00a50_4964,RIdc0fe88_4965,RIdc16080_4966,RIdc1c098_4967,RIdc25080_4968,RIdb67810_4969,RIdda8518_4970,RIdd9d5c8_4971,RIdd8f270_4972,
        RIdd82fe8_4973,RIdd74150_4974,RIdc641b8_4975,RIdc54600_4976,RIdc46848_4977,RIdc3b970_4978,RIdf77220_4979,RIdf79f98_4980,RIdf7c860_4981,RIdf7ff38_4982,
        RIdf82800_4983,RIdf85ed8_4984,RIdf887a0_4985,RIdf8be78_4986,RIdf8e740_4987,RIdf91008_4988,RIdf946e0_4989,RIdf96fa8_4990,RIdf9a680_4991,RIdf9ccf0_4992,
        RIdf9ec58_4993,RIdfa04b8_4994,RIdfa1bb0_4995,RIdfa3b18_4996,RIdfa4dd8_4997,RIdfa6110_4998,RIdfa75b0_4999,RIdfa88e8_5000,RIdfa9d10_5001,RIdfab048_5002,
        RIdfac218_5003,RIdfad460_5004,RIdfaecc0_5005,RIdfb0610_5006,RIdfb1c90_5007,RIdfb3310_5008,RIdfb4828_5009,RIdfb5d40_5010,RIdfb77f8_5011,RIdfb92b0_5012,
        RIdfba9a8_5013,RIddf2ca8_5014,RIddf4580_5015,RIddf6308_5016,RIddf8270_5017,RIddf9e90_5018,RIddfbdf8_5019,RIddfdb08_5020,RIddff548_5021,RIde015a0_5022,
        RIde03508_5023,RIde04fc0_5024,RIe03bbe8_5025,RIe039cf8_5026,RIe038600_5027,RIe0363c8_5028,RIe033b78_5029,RIe031580_5030,RIe02ee98_5031,RIe02c4e0_5032,
        RIe02a488_5033,RIe028958_5034,RIe026b58_5035,RIe025460_5036,RIe023b88_5037,RIe021fe0_5038,RIe020168_5039,RIe01dcd8_5040,RIe01b758_5041,RIe018440_5042,
        RIe0157b8_5043,RIe012590_5044,RIe010628_5045,RIe00d298_5046,RIe00a778_5047,RIe007e38_5048,RIe004df0_5049,RIe0024b0_5050,RIdfff558_5051,RIdffcd08_5052,
        RIdffa260_5053,RIdff7b78_5054,RIdff4f68_5055,RIdff1ea8_5056;
output R_25610_96cc360,R_25642_95f0d48,R_25644_9598060,R_25646_95984f8,R_25614_953c348,R_25616_96251f8,R_25618_96ed6b0,R_2561a_95f00d0,R_2561c_95f0418,
        R_2561e_95f0760,R_25620_953c3f0,R_25622_953c690,R_25612_953c9d8,R_25624_95f08b0,R_25626_953ca80,R_25628_96253f0,R_2562a_9632be8,R_253fc_9d20ef0,R_25412_9530108,
        R_25428_95f75a0,R_2543e_95301b0,R_25454_95304f8,R_2546a_9533198,R_25474_95332e8,R_25476_96dee60,R_25478_95f7798,R_2547a_96def08,R_253fe_95f7990,R_25400_9d21190,
        R_25402_9d21388,R_25404_9589e90,R_25406_9d21430,R_25408_9533780,R_2540a_9533b70,R_2540c_9d216d0,R_2540e_958a5c8,R_25410_96defb0,R_25414_9d21778,R_25416_9d21cb8,
        R_25418_95f7ae0,R_2541a_9d21d60,R_2541c_96df100,R_2541e_9d221f8,R_25420_958ac58,R_25422_95f7b88,R_25424_9533c18,R_25426_958b630,R_2542a_9d222a0,R_2542c_9533d68,
        R_2542e_95f7c30,R_25430_9d22498,R_25432_9d22540,R_25434_9533f60,R_25436_96df1a8,R_25438_95f7f78,R_2543a_9534008,R_2543c_9534200,R_25440_95f80c8,R_25442_96df250,
        R_25444_9d22690,R_25446_95fa438,R_25448_95fa4e0,R_2544a_958bcc0,R_2544c_9d22738,R_2544e_9d227e0,R_25450_9d22888,R_25452_9d22930,R_25456_9d229d8,R_25458_95fa588,
        R_2545a_9534350,R_2545c_95fa828,R_2545e_9d22a80,R_25460_96df2f8,R_25462_96df3a0,R_25464_95343f8,R_25466_95fa8d0,R_25468_95faac8,R_2546c_958bd68,R_2546e_958be10,
        R_25470_95fab70,R_25472_9d22b28,R_2547c_958beb8,R_25492_9d22bd0,R_254a8_958bf60,R_254be_9d22c78,R_254d4_9d22dc8,R_254ea_9d22e70,R_254f4_958c0b0,R_254f6_9d22f18,
        R_254f8_958c158,R_254fa_9d22fc0,R_2547e_958c200,R_25480_9d23068,R_25482_9d231b8,R_25484_958c2a8,R_25486_958c350,R_25488_9d23458,R_2548a_958c4a0,R_2548c_9d235a8,
        R_2548e_9d236f8,R_25490_958c548,R_25494_958c5f0,R_25496_9d237a0,R_25498_958c698,R_2549a_958f728,R_2549c_9d23848,R_2549e_958f7d0,R_254a0_958f878,R_254a2_9d23998,
        R_254a4_9d23ae8,R_254a6_9d23c38,R_254aa_9d23d88,R_254ac_9d23e30,R_254ae_9d23f80,R_254b0_9d24028,R_254b2_9d240d0,R_254b4_9d24220,R_254b6_9d242c8,R_254b8_9590988,
        R_254ba_9590a30,R_254bc_9590cd0,R_254c0_9d24418,R_254c2_9590d78,R_254c4_9590f70,R_254c6_9591178,R_254c8_9d24568,R_254ca_9d24bf8,R_254cc_9d25090,R_254ce_95916b8,
        R_254d0_9591808,R_254d2_9d251e0,R_254d6_9d25f10,R_254d8_9d25fb8,R_254da_95918b0,R_254dc_9d265a0,R_254de_9591958,R_254e0_9d26990,R_254e2_9d26c30,R_254e4_9591a00,
        R_254e6_95347e8,R_254e8_9591b50,R_254ec_9591bf8,R_254ee_9d26d80,R_254f0_9d27368,R_254f2_9d27410,R_254fc_96df4f0,R_25512_9d276b0,R_25528_96df598,R_2553e_9534890,
        R_25554_9d27c98,R_2556a_96df640,R_25574_9d27de8,R_25576_96df6e8,R_25578_9534bd8,R_2557a_96df838,R_254fe_96dfad8,R_25500_9534d28,R_25502_9534dd0,R_25504_9534f20,
        R_25506_9d281d8,R_25508_96dfb80,R_2550a_9d28328,R_2550c_9d283d0,R_2550e_96dfc28,R_25510_9534fc8,R_25514_96dfcd0,R_25516_9d28520,R_25518_96dfe20,R_2551a_96dfec8,
        R_2551c_9535070,R_2551e_95351c0,R_25520_9535268,R_25522_96dff70,R_25524_96e0018,R_25526_96e00c0,R_2552a_9535310,R_2552c_96e0168,R_2552e_96e0210,R_25530_96e02b8,
        R_25532_96e0408,R_25534_96e0558,R_25536_96e0600,R_25538_9535658,R_2553a_9d289b8,R_2553c_96e06a8,R_25540_95358f8,R_25542_96e0750,R_25544_96e0b40,R_25546_96e0be8,
        R_25548_96e0c90,R_2554a_96e0d38,R_2554c_95359a0,R_2554e_9d28a60,R_25550_96e0e88,R_25552_9535a48,R_25556_96e0f30,R_25558_9535b98,R_2555a_9d28c58,R_2555c_96e0fd8,
        R_2555e_9d28d00,R_25560_9535c40,R_25562_95362d0,R_25564_9536810,R_25566_9536a08,R_25568_96e1080,R_2556c_96e1128,R_2556e_9d28ef8,R_25570_96e11d0,R_25572_96e1c50,
        R_2557c_9591d48,R_25592_9591df0,R_255a8_96e2e08,R_255be_9591e98,R_255d4_9591f40,R_255ea_96e3690,R_255f4_96e6918,R_255f6_96e69c0,R_255f8_9d29048,R_255fa_9d28718,
        R_2557e_9591fe8,R_25580_96e6fa8,R_25582_96e72f0,R_25584_9d287c0,R_25586_9592090,R_25588_9592138,R_2558a_96e7398,R_2558c_9d28868,R_2558e_9d290f0,R_25590_9d29240,
        R_25594_96e7cc8,R_25596_95921e0,R_25598_9592288,R_2559a_9592330,R_2559c_96e82b0,R_2559e_9d292e8,R_255a0_9d2dfb0,R_255a2_9592528,R_255a4_9592678,R_255a6_9d2e058,
        R_255aa_96e8358,R_255ac_9592918,R_255ae_96e86a0,R_255b0_9d2e988,R_255b2_9d29390,R_255b4_9d2ec28,R_255b6_9d294e0,R_255b8_9d2f360,R_255ba_9592a68,R_255bc_9592b10,
        R_255c0_9d30128,R_255c2_9592c60,R_255c4_96e8940,R_255c6_96e89e8,R_255c8_9d30278,R_255ca_96e8be0,R_255cc_9592f00,R_255ce_9d29588,R_255d0_9d296d8,R_255d2_9d30518,
        R_255d6_9d29828,R_255d8_96e9120,R_255da_96e93c0,R_255dc_96e9510,R_255de_9d307b8,R_255e0_9d29cc0,R_255e2_9592fa8,R_255e4_9593050,R_255e6_96e9858,R_255e8_96e9a50,
        R_255ec_95930f8,R_255ee_9d29eb8,R_255f0_96ea038,R_255f2_95931a0,R_253bc_96eacb0,R_253be_9593248,R_253c0_9d29f60,R_253c2_95932f0,R_253c4_96eae00,R_253c6_9536b58,
        R_253c8_9593398,R_253ca_9d2a350,R_253cc_b7dc210,R_253ce_b7dcd38,R_253d0_b7dcde0,R_253d2_9593590,R_253d4_96376b8,R_253d6_9d2a4a0,R_253d8_9596038,R_253da_b7dc2b8,
        R_253dc_96eb0a0,R_253de_9596578,R_253e0_9536f48,R_253e2_96eb298,R_253e4_9537098,R_253e6_96eb340,R_253e8_95373e0,R_253ea_9596a10,R_253ec_9d30860,R_253ee_9ef0090,
        R_253f0_9d30f98,R_253f2_9ef05d0,R_253f4_9d31040,R_253f6_9d31238,R_253f8_9d314d8,R_253fa_9d316d0,R_25666_96346d0,R_1a4_b821b50,R_1a3_b821aa8,R_23ca4_96329f0,
        R_23cba_9f596e0,R_23cd0_962b7c0,R_23ce6_955f268,R_23cfc_9f5c4d0,R_23d12_9d225e8,R_23d1c_962b910,R_23d1e_95a3470,R_23d20_9632c90,R_23d22_95a3710,R_23ca6_9ee76c0,
        R_23ca8_9ee7810,R_23caa_9ee78b8,R_23cac_9ee8140,R_23cae_962bbb0,R_23cb0_9ee8920,R_23cb2_9d22d20,R_23cb4_9ee8bc0,R_23cb6_9632d38,R_23cb8_9d23110,R_23cbc_962bc58,
        R_23cbe_9ee9ad8,R_23cc0_9d23260,R_23cc2_9632f30,R_23cc4_9eec430,R_23cc6_9d23308,R_23cc8_9eef4c0,R_23cca_9eefca0,R_23ccc_9d23650,R_23cce_9ef0678,R_23cd2_95a3908,
        R_23cd4_962bd00,R_23cd6_9632fd8,R_23cd8_962be50,R_23cda_96331d0,R_23cdc_962bef8,R_23cde_9d30ef0,R_23ce0_9d238f0,R_23ce2_9d23b90,R_23ce4_962bfa0,R_23ce8_962c048,
        R_23cea_95a3a58,R_23cec_9d23ed8,R_23cee_9ef09c0,R_23cf0_9ef4380,R_23cf2_95a3ba8,R_23cf4_9ef4a10,R_23cf6_962c0f0,R_23cf8_96c3060,R_23cfa_96c6d68,R_23cfe_9d310e8,
        R_23d00_96c72a8,R_23d02_962c390,R_23d04_96c74a0,R_23d06_962da88,R_23d08_9d24178,R_23d0a_962df20,R_23d0c_9633278,R_23d0e_9633320,R_23d10_95a3e48,R_23d14_95a4040,
        R_23d16_9d24370,R_23d18_96c7e78,R_23d1a_96333c8,R_23d24_9633470,R_23d3a_9633518,R_23d50_962dfc8,R_23d66_9629b88,R_23d7c_95547c8,R_23d92_96335c0,R_23d9c_96337b8,
        R_23d9e_9633908,R_23da0_9633a58,R_23da2_962e7a8,R_23d26_9554870,R_23d28_962a560,R_23d2a_962ee38,R_23d2c_962a8a8,R_23d2e_962f2d0,R_23d30_95549c0,R_23d32_9633cf8,
        R_23d34_962f4c8,R_23d36_9633da0,R_23d38_9633e48,R_23d3c_9633ef0,R_23d3e_962c4e0,R_23d40_9554bb8,R_23d42_9554d08,R_23d44_9634040,R_23d46_962f6c0,R_23d48_9554f00,
        R_23d4a_962c8d0,R_23d4c_9635000,R_23d4e_962fab0,R_23d52_95552f0,R_23d54_96350a8,R_23d56_96351f8,R_23d58_962fc00,R_23d5a_95554e8,R_23d5c_9555638,R_23d5e_9635540,
        R_23d60_96355e8,R_23d62_9635738,R_23d64_96359d8,R_23d68_962ca20,R_23d6a_9635f18,R_23d6c_962ff48,R_23d6e_9636068,R_23d70_96363b0,R_23d72_9636ae8,R_23d74_9637220,
        R_23d76_9637e98,R_23d78_9638b10,R_23d7a_962d4a0,R_23d7e_96305d8,R_23d80_9638bb8,R_23d82_9638fa8,R_23d84_962d548,R_23d86_9639398,R_23d88_95556e0,R_23d8a_9639440,
        R_23d8c_9d18d00,R_23d8e_9d19d68,R_23d90_9630a70,R_23d94_9d1a008,R_23d96_9d1a350,R_23d98_9d1a9e0,R_23d9a_96314f0,R_23da4_9634430,R_23dba_95558d8,R_23dd0_9555a28,
        R_23de6_9d1ac80,R_23dfc_962d9e0,R_23e12_9555b78,R_23e1c_96344d8,R_23e1e_9555e18,R_23e20_9d1b070,R_23e22_9d1b8f8,R_23da6_9634a18,R_23da8_9555f68,R_23daa_9635150,
        R_23dac_96352a0,R_23dae_9556010,R_23db0_9557078,R_23db2_96353f0,R_23db4_9d1ba48,R_23db6_962db30,R_23db8_96357e0,R_23dbc_9559730,R_23dbe_955bde8,R_23dc0_955dd68,
        R_23dc2_9d1baf0,R_23dc4_955e158,R_23dc6_9638db0,R_23dc8_9d1bb98,R_23dca_9639248,R_23dcc_9d1bce8,R_23dce_96c81c0,R_23dd2_955e4a0,R_23dd4_955ea88,R_23dd6_96392f0,
        R_23dd8_9d15d18,R_23dda_955ee78,R_23ddc_9d168e8,R_23dde_9d16ae0,R_23de0_962e310,R_23de2_9d16c30,R_23de4_9d16e28,R_23de8_9d170c8,R_23dea_955f1c0,R_23dec_96c87a8,
        R_23dee_955f310,R_23df0_9d1bee0,R_23df2_955f3b8,R_23df4_95a39b0,R_23df6_96c8af0,R_23df8_95a3b00,R_23dfa_95a40e8,R_23dfe_95a44d8,R_23e00_9d1bf88,R_23e02_95a4580,
        R_23e04_95a4c10,R_23e06_9d17218,R_23e08_95a5348,R_23e0a_962ec40,R_23e0c_9d17608,R_23e0e_95a57e0,R_23e10_95a5930,R_23e14_9d18910,R_23e16_9d19630,R_23e18_95a5c78,
        R_23e1a_95a6260,R_23e24_9d1c030,R_23e3a_95a4628,R_23e50_95a48c8,R_23e66_95a4b68,R_23e7c_95b1438,R_23e92_9d19780,R_23e9c_95a6d88,R_23e9e_95b1780,R_23ea0_95a7028,
        R_23ea2_95a70d0,R_23e26_95b1828,R_23e28_95a7220,R_23e2a_95b2bd8,R_23e2c_95b3310,R_23e2e_95818b0,R_23e30_9582138,R_23e32_9582288,R_23e34_95a7760,R_23e36_9582870,
        R_23e38_95a78b0,R_23e3c_9d1c0d8,R_23e3e_9582a68,R_23e40_9d1b118,R_23e42_9582e58,R_23e44_9582f00,R_23e46_95830f8,R_23e48_958cbd8,R_23e4a_958cc80,R_23e4c_95a7aa8,
        R_23e4e_958f5d8,R_23e52_958f920,R_23e54_9590058,R_23e56_95a7bf8,R_23e58_95a7ca0,R_23e5a_95901a8,R_23e5c_959fdb8,R_23e5e_95a0b80,R_23e60_9d1c4c8,R_23e62_9625b28,
        R_23e64_96261b8,R_23e68_9d1b268,R_23e6a_9d1c570,R_23e6c_95a7d48,R_23e6e_9626458,R_23e70_95a8090,R_23e72_9628330,R_23e74_9628480,R_23e76_9628528,R_23e78_95a8138,
        R_23e7a_96285d0,R_23e7e_9628720,R_23e80_9628bb8,R_23e82_962c198,R_23e84_9d1c618,R_23e86_95a8288,R_23e88_9634238,R_23e8a_9d1c6c0,R_23e8c_96342e0,R_23e8e_9634970,
        R_23e90_9d1c8b8,R_23e94_9639830,R_23e96_9d159d0,R_23e98_9d15e68,R_23e9a_95a83d8,R_23c64_96c9a08,R_23c66_9d1b658,R_23c68_96ca920,R_23c6a_9d244c0,R_23c6c_96cb4f0,
        R_23c6e_9d1b700,R_23c70_9d1ca08,R_23c72_96cb640,R_23c74_962f030,R_23c76_9d1cc00,R_23c78_9d1cd50,R_23c7a_9d1cdf8,R_23c7c_9d1b7a8,R_23c7e_9d1cf48,R_23c80_9d1d098,
        R_23c82_9d1d1e8,R_23c84_95a8528,R_23c86_9d1b9a0,R_23c88_95a8720,R_23c8a_9d1be38,R_23c8c_9d246b8,R_23c8e_96cb838,R_23c90_9d24760,R_23c92_9d1c2d0,R_23c94_9d1d3e0,
        R_23c96_95a87c8,R_23c98_9d19438,R_23c9a_9d1c378,R_23c9c_9d1c768,R_23c9e_9d1d488,R_23ca0_9d1c960,R_23ca2_9d1e8e0,R_23ebc_9667ae0,R_23ebe_965f6f8,R_23ec0_9667b88,
        R_23ec2_96688a8,R_23ec4_95ac230,R_23ec6_95ac428,R_23ec8_966a780,R_23eca_966a8d0,R_23eba_965f8f0,R_23ecc_95ac620,R_23ece_95ac770,R_23ed0_966a978,R_23ed2_966aa20,
        R_23eb8_966aac8,R_23eea_95b1588,R_23eec_9d1e448,R_23eee_9d1e790,R_23a0c_95b1630,R_23a22_95b1c18,R_23a38_966acc0,R_23a4e_95b1d68,R_23a64_966ad68,R_23a7a_95b2c80,
        R_23a84_9661a68,R_23a86_9d1d7d0,R_23a88_966ae10,R_23a8a_966b0b0,R_23a0e_962f420,R_23a10_966ba88,R_23a12_95b2fc8,R_23a14_9d1f6a8,R_23a16_952daf8,R_23a18_95b3268,
        R_23a1a_9581220,R_23a1c_9d1d878,R_23a1e_9663160,R_23a20_9d1e250,R_23a24_9d1fb40,R_23a26_95305a0,R_23a28_95812c8,R_23a2a_9530798,R_23a2c_95816b8,R_23a2e_9663550,
        R_23a30_9531e90,R_23a32_9531f38,R_23a34_9532130,R_23a36_9532280,R_23a3a_9532328,R_23a3c_9581760,R_23a3e_9581f40,R_23a40_95323d0,R_23a42_9532868,R_23a44_9582720,
        R_23a46_9532b08,R_23a48_9532c58,R_23a4a_9582918,R_23a4c_966a4e0,R_23a50_9532e50,R_23a52_9d24808,R_23a54_9533390,R_23a56_9d20668,R_23a58_9582db0,R_23a5a_9583050,
        R_23a5c_9533978,R_23a5e_9534158,R_23a60_9d20710,R_23a62_95349e0,R_23a66_9537290,R_23a68_9d1f750,R_23a6a_966a6d8,R_23a6c_966aeb8,R_23a6e_966b158,R_23a70_9537a70,
        R_23a72_9539f30,R_23a74_95831a0,R_23a76_9537c68,R_23a78_9d20a58,R_23a7c_9537d10,R_23a7e_9537e60,R_23a80_9538250,R_23a82_95382f8,R_23a8c_9d21e08,R_23aa2_9583440,
        R_23ab8_9d1f8a0,R_23ace_9d1ff30,R_23ae4_9d23ce0,R_23afa_95834e8,R_23b04_9583590,R_23b06_9d20860,R_23b08_9d24958,R_23b0a_9d24ca0,R_23a8e_95836e0,R_23a90_9583e18,
        R_23a92_9d25288,R_23a94_9d20908,R_23a96_9d25330,R_23a98_9d22348,R_23a9a_9d253d8,R_23a9c_9d233b0,R_23a9e_9d25528,R_23aa0_9d255d0,R_23aa4_9d23500,R_23aa6_9d25678,
        R_23aa8_9d23a40,R_23aaa_9d24610,R_23aac_9d25880,R_23aae_9d248b0,R_23ab0_9d26258,R_23ab2_9584898,R_23ab4_9d24a00,R_23ab6_9d26450,R_23aba_9d26648,R_23abc_9d26e28,
        R_23abe_9d270c8,R_23ac0_9584c88,R_23ac2_9d24aa8,R_23ac4_9d24d48,R_23ac6_9585270,R_23ac8_9585708,R_23aca_9d27bf0,R_23acc_9d28910,R_23ad0_9d29198,R_23ad2_9d29630,
        R_23ad4_9d24fe8,R_23ad6_95857b0,R_23ad8_9d2a0b0,R_23ada_9585900,R_23adc_9d2a200,R_23ade_9d2a3f8,R_23ae0_9d2a7e8,R_23ae2_9d25138,R_23ae6_9d2ad28,R_23ae8_95860e0,
        R_23aea_9d25480,R_23aec_9d25928,R_23aee_9d25bc8,R_23af0_95864d0,R_23af2_9d25e68,R_23af4_95866c8,R_23af6_9586770,R_23af8_9587688,R_23afc_9d26ed0,R_23afe_9587730,
        R_23b00_9d27aa0,R_23b02_9d2add0,R_23b0c_95877d8,R_23b22_95386e8,R_23b38_95388e0,R_23b4e_9588108,R_23b64_9538ad8,R_23b7a_9d2b118,R_23b84_95881b0,R_23b86_95899f8,
        R_23b88_9589aa0,R_23b8a_9d2b460,R_23b0e_958d268,R_23b10_95390c0,R_23b12_9539168,R_23b14_95394b0,R_23b16_95399f0,R_23b18_9539c90,R_23b1a_953ba18,R_23b1c_953bac0,
        R_23b1e_958d460,R_23b20_9d2b508,R_23b24_953bf58,R_23b26_953c0a8,R_23b28_953c1f8,R_23b2a_953c540,R_23b2c_9d2b5b0,R_23b2e_953c888,R_23b30_953cdc8,R_23b32_958da48,
        R_23b34_9d2b700,R_23b36_953cf18,R_23b3a_958de38,R_23b3c_958e180,R_23b3e_96ddca8,R_23b40_96dddf8,R_23b42_958e570,R_23b44_958e810,R_23b46_96de098,R_23b48_9d285c8,
        R_23b4a_96de3e0,R_23b4c_9d28b08,R_23b50_96de530,R_23b52_958ef48,R_23b54_9d24b50,R_23b56_9d25d18,R_23b58_958ff08,R_23b5a_96e6c60,R_23b5c_96e8160,R_23b5e_96ebc70,
        R_23b60_95903a0,R_23b62_95906e8,R_23b66_96ebdc0,R_23b68_95efb90,R_23b6a_9596d58,R_23b6c_9d2b7a8,R_23b6e_9598c30,R_23b70_95f0220,R_23b72_9598cd8,R_23b74_95f1918,
        R_23b76_9599170,R_23b78_9d28bb0,R_23b7c_95f37f0,R_23b7e_95f41c8,R_23b80_95f4318,R_23b82_95992c0,R_23b8c_9599608,R_23ba2_9599758,R_23bb8_9599800,R_23bce_9599950,
        R_23be4_962f570,R_23bfa_9599b48,R_23c04_959a088,R_23c06_959a130,R_23c08_959a1d8,R_23c0a_962f618,R_23b8e_959a5c8,R_23b90_959a9b8,R_23b92_959ac58,R_23b94_959aef8,
        R_23b96_962f8b8,R_23b98_959afa0,R_23b9a_959b048,R_23b9c_959b0f0,R_23b9e_959b198,R_23ba0_959b240,R_23ba4_959b6d8,R_23ba6_959b828,R_23ba8_959b8d0,R_23baa_959ba20,
        R_23bac_9d28da8,R_23bae_959bac8,R_23bb0_959d268,R_23bb2_959d508,R_23bb4_959dce8,R_23bb6_959e420,R_23bba_9d28fa0,R_23bbc_962f960,R_23bbe_9d298d0,R_23bc0_959e618,
        R_23bc2_959eea0,R_23bc4_959f098,R_23bc6_9d29978,R_23bc8_9d25dc0,R_23bca_959f9c8,R_23bcc_9d29a20,R_23bd0_95a0e20,R_23bd2_9d29b70,R_23bd4_962fb58,R_23bd6_95a0f70,
        R_23bd8_9d29c18,R_23bda_9619ae0,R_23bdc_9619b88,R_23bde_9619d80,R_23be0_9619e28,R_23be2_961a020,R_23be6_961a0c8,R_23be8_961a218,R_23bea_961a4b8,R_23bec_961a800,
        R_23bee_961a8a8,R_23bf0_961a950,R_23bf2_961ad40,R_23bf4_961ade8,R_23bf6_961ae90,R_23bf8_961af38,R_23bfc_9d26060,R_23bfe_961b088,R_23c00_9d29d68,R_23c02_961b1d8,
        R_239cc_95f4af8,R_239ce_962fd50,R_239d0_9558e00,R_239d2_9d261b0,R_239d4_95f52d8,R_239d6_9558ea8,R_239d8_961b670,R_239da_95f5620,R_239dc_961b910,R_239de_9d2b850,
        R_239e0_9d2b9a0,R_239e2_9d29e10,R_239e4_9d2a158,R_239e6_961bb08,R_239e8_961c978,R_239ea_961cd68,R_239ec_9d2baf0,R_239ee_95f5968,R_239f0_95f5ab8,R_239f2_9d2a2a8,
        R_239f4_961ce10,R_239f6_9634e08,R_239f8_9d2bb98,R_239fa_9d2bd90,R_239fc_962fdf8,R_239fe_962fea0,R_23a00_961d200,R_23a02_961d5f0,R_23a04_961d698,R_23a06_962fff0,
        R_23a08_961d740,R_23a0a_961d938,R_23c24_9d2a698,R_23c26_9d2c420,R_23c28_962ac98,R_23c2a_9d2c4c8,R_23c2c_9d2c570,R_23c2e_95f63e8,R_23c30_9d2a890,R_23c32_962ad40,
        R_23c22_9d2aa88,R_23c34_9d2c810,R_23c36_9d2ab30,R_23c38_9d2c8b8,R_23c3a_9d2cab0,R_23c20_9635e70,R_23c52_962b868,R_23c54_9d2af20,R_23c56_9d2b310,R_23774_9630098,
        R_2378a_962b9b8,R_237a0_9d2cd50,R_237b6_962bb08,R_237cc_9d2cff0,R_237e2_9d2d098,R_237ec_9d2d140,R_237ee_9d2d290,R_237f0_962c240,R_237f2_9559688,R_23776_96301e8,
        R_23778_9d2d7d0,R_2377a_962c2e8,R_2377c_9d2d878,R_2377e_962ce10,R_23780_9d2d920,R_23782_962d938,R_23784_962e5b0,R_23786_9d2d9c8,R_23788_9d2dc68,R_2378c_9d2dd10,
        R_2378e_9d2ddb8,R_23790_9d2e100,R_23792_9d2e1a8,R_23794_9d2f0c0,R_23796_9630290,R_23798_96303e0,R_2379a_9d2f210,R_2379c_9d2f7f8,R_2379e_9630728,R_237a2_96307d0,
        R_237a4_9d2fb40,R_237a6_9d301d0,R_237a8_9559bc8,R_237aa_9630140,R_237ac_96312f8,R_237ae_9d30710,R_237b0_9630b18,R_237b2_9630c68,R_237b4_9d309b0,R_237b8_9630d10,
        R_237ba_9630fb0,R_237bc_9631100,R_237be_9d30a58,R_237c0_9d30da0,R_237c2_96311a8,R_237c4_96313a0,R_237c6_96318e0,R_237c8_9631a30,R_237ca_9d30e48,R_237ce_9d31190,
        R_237d0_9631b80,R_237d2_9d31f58,R_237d4_9631448,R_237d6_9631790,R_237d8_9d323f0,R_237da_9631ad8,R_237dc_9d32540,R_237de_9632018,R_237e0_9631cd0,R_237e4_9632210,
        R_237e6_9d32690,R_237e8_96322b8,R_237ea_9d32888,R_237f4_9631e20,R_2380a_9d329d8,R_23820_9d32a80,R_23836_9d32f18,R_2384c_9d2b3b8,R_23862_9631ec8,R_2386c_9632360,
        R_2386e_9632a98,R_23870_9d32fc0,R_23872_9632408,R_237f6_9632600,R_237f8_9d33500,R_237fa_96326a8,R_237fc_9d33650,R_237fe_9d336f8,R_23800_9d33a40,R_23802_9632750,
        R_23804_96328a0,R_23806_9d340d0,R_23808_9632948,R_2380c_9d2b658,R_2380e_9d34418,R_23810_9d34760,R_23812_9d34fe8,R_23814_9632de0,R_23816_9632e88,R_23818_9d35720,
        R_2381a_9d2bc40,R_2381c_b805670,R_2381e_b805868,R_23822_9633080,R_23824_b8060f0,R_23826_9633128,R_23828_9633b00,R_2382a_9632b40,R_2382c_9634190,R_2382e_9638720,
        R_23830_9d2c180,R_23832_96389c0,R_23834_9638a68,R_23838_9d15880,R_2383a_b806198,R_2383c_9d2c768,R_2383e_9d16a38,R_23840_9d2ca08,R_23842_b806240,R_23844_9d17170,
        R_23846_9d17c98,R_23848_b8062e8,R_2384a_b806390,R_2384e_9d2cca8,R_23850_9d17fe0,R_23852_9d18328,R_23854_9d2d1e8,R_23856_9d1fd38,R_23858_b8064e0,R_2385a_9d2d3e0,
        R_2385c_9d220a8,R_2385e_9535d90,R_23860_b806588,R_23864_9d25720,R_23866_b8066d8,R_23868_b806780,R_2386a_9d2d530,R_23874_95f7840,R_2388a_95f7e28,R_238a0_9d28e50,
        R_238b6_95f8170,R_238cc_95fcd90,R_238e2_95fda08,R_238ec_95fdb58,R_238ee_95fdca8,R_238f0_95fdd50,R_238f2_9d2d728,R_23876_95ff6e8,R_23878_9535e38,R_2387a_9633668,
        R_2387c_9f4ddd0,R_2387e_9f51b80,R_23880_9f51e20,R_23882_9d29ac8,R_23884_9f53278,R_23886_9f53320,R_23888_9f54580,R_2388c_9f54778,R_2388e_9d2dbc0,R_23890_9d2e250,
        R_23892_9f548c8,R_23894_9f54970,R_23896_9f54c10,R_23898_9f55348,R_2389a_9f55498,R_2389c_9d2a740,R_2389e_9d2e3a0,R_238a2_9d2b070,R_238a4_9633710,R_238a6_9f55b28,
        R_238a8_9f56260,R_238aa_9f56500,R_238ac_9f5baf8,R_238ae_9ee9d78,R_238b0_9d2ba48,R_238b2_9d2bce8,R_238b4_9eea0c0,R_238b8_9eeb518,R_238ba_9eedf18,R_238bc_9eee6f8,
        R_238be_9ef2010,R_238c0_9537530,R_238c2_9ef2208,R_238c4_9ef3660,R_238c6_9ef3858,R_238c8_9633860,R_238ca_9ef3a50,R_238ce_9ef3af8,R_238d0_9ef3ba0,R_238d2_9ef3c48,
        R_238d4_9ef4620,R_238d6_9d2c2d0,R_238d8_9ef4770,R_238da_9d2cb58,R_238dc_9ef4ab8,R_238de_9ef4c08,R_238e0_9ef4ff8,R_238e4_9ef5148,R_238e6_9ef51f0,R_238e8_9d2cf48,
        R_238ea_9ef53e8,R_238f4_9d2e4f0,R_2390a_96339b0,R_23920_9633c50,R_23936_9d266f0,R_2394c_9d2e838,R_23962_9d2ecd0,R_2396c_9d2ed78,R_2396e_9d2f018,R_23970_9d2f168,
        R_23972_b8068d0,R_238f6_9d2f2b8,R_238f8_9d2f9f0,R_238fa_9d2fde0,R_238fc_9633f98,R_238fe_b806a20,R_23900_96340e8,R_23902_9d30320,R_23904_9634580,R_23906_9d305c0,
        R_23908_9634b68,R_2390c_9d30ba8,R_2390e_9d30c50,R_23910_b806ac8,R_23912_9d32000,R_23914_b806b70,R_23916_9d320a8,R_23918_9634c10,R_2391a_9d32150,R_2391c_9634cb8,
        R_2391e_9d32498,R_23922_9d32738,R_23924_9d327e0,R_23926_9d32b28,R_23928_9d32bd0,R_2392a_9635348,R_2392c_9635690,R_2392e_9d32c78,R_23930_9d32d20,R_23932_9635a80,
        R_23934_9d32dc8,R_23938_9d331b8,R_2393a_9d2d488,R_2393c_9d333b0,R_2393e_9d335a8,R_23940_9d337a0,R_23942_9635b28,R_23944_9d2d5d8,R_23946_9d338f0,R_23948_9635bd0,
        R_2394a_9d33998,R_2394e_9d33ae8,R_23950_9d33b90,R_23952_9636110,R_23954_9d33ce0,R_23956_b806c18,R_23958_9d33ed8,R_2395a_9d33f80,R_2395c_9636308,R_2395e_b806cc0,
        R_23960_9d34028,R_23964_9d34178,R_23966_9d2db18,R_23968_96365a8,R_2396a_9636848,R_23734_96368f0,R_23736_9636998,R_23738_9636a40,R_2373a_b7dc0c0,R_2373c_9636b90,
        R_2373e_9636c38,R_23740_b7dc168,R_23742_b806d68,R_23744_b806e10,R_23746_9636ed8,R_23748_b806eb8,R_2374a_9637028,R_2374c_b806f60,R_2374e_b8070b0,R_23750_9d33308,
        R_23752_b807158,R_23754_9ef5880,R_23756_9d26798,R_23758_9d342c8,R_2375a_9ef5928,R_2375c_96c2b20,R_2375e_9d31820,R_23760_9d31970,R_23762_9637178,R_23764_9d26840,
        R_23766_96372c8,R_23768_9d268e8,R_2376a_9d26a38,R_2376c_9d26ae0,R_2376e_9637370,R_23770_9d26b88,R_23772_9637418,R_2398c_96c2fb8,R_2398e_9559c70,R_23990_96c35a0,
        R_23992_96e8010,R_23994_955a300,R_23996_955a450,R_23998_9d34ca0,R_2399a_96c3840,R_2398a_9d34d48,R_2399c_96c3a38,R_2399e_96c3d80,R_239a0_955a840,R_239a2_96c59b8,
        R_23988_96eaf50,R_239ba_96ca728,R_239bc_955b8a8,R_239be_b7db6e8,R_234dc_b8085b0,R_234f2_b80b988,R_23508_b808658,R_2351e_b808700,R_23534_b8087a8,R_2354a_b8088f8,
        R_23554_b80ba30,R_23556_b80bb80,R_23558_b80bec8,R_2355a_b80bf70,R_234de_b8089a0,R_234e0_b808a48,R_234e2_b809768,R_234e4_b809df8,R_234e6_b80c2b8,R_234e8_b80e040,
        R_234ea_b80e580,R_234ec_b80c600,R_234ee_b80f0a8,R_234f0_b80fd20,R_234f4_b80c750,R_234f6_b80ffc0,R_234f8_b7ddf98,R_234fa_b80c7f8,R_234fc_b7de0e8,R_234fe_b7de388,
        R_23500_b7de430,R_23502_b80c9f0,R_23504_b7de580,R_23506_b80ca98,R_2350a_b7de820,R_2350c_b7dea18,R_2350e_b7dee08,R_23510_b80cc90,R_23512_b80cd38,R_23514_b7df1f8,
        R_23516_b80ce88,R_23518_b7df348,R_2351a_b7df540,R_2351c_b80cf30,R_23520_b7dfc78,R_23522_b80d080,R_23524_b80d278,R_23526_b7dff18,R_23528_b80d320,R_2352a_b7e0068,
        R_2352c_b80d5c0,R_2352e_b7e01b8,R_23530_b80d668,R_23532_b7e0458,R_23536_b7e05a8,R_23538_b80d7b8,R_2353a_b80de48,R_2353c_b7e0998,R_2353e_b7e0b90,R_23540_b7e1178,
        R_23542_b80e430,R_23544_b80e628,R_23546_b80e778,R_23548_b7e1568,R_2354c_b80e970,R_2354e_b7e16b8,R_23550_b80eb68,R_23552_b7e1808,R_2355c_b7e18b0,R_23572_b805c58,
        R_23588_b7e1958,R_2359e_b80ed60,R_235b4_95ad7d8,R_235ca_b806438,R_235d4_b7e1a00,R_235d6_b80f000,R_235d8_b7e1bf8,R_235da_b7e1ca0,R_2355e_b7e1e98,R_23560_95ad9d0,
        R_23562_b7e1f40,R_23564_95adb20,R_23566_b7e1fe8,R_23568_b80f3f0,R_2356a_b80f5e8,R_2356c_b806630,R_2356e_b7e2090,R_23570_b80f690,R_23574_b7e2138,R_23576_b7e21e0,
        R_23578_b7e23d8,R_2357a_b7e2720,R_2357c_b7e2870,R_2357e_b7e29c0,R_23580_b806828,R_23582_b7e2a68,R_23584_b7e2c60,R_23586_b7e2f00,R_2358a_b80f7e0,R_2358c_96cb8e0,
        R_2358e_b7e2fa8,R_23590_b7e30f8,R_23592_b806978,R_23594_b807008,R_23596_b7e32f0,R_23598_b80fb28,R_2359a_b7e3398,R_2359c_b807698,R_235a0_b7e34e8,R_235a2_96cbb80,
        R_235a4_b80fbd0,R_235a6_96cc018,R_235a8_95adf10,R_235aa_b7e36e0,R_235ac_b807890,R_235ae_b7e3788,R_235b0_b7e38d8,R_235b2_b7e3ad0,R_235b6_b7e3cc8,R_235b8_b7e3f68,
        R_235ba_b807f20,R_235bc_b807fc8,R_235be_b8101b8,R_235c0_b7e40b8,R_235c2_b7e4208,R_235c4_b8105a8,R_235c6_b810650,R_235c8_96cc210,R_235cc_b7e42b0,R_235ce_b7e4400,
        R_235d0_b7e4550,R_235d2_b7e45f8,R_235dc_b8106f8,R_235f2_b7e46a0,R_23608_b808118,R_2361e_b7e47f0,R_23634_b7e49e8,R_2364a_b7dd860,R_23654_95ae060,R_23656_b7dd908,
        R_23658_b7ddda0,R_2365a_b7dde48,R_235de_9637b50,R_235e0_95ae1b0,R_235e2_b7ddef0,R_235e4_b7de238,R_235e6_b7e4b38,R_235e8_9637fe8,R_235ea_b7de2e0,R_235ec_b808310,
        R_235ee_9638138,R_235f0_96381e0,R_235f4_b7e4d30,R_235f6_96383d8,R_235f8_b7de6d0,R_235fa_9638480,R_235fc_b7de8c8,R_235fe_9638528,R_23600_96385d0,R_23602_b7de970,
        R_23604_b7deac0,R_23606_9638678,R_2360a_96387c8;

wire \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 ,
         \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 ,
         \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 ,
         \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 ,
         \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 ,
         \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 ,
         \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 ,
         \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 ,
         \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 ,
         \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 ,
         \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 ,
         \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 ,
         \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 ,
         \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 ,
         \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 ,
         \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 ,
         \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 ,
         \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 ,
         \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 ,
         \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 ,
         \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 ,
         \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 ,
         \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 ,
         \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 ,
         \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 ,
         \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 ,
         \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 ,
         \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 ,
         \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 ,
         \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 ,
         \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 ,
         \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 ,
         \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 ,
         \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 ,
         \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 ,
         \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 ,
         \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 ,
         \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 ,
         \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 ,
         \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 ,
         \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 ,
         \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 ,
         \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 ,
         \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 ,
         \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 ,
         \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 ,
         \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 ,
         \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 ,
         \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 ,
         \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 ,
         \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 ,
         \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 ,
         \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 ,
         \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 ,
         \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 ,
         \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 ,
         \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 ,
         \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 ,
         \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 ,
         \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 ,
         \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 ,
         \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 ,
         \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 ,
         \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 ,
         \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 ,
         \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 ,
         \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 ,
         \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 ,
         \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 ,
         \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 ,
         \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 ,
         \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 ,
         \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 ,
         \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 ,
         \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 ,
         \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 ,
         \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 ,
         \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 ,
         \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 ,
         \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 ,
         \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 ,
         \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 ,
         \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 ,
         \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 ,
         \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 ,
         \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 ,
         \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 ,
         \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 ,
         \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 ,
         \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 ,
         \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 ,
         \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 ,
         \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 ,
         \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 ,
         \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 ,
         \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 ,
         \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 ,
         \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 ,
         \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 ,
         \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 ,
         \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 ,
         \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 ,
         \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 ,
         \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 ,
         \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 ,
         \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 ,
         \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 ,
         \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 ,
         \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 ,
         \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 ,
         \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 ,
         \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 ,
         \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 ,
         \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 ,
         \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 ,
         \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 ,
         \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 ,
         \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 ,
         \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 ,
         \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 ,
         \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 ,
         \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 ,
         \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 ,
         \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 ,
         \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 ,
         \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 ,
         \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 ,
         \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 ,
         \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 ,
         \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 ,
         \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 ,
         \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 ,
         \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 ,
         \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 ,
         \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 ,
         \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 ,
         \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 ,
         \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 ,
         \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671_N$1 , \4672_N$3 , \4673_N$5 , \4674_N$7 ,
         \4675_N$9 , \4676_N$11 , \4677_N$13 , \4678_N$15 , \4679_N$17 , \4680_N$19 , \4681_N$21 , \4682_N$23 , \4683_N$25 , \4684_N$27 ,
         \4685_N$29 , \4686_N$31 , \4687_N$33 , \4688_N$35 , \4689_N$37 , \4690_N$39 , \4691_N$41 , \4692_N$43 , \4693_N$45 , \4694_N$47 ,
         \4695_N$49 , \4696_N$51 , \4697_N$53 , \4698_N$55 , \4699_N$57 , \4700_N$59 , \4701_N$61 , \4702_N$63 , \4703_N$65 , \4704_N$67 ,
         \4705_N$69 , \4706_N$71 , \4707_N$73 , \4708_N$75 , \4709_N$77 , \4710_N$79 , \4711_N$81 , \4712_N$83 , \4713_N$85 , \4714_N$87 ,
         \4715_N$89 , \4716_N$91 , \4717_N$93 , \4718_N$95 , \4719_N$97 , \4720_N$99 , \4721_N$101 , \4722_N$103 , \4723_N$105 , \4724_N$107 ,
         \4725_N$109 , \4726_N$111 , \4727_N$113 , \4728_N$115 , \4729_N$117 , \4730_N$119 , \4731_N$121 , \4732_N$123 , \4733_N$125 , \4734_N$127 ,
         \4735_N$129 , \4736_N$131 , \4737_N$133 , \4738_N$135 , \4739_N$137 , \4740_N$139 , \4741_N$141 , \4742_N$143 , \4743_N$145 , \4744_N$147 ,
         \4745_N$149 , \4746_N$151 , \4747_N$153 , \4748_N$155 , \4749_N$157 , \4750_N$159 , \4751_N$161 , \4752_N$163 , \4753_N$165 , \4754_N$167 ,
         \4755_N$169 , \4756_N$171 , \4757_N$173 , \4758_N$175 , \4759_N$177 , \4760_N$179 , \4761_N$181 , \4762_N$183 , \4763_N$185 , \4764_N$187 ,
         \4765_N$189 , \4766_N$191 , \4767_N$193 , \4768_N$195 , \4769_N$197 , \4770_N$199 , \4771_N$201 , \4772_N$203 , \4773_N$205 , \4774_N$207 ,
         \4775_N$209 , \4776_N$211 , \4777_N$213 , \4778_N$215 , \4779_N$217 , \4780_N$219 , \4781_N$221 , \4782_N$223 , \4783_N$225 , \4784_N$227 ,
         \4785_N$229 , \4786_N$231 , \4787_N$233 , \4788_N$235 , \4789_N$237 , \4790_N$239 , \4791_N$241 , \4792_N$243 , \4793_N$245 , \4794_N$247 ,
         \4795_N$249 , \4796_N$251 , \4797_N$253 , \4798_N$255 , \4799_N$257 , \4800_N$259 , \4801_N$261 , \4802_N$263 , \4803_N$265 , \4804_N$267 ,
         \4805_N$269 , \4806_N$271 , \4807_N$273 , \4808_N$275 , \4809_N$277 , \4810_N$279 , \4811_N$281 , \4812_N$283 , \4813_N$285 , \4814_N$287 ,
         \4815_N$289 , \4816_N$291 , \4817_N$293 , \4818_N$295 , \4819_N$297 , \4820_N$299 , \4821_N$301 , \4822_N$303 , \4823_N$305 , \4824_N$307 ,
         \4825_N$309 , \4826_N$311 , \4827_N$313 , \4828_N$315 , \4829_N$317 , \4830_N$319 , \4831_N$321 , \4832_N$323 , \4833_N$325 , \4834_N$327 ,
         \4835_N$329 , \4836_N$331 , \4837_N$333 , \4838_N$335 , \4839_N$337 , \4840_N$339 , \4841_N$341 , \4842_N$343 , \4843_N$345 , \4844_N$347 ,
         \4845_N$349 , \4846_N$351 , \4847_N$353 , \4848_N$355 , \4849_N$357 , \4850_N$359 , \4851_N$361 , \4852_N$363 , \4853_N$365 , \4854_N$367 ,
         \4855_N$369 , \4856_N$371 , \4857_N$373 , \4858_N$375 , \4859_N$377 , \4860_N$379 , \4861_N$381 , \4862_N$383 , \4863_N$385 , \4864_N$387 ,
         \4865_N$389 , \4866_N$391 , \4867_N$393 , \4868_N$395 , \4869_N$397 , \4870_N$399 , \4871_N$401 , \4872_N$403 , \4873_N$405 , \4874_N$407 ,
         \4875_N$409 , \4876_N$411 , \4877_N$413 , \4878_N$415 , \4879_N$417 , \4880_N$419 , \4881_N$421 , \4882_N$423 , \4883_N$425 , \4884_N$427 ,
         \4885_N$429 , \4886_N$431 , \4887_N$433 , \4888_N$435 , \4889_N$437 , \4890_N$439 , \4891_N$441 , \4892_N$443 , \4893_N$445 , \4894_N$447 ,
         \4895_N$449 , \4896_N$451 , \4897_N$453 , \4898_N$455 , \4899_N$457 , \4900_N$459 , \4901_N$461 , \4902_N$463 , \4903_N$465 , \4904_N$467 ,
         \4905_N$469 , \4906_N$471 , \4907_N$473 , \4908_N$475 , \4909_N$477 , \4910_N$479 , \4911_N$481 , \4912_N$483 , \4913_N$485 , \4914_N$487 ,
         \4915_N$489 , \4916_N$491 , \4917_N$493 , \4918_N$495 , \4919_N$497 , \4920_N$499 , \4921_N$501 , \4922_N$503 , \4923_N$505 , \4924_N$507 ,
         \4925_N$509 , \4926_N$511 , \4927_N$513 , \4928_N$515 , \4929_N$517 , \4930_N$519 , \4931_N$521 , \4932_N$523 , \4933_N$525 , \4934_N$527 ,
         \4935_N$529 , \4936_N$531 , \4937_N$533 , \4938_N$535 , \4939_N$537 , \4940_N$539 , \4941_N$541 , \4942_N$543 , \4943_N$545 , \4944_N$547 ,
         \4945_N$549 , \4946_N$551 , \4947_N$553 , \4948_N$555 , \4949_N$557 , \4950_N$559 , \4951_N$561 , \4952_N$563 , \4953_N$565 , \4954_N$567 ,
         \4955_N$569 , \4956_N$571 , \4957_N$573 , \4958_N$575 , \4959_N$577 , \4960_N$579 , \4961_N$581 , \4962_N$583 , \4963_N$585 , \4964_N$587 ,
         \4965_N$589 , \4966_N$591 , \4967_N$593 , \4968_N$595 , \4969_N$597 , \4970_N$599 , \4971_N$601 , \4972_N$603 , \4973_N$605 , \4974_N$607 ,
         \4975_N$609 , \4976_N$611 , \4977_N$613 , \4978_N$615 , \4979_N$617 , \4980_N$619 , \4981_N$621 , \4982_N$623 , \4983_N$625 , \4984_N$627 ,
         \4985_N$629 , \4986_N$631 , \4987_N$633 , \4988_N$635 , \4989_N$637 , \4990_N$639 , \4991_N$641 , \4992_N$643 , \4993_N$645 , \4994_N$647 ,
         \4995_N$649 , \4996_N$651 , \4997_N$653 , \4998_N$655 , \4999_N$657 , \5000_N$659 , \5001_N$661 , \5002_N$663 , \5003_N$665 , \5004_N$667 ,
         \5005_N$669 , \5006_N$671 , \5007_N$673 , \5008_N$675 , \5009_N$677 , \5010_N$679 , \5011_N$681 , \5012_N$683 , \5013_N$685 , \5014_N$687 ,
         \5015_N$689 , \5016_N$691 , \5017_N$693 , \5018_N$695 , \5019_N$697 , \5020_N$699 , \5021_N$701 , \5022_N$703 , \5023_N$705 , \5024_N$707 ,
         \5025_N$709 , \5026_N$711 , \5027_N$713 , \5028_N$715 , \5029_N$717 , \5030_N$719 , \5031_N$721 , \5032_N$723 , \5033_N$725 , \5034_N$727 ,
         \5035_N$729 , \5036_N$731 , \5037_N$733 , \5038_N$735 , \5039_N$737 , \5040_N$739 , \5041_N$741 , \5042_N$743 , \5043_N$745 , \5044_N$747 ,
         \5045_N$749 , \5046_N$751 , \5047_N$753 , \5048_N$755 , \5049_N$757 , \5050_N$759 , \5051_N$761 , \5052_N$763 , \5053_N$765 , \5054_N$767 ,
         \5055_N$769 , \5056_N$771 , \5057_N$773 , \5058_N$775 , \5059_N$777 , \5060_N$779 , \5061_N$781 , \5062_N$783 , \5063_N$785 , \5064_N$787 ,
         \5065_N$789 , \5066_N$791 , \5067_N$793 , \5068_N$795 , \5069_N$797 , \5070_N$799 , \5071_N$801 , \5072_N$803 , \5073_N$805 , \5074_N$807 ,
         \5075_N$809 , \5076_N$811 , \5077_N$813 , \5078_N$815 , \5079_N$817 , \5080_N$819 , \5081_N$821 , \5082_N$823 , \5083_N$825 , \5084_N$827 ,
         \5085_N$829 , \5086_N$831 , \5087_N$833 , \5088_N$835 , \5089_N$837 , \5090_N$839 , \5091_N$841 , \5092_N$843 , \5093_N$845 , \5094_N$847 ,
         \5095_N$849 , \5096_N$851 , \5097_N$853 , \5098_N$855 , \5099_N$857 , \5100_N$859 , \5101_N$861 , \5102_N$863 , \5103_N$865 , \5104_N$867 ,
         \5105_N$869 , \5106_N$871 , \5107_N$873 , \5108_N$875 , \5109_N$877 , \5110_N$879 , \5111_N$881 , \5112_N$883 , \5113_N$885 , \5114_N$887 ,
         \5115_N$889 , \5116_N$891 , \5117_N$893 , \5118_N$895 , \5119_N$897 , \5120_N$899 , \5121_N$901 , \5122_N$903 , \5123_N$905 , \5124_N$907 ,
         \5125_N$909 , \5126_N$911 , \5127_N$913 , \5128_N$915 , \5129_N$917 , \5130_N$919 , \5131_N$921 , \5132_N$923 , \5133_N$925 , \5134_N$927 ,
         \5135_N$929 , \5136_N$931 , \5137_N$933 , \5138_N$935 , \5139_N$937 , \5140_N$939 , \5141_N$941 , \5142_N$943 , \5143_N$945 , \5144_N$947 ,
         \5145_N$949 , \5146_N$951 , \5147_N$953 , \5148_N$955 , \5149_N$957 , \5150_N$959 , \5151_N$961 , \5152_N$963 , \5153_N$965 , \5154_N$967 ,
         \5155_N$969 , \5156_N$971 , \5157_N$973 , \5158_N$975 , \5159_N$977 , \5160_N$979 , \5161_N$981 , \5162_N$983 , \5163_N$985 , \5164_N$987 ,
         \5165_N$989 , \5166_N$991 , \5167_N$993 , \5168_N$995 , \5169_N$997 , \5170_N$999 , \5171_N$1001 , \5172_N$1003 , \5173_N$1005 , \5174_N$1007 ,
         \5175_N$1009 , \5176_N$1011 , \5177_N$1013 , \5178_N$1015 , \5179_N$1017 , \5180_N$1019 , \5181_N$1021 , \5182_N$1023 , \5183_N$1025 , \5184_N$1027 ,
         \5185_N$1029 , \5186_N$1031 , \5187_N$1033 , \5188_N$1035 , \5189_N$1037 , \5190_N$1039 , \5191_N$1041 , \5192_N$1043 , \5193_N$1045 , \5194_N$1047 ,
         \5195_N$1049 , \5196_N$1051 , \5197_N$1053 , \5198_N$1055 , \5199_N$1057 , \5200_N$1059 , \5201_N$1061 , \5202_N$1063 , \5203_N$1065 , \5204_N$1067 ,
         \5205_N$1069 , \5206_N$1071 , \5207_N$1073 , \5208_N$1075 , \5209_N$1077 , \5210_N$1079 , \5211_N$1081 , \5212_N$1083 , \5213_N$1085 , \5214_N$1087 ,
         \5215_N$1089 , \5216_N$1091 , \5217_N$1093 , \5218_N$1095 , \5219_N$1097 , \5220_N$1099 , \5221_N$1101 , \5222_N$1103 , \5223_N$1105 , \5224_N$1107 ,
         \5225_N$1109 , \5226_N$1111 , \5227_N$1113 , \5228_N$1115 , \5229_N$1117 , \5230_N$1119 , \5231_N$1121 , \5232_N$1123 , \5233_N$1125 , \5234_N$1127 ,
         \5235_N$1129 , \5236_N$1131 , \5237_N$1133 , \5238_N$1135 , \5239_N$1137 , \5240_N$1139 , \5241_N$1141 , \5242_N$1143 , \5243_N$1145 , \5244_N$1147 ,
         \5245_N$1149 , \5246_N$1151 , \5247_N$1153 , \5248_N$1155 , \5249_N$1157 , \5250_N$1159 , \5251_N$1161 , \5252_N$1163 , \5253_N$1165 , \5254_N$1167 ,
         \5255_N$1169 , \5256_N$1171 , \5257_N$1173 , \5258_N$1175 , \5259_N$1177 , \5260_N$1179 , \5261_N$1181 , \5262_N$1183 , \5263_N$1185 , \5264_N$1187 ,
         \5265_N$1189 , \5266_N$1191 , \5267_N$1193 , \5268_N$1195 , \5269_N$1197 , \5270_N$1199 , \5271_N$1201 , \5272_N$1203 , \5273_N$1205 , \5274_N$1207 ,
         \5275_N$1209 , \5276_N$1211 , \5277_N$1213 , \5278_N$1215 , \5279_N$1217 , \5280_N$1219 , \5281_N$1221 , \5282_N$1223 , \5283_N$1225 , \5284_N$1227 ,
         \5285_N$1229 , \5286_N$1231 , \5287_N$1233 , \5288_N$1235 , \5289_N$1237 , \5290_N$1239 , \5291_N$1241 , \5292_N$1243 , \5293_N$1245 , \5294_N$1247 ,
         \5295_N$1249 , \5296_N$1251 , \5297_N$1253 , \5298_N$1255 , \5299_N$1257 , \5300_N$1259 , \5301_N$1261 , \5302_N$1263 , \5303_N$1265 , \5304_N$1267 ,
         \5305_N$1269 , \5306_N$1271 , \5307_N$1273 , \5308_N$1275 , \5309_N$1277 , \5310_N$1279 , \5311_N$1281 , \5312_N$1283 , \5313_N$1285 , \5314_N$1287 ,
         \5315_N$1289 , \5316_N$1291 , \5317_N$1293 , \5318_N$1295 , \5319_N$1297 , \5320_N$1299 , \5321_N$1301 , \5322_N$1303 , \5323_N$1305 , \5324_N$1307 ,
         \5325_N$1309 , \5326_N$1311 , \5327_N$1313 , \5328_N$1315 , \5329_N$1317 , \5330_N$1319 , \5331_N$1321 , \5332_N$1323 , \5333_N$1325 , \5334_N$1327 ,
         \5335_N$1329 , \5336_N$1331 , \5337_N$1333 , \5338_N$1335 , \5339_N$1337 , \5340_N$1339 , \5341_N$1341 , \5342_N$1343 , \5343_N$1345 , \5344_N$1347 ,
         \5345_N$1349 , \5346_N$1351 , \5347_N$1353 , \5348_N$1355 , \5349_N$1357 , \5350_N$1359 , \5351_N$1361 , \5352_N$1363 , \5353_N$1365 , \5354_N$1367 ,
         \5355_N$1369 , \5356_N$1371 , \5357_N$1373 , \5358_N$1375 , \5359_N$1377 , \5360_N$1379 , \5361_N$1381 , \5362_N$1383 , \5363_N$1385 , \5364_N$1387 ,
         \5365_N$1389 , \5366_N$1391 , \5367_N$1393 , \5368_N$1395 , \5369_N$1397 , \5370_N$1399 , \5371_N$1401 , \5372_N$1403 , \5373_N$1405 , \5374_N$1407 ,
         \5375_N$1409 , \5376_N$1411 , \5377_N$1413 , \5378_N$1415 , \5379_N$1417 , \5380_N$1419 , \5381_N$1421 , \5382_N$1423 , \5383_N$1425 , \5384_N$1427 ,
         \5385_N$1429 , \5386_N$1431 , \5387_N$1433 , \5388_N$1435 , \5389_N$1437 , \5390_N$1439 , \5391_N$1441 , \5392_N$1443 , \5393_N$1445 , \5394_N$1447 ,
         \5395_N$1449 , \5396_N$1451 , \5397_N$1453 , \5398_N$1455 , \5399_N$1457 , \5400_N$1459 , \5401_N$1461 , \5402_N$1463 , \5403_N$1465 , \5404_N$1467 ,
         \5405_N$1469 , \5406_N$1471 , \5407_N$1473 , \5408_N$1475 , \5409_N$1477 , \5410_N$1479 , \5411_N$1481 , \5412_N$1483 , \5413_N$1485 , \5414_N$1487 ,
         \5415_N$1489 , \5416_N$1491 , \5417_N$1493 , \5418_N$1495 , \5419_N$1497 , \5420_N$1499 , \5421_N$1501 , \5422_N$1503 , \5423_N$1505 , \5424_N$1507 ,
         \5425_N$1509 , \5426_N$1511 , \5427_N$1513 , \5428_N$1515 , \5429_N$1517 , \5430_N$1519 , \5431_N$1521 , \5432_N$1523 , \5433_N$1525 , \5434_N$1527 ,
         \5435_N$1529 , \5436_N$1531 , \5437_N$1533 , \5438_N$1535 , \5439_N$1537 , \5440_N$1539 , \5441_N$1541 , \5442_N$1543 , \5443_N$1545 , \5444_N$1547 ,
         \5445_N$1549 , \5446_N$1551 , \5447_N$1553 , \5448_N$1555 , \5449_N$1557 , \5450_N$1559 , \5451_N$1561 , \5452_N$1563 , \5453_N$1565 , \5454_N$1567 ,
         \5455_N$1569 , \5456_N$1571 , \5457_N$1573 , \5458_N$1575 , \5459_N$1577 , \5460_N$1579 , \5461_N$1581 , \5462_N$1583 , \5463_N$1585 , \5464_N$1587 ,
         \5465_N$1589 , \5466_N$1591 , \5467_N$1593 , \5468_N$1595 , \5469_N$1597 , \5470_N$1599 , \5471_N$1601 , \5472_N$1603 , \5473_N$1605 , \5474_N$1607 ,
         \5475_N$1609 , \5476_N$1611 , \5477_N$1613 , \5478_N$1615 , \5479_N$1617 , \5480_N$1619 , \5481_N$1621 , \5482_N$1623 , \5483_N$1625 , \5484_N$1627 ,
         \5485_N$1629 , \5486_N$1631 , \5487_N$1633 , \5488_N$1635 , \5489_N$1637 , \5490_N$1639 , \5491_N$1641 , \5492_N$1643 , \5493_N$1645 , \5494_N$1647 ,
         \5495_N$1649 , \5496_N$1651 , \5497_N$1653 , \5498_N$1655 , \5499_N$1657 , \5500_N$1659 , \5501_N$1661 , \5502_N$1663 , \5503_N$1665 , \5504_N$1667 ,
         \5505_N$1669 , \5506_N$1671 , \5507_N$1673 , \5508_N$1675 , \5509_N$1677 , \5510_N$1679 , \5511_N$1681 , \5512_N$1683 , \5513_N$1685 , \5514_N$1687 ,
         \5515_N$1689 , \5516_N$1691 , \5517_N$1693 , \5518_N$1695 , \5519_N$1697 , \5520_N$1699 , \5521_N$1701 , \5522_N$1703 , \5523_N$1705 , \5524_N$1707 ,
         \5525_N$1709 , \5526_N$1711 , \5527_N$1713 , \5528_N$1715 , \5529_N$1717 , \5530_N$1719 , \5531_N$1721 , \5532_N$1723 , \5533_N$1725 , \5534_N$1727 ,
         \5535_N$1729 , \5536_N$1731 , \5537_N$1733 , \5538_N$1735 , \5539_N$1737 , \5540_N$1739 , \5541_N$1741 , \5542_N$1743 , \5543_N$1745 , \5544_N$1747 ,
         \5545_N$1749 , \5546_N$1751 , \5547_N$1753 , \5548_N$1755 , \5549_N$1757 , \5550_N$1759 , \5551_N$1761 , \5552_N$1763 , \5553_N$1765 , \5554_N$1767 ,
         \5555_N$1769 , \5556_N$1771 , \5557_N$1773 , \5558_N$1775 , \5559_N$1777 , \5560_N$1779 , \5561_N$1781 , \5562_N$1783 , \5563_N$1785 , \5564_N$1787 ,
         \5565_N$1789 , \5566_N$1791 , \5567_N$1793 , \5568_N$1795 , \5569_N$1797 , \5570_N$1799 , \5571_N$1801 , \5572_N$1803 , \5573_N$1805 , \5574_N$1807 ,
         \5575_N$1809 , \5576_N$1811 , \5577_N$1813 , \5578_N$1815 , \5579_N$1817 , \5580_N$1819 , \5581_N$1821 , \5582_N$1823 , \5583_N$1825 , \5584_N$1827 ,
         \5585_N$1829 , \5586_N$1831 , \5587_N$1833 , \5588_N$1835 , \5589_N$1837 , \5590_N$1839 , \5591_N$1841 , \5592_N$1843 , \5593_N$1845 , \5594_N$1847 ,
         \5595_N$1849 , \5596_N$1851 , \5597_N$1853 , \5598_N$1855 , \5599_N$1857 , \5600_N$1859 , \5601_N$1861 , \5602_N$1863 , \5603_N$1865 , \5604_N$1867 ,
         \5605_N$1869 , \5606_N$1871 , \5607_N$1873 , \5608_N$1875 , \5609_N$1877 , \5610_N$1879 , \5611_N$1881 , \5612_N$1883 , \5613_N$1885 , \5614_N$1887 ,
         \5615_N$1889 , \5616_N$1891 , \5617_N$1893 , \5618_N$1895 , \5619_N$1897 , \5620_N$1899 , \5621_N$1901 , \5622_N$1903 , \5623_N$1905 , \5624_N$1907 ,
         \5625_N$1909 , \5626_N$1911 , \5627_N$1913 , \5628_N$1915 , \5629_N$1917 , \5630_N$1919 , \5631_N$1921 , \5632_N$1923 , \5633_N$1925 , \5634_N$1927 ,
         \5635_N$1929 , \5636_N$1931 , \5637_N$1933 , \5638_N$1935 , \5639_N$1937 , \5640_N$1939 , \5641_N$1941 , \5642_N$1943 , \5643_N$1945 , \5644_N$1947 ,
         \5645_N$1949 , \5646_N$1951 , \5647_N$1953 , \5648_N$1955 , \5649_N$1957 , \5650_N$1959 , \5651_N$1961 , \5652_N$1963 , \5653_N$1965 , \5654_N$1967 ,
         \5655_N$1969 , \5656_N$1971 , \5657_N$1973 , \5658_N$1975 , \5659_N$1977 , \5660_N$1979 , \5661_N$1981 , \5662_N$1983 , \5663_N$1985 , \5664_N$1987 ,
         \5665_N$1989 , \5666_N$1991 , \5667_N$1993 , \5668_N$1995 , \5669_N$1997 , \5670_N$1999 , \5671_N$2001 , \5672_N$2003 , \5673_N$2005 , \5674_N$2007 ,
         \5675_N$2009 , \5676_N$2011 , \5677_N$2013 , \5678_N$2015 , \5679_N$2017 , \5680_N$2019 , \5681_N$2021 , \5682_N$2023 , \5683_N$2025 , \5684_N$2027 ,
         \5685_N$2029 , \5686_N$2031 , \5687_N$2033 , \5688_N$2035 , \5689_N$2037 , \5690_N$2039 , \5691_N$2041 , \5692_N$2043 , \5693_N$2045 , \5694_N$2047 ,
         \5695_N$2049 , \5696_N$2051 , \5697_N$2053 , \5698_N$2055 , \5699_N$2057 , \5700_N$2059 , \5701_N$2061 , \5702_N$2063 , \5703_N$2065 , \5704_N$2067 ,
         \5705_N$2069 , \5706_N$2071 , \5707_N$2073 , \5708_N$2075 , \5709_N$2077 , \5710_N$2079 , \5711_N$2081 , \5712_N$2083 , \5713_N$2085 , \5714_N$2087 ,
         \5715_N$2089 , \5716_N$2091 , \5717_N$2093 , \5718_N$2095 , \5719_N$2097 , \5720_N$2099 , \5721_N$2101 , \5722_N$2103 , \5723_N$2105 , \5724_N$2107 ,
         \5725_N$2109 , \5726_N$2111 , \5727_N$2113 , \5728_N$2115 , \5729_N$2117 , \5730_N$2119 , \5731_N$2121 , \5732_N$2123 , \5733_N$2125 , \5734_N$2127 ,
         \5735_N$2129 , \5736_N$2131 , \5737_N$2133 , \5738_N$2135 , \5739_N$2137 , \5740_N$2139 , \5741_N$2141 , \5742_N$2143 , \5743_N$2145 , \5744_N$2147 ,
         \5745_N$2149 , \5746_N$2151 , \5747_N$2153 , \5748_N$2155 , \5749_N$2157 , \5750_N$2159 , \5751_N$2161 , \5752_N$2163 , \5753_N$2165 , \5754_N$2167 ,
         \5755_N$2169 , \5756_N$2171 , \5757_N$2173 , \5758_N$2175 , \5759_N$2177 , \5760_N$2179 , \5761_N$2181 , \5762_N$2183 , \5763_N$2185 , \5764_N$2187 ,
         \5765_N$2189 , \5766_N$2191 , \5767_N$2193 , \5768_N$2195 , \5769_N$2197 , \5770_N$2199 , \5771_N$2201 , \5772_N$2203 , \5773_N$2205 , \5774_N$2207 ,
         \5775_N$2209 , \5776_N$2211 , \5777_N$2213 , \5778_N$2215 , \5779_N$2217 , \5780_N$2219 , \5781_N$2221 , \5782_N$2223 , \5783_N$2225 , \5784_N$2227 ,
         \5785_N$2229 , \5786_N$2231 , \5787_N$2233 , \5788_N$2235 , \5789_N$2237 , \5790_N$2239 , \5791_N$2241 , \5792_N$2243 , \5793_N$2245 , \5794_N$2247 ,
         \5795_N$2249 , \5796_N$2251 , \5797_N$2253 , \5798_N$2255 , \5799_N$2257 , \5800_N$2259 , \5801_N$2261 , \5802_N$2263 , \5803_N$2265 , \5804_N$2267 ,
         \5805_N$2269 , \5806_N$2271 , \5807_N$2273 , \5808_N$2275 , \5809_N$2277 , \5810_N$2279 , \5811_N$2281 , \5812_N$2283 , \5813_N$2285 , \5814_N$2287 ,
         \5815_N$2289 , \5816_N$2291 , \5817_N$2293 , \5818_N$2295 , \5819_N$2297 , \5820_N$2299 , \5821_N$2301 , \5822_N$2303 , \5823_N$2305 , \5824_N$2307 ,
         \5825_N$2309 , \5826_N$2311 , \5827_N$2313 , \5828_N$2315 , \5829_N$2317 , \5830_N$2319 , \5831_N$2321 , \5832_N$2323 , \5833_N$2325 , \5834_N$2327 ,
         \5835_N$2329 , \5836_N$2331 , \5837_N$2333 , \5838_N$2335 , \5839_N$2337 , \5840_N$2339 , \5841_N$2341 , \5842_N$2343 , \5843_N$2345 , \5844_N$2347 ,
         \5845_N$2349 , \5846_N$2351 , \5847_N$2353 , \5848_N$2355 , \5849_N$2357 , \5850_N$2359 , \5851_N$2361 , \5852_N$2363 , \5853_N$2365 , \5854_N$2367 ,
         \5855_N$2369 , \5856_N$2371 , \5857_N$2373 , \5858_N$2375 , \5859_N$2377 , \5860_N$2379 , \5861_N$2381 , \5862_N$2383 , \5863_N$2385 , \5864_N$2387 ,
         \5865_N$2389 , \5866_N$2391 , \5867_N$2393 , \5868_N$2395 , \5869_N$2397 , \5870_N$2399 , \5871_N$2401 , \5872_N$2403 , \5873_N$2405 , \5874_N$2407 ,
         \5875_N$2409 , \5876_N$2411 , \5877_N$2413 , \5878_N$2415 , \5879_N$2417 , \5880_N$2419 , \5881_N$2421 , \5882_N$2423 , \5883_N$2425 , \5884_N$2427 ,
         \5885_N$2429 , \5886_N$2431 , \5887_N$2433 , \5888_N$2435 , \5889_N$2437 , \5890_N$2439 , \5891_N$2441 , \5892_N$2443 , \5893_N$2445 , \5894_N$2447 ,
         \5895_N$2449 , \5896_N$2451 , \5897_N$2453 , \5898_N$2455 , \5899_N$2457 , \5900_N$2459 , \5901_N$2461 , \5902_N$2463 , \5903_N$2465 , \5904_N$2467 ,
         \5905_N$2469 , \5906_N$2471 , \5907_N$2473 , \5908_N$2475 , \5909_N$2477 , \5910_N$2479 , \5911_N$2481 , \5912_N$2483 , \5913_N$2485 , \5914_N$2487 ,
         \5915_N$2489 , \5916_N$2491 , \5917_N$2493 , \5918_N$2495 , \5919_N$2497 , \5920_N$2499 , \5921_N$2501 , \5922_N$2503 , \5923_N$2505 , \5924_N$2507 ,
         \5925_N$2509 , \5926_N$2511 , \5927_N$2513 , \5928_N$2515 , \5929_N$2517 , \5930_N$2519 , \5931_N$2521 , \5932_N$2523 , \5933_N$2525 , \5934_N$2527 ,
         \5935_N$2529 , \5936_N$2531 , \5937_N$2533 , \5938_N$2535 , \5939_N$2537 , \5940_N$2539 , \5941_N$2541 , \5942_N$2543 , \5943_N$2545 , \5944_N$2547 ,
         \5945_N$2549 , \5946_N$2551 , \5947_N$2553 , \5948_N$2555 , \5949_N$2557 , \5950_N$2559 , \5951_N$2561 , \5952_N$2563 , \5953_N$2565 , \5954_N$2567 ,
         \5955_N$2569 , \5956_N$2571 , \5957_N$2573 , \5958_N$2575 , \5959_N$2577 , \5960_N$2579 , \5961_N$2581 , \5962_N$2583 , \5963_N$2585 , \5964_N$2587 ,
         \5965_N$2589 , \5966_N$2591 , \5967_N$2593 , \5968_N$2595 , \5969_N$2597 , \5970_N$2599 , \5971_N$2601 , \5972_N$2603 , \5973_N$2605 , \5974_N$2607 ,
         \5975_N$2609 , \5976_N$2611 , \5977_N$2613 , \5978_N$2615 , \5979_N$2617 , \5980_N$2619 , \5981_N$2621 , \5982_N$2623 , \5983_N$2625 , \5984_N$2627 ,
         \5985_N$2629 , \5986_N$2631 , \5987_N$2633 , \5988_N$2635 , \5989_N$2637 , \5990_N$2639 , \5991_N$2641 , \5992_N$2643 , \5993_N$2645 , \5994_N$2647 ,
         \5995_N$2649 , \5996_N$2651 , \5997_N$2653 , \5998_N$2655 , \5999_N$2657 , \6000_N$2659 , \6001_N$2661 , \6002_N$2663 , \6003_N$2665 , \6004_N$2667 ,
         \6005_N$2669 , \6006_N$2671 , \6007_N$2673 , \6008_N$2675 , \6009_N$2677 , \6010_N$2679 , \6011_N$2681 , \6012_N$2683 , \6013_N$2685 , \6014_N$2687 ,
         \6015_N$2689 , \6016_N$2691 , \6017_N$2693 , \6018_N$2695 , \6019_N$2697 , \6020_N$2699 , \6021_N$2701 , \6022_N$2703 , \6023_N$2705 , \6024_N$2707 ,
         \6025_N$2709 , \6026_N$2711 , \6027_N$2713 , \6028_N$2715 , \6029_N$2717 , \6030_N$2719 , \6031_N$2721 , \6032_N$2723 , \6033_N$2725 , \6034_N$2727 ,
         \6035_N$2729 , \6036_N$2731 , \6037_N$2733 , \6038_N$2735 , \6039_N$2737 , \6040_N$2739 , \6041_N$2741 , \6042_N$2743 , \6043_N$2745 , \6044_N$2747 ,
         \6045_N$2749 , \6046_N$2751 , \6047_N$2753 , \6048_N$2755 , \6049_N$2757 , \6050_N$2759 , \6051_N$2761 , \6052_N$2762 , \6053_N$2764 , \6054_N$2765 ,
         \6055_N$2766 , \6056_ZERO , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 ,
         \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 ,
         \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 ,
         \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 ,
         \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 ,
         \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 ,
         \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 ,
         \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 ,
         \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 ,
         \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 ,
         \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 ,
         \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 ,
         \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 ,
         \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 ,
         \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 ,
         \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 ,
         \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 ,
         \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 ,
         \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 ,
         \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 ,
         \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 ,
         \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 ,
         \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 ,
         \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 ,
         \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 ,
         \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 ,
         \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 ,
         \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 ,
         \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 ,
         \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 ,
         \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 ,
         \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 ,
         \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 ,
         \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 ,
         \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 ,
         \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 ,
         \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 ,
         \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 ,
         \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 ,
         \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 ,
         \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 ,
         \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 ,
         \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 ,
         \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 ,
         \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 ,
         \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 ,
         \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 ,
         \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 ,
         \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 ,
         \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 ,
         \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 ,
         \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 ,
         \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 ,
         \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 ,
         \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 ,
         \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 ,
         \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 ,
         \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 ,
         \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 ,
         \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 ,
         \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 ,
         \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 ,
         \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 ,
         \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 ,
         \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 ,
         \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 ,
         \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 ,
         \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 ,
         \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 ,
         \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 ,
         \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 ,
         \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 ,
         \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 ,
         \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 ,
         \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 ,
         \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 ,
         \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 ,
         \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 ,
         \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 ,
         \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 ,
         \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 ,
         \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 ,
         \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 ,
         \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 ,
         \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 ,
         \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 ,
         \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 ,
         \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 ,
         \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 ,
         \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 ,
         \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 ,
         \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 ,
         \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 ,
         \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 ,
         \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 ,
         \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 ,
         \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 ,
         \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 ,
         \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 ,
         \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 ,
         \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 ,
         \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 ,
         \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 ,
         \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 ,
         \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 ,
         \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 ,
         \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 ,
         \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 ,
         \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 ,
         \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 ,
         \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 ,
         \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 ,
         \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 ,
         \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 ,
         \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 ,
         \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 ,
         \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 ,
         \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 ,
         \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 ,
         \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 ,
         \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 ,
         \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 ,
         \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 ,
         \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 ,
         \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 ,
         \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 ,
         \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 ,
         \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 ,
         \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 ,
         \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 ,
         \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 ,
         \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 ,
         \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 ,
         \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 ,
         \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 ,
         \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 ,
         \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 ,
         \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 ,
         \7435 , \7436 , \7437 , \7438_N$2 , \7439_N$4 , \7440_N$6 , \7441_N$8 , \7442_N$10 , \7443_N$12 , \7444_N$14 ,
         \7445_N$16 , \7446_N$18 , \7447_N$20 , \7448_N$22 , \7449_N$24 , \7450_N$26 , \7451_N$28 , \7452_N$30 , \7453_N$32 , \7454_N$34 ,
         \7455_N$36 , \7456_N$38 , \7457_N$40 , \7458_N$42 , \7459_N$44 , \7460_N$46 , \7461_N$48 , \7462_N$50 , \7463_N$52 , \7464_N$54 ,
         \7465_N$56 , \7466_N$58 , \7467_N$60 , \7468_N$62 , \7469_N$64 , \7470_N$66 , \7471_N$68 , \7472_N$70 , \7473_N$72 , \7474_N$74 ,
         \7475_N$76 , \7476_N$78 , \7477_N$80 , \7478_N$82 , \7479_N$84 , \7480_N$86 , \7481_N$88 , \7482_N$90 , \7483_N$92 , \7484_N$94 ,
         \7485_N$96 , \7486_N$98 , \7487_N$100 , \7488_N$102 , \7489_N$104 , \7490_N$106 , \7491_N$108 , \7492_N$110 , \7493_N$112 , \7494_N$114 ,
         \7495_N$116 , \7496_N$118 , \7497_N$120 , \7498_N$122 , \7499_N$124 , \7500_N$126 , \7501_N$128 , \7502_N$130 , \7503_N$132 , \7504_N$134 ,
         \7505_N$136 , \7506_N$138 , \7507_N$140 , \7508_N$142 , \7509_N$144 , \7510_N$146 , \7511_N$148 , \7512_N$150 , \7513_N$152 , \7514_N$154 ,
         \7515_N$156 , \7516_N$158 , \7517_N$160 , \7518_N$162 , \7519_N$164 , \7520_N$166 , \7521_N$168 , \7522_N$170 , \7523_N$172 , \7524_N$174 ,
         \7525_N$176 , \7526_N$178 , \7527_N$180 , \7528_N$182 , \7529_N$184 , \7530_N$186 , \7531_N$188 , \7532_N$190 , \7533_N$192 , \7534_N$194 ,
         \7535_N$196 , \7536_N$198 , \7537_N$200 , \7538_N$202 , \7539_N$204 , \7540_N$206 , \7541_N$208 , \7542_N$210 , \7543_N$212 , \7544_N$214 ,
         \7545_N$216 , \7546_N$218 , \7547_N$220 , \7548_N$222 , \7549_N$224 , \7550_N$226 , \7551_N$228 , \7552_N$230 , \7553_N$232 , \7554_N$234 ,
         \7555_N$236 , \7556_N$238 , \7557_N$240 , \7558_N$242 , \7559_N$244 , \7560_N$246 , \7561_N$248 , \7562_N$250 , \7563_N$252 , \7564_N$254 ,
         \7565_N$256 , \7566_N$258 , \7567_N$260 , \7568_N$262 , \7569_N$264 , \7570_N$266 , \7571_N$268 , \7572_N$270 , \7573_N$272 , \7574_N$274 ,
         \7575_N$276 , \7576_N$278 , \7577_N$280 , \7578_N$282 , \7579_N$284 , \7580_N$286 , \7581_N$288 , \7582_N$290 , \7583_N$292 , \7584_N$294 ,
         \7585_N$296 , \7586_N$298 , \7587_N$300 , \7588_N$302 , \7589_N$304 , \7590_N$306 , \7591_N$308 , \7592_N$310 , \7593_N$312 , \7594_N$314 ,
         \7595_N$316 , \7596_N$318 , \7597_N$320 , \7598_N$322 , \7599_N$324 , \7600_N$326 , \7601_N$328 , \7602_N$330 , \7603_N$332 , \7604_N$334 ,
         \7605_N$336 , \7606_N$338 , \7607_N$340 , \7608_N$342 , \7609_N$344 , \7610_N$346 , \7611_N$348 , \7612_N$350 , \7613_N$352 , \7614_N$354 ,
         \7615_N$356 , \7616_N$358 , \7617_N$360 , \7618_N$362 , \7619_N$364 , \7620_N$366 , \7621_N$368 , \7622_N$370 , \7623_N$372 , \7624_N$374 ,
         \7625_N$376 , \7626_N$378 , \7627_N$380 , \7628_N$382 , \7629_N$384 , \7630_N$386 , \7631_N$388 , \7632_N$390 , \7633_N$392 , \7634_N$394 ,
         \7635_N$396 , \7636_N$398 , \7637_N$400 , \7638_N$402 , \7639_N$404 , \7640_N$406 , \7641_N$408 , \7642_N$410 , \7643_N$412 , \7644_N$414 ,
         \7645_N$416 , \7646_N$418 , \7647_N$420 , \7648_N$422 , \7649_N$424 , \7650_N$426 , \7651_N$428 , \7652_N$430 , \7653_N$432 , \7654_N$434 ,
         \7655_N$436 , \7656_N$438 , \7657_N$440 , \7658_N$442 , \7659_N$444 , \7660_N$446 , \7661_N$448 , \7662_N$450 , \7663_N$452 , \7664_N$454 ,
         \7665_N$456 , \7666_N$458 , \7667_N$460 , \7668_N$462 , \7669_N$464 , \7670_N$466 , \7671_N$468 , \7672_N$470 , \7673_N$472 , \7674_N$474 ,
         \7675_N$476 , \7676_N$478 , \7677_N$480 , \7678_N$482 , \7679_N$484 , \7680_N$486 , \7681_N$488 , \7682_N$490 , \7683_N$492 , \7684_N$494 ,
         \7685_N$496 , \7686_N$498 , \7687_N$500 , \7688_N$502 , \7689_N$504 , \7690_N$506 , \7691_N$508 , \7692_N$510 , \7693_N$512 , \7694_N$514 ,
         \7695_N$516 , \7696_N$518 , \7697_N$520 , \7698_N$522 , \7699_N$524 , \7700_N$526 , \7701_N$528 , \7702_N$530 , \7703_N$532 , \7704_N$534 ,
         \7705_N$536 , \7706_N$538 , \7707_N$540 , \7708_N$542 , \7709_N$544 , \7710_N$546 , \7711_N$548 , \7712_N$550 , \7713_N$552 , \7714_N$554 ,
         \7715_N$556 , \7716_N$558 , \7717_N$560 , \7718_N$562 , \7719_N$564 , \7720_N$566 , \7721_N$568 , \7722_N$570 , \7723_N$572 , \7724_N$574 ,
         \7725_N$576 , \7726_N$578 , \7727_N$580 , \7728_N$582 , \7729_N$584 , \7730_N$586 , \7731_N$588 , \7732_N$590 , \7733_N$592 , \7734_N$594 ,
         \7735_N$596 , \7736_N$598 , \7737_N$600 , \7738_N$602 , \7739_N$604 , \7740_N$606 , \7741_N$608 , \7742_N$610 , \7743_N$612 , \7744_N$614 ,
         \7745_N$616 , \7746_N$618 , \7747_N$620 , \7748_N$622 , \7749_N$624 , \7750_N$626 , \7751_N$628 , \7752_N$630 , \7753_N$632 , \7754_N$634 ,
         \7755_N$636 , \7756_N$638 , \7757_N$640 , \7758_N$642 , \7759_N$644 , \7760_N$646 , \7761_N$648 , \7762_N$650 , \7763_N$652 , \7764_N$654 ,
         \7765_N$656 , \7766_N$658 , \7767_N$660 , \7768_N$662 , \7769_N$664 , \7770_N$666 , \7771_N$668 , \7772_N$670 , \7773_N$672 , \7774_N$674 ,
         \7775_N$676 , \7776_N$678 , \7777_N$680 , \7778_N$682 , \7779_N$684 , \7780_N$686 , \7781_N$688 , \7782_N$690 , \7783_N$692 , \7784_N$694 ,
         \7785_N$696 , \7786_N$698 , \7787_N$700 , \7788_N$702 , \7789_N$704 , \7790_N$706 , \7791_N$708 , \7792_N$710 , \7793_N$712 , \7794_N$714 ,
         \7795_N$716 , \7796_N$718 , \7797_N$720 , \7798_N$722 , \7799_N$724 , \7800_N$726 , \7801_N$728 , \7802_N$730 , \7803_N$732 , \7804_N$734 ,
         \7805_N$736 , \7806_N$738 , \7807_N$740 , \7808_N$742 , \7809_N$744 , \7810_N$746 , \7811_N$748 , \7812_N$750 , \7813_N$752 , \7814_N$754 ,
         \7815_N$756 , \7816_N$758 , \7817_N$760 , \7818_N$762 , \7819_N$764 , \7820_N$766 , \7821_N$768 , \7822_N$770 , \7823_N$772 , \7824_N$774 ,
         \7825_N$776 , \7826_N$778 , \7827_N$780 , \7828_N$782 , \7829_N$784 , \7830_N$786 , \7831_N$788 , \7832_N$790 , \7833_N$792 , \7834_N$794 ,
         \7835_N$796 , \7836_N$798 , \7837_N$800 , \7838_N$802 , \7839_N$804 , \7840_N$806 , \7841_N$808 , \7842_N$810 , \7843_N$812 , \7844_N$814 ,
         \7845_N$816 , \7846_N$818 , \7847_N$820 , \7848_N$822 , \7849_N$824 , \7850_N$826 , \7851_N$828 , \7852_N$830 , \7853_N$832 , \7854_N$834 ,
         \7855_N$836 , \7856_N$838 , \7857_N$840 , \7858_N$842 , \7859_N$844 , \7860_N$846 , \7861_N$848 , \7862_N$850 , \7863_N$852 , \7864_N$854 ,
         \7865_N$856 , \7866_N$858 , \7867_N$860 , \7868_N$862 , \7869_N$864 , \7870_N$866 , \7871_N$868 , \7872_N$870 , \7873_N$872 , \7874_N$874 ,
         \7875_N$876 , \7876_N$878 , \7877_N$880 , \7878_N$882 , \7879_N$884 , \7880_N$886 , \7881_N$888 , \7882_N$890 , \7883_N$892 , \7884_N$894 ,
         \7885_N$896 , \7886_N$898 , \7887_N$900 , \7888_N$902 , \7889_N$904 , \7890_N$906 , \7891_N$908 , \7892_N$910 , \7893_N$912 , \7894_N$914 ,
         \7895_N$916 , \7896_N$918 , \7897_N$920 , \7898_N$922 , \7899_N$924 , \7900_N$926 , \7901_N$928 , \7902_N$930 , \7903_N$932 , \7904_N$934 ,
         \7905_N$936 , \7906_N$938 , \7907_N$940 , \7908_N$942 , \7909_N$944 , \7910_N$946 , \7911_N$948 , \7912_N$950 , \7913_N$952 , \7914_N$954 ,
         \7915_N$956 , \7916_N$958 , \7917_N$960 , \7918_N$962 , \7919_N$964 , \7920_N$966 , \7921_N$968 , \7922_N$970 , \7923_N$972 , \7924_N$974 ,
         \7925_N$976 , \7926_N$978 , \7927_N$980 , \7928_N$982 , \7929_N$984 , \7930_N$986 , \7931_N$988 , \7932_N$990 , \7933_N$992 , \7934_N$994 ,
         \7935_N$996 , \7936_N$998 , \7937_N$1000 , \7938_N$1002 , \7939_N$1004 , \7940_N$1006 , \7941_N$1008 , \7942_N$1010 , \7943_N$1012 , \7944_N$1014 ,
         \7945_N$1016 , \7946_N$1018 , \7947_N$1020 , \7948_N$1022 , \7949_N$1024 , \7950_N$1026 , \7951_N$1028 , \7952_N$1030 , \7953_N$1032 , \7954_N$1034 ,
         \7955_N$1036 , \7956_N$1038 , \7957_N$1040 , \7958_N$1042 , \7959_N$1044 , \7960_N$1046 , \7961_N$1048 , \7962_N$1050 , \7963_N$1052 , \7964_N$1054 ,
         \7965_N$1056 , \7966_N$1058 , \7967_N$1060 , \7968_N$1062 , \7969_N$1064 , \7970_N$1066 , \7971_N$1068 , \7972_N$1070 , \7973_N$1072 , \7974_N$1074 ,
         \7975_N$1076 , \7976_N$1078 , \7977_N$1080 , \7978_N$1082 , \7979_N$1084 , \7980_N$1086 , \7981_N$1088 , \7982_N$1090 , \7983_N$1092 , \7984_N$1094 ,
         \7985_N$1096 , \7986_N$1098 , \7987_N$1100 , \7988_N$1102 , \7989_N$1104 , \7990_N$1106 , \7991_N$1108 , \7992_N$1110 , \7993_N$1112 , \7994_N$1114 ,
         \7995_N$1116 , \7996_N$1118 , \7997_N$1120 , \7998_N$1122 , \7999_N$1124 , \8000_N$1126 , \8001_N$1128 , \8002_N$1130 , \8003_N$1132 , \8004_N$1134 ,
         \8005_N$1136 , \8006_N$1138 , \8007_N$1140 , \8008_N$1142 , \8009_N$1144 , \8010_N$1146 , \8011_N$1148 , \8012_N$1150 , \8013_N$1152 , \8014_N$1154 ,
         \8015_N$1156 , \8016_N$1158 , \8017_N$1160 , \8018_N$1162 , \8019_N$1164 , \8020_N$1166 , \8021_N$1168 , \8022_N$1170 , \8023_N$1172 , \8024_N$1174 ,
         \8025_N$1176 , \8026_N$1178 , \8027_N$1180 , \8028_N$1182 , \8029_N$1184 , \8030_N$1186 , \8031_N$1188 , \8032_N$1190 , \8033_N$1192 , \8034_N$1194 ,
         \8035_N$1196 , \8036_N$1198 , \8037_N$1200 , \8038_N$1202 , \8039_N$1204 , \8040_N$1206 , \8041_N$1208 , \8042_N$1210 , \8043_N$1212 , \8044_N$1214 ,
         \8045_N$1216 , \8046_N$1218 , \8047_N$1220 , \8048_N$1222 , \8049_N$1224 , \8050_N$1226 , \8051_N$1228 , \8052_N$1230 , \8053_N$1232 , \8054_N$1234 ,
         \8055_N$1236 , \8056_N$1238 , \8057_N$1240 , \8058_N$1242 , \8059_N$1244 , \8060_N$1246 , \8061_N$1248 , \8062_N$1250 , \8063_N$1252 , \8064_N$1254 ,
         \8065_N$1256 , \8066_N$1258 , \8067_N$1260 , \8068_N$1262 , \8069_N$1264 , \8070_N$1266 , \8071_N$1268 , \8072_N$1270 , \8073_N$1272 , \8074_N$1274 ,
         \8075_N$1276 , \8076_N$1278 , \8077_N$1280 , \8078_N$1282 , \8079_N$1284 , \8080_N$1286 , \8081_N$1288 , \8082_N$1290 , \8083_N$1292 , \8084_N$1294 ,
         \8085_N$1296 , \8086_N$1298 , \8087_N$1300 , \8088_N$1302 , \8089_N$1304 , \8090_N$1306 , \8091_N$1308 , \8092_N$1310 , \8093_N$1312 , \8094_N$1314 ,
         \8095_N$1316 , \8096_N$1318 , \8097_N$1320 , \8098_N$1322 , \8099_N$1324 , \8100_N$1326 , \8101_N$1328 , \8102_N$1330 , \8103_N$1332 , \8104_N$1334 ,
         \8105_N$1336 , \8106_N$1338 , \8107_N$1340 , \8108_N$1342 , \8109_N$1344 , \8110_N$1346 , \8111_N$1348 , \8112_N$1350 , \8113_N$1352 , \8114_N$1354 ,
         \8115_N$1356 , \8116_N$1358 , \8117_N$1360 , \8118_N$1362 , \8119_N$1364 , \8120_N$1366 , \8121_N$1368 , \8122_N$1370 , \8123_N$1372 , \8124_N$1374 ,
         \8125_N$1376 , \8126_N$1378 , \8127_N$1380 , \8128_N$1382 , \8129_N$1384 , \8130_N$1386 , \8131_N$1388 , \8132_N$1390 , \8133_N$1392 , \8134_N$1394 ,
         \8135_N$1396 , \8136_N$1398 , \8137_N$1400 , \8138_N$1402 , \8139_N$1404 , \8140_N$1406 , \8141_N$1408 , \8142_N$1410 , \8143_N$1412 , \8144_N$1414 ,
         \8145_N$1416 , \8146_N$1418 , \8147_N$1420 , \8148_N$1422 , \8149_N$1424 , \8150_N$1426 , \8151_N$1428 , \8152_N$1430 , \8153_N$1432 , \8154_N$1434 ,
         \8155_N$1436 , \8156_N$1438 , \8157_N$1440 , \8158_N$1442 , \8159_N$1444 , \8160_N$1446 , \8161_N$1448 , \8162_N$1450 , \8163_N$1452 , \8164_N$1454 ,
         \8165_N$1456 , \8166_N$1458 , \8167_N$1460 , \8168_N$1462 , \8169_N$1464 , \8170_N$1466 , \8171_N$1468 , \8172_N$1470 , \8173_N$1472 , \8174_N$1474 ,
         \8175_N$1476 , \8176_N$1478 , \8177_N$1480 , \8178_N$1482 , \8179_N$1484 , \8180_N$1486 , \8181_N$1488 , \8182_N$1490 , \8183_N$1492 , \8184_N$1494 ,
         \8185_N$1496 , \8186_N$1498 , \8187_N$1500 , \8188_N$1502 , \8189_N$1504 , \8190_N$1506 , \8191_N$1508 , \8192_N$1510 , \8193_N$1512 , \8194_N$1514 ,
         \8195_N$1516 , \8196_N$1518 , \8197_N$1520 , \8198_N$1522 , \8199_N$1524 , \8200_N$1526 , \8201_N$1528 , \8202_N$1530 , \8203_N$1532 , \8204_N$1534 ,
         \8205_N$1536 , \8206_N$1538 , \8207_N$1540 , \8208_N$1542 , \8209_N$1544 , \8210_N$1546 , \8211_N$1548 , \8212_N$1550 , \8213_N$1552 , \8214_N$1554 ,
         \8215_N$1556 , \8216_N$1558 , \8217_N$1560 , \8218_N$1562 , \8219_N$1564 , \8220_N$1566 , \8221_N$1568 , \8222_N$1570 , \8223_N$1572 , \8224_N$1574 ,
         \8225_N$1576 , \8226_N$1578 , \8227_N$1580 , \8228_N$1582 , \8229_N$1584 , \8230_N$1586 , \8231_N$1588 , \8232_N$1590 , \8233_N$1592 , \8234_N$1594 ,
         \8235_N$1596 , \8236_N$1598 , \8237_N$1600 , \8238_N$1602 , \8239_N$1604 , \8240_N$1606 , \8241_N$1608 , \8242_N$1610 , \8243_N$1612 , \8244_N$1614 ,
         \8245_N$1616 , \8246_N$1618 , \8247_N$1620 , \8248_N$1622 , \8249_N$1624 , \8250_N$1626 , \8251_N$1628 , \8252_N$1630 , \8253_N$1632 , \8254_N$1634 ,
         \8255_N$1636 , \8256_N$1638 , \8257_N$1640 , \8258_N$1642 , \8259_N$1644 , \8260_N$1646 , \8261_N$1648 , \8262_N$1650 , \8263_N$1652 , \8264_N$1654 ,
         \8265_N$1656 , \8266_N$1658 , \8267_N$1660 , \8268_N$1662 , \8269_N$1664 , \8270_N$1666 , \8271_N$1668 , \8272_N$1670 , \8273_N$1672 , \8274_N$1674 ,
         \8275_N$1676 , \8276_N$1678 , \8277_N$1680 , \8278_N$1682 , \8279_N$1684 , \8280_N$1686 , \8281_N$1688 , \8282_N$1690 , \8283_N$1692 , \8284_N$1694 ,
         \8285_N$1696 , \8286_N$1698 , \8287_N$1700 , \8288_N$1702 , \8289_N$1704 , \8290_N$1706 , \8291_N$1708 , \8292_N$1710 , \8293_N$1712 , \8294_N$1714 ,
         \8295_N$1716 , \8296_N$1718 , \8297_N$1720 , \8298_N$1722 , \8299_N$1724 , \8300_N$1726 , \8301_N$1728 , \8302_N$1730 , \8303_N$1732 , \8304_N$1734 ,
         \8305_N$1736 , \8306_N$1738 , \8307_N$1740 , \8308_N$1742 , \8309_N$1744 , \8310_N$1746 , \8311_N$1748 , \8312_N$1750 , \8313_N$1752 , \8314_N$1754 ,
         \8315_N$1756 , \8316_N$1758 , \8317_N$1760 , \8318_N$1762 , \8319_N$1764 , \8320_N$1766 , \8321_N$1768 , \8322_N$1770 , \8323_N$1772 , \8324_N$1774 ,
         \8325_N$1776 , \8326_N$1778 , \8327_N$1780 , \8328_N$1782 , \8329_N$1784 , \8330_N$1786 , \8331_N$1788 , \8332_N$1790 , \8333_N$1792 , \8334_N$1794 ,
         \8335_N$1796 , \8336_N$1798 , \8337_N$1800 , \8338_N$1802 , \8339_N$1804 , \8340_N$1806 , \8341_N$1808 , \8342_N$1810 , \8343_N$1812 , \8344_N$1814 ,
         \8345_N$1816 , \8346_N$1818 , \8347_N$1820 , \8348_N$1822 , \8349_N$1824 , \8350_N$1826 , \8351_N$1828 , \8352_N$1830 , \8353_N$1832 , \8354_N$1834 ,
         \8355_N$1836 , \8356_N$1838 , \8357_N$1840 , \8358_N$1842 , \8359_N$1844 , \8360_N$1846 , \8361_N$1848 , \8362_N$1850 , \8363_N$1852 , \8364_N$1854 ,
         \8365_N$1856 , \8366_N$1858 , \8367_N$1860 , \8368_N$1862 , \8369_N$1864 , \8370_N$1866 , \8371_N$1868 , \8372_N$1870 , \8373_N$1872 , \8374_N$1874 ,
         \8375_N$1876 , \8376_N$1878 , \8377_N$1880 , \8378_N$1882 , \8379_N$1884 , \8380_N$1886 , \8381_N$1888 , \8382_N$1890 , \8383_N$1892 , \8384_N$1894 ,
         \8385_N$1896 , \8386_N$1898 , \8387_N$1900 , \8388_N$1902 , \8389_N$1904 , \8390_N$1906 , \8391_N$1908 , \8392_N$1910 , \8393_N$1912 , \8394_N$1914 ,
         \8395_N$1916 , \8396_N$1918 , \8397_N$1920 , \8398_N$1922 , \8399_N$1924 , \8400_N$1926 , \8401_N$1928 , \8402_N$1930 , \8403_N$1932 , \8404_N$1934 ,
         \8405_N$1936 , \8406_N$1938 , \8407_N$1940 , \8408_N$1942 , \8409_N$1944 , \8410_N$1946 , \8411_N$1948 , \8412_N$1950 , \8413_N$1952 , \8414_N$1954 ,
         \8415_N$1956 , \8416_N$1958 , \8417_N$1960 , \8418_N$1962 , \8419_N$1964 , \8420_N$1966 , \8421_N$1968 , \8422_N$1970 , \8423_N$1972 , \8424_N$1974 ,
         \8425_N$1976 , \8426_N$1978 , \8427_N$1980 , \8428_N$1982 , \8429_N$1984 , \8430_N$1986 , \8431_N$1988 , \8432_N$1990 , \8433_N$1992 , \8434_N$1994 ,
         \8435_N$1996 , \8436_N$1998 , \8437_N$2000 , \8438_N$2002 , \8439_N$2004 , \8440_N$2006 , \8441_N$2008 , \8442_N$2010 , \8443_N$2012 , \8444_N$2014 ,
         \8445_N$2016 , \8446_N$2018 , \8447_N$2020 , \8448_N$2022 , \8449_N$2024 , \8450_N$2026 , \8451_N$2028 , \8452_N$2030 , \8453_N$2032 , \8454_N$2034 ,
         \8455_N$2036 , \8456_N$2038 , \8457_N$2040 , \8458_N$2042 , \8459_N$2044 , \8460_N$2046 , \8461_N$2048 , \8462_N$2050 , \8463_N$2052 , \8464_N$2054 ,
         \8465_N$2056 , \8466_N$2058 , \8467_N$2060 , \8468_N$2062 , \8469_N$2064 , \8470_N$2066 , \8471_N$2068 , \8472_N$2070 , \8473_N$2072 , \8474_N$2074 ,
         \8475_N$2076 , \8476_N$2078 , \8477_N$2080 , \8478_N$2082 , \8479_N$2084 , \8480_N$2086 , \8481_N$2088 , \8482_N$2090 , \8483_N$2092 , \8484_N$2094 ,
         \8485_N$2096 , \8486_N$2098 , \8487_N$2100 , \8488_N$2102 , \8489_N$2104 , \8490_N$2106 , \8491_N$2108 , \8492_N$2110 , \8493_N$2112 , \8494_N$2114 ,
         \8495_N$2116 , \8496_N$2118 , \8497_N$2120 , \8498_N$2122 , \8499_N$2124 , \8500_N$2126 , \8501_N$2128 , \8502_N$2130 , \8503_N$2132 , \8504_N$2134 ,
         \8505_N$2136 , \8506_N$2138 , \8507_N$2140 , \8508_N$2142 , \8509_N$2144 , \8510_N$2146 , \8511_N$2148 , \8512_N$2150 , \8513_N$2152 , \8514_N$2154 ,
         \8515_N$2156 , \8516_N$2158 , \8517_N$2160 , \8518_N$2162 , \8519_N$2164 , \8520_N$2166 , \8521_N$2168 , \8522_N$2170 , \8523_N$2172 , \8524_N$2174 ,
         \8525_N$2176 , \8526_N$2178 , \8527_N$2180 , \8528_N$2182 , \8529_N$2184 , \8530_N$2186 , \8531_N$2188 , \8532_N$2190 , \8533_N$2192 , \8534_N$2194 ,
         \8535_N$2196 , \8536_N$2198 , \8537_N$2200 , \8538_N$2202 , \8539_N$2204 , \8540_N$2206 , \8541_N$2208 , \8542_N$2210 , \8543_N$2212 , \8544_N$2214 ,
         \8545_N$2216 , \8546_N$2218 , \8547_N$2220 , \8548_N$2222 , \8549_N$2224 , \8550_N$2226 , \8551_N$2228 , \8552_N$2230 , \8553_N$2232 , \8554_N$2234 ,
         \8555_N$2236 , \8556_N$2238 , \8557_N$2240 , \8558_N$2242 , \8559_N$2244 , \8560_N$2246 , \8561_N$2248 , \8562_N$2250 , \8563_N$2252 , \8564_N$2254 ,
         \8565_N$2256 , \8566_N$2258 , \8567_N$2260 , \8568_N$2262 , \8569_N$2264 , \8570_N$2266 , \8571_N$2268 , \8572_N$2270 , \8573_N$2272 , \8574_N$2274 ,
         \8575_N$2276 , \8576_N$2278 , \8577_N$2280 , \8578_N$2282 , \8579_N$2284 , \8580_N$2286 , \8581_N$2288 , \8582_N$2290 , \8583_N$2292 , \8584_N$2294 ,
         \8585_N$2296 , \8586_N$2298 , \8587_N$2300 , \8588_N$2302 , \8589_N$2304 , \8590_N$2306 , \8591_N$2308 , \8592_N$2310 , \8593_N$2312 , \8594_N$2314 ,
         \8595_N$2316 , \8596_N$2318 , \8597_N$2320 , \8598_N$2322 , \8599_N$2324 , \8600_N$2326 , \8601_N$2328 , \8602_N$2330 , \8603_N$2332 , \8604_N$2334 ,
         \8605_N$2336 , \8606_N$2338 , \8607_N$2340 , \8608_N$2342 , \8609_N$2344 , \8610_N$2346 , \8611_N$2348 , \8612_N$2350 , \8613_N$2352 , \8614_N$2354 ,
         \8615_N$2356 , \8616_N$2358 , \8617_N$2360 , \8618_N$2362 , \8619_N$2364 , \8620_N$2366 , \8621_N$2368 , \8622_N$2370 , \8623_N$2372 , \8624_N$2374 ,
         \8625_N$2376 , \8626_N$2378 , \8627_N$2380 , \8628_N$2382 , \8629_N$2384 , \8630_N$2386 , \8631_N$2388 , \8632_N$2390 , \8633_N$2392 , \8634_N$2394 ,
         \8635_N$2396 , \8636_N$2398 , \8637_N$2400 , \8638_N$2402 , \8639_N$2404 , \8640_N$2406 , \8641_N$2408 , \8642_N$2410 , \8643_N$2412 , \8644_N$2414 ,
         \8645_N$2416 , \8646_N$2418 , \8647_N$2420 , \8648_N$2422 , \8649_N$2424 , \8650_N$2426 , \8651_N$2428 , \8652_N$2430 , \8653_N$2432 , \8654_N$2434 ,
         \8655_N$2436 , \8656_N$2438 , \8657_N$2440 , \8658_N$2442 , \8659_N$2444 , \8660_N$2446 , \8661_N$2448 , \8662_N$2450 , \8663_N$2452 , \8664_N$2454 ,
         \8665_N$2456 , \8666_N$2458 , \8667_N$2460 , \8668_N$2462 , \8669_N$2464 , \8670_N$2466 , \8671_N$2468 , \8672_N$2470 , \8673_N$2472 , \8674_N$2474 ,
         \8675_N$2476 , \8676_N$2478 , \8677_N$2480 , \8678_N$2482 , \8679_N$2484 , \8680_N$2486 , \8681_N$2488 , \8682_N$2490 , \8683_N$2492 , \8684_N$2494 ,
         \8685_N$2496 , \8686_N$2498 , \8687_N$2500 , \8688_N$2502 , \8689_N$2504 , \8690_N$2506 , \8691_N$2508 , \8692_N$2510 , \8693_N$2512 , \8694_N$2514 ,
         \8695_N$2516 , \8696_N$2518 , \8697_N$2520 , \8698_N$2522 , \8699_N$2524 , \8700_N$2526 , \8701_N$2528 , \8702_N$2530 , \8703_N$2532 , \8704_N$2534 ,
         \8705_N$2536 , \8706_N$2538 , \8707_N$2540 , \8708_N$2542 , \8709_N$2544 , \8710_N$2546 , \8711_N$2548 , \8712_N$2550 , \8713_N$2552 , \8714_N$2554 ,
         \8715_N$2556 , \8716_N$2558 , \8717_N$2560 , \8718_N$2562 , \8719_N$2564 , \8720_N$2566 , \8721_N$2568 , \8722_N$2570 , \8723_N$2572 , \8724_N$2574 ,
         \8725_N$2576 , \8726_N$2578 , \8727_N$2580 , \8728_N$2582 , \8729_N$2584 , \8730_N$2586 , \8731_N$2588 , \8732_N$2590 , \8733_N$2592 , \8734_N$2594 ,
         \8735_N$2596 , \8736_N$2598 , \8737_N$2600 , \8738_N$2602 , \8739_N$2604 , \8740_N$2606 , \8741_N$2608 , \8742_N$2610 , \8743_N$2612 , \8744_N$2614 ,
         \8745_N$2616 , \8746_N$2618 , \8747_N$2620 , \8748_N$2622 , \8749_N$2624 , \8750_N$2626 , \8751_N$2628 , \8752_N$2630 , \8753_N$2632 , \8754_N$2634 ,
         \8755_N$2636 , \8756_N$2638 , \8757_N$2640 , \8758_N$2642 , \8759_N$2644 , \8760_N$2646 , \8761_N$2648 , \8762_N$2650 , \8763_N$2652 , \8764_N$2654 ,
         \8765_N$2656 , \8766_N$2658 , \8767_N$2660 , \8768_N$2662 , \8769_N$2664 , \8770_N$2666 , \8771_N$2668 , \8772_N$2670 , \8773_N$2672 , \8774_N$2674 ,
         \8775_N$2676 , \8776_N$2678 , \8777_N$2680 , \8778_N$2682 , \8779_N$2684 , \8780_N$2686 , \8781_N$2688 , \8782_N$2690 , \8783_N$2692 , \8784_N$2694 ,
         \8785_N$2696 , \8786_N$2698 , \8787_N$2700 , \8788_N$2702 , \8789_N$2704 , \8790_N$2706 , \8791_N$2708 , \8792_N$2710 , \8793_N$2712 , \8794_N$2714 ,
         \8795_N$2716 , \8796_N$2718 , \8797_N$2720 , \8798_N$2722 , \8799_N$2724 , \8800_N$2726 , \8801_N$2728 , \8802_N$2730 , \8803_N$2732 , \8804_N$2734 ,
         \8805_N$2736 , \8806_N$2738 , \8807_N$2740 , \8808_N$2742 , \8809_N$2744 , \8810_N$2746 , \8811_N$2748 , \8812_N$2750 , \8813_N$2752 , \8814_N$2754 ,
         \8815_N$2756 , \8816_N$2758 , \8817_N$2760 , \8818_N$2763 , \8819_ONE , \8820 , \8821 , \8822 , \8823 , \8824 ,
         \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 ,
         \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 ,
         \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 ,
         \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 ,
         \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 ,
         \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 ,
         \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 ,
         \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 ,
         \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 ,
         \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 ,
         \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 ,
         \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 ,
         \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 ,
         \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 ,
         \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 ,
         \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 ,
         \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 ,
         \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 ,
         \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 ,
         \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 ,
         \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 ,
         \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 ,
         \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 ,
         \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 ,
         \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 ,
         \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 ,
         \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 ,
         \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 ,
         \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 ,
         \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 ,
         \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 ,
         \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 ,
         \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 ,
         \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 ,
         \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 ,
         \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 ,
         \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 ,
         \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 ,
         \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 ,
         \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 ,
         \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 ,
         \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 ,
         \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 ,
         \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 ,
         \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 ,
         \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 ,
         \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 ,
         \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 ,
         \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 ,
         \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 ,
         \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 ,
         \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 ,
         \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 ,
         \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 ,
         \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 ,
         \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 ,
         \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 ,
         \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 ,
         \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 ,
         \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 ,
         \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 ,
         \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 ,
         \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 ,
         \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 ,
         \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 ,
         \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 ,
         \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 ,
         \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 ,
         \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 ,
         \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 ,
         \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 ,
         \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 ,
         \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 ,
         \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 ,
         \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 ,
         \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 ,
         \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 ,
         \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 ,
         \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 ,
         \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 ,
         \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 ,
         \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 ,
         \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 ,
         \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 ,
         \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 ,
         \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 ,
         \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 ,
         \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 ,
         \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 ,
         \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 ,
         \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 ,
         \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 ,
         \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 ,
         \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 ,
         \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 ,
         \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 ,
         \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 ,
         \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 ,
         \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 ,
         \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 ,
         \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 ,
         \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 ,
         \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 ,
         \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 ,
         \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 ,
         \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 ,
         \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 ,
         \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 ,
         \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 ,
         \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 ,
         \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 ,
         \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 ,
         \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 ,
         \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 ,
         \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 ,
         \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 ,
         \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 ,
         \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 ,
         \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 ,
         \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 ,
         \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 ,
         \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 ,
         \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 ,
         \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 ,
         \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 ,
         \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 ,
         \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 ,
         \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 ,
         \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 ,
         \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 ,
         \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 ,
         \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 ,
         \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 ,
         \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 ,
         \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 ,
         \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 ,
         \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 ,
         \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 ,
         \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 ,
         \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 ,
         \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 ,
         \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 ,
         \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 ,
         \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 ,
         \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 ,
         \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 ,
         \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 ,
         \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 ,
         \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 ,
         \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 ,
         \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 ,
         \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 ,
         \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 ,
         \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 ,
         \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 ,
         \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 ,
         \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 ,
         \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 ,
         \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 ,
         \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 ,
         \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 ,
         \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 ,
         \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 ,
         \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 ,
         \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 ,
         \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 ,
         \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 ,
         \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 ,
         \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 ,
         \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 ,
         \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 ,
         \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 ,
         \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 ,
         \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 ,
         \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 ,
         \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 ,
         \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 ,
         \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 ,
         \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 ,
         \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 ,
         \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 ,
         \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 ,
         \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 ,
         \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 ,
         \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 ,
         \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 ,
         \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 ,
         \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 ,
         \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 ,
         \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 ,
         \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 ,
         \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 ,
         \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 ,
         \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 ,
         \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 ,
         \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 ,
         \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 ,
         \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 ,
         \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 ,
         \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 ,
         \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 ,
         \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 ,
         \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 ,
         \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 ,
         \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 ,
         \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 ,
         \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 ,
         \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 ,
         \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 ,
         \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 ,
         \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 ,
         \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 ,
         \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 ,
         \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 ,
         \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 ,
         \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 ,
         \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 ,
         \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 ,
         \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 ,
         \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 ,
         \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 ,
         \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 ,
         \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 ,
         \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 ,
         \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 ,
         \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 ,
         \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 ,
         \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 ,
         \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 ,
         \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 ,
         \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 ,
         \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 ,
         \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 ,
         \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 ,
         \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 ,
         \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 ,
         \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 ,
         \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 ,
         \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 ,
         \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 ,
         \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 ,
         \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 ,
         \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 ,
         \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 ,
         \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 ,
         \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 ,
         \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 ,
         \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 ,
         \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 ,
         \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 ,
         \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 ,
         \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 ,
         \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 ,
         \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 ,
         \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 ,
         \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 ,
         \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 ,
         \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 ,
         \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 ,
         \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 ,
         \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 ,
         \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 ,
         \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 ,
         \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 ,
         \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 ,
         \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 ,
         \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 ,
         \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 ,
         \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 ,
         \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 ,
         \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 ,
         \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 ,
         \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 ,
         \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 ,
         \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 ,
         \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 ,
         \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 ,
         \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 ,
         \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 ,
         \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 ,
         \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 ,
         \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 ,
         \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 ,
         \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 ,
         \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 ,
         \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 ,
         \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 ,
         \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 ,
         \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 ,
         \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 ,
         \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 ,
         \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 ,
         \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 ,
         \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 ,
         \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 ,
         \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 ,
         \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 ,
         \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 ,
         \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 ,
         \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 ,
         \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 ,
         \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 ,
         \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 ,
         \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 ,
         \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 ,
         \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 ,
         \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 ,
         \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 ,
         \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 ,
         \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 ,
         \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 ,
         \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 ,
         \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 ,
         \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 ,
         \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 ,
         \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 ,
         \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 ,
         \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 ,
         \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 ,
         \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 ,
         \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 ,
         \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 ,
         \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 ,
         \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 ,
         \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 ,
         \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 ,
         \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 ,
         \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 ,
         \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 ,
         \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 ,
         \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 ,
         \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 ,
         \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 ,
         \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 ,
         \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 ,
         \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 ,
         \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 ,
         \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 ,
         \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 ,
         \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 ,
         \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 ,
         \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 ,
         \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 ,
         \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 ,
         \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 ,
         \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 ,
         \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 ,
         \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 ,
         \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 ,
         \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 ,
         \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 ,
         \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 ,
         \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 ,
         \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 ,
         \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 ,
         \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 ,
         \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 ,
         \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 ,
         \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 ,
         \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 ,
         \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 ,
         \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 ,
         \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 ,
         \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 ,
         \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 ,
         \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 ,
         \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 ,
         \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 ,
         \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 ,
         \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 ,
         \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 ,
         \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 ,
         \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 ,
         \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 ,
         \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 ,
         \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 ,
         \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 ,
         \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 ,
         \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 ,
         \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 ,
         \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 ,
         \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 ,
         \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 ,
         \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 ,
         \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 ,
         \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 ,
         \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 ,
         \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 ,
         \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 ,
         \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 ,
         \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 ,
         \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 ,
         \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 ,
         \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 ,
         \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 ,
         \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 ,
         \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 ,
         \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 ,
         \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 ,
         \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 ,
         \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 ,
         \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 ,
         \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 ,
         \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 ,
         \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 ,
         \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 ,
         \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 ,
         \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 ,
         \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 ,
         \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 ,
         \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 ,
         \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 ,
         \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 ,
         \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 ,
         \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 ,
         \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 ,
         \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 ,
         \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 ,
         \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 ,
         \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 ,
         \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 ,
         \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 ,
         \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 ,
         \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 ,
         \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 ,
         \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 ,
         \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 ,
         \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 ,
         \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 ,
         \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 ,
         \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 ,
         \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 ,
         \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 ,
         \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 ,
         \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 ,
         \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 ,
         \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 ,
         \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 ,
         \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 ,
         \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 ,
         \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 ,
         \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 ,
         \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 ,
         \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 ,
         \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 ,
         \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 ,
         \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 ,
         \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 ,
         \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 ,
         \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 ,
         \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 ,
         \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 ,
         \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 ,
         \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 ,
         \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 ,
         \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 ,
         \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 ,
         \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 ,
         \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 ,
         \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 ,
         \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 ,
         \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 ,
         \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 ,
         \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 ,
         \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 ,
         \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 ,
         \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 ,
         \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 ,
         \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 ,
         \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 ,
         \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 ,
         \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 ,
         \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 ,
         \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 ,
         \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 ,
         \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 ,
         \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 ,
         \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 ,
         \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 ,
         \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 ,
         \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 ,
         \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 ,
         \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 ,
         \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 ,
         \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 ,
         \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 ,
         \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 ,
         \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 ,
         \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 ,
         \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 ,
         \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 ,
         \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 ,
         \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 ,
         \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 ,
         \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 ,
         \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 ,
         \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 ,
         \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 ,
         \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 ,
         \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 ,
         \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 ,
         \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 ,
         \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 ,
         \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 ,
         \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 ,
         \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 ,
         \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 ,
         \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 ,
         \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 ,
         \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 ,
         \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 ,
         \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 ,
         \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 ,
         \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 ,
         \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 ,
         \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 ,
         \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 ,
         \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 ,
         \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 ,
         \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 ,
         \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 ,
         \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 ,
         \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 ,
         \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 ,
         \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 ,
         \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 ,
         \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 ,
         \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 ,
         \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 ,
         \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 ,
         \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 ,
         \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 ,
         \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 ,
         \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 ,
         \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 ,
         \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 ,
         \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 ,
         \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 ,
         \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 ,
         \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 ,
         \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 ,
         \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 ,
         \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 ,
         \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 ,
         \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 ,
         \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 ,
         \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 ,
         \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 ,
         \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 ,
         \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 ,
         \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 ,
         \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 ,
         \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 ,
         \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 ,
         \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 ,
         \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 ,
         \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 ,
         \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 ,
         \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 ,
         \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 ,
         \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 ,
         \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 ,
         \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 ,
         \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 ,
         \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 ,
         \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 ,
         \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 ,
         \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 ,
         \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 ,
         \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 ,
         \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 ,
         \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 ,
         \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 ,
         \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 ,
         \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 ,
         \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 ,
         \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 ,
         \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 ,
         \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 ,
         \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 ,
         \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 ,
         \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 ,
         \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 ,
         \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 ,
         \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 ,
         \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 ,
         \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 ,
         \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 ,
         \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 ,
         \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 ,
         \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 ,
         \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 ,
         \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 ,
         \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 ,
         \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 ,
         \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 ,
         \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 ,
         \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 ,
         \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 ,
         \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 ,
         \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 ,
         \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 ,
         \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 ,
         \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 ,
         \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 ,
         \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 ,
         \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 ,
         \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 ,
         \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 ,
         \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 ,
         \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 ,
         \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 ,
         \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 ,
         \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 ,
         \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 ,
         \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 ,
         \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 ,
         \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 ,
         \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 ,
         \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 ,
         \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 ,
         \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 ,
         \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 ,
         \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 ,
         \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 ,
         \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 ,
         \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 ,
         \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 ,
         \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 ,
         \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 ,
         \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 ,
         \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 ,
         \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 ,
         \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 ,
         \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 ,
         \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 ,
         \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 ,
         \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 ,
         \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 ,
         \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 ,
         \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 ,
         \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 ,
         \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 ,
         \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 ,
         \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 ,
         \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 ,
         \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 ,
         \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 ,
         \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 ,
         \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 ,
         \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 ,
         \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 ,
         \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 ,
         \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 ,
         \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 ,
         \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 ,
         \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 ,
         \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 ,
         \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 ,
         \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 ,
         \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 ,
         \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 ,
         \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 ,
         \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 ,
         \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 ,
         \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 ,
         \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 ,
         \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 ,
         \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 ,
         \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 ,
         \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 ,
         \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 ,
         \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 ,
         \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 ,
         \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 ,
         \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 ,
         \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 ,
         \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 ,
         \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 ,
         \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 ,
         \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 ,
         \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 ,
         \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 ,
         \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 ,
         \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 ,
         \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 ,
         \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 ,
         \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 ,
         \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 ,
         \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 ,
         \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 ,
         \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 ,
         \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 ,
         \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 ,
         \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 ,
         \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 ,
         \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 ,
         \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 ,
         \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 ,
         \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 ,
         \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 ,
         \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 ,
         \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 ,
         \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 ,
         \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 ,
         \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 ,
         \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 ,
         \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 ,
         \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 ,
         \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 ,
         \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 ,
         \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 ,
         \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 ,
         \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 ,
         \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 ,
         \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 ,
         \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 ,
         \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 ,
         \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 ,
         \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 ,
         \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 ,
         \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 ,
         \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 ,
         \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 ,
         \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 ,
         \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 ,
         \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 ,
         \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 ,
         \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 ,
         \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 ,
         \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 ,
         \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 ,
         \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 ,
         \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 ,
         \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 ,
         \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 ,
         \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 ,
         \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 ,
         \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 ,
         \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 ,
         \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 ,
         \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 ,
         \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 ,
         \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 ,
         \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 ,
         \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 ,
         \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 ,
         \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 ,
         \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 ,
         \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 ,
         \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 ,
         \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 ,
         \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 ,
         \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 ,
         \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 ,
         \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 ,
         \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 ,
         \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 ,
         \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 ,
         \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 ,
         \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 ,
         \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 ,
         \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 ,
         \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 ,
         \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 ,
         \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 ,
         \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 ,
         \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 ,
         \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 ,
         \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 ,
         \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 ,
         \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 ,
         \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 ,
         \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 ,
         \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 ,
         \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 ,
         \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 ,
         \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 ,
         \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 ,
         \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 ,
         \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 ,
         \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 ,
         \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 ,
         \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 ,
         \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 ,
         \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 ,
         \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 ,
         \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 ,
         \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 ,
         \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 ,
         \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 ,
         \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 ,
         \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 ,
         \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 ,
         \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 ,
         \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 ,
         \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 ,
         \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 ,
         \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 ,
         \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 ,
         \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 ,
         \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 ,
         \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 ,
         \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 ,
         \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 ,
         \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 ,
         \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 ,
         \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 ,
         \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 ,
         \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 ,
         \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 ,
         \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 ,
         \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 ,
         \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 ,
         \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 ,
         \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 ,
         \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 ,
         \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 ,
         \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 ,
         \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 ,
         \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 ,
         \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 ,
         \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 ,
         \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 ,
         \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 ,
         \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 ,
         \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 ,
         \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 ,
         \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 ,
         \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 ,
         \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 ,
         \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 ,
         \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 ,
         \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 ,
         \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 ,
         \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 ,
         \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 ,
         \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 ,
         \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 ,
         \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 ,
         \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 ,
         \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 ,
         \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 ,
         \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 ,
         \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 ,
         \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 ,
         \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 ,
         \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 ,
         \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 ,
         \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 ,
         \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 ,
         \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 ,
         \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 ,
         \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 ,
         \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 ,
         \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 ,
         \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 ,
         \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 ,
         \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 ,
         \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 ,
         \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 ,
         \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 ,
         \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 ,
         \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 ,
         \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 ,
         \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 ,
         \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 ,
         \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 ,
         \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 ,
         \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 ,
         \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 ,
         \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 ,
         \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 ,
         \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 ,
         \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 ,
         \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 ,
         \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 ,
         \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 ,
         \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 ,
         \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 ,
         \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 ,
         \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 ,
         \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 ,
         \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 ,
         \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 ,
         \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 ,
         \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 ,
         \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 ,
         \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 ,
         \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 ,
         \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 ,
         \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 ,
         \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 ,
         \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 ,
         \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 ,
         \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 ,
         \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 ,
         \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 ,
         \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 ,
         \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 ,
         \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 ,
         \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 ,
         \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 ,
         \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 ,
         \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 ,
         \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 ,
         \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 ,
         \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 ,
         \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 ,
         \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 ,
         \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 ,
         \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 ,
         \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 ,
         \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 ,
         \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 ,
         \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 ,
         \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 ,
         \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 ,
         \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 ,
         \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 ,
         \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 , \18033 , \18034 ,
         \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 ,
         \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 ,
         \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 ,
         \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 ,
         \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 ,
         \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 ,
         \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 ,
         \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 ,
         \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 ,
         \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 ,
         \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 ,
         \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 ,
         \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 ,
         \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 ,
         \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 ,
         \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 ,
         \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 ,
         \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 ,
         \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 ,
         \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 ,
         \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 ,
         \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 ,
         \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 ,
         \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 ,
         \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 ,
         \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 ,
         \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 ,
         \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 ,
         \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 ,
         \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 ,
         \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 ,
         \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 ,
         \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 ,
         \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 ,
         \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 ,
         \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 ,
         \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 ,
         \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 ,
         \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 ,
         \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 ,
         \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 ,
         \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 ,
         \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 ,
         \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 ,
         \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 ,
         \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 ,
         \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 ,
         \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 ,
         \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 ,
         \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 ,
         \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 ,
         \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 ,
         \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 ,
         \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 ,
         \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 ,
         \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 ,
         \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 ,
         \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 ,
         \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 ,
         \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 ,
         \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 ,
         \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 ,
         \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 ,
         \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 ,
         \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 ,
         \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 ,
         \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 ,
         \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 ,
         \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 ,
         \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 ,
         \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 ,
         \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 ,
         \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 ,
         \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 ,
         \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 ,
         \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 ,
         \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 ,
         \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 ,
         \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 ,
         \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 ,
         \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 ,
         \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 ,
         \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 ,
         \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 ,
         \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 ,
         \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 ,
         \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 ,
         \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 ,
         \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 ,
         \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 ,
         \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 ,
         \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 ,
         \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 ,
         \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 ,
         \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 ,
         \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 ,
         \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 ,
         \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 ,
         \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 ,
         \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 ,
         \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 ,
         \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 ,
         \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 ,
         \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 ,
         \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 ,
         \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 , \19093 , \19094 ,
         \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 ,
         \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 ,
         \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 ,
         \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 ,
         \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 ,
         \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 ,
         \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 ,
         \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 ,
         \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 ,
         \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 ,
         \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 ,
         \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 ,
         \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 ,
         \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 ,
         \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 ,
         \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 ,
         \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 ,
         \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 ,
         \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 ,
         \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 ,
         \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 ,
         \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 ,
         \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 ,
         \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 ,
         \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 ,
         \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 ,
         \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 ,
         \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 ,
         \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 ,
         \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 ,
         \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 ,
         \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 ,
         \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 ,
         \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 ,
         \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 ,
         \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 ,
         \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 ,
         \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 ,
         \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 ,
         \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 ,
         \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 ,
         \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 ,
         \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 ,
         \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 ,
         \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 ,
         \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 ,
         \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 ,
         \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 ,
         \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 ,
         \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 ,
         \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 ,
         \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 ,
         \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 ,
         \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 ,
         \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 ,
         \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 ,
         \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 ,
         \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 ,
         \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 ,
         \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 ,
         \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 ,
         \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 ,
         \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 ,
         \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 ,
         \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 ,
         \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 ,
         \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 ,
         \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 ,
         \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 ,
         \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 ,
         \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 ,
         \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 ,
         \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 ,
         \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 ,
         \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 ,
         \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 ,
         \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 ,
         \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 ,
         \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 ,
         \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 ,
         \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 ,
         \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 ,
         \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 ,
         \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 ,
         \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 ,
         \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 ,
         \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 ,
         \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 ,
         \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 ,
         \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 ,
         \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 , \20003 , \20004 ,
         \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 ,
         \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 ,
         \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 ,
         \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 ,
         \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 ,
         \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 ,
         \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 ,
         \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 ,
         \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 ,
         \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 ,
         \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 ,
         \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 ,
         \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 ,
         \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 ,
         \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 ,
         \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 ,
         \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 ,
         \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 ,
         \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 ,
         \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 ,
         \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 ,
         \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 ,
         \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 ,
         \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 ,
         \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 ,
         \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 ,
         \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 ,
         \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 ,
         \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 ,
         \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 ,
         \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 ,
         \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 ,
         \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 ,
         \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 ,
         \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 ,
         \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 ,
         \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 ,
         \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 ,
         \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 ,
         \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 ,
         \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 ,
         \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 ,
         \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 ,
         \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 ,
         \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 ,
         \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 ,
         \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 ,
         \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 ,
         \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 ,
         \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 ,
         \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 ,
         \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 ,
         \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 ,
         \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 ,
         \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 ,
         \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 ,
         \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 ,
         \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 ,
         \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 ,
         \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 ,
         \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 ,
         \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 ,
         \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 ,
         \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 ,
         \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 ,
         \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 ,
         \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 ,
         \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 ,
         \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 ,
         \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 ,
         \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 ,
         \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 , \20723 , \20724 ,
         \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 ,
         \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 ,
         \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 ,
         \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 ,
         \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 ,
         \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 ,
         \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 ,
         \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 ,
         \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 ,
         \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 ,
         \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 ,
         \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 ,
         \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 ,
         \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 ,
         \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 ,
         \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 ,
         \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 ,
         \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 ,
         \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 ,
         \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 ,
         \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 ,
         \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 ,
         \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 ,
         \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 ,
         \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 ,
         \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 ,
         \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 ,
         \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 ,
         \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 ,
         \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 ,
         \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 ,
         \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 ,
         \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 ,
         \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 ,
         \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 ,
         \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 ,
         \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 ,
         \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 ,
         \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 ,
         \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 ,
         \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 ,
         \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 ,
         \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 ,
         \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 ,
         \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 ,
         \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 ,
         \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 ,
         \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 ,
         \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 ,
         \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 ,
         \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 ,
         \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 ,
         \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 ,
         \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 ,
         \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 ,
         \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 ,
         \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 ,
         \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 ,
         \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 ,
         \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 ,
         \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 ,
         \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 ,
         \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 ,
         \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 ,
         \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 ,
         \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 ,
         \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 ,
         \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 ,
         \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 ,
         \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 ,
         \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 ,
         \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 ,
         \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 ,
         \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 ,
         \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 ,
         \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 ,
         \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 ,
         \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 ,
         \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 ,
         \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 ,
         \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 ,
         \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 ,
         \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 ,
         \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 ,
         \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 ,
         \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 ,
         \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 ,
         \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 ,
         \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 ,
         \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 ,
         \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 ,
         \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 ,
         \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 , \21653 , \21654 ,
         \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 ,
         \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 ,
         \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 ,
         \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 ,
         \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 ,
         \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 ,
         \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 ,
         \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 ,
         \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 ,
         \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 ,
         \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 ,
         \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 ,
         \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 ,
         \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 ,
         \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 ,
         \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 ,
         \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 ,
         \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 ,
         \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 ,
         \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 ,
         \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 ,
         \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 ,
         \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 ,
         \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 ,
         \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 ,
         \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 ,
         \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 ,
         \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 ,
         \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 ,
         \21945_nR25610 , \21946 , \21947 , \21948 , \21949 , \21950_nR25642 , \21951 , \21952 , \21953 , \21954 ,
         \21955_nR25644 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961_nR25646 , \21962 , \21963 , \21964 ,
         \21965 , \21966 , \21967_nR25614 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 ,
         \21975 , \21976 , \21977 , \21978_nR25616 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 ,
         \21985 , \21986 , \21987 , \21988_nR25618 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 ,
         \21995 , \21996 , \21997 , \21998_nR2561a , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 ,
         \22005 , \22006 , \22007 , \22008_nR2561c , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 ,
         \22015 , \22016 , \22017 , \22018_nR2561e , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 ,
         \22025 , \22026 , \22027 , \22028_nR25620 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 ,
         \22035 , \22036 , \22037 , \22038_nR25622 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 ,
         \22045 , \22046 , \22047 , \22048_nR25612 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 ,
         \22055 , \22056 , \22057 , \22058_nR25624 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 ,
         \22065 , \22066 , \22067 , \22068_nR25626 , \22069 , \22070 , \22071 , \22072 , \22073 , \22074 ,
         \22075 , \22076 , \22077 , \22078_nR25628 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 ,
         \22085 , \22086 , \22087 , \22088_nR2562a , \22089 , \22090 , \22091 , \22092 , \22093 , \22094 ,
         \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 , \22103 , \22104 ,
         \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 , \22113 , \22114 ,
         \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 , \22123 , \22124 ,
         \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 , \22133 , \22134 ,
         \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 ,
         \22145_nR253fc , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 , \22153 , \22154 ,
         \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , \22163 , \22164 ,
         \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 , \22173_nR25412 , \22174 ,
         \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 , \22183 , \22184 ,
         \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , \22193_nR25428 , \22194 ,
         \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 ,
         \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 , \22213 , \22214 ,
         \22215 , \22216_nR2543e , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , \22223 , \22224 ,
         \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 ,
         \22235 , \22236 , \22237_nR25454 , \22238 , \22239 , \22240 , \22241 , \22242 , \22243 , \22244 ,
         \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 ,
         \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 , \22263 , \22264_nR2546a ,
         \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 , \22273 , \22274 ,
         \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 ,
         \22285_nR25474 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 ,
         \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 , \22303 , \22304 ,
         \22305 , \22306_nR25476 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 ,
         \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 ,
         \22325 , \22326 , \22327 , \22328_nR25478 , \22329 , \22330 , \22331 , \22332 , \22333 , \22334 ,
         \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 ,
         \22345 , \22346 , \22347 , \22348 , \22349_nR2547a , \22350 , \22351 , \22352 , \22353 , \22354 ,
         \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 , \22363 , \22364 ,
         \22365 , \22366 , \22367 , \22368 , \22369 , \22370_nR253fe , \22371 , \22372 , \22373 , \22374 ,
         \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 ,
         \22385 , \22386 , \22387 , \22388 , \22389 , \22390_nR25400 , \22391 , \22392 , \22393 , \22394 ,
         \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 ,
         \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411_nR25402 , \22412 , \22413 , \22414 ,
         \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 ,
         \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432_nR25404 , \22433 , \22434 ,
         \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 ,
         \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451_nR25406 , \22452 , \22453 , \22454 ,
         \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 ,
         \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471_nR25408 , \22472 , \22473 , \22474 ,
         \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 ,
         \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491_nR2540a , \22492 , \22493 , \22494 ,
         \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 ,
         \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512_nR2540c , \22513 , \22514 ,
         \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 ,
         \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532_nR2540e , \22533 , \22534 ,
         \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 ,
         \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552_nR25410 , \22553 , \22554 ,
         \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 ,
         \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572_nR25414 , \22573 , \22574 ,
         \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 ,
         \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592_nR25416 , \22593 , \22594 ,
         \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 , \22603 , \22604 ,
         \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612_nR25418 , \22613 , \22614 ,
         \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 ,
         \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632_nR2541a , \22633 , \22634 ,
         \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 ,
         \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653_nR2541c , \22654 ,
         \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 ,
         \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673_nR2541e , \22674 ,
         \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 ,
         \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694_nR25420 ,
         \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 ,
         \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 , \22714_nR25422 ,
         \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 ,
         \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734_nR25424 ,
         \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 ,
         \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754_nR25426 ,
         \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 ,
         \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 ,
         \22775 , \22776_nR2542a , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 , \22783 , \22784 ,
         \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 ,
         \22795 , \22796_nR2542c , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 ,
         \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 ,
         \22815 , \22816_nR2542e , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 ,
         \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 ,
         \22835 , \22836_nR25430 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 ,
         \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 ,
         \22855 , \22856_nR25432 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 ,
         \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 ,
         \22875 , \22876_nR25434 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 ,
         \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 ,
         \22895 , \22896_nR25436 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 ,
         \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914 ,
         \22915 , \22916 , \22917 , \22918_nR25438 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 ,
         \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 ,
         \22935 , \22936 , \22937 , \22938_nR2543a , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 ,
         \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 ,
         \22955 , \22956 , \22957 , \22958_nR2543c , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 ,
         \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 ,
         \22975 , \22976 , \22977 , \22978_nR25440 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 ,
         \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 ,
         \22995 , \22996 , \22997_nR25442 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 ,
         \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 ,
         \23015 , \23016_nR25444 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 ,
         \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 ,
         \23035 , \23036_nR25446 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 ,
         \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 ,
         \23055 , \23056 , \23057 , \23058_nR25448 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 ,
         \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 ,
         \23075 , \23076 , \23077 , \23078_nR2544a , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 ,
         \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 ,
         \23095 , \23096 , \23097 , \23098_nR2544c , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 ,
         \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 , \23114 ,
         \23115 , \23116 , \23117 , \23118_nR2544e , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 ,
         \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 ,
         \23135 , \23136 , \23137 , \23138_nR25450 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 ,
         \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 ,
         \23155 , \23156 , \23157 , \23158_nR25452 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 ,
         \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 ,
         \23175 , \23176 , \23177 , \23178_nR25456 , \23179 , \23180 , \23181 , \23182 , \23183 , \23184 ,
         \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 , \23193 , \23194 ,
         \23195 , \23196 , \23197_nR25458 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 ,
         \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 ,
         \23215 , \23216 , \23217_nR2545a , \23218 , \23219 , \23220 , \23221 , \23222 , \23223 , \23224 ,
         \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 ,
         \23235 , \23236 , \23237_nR2545c , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 ,
         \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 ,
         \23255 , \23256 , \23257_nR2545e , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 ,
         \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 , \23274 ,
         \23275 , \23276 , \23277_nR25460 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 ,
         \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 ,
         \23295 , \23296 , \23297_nR25462 , \23298 , \23299 , \23300 , \23301 , \23302 , \23303 , \23304 ,
         \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 ,
         \23315 , \23316_nR25464 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 ,
         \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 , \23333 , \23334 ,
         \23335 , \23336_nR25466 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 ,
         \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 ,
         \23355 , \23356_nR25468 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 ,
         \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 ,
         \23375 , \23376 , \23377_nR2546c , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 ,
         \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 ,
         \23395 , \23396 , \23397_nR2546e , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 ,
         \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 ,
         \23415 , \23416 , \23417_nR25470 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 ,
         \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 ,
         \23435 , \23436 , \23437_nR25472 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 ,
         \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 , \23453 , \23454 ,
         \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 ,
         \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471_nR2547c , \23472 , \23473 , \23474 ,
         \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483 , \23484 ,
         \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491_nR25492 , \23492 , \23493 , \23494 ,
         \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 ,
         \23505 , \23506 , \23507 , \23508 , \23509_nR254a8 , \23510 , \23511 , \23512 , \23513 , \23514 ,
         \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 ,
         \23525 , \23526 , \23527_nR254be , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 ,
         \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 ,
         \23545 , \23546 , \23547_nR254d4 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 ,
         \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 , \23563 , \23564 ,
         \23565 , \23566 , \23567 , \23568_nR254ea , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 ,
         \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 ,
         \23585 , \23586_nR254f4 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 ,
         \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 ,
         \23605_nR254f6 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 ,
         \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 , \23623_nR254f8 , \23624 ,
         \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 ,
         \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643_nR254fa , \23644 ,
         \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 ,
         \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662_nR2547e , \23663 , \23664 ,
         \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 , \23673 , \23674 ,
         \23675 , \23676 , \23677 , \23678 , \23679 , \23680_nR25480 , \23681 , \23682 , \23683 , \23684 ,
         \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 ,
         \23695 , \23696 , \23697 , \23698 , \23699_nR25482 , \23700 , \23701 , \23702 , \23703 , \23704 ,
         \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 ,
         \23715 , \23716 , \23717_nR25484 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 ,
         \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 ,
         \23735_nR25486 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 ,
         \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753_nR25488 , \23754 ,
         \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 ,
         \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772_nR2548a , \23773 , \23774 ,
         \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 , \23783 , \23784 ,
         \23785 , \23786 , \23787 , \23788 , \23789 , \23790_nR2548c , \23791 , \23792 , \23793 , \23794 ,
         \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 ,
         \23805 , \23806 , \23807 , \23808_nR2548e , \23809 , \23810 , \23811 , \23812 , \23813 , \23814 ,
         \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 ,
         \23825 , \23826_nR25490 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 ,
         \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844_nR25494 ,
         \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 ,
         \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862_nR25496 , \23863 , \23864 ,
         \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 ,
         \23875 , \23876 , \23877 , \23878 , \23879 , \23880_nR25498 , \23881 , \23882 , \23883 , \23884 ,
         \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 ,
         \23895 , \23896 , \23897 , \23898_nR2549a , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 ,
         \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 ,
         \23915 , \23916_nR2549c , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 ,
         \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934_nR2549e ,
         \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 ,
         \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953_nR254a0 , \23954 ,
         \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 ,
         \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971_nR254a2 , \23972 , \23973 , \23974 ,
         \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 ,
         \23985 , \23986 , \23987 , \23988 , \23989_nR254a4 , \23990 , \23991 , \23992 , \23993 , \23994 ,
         \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 , \24003 , \24004 ,
         \24005 , \24006 , \24007_nR254a6 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 ,
         \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 ,
         \24025_nR254aa , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 ,
         \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043_nR254ac , \24044 ,
         \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 ,
         \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061_nR254ae , \24062 , \24063 , \24064 ,
         \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 ,
         \24075 , \24076 , \24077 , \24078 , \24079_nR254b0 , \24080 , \24081 , \24082 , \24083 , \24084 ,
         \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 ,
         \24095 , \24096 , \24097_nR254b2 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 ,
         \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 ,
         \24115_nR254b4 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 ,
         \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133 , \24134 ,
         \24135_nR254b6 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 , \24143 , \24144 ,
         \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153_nR254b8 , \24154 ,
         \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 , \24163 , \24164 ,
         \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173_nR254ba , \24174 ,
         \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 , \24183 , \24184 ,
         \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191_nR254bc , \24192 , \24193 , \24194 ,
         \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 ,
         \24205 , \24206 , \24207 , \24208 , \24209_nR254c0 , \24210 , \24211 , \24212 , \24213 , \24214 ,
         \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 ,
         \24225 , \24226 , \24227_nR254c2 , \24228 , \24229 , \24230 , \24231 , \24232 , \24233 , \24234 ,
         \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 , \24243 , \24244 ,
         \24245_nR254c4 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 ,
         \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263_nR254c6 , \24264 ,
         \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 ,
         \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281_nR254c8 , \24282 , \24283 , \24284 ,
         \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 ,
         \24295 , \24296 , \24297 , \24298 , \24299_nR254ca , \24300 , \24301 , \24302 , \24303 , \24304 ,
         \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 ,
         \24315 , \24316 , \24317_nR254cc , \24318 , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 ,
         \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333 , \24334 ,
         \24335_nR254ce , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 ,
         \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 , \24353_nR254d0 , \24354 ,
         \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 ,
         \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371_nR254d2 , \24372 , \24373 , \24374 ,
         \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 , \24383 , \24384 ,
         \24385 , \24386 , \24387 , \24388 , \24389_nR254d6 , \24390 , \24391 , \24392 , \24393 , \24394 ,
         \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 ,
         \24405 , \24406 , \24407_nR254d8 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413 , \24414 ,
         \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 ,
         \24425 , \24426_nR254da , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 , \24433 , \24434 ,
         \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444_nR254dc ,
         \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 ,
         \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462_nR254de , \24463 , \24464 ,
         \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 ,
         \24475 , \24476 , \24477 , \24478 , \24479 , \24480_nR254e0 , \24481 , \24482 , \24483 , \24484 ,
         \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494 ,
         \24495 , \24496 , \24497 , \24498_nR254e2 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 ,
         \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 , \24513 , \24514 ,
         \24515 , \24516_nR254e4 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 ,
         \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534_nR254e6 ,
         \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 , \24543 , \24544 ,
         \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552_nR254e8 , \24553 , \24554 ,
         \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 ,
         \24565 , \24566 , \24567 , \24568 , \24569 , \24570_nR254ec , \24571 , \24572 , \24573 , \24574 ,
         \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 ,
         \24585 , \24586 , \24587 , \24588_nR254ee , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 ,
         \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 ,
         \24605 , \24606_nR254f0 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 ,
         \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624_nR254f2 ,
         \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 ,
         \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 , \24643 , \24644 ,
         \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 ,
         \24655 , \24656_nR254fc , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 ,
         \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 ,
         \24675_nR25512 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 ,
         \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692_nR25528 , \24693 , \24694 ,
         \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 ,
         \24705 , \24706 , \24707 , \24708 , \24709 , \24710_nR2553e , \24711 , \24712 , \24713 , \24714 ,
         \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 ,
         \24725 , \24726 , \24727 , \24728 , \24729_nR25554 , \24730 , \24731 , \24732 , \24733 , \24734 ,
         \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 ,
         \24745 , \24746 , \24747_nR2556a , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 ,
         \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764_nR25574 ,
         \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 , \24773 , \24774 ,
         \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781_nR25576 , \24782 , \24783 , \24784 ,
         \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 ,
         \24795 , \24796 , \24797 , \24798_nR25578 , \24799 , \24800 , \24801 , \24802 , \24803 , \24804 ,
         \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 ,
         \24815 , \24816_nR2557a , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 ,
         \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834_nR254fe ,
         \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 ,
         \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851_nR25500 , \24852 , \24853 , \24854 ,
         \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 ,
         \24865 , \24866 , \24867 , \24868_nR25502 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 ,
         \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 , \24883 , \24884 ,
         \24885_nR25504 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 ,
         \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902_nR25506 , \24903 , \24904 ,
         \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 ,
         \24915 , \24916 , \24917 , \24918 , \24919 , \24920_nR25508 , \24921 , \24922 , \24923 , \24924 ,
         \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 , \24934 ,
         \24935 , \24936 , \24937_nR2550a , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 ,
         \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954_nR2550c ,
         \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 , \24963 , \24964 ,
         \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971_nR2550e , \24972 , \24973 , \24974 ,
         \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 ,
         \24985 , \24986 , \24987 , \24988_nR25510 , \24989 , \24990 , \24991 , \24992 , \24993 , \24994 ,
         \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 ,
         \25005_nR25514 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 ,
         \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022_nR25516 , \25023 , \25024 ,
         \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 ,
         \25035 , \25036 , \25037 , \25038 , \25039_nR25518 , \25040 , \25041 , \25042 , \25043 , \25044 ,
         \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 ,
         \25055 , \25056_nR2551a , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 ,
         \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073_nR2551c , \25074 ,
         \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 ,
         \25085 , \25086 , \25087 , \25088 , \25089 , \25090_nR2551e , \25091 , \25092 , \25093 , \25094 ,
         \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 ,
         \25105 , \25106 , \25107_nR25520 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 ,
         \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124_nR25522 ,
         \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 , \25133 , \25134 ,
         \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141_nR25524 , \25142 , \25143 , \25144 ,
         \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 ,
         \25155 , \25156 , \25157 , \25158_nR25526 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 ,
         \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 ,
         \25175_nR2552a , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 ,
         \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192_nR2552c , \25193 , \25194 ,
         \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 ,
         \25205 , \25206 , \25207 , \25208 , \25209_nR2552e , \25210 , \25211 , \25212 , \25213 , \25214 ,
         \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 ,
         \25225 , \25226_nR25530 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 ,
         \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243_nR25532 , \25244 ,
         \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 ,
         \25255 , \25256 , \25257 , \25258 , \25259 , \25260_nR25534 , \25261 , \25262 , \25263 , \25264 ,
         \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 , \25273 , \25274 ,
         \25275 , \25276 , \25277_nR25536 , \25278 , \25279 , \25280 , \25281 , \25282 , \25283 , \25284 ,
         \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294_nR25538 ,
         \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 ,
         \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311_nR2553a , \25312 , \25313 , \25314 ,
         \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 ,
         \25325 , \25326 , \25327 , \25328_nR2553c , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 ,
         \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 ,
         \25345_nR25540 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 ,
         \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362_nR25542 , \25363 , \25364 ,
         \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 ,
         \25375 , \25376 , \25377 , \25378 , \25379_nR25544 , \25380 , \25381 , \25382 , \25383 , \25384 ,
         \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 , \25393 , \25394 ,
         \25395 , \25396_nR25546 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 ,
         \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413_nR25548 , \25414 ,
         \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 , \25423 , \25424 ,
         \25425 , \25426 , \25427 , \25428 , \25429 , \25430_nR2554a , \25431 , \25432 , \25433 , \25434 ,
         \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 ,
         \25445 , \25446 , \25447_nR2554c , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 ,
         \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 ,
         \25465_nR2554e , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 , \25473 , \25474 ,
         \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482_nR25550 , \25483 , \25484 ,
         \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 ,
         \25495 , \25496 , \25497 , \25498 , \25499_nR25552 , \25500 , \25501 , \25502 , \25503 , \25504 ,
         \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 ,
         \25515 , \25516_nR25556 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 ,
         \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533_nR25558 , \25534 ,
         \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 ,
         \25545 , \25546 , \25547 , \25548 , \25549 , \25550_nR2555a , \25551 , \25552 , \25553 , \25554 ,
         \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 ,
         \25565 , \25566 , \25567_nR2555c , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 ,
         \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584_nR2555e ,
         \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 ,
         \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601_nR25560 , \25602 , \25603 , \25604 ,
         \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 ,
         \25615 , \25616 , \25617 , \25618_nR25562 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 ,
         \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 , \25634 ,
         \25635_nR25564 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 ,
         \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653_nR25566 , \25654 ,
         \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 ,
         \25665 , \25666 , \25667 , \25668 , \25669 , \25670_nR25568 , \25671 , \25672 , \25673 , \25674 ,
         \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 ,
         \25685 , \25686 , \25687_nR2556c , \25688 , \25689 , \25690 , \25691 , \25692 , \25693 , \25694 ,
         \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704_nR2556e ,
         \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713 , \25714 ,
         \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721_nR25570 , \25722 , \25723 , \25724 ,
         \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 ,
         \25735 , \25736 , \25737 , \25738_nR25572 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 ,
         \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 ,
         \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 ,
         \25765_nR2557c , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 , \25773 , \25774 ,
         \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781_nR25592 , \25782 , \25783 , \25784 ,
         \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 , \25793 , \25794 ,
         \25795 , \25796 , \25797 , \25798_nR255a8 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 ,
         \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 , \25813 , \25814_nR255be ,
         \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 ,
         \25825 , \25826 , \25827 , \25828_nR255d4 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 ,
         \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843_nR255ea , \25844 ,
         \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 ,
         \25855 , \25856 , \25857_nR255f4 , \25858 , \25859 , \25860 , \25861 , \25862 , \25863 , \25864 ,
         \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871_nR255f6 , \25872 , \25873 , \25874 ,
         \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 ,
         \25885_nR255f8 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 ,
         \25895 , \25896 , \25897 , \25898 , \25899 , \25900_nR255fa , \25901 , \25902 , \25903 , \25904 ,
         \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914_nR2557e ,
         \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 ,
         \25925 , \25926 , \25927 , \25928_nR25580 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 ,
         \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942_nR25582 , \25943 , \25944 ,
         \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 ,
         \25955 , \25956_nR25584 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 ,
         \25965 , \25966 , \25967 , \25968 , \25969 , \25970_nR25586 , \25971 , \25972 , \25973 , \25974 ,
         \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984_nR25588 ,
         \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 ,
         \25995 , \25996 , \25997 , \25998_nR2558a , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 ,
         \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012_nR2558c , \26013 , \26014 ,
         \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 ,
         \26025 , \26026_nR2558e , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 ,
         \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041_nR25590 , \26042 , \26043 , \26044 ,
         \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 ,
         \26055_nR25594 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 ,
         \26065 , \26066 , \26067 , \26068 , \26069_nR25596 , \26070 , \26071 , \26072 , \26073 , \26074 ,
         \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083_nR25598 , \26084 ,
         \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 ,
         \26095 , \26096 , \26097_nR2559a , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 ,
         \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111_nR2559c , \26112 , \26113 , \26114 ,
         \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 ,
         \26125_nR2559e , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 ,
         \26135 , \26136 , \26137 , \26138 , \26139_nR255a0 , \26140 , \26141 , \26142 , \26143 , \26144 ,
         \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153_nR255a2 , \26154 ,
         \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 ,
         \26165 , \26166 , \26167_nR255a4 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 ,
         \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181_nR255a6 , \26182 , \26183 , \26184 ,
         \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 ,
         \26195 , \26196_nR255aa , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 ,
         \26205 , \26206 , \26207 , \26208 , \26209 , \26210_nR255ac , \26211 , \26212 , \26213 , \26214 ,
         \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224_nR255ae ,
         \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 ,
         \26235 , \26236 , \26237 , \26238_nR255b0 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 ,
         \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252_nR255b2 , \26253 , \26254 ,
         \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 ,
         \26265 , \26266_nR255b4 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273 , \26274 ,
         \26275 , \26276 , \26277 , \26278 , \26279 , \26280_nR255b6 , \26281 , \26282 , \26283 , \26284 ,
         \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294_nR255b8 ,
         \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 ,
         \26305 , \26306 , \26307 , \26308_nR255ba , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 ,
         \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322_nR255bc , \26323 , \26324 ,
         \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 ,
         \26335 , \26336_nR255c0 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 , \26343 , \26344 ,
         \26345 , \26346 , \26347 , \26348 , \26349 , \26350_nR255c2 , \26351 , \26352 , \26353 , \26354 ,
         \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 , \26363 , \26364_nR255c4 ,
         \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 ,
         \26375 , \26376 , \26377 , \26378_nR255c6 , \26379 , \26380 , \26381 , \26382 , \26383 , \26384 ,
         \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392_nR255c8 , \26393 , \26394 ,
         \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404 ,
         \26405 , \26406_nR255ca , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 , \26413 , \26414 ,
         \26415 , \26416 , \26417 , \26418 , \26419 , \26420_nR255cc , \26421 , \26422 , \26423 , \26424 ,
         \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 , \26433 , \26434_nR255ce ,
         \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 , \26443 , \26444 ,
         \26445 , \26446 , \26447 , \26448_nR255d0 , \26449 , \26450 , \26451 , \26452 , \26453 , \26454 ,
         \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462_nR255d2 , \26463 , \26464 ,
         \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 , \26473 , \26474 ,
         \26475 , \26476_nR255d6 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 , \26483 , \26484 ,
         \26485 , \26486 , \26487 , \26488 , \26489 , \26490_nR255d8 , \26491 , \26492 , \26493 , \26494 ,
         \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 , \26503 , \26504_nR255da ,
         \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 ,
         \26515 , \26516 , \26517 , \26518_nR255dc , \26519 , \26520 , \26521 , \26522 , \26523 , \26524 ,
         \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532_nR255de , \26533 , \26534 ,
         \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 ,
         \26545 , \26546_nR255e0 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 , \26553 , \26554 ,
         \26555 , \26556 , \26557 , \26558 , \26559 , \26560_nR255e2 , \26561 , \26562 , \26563 , \26564 ,
         \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574_nR255e4 ,
         \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584 ,
         \26585 , \26586 , \26587 , \26588_nR255e6 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 ,
         \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602_nR255e8 , \26603 , \26604 ,
         \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 ,
         \26615 , \26616_nR255ec , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 ,
         \26625 , \26626 , \26627 , \26628 , \26629 , \26630_nR255ee , \26631 , \26632 , \26633 , \26634 ,
         \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644_nR255f0 ,
         \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654 ,
         \26655 , \26656 , \26657 , \26658_nR255f2 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 ,
         \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 , \26673 , \26674 ,
         \26675 , \26676 , \26677_nR253bc , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 ,
         \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 ,
         \26695_nR253be , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704 ,
         \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712_nR253c0 , \26713 , \26714 ,
         \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 , \26723 , \26724 ,
         \26725 , \26726 , \26727 , \26728 , \26729_nR253c2 , \26730 , \26731 , \26732 , \26733 , \26734 ,
         \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 ,
         \26745 , \26746_nR253c4 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 ,
         \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763_nR253c6 , \26764 ,
         \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 , \26773 , \26774 ,
         \26775 , \26776 , \26777 , \26778 , \26779 , \26780_nR253c8 , \26781 , \26782 , \26783 , \26784 ,
         \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 ,
         \26795 , \26796 , \26797_nR253ca , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804 ,
         \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812_nR253cc , \26813 , \26814 ,
         \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 , \26823 , \26824 ,
         \26825 , \26826 , \26827_nR253ce , \26828 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 ,
         \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842_nR253d0 , \26843 , \26844 ,
         \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 , \26853 , \26854 ,
         \26855 , \26856 , \26857_nR253d2 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 ,
         \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872_nR253d4 , \26873 , \26874 ,
         \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 , \26883 , \26884 ,
         \26885 , \26886 , \26887_nR253d6 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 ,
         \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902_nR253d8 , \26903 , \26904 ,
         \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 ,
         \26915 , \26916 , \26917_nR253da , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 ,
         \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932_nR253dc , \26933 , \26934 ,
         \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 ,
         \26945 , \26946 , \26947_nR253de , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 ,
         \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962_nR253e0 , \26963 , \26964 ,
         \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 ,
         \26975 , \26976 , \26977_nR253e2 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 ,
         \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992_nR253e4 , \26993 , \26994 ,
         \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 ,
         \27005 , \27006 , \27007_nR253e6 , \27008 , \27009 , \27010 , \27011 , \27012 , \27013 , \27014 ,
         \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022_nR253e8 , \27023 , \27024 ,
         \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 ,
         \27035 , \27036 , \27037_nR253ea , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 ,
         \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052_nR253ec , \27053 , \27054 ,
         \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 ,
         \27065 , \27066 , \27067_nR253ee , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 ,
         \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082_nR253f0 , \27083 , \27084 ,
         \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 , \27094 ,
         \27095 , \27096 , \27097_nR253f2 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 ,
         \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112_nR253f4 , \27113 , \27114 ,
         \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 ,
         \27125 , \27126 , \27127_nR253f6 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 ,
         \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142_nR253f8 , \27143 , \27144 ,
         \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 ,
         \27155 , \27156 , \27157_nR253fa , \27158 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 ,
         \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174_nR25666 ,
         \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 ,
         \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 ,
         \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 ,
         \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 ,
         \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 ,
         \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 ,
         \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 ,
         \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 ,
         \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 ,
         \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 ,
         \27275 , \27276 , \27277 , \27278 , \27279_nR22c68 , \27280 , \27281 , \27282 , \27283 , \27284 ,
         \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 , \27293 , \27294 ,
         \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 , \27303 , \27304 ,
         \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 , \27313 , \27314 ,
         \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 ,
         \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 ,
         \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344_nR22c59 ,
         \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 ,
         \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 , \27363 , \27364 ,
         \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 ,
         \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 ,
         \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 , \27393 , \27394 ,
         \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 ,
         \27405 , \27406 , \27407 , \27408 , \27409 , \27410_nR23ca4 , \27411 , \27412 , \27413 , \27414 ,
         \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 ,
         \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 ,
         \27435 , \27436 , \27437 , \27438_nR23cba , \27439 , \27440 , \27441 , \27442 , \27443 , \27444 ,
         \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 ,
         \27455 , \27456_nR23cd0 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 ,
         \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 , \27473 , \27474 ,
         \27475 , \27476 , \27477_nR23ce6 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 ,
         \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 ,
         \27495 , \27496 , \27497_nR23cfc , \27498 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 ,
         \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 ,
         \27515 , \27516 , \27517 , \27518_nR23d12 , \27519 , \27520 , \27521 , \27522 , \27523 , \27524 ,
         \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 ,
         \27535 , \27536 , \27537_nR23d1c , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 ,
         \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 , \27553 , \27554 ,
         \27555 , \27556_nR23d1e , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 ,
         \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 ,
         \27575 , \27576 , \27577 , \27578_nR23d20 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 ,
         \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 ,
         \27595 , \27596 , \27597 , \27598 , \27599_nR23d22 , \27600 , \27601 , \27602 , \27603 , \27604 ,
         \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 ,
         \27615 , \27616 , \27617 , \27618 , \27619_nR23ca6 , \27620 , \27621 , \27622 , \27623 , \27624 ,
         \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 , \27633 , \27634 ,
         \27635 , \27636 , \27637 , \27638_nR23ca8 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 ,
         \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 ,
         \27655 , \27656 , \27657 , \27658_nR23caa , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 ,
         \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 ,
         \27675 , \27676 , \27677 , \27678_nR23cac , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 ,
         \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 ,
         \27695 , \27696_nR23cae , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 ,
         \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714_nR23cb0 ,
         \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 ,
         \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732_nR23cb2 , \27733 , \27734 ,
         \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 ,
         \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751_nR23cb4 , \27752 , \27753 , \27754 ,
         \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 ,
         \27765 , \27766 , \27767 , \27768 , \27769 , \27770_nR23cb6 , \27771 , \27772 , \27773 , \27774 ,
         \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 ,
         \27785 , \27786 , \27787 , \27788 , \27789_nR23cb8 , \27790 , \27791 , \27792 , \27793 , \27794 ,
         \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 ,
         \27805 , \27806 , \27807 , \27808 , \27809_nR23cbc , \27810 , \27811 , \27812 , \27813 , \27814 ,
         \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 ,
         \27825 , \27826 , \27827_nR23cbe , \27828 , \27829 , \27830 , \27831 , \27832 , \27833 , \27834 ,
         \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 , \27843 , \27844 ,
         \27845_nR23cc0 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 ,
         \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 , \27863 , \27864_nR23cc2 ,
         \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 ,
         \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883_nR23cc4 , \27884 ,
         \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 ,
         \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902_nR23cc6 , \27903 , \27904 ,
         \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 ,
         \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921_nR23cc8 , \27922 , \27923 , \27924 ,
         \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 ,
         \27935 , \27936 , \27937 , \27938 , \27939 , \27940_nR23cca , \27941 , \27942 , \27943 , \27944 ,
         \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 , \27953 , \27954 ,
         \27955 , \27956 , \27957 , \27958 , \27959_nR23ccc , \27960 , \27961 , \27962 , \27963 , \27964 ,
         \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 , \27973 , \27974 ,
         \27975 , \27976 , \27977 , \27978_nR23cce , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 ,
         \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 ,
         \27995 , \27996 , \27997 , \27998_nR23cd2 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 ,
         \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 ,
         \28015 , \28016 , \28017 , \28018 , \28019_nR23cd4 , \28020 , \28021 , \28022 , \28023 , \28024 ,
         \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 , \28033 , \28034 ,
         \28035 , \28036 , \28037 , \28038 , \28039_nR23cd6 , \28040 , \28041 , \28042 , \28043 , \28044 ,
         \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 ,
         \28055 , \28056 , \28057 , \28058_nR23cd8 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 ,
         \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 ,
         \28075 , \28076_nR23cda , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 ,
         \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 ,
         \28095_nR23cdc , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 ,
         \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 , \28113 , \28114_nR23cde ,
         \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 ,
         \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133_nR23ce0 , \28134 ,
         \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 , \28143 , \28144 ,
         \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152_nR23ce2 , \28153 , \28154 ,
         \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 ,
         \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171_nR23ce4 , \28172 , \28173 , \28174 ,
         \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 ,
         \28185 , \28186 , \28187 , \28188 , \28189 , \28190_nR23ce8 , \28191 , \28192 , \28193 , \28194 ,
         \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 ,
         \28205 , \28206 , \28207 , \28208 , \28209_nR23cea , \28210 , \28211 , \28212 , \28213 , \28214 ,
         \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 , \28223 , \28224 ,
         \28225 , \28226 , \28227 , \28228_nR23cec , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 ,
         \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 ,
         \28245 , \28246 , \28247_nR23cee , \28248 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 ,
         \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 ,
         \28265 , \28266 , \28267_nR23cf0 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 ,
         \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 ,
         \28285 , \28286_nR23cf2 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 ,
         \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 ,
         \28305_nR23cf4 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 ,
         \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324_nR23cf6 ,
         \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 ,
         \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343_nR23cf8 , \28344 ,
         \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 ,
         \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362_nR23cfa , \28363 , \28364 ,
         \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 ,
         \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382_nR23cfe , \28383 , \28384 ,
         \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 , \28393 , \28394 ,
         \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402_nR23d00 , \28403 , \28404 ,
         \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 ,
         \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422_nR23d02 , \28423 , \28424 ,
         \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 ,
         \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442_nR23d04 , \28443 , \28444 ,
         \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 ,
         \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462_nR23d06 , \28463 , \28464 ,
         \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 ,
         \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481_nR23d08 , \28482 , \28483 , \28484 ,
         \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 ,
         \28495 , \28496 , \28497 , \28498 , \28499 , \28500_nR23d0a , \28501 , \28502 , \28503 , \28504 ,
         \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 ,
         \28515 , \28516 , \28517 , \28518 , \28519 , \28520_nR23d0c , \28521 , \28522 , \28523 , \28524 ,
         \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 , \28533 , \28534 ,
         \28535 , \28536 , \28537 , \28538 , \28539_nR23d0e , \28540 , \28541 , \28542 , \28543 , \28544 ,
         \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 , \28553 , \28554 ,
         \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561_nR23d10 , \28562 , \28563 , \28564 ,
         \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 , \28573 , \28574 ,
         \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581_nR23d14 , \28582 , \28583 , \28584 ,
         \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 ,
         \28595 , \28596 , \28597 , \28598 , \28599_nR23d16 , \28600 , \28601 , \28602 , \28603 , \28604 ,
         \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 ,
         \28615 , \28616 , \28617 , \28618_nR23d18 , \28619 , \28620 , \28621 , \28622 , \28623 , \28624 ,
         \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 ,
         \28635 , \28636_nR23d1a , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 , \28643 , \28644 ,
         \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 , \28653 , \28654 ,
         \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 , \28663 , \28664 ,
         \28665 , \28666 , \28667 , \28668_nR23d24 , \28669 , \28670 , \28671 , \28672 , \28673 , \28674 ,
         \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 , \28683 , \28684 ,
         \28685 , \28686 , \28687 , \28688 , \28689_nR23d3a , \28690 , \28691 , \28692 , \28693 , \28694 ,
         \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 , \28703 , \28704 ,
         \28705 , \28706 , \28707 , \28708_nR23d50 , \28709 , \28710 , \28711 , \28712 , \28713 , \28714 ,
         \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 , \28723 , \28724 ,
         \28725 , \28726 , \28727 , \28728_nR23d66 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 ,
         \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 , \28743 , \28744 ,
         \28745 , \28746 , \28747_nR23d7c , \28748 , \28749 , \28750 , \28751 , \28752 , \28753 , \28754 ,
         \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 ,
         \28765 , \28766 , \28767_nR23d92 , \28768 , \28769 , \28770 , \28771 , \28772 , \28773 , \28774 ,
         \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 ,
         \28785 , \28786_nR23d9c , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 , \28793 , \28794 ,
         \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804_nR23d9e ,
         \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 ,
         \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822_nR23da0 , \28823 , \28824 ,
         \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 ,
         \28835 , \28836 , \28837 , \28838_nR23da2 , \28839 , \28840 , \28841 , \28842 , \28843 , \28844 ,
         \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 ,
         \28855_nR23d26 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 , \28863 , \28864 ,
         \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871_nR23d28 , \28872 , \28873 , \28874 ,
         \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 , \28883 , \28884 ,
         \28885 , \28886 , \28887_nR23d2a , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 ,
         \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904_nR23d2c ,
         \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 ,
         \28915 , \28916 , \28917 , \28918 , \28919 , \28920_nR23d2e , \28921 , \28922 , \28923 , \28924 ,
         \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , \28933 , \28934 ,
         \28935 , \28936 , \28937_nR23d30 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 ,
         \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 , \28953 , \28954_nR23d32 ,
         \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 ,
         \28965 , \28966 , \28967 , \28968 , \28969 , \28970_nR23d34 , \28971 , \28972 , \28973 , \28974 ,
         \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 ,
         \28985 , \28986_nR23d36 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 ,
         \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004_nR23d38 ,
         \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014 ,
         \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022_nR23d3c , \29023 , \29024 ,
         \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 ,
         \29035 , \29036 , \29037 , \29038 , \29039 , \29040_nR23d3e , \29041 , \29042 , \29043 , \29044 ,
         \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 ,
         \29055 , \29056 , \29057 , \29058_nR23d40 , \29059 , \29060 , \29061 , \29062 , \29063 , \29064 ,
         \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 ,
         \29075 , \29076_nR23d42 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 , \29083 , \29084 ,
         \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094_nR23d44 ,
         \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 ,
         \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112_nR23d46 , \29113 , \29114 ,
         \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 ,
         \29125 , \29126 , \29127 , \29128 , \29129 , \29130_nR23d48 , \29131 , \29132 , \29133 , \29134 ,
         \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 , \29143 , \29144 ,
         \29145 , \29146 , \29147 , \29148_nR23d4a , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 ,
         \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 ,
         \29165 , \29166_nR23d4c , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 ,
         \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 , \29183 , \29184_nR23d4e ,
         \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 , \29193 , \29194 ,
         \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202_nR23d52 , \29203 , \29204 ,
         \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 ,
         \29215 , \29216 , \29217 , \29218 , \29219 , \29220_nR23d54 , \29221 , \29222 , \29223 , \29224 ,
         \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 ,
         \29235 , \29236 , \29237 , \29238_nR23d56 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 ,
         \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 ,
         \29255 , \29256_nR23d58 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 ,
         \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 , \29274_nR23d5a ,
         \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 ,
         \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292_nR23d5c , \29293 , \29294 ,
         \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 , \29303 , \29304 ,
         \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311_nR23d5e , \29312 , \29313 , \29314 ,
         \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 ,
         \29325 , \29326 , \29327_nR23d60 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 ,
         \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 ,
         \29345_nR23d62 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 ,
         \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361_nR23d64 , \29362 , \29363 , \29364 ,
         \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 ,
         \29375 , \29376 , \29377_nR23d68 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 ,
         \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393_nR23d6a , \29394 ,
         \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 ,
         \29405 , \29406 , \29407 , \29408 , \29409_nR23d6c , \29410 , \29411 , \29412 , \29413 , \29414 ,
         \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 ,
         \29425_nR23d6e , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433 , \29434 ,
         \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443_nR23d70 , \29444 ,
         \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 ,
         \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461_nR23d72 , \29462 , \29463 , \29464 ,
         \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 ,
         \29475 , \29476 , \29477 , \29478 , \29479_nR23d74 , \29480 , \29481 , \29482 , \29483 , \29484 ,
         \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 ,
         \29495 , \29496 , \29497_nR23d76 , \29498 , \29499 , \29500 , \29501 , \29502 , \29503 , \29504 ,
         \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 ,
         \29515_nR23d78 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 ,
         \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533_nR23d7a , \29534 ,
         \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 , \29543 , \29544 ,
         \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551_nR23d7e , \29552 , \29553 , \29554 ,
         \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 ,
         \29565 , \29566 , \29567 , \29568 , \29569_nR23d80 , \29570 , \29571 , \29572 , \29573 , \29574 ,
         \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 ,
         \29585 , \29586 , \29587 , \29588_nR23d82 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 ,
         \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 ,
         \29605 , \29606_nR23d84 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 ,
         \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624_nR23d86 ,
         \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 ,
         \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642_nR23d88 , \29643 , \29644 ,
         \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 ,
         \29655 , \29656 , \29657 , \29658 , \29659 , \29660_nR23d8a , \29661 , \29662 , \29663 , \29664 ,
         \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 ,
         \29675 , \29676 , \29677 , \29678_nR23d8c , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 ,
         \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 ,
         \29695 , \29696_nR23d8e , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 , \29703 , \29704 ,
         \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714_nR23d90 ,
         \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 ,
         \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732_nR23d94 , \29733 , \29734 ,
         \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 ,
         \29745 , \29746 , \29747 , \29748 , \29749 , \29750_nR23d96 , \29751 , \29752 , \29753 , \29754 ,
         \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 ,
         \29765 , \29766 , \29767 , \29768_nR23d98 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 ,
         \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 ,
         \29785 , \29786_nR23d9a , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 ,
         \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 ,
         \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 ,
         \29815 , \29816 , \29817_nR23da4 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 ,
         \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833 , \29834 ,
         \29835 , \29836 , \29837_nR23dba , \29838 , \29839 , \29840 , \29841 , \29842 , \29843 , \29844 ,
         \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 ,
         \29855_nR23dd0 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 ,
         \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873_nR23de6 , \29874 ,
         \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 ,
         \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891_nR23dfc , \29892 , \29893 , \29894 ,
         \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 ,
         \29905 , \29906 , \29907 , \29908 , \29909 , \29910_nR23e12 , \29911 , \29912 , \29913 , \29914 ,
         \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 , \29923 , \29924 ,
         \29925 , \29926 , \29927 , \29928_nR23e1c , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 ,
         \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 ,
         \29945_nR23e1e , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 ,
         \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962_nR23e20 , \29963 , \29964 ,
         \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 , \29974 ,
         \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981_nR23e22 , \29982 , \29983 , \29984 ,
         \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 ,
         \29995 , \29996 , \29997 , \29998_nR23da6 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 ,
         \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 ,
         \30015_nR23da8 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 ,
         \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031_nR23daa , \30032 , \30033 , \30034 ,
         \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 , \30044 ,
         \30045 , \30046 , \30047_nR23dac , \30048 , \30049 , \30050 , \30051 , \30052 , \30053 , \30054 ,
         \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063_nR23dae , \30064 ,
         \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073 , \30074 ,
         \30075 , \30076 , \30077 , \30078 , \30079_nR23db0 , \30080 , \30081 , \30082 , \30083 , \30084 ,
         \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 ,
         \30095_nR23db2 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 ,
         \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111_nR23db4 , \30112 , \30113 , \30114 ,
         \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 ,
         \30125 , \30126 , \30127 , \30128_nR23db6 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 ,
         \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 , \30143 , \30144_nR23db8 ,
         \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 ,
         \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161_nR23dbc , \30162 , \30163 , \30164 ,
         \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 ,
         \30175 , \30176 , \30177 , \30178_nR23dbe , \30179 , \30180 , \30181 , \30182 , \30183 , \30184 ,
         \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 ,
         \30195_nR23dc0 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 ,
         \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212_nR23dc2 , \30213 , \30214 ,
         \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 ,
         \30225 , \30226 , \30227 , \30228 , \30229_nR23dc4 , \30230 , \30231 , \30232 , \30233 , \30234 ,
         \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 , \30243 , \30244 ,
         \30245 , \30246_nR23dc6 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 ,
         \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263_nR23dc8 , \30264 ,
         \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 ,
         \30275 , \30276 , \30277 , \30278 , \30279 , \30280_nR23dca , \30281 , \30282 , \30283 , \30284 ,
         \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 , \30293 , \30294 ,
         \30295 , \30296 , \30297_nR23dcc , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 ,
         \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314_nR23dce ,
         \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 , \30323 , \30324 ,
         \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331_nR23dd2 , \30332 , \30333 , \30334 ,
         \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 ,
         \30345 , \30346 , \30347 , \30348_nR23dd4 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 ,
         \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 ,
         \30365_nR23dd6 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 , \30373 , \30374 ,
         \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382_nR23dd8 , \30383 , \30384 ,
         \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 ,
         \30395 , \30396 , \30397 , \30398 , \30399_nR23dda , \30400 , \30401 , \30402 , \30403 , \30404 ,
         \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 ,
         \30415_nR23ddc , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 ,
         \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431_nR23dde , \30432 , \30433 , \30434 ,
         \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 ,
         \30445 , \30446 , \30447_nR23de0 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 , \30454 ,
         \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463_nR23de2 , \30464 ,
         \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 ,
         \30475 , \30476 , \30477 , \30478 , \30479_nR23de4 , \30480 , \30481 , \30482 , \30483 , \30484 ,
         \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 ,
         \30495_nR23de8 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 ,
         \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511_nR23dea , \30512 , \30513 , \30514 ,
         \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 ,
         \30525 , \30526 , \30527 , \30528 , \30529_nR23dec , \30530 , \30531 , \30532 , \30533 , \30534 ,
         \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 ,
         \30545 , \30546 , \30547_nR23dee , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 ,
         \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564_nR23df0 ,
         \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 ,
         \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582_nR23df2 , \30583 , \30584 ,
         \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 ,
         \30595 , \30596 , \30597 , \30598 , \30599_nR23df4 , \30600 , \30601 , \30602 , \30603 , \30604 ,
         \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 ,
         \30615 , \30616 , \30617_nR23df6 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 ,
         \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634_nR23df8 ,
         \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 ,
         \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651_nR23dfa , \30652 , \30653 , \30654 ,
         \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 ,
         \30665 , \30666 , \30667 , \30668_nR23dfe , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 ,
         \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 ,
         \30685_nR23e00 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 ,
         \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702_nR23e02 , \30703 , \30704 ,
         \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 ,
         \30715 , \30716 , \30717 , \30718 , \30719_nR23e04 , \30720 , \30721 , \30722 , \30723 , \30724 ,
         \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 ,
         \30735 , \30736_nR23e06 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 , \30743 , \30744 ,
         \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753_nR23e08 , \30754 ,
         \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764 ,
         \30765 , \30766 , \30767 , \30768 , \30769 , \30770_nR23e0a , \30771 , \30772 , \30773 , \30774 ,
         \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 ,
         \30785 , \30786 , \30787_nR23e0c , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 ,
         \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 , \30803 , \30804 ,
         \30805_nR23e0e , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 , \30813 , \30814 ,
         \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822_nR23e10 , \30823 , \30824 ,
         \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 , \30833 , \30834 ,
         \30835 , \30836 , \30837 , \30838 , \30839_nR23e14 , \30840 , \30841 , \30842 , \30843 , \30844 ,
         \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 , \30853 , \30854 ,
         \30855 , \30856_nR23e16 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 ,
         \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 , \30873_nR23e18 , \30874 ,
         \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 , \30883 , \30884 ,
         \30885 , \30886 , \30887 , \30888 , \30889 , \30890_nR23e1a , \30891 , \30892 , \30893 , \30894 ,
         \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 , \30903 , \30904 ,
         \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 , \30913 , \30914 ,
         \30915 , \30916_nR23e24 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 , \30923 , \30924 ,
         \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932_nR23e3a , \30933 , \30934 ,
         \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 , \30943 , \30944 ,
         \30945 , \30946 , \30947 , \30948_nR23e50 , \30949 , \30950 , \30951 , \30952 , \30953 , \30954 ,
         \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 ,
         \30965_nR23e66 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 , \30973 , \30974 ,
         \30975 , \30976 , \30977 , \30978 , \30979 , \30980_nR23e7c , \30981 , \30982 , \30983 , \30984 ,
         \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 , \30993 , \30994 ,
         \30995_nR23e92 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 ,
         \31005 , \31006 , \31007 , \31008 , \31009_nR23e9c , \31010 , \31011 , \31012 , \31013 , \31014 ,
         \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023_nR23e9e , \31024 ,
         \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 , \31033 , \31034 ,
         \31035 , \31036 , \31037_nR23ea0 , \31038 , \31039 , \31040 , \31041 , \31042 , \31043 , \31044 ,
         \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052_nR23ea2 , \31053 , \31054 ,
         \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 , \31063 , \31064 ,
         \31065 , \31066_nR23e26 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 ,
         \31075 , \31076 , \31077 , \31078 , \31079 , \31080_nR23e28 , \31081 , \31082 , \31083 , \31084 ,
         \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094_nR23e2a ,
         \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 , \31103 , \31104 ,
         \31105 , \31106 , \31107 , \31108_nR23e2c , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 ,
         \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122_nR23e2e , \31123 , \31124 ,
         \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 ,
         \31135 , \31136_nR23e30 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 , \31143 , \31144 ,
         \31145 , \31146 , \31147 , \31148 , \31149 , \31150_nR23e32 , \31151 , \31152 , \31153 , \31154 ,
         \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 , \31163 , \31164_nR23e34 ,
         \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 ,
         \31175 , \31176 , \31177 , \31178_nR23e36 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 ,
         \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193_nR23e38 , \31194 ,
         \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 ,
         \31205 , \31206 , \31207_nR23e3c , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 ,
         \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221_nR23e3e , \31222 , \31223 , \31224 ,
         \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 ,
         \31235_nR23e40 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 ,
         \31245 , \31246 , \31247 , \31248 , \31249_nR23e42 , \31250 , \31251 , \31252 , \31253 , \31254 ,
         \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 , \31263_nR23e44 , \31264 ,
         \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 ,
         \31275 , \31276 , \31277_nR23e46 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 ,
         \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291_nR23e48 , \31292 , \31293 , \31294 ,
         \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 ,
         \31305_nR23e4a , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 ,
         \31315 , \31316 , \31317 , \31318 , \31319_nR23e4c , \31320 , \31321 , \31322 , \31323 , \31324 ,
         \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333_nR23e4e , \31334 ,
         \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 ,
         \31345 , \31346 , \31347 , \31348_nR23e52 , \31349 , \31350 , \31351 , \31352 , \31353 , \31354 ,
         \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362_nR23e54 , \31363 , \31364 ,
         \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 ,
         \31375 , \31376_nR23e56 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 ,
         \31385 , \31386 , \31387 , \31388 , \31389 , \31390_nR23e58 , \31391 , \31392 , \31393 , \31394 ,
         \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404_nR23e5a ,
         \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 ,
         \31415 , \31416 , \31417 , \31418_nR23e5c , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 ,
         \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432_nR23e5e , \31433 , \31434 ,
         \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 ,
         \31445 , \31446_nR23e60 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 ,
         \31455 , \31456 , \31457 , \31458 , \31459 , \31460_nR23e62 , \31461 , \31462 , \31463 , \31464 ,
         \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474_nR23e64 ,
         \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483 , \31484 ,
         \31485 , \31486 , \31487 , \31488_nR23e68 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 ,
         \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502_nR23e6a , \31503 , \31504 ,
         \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 ,
         \31515 , \31516_nR23e6c , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 ,
         \31525 , \31526 , \31527 , \31528 , \31529 , \31530_nR23e6e , \31531 , \31532 , \31533 , \31534 ,
         \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544_nR23e70 ,
         \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 , \31553 , \31554 ,
         \31555 , \31556 , \31557 , \31558_nR23e72 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 ,
         \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572_nR23e74 , \31573 , \31574 ,
         \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 ,
         \31585 , \31586_nR23e76 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 ,
         \31595 , \31596 , \31597 , \31598 , \31599 , \31600_nR23e78 , \31601 , \31602 , \31603 , \31604 ,
         \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614_nR23e7a ,
         \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 ,
         \31625 , \31626 , \31627 , \31628_nR23e7e , \31629 , \31630 , \31631 , \31632 , \31633 , \31634 ,
         \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642_nR23e80 , \31643 , \31644 ,
         \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 ,
         \31655 , \31656_nR23e82 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 ,
         \31665 , \31666 , \31667 , \31668 , \31669 , \31670_nR23e84 , \31671 , \31672 , \31673 , \31674 ,
         \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 , \31684_nR23e86 ,
         \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 ,
         \31695 , \31696 , \31697 , \31698_nR23e88 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 ,
         \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712_nR23e8a , \31713 , \31714 ,
         \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 ,
         \31725 , \31726_nR23e8c , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 ,
         \31735 , \31736 , \31737 , \31738 , \31739 , \31740_nR23e8e , \31741 , \31742 , \31743 , \31744 ,
         \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 , \31753 , \31754_nR23e90 ,
         \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 ,
         \31765 , \31766 , \31767 , \31768_nR23e94 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 ,
         \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782_nR23e96 , \31783 , \31784 ,
         \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 , \31793 , \31794 ,
         \31795 , \31796_nR23e98 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 ,
         \31805 , \31806 , \31807 , \31808 , \31809 , \31810_nR23e9a , \31811 , \31812 , \31813 , \31814 ,
         \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 ,
         \31825 , \31826 , \31827 , \31828 , \31829_nR23c64 , \31830 , \31831 , \31832 , \31833 , \31834 ,
         \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 ,
         \31845 , \31846_nR23c66 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 ,
         \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862_nR23c68 , \31863 , \31864 ,
         \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 ,
         \31875 , \31876 , \31877 , \31878_nR23c6a , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 ,
         \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894_nR23c6c ,
         \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 ,
         \31905 , \31906 , \31907 , \31908 , \31909 , \31910_nR23c6e , \31911 , \31912 , \31913 , \31914 ,
         \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 , \31923 , \31924 ,
         \31925 , \31926_nR23c70 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 ,
         \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942_nR23c72 , \31943 , \31944 ,
         \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 ,
         \31955 , \31956 , \31957_nR23c74 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 ,
         \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972_nR23c76 , \31973 , \31974 ,
         \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 ,
         \31985 , \31986 , \31987_nR23c78 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 ,
         \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002_nR23c7a , \32003 , \32004 ,
         \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 ,
         \32015 , \32016 , \32017_nR23c7c , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 ,
         \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032_nR23c7e , \32033 , \32034 ,
         \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 ,
         \32045 , \32046 , \32047_nR23c80 , \32048 , \32049 , \32050 , \32051 , \32052 , \32053 , \32054 ,
         \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062_nR23c82 , \32063 , \32064 ,
         \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 ,
         \32075 , \32076 , \32077_nR23c84 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 ,
         \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092_nR23c86 , \32093 , \32094 ,
         \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 ,
         \32105 , \32106 , \32107_nR23c88 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 , \32114 ,
         \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122_nR23c8a , \32123 , \32124 ,
         \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 ,
         \32135 , \32136 , \32137_nR23c8c , \32138 , \32139 , \32140 , \32141 , \32142 , \32143 , \32144 ,
         \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152_nR23c8e , \32153 , \32154 ,
         \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 ,
         \32165 , \32166 , \32167_nR23c90 , \32168 , \32169 , \32170 , \32171 , \32172 , \32173 , \32174 ,
         \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182_nR23c92 , \32183 , \32184 ,
         \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 ,
         \32195 , \32196 , \32197_nR23c94 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 ,
         \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212_nR23c96 , \32213 , \32214 ,
         \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 , \32223 , \32224 ,
         \32225 , \32226 , \32227_nR23c98 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 ,
         \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242_nR23c9a , \32243 , \32244 ,
         \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 ,
         \32255 , \32256 , \32257_nR23c9c , \32258 , \32259 , \32260 , \32261 , \32262 , \32263 , \32264 ,
         \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272_nR23c9e , \32273 , \32274 ,
         \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 ,
         \32285 , \32286 , \32287_nR23ca0 , \32288 , \32289 , \32290 , \32291 , \32292 , \32293 , \32294 ,
         \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302_nR23ca2 , \32303 , \32304 ,
         \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314_nR23ebc ,
         \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 , \32323 , \32324 ,
         \32325_nR23ebe , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 ,
         \32335_nR23ec0 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 , \32343 , \32344 ,
         \32345_nR23ec2 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 ,
         \32355_nR23ec4 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 , \32364 ,
         \32365_nR23ec6 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 , \32373 , \32374 ,
         \32375_nR23ec8 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 ,
         \32385_nR23eca , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 , \32393 , \32394 ,
         \32395_nR23eba , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 ,
         \32405_nR23ecc , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 , \32413 , \32414 ,
         \32415_nR23ece , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 ,
         \32425_nR23ed0 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 , \32433 , \32434 ,
         \32435_nR23ed2 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 ,
         \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 , \32453 , \32454 ,
         \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 , \32463 , \32464 ,
         \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 ,
         \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 ,
         \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 ,
         \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 ,
         \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 , \32513 , \32514 ,
         \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 ,
         \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 ,
         \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 ,
         \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 ,
         \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 ,
         \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 ,
         \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 ,
         \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 , \32594 ,
         \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 ,
         \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 ,
         \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 ,
         \32625 , \32626 , \32627 , \32628 , \32629_nR23eb8 , \32630 , \32631 , \32632 , \32633 , \32634_nR23eea ,
         \32635 , \32636 , \32637 , \32638 , \32639_nR23eec , \32640 , \32641 , \32642 , \32643 , \32644 ,
         \32645 , \32646 , \32647_nR23eee , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 ,
         \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 , \32663 , \32664 ,
         \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 ,
         \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 ,
         \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 ,
         \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704_nR23a0c ,
         \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 ,
         \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 ,
         \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733_nR23a22 , \32734 ,
         \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 ,
         \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753_nR23a38 , \32754 ,
         \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 ,
         \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774_nR23a4e ,
         \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 ,
         \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 , \32793 , \32794 ,
         \32795 , \32796_nR23a64 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 , \32803 , \32804 ,
         \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 , \32813 , \32814 ,
         \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821_nR23a7a , \32822 , \32823 , \32824 ,
         \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 ,
         \32835 , \32836 , \32837 , \32838 , \32839_nR23a84 , \32840 , \32841 , \32842 , \32843 , \32844 ,
         \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 ,
         \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862_nR23a86 , \32863 , \32864 ,
         \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 ,
         \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884_nR23a88 ,
         \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 , \32893 , \32894 ,
         \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 ,
         \32905_nR23a8a , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 ,
         \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924_nR23a0e ,
         \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 , \32933 , \32934 ,
         \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944_nR23a10 ,
         \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 ,
         \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 , \32963_nR23a12 , \32964 ,
         \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 , \32973 , \32974 ,
         \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984_nR23a14 ,
         \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 , \32993 , \32994 ,
         \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004_nR23a16 ,
         \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 , \33013 , \33014 ,
         \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024_nR23a18 ,
         \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 , \33033 , \33034 ,
         \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 , \33043_nR23a1a , \33044 ,
         \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 ,
         \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 , \33063_nR23a1c , \33064 ,
         \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 ,
         \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081_nR23a1e , \33082 , \33083 , \33084 ,
         \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 ,
         \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101_nR23a20 , \33102 , \33103 , \33104 ,
         \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 ,
         \33115 , \33116 , \33117 , \33118 , \33119 , \33120_nR23a24 , \33121 , \33122 , \33123 , \33124 ,
         \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 , \33133 , \33134 ,
         \33135 , \33136 , \33137 , \33138 , \33139_nR23a26 , \33140 , \33141 , \33142 , \33143 , \33144 ,
         \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 , \33153 , \33154 ,
         \33155 , \33156 , \33157 , \33158 , \33159_nR23a28 , \33160 , \33161 , \33162 , \33163 , \33164 ,
         \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 , \33173 , \33174 ,
         \33175 , \33176 , \33177_nR23a2a , \33178 , \33179 , \33180 , \33181 , \33182 , \33183 , \33184 ,
         \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 , \33193 , \33194 ,
         \33195 , \33196 , \33197_nR23a2c , \33198 , \33199 , \33200 , \33201 , \33202 , \33203 , \33204 ,
         \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 ,
         \33215_nR23a2e , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , \33223 , \33224 ,
         \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 ,
         \33235 , \33236_nR23a30 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 , \33243 , \33244 ,
         \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 ,
         \33255_nR23a32 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 , \33263 , \33264 ,
         \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 ,
         \33275_nR23a34 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 , \33283 , \33284 ,
         \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294_nR23a36 ,
         \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 , \33303 , \33304 ,
         \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 ,
         \33315_nR23a3a , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 , \33323 , \33324 ,
         \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334_nR23a3c ,
         \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 , \33343 , \33344 ,
         \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354_nR23a3e ,
         \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 , \33363 , \33364 ,
         \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 , \33373_nR23a40 , \33374 ,
         \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , \33384 ,
         \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392_nR23a42 , \33393 , \33394 ,
         \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , \33403 , \33404 ,
         \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412_nR23a44 , \33413 , \33414 ,
         \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , \33423 , \33424 ,
         \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432_nR23a46 , \33433 , \33434 ,
         \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , \33443 , \33444 ,
         \33445 , \33446 , \33447 , \33448 , \33449 , \33450_nR23a48 , \33451 , \33452 , \33453 , \33454 ,
         \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , \33463 , \33464 ,
         \33465 , \33466 , \33467 , \33468 , \33469_nR23a4a , \33470 , \33471 , \33472 , \33473 , \33474 ,
         \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , \33483 , \33484 ,
         \33485 , \33486 , \33487 , \33488_nR23a4c , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 ,
         \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , \33503 , \33504 ,
         \33505 , \33506 , \33507_nR23a50 , \33508 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 ,
         \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , \33523 , \33524 ,
         \33525 , \33526 , \33527_nR23a52 , \33528 , \33529 , \33530 , \33531 , \33532 , \33533 , \33534 ,
         \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 , \33543 , \33544 ,
         \33545 , \33546 , \33547_nR23a54 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 ,
         \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 ,
         \33565 , \33566_nR23a56 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 , \33573 , \33574 ,
         \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 ,
         \33585 , \33586_nR23a58 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 ,
         \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 , \33603 , \33604_nR23a5a ,
         \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613 , \33614 ,
         \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622_nR23a5c , \33623 , \33624 ,
         \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 , \33633 , \33634 ,
         \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642_nR23a5e , \33643 , \33644 ,
         \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 ,
         \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661_nR23a60 , \33662 , \33663 , \33664 ,
         \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 ,
         \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681_nR23a62 , \33682 , \33683 , \33684 ,
         \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 ,
         \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701_nR23a66 , \33702 , \33703 , \33704 ,
         \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 , \33713 , \33714 ,
         \33715 , \33716 , \33717 , \33718 , \33719_nR23a68 , \33720 , \33721 , \33722 , \33723 , \33724 ,
         \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 ,
         \33735 , \33736 , \33737 , \33738_nR23a6a , \33739 , \33740 , \33741 , \33742 , \33743 , \33744 ,
         \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 ,
         \33755 , \33756_nR23a6c , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 ,
         \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 ,
         \33775 , \33776_nR23a6e , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 ,
         \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 , \33793 , \33794 ,
         \33795 , \33796_nR23a70 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 ,
         \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 ,
         \33815_nR23a72 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 , \33823 , \33824 ,
         \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834_nR23a74 ,
         \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 ,
         \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853_nR23a76 , \33854 ,
         \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 ,
         \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872_nR23a78 , \33873 , \33874 ,
         \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 ,
         \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892_nR23a7c , \33893 , \33894 ,
         \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 , \33903 , \33904 ,
         \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912_nR23a7e , \33913 , \33914 ,
         \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 ,
         \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931_nR23a80 , \33932 , \33933 , \33934 ,
         \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 ,
         \33945 , \33946 , \33947 , \33948 , \33949 , \33950_nR23a82 , \33951 , \33952 , \33953 , \33954 ,
         \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 ,
         \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 ,
         \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 , \33983 , \33984_nR23a8c ,
         \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 ,
         \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004_nR23aa2 ,
         \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 ,
         \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022_nR23ab8 , \34023 , \34024 ,
         \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 ,
         \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042_nR23ace , \34043 , \34044 ,
         \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 , \34053 , \34054 ,
         \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061_nR23ae4 , \34062 , \34063 , \34064 ,
         \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 ,
         \34075 , \34076 , \34077 , \34078 , \34079 , \34080_nR23afa , \34081 , \34082 , \34083 , \34084 ,
         \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 ,
         \34095 , \34096 , \34097 , \34098 , \34099_nR23b04 , \34100 , \34101 , \34102 , \34103 , \34104 ,
         \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 , \34114 ,
         \34115 , \34116 , \34117_nR23b06 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 ,
         \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 ,
         \34135_nR23b08 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 , \34143 , \34144 ,
         \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153_nR23b0a , \34154 ,
         \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 ,
         \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171_nR23a8e , \34172 , \34173 , \34174 ,
         \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 ,
         \34185 , \34186 , \34187 , \34188 , \34189_nR23a90 , \34190 , \34191 , \34192 , \34193 , \34194 ,
         \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 ,
         \34205 , \34206 , \34207_nR23a92 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 ,
         \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 , \34223 , \34224 ,
         \34225_nR23a94 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 ,
         \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243_nR23a96 , \34244 ,
         \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 , \34253 , \34254 ,
         \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261_nR23a98 , \34262 , \34263 , \34264 ,
         \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 ,
         \34275 , \34276 , \34277 , \34278 , \34279_nR23a9a , \34280 , \34281 , \34282 , \34283 , \34284 ,
         \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294 ,
         \34295 , \34296 , \34297_nR23a9c , \34298 , \34299 , \34300 , \34301 , \34302 , \34303 , \34304 ,
         \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 ,
         \34315 , \34316_nR23a9e , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 ,
         \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 , \34333 , \34334 ,
         \34335_nR23aa0 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 ,
         \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353_nR23aa4 , \34354 ,
         \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 ,
         \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371_nR23aa6 , \34372 , \34373 , \34374 ,
         \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 , \34384 ,
         \34385 , \34386 , \34387 , \34388 , \34389_nR23aa8 , \34390 , \34391 , \34392 , \34393 , \34394 ,
         \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 ,
         \34405 , \34406 , \34407_nR23aaa , \34408 , \34409 , \34410 , \34411 , \34412 , \34413 , \34414 ,
         \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 ,
         \34425_nR23aac , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 ,
         \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 , \34443_nR23aae , \34444 ,
         \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 ,
         \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461_nR23ab0 , \34462 , \34463 , \34464 ,
         \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 ,
         \34475 , \34476 , \34477 , \34478 , \34479_nR23ab2 , \34480 , \34481 , \34482 , \34483 , \34484 ,
         \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 , \34493 , \34494 ,
         \34495 , \34496 , \34497_nR23ab4 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 ,
         \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 ,
         \34515_nR23ab6 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 ,
         \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 , \34533_nR23aba , \34534 ,
         \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 ,
         \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551_nR23abc , \34552 , \34553 , \34554 ,
         \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 , \34563 , \34564 ,
         \34565 , \34566 , \34567 , \34568 , \34569_nR23abe , \34570 , \34571 , \34572 , \34573 , \34574 ,
         \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 ,
         \34585 , \34586 , \34587_nR23ac0 , \34588 , \34589 , \34590 , \34591 , \34592 , \34593 , \34594 ,
         \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 ,
         \34605_nR23ac2 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 , \34613 , \34614 ,
         \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623_nR23ac4 , \34624 ,
         \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 , \34634 ,
         \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641_nR23ac6 , \34642 , \34643 , \34644 ,
         \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 ,
         \34655 , \34656 , \34657 , \34658 , \34659_nR23ac8 , \34660 , \34661 , \34662 , \34663 , \34664 ,
         \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 ,
         \34675 , \34676 , \34677 , \34678_nR23aca , \34679 , \34680 , \34681 , \34682 , \34683 , \34684 ,
         \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 ,
         \34695 , \34696_nR23acc , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 , \34703 , \34704 ,
         \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 ,
         \34715_nR23ad0 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 , \34723 , \34724 ,
         \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 , \34733_nR23ad2 , \34734 ,
         \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 ,
         \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751_nR23ad4 , \34752 , \34753 , \34754 ,
         \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 ,
         \34765 , \34766 , \34767 , \34768 , \34769_nR23ad6 , \34770 , \34771 , \34772 , \34773 , \34774 ,
         \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 , \34783 , \34784 ,
         \34785 , \34786 , \34787_nR23ad8 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 ,
         \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 ,
         \34805_nR23ada , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 , \34813 , \34814 ,
         \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823_nR23adc , \34824 ,
         \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 ,
         \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841_nR23ade , \34842 , \34843 , \34844 ,
         \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 ,
         \34855 , \34856 , \34857 , \34858 , \34859_nR23ae0 , \34860 , \34861 , \34862 , \34863 , \34864 ,
         \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 ,
         \34875 , \34876 , \34877_nR23ae2 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 ,
         \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 , \34893 , \34894 ,
         \34895_nR23ae6 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 ,
         \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913_nR23ae8 , \34914 ,
         \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 , \34923 , \34924 ,
         \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933_nR23aea , \34934 ,
         \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 ,
         \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951_nR23aec , \34952 , \34953 , \34954 ,
         \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 ,
         \34965 , \34966 , \34967 , \34968 , \34969_nR23aee , \34970 , \34971 , \34972 , \34973 , \34974 ,
         \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 ,
         \34985 , \34986 , \34987_nR23af0 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 ,
         \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 , \35003 , \35004 ,
         \35005_nR23af2 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 ,
         \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023_nR23af4 , \35024 ,
         \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 ,
         \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041_nR23af6 , \35042 , \35043 , \35044 ,
         \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 , \35053 , \35054 ,
         \35055 , \35056 , \35057 , \35058 , \35059_nR23af8 , \35060 , \35061 , \35062 , \35063 , \35064 ,
         \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 ,
         \35075 , \35076 , \35077_nR23afc , \35078 , \35079 , \35080 , \35081 , \35082 , \35083 , \35084 ,
         \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094 ,
         \35095_nR23afe , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 ,
         \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 , \35113_nR23b00 , \35114 ,
         \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 ,
         \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131_nR23b02 , \35132 , \35133 , \35134 ,
         \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 ,
         \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 ,
         \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 , \35163 , \35164_nR23b0c ,
         \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 ,
         \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182_nR23b22 , \35183 , \35184 ,
         \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 ,
         \35195 , \35196 , \35197 , \35198 , \35199 , \35200_nR23b38 , \35201 , \35202 , \35203 , \35204 ,
         \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 ,
         \35215 , \35216 , \35217 , \35218_nR23b4e , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 ,
         \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 , \35233 , \35234 ,
         \35235 , \35236_nR23b64 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 , \35243 , \35244 ,
         \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 ,
         \35255 , \35256_nR23b7a , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 , \35263 , \35264 ,
         \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272_nR23b84 , \35273 , \35274 ,
         \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 , \35283 , \35284 ,
         \35285 , \35286 , \35287 , \35288 , \35289_nR23b86 , \35290 , \35291 , \35292 , \35293 , \35294 ,
         \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 , \35303 , \35304 ,
         \35305 , \35306_nR23b88 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 ,
         \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 ,
         \35325_nR23b8a , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 , \35333 , \35334 ,
         \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342_nR23b0e , \35343 , \35344 ,
         \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 , \35353 , \35354 ,
         \35355 , \35356 , \35357 , \35358 , \35359_nR23b10 , \35360 , \35361 , \35362 , \35363 , \35364 ,
         \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 , \35373 , \35374 ,
         \35375 , \35376 , \35377_nR23b12 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 ,
         \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 , \35393 , \35394_nR23b14 ,
         \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 , \35403 , \35404 ,
         \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411_nR23b16 , \35412 , \35413 , \35414 ,
         \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 , \35423 , \35424 ,
         \35425 , \35426 , \35427 , \35428_nR23b18 , \35429 , \35430 , \35431 , \35432 , \35433 , \35434 ,
         \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 , \35443 , \35444 ,
         \35445_nR23b1a , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 , \35453 , \35454 ,
         \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462_nR23b1c , \35463 , \35464 ,
         \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 , \35473 , \35474 ,
         \35475 , \35476 , \35477 , \35478 , \35479_nR23b1e , \35480 , \35481 , \35482 , \35483 , \35484 ,
         \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , \35494 ,
         \35495 , \35496_nR23b20 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 ,
         \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513_nR23b24 , \35514 ,
         \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 , \35523 , \35524 ,
         \35525 , \35526 , \35527 , \35528 , \35529 , \35530_nR23b26 , \35531 , \35532 , \35533 , \35534 ,
         \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 , \35543 , \35544 ,
         \35545 , \35546 , \35547 , \35548_nR23b28 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 ,
         \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 , \35563 , \35564 ,
         \35565_nR23b2a , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 , \35573 , \35574 ,
         \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582_nR23b2c , \35583 , \35584 ,
         \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 ,
         \35595 , \35596 , \35597 , \35598 , \35599_nR23b2e , \35600 , \35601 , \35602 , \35603 , \35604 ,
         \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 ,
         \35615 , \35616_nR23b30 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 , \35623 , \35624 ,
         \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633_nR23b32 , \35634 ,
         \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 , \35643 , \35644 ,
         \35645 , \35646 , \35647 , \35648 , \35649 , \35650_nR23b34 , \35651 , \35652 , \35653 , \35654 ,
         \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , \35663 , \35664 ,
         \35665 , \35666 , \35667_nR23b36 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 ,
         \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , \35683 , \35684_nR23b3a ,
         \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 ,
         \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701_nR23b3c , \35702 , \35703 , \35704 ,
         \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 , \35713 , \35714 ,
         \35715 , \35716 , \35717 , \35718_nR23b3e , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 ,
         \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 , \35733 , \35734 ,
         \35735_nR23b40 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 ,
         \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752_nR23b42 , \35753 , \35754 ,
         \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 ,
         \35765 , \35766 , \35767 , \35768 , \35769_nR23b44 , \35770 , \35771 , \35772 , \35773 , \35774 ,
         \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 ,
         \35785 , \35786_nR23b46 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 , \35793 , \35794 ,
         \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 , \35803_nR23b48 , \35804 ,
         \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 , \35813 , \35814 ,
         \35815 , \35816 , \35817 , \35818 , \35819 , \35820_nR23b4a , \35821 , \35822 , \35823 , \35824 ,
         \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 , \35833 , \35834 ,
         \35835 , \35836 , \35837_nR23b4c , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 ,
         \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854_nR23b50 ,
         \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 , \35863 , \35864 ,
         \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871_nR23b52 , \35872 , \35873 , \35874 ,
         \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 ,
         \35885 , \35886 , \35887 , \35888_nR23b54 , \35889 , \35890 , \35891 , \35892 , \35893 , \35894 ,
         \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 ,
         \35905_nR23b56 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 ,
         \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922_nR23b58 , \35923 , \35924 ,
         \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 ,
         \35935 , \35936 , \35937 , \35938 , \35939_nR23b5a , \35940 , \35941 , \35942 , \35943 , \35944 ,
         \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 ,
         \35955 , \35956_nR23b5c , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 ,
         \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 , \35973_nR23b5e , \35974 ,
         \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 ,
         \35985 , \35986 , \35987 , \35988 , \35989 , \35990_nR23b60 , \35991 , \35992 , \35993 , \35994 ,
         \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 ,
         \36005 , \36006 , \36007_nR23b62 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 ,
         \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 , \36024_nR23b66 ,
         \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 ,
         \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041_nR23b68 , \36042 , \36043 , \36044 ,
         \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 , \36053 , \36054 ,
         \36055 , \36056 , \36057 , \36058_nR23b6a , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 ,
         \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 ,
         \36075_nR23b6c , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 , \36083 , \36084 ,
         \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092_nR23b6e , \36093 , \36094 ,
         \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 ,
         \36105 , \36106 , \36107 , \36108 , \36109_nR23b70 , \36110 , \36111 , \36112 , \36113 , \36114 ,
         \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 ,
         \36125 , \36126_nR23b72 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 , \36133 , \36134 ,
         \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143_nR23b74 , \36144 ,
         \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 ,
         \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161_nR23b76 , \36162 , \36163 , \36164 ,
         \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 , \36173 , \36174 ,
         \36175 , \36176 , \36177 , \36178_nR23b78 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 ,
         \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 ,
         \36195_nR23b7c , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 ,
         \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212_nR23b7e , \36213 , \36214 ,
         \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 ,
         \36225 , \36226 , \36227 , \36228 , \36229_nR23b80 , \36230 , \36231 , \36232 , \36233 , \36234 ,
         \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 , \36243 , \36244 ,
         \36245 , \36246_nR23b82 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 ,
         \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 ,
         \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 , \36273_nR23b8c , \36274 ,
         \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 ,
         \36285 , \36286 , \36287 , \36288 , \36289_nR23ba2 , \36290 , \36291 , \36292 , \36293 , \36294 ,
         \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 , \36303 , \36304 ,
         \36305_nR23bb8 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 ,
         \36315 , \36316 , \36317 , \36318 , \36319 , \36320_nR23bce , \36321 , \36322 , \36323 , \36324 ,
         \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36334 ,
         \36335_nR23be4 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 , \36343 , \36344 ,
         \36345 , \36346 , \36347 , \36348 , \36349 , \36350_nR23bfa , \36351 , \36352 , \36353 , \36354 ,
         \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364_nR23c04 ,
         \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 , \36373 , \36374 ,
         \36375 , \36376 , \36377 , \36378 , \36379_nR23c06 , \36380 , \36381 , \36382 , \36383 , \36384 ,
         \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393_nR23c08 , \36394 ,
         \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 , \36403 , \36404 ,
         \36405 , \36406 , \36407 , \36408_nR23c0a , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 ,
         \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422_nR23b8e , \36423 , \36424 ,
         \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 ,
         \36435 , \36436_nR23b90 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 ,
         \36445 , \36446 , \36447 , \36448 , \36449 , \36450_nR23b92 , \36451 , \36452 , \36453 , \36454 ,
         \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464_nR23b94 ,
         \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 ,
         \36475 , \36476 , \36477 , \36478_nR23b96 , \36479 , \36480 , \36481 , \36482 , \36483 , \36484 ,
         \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492_nR23b98 , \36493 , \36494 ,
         \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 ,
         \36505 , \36506_nR23b9a , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 , \36513 , \36514 ,
         \36515 , \36516 , \36517 , \36518 , \36519 , \36520_nR23b9c , \36521 , \36522 , \36523 , \36524 ,
         \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534_nR23b9e ,
         \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 ,
         \36545 , \36546 , \36547 , \36548 , \36549_nR23ba0 , \36550 , \36551 , \36552 , \36553 , \36554 ,
         \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 , \36563_nR23ba4 , \36564 ,
         \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 ,
         \36575 , \36576 , \36577_nR23ba6 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 ,
         \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591_nR23ba8 , \36592 , \36593 , \36594 ,
         \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 ,
         \36605_nR23baa , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 ,
         \36615 , \36616 , \36617 , \36618 , \36619_nR23bac , \36620 , \36621 , \36622 , \36623 , \36624 ,
         \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633_nR23bae , \36634 ,
         \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 , \36643 , \36644 ,
         \36645 , \36646 , \36647_nR23bb0 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 ,
         \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661_nR23bb2 , \36662 , \36663 , \36664 ,
         \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 , \36673 , \36674 ,
         \36675_nR23bb4 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 ,
         \36685 , \36686 , \36687 , \36688 , \36689_nR23bb6 , \36690 , \36691 , \36692 , \36693 , \36694 ,
         \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704_nR23bba ,
         \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 ,
         \36715 , \36716 , \36717 , \36718_nR23bbc , \36719 , \36720 , \36721 , \36722 , \36723 , \36724 ,
         \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732_nR23bbe , \36733 , \36734 ,
         \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 ,
         \36745 , \36746_nR23bc0 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 , \36753 , \36754 ,
         \36755 , \36756 , \36757 , \36758 , \36759 , \36760_nR23bc2 , \36761 , \36762 , \36763 , \36764 ,
         \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774_nR23bc4 ,
         \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 , \36783 , \36784 ,
         \36785 , \36786 , \36787 , \36788_nR23bc6 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 ,
         \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802_nR23bc8 , \36803 , \36804 ,
         \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 , \36814 ,
         \36815 , \36816_nR23bca , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 ,
         \36825 , \36826 , \36827 , \36828 , \36829 , \36830_nR23bcc , \36831 , \36832 , \36833 , \36834 ,
         \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844_nR23bd0 ,
         \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 , \36853 , \36854 ,
         \36855 , \36856 , \36857 , \36858_nR23bd2 , \36859 , \36860 , \36861 , \36862 , \36863 , \36864 ,
         \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872_nR23bd4 , \36873 , \36874 ,
         \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 , \36883 , \36884 ,
         \36885 , \36886_nR23bd6 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 ,
         \36895 , \36896 , \36897 , \36898 , \36899 , \36900_nR23bd8 , \36901 , \36902 , \36903 , \36904 ,
         \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914_nR23bda ,
         \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 , \36923 , \36924 ,
         \36925 , \36926 , \36927 , \36928_nR23bdc , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 ,
         \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942_nR23bde , \36943 , \36944 ,
         \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 ,
         \36955 , \36956_nR23be0 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 , \36964 ,
         \36965 , \36966 , \36967 , \36968 , \36969 , \36970_nR23be2 , \36971 , \36972 , \36973 , \36974 ,
         \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984_nR23be6 ,
         \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 , \36993 , \36994 ,
         \36995 , \36996 , \36997 , \36998_nR23be8 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 ,
         \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012_nR23bea , \37013 , \37014 ,
         \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 ,
         \37025 , \37026_nR23bec , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 ,
         \37035 , \37036 , \37037 , \37038 , \37039 , \37040_nR23bee , \37041 , \37042 , \37043 , \37044 ,
         \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054_nR23bf0 ,
         \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 ,
         \37065 , \37066 , \37067 , \37068_nR23bf2 , \37069 , \37070 , \37071 , \37072 , \37073 , \37074 ,
         \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082_nR23bf4 , \37083 , \37084 ,
         \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 ,
         \37095 , \37096_nR23bf6 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 ,
         \37105 , \37106 , \37107 , \37108 , \37109 , \37110_nR23bf8 , \37111 , \37112 , \37113 , \37114 ,
         \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 , \37123 , \37124_nR23bfc ,
         \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 ,
         \37135 , \37136 , \37137 , \37138_nR23bfe , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 ,
         \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152_nR23c00 , \37153 , \37154 ,
         \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 ,
         \37165 , \37166_nR23c02 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 ,
         \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 ,
         \37185_nR239cc , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 ,
         \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203_nR239ce , \37204 ,
         \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 ,
         \37215 , \37216 , \37217 , \37218 , \37219_nR239d0 , \37220 , \37221 , \37222 , \37223 , \37224 ,
         \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 , \37233 , \37234 ,
         \37235 , \37236_nR239d2 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 ,
         \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 , \37253_nR239d4 , \37254 ,
         \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 , \37263 , \37264 ,
         \37265 , \37266 , \37267 , \37268 , \37269 , \37270_nR239d6 , \37271 , \37272 , \37273 , \37274 ,
         \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 ,
         \37285 , \37286 , \37287_nR239d8 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 ,
         \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304_nR239da ,
         \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 , \37313 , \37314 ,
         \37315 , \37316 , \37317 , \37318 , \37319_nR239dc , \37320 , \37321 , \37322 , \37323 , \37324 ,
         \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334_nR239de ,
         \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 , \37343 , \37344 ,
         \37345 , \37346 , \37347 , \37348 , \37349_nR239e0 , \37350 , \37351 , \37352 , \37353 , \37354 ,
         \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364_nR239e2 ,
         \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 ,
         \37375 , \37376 , \37377 , \37378 , \37379_nR239e4 , \37380 , \37381 , \37382 , \37383 , \37384 ,
         \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 , \37393 , \37394_nR239e6 ,
         \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 ,
         \37405 , \37406 , \37407 , \37408 , \37409_nR239e8 , \37410 , \37411 , \37412 , \37413 , \37414 ,
         \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 , \37423 , \37424_nR239ea ,
         \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 ,
         \37435 , \37436 , \37437 , \37438 , \37439_nR239ec , \37440 , \37441 , \37442 , \37443 , \37444 ,
         \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 , \37453 , \37454_nR239ee ,
         \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 ,
         \37465 , \37466 , \37467 , \37468 , \37469_nR239f0 , \37470 , \37471 , \37472 , \37473 , \37474 ,
         \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 , \37483 , \37484_nR239f2 ,
         \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 ,
         \37495 , \37496 , \37497 , \37498 , \37499_nR239f4 , \37500 , \37501 , \37502 , \37503 , \37504 ,
         \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37514_nR239f6 ,
         \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 , \37523 , \37524 ,
         \37525 , \37526 , \37527 , \37528 , \37529_nR239f8 , \37530 , \37531 , \37532 , \37533 , \37534 ,
         \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544_nR239fa ,
         \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 , \37553 , \37554 ,
         \37555 , \37556 , \37557 , \37558 , \37559_nR239fc , \37560 , \37561 , \37562 , \37563 , \37564 ,
         \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 , \37573 , \37574_nR239fe ,
         \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 ,
         \37585 , \37586 , \37587 , \37588 , \37589_nR23a00 , \37590 , \37591 , \37592 , \37593 , \37594 ,
         \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604_nR23a02 ,
         \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 , \37613 , \37614 ,
         \37615 , \37616 , \37617 , \37618 , \37619_nR23a04 , \37620 , \37621 , \37622 , \37623 , \37624 ,
         \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 , \37633 , \37634_nR23a06 ,
         \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 ,
         \37645 , \37646 , \37647 , \37648 , \37649_nR23a08 , \37650 , \37651 , \37652 , \37653 , \37654 ,
         \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 , \37663 , \37664_nR23a0a ,
         \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 ,
         \37675 , \37676_nR23c24 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 , \37683 , \37684 ,
         \37685 , \37686 , \37687_nR23c26 , \37688 , \37689 , \37690 , \37691 , \37692 , \37693 , \37694 ,
         \37695 , \37696 , \37697_nR23c28 , \37698 , \37699 , \37700 , \37701 , \37702 , \37703 , \37704 ,
         \37705 , \37706 , \37707_nR23c2a , \37708 , \37709 , \37710 , \37711 , \37712 , \37713 , \37714 ,
         \37715 , \37716 , \37717_nR23c2c , \37718 , \37719 , \37720 , \37721 , \37722 , \37723 , \37724 ,
         \37725 , \37726 , \37727_nR23c2e , \37728 , \37729 , \37730 , \37731 , \37732 , \37733 , \37734 ,
         \37735 , \37736 , \37737_nR23c30 , \37738 , \37739 , \37740 , \37741 , \37742 , \37743 , \37744 ,
         \37745 , \37746 , \37747_nR23c32 , \37748 , \37749 , \37750 , \37751 , \37752 , \37753 , \37754 ,
         \37755 , \37756 , \37757_nR23c22 , \37758 , \37759 , \37760 , \37761 , \37762 , \37763 , \37764 ,
         \37765 , \37766 , \37767_nR23c34 , \37768 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 ,
         \37775 , \37776 , \37777_nR23c36 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 ,
         \37785 , \37786 , \37787_nR23c38 , \37788 , \37789 , \37790 , \37791 , \37792 , \37793 , \37794 ,
         \37795 , \37796 , \37797_nR23c3a , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 ,
         \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 , \37813 , \37814 ,
         \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 ,
         \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 , \37833 , \37834 ,
         \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 ,
         \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 , \37853 , \37854 ,
         \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 ,
         \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 , \37873 , \37874 ,
         \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 ,
         \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 , \37894 ,
         \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 , \37903 , \37904 ,
         \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 ,
         \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 , \37923 , \37924 ,
         \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 ,
         \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 , \37943 , \37944 ,
         \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 ,
         \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 , \37963 , \37964 ,
         \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974 ,
         \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 , \37983 , \37984 ,
         \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 ,
         \37995 , \37996 , \37997_nR23c20 , \37998 , \37999 , \38000 , \38001 , \38002_nR23c52 , \38003 , \38004 ,
         \38005 , \38006 , \38007_nR23c54 , \38008 , \38009 , \38010 , \38011 , \38012_nR23c56 , \38013 , \38014 ,
         \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 ,
         \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 , \38033 , \38034 ,
         \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 ,
         \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 , \38053 , \38054 ,
         \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 ,
         \38065 , \38066 , \38067 , \38068_nR23774 , \38069 , \38070 , \38071 , \38072 , \38073 , \38074 ,
         \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 ,
         \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 , \38093 , \38094 ,
         \38095 , \38096_nR2378a , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 ,
         \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 ,
         \38115_nR237a0 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 , \38123 , \38124 ,
         \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 , \38133 , \38134 ,
         \38135 , \38136_nR237b6 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 ,
         \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 ,
         \38155_nR237cc , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 , \38164 ,
         \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 , \38173 , \38174 ,
         \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181_nR237e2 , \38182 , \38183 , \38184 ,
         \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 ,
         \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201_nR237ec , \38202 , \38203 , \38204 ,
         \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 ,
         \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221_nR237ee , \38222 , \38223 , \38224 ,
         \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 ,
         \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241_nR237f0 , \38242 , \38243 , \38244 ,
         \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 , \38253 , \38254 ,
         \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261_nR237f2 , \38262 , \38263 , \38264 ,
         \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 ,
         \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281_nR23776 , \38282 , \38283 , \38284 ,
         \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 ,
         \38295 , \38296 , \38297 , \38298 , \38299 , \38300_nR23778 , \38301 , \38302 , \38303 , \38304 ,
         \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 ,
         \38315 , \38316 , \38317 , \38318 , \38319_nR2377a , \38320 , \38321 , \38322 , \38323 , \38324 ,
         \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 , \38333 , \38334 ,
         \38335 , \38336 , \38337 , \38338 , \38339_nR2377c , \38340 , \38341 , \38342 , \38343 , \38344 ,
         \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 ,
         \38355 , \38356 , \38357 , \38358 , \38359_nR2377e , \38360 , \38361 , \38362 , \38363 , \38364 ,
         \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 ,
         \38375 , \38376 , \38377 , \38378_nR23780 , \38379 , \38380 , \38381 , \38382 , \38383 , \38384 ,
         \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 ,
         \38395 , \38396 , \38397_nR23782 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 ,
         \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 , \38413 , \38414 ,
         \38415 , \38416 , \38417_nR23784 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 ,
         \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 ,
         \38435_nR23786 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 , \38443 , \38444 ,
         \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453_nR23788 , \38454 ,
         \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 ,
         \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472_nR2378c , \38473 , \38474 ,
         \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 ,
         \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491_nR2378e , \38492 , \38493 , \38494 ,
         \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 ,
         \38505 , \38506 , \38507 , \38508 , \38509 , \38510_nR23790 , \38511 , \38512 , \38513 , \38514 ,
         \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 , \38523 , \38524 ,
         \38525 , \38526 , \38527 , \38528_nR23792 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 ,
         \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 ,
         \38545 , \38546 , \38547_nR23794 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 ,
         \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 ,
         \38565_nR23796 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 , \38573 , \38574 ,
         \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583_nR23798 , \38584 ,
         \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 ,
         \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601_nR2379a , \38602 , \38603 , \38604 ,
         \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 , \38613 , \38614 ,
         \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622_nR2379c , \38623 , \38624 ,
         \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 ,
         \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 , \38643_nR2379e , \38644 ,
         \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 , \38653 , \38654 ,
         \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663_nR237a2 , \38664 ,
         \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 ,
         \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 , \38683_nR237a4 , \38684 ,
         \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 ,
         \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703_nR237a6 , \38704 ,
         \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 ,
         \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723_nR237a8 , \38724 ,
         \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 , \38733 , \38734 ,
         \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744_nR237aa ,
         \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 ,
         \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 , \38763 , \38764_nR237ac ,
         \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 ,
         \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783_nR237ae , \38784 ,
         \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 ,
         \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802_nR237b0 , \38803 , \38804 ,
         \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 , \38814 ,
         \38815 , \38816 , \38817 , \38818 , \38819 , \38820_nR237b2 , \38821 , \38822 , \38823 , \38824 ,
         \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 ,
         \38835 , \38836 , \38837 , \38838 , \38839_nR237b4 , \38840 , \38841 , \38842 , \38843 , \38844 ,
         \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 ,
         \38855 , \38856 , \38857_nR237b8 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 ,
         \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 , \38873 , \38874 ,
         \38875_nR237ba , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 ,
         \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893_nR237bc , \38894 ,
         \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 ,
         \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912_nR237be , \38913 , \38914 ,
         \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 , \38923 , \38924 ,
         \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931_nR237c0 , \38932 , \38933 , \38934 ,
         \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 ,
         \38945 , \38946 , \38947 , \38948 , \38949 , \38950_nR237c2 , \38951 , \38952 , \38953 , \38954 ,
         \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 ,
         \38965 , \38966 , \38967 , \38968_nR237c4 , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 ,
         \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 ,
         \38985 , \38986 , \38987_nR237c6 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 ,
         \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 , \39003 , \39004 ,
         \39005_nR237c8 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 ,
         \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024_nR237ca ,
         \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 , \39033 , \39034 ,
         \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043_nR237ce , \39044 ,
         \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 ,
         \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064_nR237d0 ,
         \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 ,
         \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 , \39084_nR237d2 ,
         \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 ,
         \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103_nR237d4 , \39104 ,
         \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 ,
         \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122_nR237d6 , \39123 , \39124 ,
         \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 ,
         \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141_nR237d8 , \39142 , \39143 , \39144 ,
         \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 , \39153 , \39154 ,
         \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161_nR237da , \39162 , \39163 , \39164 ,
         \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 ,
         \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181_nR237dc , \39182 , \39183 , \39184 ,
         \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 ,
         \39195 , \39196 , \39197 , \39198 , \39199 , \39200_nR237de , \39201 , \39202 , \39203 , \39204 ,
         \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 , \39213 , \39214 ,
         \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221_nR237e0 , \39222 , \39223 , \39224 ,
         \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 , \39233 , \39234 ,
         \39235 , \39236 , \39237 , \39238 , \39239 , \39240_nR237e4 , \39241 , \39242 , \39243 , \39244 ,
         \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 , \39253 , \39254 ,
         \39255 , \39256 , \39257 , \39258 , \39259 , \39260_nR237e6 , \39261 , \39262 , \39263 , \39264 ,
         \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 , \39273 , \39274 ,
         \39275 , \39276 , \39277 , \39278 , \39279_nR237e8 , \39280 , \39281 , \39282 , \39283 , \39284 ,
         \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 , \39293 , \39294 ,
         \39295 , \39296 , \39297 , \39298_nR237ea , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 ,
         \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 , \39314 ,
         \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 , \39323 , \39324 ,
         \39325 , \39326 , \39327 , \39328 , \39329 , \39330_nR237f4 , \39331 , \39332 , \39333 , \39334 ,
         \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 ,
         \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351_nR2380a , \39352 , \39353 , \39354 ,
         \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 ,
         \39365 , \39366 , \39367 , \39368 , \39369 , \39370_nR23820 , \39371 , \39372 , \39373 , \39374 ,
         \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 ,
         \39385 , \39386 , \39387 , \39388 , \39389 , \39390_nR23836 , \39391 , \39392 , \39393 , \39394 ,
         \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 , \39403 , \39404 ,
         \39405 , \39406 , \39407 , \39408 , \39409_nR2384c , \39410 , \39411 , \39412 , \39413 , \39414 ,
         \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 ,
         \39425 , \39426 , \39427 , \39428_nR23862 , \39429 , \39430 , \39431 , \39432 , \39433 , \39434 ,
         \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 ,
         \39445 , \39446 , \39447_nR2386c , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 ,
         \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 ,
         \39465_nR2386e , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 ,
         \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 , \39483_nR23870 , \39484 ,
         \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 ,
         \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501_nR23872 , \39502 , \39503 , \39504 ,
         \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 , \39513 , \39514 ,
         \39515 , \39516 , \39517 , \39518 , \39519 , \39520_nR237f6 , \39521 , \39522 , \39523 , \39524 ,
         \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 ,
         \39535 , \39536 , \39537 , \39538_nR237f8 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 ,
         \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 ,
         \39555 , \39556_nR237fa , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 , \39564 ,
         \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574_nR237fc ,
         \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 ,
         \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592_nR237fe , \39593 , \39594 ,
         \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 ,
         \39605 , \39606 , \39607 , \39608 , \39609 , \39610_nR23800 , \39611 , \39612 , \39613 , \39614 ,
         \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 , \39623 , \39624 ,
         \39625 , \39626 , \39627 , \39628_nR23802 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 ,
         \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 ,
         \39645 , \39646_nR23804 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 ,
         \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664_nR23806 ,
         \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 , \39673 , \39674 ,
         \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682_nR23808 , \39683 , \39684 ,
         \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 ,
         \39695 , \39696 , \39697 , \39698 , \39699 , \39700_nR2380c , \39701 , \39702 , \39703 , \39704 ,
         \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 ,
         \39715 , \39716 , \39717 , \39718_nR2380e , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 ,
         \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 ,
         \39735 , \39736_nR23810 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 ,
         \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 , \39753 , \39754_nR23812 ,
         \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 ,
         \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772_nR23814 , \39773 , \39774 ,
         \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 ,
         \39785 , \39786 , \39787 , \39788 , \39789 , \39790_nR23816 , \39791 , \39792 , \39793 , \39794 ,
         \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 ,
         \39805 , \39806 , \39807 , \39808_nR23818 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 ,
         \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 , \39823 , \39824 ,
         \39825 , \39826_nR2381a , \39827 , \39828 , \39829 , \39830 , \39831 , \39832 , \39833 , \39834 ,
         \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844_nR2381c ,
         \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852 , \39853 , \39854 ,
         \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862_nR2381e , \39863 , \39864 ,
         \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 , \39873 , \39874 ,
         \39875 , \39876 , \39877 , \39878 , \39879 , \39880_nR23822 , \39881 , \39882 , \39883 , \39884 ,
         \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 ,
         \39895 , \39896 , \39897 , \39898_nR23824 , \39899 , \39900 , \39901 , \39902 , \39903 , \39904 ,
         \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 ,
         \39915 , \39916_nR23826 , \39917 , \39918 , \39919 , \39920 , \39921 , \39922 , \39923 , \39924 ,
         \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934_nR23828 ,
         \39935 , \39936 , \39937 , \39938 , \39939 , \39940 , \39941 , \39942 , \39943 , \39944 ,
         \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952_nR2382a , \39953 , \39954 ,
         \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962 , \39963 , \39964 ,
         \39965 , \39966 , \39967 , \39968 , \39969 , \39970_nR2382c , \39971 , \39972 , \39973 , \39974 ,
         \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 , \39983 , \39984 ,
         \39985 , \39986 , \39987 , \39988_nR2382e , \39989 , \39990 , \39991 , \39992 , \39993 , \39994 ,
         \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002 , \40003 , \40004 ,
         \40005 , \40006_nR23830 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 , \40013 , \40014 ,
         \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 , \40023 , \40024 ,
         \40025_nR23832 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 , \40033 , \40034 ,
         \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 , \40043_nR23834 , \40044 ,
         \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 , \40053 , \40054 ,
         \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061_nR23838 , \40062 , \40063 , \40064 ,
         \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 , \40073 , \40074 ,
         \40075 , \40076 , \40077 , \40078 , \40079_nR2383a , \40080 , \40081 , \40082 , \40083 , \40084 ,
         \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 , \40093 , \40094 ,
         \40095 , \40096 , \40097_nR2383c , \40098 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 ,
         \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 ,
         \40115_nR2383e , \40116 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 , \40123 , \40124 ,
         \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133_nR23840 , \40134 ,
         \40135 , \40136 , \40137 , \40138 , \40139 , \40140 , \40141 , \40142 , \40143 , \40144 ,
         \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151_nR23842 , \40152 , \40153 , \40154 ,
         \40155 , \40156 , \40157 , \40158 , \40159 , \40160 , \40161 , \40162 , \40163 , \40164 ,
         \40165 , \40166 , \40167 , \40168 , \40169_nR23844 , \40170 , \40171 , \40172 , \40173 , \40174 ,
         \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182 , \40183 , \40184 ,
         \40185 , \40186 , \40187_nR23846 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 ,
         \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 , \40203 , \40204 ,
         \40205_nR23848 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 ,
         \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223_nR2384a , \40224 ,
         \40225 , \40226 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 , \40233 , \40234 ,
         \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241_nR2384e , \40242 , \40243 , \40244 ,
         \40245 , \40246 , \40247 , \40248 , \40249 , \40250 , \40251 , \40252 , \40253 , \40254 ,
         \40255 , \40256 , \40257 , \40258 , \40259_nR23850 , \40260 , \40261 , \40262 , \40263 , \40264 ,
         \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271 , \40272 , \40273 , \40274 ,
         \40275 , \40276 , \40277 , \40278_nR23852 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 ,
         \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 , \40293 , \40294 ,
         \40295 , \40296_nR23854 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 ,
         \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 , \40314_nR23856 ,
         \40315 , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 , \40323 , \40324 ,
         \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332_nR23858 , \40333 , \40334 ,
         \40335 , \40336 , \40337 , \40338 , \40339 , \40340 , \40341 , \40342 , \40343 , \40344 ,
         \40345 , \40346 , \40347 , \40348 , \40349 , \40350_nR2385a , \40351 , \40352 , \40353 , \40354 ,
         \40355 , \40356 , \40357 , \40358 , \40359 , \40360 , \40361 , \40362 , \40363 , \40364 ,
         \40365 , \40366 , \40367 , \40368_nR2385c , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 ,
         \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381 , \40382 , \40383 , \40384 ,
         \40385 , \40386_nR2385e , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 ,
         \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 , \40403 , \40404_nR23860 ,
         \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411 , \40412 , \40413 , \40414 ,
         \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422_nR23864 , \40423 , \40424 ,
         \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 ,
         \40435 , \40436 , \40437 , \40438 , \40439 , \40440_nR23866 , \40441 , \40442 , \40443 , \40444 ,
         \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 , \40453 , \40454 ,
         \40455 , \40456 , \40457 , \40458_nR23868 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 ,
         \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 ,
         \40475 , \40476_nR2386a , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 , \40483 , \40484 ,
         \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 ,
         \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 ,
         \40505 , \40506 , \40507_nR23874 , \40508 , \40509 , \40510 , \40511 , \40512 , \40513 , \40514 ,
         \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 ,
         \40525 , \40526 , \40527_nR2388a , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 ,
         \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 , \40543 , \40544 ,
         \40545_nR238a0 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 ,
         \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563_nR238b6 , \40564 ,
         \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 ,
         \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581_nR238cc , \40582 , \40583 , \40584 ,
         \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 , \40594 ,
         \40595 , \40596 , \40597 , \40598 , \40599_nR238e2 , \40600 , \40601 , \40602 , \40603 , \40604 ,
         \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 ,
         \40615 , \40616_nR238ec , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 , \40623 , \40624 ,
         \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633_nR238ee , \40634 ,
         \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 ,
         \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651_nR238f0 , \40652 , \40653 , \40654 ,
         \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 ,
         \40665 , \40666 , \40667 , \40668 , \40669_nR238f2 , \40670 , \40671 , \40672 , \40673 , \40674 ,
         \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 , \40683 , \40684 ,
         \40685 , \40686 , \40687 , \40688_nR23876 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 ,
         \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 ,
         \40705 , \40706_nR23878 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 ,
         \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724_nR2387a ,
         \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 , \40734 ,
         \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741_nR2387c , \40742 , \40743 , \40744 ,
         \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 ,
         \40755 , \40756 , \40757 , \40758_nR2387e , \40759 , \40760 , \40761 , \40762 , \40763 , \40764 ,
         \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 ,
         \40775_nR23880 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 ,
         \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792_nR23882 , \40793 , \40794 ,
         \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 ,
         \40805 , \40806 , \40807 , \40808 , \40809_nR23884 , \40810 , \40811 , \40812 , \40813 , \40814 ,
         \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 , \40823 , \40824 ,
         \40825 , \40826_nR23886 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 ,
         \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843_nR23888 , \40844 ,
         \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 , \40853 , \40854 ,
         \40855 , \40856 , \40857 , \40858 , \40859 , \40860_nR2388c , \40861 , \40862 , \40863 , \40864 ,
         \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 ,
         \40875 , \40876 , \40877_nR2388e , \40878 , \40879 , \40880 , \40881 , \40882 , \40883 , \40884 ,
         \40885 , \40886 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 ,
         \40895_nR23890 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 ,
         \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912_nR23892 , \40913 , \40914 ,
         \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 ,
         \40925 , \40926 , \40927 , \40928 , \40929_nR23894 , \40930 , \40931 , \40932 , \40933 , \40934 ,
         \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 , \40943 , \40944 ,
         \40945 , \40946_nR23896 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 ,
         \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963_nR23898 , \40964 ,
         \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 , \40973 , \40974 ,
         \40975 , \40976 , \40977 , \40978 , \40979 , \40980_nR2389a , \40981 , \40982 , \40983 , \40984 ,
         \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 ,
         \40995 , \40996 , \40997_nR2389c , \40998 , \40999 , \41000 , \41001 , \41002 , \41003 , \41004 ,
         \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014_nR2389e ,
         \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 ,
         \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031_nR238a2 , \41032 , \41033 , \41034 ,
         \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 , \41043 , \41044 ,
         \41045 , \41046 , \41047 , \41048_nR238a4 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 ,
         \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 ,
         \41065_nR238a6 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 ,
         \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082_nR238a8 , \41083 , \41084 ,
         \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 ,
         \41095 , \41096 , \41097 , \41098 , \41099_nR238aa , \41100 , \41101 , \41102 , \41103 , \41104 ,
         \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 , \41113 , \41114 ,
         \41115 , \41116_nR238ac , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 ,
         \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133_nR238ae , \41134 ,
         \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 , \41143 , \41144 ,
         \41145 , \41146 , \41147 , \41148 , \41149 , \41150_nR238b0 , \41151 , \41152 , \41153 , \41154 ,
         \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 ,
         \41165 , \41166 , \41167_nR238b2 , \41168 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 ,
         \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184_nR238b4 ,
         \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 ,
         \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201_nR238b8 , \41202 , \41203 , \41204 ,
         \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 ,
         \41215 , \41216 , \41217 , \41218_nR238ba , \41219 , \41220 , \41221 , \41222 , \41223 , \41224 ,
         \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 ,
         \41235_nR238bc , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 ,
         \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252_nR238be , \41253 , \41254 ,
         \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 ,
         \41265 , \41266 , \41267 , \41268 , \41269_nR238c0 , \41270 , \41271 , \41272 , \41273 , \41274 ,
         \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 , \41283 , \41284 ,
         \41285 , \41286 , \41287_nR238c2 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 ,
         \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304_nR238c4 ,
         \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 , \41313 , \41314 ,
         \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322_nR238c6 , \41323 , \41324 ,
         \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 ,
         \41335 , \41336 , \41337 , \41338 , \41339_nR238c8 , \41340 , \41341 , \41342 , \41343 , \41344 ,
         \41345 , \41346 , \41347 , \41348 , \41349 , \41350 , \41351 , \41352 , \41353 , \41354 ,
         \41355 , \41356_nR238ca , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 ,
         \41365 , \41366 , \41367 , \41368 , \41369 , \41370 , \41371 , \41372 , \41373_nR238ce , \41374 ,
         \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 , \41383 , \41384 ,
         \41385 , \41386 , \41387 , \41388 , \41389 , \41390_nR238d0 , \41391 , \41392 , \41393 , \41394 ,
         \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 ,
         \41405 , \41406 , \41407_nR238d2 , \41408 , \41409 , \41410 , \41411 , \41412 , \41413 , \41414 ,
         \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424_nR238d4 ,
         \41425 , \41426 , \41427 , \41428 , \41429 , \41430 , \41431 , \41432 , \41433 , \41434 ,
         \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441_nR238d6 , \41442 , \41443 , \41444 ,
         \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451 , \41452 , \41453 , \41454 ,
         \41455 , \41456 , \41457 , \41458_nR238d8 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 ,
         \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472 , \41473 , \41474 ,
         \41475_nR238da , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 ,
         \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492_nR238dc , \41493 , \41494 ,
         \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 , \41503 , \41504 ,
         \41505 , \41506 , \41507 , \41508 , \41509 , \41510_nR238de , \41511 , \41512 , \41513 , \41514 ,
         \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 ,
         \41525 , \41526 , \41527_nR238e0 , \41528 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 ,
         \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544_nR238e4 ,
         \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 ,
         \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561_nR238e6 , \41562 , \41563 , \41564 ,
         \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 ,
         \41575 , \41576 , \41577 , \41578_nR238e8 , \41579 , \41580 , \41581 , \41582 , \41583 , \41584 ,
         \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 ,
         \41595_nR238ea , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 ,
         \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 , \41613 , \41614 ,
         \41615 , \41616 , \41617 , \41618 , \41619 , \41620_nR238f4 , \41621 , \41622 , \41623 , \41624 ,
         \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 ,
         \41635 , \41636_nR2390a , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 , \41643 , \41644 ,
         \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653_nR23920 , \41654 ,
         \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 ,
         \41665 , \41666 , \41667 , \41668 , \41669_nR23936 , \41670 , \41671 , \41672 , \41673 , \41674 ,
         \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683_nR2394c , \41684 ,
         \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 ,
         \41695 , \41696 , \41697 , \41698_nR23962 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 ,
         \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712_nR2396c , \41713 , \41714 ,
         \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 , \41723 , \41724 ,
         \41725 , \41726_nR2396e , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 ,
         \41735 , \41736 , \41737 , \41738 , \41739 , \41740_nR23970 , \41741 , \41742 , \41743 , \41744 ,
         \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 , \41753 , \41754 ,
         \41755_nR23972 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 ,
         \41765 , \41766 , \41767 , \41768 , \41769_nR238f6 , \41770 , \41771 , \41772 , \41773 , \41774 ,
         \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 , \41783_nR238f8 , \41784 ,
         \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 ,
         \41795 , \41796 , \41797_nR238fa , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 ,
         \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811_nR238fc , \41812 , \41813 , \41814 ,
         \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 ,
         \41825 , \41826_nR238fe , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 ,
         \41835 , \41836 , \41837 , \41838 , \41839 , \41840_nR23900 , \41841 , \41842 , \41843 , \41844 ,
         \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854_nR23902 ,
         \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 , \41863 , \41864 ,
         \41865 , \41866 , \41867 , \41868_nR23904 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 ,
         \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882_nR23906 , \41883 , \41884 ,
         \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 , \41893 , \41894 ,
         \41895 , \41896_nR23908 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 ,
         \41905 , \41906 , \41907 , \41908 , \41909 , \41910_nR2390c , \41911 , \41912 , \41913 , \41914 ,
         \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 , \41923 , \41924_nR2390e ,
         \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 ,
         \41935 , \41936 , \41937 , \41938_nR23910 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 ,
         \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952_nR23912 , \41953 , \41954 ,
         \41955 , \41956 , \41957 , \41958 , \41959 , \41960 , \41961 , \41962 , \41963 , \41964 ,
         \41965 , \41966_nR23914 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 ,
         \41975 , \41976 , \41977 , \41978 , \41979 , \41980_nR23916 , \41981 , \41982 , \41983 , \41984 ,
         \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994_nR23918 ,
         \41995 , \41996 , \41997 , \41998 , \41999 , \42000 , \42001 , \42002 , \42003 , \42004 ,
         \42005 , \42006 , \42007 , \42008_nR2391a , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 ,
         \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021 , \42022_nR2391c , \42023 , \42024 ,
         \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 ,
         \42035 , \42036_nR2391e , \42037 , \42038 , \42039 , \42040 , \42041 , \42042 , \42043 , \42044 ,
         \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051_nR23922 , \42052 , \42053 , \42054 ,
         \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 , \42063 , \42064 ,
         \42065_nR23924 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 ,
         \42075 , \42076 , \42077 , \42078 , \42079_nR23926 , \42080 , \42081 , \42082 , \42083 , \42084 ,
         \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 , \42093_nR23928 , \42094 ,
         \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 , \42104 ,
         \42105 , \42106 , \42107_nR2392a , \42108 , \42109 , \42110 , \42111 , \42112 , \42113 , \42114 ,
         \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121_nR2392c , \42122 , \42123 , \42124 ,
         \42125 , \42126 , \42127 , \42128 , \42129 , \42130 , \42131 , \42132 , \42133 , \42134 ,
         \42135_nR2392e , \42136 , \42137 , \42138 , \42139 , \42140 , \42141 , \42142 , \42143 , \42144 ,
         \42145 , \42146 , \42147 , \42148 , \42149_nR23930 , \42150 , \42151 , \42152 , \42153 , \42154 ,
         \42155 , \42156 , \42157 , \42158 , \42159 , \42160 , \42161 , \42162 , \42163_nR23932 , \42164 ,
         \42165 , \42166 , \42167 , \42168 , \42169 , \42170 , \42171 , \42172 , \42173 , \42174 ,
         \42175 , \42176 , \42177_nR23934 , \42178 , \42179 , \42180 , \42181 , \42182 , \42183 , \42184 ,
         \42185 , \42186 , \42187 , \42188 , \42189 , \42190 , \42191_nR23938 , \42192 , \42193 , \42194 ,
         \42195 , \42196 , \42197 , \42198 , \42199 , \42200 , \42201 , \42202 , \42203 , \42204 ,
         \42205_nR2393a , \42206 , \42207 , \42208 , \42209 , \42210 , \42211 , \42212 , \42213 , \42214 ,
         \42215 , \42216 , \42217 , \42218 , \42219_nR2393c , \42220 , \42221 , \42222 , \42223 , \42224 ,
         \42225 , \42226 , \42227 , \42228 , \42229 , \42230 , \42231 , \42232 , \42233_nR2393e , \42234 ,
         \42235 , \42236 , \42237 , \42238 , \42239 , \42240 , \42241 , \42242 , \42243 , \42244 ,
         \42245 , \42246 , \42247_nR23940 , \42248 , \42249 , \42250 , \42251 , \42252 , \42253 , \42254 ,
         \42255 , \42256 , \42257 , \42258 , \42259 , \42260 , \42261_nR23942 , \42262 , \42263 , \42264 ,
         \42265 , \42266 , \42267 , \42268 , \42269 , \42270 , \42271 , \42272 , \42273 , \42274 ,
         \42275_nR23944 , \42276 , \42277 , \42278 , \42279 , \42280 , \42281 , \42282 , \42283 , \42284 ,
         \42285 , \42286 , \42287 , \42288 , \42289_nR23946 , \42290 , \42291 , \42292 , \42293 , \42294 ,
         \42295 , \42296 , \42297 , \42298 , \42299 , \42300 , \42301 , \42302 , \42303_nR23948 , \42304 ,
         \42305 , \42306 , \42307 , \42308 , \42309 , \42310 , \42311 , \42312 , \42313 , \42314 ,
         \42315 , \42316 , \42317_nR2394a , \42318 , \42319 , \42320 , \42321 , \42322 , \42323 , \42324 ,
         \42325 , \42326 , \42327 , \42328 , \42329 , \42330 , \42331_nR2394e , \42332 , \42333 , \42334 ,
         \42335 , \42336 , \42337 , \42338 , \42339 , \42340 , \42341 , \42342 , \42343 , \42344 ,
         \42345_nR23950 , \42346 , \42347 , \42348 , \42349 , \42350 , \42351 , \42352 , \42353 , \42354 ,
         \42355 , \42356 , \42357 , \42358 , \42359_nR23952 , \42360 , \42361 , \42362 , \42363 , \42364 ,
         \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 , \42373_nR23954 , \42374 ,
         \42375 , \42376 , \42377 , \42378 , \42379 , \42380 , \42381 , \42382 , \42383 , \42384 ,
         \42385 , \42386 , \42387_nR23956 , \42388 , \42389 , \42390 , \42391 , \42392 , \42393 , \42394 ,
         \42395 , \42396 , \42397 , \42398 , \42399 , \42400 , \42401_nR23958 , \42402 , \42403 , \42404 ,
         \42405 , \42406 , \42407 , \42408 , \42409 , \42410 , \42411 , \42412 , \42413 , \42414 ,
         \42415_nR2395a , \42416 , \42417 , \42418 , \42419 , \42420 , \42421 , \42422 , \42423 , \42424 ,
         \42425 , \42426 , \42427 , \42428 , \42429_nR2395c , \42430 , \42431 , \42432 , \42433 , \42434 ,
         \42435 , \42436 , \42437 , \42438 , \42439 , \42440 , \42441 , \42442 , \42443_nR2395e , \42444 ,
         \42445 , \42446 , \42447 , \42448 , \42449 , \42450 , \42451 , \42452 , \42453 , \42454 ,
         \42455 , \42456 , \42457_nR23960 , \42458 , \42459 , \42460 , \42461 , \42462 , \42463 , \42464 ,
         \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471_nR23964 , \42472 , \42473 , \42474 ,
         \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 , \42483 , \42484 ,
         \42485_nR23966 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 , \42493 , \42494 ,
         \42495 , \42496 , \42497 , \42498 , \42499_nR23968 , \42500 , \42501 , \42502 , \42503 , \42504 ,
         \42505 , \42506 , \42507 , \42508 , \42509 , \42510 , \42511 , \42512 , \42513_nR2396a , \42514 ,
         \42515 , \42516 , \42517 , \42518 , \42519 , \42520 , \42521 , \42522 , \42523 , \42524 ,
         \42525 , \42526 , \42527 , \42528 , \42529 , \42530 , \42531 , \42532 , \42533_nR23734 , \42534 ,
         \42535 , \42536 , \42537 , \42538 , \42539 , \42540 , \42541 , \42542 , \42543 , \42544 ,
         \42545 , \42546 , \42547 , \42548 , \42549 , \42550_nR23736 , \42551 , \42552 , \42553 , \42554 ,
         \42555 , \42556 , \42557 , \42558 , \42559 , \42560 , \42561 , \42562 , \42563 , \42564 ,
         \42565 , \42566 , \42567_nR23738 , \42568 , \42569 , \42570 , \42571 , \42572 , \42573 , \42574 ,
         \42575 , \42576 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582 , \42583 , \42584_nR2373a ,
         \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591 , \42592 , \42593 , \42594 ,
         \42595 , \42596 , \42597 , \42598 , \42599 , \42600 , \42601_nR2373c , \42602 , \42603 , \42604 ,
         \42605 , \42606 , \42607 , \42608 , \42609 , \42610 , \42611 , \42612 , \42613 , \42614 ,
         \42615 , \42616 , \42617 , \42618_nR2373e , \42619 , \42620 , \42621 , \42622 , \42623 , \42624 ,
         \42625 , \42626 , \42627 , \42628 , \42629 , \42630 , \42631 , \42632 , \42633 , \42634 ,
         \42635_nR23740 , \42636 , \42637 , \42638 , \42639 , \42640 , \42641 , \42642 , \42643 , \42644 ,
         \42645 , \42646 , \42647 , \42648 , \42649 , \42650 , \42651 , \42652_nR23742 , \42653 , \42654 ,
         \42655 , \42656 , \42657 , \42658 , \42659 , \42660 , \42661 , \42662 , \42663 , \42664 ,
         \42665 , \42666 , \42667_nR23744 , \42668 , \42669 , \42670 , \42671 , \42672 , \42673 , \42674 ,
         \42675 , \42676 , \42677 , \42678 , \42679 , \42680 , \42681 , \42682_nR23746 , \42683 , \42684 ,
         \42685 , \42686 , \42687 , \42688 , \42689 , \42690 , \42691 , \42692 , \42693 , \42694 ,
         \42695 , \42696 , \42697_nR23748 , \42698 , \42699 , \42700 , \42701 , \42702 , \42703 , \42704 ,
         \42705 , \42706 , \42707 , \42708 , \42709 , \42710 , \42711 , \42712_nR2374a , \42713 , \42714 ,
         \42715 , \42716 , \42717 , \42718 , \42719 , \42720 , \42721 , \42722 , \42723 , \42724 ,
         \42725 , \42726 , \42727_nR2374c , \42728 , \42729 , \42730 , \42731 , \42732 , \42733 , \42734 ,
         \42735 , \42736 , \42737 , \42738 , \42739 , \42740 , \42741 , \42742_nR2374e , \42743 , \42744 ,
         \42745 , \42746 , \42747 , \42748 , \42749 , \42750 , \42751 , \42752 , \42753 , \42754 ,
         \42755 , \42756 , \42757_nR23750 , \42758 , \42759 , \42760 , \42761 , \42762 , \42763 , \42764 ,
         \42765 , \42766 , \42767 , \42768 , \42769 , \42770 , \42771 , \42772_nR23752 , \42773 , \42774 ,
         \42775 , \42776 , \42777 , \42778 , \42779 , \42780 , \42781 , \42782 , \42783 , \42784 ,
         \42785 , \42786 , \42787_nR23754 , \42788 , \42789 , \42790 , \42791 , \42792 , \42793 , \42794 ,
         \42795 , \42796 , \42797 , \42798 , \42799 , \42800 , \42801 , \42802_nR23756 , \42803 , \42804 ,
         \42805 , \42806 , \42807 , \42808 , \42809 , \42810 , \42811 , \42812 , \42813 , \42814 ,
         \42815 , \42816 , \42817_nR23758 , \42818 , \42819 , \42820 , \42821 , \42822 , \42823 , \42824 ,
         \42825 , \42826 , \42827 , \42828 , \42829 , \42830 , \42831 , \42832_nR2375a , \42833 , \42834 ,
         \42835 , \42836 , \42837 , \42838 , \42839 , \42840 , \42841 , \42842 , \42843 , \42844 ,
         \42845 , \42846 , \42847_nR2375c , \42848 , \42849 , \42850 , \42851 , \42852 , \42853 , \42854 ,
         \42855 , \42856 , \42857 , \42858 , \42859 , \42860 , \42861 , \42862_nR2375e , \42863 , \42864 ,
         \42865 , \42866 , \42867 , \42868 , \42869 , \42870 , \42871 , \42872 , \42873 , \42874 ,
         \42875 , \42876 , \42877_nR23760 , \42878 , \42879 , \42880 , \42881 , \42882 , \42883 , \42884 ,
         \42885 , \42886 , \42887 , \42888 , \42889 , \42890 , \42891 , \42892_nR23762 , \42893 , \42894 ,
         \42895 , \42896 , \42897 , \42898 , \42899 , \42900 , \42901 , \42902 , \42903 , \42904 ,
         \42905 , \42906 , \42907_nR23764 , \42908 , \42909 , \42910 , \42911 , \42912 , \42913 , \42914 ,
         \42915 , \42916 , \42917 , \42918 , \42919 , \42920 , \42921 , \42922_nR23766 , \42923 , \42924 ,
         \42925 , \42926 , \42927 , \42928 , \42929 , \42930 , \42931 , \42932 , \42933 , \42934 ,
         \42935 , \42936 , \42937_nR23768 , \42938 , \42939 , \42940 , \42941 , \42942 , \42943 , \42944 ,
         \42945 , \42946 , \42947 , \42948 , \42949 , \42950 , \42951 , \42952_nR2376a , \42953 , \42954 ,
         \42955 , \42956 , \42957 , \42958 , \42959 , \42960 , \42961 , \42962 , \42963 , \42964 ,
         \42965 , \42966 , \42967_nR2376c , \42968 , \42969 , \42970 , \42971 , \42972 , \42973 , \42974 ,
         \42975 , \42976 , \42977 , \42978 , \42979 , \42980 , \42981 , \42982_nR2376e , \42983 , \42984 ,
         \42985 , \42986 , \42987 , \42988 , \42989 , \42990 , \42991 , \42992 , \42993 , \42994 ,
         \42995 , \42996 , \42997_nR23770 , \42998 , \42999 , \43000 , \43001 , \43002 , \43003 , \43004 ,
         \43005 , \43006 , \43007 , \43008 , \43009 , \43010 , \43011 , \43012_nR23772 , \43013 , \43014 ,
         \43015 , \43016 , \43017 , \43018 , \43019 , \43020 , \43021 , \43022 , \43023 , \43024 ,
         \43025 , \43026 , \43027_nR2398c , \43028 , \43029 , \43030 , \43031 , \43032 , \43033 , \43034 ,
         \43035 , \43036 , \43037 , \43038_nR2398e , \43039 , \43040 , \43041 , \43042 , \43043 , \43044 ,
         \43045 , \43046 , \43047 , \43048_nR23990 , \43049 , \43050 , \43051 , \43052 , \43053 , \43054 ,
         \43055 , \43056 , \43057 , \43058_nR23992 , \43059 , \43060 , \43061 , \43062 , \43063 , \43064 ,
         \43065 , \43066 , \43067 , \43068_nR23994 , \43069 , \43070 , \43071 , \43072 , \43073 , \43074 ,
         \43075 , \43076 , \43077 , \43078_nR23996 , \43079 , \43080 , \43081 , \43082 , \43083 , \43084 ,
         \43085 , \43086 , \43087 , \43088_nR23998 , \43089 , \43090 , \43091 , \43092 , \43093 , \43094 ,
         \43095 , \43096 , \43097 , \43098_nR2399a , \43099 , \43100 , \43101 , \43102 , \43103 , \43104 ,
         \43105 , \43106 , \43107 , \43108_nR2398a , \43109 , \43110 , \43111 , \43112 , \43113 , \43114 ,
         \43115 , \43116 , \43117 , \43118_nR2399c , \43119 , \43120 , \43121 , \43122 , \43123 , \43124 ,
         \43125 , \43126 , \43127 , \43128_nR2399e , \43129 , \43130 , \43131 , \43132 , \43133 , \43134 ,
         \43135 , \43136 , \43137 , \43138_nR239a0 , \43139 , \43140 , \43141 , \43142 , \43143 , \43144 ,
         \43145 , \43146 , \43147 , \43148_nR239a2 , \43149 , \43150 , \43151 , \43152 , \43153 , \43154 ,
         \43155 , \43156 , \43157 , \43158 , \43159 , \43160 , \43161 , \43162 , \43163 , \43164 ,
         \43165 , \43166 , \43167 , \43168 , \43169 , \43170 , \43171 , \43172 , \43173 , \43174 ,
         \43175 , \43176 , \43177 , \43178 , \43179 , \43180 , \43181 , \43182 , \43183 , \43184 ,
         \43185 , \43186 , \43187 , \43188 , \43189 , \43190 , \43191 , \43192 , \43193 , \43194 ,
         \43195 , \43196 , \43197 , \43198 , \43199 , \43200 , \43201 , \43202 , \43203 , \43204 ,
         \43205 , \43206 , \43207 , \43208 , \43209 , \43210 , \43211 , \43212 , \43213 , \43214 ,
         \43215 , \43216 , \43217 , \43218 , \43219 , \43220 , \43221 , \43222 , \43223 , \43224 ,
         \43225 , \43226 , \43227 , \43228 , \43229 , \43230 , \43231 , \43232 , \43233 , \43234 ,
         \43235 , \43236 , \43237 , \43238 , \43239 , \43240 , \43241 , \43242 , \43243 , \43244 ,
         \43245 , \43246 , \43247 , \43248 , \43249 , \43250 , \43251 , \43252 , \43253 , \43254 ,
         \43255 , \43256 , \43257 , \43258 , \43259 , \43260 , \43261 , \43262 , \43263 , \43264 ,
         \43265 , \43266 , \43267 , \43268 , \43269 , \43270 , \43271 , \43272 , \43273 , \43274 ,
         \43275 , \43276 , \43277 , \43278 , \43279 , \43280 , \43281 , \43282 , \43283 , \43284 ,
         \43285 , \43286 , \43287 , \43288 , \43289 , \43290 , \43291 , \43292 , \43293 , \43294 ,
         \43295 , \43296 , \43297 , \43298 , \43299 , \43300 , \43301 , \43302 , \43303 , \43304 ,
         \43305 , \43306 , \43307 , \43308 , \43309 , \43310 , \43311 , \43312 , \43313 , \43314 ,
         \43315 , \43316 , \43317 , \43318 , \43319 , \43320 , \43321 , \43322 , \43323 , \43324 ,
         \43325 , \43326 , \43327 , \43328 , \43329 , \43330 , \43331 , \43332 , \43333 , \43334 ,
         \43335 , \43336 , \43337 , \43338 , \43339 , \43340 , \43341 , \43342 , \43343_nR23988 , \43344 ,
         \43345 , \43346 , \43347 , \43348_nR239ba , \43349 , \43350 , \43351 , \43352 , \43353_nR239bc , \43354 ,
         \43355 , \43356 , \43357 , \43358 , \43359_nR239be , \43360 , \43361 , \43362 , \43363 , \43364 ,
         \43365 , \43366 , \43367 , \43368 , \43369 , \43370 , \43371 , \43372 , \43373 , \43374 ,
         \43375 , \43376 , \43377 , \43378 , \43379 , \43380 , \43381 , \43382 , \43383 , \43384 ,
         \43385 , \43386 , \43387 , \43388 , \43389 , \43390 , \43391 , \43392 , \43393 , \43394 ,
         \43395 , \43396 , \43397 , \43398 , \43399 , \43400 , \43401 , \43402 , \43403 , \43404 ,
         \43405 , \43406 , \43407 , \43408 , \43409 , \43410 , \43411 , \43412 , \43413 , \43414 ,
         \43415 , \43416 , \43417 , \43418 , \43419_nR234dc , \43420 , \43421 , \43422 , \43423 , \43424 ,
         \43425 , \43426 , \43427 , \43428 , \43429 , \43430 , \43431 , \43432 , \43433 , \43434 ,
         \43435 , \43436 , \43437 , \43438 , \43439 , \43440 , \43441_nR234f2 , \43442 , \43443 , \43444 ,
         \43445 , \43446 , \43447 , \43448 , \43449 , \43450 , \43451 , \43452 , \43453 , \43454 ,
         \43455 , \43456 , \43457 , \43458 , \43459 , \43460_nR23508 , \43461 , \43462 , \43463 , \43464 ,
         \43465 , \43466 , \43467 , \43468 , \43469 , \43470 , \43471 , \43472 , \43473 , \43474 ,
         \43475 , \43476 , \43477 , \43478 , \43479 , \43480_nR2351e , \43481 , \43482 , \43483 , \43484 ,
         \43485 , \43486 , \43487 , \43488 , \43489 , \43490 , \43491 , \43492 , \43493 , \43494 ,
         \43495 , \43496 , \43497 , \43498 , \43499 , \43500 , \43501_nR23534 , \43502 , \43503 , \43504 ,
         \43505 , \43506 , \43507 , \43508 , \43509 , \43510 , \43511 , \43512 , \43513 , \43514 ,
         \43515 , \43516 , \43517 , \43518 , \43519 , \43520 , \43521 , \43522 , \43523 , \43524_nR2354a ,
         \43525 , \43526 , \43527 , \43528 , \43529 , \43530 , \43531 , \43532 , \43533 , \43534 ,
         \43535 , \43536 , \43537 , \43538 , \43539 , \43540 , \43541 , \43542 , \43543 , \43544 ,
         \43545_nR23554 , \43546 , \43547 , \43548 , \43549 , \43550 , \43551 , \43552 , \43553 , \43554 ,
         \43555 , \43556 , \43557 , \43558 , \43559 , \43560 , \43561 , \43562 , \43563 , \43564 ,
         \43565 , \43566_nR23556 , \43567 , \43568 , \43569 , \43570 , \43571 , \43572 , \43573 , \43574 ,
         \43575 , \43576 , \43577 , \43578 , \43579 , \43580 , \43581 , \43582 , \43583 , \43584 ,
         \43585 , \43586 , \43587_nR23558 , \43588 , \43589 , \43590 , \43591 , \43592 , \43593 , \43594 ,
         \43595 , \43596 , \43597 , \43598 , \43599 , \43600 , \43601 , \43602 , \43603 , \43604 ,
         \43605 , \43606 , \43607 , \43608 , \43609 , \43610 , \43611_nR2355a , \43612 , \43613 , \43614 ,
         \43615 , \43616 , \43617 , \43618 , \43619 , \43620 , \43621 , \43622 , \43623 , \43624 ,
         \43625 , \43626 , \43627 , \43628 , \43629 , \43630 , \43631 , \43632_nR234de , \43633 , \43634 ,
         \43635 , \43636 , \43637 , \43638 , \43639 , \43640 , \43641 , \43642 , \43643 , \43644 ,
         \43645 , \43646 , \43647 , \43648 , \43649 , \43650_nR234e0 , \43651 , \43652 , \43653 , \43654 ,
         \43655 , \43656 , \43657 , \43658 , \43659 , \43660 , \43661 , \43662 , \43663 , \43664 ,
         \43665 , \43666 , \43667 , \43668 , \43669 , \43670 , \43671_nR234e2 , \43672 , \43673 , \43674 ,
         \43675 , \43676 , \43677 , \43678 , \43679 , \43680 , \43681 , \43682 , \43683 , \43684 ,
         \43685 , \43686 , \43687 , \43688 , \43689 , \43690_nR234e4 , \43691 , \43692 , \43693 , \43694 ,
         \43695 , \43696 , \43697 , \43698 , \43699 , \43700 , \43701 , \43702 , \43703 , \43704 ,
         \43705 , \43706 , \43707 , \43708_nR234e6 , \43709 , \43710 , \43711 , \43712 , \43713 , \43714 ,
         \43715 , \43716 , \43717 , \43718 , \43719 , \43720 , \43721 , \43722 , \43723 , \43724 ,
         \43725 , \43726 , \43727 , \43728_nR234e8 , \43729 , \43730 , \43731 , \43732 , \43733 , \43734 ,
         \43735 , \43736 , \43737 , \43738 , \43739 , \43740 , \43741 , \43742 , \43743 , \43744 ,
         \43745 , \43746 , \43747 , \43748_nR234ea , \43749 , \43750 , \43751 , \43752 , \43753 , \43754 ,
         \43755 , \43756 , \43757 , \43758 , \43759 , \43760 , \43761 , \43762 , \43763 , \43764 ,
         \43765 , \43766_nR234ec , \43767 , \43768 , \43769 , \43770 , \43771 , \43772 , \43773 , \43774 ,
         \43775 , \43776 , \43777 , \43778 , \43779 , \43780 , \43781 , \43782 , \43783 , \43784 ,
         \43785 , \43786_nR234ee , \43787 , \43788 , \43789 , \43790 , \43791 , \43792 , \43793 , \43794 ,
         \43795 , \43796 , \43797 , \43798 , \43799 , \43800 , \43801 , \43802 , \43803 , \43804 ,
         \43805_nR234f0 , \43806 , \43807 , \43808 , \43809 , \43810 , \43811 , \43812 , \43813 , \43814 ,
         \43815 , \43816 , \43817 , \43818 , \43819 , \43820 , \43821 , \43822 , \43823_nR234f4 , \43824 ,
         \43825 , \43826 , \43827 , \43828 , \43829 , \43830 , \43831 , \43832 , \43833 , \43834 ,
         \43835 , \43836 , \43837 , \43838 , \43839 , \43840 , \43841 , \43842_nR234f6 , \43843 , \43844 ,
         \43845 , \43846 , \43847 , \43848 , \43849 , \43850 , \43851 , \43852 , \43853 , \43854 ,
         \43855 , \43856 , \43857 , \43858 , \43859 , \43860 , \43861 , \43862_nR234f8 , \43863 , \43864 ,
         \43865 , \43866 , \43867 , \43868 , \43869 , \43870 , \43871 , \43872 , \43873 , \43874 ,
         \43875 , \43876 , \43877 , \43878 , \43879 , \43880 , \43881 , \43882_nR234fa , \43883 , \43884 ,
         \43885 , \43886 , \43887 , \43888 , \43889 , \43890 , \43891 , \43892 , \43893 , \43894 ,
         \43895 , \43896 , \43897 , \43898 , \43899 , \43900_nR234fc , \43901 , \43902 , \43903 , \43904 ,
         \43905 , \43906 , \43907 , \43908 , \43909 , \43910 , \43911 , \43912 , \43913 , \43914 ,
         \43915 , \43916 , \43917 , \43918 , \43919 , \43920_nR234fe , \43921 , \43922 , \43923 , \43924 ,
         \43925 , \43926 , \43927 , \43928 , \43929 , \43930 , \43931 , \43932 , \43933 , \43934 ,
         \43935 , \43936 , \43937 , \43938 , \43939_nR23500 , \43940 , \43941 , \43942 , \43943 , \43944 ,
         \43945 , \43946 , \43947 , \43948 , \43949 , \43950 , \43951 , \43952 , \43953 , \43954 ,
         \43955 , \43956 , \43957 , \43958 , \43959_nR23502 , \43960 , \43961 , \43962 , \43963 , \43964 ,
         \43965 , \43966 , \43967 , \43968 , \43969 , \43970 , \43971 , \43972 , \43973 , \43974 ,
         \43975 , \43976 , \43977 , \43978 , \43979_nR23504 , \43980 , \43981 , \43982 , \43983 , \43984 ,
         \43985 , \43986 , \43987 , \43988 , \43989 , \43990 , \43991 , \43992 , \43993 , \43994 ,
         \43995 , \43996 , \43997_nR23506 , \43998 , \43999 , \44000 , \44001 , \44002 , \44003 , \44004 ,
         \44005 , \44006 , \44007 , \44008 , \44009 , \44010 , \44011 , \44012 , \44013 , \44014 ,
         \44015 , \44016_nR2350a , \44017 , \44018 , \44019 , \44020 , \44021 , \44022 , \44023 , \44024 ,
         \44025 , \44026 , \44027 , \44028 , \44029 , \44030 , \44031 , \44032 , \44033 , \44034 ,
         \44035_nR2350c , \44036 , \44037 , \44038 , \44039 , \44040 , \44041 , \44042 , \44043 , \44044 ,
         \44045 , \44046 , \44047 , \44048 , \44049 , \44050 , \44051 , \44052 , \44053_nR2350e , \44054 ,
         \44055 , \44056 , \44057 , \44058 , \44059 , \44060 , \44061 , \44062 , \44063 , \44064 ,
         \44065 , \44066 , \44067 , \44068 , \44069 , \44070 , \44071 , \44072_nR23510 , \44073 , \44074 ,
         \44075 , \44076 , \44077 , \44078 , \44079 , \44080 , \44081 , \44082 , \44083 , \44084 ,
         \44085 , \44086 , \44087 , \44088 , \44089 , \44090 , \44091 , \44092_nR23512 , \44093 , \44094 ,
         \44095 , \44096 , \44097 , \44098 , \44099 , \44100 , \44101 , \44102 , \44103 , \44104 ,
         \44105 , \44106 , \44107 , \44108 , \44109 , \44110 , \44111_nR23514 , \44112 , \44113 , \44114 ,
         \44115 , \44116 , \44117 , \44118 , \44119 , \44120 , \44121 , \44122 , \44123 , \44124 ,
         \44125 , \44126 , \44127 , \44128 , \44129_nR23516 , \44130 , \44131 , \44132 , \44133 , \44134 ,
         \44135 , \44136 , \44137 , \44138 , \44139 , \44140 , \44141 , \44142 , \44143 , \44144 ,
         \44145 , \44146 , \44147 , \44148 , \44149_nR23518 , \44150 , \44151 , \44152 , \44153 , \44154 ,
         \44155 , \44156 , \44157 , \44158 , \44159 , \44160 , \44161 , \44162 , \44163 , \44164 ,
         \44165 , \44166 , \44167 , \44168 , \44169_nR2351a , \44170 , \44171 , \44172 , \44173 , \44174 ,
         \44175 , \44176 , \44177 , \44178 , \44179 , \44180 , \44181 , \44182 , \44183 , \44184 ,
         \44185 , \44186 , \44187 , \44188 , \44189_nR2351c , \44190 , \44191 , \44192 , \44193 , \44194 ,
         \44195 , \44196 , \44197 , \44198 , \44199 , \44200 , \44201 , \44202 , \44203 , \44204 ,
         \44205 , \44206 , \44207 , \44208_nR23520 , \44209 , \44210 , \44211 , \44212 , \44213 , \44214 ,
         \44215 , \44216 , \44217 , \44218 , \44219 , \44220 , \44221 , \44222 , \44223 , \44224 ,
         \44225 , \44226_nR23522 , \44227 , \44228 , \44229 , \44230 , \44231 , \44232 , \44233 , \44234 ,
         \44235 , \44236 , \44237 , \44238 , \44239 , \44240 , \44241 , \44242 , \44243 , \44244_nR23524 ,
         \44245 , \44246 , \44247 , \44248 , \44249 , \44250 , \44251 , \44252 , \44253 , \44254 ,
         \44255 , \44256 , \44257 , \44258 , \44259 , \44260 , \44261 , \44262 , \44263_nR23526 , \44264 ,
         \44265 , \44266 , \44267 , \44268 , \44269 , \44270 , \44271 , \44272 , \44273 , \44274 ,
         \44275 , \44276 , \44277 , \44278 , \44279 , \44280 , \44281 , \44282 , \44283 , \44284_nR23528 ,
         \44285 , \44286 , \44287 , \44288 , \44289 , \44290 , \44291 , \44292 , \44293 , \44294 ,
         \44295 , \44296 , \44297 , \44298 , \44299 , \44300 , \44301 , \44302 , \44303 , \44304_nR2352a ,
         \44305 , \44306 , \44307 , \44308 , \44309 , \44310 , \44311 , \44312 , \44313 , \44314 ,
         \44315 , \44316 , \44317 , \44318 , \44319 , \44320 , \44321 , \44322 , \44323 , \44324_nR2352c ,
         \44325 , \44326 , \44327 , \44328 , \44329 , \44330 , \44331 , \44332 , \44333 , \44334 ,
         \44335 , \44336 , \44337 , \44338 , \44339 , \44340 , \44341 , \44342_nR2352e , \44343 , \44344 ,
         \44345 , \44346 , \44347 , \44348 , \44349 , \44350 , \44351 , \44352 , \44353 , \44354 ,
         \44355 , \44356 , \44357 , \44358 , \44359 , \44360 , \44361 , \44362_nR23530 , \44363 , \44364 ,
         \44365 , \44366 , \44367 , \44368 , \44369 , \44370 , \44371 , \44372 , \44373 , \44374 ,
         \44375 , \44376 , \44377 , \44378 , \44379 , \44380_nR23532 , \44381 , \44382 , \44383 , \44384 ,
         \44385 , \44386 , \44387 , \44388 , \44389 , \44390 , \44391 , \44392 , \44393 , \44394 ,
         \44395 , \44396 , \44397 , \44398_nR23536 , \44399 , \44400 , \44401 , \44402 , \44403 , \44404 ,
         \44405 , \44406 , \44407 , \44408 , \44409 , \44410 , \44411 , \44412 , \44413 , \44414 ,
         \44415 , \44416 , \44417_nR23538 , \44418 , \44419 , \44420 , \44421 , \44422 , \44423 , \44424 ,
         \44425 , \44426 , \44427 , \44428 , \44429 , \44430 , \44431 , \44432 , \44433 , \44434 ,
         \44435_nR2353a , \44436 , \44437 , \44438 , \44439 , \44440 , \44441 , \44442 , \44443 , \44444 ,
         \44445 , \44446 , \44447 , \44448 , \44449 , \44450 , \44451 , \44452 , \44453 , \44454 ,
         \44455_nR2353c , \44456 , \44457 , \44458 , \44459 , \44460 , \44461 , \44462 , \44463 , \44464 ,
         \44465 , \44466 , \44467 , \44468 , \44469 , \44470 , \44471 , \44472 , \44473_nR2353e , \44474 ,
         \44475 , \44476 , \44477 , \44478 , \44479 , \44480 , \44481 , \44482 , \44483 , \44484 ,
         \44485 , \44486 , \44487 , \44488 , \44489 , \44490 , \44491_nR23540 , \44492 , \44493 , \44494 ,
         \44495 , \44496 , \44497 , \44498 , \44499 , \44500 , \44501 , \44502 , \44503 , \44504 ,
         \44505 , \44506 , \44507 , \44508 , \44509 , \44510 , \44511 , \44512 , \44513_nR23542 , \44514 ,
         \44515 , \44516 , \44517 , \44518 , \44519 , \44520 , \44521 , \44522 , \44523 , \44524 ,
         \44525 , \44526 , \44527 , \44528 , \44529 , \44530 , \44531 , \44532 , \44533 , \44534_nR23544 ,
         \44535 , \44536 , \44537 , \44538 , \44539 , \44540 , \44541 , \44542 , \44543 , \44544 ,
         \44545 , \44546 , \44547 , \44548 , \44549 , \44550 , \44551 , \44552 , \44553_nR23546 , \44554 ,
         \44555 , \44556 , \44557 , \44558 , \44559 , \44560 , \44561 , \44562 , \44563 , \44564 ,
         \44565 , \44566 , \44567 , \44568 , \44569 , \44570 , \44571_nR23548 , \44572 , \44573 , \44574 ,
         \44575 , \44576 , \44577 , \44578 , \44579 , \44580 , \44581 , \44582 , \44583 , \44584 ,
         \44585 , \44586 , \44587 , \44588 , \44589_nR2354c , \44590 , \44591 , \44592 , \44593 , \44594 ,
         \44595 , \44596 , \44597 , \44598 , \44599 , \44600 , \44601 , \44602 , \44603 , \44604 ,
         \44605 , \44606 , \44607 , \44608 , \44609_nR2354e , \44610 , \44611 , \44612 , \44613 , \44614 ,
         \44615 , \44616 , \44617 , \44618 , \44619 , \44620 , \44621 , \44622 , \44623 , \44624 ,
         \44625 , \44626 , \44627 , \44628_nR23550 , \44629 , \44630 , \44631 , \44632 , \44633 , \44634 ,
         \44635 , \44636 , \44637 , \44638 , \44639 , \44640 , \44641 , \44642 , \44643 , \44644 ,
         \44645 , \44646_nR23552 , \44647 , \44648 , \44649 , \44650 , \44651 , \44652 , \44653 , \44654 ,
         \44655 , \44656 , \44657 , \44658 , \44659 , \44660 , \44661 , \44662 , \44663 , \44664 ,
         \44665 , \44666 , \44667 , \44668 , \44669 , \44670 , \44671 , \44672 , \44673 , \44674 ,
         \44675 , \44676 , \44677 , \44678 , \44679 , \44680_nR2355c , \44681 , \44682 , \44683 , \44684 ,
         \44685 , \44686 , \44687 , \44688 , \44689 , \44690 , \44691 , \44692 , \44693 , \44694 ,
         \44695 , \44696 , \44697 , \44698 , \44699 , \44700_nR23572 , \44701 , \44702 , \44703 , \44704 ,
         \44705 , \44706 , \44707 , \44708 , \44709 , \44710 , \44711 , \44712 , \44713 , \44714 ,
         \44715 , \44716 , \44717 , \44718 , \44719_nR23588 , \44720 , \44721 , \44722 , \44723 , \44724 ,
         \44725 , \44726 , \44727 , \44728 , \44729 , \44730 , \44731 , \44732 , \44733 , \44734 ,
         \44735 , \44736 , \44737 , \44738_nR2359e , \44739 , \44740 , \44741 , \44742 , \44743 , \44744 ,
         \44745 , \44746 , \44747 , \44748 , \44749 , \44750 , \44751 , \44752 , \44753 , \44754 ,
         \44755 , \44756_nR235b4 , \44757 , \44758 , \44759 , \44760 , \44761 , \44762 , \44763 , \44764 ,
         \44765 , \44766 , \44767 , \44768 , \44769 , \44770 , \44771 , \44772 , \44773 , \44774 ,
         \44775 , \44776 , \44777_nR235ca , \44778 , \44779 , \44780 , \44781 , \44782 , \44783 , \44784 ,
         \44785 , \44786 , \44787 , \44788 , \44789 , \44790 , \44791 , \44792 , \44793 , \44794 ,
         \44795 , \44796_nR235d4 , \44797 , \44798 , \44799 , \44800 , \44801 , \44802 , \44803 , \44804 ,
         \44805 , \44806 , \44807 , \44808 , \44809 , \44810 , \44811 , \44812 , \44813 , \44814 ,
         \44815_nR235d6 , \44816 , \44817 , \44818 , \44819 , \44820 , \44821 , \44822 , \44823 , \44824 ,
         \44825 , \44826 , \44827 , \44828 , \44829 , \44830 , \44831 , \44832 , \44833_nR235d8 , \44834 ,
         \44835 , \44836 , \44837 , \44838 , \44839 , \44840 , \44841 , \44842 , \44843 , \44844 ,
         \44845 , \44846 , \44847 , \44848 , \44849 , \44850 , \44851 , \44852_nR235da , \44853 , \44854 ,
         \44855 , \44856 , \44857 , \44858 , \44859 , \44860 , \44861 , \44862 , \44863 , \44864 ,
         \44865 , \44866 , \44867 , \44868 , \44869 , \44870_nR2355e , \44871 , \44872 , \44873 , \44874 ,
         \44875 , \44876 , \44877 , \44878 , \44879 , \44880 , \44881 , \44882 , \44883 , \44884 ,
         \44885 , \44886 , \44887 , \44888 , \44889_nR23560 , \44890 , \44891 , \44892 , \44893 , \44894 ,
         \44895 , \44896 , \44897 , \44898 , \44899 , \44900 , \44901 , \44902 , \44903 , \44904 ,
         \44905 , \44906 , \44907 , \44908_nR23562 , \44909 , \44910 , \44911 , \44912 , \44913 , \44914 ,
         \44915 , \44916 , \44917 , \44918 , \44919 , \44920 , \44921 , \44922 , \44923 , \44924 ,
         \44925 , \44926_nR23564 , \44927 , \44928 , \44929 , \44930 , \44931 , \44932 , \44933 , \44934 ,
         \44935 , \44936 , \44937 , \44938 , \44939 , \44940 , \44941 , \44942 , \44943 , \44944_nR23566 ,
         \44945 , \44946 , \44947 , \44948 , \44949 , \44950 , \44951 , \44952 , \44953 , \44954 ,
         \44955 , \44956 , \44957 , \44958 , \44959 , \44960 , \44961 , \44962_nR23568 , \44963 , \44964 ,
         \44965 , \44966 , \44967 , \44968 , \44969 , \44970 , \44971 , \44972 , \44973 , \44974 ,
         \44975 , \44976 , \44977 , \44978 , \44979 , \44980_nR2356a , \44981 , \44982 , \44983 , \44984 ,
         \44985 , \44986 , \44987 , \44988 , \44989 , \44990 , \44991 , \44992 , \44993 , \44994 ,
         \44995 , \44996 , \44997 , \44998_nR2356c , \44999 , \45000 , \45001 , \45002 , \45003 , \45004 ,
         \45005 , \45006 , \45007 , \45008 , \45009 , \45010 , \45011 , \45012 , \45013 , \45014 ,
         \45015 , \45016_nR2356e , \45017 , \45018 , \45019 , \45020 , \45021 , \45022 , \45023 , \45024 ,
         \45025 , \45026 , \45027 , \45028 , \45029 , \45030 , \45031 , \45032 , \45033 , \45034_nR23570 ,
         \45035 , \45036 , \45037 , \45038 , \45039 , \45040 , \45041 , \45042 , \45043 , \45044 ,
         \45045 , \45046 , \45047 , \45048 , \45049 , \45050 , \45051 , \45052_nR23574 , \45053 , \45054 ,
         \45055 , \45056 , \45057 , \45058 , \45059 , \45060 , \45061 , \45062 , \45063 , \45064 ,
         \45065 , \45066 , \45067 , \45068 , \45069 , \45070_nR23576 , \45071 , \45072 , \45073 , \45074 ,
         \45075 , \45076 , \45077 , \45078 , \45079 , \45080 , \45081 , \45082 , \45083 , \45084 ,
         \45085 , \45086 , \45087 , \45088_nR23578 , \45089 , \45090 , \45091 , \45092 , \45093 , \45094 ,
         \45095 , \45096 , \45097 , \45098 , \45099 , \45100 , \45101 , \45102 , \45103 , \45104 ,
         \45105 , \45106_nR2357a , \45107 , \45108 , \45109 , \45110 , \45111 , \45112 , \45113 , \45114 ,
         \45115 , \45116 , \45117 , \45118 , \45119 , \45120 , \45121 , \45122 , \45123 , \45124_nR2357c ,
         \45125 , \45126 , \45127 , \45128 , \45129 , \45130 , \45131 , \45132 , \45133 , \45134 ,
         \45135 , \45136 , \45137 , \45138 , \45139 , \45140 , \45141 , \45142_nR2357e , \45143 , \45144 ,
         \45145 , \45146 , \45147 , \45148 , \45149 , \45150 , \45151 , \45152 , \45153 , \45154 ,
         \45155 , \45156 , \45157 , \45158 , \45159 , \45160_nR23580 , \45161 , \45162 , \45163 , \45164 ,
         \45165 , \45166 , \45167 , \45168 , \45169 , \45170 , \45171 , \45172 , \45173 , \45174 ,
         \45175 , \45176 , \45177 , \45178_nR23582 , \45179 , \45180 , \45181 , \45182 , \45183 , \45184 ,
         \45185 , \45186 , \45187 , \45188 , \45189 , \45190 , \45191 , \45192 , \45193 , \45194 ,
         \45195 , \45196_nR23584 , \45197 , \45198 , \45199 , \45200 , \45201 , \45202 , \45203 , \45204 ,
         \45205 , \45206 , \45207 , \45208 , \45209 , \45210 , \45211 , \45212 , \45213 , \45214_nR23586 ,
         \45215 , \45216 , \45217 , \45218 , \45219 , \45220 , \45221 , \45222 , \45223 , \45224 ,
         \45225 , \45226 , \45227 , \45228 , \45229 , \45230 , \45231 , \45232_nR2358a , \45233 , \45234 ,
         \45235 , \45236 , \45237 , \45238 , \45239 , \45240 , \45241 , \45242 , \45243 , \45244 ,
         \45245 , \45246 , \45247 , \45248 , \45249 , \45250_nR2358c , \45251 , \45252 , \45253 , \45254 ,
         \45255 , \45256 , \45257 , \45258 , \45259 , \45260 , \45261 , \45262 , \45263 , \45264 ,
         \45265 , \45266 , \45267 , \45268_nR2358e , \45269 , \45270 , \45271 , \45272 , \45273 , \45274 ,
         \45275 , \45276 , \45277 , \45278 , \45279 , \45280 , \45281 , \45282 , \45283 , \45284 ,
         \45285 , \45286_nR23590 , \45287 , \45288 , \45289 , \45290 , \45291 , \45292 , \45293 , \45294 ,
         \45295 , \45296 , \45297 , \45298 , \45299 , \45300 , \45301 , \45302 , \45303 , \45304_nR23592 ,
         \45305 , \45306 , \45307 , \45308 , \45309 , \45310 , \45311 , \45312 , \45313 , \45314 ,
         \45315 , \45316 , \45317 , \45318 , \45319 , \45320 , \45321 , \45322_nR23594 , \45323 , \45324 ,
         \45325 , \45326 , \45327 , \45328 , \45329 , \45330 , \45331 , \45332 , \45333 , \45334 ,
         \45335 , \45336 , \45337 , \45338 , \45339 , \45340 , \45341_nR23596 , \45342 , \45343 , \45344 ,
         \45345 , \45346 , \45347 , \45348 , \45349 , \45350 , \45351 , \45352 , \45353 , \45354 ,
         \45355 , \45356 , \45357 , \45358 , \45359_nR23598 , \45360 , \45361 , \45362 , \45363 , \45364 ,
         \45365 , \45366 , \45367 , \45368 , \45369 , \45370 , \45371 , \45372 , \45373 , \45374 ,
         \45375 , \45376 , \45377 , \45378_nR2359a , \45379 , \45380 , \45381 , \45382 , \45383 , \45384 ,
         \45385 , \45386 , \45387 , \45388 , \45389 , \45390 , \45391 , \45392 , \45393 , \45394 ,
         \45395 , \45396_nR2359c , \45397 , \45398 , \45399 , \45400 , \45401 , \45402 , \45403 , \45404 ,
         \45405 , \45406 , \45407 , \45408 , \45409 , \45410 , \45411 , \45412 , \45413 , \45414_nR235a0 ,
         \45415 , \45416 , \45417 , \45418 , \45419 , \45420 , \45421 , \45422 , \45423 , \45424 ,
         \45425 , \45426 , \45427 , \45428 , \45429 , \45430 , \45431 , \45432_nR235a2 , \45433 , \45434 ,
         \45435 , \45436 , \45437 , \45438 , \45439 , \45440 , \45441 , \45442 , \45443 , \45444 ,
         \45445 , \45446 , \45447 , \45448 , \45449 , \45450_nR235a4 , \45451 , \45452 , \45453 , \45454 ,
         \45455 , \45456 , \45457 , \45458 , \45459 , \45460 , \45461 , \45462 , \45463 , \45464 ,
         \45465 , \45466 , \45467 , \45468_nR235a6 , \45469 , \45470 , \45471 , \45472 , \45473 , \45474 ,
         \45475 , \45476 , \45477 , \45478 , \45479 , \45480 , \45481 , \45482 , \45483 , \45484 ,
         \45485 , \45486_nR235a8 , \45487 , \45488 , \45489 , \45490 , \45491 , \45492 , \45493 , \45494 ,
         \45495 , \45496 , \45497 , \45498 , \45499 , \45500 , \45501 , \45502 , \45503 , \45504_nR235aa ,
         \45505 , \45506 , \45507 , \45508 , \45509 , \45510 , \45511 , \45512 , \45513 , \45514 ,
         \45515 , \45516 , \45517 , \45518 , \45519 , \45520 , \45521 , \45522_nR235ac , \45523 , \45524 ,
         \45525 , \45526 , \45527 , \45528 , \45529 , \45530 , \45531 , \45532 , \45533 , \45534 ,
         \45535 , \45536 , \45537 , \45538 , \45539 , \45540_nR235ae , \45541 , \45542 , \45543 , \45544 ,
         \45545 , \45546 , \45547 , \45548 , \45549 , \45550 , \45551 , \45552 , \45553 , \45554 ,
         \45555 , \45556 , \45557 , \45558_nR235b0 , \45559 , \45560 , \45561 , \45562 , \45563 , \45564 ,
         \45565 , \45566 , \45567 , \45568 , \45569 , \45570 , \45571 , \45572 , \45573 , \45574 ,
         \45575 , \45576_nR235b2 , \45577 , \45578 , \45579 , \45580 , \45581 , \45582 , \45583 , \45584 ,
         \45585 , \45586 , \45587 , \45588 , \45589 , \45590 , \45591 , \45592 , \45593 , \45594_nR235b6 ,
         \45595 , \45596 , \45597 , \45598 , \45599 , \45600 , \45601 , \45602 , \45603 , \45604 ,
         \45605 , \45606 , \45607 , \45608 , \45609 , \45610 , \45611 , \45612_nR235b8 , \45613 , \45614 ,
         \45615 , \45616 , \45617 , \45618 , \45619 , \45620 , \45621 , \45622 , \45623 , \45624 ,
         \45625 , \45626 , \45627 , \45628 , \45629 , \45630 , \45631_nR235ba , \45632 , \45633 , \45634 ,
         \45635 , \45636 , \45637 , \45638 , \45639 , \45640 , \45641 , \45642 , \45643 , \45644 ,
         \45645 , \45646 , \45647 , \45648 , \45649_nR235bc , \45650 , \45651 , \45652 , \45653 , \45654 ,
         \45655 , \45656 , \45657 , \45658 , \45659 , \45660 , \45661 , \45662 , \45663 , \45664 ,
         \45665 , \45666 , \45667_nR235be , \45668 , \45669 , \45670 , \45671 , \45672 , \45673 , \45674 ,
         \45675 , \45676 , \45677 , \45678 , \45679 , \45680 , \45681 , \45682 , \45683 , \45684 ,
         \45685_nR235c0 , \45686 , \45687 , \45688 , \45689 , \45690 , \45691 , \45692 , \45693 , \45694 ,
         \45695 , \45696 , \45697 , \45698 , \45699 , \45700 , \45701 , \45702 , \45703_nR235c2 , \45704 ,
         \45705 , \45706 , \45707 , \45708 , \45709 , \45710 , \45711 , \45712 , \45713 , \45714 ,
         \45715 , \45716 , \45717 , \45718 , \45719 , \45720 , \45721_nR235c4 , \45722 , \45723 , \45724 ,
         \45725 , \45726 , \45727 , \45728 , \45729 , \45730 , \45731 , \45732 , \45733 , \45734 ,
         \45735 , \45736 , \45737 , \45738 , \45739_nR235c6 , \45740 , \45741 , \45742 , \45743 , \45744 ,
         \45745 , \45746 , \45747 , \45748 , \45749 , \45750 , \45751 , \45752 , \45753 , \45754 ,
         \45755 , \45756 , \45757_nR235c8 , \45758 , \45759 , \45760 , \45761 , \45762 , \45763 , \45764 ,
         \45765 , \45766 , \45767 , \45768 , \45769 , \45770 , \45771 , \45772 , \45773 , \45774 ,
         \45775_nR235cc , \45776 , \45777 , \45778 , \45779 , \45780 , \45781 , \45782 , \45783 , \45784 ,
         \45785 , \45786 , \45787 , \45788 , \45789 , \45790 , \45791 , \45792 , \45793_nR235ce , \45794 ,
         \45795 , \45796 , \45797 , \45798 , \45799 , \45800 , \45801 , \45802 , \45803 , \45804 ,
         \45805 , \45806 , \45807 , \45808 , \45809 , \45810 , \45811_nR235d0 , \45812 , \45813 , \45814 ,
         \45815 , \45816 , \45817 , \45818 , \45819 , \45820 , \45821 , \45822 , \45823 , \45824 ,
         \45825 , \45826 , \45827 , \45828 , \45829_nR235d2 , \45830 , \45831 , \45832 , \45833 , \45834 ,
         \45835 , \45836 , \45837 , \45838 , \45839 , \45840 , \45841 , \45842 , \45843 , \45844 ,
         \45845 , \45846 , \45847 , \45848 , \45849 , \45850 , \45851 , \45852 , \45853 , \45854 ,
         \45855 , \45856 , \45857 , \45858 , \45859 , \45860 , \45861 , \45862_nR235dc , \45863 , \45864 ,
         \45865 , \45866 , \45867 , \45868 , \45869 , \45870 , \45871 , \45872 , \45873 , \45874 ,
         \45875 , \45876 , \45877 , \45878 , \45879 , \45880 , \45881_nR235f2 , \45882 , \45883 , \45884 ,
         \45885 , \45886 , \45887 , \45888 , \45889 , \45890 , \45891 , \45892 , \45893 , \45894 ,
         \45895 , \45896 , \45897 , \45898_nR23608 , \45899 , \45900 , \45901 , \45902 , \45903 , \45904 ,
         \45905 , \45906 , \45907 , \45908 , \45909 , \45910 , \45911 , \45912 , \45913 , \45914 ,
         \45915 , \45916_nR2361e , \45917 , \45918 , \45919 , \45920 , \45921 , \45922 , \45923 , \45924 ,
         \45925 , \45926 , \45927 , \45928 , \45929 , \45930 , \45931 , \45932 , \45933 , \45934_nR23634 ,
         \45935 , \45936 , \45937 , \45938 , \45939 , \45940 , \45941 , \45942 , \45943 , \45944 ,
         \45945 , \45946 , \45947 , \45948 , \45949 , \45950 , \45951 , \45952 , \45953_nR2364a , \45954 ,
         \45955 , \45956 , \45957 , \45958 , \45959 , \45960 , \45961 , \45962 , \45963 , \45964 ,
         \45965 , \45966 , \45967 , \45968 , \45969 , \45970 , \45971_nR23654 , \45972 , \45973 , \45974 ,
         \45975 , \45976 , \45977 , \45978 , \45979 , \45980 , \45981 , \45982 , \45983 , \45984 ,
         \45985 , \45986 , \45987 , \45988 , \45989_nR23656 , \45990 , \45991 , \45992 , \45993 , \45994 ,
         \45995 , \45996 , \45997 , \45998 , \45999 , \46000 , \46001 , \46002 , \46003 , \46004 ,
         \46005 , \46006_nR23658 , \46007 , \46008 , \46009 , \46010 , \46011 , \46012 , \46013 , \46014 ,
         \46015 , \46016 , \46017 , \46018 , \46019 , \46020 , \46021 , \46022 , \46023 , \46024 ,
         \46025_nR2365a , \46026 , \46027 , \46028 , \46029 , \46030 , \46031 , \46032 , \46033 , \46034 ,
         \46035 , \46036 , \46037 , \46038 , \46039 , \46040 , \46041 , \46042_nR235de , \46043 , \46044 ,
         \46045 , \46046 , \46047 , \46048 , \46049 , \46050 , \46051 , \46052 , \46053 , \46054 ,
         \46055 , \46056 , \46057 , \46058 , \46059 , \46060 , \46061_nR235e0 , \46062 , \46063 , \46064 ,
         \46065 , \46066 , \46067 , \46068 , \46069 , \46070 , \46071 , \46072 , \46073 , \46074 ,
         \46075 , \46076 , \46077 , \46078 , \46079_nR235e2 , \46080 , \46081 , \46082 , \46083 , \46084 ,
         \46085 , \46086 , \46087 , \46088 , \46089 , \46090 , \46091 , \46092 , \46093 , \46094 ,
         \46095 , \46096 , \46097_nR235e4 , \46098 , \46099 , \46100 , \46101 , \46102 , \46103 , \46104 ,
         \46105 , \46106 , \46107 , \46108 , \46109 , \46110 , \46111 , \46112 , \46113 , \46114_nR235e6 ,
         \46115 , \46116 , \46117 , \46118 , \46119 , \46120 , \46121 , \46122 , \46123 , \46124 ,
         \46125 , \46126 , \46127 , \46128 , \46129 , \46130 , \46131_nR235e8 , \46132 , \46133 , \46134 ,
         \46135 , \46136 , \46137 , \46138 , \46139 , \46140 , \46141 , \46142 , \46143 , \46144 ,
         \46145 , \46146 , \46147 , \46148_nR235ea , \46149 , \46150 , \46151 , \46152 , \46153 , \46154 ,
         \46155 , \46156 , \46157 , \46158 , \46159 , \46160 , \46161 , \46162 , \46163 , \46164 ,
         \46165_nR235ec , \46166 , \46167 , \46168 , \46169 , \46170 , \46171 , \46172 , \46173 , \46174 ,
         \46175 , \46176 , \46177 , \46178 , \46179 , \46180 , \46181 , \46182_nR235ee , \46183 , \46184 ,
         \46185 , \46186 , \46187 , \46188 , \46189 , \46190 , \46191 , \46192 , \46193 , \46194 ,
         \46195 , \46196 , \46197 , \46198 , \46199_nR235f0 , \46200 , \46201 , \46202 , \46203 , \46204 ,
         \46205 , \46206 , \46207 , \46208 , \46209 , \46210 , \46211 , \46212 , \46213 , \46214 ,
         \46215 , \46216_nR235f4 , \46217 , \46218 , \46219 , \46220 , \46221 , \46222 , \46223 , \46224 ,
         \46225 , \46226 , \46227 , \46228 , \46229 , \46230 , \46231 , \46232 , \46233_nR235f6 , \46234 ,
         \46235 , \46236 , \46237 , \46238 , \46239 , \46240 , \46241 , \46242 , \46243 , \46244 ,
         \46245 , \46246 , \46247 , \46248 , \46249 , \46250 , \46251_nR235f8 , \46252 , \46253 , \46254 ,
         \46255 , \46256 , \46257 , \46258 , \46259 , \46260 , \46261 , \46262 , \46263 , \46264 ,
         \46265 , \46266 , \46267 , \46268_nR235fa , \46269 , \46270 , \46271 , \46272 , \46273 , \46274 ,
         \46275 , \46276 , \46277 , \46278 , \46279 , \46280 , \46281 , \46282 , \46283 , \46284 ,
         \46285_nR235fc , \46286 , \46287 , \46288 , \46289 , \46290 , \46291 , \46292 , \46293 , \46294 ,
         \46295 , \46296 , \46297 , \46298 , \46299 , \46300 , \46301 , \46302_nR235fe , \46303 , \46304 ,
         \46305 , \46306 , \46307 , \46308 , \46309 , \46310 , \46311 , \46312 , \46313 , \46314 ,
         \46315 , \46316 , \46317 , \46318 , \46319_nR23600 , \46320 , \46321 , \46322 , \46323 , \46324 ,
         \46325 , \46326 , \46327 , \46328 , \46329 , \46330 , \46331 , \46332 , \46333 , \46334 ,
         \46335 , \46336_nR23602 , \46337 , \46338 , \46339 , \46340 , \46341 , \46342 , \46343 , \46344 ,
         \46345 , \46346 , \46347 , \46348 , \46349 , \46350 , \46351 , \46352 , \46353_nR23604 , \46354 ,
         \46355 , \46356 , \46357 , \46358 , \46359 , \46360 , \46361 , \46362 , \46363 , \46364 ,
         \46365 , \46366 , \46367 , \46368 , \46369 , \46370_nR23606 , \46371 , \46372 , \46373 , \46374 ,
         \46375 , \46376 , \46377 , \46378 , \46379 , \46380 , \46381 , \46382 , \46383 , \46384 ,
         \46385 , \46386 , \46387_nR2360a , \46388 ;
buf \U$labaj4975 ( R_25610_96cc360, \21946 );
buf \U$labaj4976 ( R_25642_95f0d48, \21951 );
buf \U$labaj4977 ( R_25644_9598060, \21956 );
buf \U$labaj4978 ( R_25646_95984f8, \21962 );
buf \U$labaj4979 ( R_25614_953c348, \21968 );
buf \U$labaj4980 ( R_25616_96251f8, \21979 );
buf \U$labaj4981 ( R_25618_96ed6b0, \21989 );
buf \U$labaj4982 ( R_2561a_95f00d0, \21999 );
buf \U$labaj4983 ( R_2561c_95f0418, \22009 );
buf \U$labaj4984 ( R_2561e_95f0760, \22019 );
buf \U$labaj4985 ( R_25620_953c3f0, \22029 );
buf \U$labaj4986 ( R_25622_953c690, \22039 );
buf \U$labaj4987 ( R_25612_953c9d8, \22049 );
buf \U$labaj4988 ( R_25624_95f08b0, \22059 );
buf \U$labaj4989 ( R_25626_953ca80, \22069 );
buf \U$labaj4990 ( R_25628_96253f0, \22079 );
buf \U$labaj4991 ( R_2562a_9632be8, \22089 );
buf \U$labaj4992 ( R_253fc_9d20ef0, \22146 );
buf \U$labaj4993 ( R_25412_9530108, \22174 );
buf \U$labaj4994 ( R_25428_95f75a0, \22194 );
buf \U$labaj4995 ( R_2543e_95301b0, \22217 );
buf \U$labaj4996 ( R_25454_95304f8, \22238 );
buf \U$labaj4997 ( R_2546a_9533198, \22265 );
buf \U$labaj4998 ( R_25474_95332e8, \22286 );
buf \U$labaj4999 ( R_25476_96dee60, \22307 );
buf \U$labaj5000 ( R_25478_95f7798, \22329 );
buf \U$labaj5001 ( R_2547a_96def08, \22350 );
buf \U$labaj5002 ( R_253fe_95f7990, \22371 );
buf \U$labaj5003 ( R_25400_9d21190, \22391 );
buf \U$labaj5004 ( R_25402_9d21388, \22412 );
buf \U$labaj5005 ( R_25404_9589e90, \22433 );
buf \U$labaj5006 ( R_25406_9d21430, \22452 );
buf \U$labaj5007 ( R_25408_9533780, \22472 );
buf \U$labaj5008 ( R_2540a_9533b70, \22492 );
buf \U$labaj5009 ( R_2540c_9d216d0, \22513 );
buf \U$labaj5010 ( R_2540e_958a5c8, \22533 );
buf \U$labaj5011 ( R_25410_96defb0, \22553 );
buf \U$labaj5012 ( R_25414_9d21778, \22573 );
buf \U$labaj5013 ( R_25416_9d21cb8, \22593 );
buf \U$labaj5014 ( R_25418_95f7ae0, \22613 );
buf \U$labaj5015 ( R_2541a_9d21d60, \22633 );
buf \U$labaj5016 ( R_2541c_96df100, \22654 );
buf \U$labaj5017 ( R_2541e_9d221f8, \22674 );
buf \U$labaj5018 ( R_25420_958ac58, \22695 );
buf \U$labaj5019 ( R_25422_95f7b88, \22715 );
buf \U$labaj5020 ( R_25424_9533c18, \22735 );
buf \U$labaj5021 ( R_25426_958b630, \22755 );
buf \U$labaj5022 ( R_2542a_9d222a0, \22777 );
buf \U$labaj5023 ( R_2542c_9533d68, \22797 );
buf \U$labaj5024 ( R_2542e_95f7c30, \22817 );
buf \U$labaj5025 ( R_25430_9d22498, \22837 );
buf \U$labaj5026 ( R_25432_9d22540, \22857 );
buf \U$labaj5027 ( R_25434_9533f60, \22877 );
buf \U$labaj5028 ( R_25436_96df1a8, \22897 );
buf \U$labaj5029 ( R_25438_95f7f78, \22919 );
buf \U$labaj5030 ( R_2543a_9534008, \22939 );
buf \U$labaj5031 ( R_2543c_9534200, \22959 );
buf \U$labaj5032 ( R_25440_95f80c8, \22979 );
buf \U$labaj5033 ( R_25442_96df250, \22998 );
buf \U$labaj5034 ( R_25444_9d22690, \23017 );
buf \U$labaj5035 ( R_25446_95fa438, \23037 );
buf \U$labaj5036 ( R_25448_95fa4e0, \23059 );
buf \U$labaj5037 ( R_2544a_958bcc0, \23079 );
buf \U$labaj5038 ( R_2544c_9d22738, \23099 );
buf \U$labaj5039 ( R_2544e_9d227e0, \23119 );
buf \U$labaj5040 ( R_25450_9d22888, \23139 );
buf \U$labaj5041 ( R_25452_9d22930, \23159 );
buf \U$labaj5042 ( R_25456_9d229d8, \23179 );
buf \U$labaj5043 ( R_25458_95fa588, \23198 );
buf \U$labaj5044 ( R_2545a_9534350, \23218 );
buf \U$labaj5045 ( R_2545c_95fa828, \23238 );
buf \U$labaj5046 ( R_2545e_9d22a80, \23258 );
buf \U$labaj5047 ( R_25460_96df2f8, \23278 );
buf \U$labaj5048 ( R_25462_96df3a0, \23298 );
buf \U$labaj5049 ( R_25464_95343f8, \23317 );
buf \U$labaj5050 ( R_25466_95fa8d0, \23337 );
buf \U$labaj5051 ( R_25468_95faac8, \23357 );
buf \U$labaj5052 ( R_2546c_958bd68, \23378 );
buf \U$labaj5053 ( R_2546e_958be10, \23398 );
buf \U$labaj5054 ( R_25470_95fab70, \23418 );
buf \U$labaj5055 ( R_25472_9d22b28, \23438 );
buf \U$labaj5056 ( R_2547c_958beb8, \23472 );
buf \U$labaj5057 ( R_25492_9d22bd0, \23492 );
buf \U$labaj5058 ( R_254a8_958bf60, \23510 );
buf \U$labaj5059 ( R_254be_9d22c78, \23528 );
buf \U$labaj5060 ( R_254d4_9d22dc8, \23548 );
buf \U$labaj5061 ( R_254ea_9d22e70, \23569 );
buf \U$labaj5062 ( R_254f4_958c0b0, \23587 );
buf \U$labaj5063 ( R_254f6_9d22f18, \23606 );
buf \U$labaj5064 ( R_254f8_958c158, \23624 );
buf \U$labaj5065 ( R_254fa_9d22fc0, \23644 );
buf \U$labaj5066 ( R_2547e_958c200, \23663 );
buf \U$labaj5067 ( R_25480_9d23068, \23681 );
buf \U$labaj5068 ( R_25482_9d231b8, \23700 );
buf \U$labaj5069 ( R_25484_958c2a8, \23718 );
buf \U$labaj5070 ( R_25486_958c350, \23736 );
buf \U$labaj5071 ( R_25488_9d23458, \23754 );
buf \U$labaj5072 ( R_2548a_958c4a0, \23773 );
buf \U$labaj5073 ( R_2548c_9d235a8, \23791 );
buf \U$labaj5074 ( R_2548e_9d236f8, \23809 );
buf \U$labaj5075 ( R_25490_958c548, \23827 );
buf \U$labaj5076 ( R_25494_958c5f0, \23845 );
buf \U$labaj5077 ( R_25496_9d237a0, \23863 );
buf \U$labaj5078 ( R_25498_958c698, \23881 );
buf \U$labaj5079 ( R_2549a_958f728, \23899 );
buf \U$labaj5080 ( R_2549c_9d23848, \23917 );
buf \U$labaj5081 ( R_2549e_958f7d0, \23935 );
buf \U$labaj5082 ( R_254a0_958f878, \23954 );
buf \U$labaj5083 ( R_254a2_9d23998, \23972 );
buf \U$labaj5084 ( R_254a4_9d23ae8, \23990 );
buf \U$labaj5085 ( R_254a6_9d23c38, \24008 );
buf \U$labaj5086 ( R_254aa_9d23d88, \24026 );
buf \U$labaj5087 ( R_254ac_9d23e30, \24044 );
buf \U$labaj5088 ( R_254ae_9d23f80, \24062 );
buf \U$labaj5089 ( R_254b0_9d24028, \24080 );
buf \U$labaj5090 ( R_254b2_9d240d0, \24098 );
buf \U$labaj5091 ( R_254b4_9d24220, \24116 );
buf \U$labaj5092 ( R_254b6_9d242c8, \24136 );
buf \U$labaj5093 ( R_254b8_9590988, \24154 );
buf \U$labaj5094 ( R_254ba_9590a30, \24174 );
buf \U$labaj5095 ( R_254bc_9590cd0, \24192 );
buf \U$labaj5096 ( R_254c0_9d24418, \24210 );
buf \U$labaj5097 ( R_254c2_9590d78, \24228 );
buf \U$labaj5098 ( R_254c4_9590f70, \24246 );
buf \U$labaj5099 ( R_254c6_9591178, \24264 );
buf \U$labaj5100 ( R_254c8_9d24568, \24282 );
buf \U$labaj5101 ( R_254ca_9d24bf8, \24300 );
buf \U$labaj5102 ( R_254cc_9d25090, \24318 );
buf \U$labaj5103 ( R_254ce_95916b8, \24336 );
buf \U$labaj5104 ( R_254d0_9591808, \24354 );
buf \U$labaj5105 ( R_254d2_9d251e0, \24372 );
buf \U$labaj5106 ( R_254d6_9d25f10, \24390 );
buf \U$labaj5107 ( R_254d8_9d25fb8, \24408 );
buf \U$labaj5108 ( R_254da_95918b0, \24427 );
buf \U$labaj5109 ( R_254dc_9d265a0, \24445 );
buf \U$labaj5110 ( R_254de_9591958, \24463 );
buf \U$labaj5111 ( R_254e0_9d26990, \24481 );
buf \U$labaj5112 ( R_254e2_9d26c30, \24499 );
buf \U$labaj5113 ( R_254e4_9591a00, \24517 );
buf \U$labaj5114 ( R_254e6_95347e8, \24535 );
buf \U$labaj5115 ( R_254e8_9591b50, \24553 );
buf \U$labaj5116 ( R_254ec_9591bf8, \24571 );
buf \U$labaj5117 ( R_254ee_9d26d80, \24589 );
buf \U$labaj5118 ( R_254f0_9d27368, \24607 );
buf \U$labaj5119 ( R_254f2_9d27410, \24625 );
buf \U$labaj5120 ( R_254fc_96df4f0, \24657 );
buf \U$labaj5121 ( R_25512_9d276b0, \24676 );
buf \U$labaj5122 ( R_25528_96df598, \24693 );
buf \U$labaj5123 ( R_2553e_9534890, \24711 );
buf \U$labaj5124 ( R_25554_9d27c98, \24730 );
buf \U$labaj5125 ( R_2556a_96df640, \24748 );
buf \U$labaj5126 ( R_25574_9d27de8, \24765 );
buf \U$labaj5127 ( R_25576_96df6e8, \24782 );
buf \U$labaj5128 ( R_25578_9534bd8, \24799 );
buf \U$labaj5129 ( R_2557a_96df838, \24817 );
buf \U$labaj5130 ( R_254fe_96dfad8, \24835 );
buf \U$labaj5131 ( R_25500_9534d28, \24852 );
buf \U$labaj5132 ( R_25502_9534dd0, \24869 );
buf \U$labaj5133 ( R_25504_9534f20, \24886 );
buf \U$labaj5134 ( R_25506_9d281d8, \24903 );
buf \U$labaj5135 ( R_25508_96dfb80, \24921 );
buf \U$labaj5136 ( R_2550a_9d28328, \24938 );
buf \U$labaj5137 ( R_2550c_9d283d0, \24955 );
buf \U$labaj5138 ( R_2550e_96dfc28, \24972 );
buf \U$labaj5139 ( R_25510_9534fc8, \24989 );
buf \U$labaj5140 ( R_25514_96dfcd0, \25006 );
buf \U$labaj5141 ( R_25516_9d28520, \25023 );
buf \U$labaj5142 ( R_25518_96dfe20, \25040 );
buf \U$labaj5143 ( R_2551a_96dfec8, \25057 );
buf \U$labaj5144 ( R_2551c_9535070, \25074 );
buf \U$labaj5145 ( R_2551e_95351c0, \25091 );
buf \U$labaj5146 ( R_25520_9535268, \25108 );
buf \U$labaj5147 ( R_25522_96dff70, \25125 );
buf \U$labaj5148 ( R_25524_96e0018, \25142 );
buf \U$labaj5149 ( R_25526_96e00c0, \25159 );
buf \U$labaj5150 ( R_2552a_9535310, \25176 );
buf \U$labaj5151 ( R_2552c_96e0168, \25193 );
buf \U$labaj5152 ( R_2552e_96e0210, \25210 );
buf \U$labaj5153 ( R_25530_96e02b8, \25227 );
buf \U$labaj5154 ( R_25532_96e0408, \25244 );
buf \U$labaj5155 ( R_25534_96e0558, \25261 );
buf \U$labaj5156 ( R_25536_96e0600, \25278 );
buf \U$labaj5157 ( R_25538_9535658, \25295 );
buf \U$labaj5158 ( R_2553a_9d289b8, \25312 );
buf \U$labaj5159 ( R_2553c_96e06a8, \25329 );
buf \U$labaj5160 ( R_25540_95358f8, \25346 );
buf \U$labaj5161 ( R_25542_96e0750, \25363 );
buf \U$labaj5162 ( R_25544_96e0b40, \25380 );
buf \U$labaj5163 ( R_25546_96e0be8, \25397 );
buf \U$labaj5164 ( R_25548_96e0c90, \25414 );
buf \U$labaj5165 ( R_2554a_96e0d38, \25431 );
buf \U$labaj5166 ( R_2554c_95359a0, \25448 );
buf \U$labaj5167 ( R_2554e_9d28a60, \25466 );
buf \U$labaj5168 ( R_25550_96e0e88, \25483 );
buf \U$labaj5169 ( R_25552_9535a48, \25500 );
buf \U$labaj5170 ( R_25556_96e0f30, \25517 );
buf \U$labaj5171 ( R_25558_9535b98, \25534 );
buf \U$labaj5172 ( R_2555a_9d28c58, \25551 );
buf \U$labaj5173 ( R_2555c_96e0fd8, \25568 );
buf \U$labaj5174 ( R_2555e_9d28d00, \25585 );
buf \U$labaj5175 ( R_25560_9535c40, \25602 );
buf \U$labaj5176 ( R_25562_95362d0, \25619 );
buf \U$labaj5177 ( R_25564_9536810, \25636 );
buf \U$labaj5178 ( R_25566_9536a08, \25654 );
buf \U$labaj5179 ( R_25568_96e1080, \25671 );
buf \U$labaj5180 ( R_2556c_96e1128, \25688 );
buf \U$labaj5181 ( R_2556e_9d28ef8, \25705 );
buf \U$labaj5182 ( R_25570_96e11d0, \25722 );
buf \U$labaj5183 ( R_25572_96e1c50, \25739 );
buf \U$labaj5184 ( R_2557c_9591d48, \25766 );
buf \U$labaj5185 ( R_25592_9591df0, \25782 );
buf \U$labaj5186 ( R_255a8_96e2e08, \25799 );
buf \U$labaj5187 ( R_255be_9591e98, \25815 );
buf \U$labaj5188 ( R_255d4_9591f40, \25829 );
buf \U$labaj5189 ( R_255ea_96e3690, \25844 );
buf \U$labaj5190 ( R_255f4_96e6918, \25858 );
buf \U$labaj5191 ( R_255f6_96e69c0, \25872 );
buf \U$labaj5192 ( R_255f8_9d29048, \25886 );
buf \U$labaj5193 ( R_255fa_9d28718, \25901 );
buf \U$labaj5194 ( R_2557e_9591fe8, \25915 );
buf \U$labaj5195 ( R_25580_96e6fa8, \25929 );
buf \U$labaj5196 ( R_25582_96e72f0, \25943 );
buf \U$labaj5197 ( R_25584_9d287c0, \25957 );
buf \U$labaj5198 ( R_25586_9592090, \25971 );
buf \U$labaj5199 ( R_25588_9592138, \25985 );
buf \U$labaj5200 ( R_2558a_96e7398, \25999 );
buf \U$labaj5201 ( R_2558c_9d28868, \26013 );
buf \U$labaj5202 ( R_2558e_9d290f0, \26027 );
buf \U$labaj5203 ( R_25590_9d29240, \26042 );
buf \U$labaj5204 ( R_25594_96e7cc8, \26056 );
buf \U$labaj5205 ( R_25596_95921e0, \26070 );
buf \U$labaj5206 ( R_25598_9592288, \26084 );
buf \U$labaj5207 ( R_2559a_9592330, \26098 );
buf \U$labaj5208 ( R_2559c_96e82b0, \26112 );
buf \U$labaj5209 ( R_2559e_9d292e8, \26126 );
buf \U$labaj5210 ( R_255a0_9d2dfb0, \26140 );
buf \U$labaj5211 ( R_255a2_9592528, \26154 );
buf \U$labaj5212 ( R_255a4_9592678, \26168 );
buf \U$labaj5213 ( R_255a6_9d2e058, \26182 );
buf \U$labaj5214 ( R_255aa_96e8358, \26197 );
buf \U$labaj5215 ( R_255ac_9592918, \26211 );
buf \U$labaj5216 ( R_255ae_96e86a0, \26225 );
buf \U$labaj5217 ( R_255b0_9d2e988, \26239 );
buf \U$labaj5218 ( R_255b2_9d29390, \26253 );
buf \U$labaj5219 ( R_255b4_9d2ec28, \26267 );
buf \U$labaj5220 ( R_255b6_9d294e0, \26281 );
buf \U$labaj5221 ( R_255b8_9d2f360, \26295 );
buf \U$labaj5222 ( R_255ba_9592a68, \26309 );
buf \U$labaj5223 ( R_255bc_9592b10, \26323 );
buf \U$labaj5224 ( R_255c0_9d30128, \26337 );
buf \U$labaj5225 ( R_255c2_9592c60, \26351 );
buf \U$labaj5226 ( R_255c4_96e8940, \26365 );
buf \U$labaj5227 ( R_255c6_96e89e8, \26379 );
buf \U$labaj5228 ( R_255c8_9d30278, \26393 );
buf \U$labaj5229 ( R_255ca_96e8be0, \26407 );
buf \U$labaj5230 ( R_255cc_9592f00, \26421 );
buf \U$labaj5231 ( R_255ce_9d29588, \26435 );
buf \U$labaj5232 ( R_255d0_9d296d8, \26449 );
buf \U$labaj5233 ( R_255d2_9d30518, \26463 );
buf \U$labaj5234 ( R_255d6_9d29828, \26477 );
buf \U$labaj5235 ( R_255d8_96e9120, \26491 );
buf \U$labaj5236 ( R_255da_96e93c0, \26505 );
buf \U$labaj5237 ( R_255dc_96e9510, \26519 );
buf \U$labaj5238 ( R_255de_9d307b8, \26533 );
buf \U$labaj5239 ( R_255e0_9d29cc0, \26547 );
buf \U$labaj5240 ( R_255e2_9592fa8, \26561 );
buf \U$labaj5241 ( R_255e4_9593050, \26575 );
buf \U$labaj5242 ( R_255e6_96e9858, \26589 );
buf \U$labaj5243 ( R_255e8_96e9a50, \26603 );
buf \U$labaj5244 ( R_255ec_95930f8, \26617 );
buf \U$labaj5245 ( R_255ee_9d29eb8, \26631 );
buf \U$labaj5246 ( R_255f0_96ea038, \26645 );
buf \U$labaj5247 ( R_255f2_95931a0, \26659 );
buf \U$labaj5248 ( R_253bc_96eacb0, \26678 );
buf \U$labaj5249 ( R_253be_9593248, \26696 );
buf \U$labaj5250 ( R_253c0_9d29f60, \26713 );
buf \U$labaj5251 ( R_253c2_95932f0, \26730 );
buf \U$labaj5252 ( R_253c4_96eae00, \26747 );
buf \U$labaj5253 ( R_253c6_9536b58, \26764 );
buf \U$labaj5254 ( R_253c8_9593398, \26781 );
buf \U$labaj5255 ( R_253ca_9d2a350, \26798 );
buf \U$labaj5256 ( R_253cc_b7dc210, \26813 );
buf \U$labaj5257 ( R_253ce_b7dcd38, \26828 );
buf \U$labaj5258 ( R_253d0_b7dcde0, \26843 );
buf \U$labaj5259 ( R_253d2_9593590, \26858 );
buf \U$labaj5260 ( R_253d4_96376b8, \26873 );
buf \U$labaj5261 ( R_253d6_9d2a4a0, \26888 );
buf \U$labaj5262 ( R_253d8_9596038, \26903 );
buf \U$labaj5263 ( R_253da_b7dc2b8, \26918 );
buf \U$labaj5264 ( R_253dc_96eb0a0, \26933 );
buf \U$labaj5265 ( R_253de_9596578, \26948 );
buf \U$labaj5266 ( R_253e0_9536f48, \26963 );
buf \U$labaj5267 ( R_253e2_96eb298, \26978 );
buf \U$labaj5268 ( R_253e4_9537098, \26993 );
buf \U$labaj5269 ( R_253e6_96eb340, \27008 );
buf \U$labaj5270 ( R_253e8_95373e0, \27023 );
buf \U$labaj5271 ( R_253ea_9596a10, \27038 );
buf \U$labaj5272 ( R_253ec_9d30860, \27053 );
buf \U$labaj5273 ( R_253ee_9ef0090, \27068 );
buf \U$labaj5274 ( R_253f0_9d30f98, \27083 );
buf \U$labaj5275 ( R_253f2_9ef05d0, \27098 );
buf \U$labaj5276 ( R_253f4_9d31040, \27113 );
buf \U$labaj5277 ( R_253f6_9d31238, \27128 );
buf \U$labaj5278 ( R_253f8_9d314d8, \27143 );
buf \U$labaj5279 ( R_253fa_9d316d0, \27158 );
buf \U$labaj5280 ( R_25666_96346d0, \27175 );
buf \U$labaj5281 ( R_1a4_b821b50, \27280 );
buf \U$labaj5282 ( R_1a3_b821aa8, \27345 );
buf \U$labaj5283 ( R_23ca4_96329f0, \27411 );
buf \U$labaj5284 ( R_23cba_9f596e0, \27439 );
buf \U$labaj5285 ( R_23cd0_962b7c0, \27457 );
buf \U$labaj5286 ( R_23ce6_955f268, \27478 );
buf \U$labaj5287 ( R_23cfc_9f5c4d0, \27498 );
buf \U$labaj5288 ( R_23d12_9d225e8, \27519 );
buf \U$labaj5289 ( R_23d1c_962b910, \27538 );
buf \U$labaj5290 ( R_23d1e_95a3470, \27557 );
buf \U$labaj5291 ( R_23d20_9632c90, \27579 );
buf \U$labaj5292 ( R_23d22_95a3710, \27600 );
buf \U$labaj5293 ( R_23ca6_9ee76c0, \27620 );
buf \U$labaj5294 ( R_23ca8_9ee7810, \27639 );
buf \U$labaj5295 ( R_23caa_9ee78b8, \27659 );
buf \U$labaj5296 ( R_23cac_9ee8140, \27679 );
buf \U$labaj5297 ( R_23cae_962bbb0, \27697 );
buf \U$labaj5298 ( R_23cb0_9ee8920, \27715 );
buf \U$labaj5299 ( R_23cb2_9d22d20, \27733 );
buf \U$labaj5300 ( R_23cb4_9ee8bc0, \27752 );
buf \U$labaj5301 ( R_23cb6_9632d38, \27771 );
buf \U$labaj5302 ( R_23cb8_9d23110, \27790 );
buf \U$labaj5303 ( R_23cbc_962bc58, \27810 );
buf \U$labaj5304 ( R_23cbe_9ee9ad8, \27828 );
buf \U$labaj5305 ( R_23cc0_9d23260, \27846 );
buf \U$labaj5306 ( R_23cc2_9632f30, \27865 );
buf \U$labaj5307 ( R_23cc4_9eec430, \27884 );
buf \U$labaj5308 ( R_23cc6_9d23308, \27903 );
buf \U$labaj5309 ( R_23cc8_9eef4c0, \27922 );
buf \U$labaj5310 ( R_23cca_9eefca0, \27941 );
buf \U$labaj5311 ( R_23ccc_9d23650, \27960 );
buf \U$labaj5312 ( R_23cce_9ef0678, \27979 );
buf \U$labaj5313 ( R_23cd2_95a3908, \27999 );
buf \U$labaj5314 ( R_23cd4_962bd00, \28020 );
buf \U$labaj5315 ( R_23cd6_9632fd8, \28040 );
buf \U$labaj5316 ( R_23cd8_962be50, \28059 );
buf \U$labaj5317 ( R_23cda_96331d0, \28077 );
buf \U$labaj5318 ( R_23cdc_962bef8, \28096 );
buf \U$labaj5319 ( R_23cde_9d30ef0, \28115 );
buf \U$labaj5320 ( R_23ce0_9d238f0, \28134 );
buf \U$labaj5321 ( R_23ce2_9d23b90, \28153 );
buf \U$labaj5322 ( R_23ce4_962bfa0, \28172 );
buf \U$labaj5323 ( R_23ce8_962c048, \28191 );
buf \U$labaj5324 ( R_23cea_95a3a58, \28210 );
buf \U$labaj5325 ( R_23cec_9d23ed8, \28229 );
buf \U$labaj5326 ( R_23cee_9ef09c0, \28248 );
buf \U$labaj5327 ( R_23cf0_9ef4380, \28268 );
buf \U$labaj5328 ( R_23cf2_95a3ba8, \28287 );
buf \U$labaj5329 ( R_23cf4_9ef4a10, \28306 );
buf \U$labaj5330 ( R_23cf6_962c0f0, \28325 );
buf \U$labaj5331 ( R_23cf8_96c3060, \28344 );
buf \U$labaj5332 ( R_23cfa_96c6d68, \28363 );
buf \U$labaj5333 ( R_23cfe_9d310e8, \28383 );
buf \U$labaj5334 ( R_23d00_96c72a8, \28403 );
buf \U$labaj5335 ( R_23d02_962c390, \28423 );
buf \U$labaj5336 ( R_23d04_96c74a0, \28443 );
buf \U$labaj5337 ( R_23d06_962da88, \28463 );
buf \U$labaj5338 ( R_23d08_9d24178, \28482 );
buf \U$labaj5339 ( R_23d0a_962df20, \28501 );
buf \U$labaj5340 ( R_23d0c_9633278, \28521 );
buf \U$labaj5341 ( R_23d0e_9633320, \28540 );
buf \U$labaj5342 ( R_23d10_95a3e48, \28562 );
buf \U$labaj5343 ( R_23d14_95a4040, \28582 );
buf \U$labaj5344 ( R_23d16_9d24370, \28600 );
buf \U$labaj5345 ( R_23d18_96c7e78, \28619 );
buf \U$labaj5346 ( R_23d1a_96333c8, \28637 );
buf \U$labaj5347 ( R_23d24_9633470, \28669 );
buf \U$labaj5348 ( R_23d3a_9633518, \28690 );
buf \U$labaj5349 ( R_23d50_962dfc8, \28709 );
buf \U$labaj5350 ( R_23d66_9629b88, \28729 );
buf \U$labaj5351 ( R_23d7c_95547c8, \28748 );
buf \U$labaj5352 ( R_23d92_96335c0, \28768 );
buf \U$labaj5353 ( R_23d9c_96337b8, \28787 );
buf \U$labaj5354 ( R_23d9e_9633908, \28805 );
buf \U$labaj5355 ( R_23da0_9633a58, \28823 );
buf \U$labaj5356 ( R_23da2_962e7a8, \28839 );
buf \U$labaj5357 ( R_23d26_9554870, \28856 );
buf \U$labaj5358 ( R_23d28_962a560, \28872 );
buf \U$labaj5359 ( R_23d2a_962ee38, \28888 );
buf \U$labaj5360 ( R_23d2c_962a8a8, \28905 );
buf \U$labaj5361 ( R_23d2e_962f2d0, \28921 );
buf \U$labaj5362 ( R_23d30_95549c0, \28938 );
buf \U$labaj5363 ( R_23d32_9633cf8, \28955 );
buf \U$labaj5364 ( R_23d34_962f4c8, \28971 );
buf \U$labaj5365 ( R_23d36_9633da0, \28987 );
buf \U$labaj5366 ( R_23d38_9633e48, \29005 );
buf \U$labaj5367 ( R_23d3c_9633ef0, \29023 );
buf \U$labaj5368 ( R_23d3e_962c4e0, \29041 );
buf \U$labaj5369 ( R_23d40_9554bb8, \29059 );
buf \U$labaj5370 ( R_23d42_9554d08, \29077 );
buf \U$labaj5371 ( R_23d44_9634040, \29095 );
buf \U$labaj5372 ( R_23d46_962f6c0, \29113 );
buf \U$labaj5373 ( R_23d48_9554f00, \29131 );
buf \U$labaj5374 ( R_23d4a_962c8d0, \29149 );
buf \U$labaj5375 ( R_23d4c_9635000, \29167 );
buf \U$labaj5376 ( R_23d4e_962fab0, \29185 );
buf \U$labaj5377 ( R_23d52_95552f0, \29203 );
buf \U$labaj5378 ( R_23d54_96350a8, \29221 );
buf \U$labaj5379 ( R_23d56_96351f8, \29239 );
buf \U$labaj5380 ( R_23d58_962fc00, \29257 );
buf \U$labaj5381 ( R_23d5a_95554e8, \29275 );
buf \U$labaj5382 ( R_23d5c_9555638, \29293 );
buf \U$labaj5383 ( R_23d5e_9635540, \29312 );
buf \U$labaj5384 ( R_23d60_96355e8, \29328 );
buf \U$labaj5385 ( R_23d62_9635738, \29346 );
buf \U$labaj5386 ( R_23d64_96359d8, \29362 );
buf \U$labaj5387 ( R_23d68_962ca20, \29378 );
buf \U$labaj5388 ( R_23d6a_9635f18, \29394 );
buf \U$labaj5389 ( R_23d6c_962ff48, \29410 );
buf \U$labaj5390 ( R_23d6e_9636068, \29426 );
buf \U$labaj5391 ( R_23d70_96363b0, \29444 );
buf \U$labaj5392 ( R_23d72_9636ae8, \29462 );
buf \U$labaj5393 ( R_23d74_9637220, \29480 );
buf \U$labaj5394 ( R_23d76_9637e98, \29498 );
buf \U$labaj5395 ( R_23d78_9638b10, \29516 );
buf \U$labaj5396 ( R_23d7a_962d4a0, \29534 );
buf \U$labaj5397 ( R_23d7e_96305d8, \29552 );
buf \U$labaj5398 ( R_23d80_9638bb8, \29570 );
buf \U$labaj5399 ( R_23d82_9638fa8, \29589 );
buf \U$labaj5400 ( R_23d84_962d548, \29607 );
buf \U$labaj5401 ( R_23d86_9639398, \29625 );
buf \U$labaj5402 ( R_23d88_95556e0, \29643 );
buf \U$labaj5403 ( R_23d8a_9639440, \29661 );
buf \U$labaj5404 ( R_23d8c_9d18d00, \29679 );
buf \U$labaj5405 ( R_23d8e_9d19d68, \29697 );
buf \U$labaj5406 ( R_23d90_9630a70, \29715 );
buf \U$labaj5407 ( R_23d94_9d1a008, \29733 );
buf \U$labaj5408 ( R_23d96_9d1a350, \29751 );
buf \U$labaj5409 ( R_23d98_9d1a9e0, \29769 );
buf \U$labaj5410 ( R_23d9a_96314f0, \29787 );
buf \U$labaj5411 ( R_23da4_9634430, \29818 );
buf \U$labaj5412 ( R_23dba_95558d8, \29838 );
buf \U$labaj5413 ( R_23dd0_9555a28, \29856 );
buf \U$labaj5414 ( R_23de6_9d1ac80, \29874 );
buf \U$labaj5415 ( R_23dfc_962d9e0, \29892 );
buf \U$labaj5416 ( R_23e12_9555b78, \29911 );
buf \U$labaj5417 ( R_23e1c_96344d8, \29929 );
buf \U$labaj5418 ( R_23e1e_9555e18, \29946 );
buf \U$labaj5419 ( R_23e20_9d1b070, \29963 );
buf \U$labaj5420 ( R_23e22_9d1b8f8, \29982 );
buf \U$labaj5421 ( R_23da6_9634a18, \29999 );
buf \U$labaj5422 ( R_23da8_9555f68, \30016 );
buf \U$labaj5423 ( R_23daa_9635150, \30032 );
buf \U$labaj5424 ( R_23dac_96352a0, \30048 );
buf \U$labaj5425 ( R_23dae_9556010, \30064 );
buf \U$labaj5426 ( R_23db0_9557078, \30080 );
buf \U$labaj5427 ( R_23db2_96353f0, \30096 );
buf \U$labaj5428 ( R_23db4_9d1ba48, \30112 );
buf \U$labaj5429 ( R_23db6_962db30, \30129 );
buf \U$labaj5430 ( R_23db8_96357e0, \30145 );
buf \U$labaj5431 ( R_23dbc_9559730, \30162 );
buf \U$labaj5432 ( R_23dbe_955bde8, \30179 );
buf \U$labaj5433 ( R_23dc0_955dd68, \30196 );
buf \U$labaj5434 ( R_23dc2_9d1baf0, \30213 );
buf \U$labaj5435 ( R_23dc4_955e158, \30230 );
buf \U$labaj5436 ( R_23dc6_9638db0, \30247 );
buf \U$labaj5437 ( R_23dc8_9d1bb98, \30264 );
buf \U$labaj5438 ( R_23dca_9639248, \30281 );
buf \U$labaj5439 ( R_23dcc_9d1bce8, \30298 );
buf \U$labaj5440 ( R_23dce_96c81c0, \30315 );
buf \U$labaj5441 ( R_23dd2_955e4a0, \30332 );
buf \U$labaj5442 ( R_23dd4_955ea88, \30349 );
buf \U$labaj5443 ( R_23dd6_96392f0, \30366 );
buf \U$labaj5444 ( R_23dd8_9d15d18, \30383 );
buf \U$labaj5445 ( R_23dda_955ee78, \30400 );
buf \U$labaj5446 ( R_23ddc_9d168e8, \30416 );
buf \U$labaj5447 ( R_23dde_9d16ae0, \30432 );
buf \U$labaj5448 ( R_23de0_962e310, \30448 );
buf \U$labaj5449 ( R_23de2_9d16c30, \30464 );
buf \U$labaj5450 ( R_23de4_9d16e28, \30480 );
buf \U$labaj5451 ( R_23de8_9d170c8, \30496 );
buf \U$labaj5452 ( R_23dea_955f1c0, \30512 );
buf \U$labaj5453 ( R_23dec_96c87a8, \30530 );
buf \U$labaj5454 ( R_23dee_955f310, \30548 );
buf \U$labaj5455 ( R_23df0_9d1bee0, \30565 );
buf \U$labaj5456 ( R_23df2_955f3b8, \30583 );
buf \U$labaj5457 ( R_23df4_95a39b0, \30600 );
buf \U$labaj5458 ( R_23df6_96c8af0, \30618 );
buf \U$labaj5459 ( R_23df8_95a3b00, \30635 );
buf \U$labaj5460 ( R_23dfa_95a40e8, \30652 );
buf \U$labaj5461 ( R_23dfe_95a44d8, \30669 );
buf \U$labaj5462 ( R_23e00_9d1bf88, \30686 );
buf \U$labaj5463 ( R_23e02_95a4580, \30703 );
buf \U$labaj5464 ( R_23e04_95a4c10, \30720 );
buf \U$labaj5465 ( R_23e06_9d17218, \30737 );
buf \U$labaj5466 ( R_23e08_95a5348, \30754 );
buf \U$labaj5467 ( R_23e0a_962ec40, \30771 );
buf \U$labaj5468 ( R_23e0c_9d17608, \30788 );
buf \U$labaj5469 ( R_23e0e_95a57e0, \30806 );
buf \U$labaj5470 ( R_23e10_95a5930, \30823 );
buf \U$labaj5471 ( R_23e14_9d18910, \30840 );
buf \U$labaj5472 ( R_23e16_9d19630, \30857 );
buf \U$labaj5473 ( R_23e18_95a5c78, \30874 );
buf \U$labaj5474 ( R_23e1a_95a6260, \30891 );
buf \U$labaj5475 ( R_23e24_9d1c030, \30917 );
buf \U$labaj5476 ( R_23e3a_95a4628, \30933 );
buf \U$labaj5477 ( R_23e50_95a48c8, \30949 );
buf \U$labaj5478 ( R_23e66_95a4b68, \30966 );
buf \U$labaj5479 ( R_23e7c_95b1438, \30981 );
buf \U$labaj5480 ( R_23e92_9d19780, \30996 );
buf \U$labaj5481 ( R_23e9c_95a6d88, \31010 );
buf \U$labaj5482 ( R_23e9e_95b1780, \31024 );
buf \U$labaj5483 ( R_23ea0_95a7028, \31038 );
buf \U$labaj5484 ( R_23ea2_95a70d0, \31053 );
buf \U$labaj5485 ( R_23e26_95b1828, \31067 );
buf \U$labaj5486 ( R_23e28_95a7220, \31081 );
buf \U$labaj5487 ( R_23e2a_95b2bd8, \31095 );
buf \U$labaj5488 ( R_23e2c_95b3310, \31109 );
buf \U$labaj5489 ( R_23e2e_95818b0, \31123 );
buf \U$labaj5490 ( R_23e30_9582138, \31137 );
buf \U$labaj5491 ( R_23e32_9582288, \31151 );
buf \U$labaj5492 ( R_23e34_95a7760, \31165 );
buf \U$labaj5493 ( R_23e36_9582870, \31179 );
buf \U$labaj5494 ( R_23e38_95a78b0, \31194 );
buf \U$labaj5495 ( R_23e3c_9d1c0d8, \31208 );
buf \U$labaj5496 ( R_23e3e_9582a68, \31222 );
buf \U$labaj5497 ( R_23e40_9d1b118, \31236 );
buf \U$labaj5498 ( R_23e42_9582e58, \31250 );
buf \U$labaj5499 ( R_23e44_9582f00, \31264 );
buf \U$labaj5500 ( R_23e46_95830f8, \31278 );
buf \U$labaj5501 ( R_23e48_958cbd8, \31292 );
buf \U$labaj5502 ( R_23e4a_958cc80, \31306 );
buf \U$labaj5503 ( R_23e4c_95a7aa8, \31320 );
buf \U$labaj5504 ( R_23e4e_958f5d8, \31334 );
buf \U$labaj5505 ( R_23e52_958f920, \31349 );
buf \U$labaj5506 ( R_23e54_9590058, \31363 );
buf \U$labaj5507 ( R_23e56_95a7bf8, \31377 );
buf \U$labaj5508 ( R_23e58_95a7ca0, \31391 );
buf \U$labaj5509 ( R_23e5a_95901a8, \31405 );
buf \U$labaj5510 ( R_23e5c_959fdb8, \31419 );
buf \U$labaj5511 ( R_23e5e_95a0b80, \31433 );
buf \U$labaj5512 ( R_23e60_9d1c4c8, \31447 );
buf \U$labaj5513 ( R_23e62_9625b28, \31461 );
buf \U$labaj5514 ( R_23e64_96261b8, \31475 );
buf \U$labaj5515 ( R_23e68_9d1b268, \31489 );
buf \U$labaj5516 ( R_23e6a_9d1c570, \31503 );
buf \U$labaj5517 ( R_23e6c_95a7d48, \31517 );
buf \U$labaj5518 ( R_23e6e_9626458, \31531 );
buf \U$labaj5519 ( R_23e70_95a8090, \31545 );
buf \U$labaj5520 ( R_23e72_9628330, \31559 );
buf \U$labaj5521 ( R_23e74_9628480, \31573 );
buf \U$labaj5522 ( R_23e76_9628528, \31587 );
buf \U$labaj5523 ( R_23e78_95a8138, \31601 );
buf \U$labaj5524 ( R_23e7a_96285d0, \31615 );
buf \U$labaj5525 ( R_23e7e_9628720, \31629 );
buf \U$labaj5526 ( R_23e80_9628bb8, \31643 );
buf \U$labaj5527 ( R_23e82_962c198, \31657 );
buf \U$labaj5528 ( R_23e84_9d1c618, \31671 );
buf \U$labaj5529 ( R_23e86_95a8288, \31685 );
buf \U$labaj5530 ( R_23e88_9634238, \31699 );
buf \U$labaj5531 ( R_23e8a_9d1c6c0, \31713 );
buf \U$labaj5532 ( R_23e8c_96342e0, \31727 );
buf \U$labaj5533 ( R_23e8e_9634970, \31741 );
buf \U$labaj5534 ( R_23e90_9d1c8b8, \31755 );
buf \U$labaj5535 ( R_23e94_9639830, \31769 );
buf \U$labaj5536 ( R_23e96_9d159d0, \31783 );
buf \U$labaj5537 ( R_23e98_9d15e68, \31797 );
buf \U$labaj5538 ( R_23e9a_95a83d8, \31811 );
buf \U$labaj5539 ( R_23c64_96c9a08, \31830 );
buf \U$labaj5540 ( R_23c66_9d1b658, \31847 );
buf \U$labaj5541 ( R_23c68_96ca920, \31863 );
buf \U$labaj5542 ( R_23c6a_9d244c0, \31879 );
buf \U$labaj5543 ( R_23c6c_96cb4f0, \31895 );
buf \U$labaj5544 ( R_23c6e_9d1b700, \31911 );
buf \U$labaj5545 ( R_23c70_9d1ca08, \31927 );
buf \U$labaj5546 ( R_23c72_96cb640, \31943 );
buf \U$labaj5547 ( R_23c74_962f030, \31958 );
buf \U$labaj5548 ( R_23c76_9d1cc00, \31973 );
buf \U$labaj5549 ( R_23c78_9d1cd50, \31988 );
buf \U$labaj5550 ( R_23c7a_9d1cdf8, \32003 );
buf \U$labaj5551 ( R_23c7c_9d1b7a8, \32018 );
buf \U$labaj5552 ( R_23c7e_9d1cf48, \32033 );
buf \U$labaj5553 ( R_23c80_9d1d098, \32048 );
buf \U$labaj5554 ( R_23c82_9d1d1e8, \32063 );
buf \U$labaj5555 ( R_23c84_95a8528, \32078 );
buf \U$labaj5556 ( R_23c86_9d1b9a0, \32093 );
buf \U$labaj5557 ( R_23c88_95a8720, \32108 );
buf \U$labaj5558 ( R_23c8a_9d1be38, \32123 );
buf \U$labaj5559 ( R_23c8c_9d246b8, \32138 );
buf \U$labaj5560 ( R_23c8e_96cb838, \32153 );
buf \U$labaj5561 ( R_23c90_9d24760, \32168 );
buf \U$labaj5562 ( R_23c92_9d1c2d0, \32183 );
buf \U$labaj5563 ( R_23c94_9d1d3e0, \32198 );
buf \U$labaj5564 ( R_23c96_95a87c8, \32213 );
buf \U$labaj5565 ( R_23c98_9d19438, \32228 );
buf \U$labaj5566 ( R_23c9a_9d1c378, \32243 );
buf \U$labaj5567 ( R_23c9c_9d1c768, \32258 );
buf \U$labaj5568 ( R_23c9e_9d1d488, \32273 );
buf \U$labaj5569 ( R_23ca0_9d1c960, \32288 );
buf \U$labaj5570 ( R_23ca2_9d1e8e0, \32303 );
buf \U$labaj5571 ( R_23ebc_9667ae0, \32315 );
buf \U$labaj5572 ( R_23ebe_965f6f8, \32326 );
buf \U$labaj5573 ( R_23ec0_9667b88, \32336 );
buf \U$labaj5574 ( R_23ec2_96688a8, \32346 );
buf \U$labaj5575 ( R_23ec4_95ac230, \32356 );
buf \U$labaj5576 ( R_23ec6_95ac428, \32366 );
buf \U$labaj5577 ( R_23ec8_966a780, \32376 );
buf \U$labaj5578 ( R_23eca_966a8d0, \32386 );
buf \U$labaj5579 ( R_23eba_965f8f0, \32396 );
buf \U$labaj5580 ( R_23ecc_95ac620, \32406 );
buf \U$labaj5581 ( R_23ece_95ac770, \32416 );
buf \U$labaj5582 ( R_23ed0_966a978, \32426 );
buf \U$labaj5583 ( R_23ed2_966aa20, \32436 );
buf \U$labaj5584 ( R_23eb8_966aac8, \32630 );
buf \U$labaj5585 ( R_23eea_95b1588, \32635 );
buf \U$labaj5586 ( R_23eec_9d1e448, \32640 );
buf \U$labaj5587 ( R_23eee_9d1e790, \32648 );
buf \U$labaj5588 ( R_23a0c_95b1630, \32705 );
buf \U$labaj5589 ( R_23a22_95b1c18, \32734 );
buf \U$labaj5590 ( R_23a38_966acc0, \32754 );
buf \U$labaj5591 ( R_23a4e_95b1d68, \32775 );
buf \U$labaj5592 ( R_23a64_966ad68, \32797 );
buf \U$labaj5593 ( R_23a7a_95b2c80, \32822 );
buf \U$labaj5594 ( R_23a84_9661a68, \32840 );
buf \U$labaj5595 ( R_23a86_9d1d7d0, \32863 );
buf \U$labaj5596 ( R_23a88_966ae10, \32885 );
buf \U$labaj5597 ( R_23a8a_966b0b0, \32906 );
buf \U$labaj5598 ( R_23a0e_962f420, \32925 );
buf \U$labaj5599 ( R_23a10_966ba88, \32945 );
buf \U$labaj5600 ( R_23a12_95b2fc8, \32964 );
buf \U$labaj5601 ( R_23a14_9d1f6a8, \32985 );
buf \U$labaj5602 ( R_23a16_952daf8, \33005 );
buf \U$labaj5603 ( R_23a18_95b3268, \33025 );
buf \U$labaj5604 ( R_23a1a_9581220, \33044 );
buf \U$labaj5605 ( R_23a1c_9d1d878, \33064 );
buf \U$labaj5606 ( R_23a1e_9663160, \33082 );
buf \U$labaj5607 ( R_23a20_9d1e250, \33102 );
buf \U$labaj5608 ( R_23a24_9d1fb40, \33121 );
buf \U$labaj5609 ( R_23a26_95305a0, \33140 );
buf \U$labaj5610 ( R_23a28_95812c8, \33160 );
buf \U$labaj5611 ( R_23a2a_9530798, \33178 );
buf \U$labaj5612 ( R_23a2c_95816b8, \33198 );
buf \U$labaj5613 ( R_23a2e_9663550, \33216 );
buf \U$labaj5614 ( R_23a30_9531e90, \33237 );
buf \U$labaj5615 ( R_23a32_9531f38, \33256 );
buf \U$labaj5616 ( R_23a34_9532130, \33276 );
buf \U$labaj5617 ( R_23a36_9532280, \33295 );
buf \U$labaj5618 ( R_23a3a_9532328, \33316 );
buf \U$labaj5619 ( R_23a3c_9581760, \33335 );
buf \U$labaj5620 ( R_23a3e_9581f40, \33355 );
buf \U$labaj5621 ( R_23a40_95323d0, \33374 );
buf \U$labaj5622 ( R_23a42_9532868, \33393 );
buf \U$labaj5623 ( R_23a44_9582720, \33413 );
buf \U$labaj5624 ( R_23a46_9532b08, \33433 );
buf \U$labaj5625 ( R_23a48_9532c58, \33451 );
buf \U$labaj5626 ( R_23a4a_9582918, \33470 );
buf \U$labaj5627 ( R_23a4c_966a4e0, \33489 );
buf \U$labaj5628 ( R_23a50_9532e50, \33508 );
buf \U$labaj5629 ( R_23a52_9d24808, \33528 );
buf \U$labaj5630 ( R_23a54_9533390, \33548 );
buf \U$labaj5631 ( R_23a56_9d20668, \33567 );
buf \U$labaj5632 ( R_23a58_9582db0, \33587 );
buf \U$labaj5633 ( R_23a5a_9583050, \33605 );
buf \U$labaj5634 ( R_23a5c_9533978, \33623 );
buf \U$labaj5635 ( R_23a5e_9534158, \33643 );
buf \U$labaj5636 ( R_23a60_9d20710, \33662 );
buf \U$labaj5637 ( R_23a62_95349e0, \33682 );
buf \U$labaj5638 ( R_23a66_9537290, \33702 );
buf \U$labaj5639 ( R_23a68_9d1f750, \33720 );
buf \U$labaj5640 ( R_23a6a_966a6d8, \33739 );
buf \U$labaj5641 ( R_23a6c_966aeb8, \33757 );
buf \U$labaj5642 ( R_23a6e_966b158, \33777 );
buf \U$labaj5643 ( R_23a70_9537a70, \33797 );
buf \U$labaj5644 ( R_23a72_9539f30, \33816 );
buf \U$labaj5645 ( R_23a74_95831a0, \33835 );
buf \U$labaj5646 ( R_23a76_9537c68, \33854 );
buf \U$labaj5647 ( R_23a78_9d20a58, \33873 );
buf \U$labaj5648 ( R_23a7c_9537d10, \33893 );
buf \U$labaj5649 ( R_23a7e_9537e60, \33913 );
buf \U$labaj5650 ( R_23a80_9538250, \33932 );
buf \U$labaj5651 ( R_23a82_95382f8, \33951 );
buf \U$labaj5652 ( R_23a8c_9d21e08, \33985 );
buf \U$labaj5653 ( R_23aa2_9583440, \34005 );
buf \U$labaj5654 ( R_23ab8_9d1f8a0, \34023 );
buf \U$labaj5655 ( R_23ace_9d1ff30, \34043 );
buf \U$labaj5656 ( R_23ae4_9d23ce0, \34062 );
buf \U$labaj5657 ( R_23afa_95834e8, \34081 );
buf \U$labaj5658 ( R_23b04_9583590, \34100 );
buf \U$labaj5659 ( R_23b06_9d20860, \34118 );
buf \U$labaj5660 ( R_23b08_9d24958, \34136 );
buf \U$labaj5661 ( R_23b0a_9d24ca0, \34154 );
buf \U$labaj5662 ( R_23a8e_95836e0, \34172 );
buf \U$labaj5663 ( R_23a90_9583e18, \34190 );
buf \U$labaj5664 ( R_23a92_9d25288, \34208 );
buf \U$labaj5665 ( R_23a94_9d20908, \34226 );
buf \U$labaj5666 ( R_23a96_9d25330, \34244 );
buf \U$labaj5667 ( R_23a98_9d22348, \34262 );
buf \U$labaj5668 ( R_23a9a_9d253d8, \34280 );
buf \U$labaj5669 ( R_23a9c_9d233b0, \34298 );
buf \U$labaj5670 ( R_23a9e_9d25528, \34317 );
buf \U$labaj5671 ( R_23aa0_9d255d0, \34336 );
buf \U$labaj5672 ( R_23aa4_9d23500, \34354 );
buf \U$labaj5673 ( R_23aa6_9d25678, \34372 );
buf \U$labaj5674 ( R_23aa8_9d23a40, \34390 );
buf \U$labaj5675 ( R_23aaa_9d24610, \34408 );
buf \U$labaj5676 ( R_23aac_9d25880, \34426 );
buf \U$labaj5677 ( R_23aae_9d248b0, \34444 );
buf \U$labaj5678 ( R_23ab0_9d26258, \34462 );
buf \U$labaj5679 ( R_23ab2_9584898, \34480 );
buf \U$labaj5680 ( R_23ab4_9d24a00, \34498 );
buf \U$labaj5681 ( R_23ab6_9d26450, \34516 );
buf \U$labaj5682 ( R_23aba_9d26648, \34534 );
buf \U$labaj5683 ( R_23abc_9d26e28, \34552 );
buf \U$labaj5684 ( R_23abe_9d270c8, \34570 );
buf \U$labaj5685 ( R_23ac0_9584c88, \34588 );
buf \U$labaj5686 ( R_23ac2_9d24aa8, \34606 );
buf \U$labaj5687 ( R_23ac4_9d24d48, \34624 );
buf \U$labaj5688 ( R_23ac6_9585270, \34642 );
buf \U$labaj5689 ( R_23ac8_9585708, \34660 );
buf \U$labaj5690 ( R_23aca_9d27bf0, \34679 );
buf \U$labaj5691 ( R_23acc_9d28910, \34697 );
buf \U$labaj5692 ( R_23ad0_9d29198, \34716 );
buf \U$labaj5693 ( R_23ad2_9d29630, \34734 );
buf \U$labaj5694 ( R_23ad4_9d24fe8, \34752 );
buf \U$labaj5695 ( R_23ad6_95857b0, \34770 );
buf \U$labaj5696 ( R_23ad8_9d2a0b0, \34788 );
buf \U$labaj5697 ( R_23ada_9585900, \34806 );
buf \U$labaj5698 ( R_23adc_9d2a200, \34824 );
buf \U$labaj5699 ( R_23ade_9d2a3f8, \34842 );
buf \U$labaj5700 ( R_23ae0_9d2a7e8, \34860 );
buf \U$labaj5701 ( R_23ae2_9d25138, \34878 );
buf \U$labaj5702 ( R_23ae6_9d2ad28, \34896 );
buf \U$labaj5703 ( R_23ae8_95860e0, \34914 );
buf \U$labaj5704 ( R_23aea_9d25480, \34934 );
buf \U$labaj5705 ( R_23aec_9d25928, \34952 );
buf \U$labaj5706 ( R_23aee_9d25bc8, \34970 );
buf \U$labaj5707 ( R_23af0_95864d0, \34988 );
buf \U$labaj5708 ( R_23af2_9d25e68, \35006 );
buf \U$labaj5709 ( R_23af4_95866c8, \35024 );
buf \U$labaj5710 ( R_23af6_9586770, \35042 );
buf \U$labaj5711 ( R_23af8_9587688, \35060 );
buf \U$labaj5712 ( R_23afc_9d26ed0, \35078 );
buf \U$labaj5713 ( R_23afe_9587730, \35096 );
buf \U$labaj5714 ( R_23b00_9d27aa0, \35114 );
buf \U$labaj5715 ( R_23b02_9d2add0, \35132 );
buf \U$labaj5716 ( R_23b0c_95877d8, \35165 );
buf \U$labaj5717 ( R_23b22_95386e8, \35183 );
buf \U$labaj5718 ( R_23b38_95388e0, \35201 );
buf \U$labaj5719 ( R_23b4e_9588108, \35219 );
buf \U$labaj5720 ( R_23b64_9538ad8, \35237 );
buf \U$labaj5721 ( R_23b7a_9d2b118, \35257 );
buf \U$labaj5722 ( R_23b84_95881b0, \35273 );
buf \U$labaj5723 ( R_23b86_95899f8, \35290 );
buf \U$labaj5724 ( R_23b88_9589aa0, \35307 );
buf \U$labaj5725 ( R_23b8a_9d2b460, \35326 );
buf \U$labaj5726 ( R_23b0e_958d268, \35343 );
buf \U$labaj5727 ( R_23b10_95390c0, \35360 );
buf \U$labaj5728 ( R_23b12_9539168, \35378 );
buf \U$labaj5729 ( R_23b14_95394b0, \35395 );
buf \U$labaj5730 ( R_23b16_95399f0, \35412 );
buf \U$labaj5731 ( R_23b18_9539c90, \35429 );
buf \U$labaj5732 ( R_23b1a_953ba18, \35446 );
buf \U$labaj5733 ( R_23b1c_953bac0, \35463 );
buf \U$labaj5734 ( R_23b1e_958d460, \35480 );
buf \U$labaj5735 ( R_23b20_9d2b508, \35497 );
buf \U$labaj5736 ( R_23b24_953bf58, \35514 );
buf \U$labaj5737 ( R_23b26_953c0a8, \35531 );
buf \U$labaj5738 ( R_23b28_953c1f8, \35549 );
buf \U$labaj5739 ( R_23b2a_953c540, \35566 );
buf \U$labaj5740 ( R_23b2c_9d2b5b0, \35583 );
buf \U$labaj5741 ( R_23b2e_953c888, \35600 );
buf \U$labaj5742 ( R_23b30_953cdc8, \35617 );
buf \U$labaj5743 ( R_23b32_958da48, \35634 );
buf \U$labaj5744 ( R_23b34_9d2b700, \35651 );
buf \U$labaj5745 ( R_23b36_953cf18, \35668 );
buf \U$labaj5746 ( R_23b3a_958de38, \35685 );
buf \U$labaj5747 ( R_23b3c_958e180, \35702 );
buf \U$labaj5748 ( R_23b3e_96ddca8, \35719 );
buf \U$labaj5749 ( R_23b40_96dddf8, \35736 );
buf \U$labaj5750 ( R_23b42_958e570, \35753 );
buf \U$labaj5751 ( R_23b44_958e810, \35770 );
buf \U$labaj5752 ( R_23b46_96de098, \35787 );
buf \U$labaj5753 ( R_23b48_9d285c8, \35804 );
buf \U$labaj5754 ( R_23b4a_96de3e0, \35821 );
buf \U$labaj5755 ( R_23b4c_9d28b08, \35838 );
buf \U$labaj5756 ( R_23b50_96de530, \35855 );
buf \U$labaj5757 ( R_23b52_958ef48, \35872 );
buf \U$labaj5758 ( R_23b54_9d24b50, \35889 );
buf \U$labaj5759 ( R_23b56_9d25d18, \35906 );
buf \U$labaj5760 ( R_23b58_958ff08, \35923 );
buf \U$labaj5761 ( R_23b5a_96e6c60, \35940 );
buf \U$labaj5762 ( R_23b5c_96e8160, \35957 );
buf \U$labaj5763 ( R_23b5e_96ebc70, \35974 );
buf \U$labaj5764 ( R_23b60_95903a0, \35991 );
buf \U$labaj5765 ( R_23b62_95906e8, \36008 );
buf \U$labaj5766 ( R_23b66_96ebdc0, \36025 );
buf \U$labaj5767 ( R_23b68_95efb90, \36042 );
buf \U$labaj5768 ( R_23b6a_9596d58, \36059 );
buf \U$labaj5769 ( R_23b6c_9d2b7a8, \36076 );
buf \U$labaj5770 ( R_23b6e_9598c30, \36093 );
buf \U$labaj5771 ( R_23b70_95f0220, \36110 );
buf \U$labaj5772 ( R_23b72_9598cd8, \36127 );
buf \U$labaj5773 ( R_23b74_95f1918, \36144 );
buf \U$labaj5774 ( R_23b76_9599170, \36162 );
buf \U$labaj5775 ( R_23b78_9d28bb0, \36179 );
buf \U$labaj5776 ( R_23b7c_95f37f0, \36196 );
buf \U$labaj5777 ( R_23b7e_95f41c8, \36213 );
buf \U$labaj5778 ( R_23b80_95f4318, \36230 );
buf \U$labaj5779 ( R_23b82_95992c0, \36247 );
buf \U$labaj5780 ( R_23b8c_9599608, \36274 );
buf \U$labaj5781 ( R_23ba2_9599758, \36290 );
buf \U$labaj5782 ( R_23bb8_9599800, \36306 );
buf \U$labaj5783 ( R_23bce_9599950, \36321 );
buf \U$labaj5784 ( R_23be4_962f570, \36336 );
buf \U$labaj5785 ( R_23bfa_9599b48, \36351 );
buf \U$labaj5786 ( R_23c04_959a088, \36365 );
buf \U$labaj5787 ( R_23c06_959a130, \36380 );
buf \U$labaj5788 ( R_23c08_959a1d8, \36394 );
buf \U$labaj5789 ( R_23c0a_962f618, \36409 );
buf \U$labaj5790 ( R_23b8e_959a5c8, \36423 );
buf \U$labaj5791 ( R_23b90_959a9b8, \36437 );
buf \U$labaj5792 ( R_23b92_959ac58, \36451 );
buf \U$labaj5793 ( R_23b94_959aef8, \36465 );
buf \U$labaj5794 ( R_23b96_962f8b8, \36479 );
buf \U$labaj5795 ( R_23b98_959afa0, \36493 );
buf \U$labaj5796 ( R_23b9a_959b048, \36507 );
buf \U$labaj5797 ( R_23b9c_959b0f0, \36521 );
buf \U$labaj5798 ( R_23b9e_959b198, \36535 );
buf \U$labaj5799 ( R_23ba0_959b240, \36550 );
buf \U$labaj5800 ( R_23ba4_959b6d8, \36564 );
buf \U$labaj5801 ( R_23ba6_959b828, \36578 );
buf \U$labaj5802 ( R_23ba8_959b8d0, \36592 );
buf \U$labaj5803 ( R_23baa_959ba20, \36606 );
buf \U$labaj5804 ( R_23bac_9d28da8, \36620 );
buf \U$labaj5805 ( R_23bae_959bac8, \36634 );
buf \U$labaj5806 ( R_23bb0_959d268, \36648 );
buf \U$labaj5807 ( R_23bb2_959d508, \36662 );
buf \U$labaj5808 ( R_23bb4_959dce8, \36676 );
buf \U$labaj5809 ( R_23bb6_959e420, \36690 );
buf \U$labaj5810 ( R_23bba_9d28fa0, \36705 );
buf \U$labaj5811 ( R_23bbc_962f960, \36719 );
buf \U$labaj5812 ( R_23bbe_9d298d0, \36733 );
buf \U$labaj5813 ( R_23bc0_959e618, \36747 );
buf \U$labaj5814 ( R_23bc2_959eea0, \36761 );
buf \U$labaj5815 ( R_23bc4_959f098, \36775 );
buf \U$labaj5816 ( R_23bc6_9d29978, \36789 );
buf \U$labaj5817 ( R_23bc8_9d25dc0, \36803 );
buf \U$labaj5818 ( R_23bca_959f9c8, \36817 );
buf \U$labaj5819 ( R_23bcc_9d29a20, \36831 );
buf \U$labaj5820 ( R_23bd0_95a0e20, \36845 );
buf \U$labaj5821 ( R_23bd2_9d29b70, \36859 );
buf \U$labaj5822 ( R_23bd4_962fb58, \36873 );
buf \U$labaj5823 ( R_23bd6_95a0f70, \36887 );
buf \U$labaj5824 ( R_23bd8_9d29c18, \36901 );
buf \U$labaj5825 ( R_23bda_9619ae0, \36915 );
buf \U$labaj5826 ( R_23bdc_9619b88, \36929 );
buf \U$labaj5827 ( R_23bde_9619d80, \36943 );
buf \U$labaj5828 ( R_23be0_9619e28, \36957 );
buf \U$labaj5829 ( R_23be2_961a020, \36971 );
buf \U$labaj5830 ( R_23be6_961a0c8, \36985 );
buf \U$labaj5831 ( R_23be8_961a218, \36999 );
buf \U$labaj5832 ( R_23bea_961a4b8, \37013 );
buf \U$labaj5833 ( R_23bec_961a800, \37027 );
buf \U$labaj5834 ( R_23bee_961a8a8, \37041 );
buf \U$labaj5835 ( R_23bf0_961a950, \37055 );
buf \U$labaj5836 ( R_23bf2_961ad40, \37069 );
buf \U$labaj5837 ( R_23bf4_961ade8, \37083 );
buf \U$labaj5838 ( R_23bf6_961ae90, \37097 );
buf \U$labaj5839 ( R_23bf8_961af38, \37111 );
buf \U$labaj5840 ( R_23bfc_9d26060, \37125 );
buf \U$labaj5841 ( R_23bfe_961b088, \37139 );
buf \U$labaj5842 ( R_23c00_9d29d68, \37153 );
buf \U$labaj5843 ( R_23c02_961b1d8, \37167 );
buf \U$labaj5844 ( R_239cc_95f4af8, \37186 );
buf \U$labaj5845 ( R_239ce_962fd50, \37204 );
buf \U$labaj5846 ( R_239d0_9558e00, \37220 );
buf \U$labaj5847 ( R_239d2_9d261b0, \37237 );
buf \U$labaj5848 ( R_239d4_95f52d8, \37254 );
buf \U$labaj5849 ( R_239d6_9558ea8, \37271 );
buf \U$labaj5850 ( R_239d8_961b670, \37288 );
buf \U$labaj5851 ( R_239da_95f5620, \37305 );
buf \U$labaj5852 ( R_239dc_961b910, \37320 );
buf \U$labaj5853 ( R_239de_9d2b850, \37335 );
buf \U$labaj5854 ( R_239e0_9d2b9a0, \37350 );
buf \U$labaj5855 ( R_239e2_9d29e10, \37365 );
buf \U$labaj5856 ( R_239e4_9d2a158, \37380 );
buf \U$labaj5857 ( R_239e6_961bb08, \37395 );
buf \U$labaj5858 ( R_239e8_961c978, \37410 );
buf \U$labaj5859 ( R_239ea_961cd68, \37425 );
buf \U$labaj5860 ( R_239ec_9d2baf0, \37440 );
buf \U$labaj5861 ( R_239ee_95f5968, \37455 );
buf \U$labaj5862 ( R_239f0_95f5ab8, \37470 );
buf \U$labaj5863 ( R_239f2_9d2a2a8, \37485 );
buf \U$labaj5864 ( R_239f4_961ce10, \37500 );
buf \U$labaj5865 ( R_239f6_9634e08, \37515 );
buf \U$labaj5866 ( R_239f8_9d2bb98, \37530 );
buf \U$labaj5867 ( R_239fa_9d2bd90, \37545 );
buf \U$labaj5868 ( R_239fc_962fdf8, \37560 );
buf \U$labaj5869 ( R_239fe_962fea0, \37575 );
buf \U$labaj5870 ( R_23a00_961d200, \37590 );
buf \U$labaj5871 ( R_23a02_961d5f0, \37605 );
buf \U$labaj5872 ( R_23a04_961d698, \37620 );
buf \U$labaj5873 ( R_23a06_962fff0, \37635 );
buf \U$labaj5874 ( R_23a08_961d740, \37650 );
buf \U$labaj5875 ( R_23a0a_961d938, \37665 );
buf \U$labaj5876 ( R_23c24_9d2a698, \37677 );
buf \U$labaj5877 ( R_23c26_9d2c420, \37688 );
buf \U$labaj5878 ( R_23c28_962ac98, \37698 );
buf \U$labaj5879 ( R_23c2a_9d2c4c8, \37708 );
buf \U$labaj5880 ( R_23c2c_9d2c570, \37718 );
buf \U$labaj5881 ( R_23c2e_95f63e8, \37728 );
buf \U$labaj5882 ( R_23c30_9d2a890, \37738 );
buf \U$labaj5883 ( R_23c32_962ad40, \37748 );
buf \U$labaj5884 ( R_23c22_9d2aa88, \37758 );
buf \U$labaj5885 ( R_23c34_9d2c810, \37768 );
buf \U$labaj5886 ( R_23c36_9d2ab30, \37778 );
buf \U$labaj5887 ( R_23c38_9d2c8b8, \37788 );
buf \U$labaj5888 ( R_23c3a_9d2cab0, \37798 );
buf \U$labaj5889 ( R_23c20_9635e70, \37998 );
buf \U$labaj5890 ( R_23c52_962b868, \38003 );
buf \U$labaj5891 ( R_23c54_9d2af20, \38008 );
buf \U$labaj5892 ( R_23c56_9d2b310, \38013 );
buf \U$labaj5893 ( R_23774_9630098, \38069 );
buf \U$labaj5894 ( R_2378a_962b9b8, \38097 );
buf \U$labaj5895 ( R_237a0_9d2cd50, \38116 );
buf \U$labaj5896 ( R_237b6_962bb08, \38137 );
buf \U$labaj5897 ( R_237cc_9d2cff0, \38156 );
buf \U$labaj5898 ( R_237e2_9d2d098, \38182 );
buf \U$labaj5899 ( R_237ec_9d2d140, \38202 );
buf \U$labaj5900 ( R_237ee_9d2d290, \38222 );
buf \U$labaj5901 ( R_237f0_962c240, \38242 );
buf \U$labaj5902 ( R_237f2_9559688, \38262 );
buf \U$labaj5903 ( R_23776_96301e8, \38282 );
buf \U$labaj5904 ( R_23778_9d2d7d0, \38301 );
buf \U$labaj5905 ( R_2377a_962c2e8, \38320 );
buf \U$labaj5906 ( R_2377c_9d2d878, \38340 );
buf \U$labaj5907 ( R_2377e_962ce10, \38360 );
buf \U$labaj5908 ( R_23780_9d2d920, \38379 );
buf \U$labaj5909 ( R_23782_962d938, \38398 );
buf \U$labaj5910 ( R_23784_962e5b0, \38418 );
buf \U$labaj5911 ( R_23786_9d2d9c8, \38436 );
buf \U$labaj5912 ( R_23788_9d2dc68, \38454 );
buf \U$labaj5913 ( R_2378c_9d2dd10, \38473 );
buf \U$labaj5914 ( R_2378e_9d2ddb8, \38492 );
buf \U$labaj5915 ( R_23790_9d2e100, \38511 );
buf \U$labaj5916 ( R_23792_9d2e1a8, \38529 );
buf \U$labaj5917 ( R_23794_9d2f0c0, \38548 );
buf \U$labaj5918 ( R_23796_9630290, \38566 );
buf \U$labaj5919 ( R_23798_96303e0, \38584 );
buf \U$labaj5920 ( R_2379a_9d2f210, \38602 );
buf \U$labaj5921 ( R_2379c_9d2f7f8, \38623 );
buf \U$labaj5922 ( R_2379e_9630728, \38644 );
buf \U$labaj5923 ( R_237a2_96307d0, \38664 );
buf \U$labaj5924 ( R_237a4_9d2fb40, \38684 );
buf \U$labaj5925 ( R_237a6_9d301d0, \38704 );
buf \U$labaj5926 ( R_237a8_9559bc8, \38724 );
buf \U$labaj5927 ( R_237aa_9630140, \38745 );
buf \U$labaj5928 ( R_237ac_96312f8, \38765 );
buf \U$labaj5929 ( R_237ae_9d30710, \38784 );
buf \U$labaj5930 ( R_237b0_9630b18, \38803 );
buf \U$labaj5931 ( R_237b2_9630c68, \38821 );
buf \U$labaj5932 ( R_237b4_9d309b0, \38840 );
buf \U$labaj5933 ( R_237b8_9630d10, \38858 );
buf \U$labaj5934 ( R_237ba_9630fb0, \38876 );
buf \U$labaj5935 ( R_237bc_9631100, \38894 );
buf \U$labaj5936 ( R_237be_9d30a58, \38913 );
buf \U$labaj5937 ( R_237c0_9d30da0, \38932 );
buf \U$labaj5938 ( R_237c2_96311a8, \38951 );
buf \U$labaj5939 ( R_237c4_96313a0, \38969 );
buf \U$labaj5940 ( R_237c6_96318e0, \38988 );
buf \U$labaj5941 ( R_237c8_9631a30, \39006 );
buf \U$labaj5942 ( R_237ca_9d30e48, \39025 );
buf \U$labaj5943 ( R_237ce_9d31190, \39044 );
buf \U$labaj5944 ( R_237d0_9631b80, \39065 );
buf \U$labaj5945 ( R_237d2_9d31f58, \39085 );
buf \U$labaj5946 ( R_237d4_9631448, \39104 );
buf \U$labaj5947 ( R_237d6_9631790, \39123 );
buf \U$labaj5948 ( R_237d8_9d323f0, \39142 );
buf \U$labaj5949 ( R_237da_9631ad8, \39162 );
buf \U$labaj5950 ( R_237dc_9d32540, \39182 );
buf \U$labaj5951 ( R_237de_9632018, \39201 );
buf \U$labaj5952 ( R_237e0_9631cd0, \39222 );
buf \U$labaj5953 ( R_237e4_9632210, \39241 );
buf \U$labaj5954 ( R_237e6_9d32690, \39261 );
buf \U$labaj5955 ( R_237e8_96322b8, \39280 );
buf \U$labaj5956 ( R_237ea_9d32888, \39299 );
buf \U$labaj5957 ( R_237f4_9631e20, \39331 );
buf \U$labaj5958 ( R_2380a_9d329d8, \39352 );
buf \U$labaj5959 ( R_23820_9d32a80, \39371 );
buf \U$labaj5960 ( R_23836_9d32f18, \39391 );
buf \U$labaj5961 ( R_2384c_9d2b3b8, \39410 );
buf \U$labaj5962 ( R_23862_9631ec8, \39429 );
buf \U$labaj5963 ( R_2386c_9632360, \39448 );
buf \U$labaj5964 ( R_2386e_9632a98, \39466 );
buf \U$labaj5965 ( R_23870_9d32fc0, \39484 );
buf \U$labaj5966 ( R_23872_9632408, \39502 );
buf \U$labaj5967 ( R_237f6_9632600, \39521 );
buf \U$labaj5968 ( R_237f8_9d33500, \39539 );
buf \U$labaj5969 ( R_237fa_96326a8, \39557 );
buf \U$labaj5970 ( R_237fc_9d33650, \39575 );
buf \U$labaj5971 ( R_237fe_9d336f8, \39593 );
buf \U$labaj5972 ( R_23800_9d33a40, \39611 );
buf \U$labaj5973 ( R_23802_9632750, \39629 );
buf \U$labaj5974 ( R_23804_96328a0, \39647 );
buf \U$labaj5975 ( R_23806_9d340d0, \39665 );
buf \U$labaj5976 ( R_23808_9632948, \39683 );
buf \U$labaj5977 ( R_2380c_9d2b658, \39701 );
buf \U$labaj5978 ( R_2380e_9d34418, \39719 );
buf \U$labaj5979 ( R_23810_9d34760, \39737 );
buf \U$labaj5980 ( R_23812_9d34fe8, \39755 );
buf \U$labaj5981 ( R_23814_9632de0, \39773 );
buf \U$labaj5982 ( R_23816_9632e88, \39791 );
buf \U$labaj5983 ( R_23818_9d35720, \39809 );
buf \U$labaj5984 ( R_2381a_9d2bc40, \39827 );
buf \U$labaj5985 ( R_2381c_b805670, \39845 );
buf \U$labaj5986 ( R_2381e_b805868, \39863 );
buf \U$labaj5987 ( R_23822_9633080, \39881 );
buf \U$labaj5988 ( R_23824_b8060f0, \39899 );
buf \U$labaj5989 ( R_23826_9633128, \39917 );
buf \U$labaj5990 ( R_23828_9633b00, \39935 );
buf \U$labaj5991 ( R_2382a_9632b40, \39953 );
buf \U$labaj5992 ( R_2382c_9634190, \39971 );
buf \U$labaj5993 ( R_2382e_9638720, \39989 );
buf \U$labaj5994 ( R_23830_9d2c180, \40007 );
buf \U$labaj5995 ( R_23832_96389c0, \40026 );
buf \U$labaj5996 ( R_23834_9638a68, \40044 );
buf \U$labaj5997 ( R_23838_9d15880, \40062 );
buf \U$labaj5998 ( R_2383a_b806198, \40080 );
buf \U$labaj5999 ( R_2383c_9d2c768, \40098 );
buf \U$labaj6000 ( R_2383e_9d16a38, \40116 );
buf \U$labaj6001 ( R_23840_9d2ca08, \40134 );
buf \U$labaj6002 ( R_23842_b806240, \40152 );
buf \U$labaj6003 ( R_23844_9d17170, \40170 );
buf \U$labaj6004 ( R_23846_9d17c98, \40188 );
buf \U$labaj6005 ( R_23848_b8062e8, \40206 );
buf \U$labaj6006 ( R_2384a_b806390, \40224 );
buf \U$labaj6007 ( R_2384e_9d2cca8, \40242 );
buf \U$labaj6008 ( R_23850_9d17fe0, \40260 );
buf \U$labaj6009 ( R_23852_9d18328, \40279 );
buf \U$labaj6010 ( R_23854_9d2d1e8, \40297 );
buf \U$labaj6011 ( R_23856_9d1fd38, \40315 );
buf \U$labaj6012 ( R_23858_b8064e0, \40333 );
buf \U$labaj6013 ( R_2385a_9d2d3e0, \40351 );
buf \U$labaj6014 ( R_2385c_9d220a8, \40369 );
buf \U$labaj6015 ( R_2385e_9535d90, \40387 );
buf \U$labaj6016 ( R_23860_b806588, \40405 );
buf \U$labaj6017 ( R_23864_9d25720, \40423 );
buf \U$labaj6018 ( R_23866_b8066d8, \40441 );
buf \U$labaj6019 ( R_23868_b806780, \40459 );
buf \U$labaj6020 ( R_2386a_9d2d530, \40477 );
buf \U$labaj6021 ( R_23874_95f7840, \40508 );
buf \U$labaj6022 ( R_2388a_95f7e28, \40528 );
buf \U$labaj6023 ( R_238a0_9d28e50, \40546 );
buf \U$labaj6024 ( R_238b6_95f8170, \40564 );
buf \U$labaj6025 ( R_238cc_95fcd90, \40582 );
buf \U$labaj6026 ( R_238e2_95fda08, \40600 );
buf \U$labaj6027 ( R_238ec_95fdb58, \40617 );
buf \U$labaj6028 ( R_238ee_95fdca8, \40634 );
buf \U$labaj6029 ( R_238f0_95fdd50, \40652 );
buf \U$labaj6030 ( R_238f2_9d2d728, \40670 );
buf \U$labaj6031 ( R_23876_95ff6e8, \40689 );
buf \U$labaj6032 ( R_23878_9535e38, \40707 );
buf \U$labaj6033 ( R_2387a_9633668, \40725 );
buf \U$labaj6034 ( R_2387c_9f4ddd0, \40742 );
buf \U$labaj6035 ( R_2387e_9f51b80, \40759 );
buf \U$labaj6036 ( R_23880_9f51e20, \40776 );
buf \U$labaj6037 ( R_23882_9d29ac8, \40793 );
buf \U$labaj6038 ( R_23884_9f53278, \40810 );
buf \U$labaj6039 ( R_23886_9f53320, \40827 );
buf \U$labaj6040 ( R_23888_9f54580, \40844 );
buf \U$labaj6041 ( R_2388c_9f54778, \40861 );
buf \U$labaj6042 ( R_2388e_9d2dbc0, \40878 );
buf \U$labaj6043 ( R_23890_9d2e250, \40896 );
buf \U$labaj6044 ( R_23892_9f548c8, \40913 );
buf \U$labaj6045 ( R_23894_9f54970, \40930 );
buf \U$labaj6046 ( R_23896_9f54c10, \40947 );
buf \U$labaj6047 ( R_23898_9f55348, \40964 );
buf \U$labaj6048 ( R_2389a_9f55498, \40981 );
buf \U$labaj6049 ( R_2389c_9d2a740, \40998 );
buf \U$labaj6050 ( R_2389e_9d2e3a0, \41015 );
buf \U$labaj6051 ( R_238a2_9d2b070, \41032 );
buf \U$labaj6052 ( R_238a4_9633710, \41049 );
buf \U$labaj6053 ( R_238a6_9f55b28, \41066 );
buf \U$labaj6054 ( R_238a8_9f56260, \41083 );
buf \U$labaj6055 ( R_238aa_9f56500, \41100 );
buf \U$labaj6056 ( R_238ac_9f5baf8, \41117 );
buf \U$labaj6057 ( R_238ae_9ee9d78, \41134 );
buf \U$labaj6058 ( R_238b0_9d2ba48, \41151 );
buf \U$labaj6059 ( R_238b2_9d2bce8, \41168 );
buf \U$labaj6060 ( R_238b4_9eea0c0, \41185 );
buf \U$labaj6061 ( R_238b8_9eeb518, \41202 );
buf \U$labaj6062 ( R_238ba_9eedf18, \41219 );
buf \U$labaj6063 ( R_238bc_9eee6f8, \41236 );
buf \U$labaj6064 ( R_238be_9ef2010, \41253 );
buf \U$labaj6065 ( R_238c0_9537530, \41270 );
buf \U$labaj6066 ( R_238c2_9ef2208, \41288 );
buf \U$labaj6067 ( R_238c4_9ef3660, \41305 );
buf \U$labaj6068 ( R_238c6_9ef3858, \41323 );
buf \U$labaj6069 ( R_238c8_9633860, \41340 );
buf \U$labaj6070 ( R_238ca_9ef3a50, \41357 );
buf \U$labaj6071 ( R_238ce_9ef3af8, \41374 );
buf \U$labaj6072 ( R_238d0_9ef3ba0, \41391 );
buf \U$labaj6073 ( R_238d2_9ef3c48, \41408 );
buf \U$labaj6074 ( R_238d4_9ef4620, \41425 );
buf \U$labaj6075 ( R_238d6_9d2c2d0, \41442 );
buf \U$labaj6076 ( R_238d8_9ef4770, \41459 );
buf \U$labaj6077 ( R_238da_9d2cb58, \41476 );
buf \U$labaj6078 ( R_238dc_9ef4ab8, \41493 );
buf \U$labaj6079 ( R_238de_9ef4c08, \41511 );
buf \U$labaj6080 ( R_238e0_9ef4ff8, \41528 );
buf \U$labaj6081 ( R_238e4_9ef5148, \41545 );
buf \U$labaj6082 ( R_238e6_9ef51f0, \41562 );
buf \U$labaj6083 ( R_238e8_9d2cf48, \41579 );
buf \U$labaj6084 ( R_238ea_9ef53e8, \41596 );
buf \U$labaj6085 ( R_238f4_9d2e4f0, \41621 );
buf \U$labaj6086 ( R_2390a_96339b0, \41637 );
buf \U$labaj6087 ( R_23920_9633c50, \41654 );
buf \U$labaj6088 ( R_23936_9d266f0, \41670 );
buf \U$labaj6089 ( R_2394c_9d2e838, \41684 );
buf \U$labaj6090 ( R_23962_9d2ecd0, \41699 );
buf \U$labaj6091 ( R_2396c_9d2ed78, \41713 );
buf \U$labaj6092 ( R_2396e_9d2f018, \41727 );
buf \U$labaj6093 ( R_23970_9d2f168, \41741 );
buf \U$labaj6094 ( R_23972_b8068d0, \41756 );
buf \U$labaj6095 ( R_238f6_9d2f2b8, \41770 );
buf \U$labaj6096 ( R_238f8_9d2f9f0, \41784 );
buf \U$labaj6097 ( R_238fa_9d2fde0, \41798 );
buf \U$labaj6098 ( R_238fc_9633f98, \41812 );
buf \U$labaj6099 ( R_238fe_b806a20, \41827 );
buf \U$labaj6100 ( R_23900_96340e8, \41841 );
buf \U$labaj6101 ( R_23902_9d30320, \41855 );
buf \U$labaj6102 ( R_23904_9634580, \41869 );
buf \U$labaj6103 ( R_23906_9d305c0, \41883 );
buf \U$labaj6104 ( R_23908_9634b68, \41897 );
buf \U$labaj6105 ( R_2390c_9d30ba8, \41911 );
buf \U$labaj6106 ( R_2390e_9d30c50, \41925 );
buf \U$labaj6107 ( R_23910_b806ac8, \41939 );
buf \U$labaj6108 ( R_23912_9d32000, \41953 );
buf \U$labaj6109 ( R_23914_b806b70, \41967 );
buf \U$labaj6110 ( R_23916_9d320a8, \41981 );
buf \U$labaj6111 ( R_23918_9634c10, \41995 );
buf \U$labaj6112 ( R_2391a_9d32150, \42009 );
buf \U$labaj6113 ( R_2391c_9634cb8, \42023 );
buf \U$labaj6114 ( R_2391e_9d32498, \42037 );
buf \U$labaj6115 ( R_23922_9d32738, \42052 );
buf \U$labaj6116 ( R_23924_9d327e0, \42066 );
buf \U$labaj6117 ( R_23926_9d32b28, \42080 );
buf \U$labaj6118 ( R_23928_9d32bd0, \42094 );
buf \U$labaj6119 ( R_2392a_9635348, \42108 );
buf \U$labaj6120 ( R_2392c_9635690, \42122 );
buf \U$labaj6121 ( R_2392e_9d32c78, \42136 );
buf \U$labaj6122 ( R_23930_9d32d20, \42150 );
buf \U$labaj6123 ( R_23932_9635a80, \42164 );
buf \U$labaj6124 ( R_23934_9d32dc8, \42178 );
buf \U$labaj6125 ( R_23938_9d331b8, \42192 );
buf \U$labaj6126 ( R_2393a_9d2d488, \42206 );
buf \U$labaj6127 ( R_2393c_9d333b0, \42220 );
buf \U$labaj6128 ( R_2393e_9d335a8, \42234 );
buf \U$labaj6129 ( R_23940_9d337a0, \42248 );
buf \U$labaj6130 ( R_23942_9635b28, \42262 );
buf \U$labaj6131 ( R_23944_9d2d5d8, \42276 );
buf \U$labaj6132 ( R_23946_9d338f0, \42290 );
buf \U$labaj6133 ( R_23948_9635bd0, \42304 );
buf \U$labaj6134 ( R_2394a_9d33998, \42318 );
buf \U$labaj6135 ( R_2394e_9d33ae8, \42332 );
buf \U$labaj6136 ( R_23950_9d33b90, \42346 );
buf \U$labaj6137 ( R_23952_9636110, \42360 );
buf \U$labaj6138 ( R_23954_9d33ce0, \42374 );
buf \U$labaj6139 ( R_23956_b806c18, \42388 );
buf \U$labaj6140 ( R_23958_9d33ed8, \42402 );
buf \U$labaj6141 ( R_2395a_9d33f80, \42416 );
buf \U$labaj6142 ( R_2395c_9636308, \42430 );
buf \U$labaj6143 ( R_2395e_b806cc0, \42444 );
buf \U$labaj6144 ( R_23960_9d34028, \42458 );
buf \U$labaj6145 ( R_23964_9d34178, \42472 );
buf \U$labaj6146 ( R_23966_9d2db18, \42486 );
buf \U$labaj6147 ( R_23968_96365a8, \42500 );
buf \U$labaj6148 ( R_2396a_9636848, \42514 );
buf \U$labaj6149 ( R_23734_96368f0, \42534 );
buf \U$labaj6150 ( R_23736_9636998, \42551 );
buf \U$labaj6151 ( R_23738_9636a40, \42568 );
buf \U$labaj6152 ( R_2373a_b7dc0c0, \42585 );
buf \U$labaj6153 ( R_2373c_9636b90, \42602 );
buf \U$labaj6154 ( R_2373e_9636c38, \42619 );
buf \U$labaj6155 ( R_23740_b7dc168, \42636 );
buf \U$labaj6156 ( R_23742_b806d68, \42653 );
buf \U$labaj6157 ( R_23744_b806e10, \42668 );
buf \U$labaj6158 ( R_23746_9636ed8, \42683 );
buf \U$labaj6159 ( R_23748_b806eb8, \42698 );
buf \U$labaj6160 ( R_2374a_9637028, \42713 );
buf \U$labaj6161 ( R_2374c_b806f60, \42728 );
buf \U$labaj6162 ( R_2374e_b8070b0, \42743 );
buf \U$labaj6163 ( R_23750_9d33308, \42758 );
buf \U$labaj6164 ( R_23752_b807158, \42773 );
buf \U$labaj6165 ( R_23754_9ef5880, \42788 );
buf \U$labaj6166 ( R_23756_9d26798, \42803 );
buf \U$labaj6167 ( R_23758_9d342c8, \42818 );
buf \U$labaj6168 ( R_2375a_9ef5928, \42833 );
buf \U$labaj6169 ( R_2375c_96c2b20, \42848 );
buf \U$labaj6170 ( R_2375e_9d31820, \42863 );
buf \U$labaj6171 ( R_23760_9d31970, \42878 );
buf \U$labaj6172 ( R_23762_9637178, \42893 );
buf \U$labaj6173 ( R_23764_9d26840, \42908 );
buf \U$labaj6174 ( R_23766_96372c8, \42923 );
buf \U$labaj6175 ( R_23768_9d268e8, \42938 );
buf \U$labaj6176 ( R_2376a_9d26a38, \42953 );
buf \U$labaj6177 ( R_2376c_9d26ae0, \42968 );
buf \U$labaj6178 ( R_2376e_9637370, \42983 );
buf \U$labaj6179 ( R_23770_9d26b88, \42998 );
buf \U$labaj6180 ( R_23772_9637418, \43013 );
buf \U$labaj6181 ( R_2398c_96c2fb8, \43028 );
buf \U$labaj6182 ( R_2398e_9559c70, \43039 );
buf \U$labaj6183 ( R_23990_96c35a0, \43049 );
buf \U$labaj6184 ( R_23992_96e8010, \43059 );
buf \U$labaj6185 ( R_23994_955a300, \43069 );
buf \U$labaj6186 ( R_23996_955a450, \43079 );
buf \U$labaj6187 ( R_23998_9d34ca0, \43089 );
buf \U$labaj6188 ( R_2399a_96c3840, \43099 );
buf \U$labaj6189 ( R_2398a_9d34d48, \43109 );
buf \U$labaj6190 ( R_2399c_96c3a38, \43119 );
buf \U$labaj6191 ( R_2399e_96c3d80, \43129 );
buf \U$labaj6192 ( R_239a0_955a840, \43139 );
buf \U$labaj6193 ( R_239a2_96c59b8, \43149 );
buf \U$labaj6194 ( R_23988_96eaf50, \43344 );
buf \U$labaj6195 ( R_239ba_96ca728, \43349 );
buf \U$labaj6196 ( R_239bc_955b8a8, \43354 );
buf \U$labaj6197 ( R_239be_b7db6e8, \43360 );
buf \U$labaj6198 ( R_234dc_b8085b0, \43420 );
buf \U$labaj6199 ( R_234f2_b80b988, \43442 );
buf \U$labaj6200 ( R_23508_b808658, \43461 );
buf \U$labaj6201 ( R_2351e_b808700, \43481 );
buf \U$labaj6202 ( R_23534_b8087a8, \43502 );
buf \U$labaj6203 ( R_2354a_b8088f8, \43525 );
buf \U$labaj6204 ( R_23554_b80ba30, \43546 );
buf \U$labaj6205 ( R_23556_b80bb80, \43567 );
buf \U$labaj6206 ( R_23558_b80bec8, \43588 );
buf \U$labaj6207 ( R_2355a_b80bf70, \43612 );
buf \U$labaj6208 ( R_234de_b8089a0, \43633 );
buf \U$labaj6209 ( R_234e0_b808a48, \43651 );
buf \U$labaj6210 ( R_234e2_b809768, \43672 );
buf \U$labaj6211 ( R_234e4_b809df8, \43691 );
buf \U$labaj6212 ( R_234e6_b80c2b8, \43709 );
buf \U$labaj6213 ( R_234e8_b80e040, \43729 );
buf \U$labaj6214 ( R_234ea_b80e580, \43749 );
buf \U$labaj6215 ( R_234ec_b80c600, \43767 );
buf \U$labaj6216 ( R_234ee_b80f0a8, \43787 );
buf \U$labaj6217 ( R_234f0_b80fd20, \43806 );
buf \U$labaj6218 ( R_234f4_b80c750, \43824 );
buf \U$labaj6219 ( R_234f6_b80ffc0, \43843 );
buf \U$labaj6220 ( R_234f8_b7ddf98, \43863 );
buf \U$labaj6221 ( R_234fa_b80c7f8, \43883 );
buf \U$labaj6222 ( R_234fc_b7de0e8, \43901 );
buf \U$labaj6223 ( R_234fe_b7de388, \43921 );
buf \U$labaj6224 ( R_23500_b7de430, \43940 );
buf \U$labaj6225 ( R_23502_b80c9f0, \43960 );
buf \U$labaj6226 ( R_23504_b7de580, \43980 );
buf \U$labaj6227 ( R_23506_b80ca98, \43998 );
buf \U$labaj6228 ( R_2350a_b7de820, \44017 );
buf \U$labaj6229 ( R_2350c_b7dea18, \44036 );
buf \U$labaj6230 ( R_2350e_b7dee08, \44054 );
buf \U$labaj6231 ( R_23510_b80cc90, \44073 );
buf \U$labaj6232 ( R_23512_b80cd38, \44093 );
buf \U$labaj6233 ( R_23514_b7df1f8, \44112 );
buf \U$labaj6234 ( R_23516_b80ce88, \44130 );
buf \U$labaj6235 ( R_23518_b7df348, \44150 );
buf \U$labaj6236 ( R_2351a_b7df540, \44170 );
buf \U$labaj6237 ( R_2351c_b80cf30, \44190 );
buf \U$labaj6238 ( R_23520_b7dfc78, \44209 );
buf \U$labaj6239 ( R_23522_b80d080, \44227 );
buf \U$labaj6240 ( R_23524_b80d278, \44245 );
buf \U$labaj6241 ( R_23526_b7dff18, \44264 );
buf \U$labaj6242 ( R_23528_b80d320, \44285 );
buf \U$labaj6243 ( R_2352a_b7e0068, \44305 );
buf \U$labaj6244 ( R_2352c_b80d5c0, \44325 );
buf \U$labaj6245 ( R_2352e_b7e01b8, \44343 );
buf \U$labaj6246 ( R_23530_b80d668, \44363 );
buf \U$labaj6247 ( R_23532_b7e0458, \44381 );
buf \U$labaj6248 ( R_23536_b7e05a8, \44399 );
buf \U$labaj6249 ( R_23538_b80d7b8, \44418 );
buf \U$labaj6250 ( R_2353a_b80de48, \44436 );
buf \U$labaj6251 ( R_2353c_b7e0998, \44456 );
buf \U$labaj6252 ( R_2353e_b7e0b90, \44474 );
buf \U$labaj6253 ( R_23540_b7e1178, \44492 );
buf \U$labaj6254 ( R_23542_b80e430, \44514 );
buf \U$labaj6255 ( R_23544_b80e628, \44535 );
buf \U$labaj6256 ( R_23546_b80e778, \44554 );
buf \U$labaj6257 ( R_23548_b7e1568, \44572 );
buf \U$labaj6258 ( R_2354c_b80e970, \44590 );
buf \U$labaj6259 ( R_2354e_b7e16b8, \44610 );
buf \U$labaj6260 ( R_23550_b80eb68, \44629 );
buf \U$labaj6261 ( R_23552_b7e1808, \44647 );
buf \U$labaj6262 ( R_2355c_b7e18b0, \44681 );
buf \U$labaj6263 ( R_23572_b805c58, \44701 );
buf \U$labaj6264 ( R_23588_b7e1958, \44720 );
buf \U$labaj6265 ( R_2359e_b80ed60, \44739 );
buf \U$labaj6266 ( R_235b4_95ad7d8, \44757 );
buf \U$labaj6267 ( R_235ca_b806438, \44778 );
buf \U$labaj6268 ( R_235d4_b7e1a00, \44797 );
buf \U$labaj6269 ( R_235d6_b80f000, \44816 );
buf \U$labaj6270 ( R_235d8_b7e1bf8, \44834 );
buf \U$labaj6271 ( R_235da_b7e1ca0, \44853 );
buf \U$labaj6272 ( R_2355e_b7e1e98, \44871 );
buf \U$labaj6273 ( R_23560_95ad9d0, \44890 );
buf \U$labaj6274 ( R_23562_b7e1f40, \44909 );
buf \U$labaj6275 ( R_23564_95adb20, \44927 );
buf \U$labaj6276 ( R_23566_b7e1fe8, \44945 );
buf \U$labaj6277 ( R_23568_b80f3f0, \44963 );
buf \U$labaj6278 ( R_2356a_b80f5e8, \44981 );
buf \U$labaj6279 ( R_2356c_b806630, \44999 );
buf \U$labaj6280 ( R_2356e_b7e2090, \45017 );
buf \U$labaj6281 ( R_23570_b80f690, \45035 );
buf \U$labaj6282 ( R_23574_b7e2138, \45053 );
buf \U$labaj6283 ( R_23576_b7e21e0, \45071 );
buf \U$labaj6284 ( R_23578_b7e23d8, \45089 );
buf \U$labaj6285 ( R_2357a_b7e2720, \45107 );
buf \U$labaj6286 ( R_2357c_b7e2870, \45125 );
buf \U$labaj6287 ( R_2357e_b7e29c0, \45143 );
buf \U$labaj6288 ( R_23580_b806828, \45161 );
buf \U$labaj6289 ( R_23582_b7e2a68, \45179 );
buf \U$labaj6290 ( R_23584_b7e2c60, \45197 );
buf \U$labaj6291 ( R_23586_b7e2f00, \45215 );
buf \U$labaj6292 ( R_2358a_b80f7e0, \45233 );
buf \U$labaj6293 ( R_2358c_96cb8e0, \45251 );
buf \U$labaj6294 ( R_2358e_b7e2fa8, \45269 );
buf \U$labaj6295 ( R_23590_b7e30f8, \45287 );
buf \U$labaj6296 ( R_23592_b806978, \45305 );
buf \U$labaj6297 ( R_23594_b807008, \45323 );
buf \U$labaj6298 ( R_23596_b7e32f0, \45342 );
buf \U$labaj6299 ( R_23598_b80fb28, \45360 );
buf \U$labaj6300 ( R_2359a_b7e3398, \45379 );
buf \U$labaj6301 ( R_2359c_b807698, \45397 );
buf \U$labaj6302 ( R_235a0_b7e34e8, \45415 );
buf \U$labaj6303 ( R_235a2_96cbb80, \45433 );
buf \U$labaj6304 ( R_235a4_b80fbd0, \45451 );
buf \U$labaj6305 ( R_235a6_96cc018, \45469 );
buf \U$labaj6306 ( R_235a8_95adf10, \45487 );
buf \U$labaj6307 ( R_235aa_b7e36e0, \45505 );
buf \U$labaj6308 ( R_235ac_b807890, \45523 );
buf \U$labaj6309 ( R_235ae_b7e3788, \45541 );
buf \U$labaj6310 ( R_235b0_b7e38d8, \45559 );
buf \U$labaj6311 ( R_235b2_b7e3ad0, \45577 );
buf \U$labaj6312 ( R_235b6_b7e3cc8, \45595 );
buf \U$labaj6313 ( R_235b8_b7e3f68, \45613 );
buf \U$labaj6314 ( R_235ba_b807f20, \45632 );
buf \U$labaj6315 ( R_235bc_b807fc8, \45650 );
buf \U$labaj6316 ( R_235be_b8101b8, \45668 );
buf \U$labaj6317 ( R_235c0_b7e40b8, \45686 );
buf \U$labaj6318 ( R_235c2_b7e4208, \45704 );
buf \U$labaj6319 ( R_235c4_b8105a8, \45722 );
buf \U$labaj6320 ( R_235c6_b810650, \45740 );
buf \U$labaj6321 ( R_235c8_96cc210, \45758 );
buf \U$labaj6322 ( R_235cc_b7e42b0, \45776 );
buf \U$labaj6323 ( R_235ce_b7e4400, \45794 );
buf \U$labaj6324 ( R_235d0_b7e4550, \45812 );
buf \U$labaj6325 ( R_235d2_b7e45f8, \45830 );
buf \U$labaj6326 ( R_235dc_b8106f8, \45863 );
buf \U$labaj6327 ( R_235f2_b7e46a0, \45882 );
buf \U$labaj6328 ( R_23608_b808118, \45899 );
buf \U$labaj6329 ( R_2361e_b7e47f0, \45917 );
buf \U$labaj6330 ( R_23634_b7e49e8, \45935 );
buf \U$labaj6331 ( R_2364a_b7dd860, \45954 );
buf \U$labaj6332 ( R_23654_95ae060, \45972 );
buf \U$labaj6333 ( R_23656_b7dd908, \45990 );
buf \U$labaj6334 ( R_23658_b7ddda0, \46007 );
buf \U$labaj6335 ( R_2365a_b7dde48, \46026 );
buf \U$labaj6336 ( R_235de_9637b50, \46043 );
buf \U$labaj6337 ( R_235e0_95ae1b0, \46062 );
buf \U$labaj6338 ( R_235e2_b7ddef0, \46080 );
buf \U$labaj6339 ( R_235e4_b7de238, \46098 );
buf \U$labaj6340 ( R_235e6_b7e4b38, \46115 );
buf \U$labaj6341 ( R_235e8_9637fe8, \46132 );
buf \U$labaj6342 ( R_235ea_b7de2e0, \46149 );
buf \U$labaj6343 ( R_235ec_b808310, \46166 );
buf \U$labaj6344 ( R_235ee_9638138, \46183 );
buf \U$labaj6345 ( R_235f0_96381e0, \46200 );
buf \U$labaj6346 ( R_235f4_b7e4d30, \46217 );
buf \U$labaj6347 ( R_235f6_96383d8, \46234 );
buf \U$labaj6348 ( R_235f8_b7de6d0, \46252 );
buf \U$labaj6349 ( R_235fa_9638480, \46269 );
buf \U$labaj6350 ( R_235fc_b7de8c8, \46286 );
buf \U$labaj6351 ( R_235fe_9638528, \46303 );
buf \U$labaj6352 ( R_23600_96385d0, \46320 );
buf \U$labaj6353 ( R_23602_b7de970, \46337 );
buf \U$labaj6354 ( R_23604_b7deac0, \46354 );
buf \U$labaj6355 ( R_23606_9638678, \46371 );
buf \U$labaj6356 ( R_2360a_96387c8, \46388 );
not \U$1 ( \8820 , RIde67cd8_3982);
not \U$2 ( \8821 , \8820 );
or \U$3 ( \8822 , RIde68638_3981, \8821 );
not \U$4 ( \8823 , \8822 );
and \U$5 ( \8824 , \8823 , RIde68f20_3980);
buf \U$6 ( \8825 , RIb79b518_270);
buf \U$7 ( \8826 , \8825 );
buf \U$8 ( \8827 , RIdbb8138_3227);
not \U$9 ( \8828 , \8827 );
not \U$10 ( \8829 , RIe549ef0_6842);
not \U$11 ( \8830 , \8829 );
not \U$12 ( \8831 , \8830 );
or \U$13 ( \8832 , RIe548ff0_6844, \8831 );
not \U$14 ( \8833 , \8832 );
not \U$15 ( \8834 , RIe5319e0_6884);
not \U$16 ( \8835 , \8834 );
not \U$17 ( \8836 , RIe549770_6843);
not \U$18 ( \8837 , \8836 );
nand \U$19 ( \8838 , \8835 , \8837 );
not \U$20 ( \8839 , \8838 );
and \U$21 ( \8840 , \8833 , \8839 );
not \U$22 ( \8841 , \8840 );
or \U$23 ( \8842 , \8828 , \8841 );
buf \U$24 ( \8843 , RIe4f85f0_6398);
not \U$25 ( \8844 , \8843 );
nand \U$26 ( \8845 , \8830 , RIe548ff0_6844);
not \U$27 ( \8846 , \8845 );
nand \U$28 ( \8847 , \8846 , \8839 );
not \U$29 ( \8848 , \8847 );
not \U$30 ( \8849 , \8848 );
or \U$31 ( \8850 , \8844 , \8849 );
nand \U$32 ( \8851 , \8842 , \8850 );
buf \U$33 ( \8852 , RIdaea590_2835);
not \U$34 ( \8853 , \8852 );
not \U$35 ( \8854 , \8837 );
or \U$36 ( \8855 , \8835 , \8854 );
not \U$37 ( \8856 , \8855 );
and \U$38 ( \8857 , \8833 , \8856 );
not \U$39 ( \8858 , \8857 );
or \U$40 ( \8859 , \8853 , \8858 );
buf \U$41 ( \8860 , RIe4301f0_6000);
not \U$42 ( \8861 , \8860 );
nand \U$43 ( \8862 , \8846 , \8856 );
not \U$44 ( \8863 , \8862 );
not \U$45 ( \8864 , \8863 );
or \U$46 ( \8865 , \8861 , \8864 );
nand \U$47 ( \8866 , \8859 , \8865 );
nor \U$48 ( \8867 , \8851 , \8866 );
buf \U$49 ( \8868 , RIde3d1e0_4027);
not \U$50 ( \8869 , \8868 );
not \U$51 ( \8870 , \8834 );
not \U$52 ( \8871 , \8870 );
or \U$53 ( \8872 , \8837 , \8871 );
not \U$54 ( \8873 , \8872 );
not \U$55 ( \8874 , RIe548ff0_6844);
or \U$56 ( \8875 , \8830 , \8874 );
not \U$57 ( \8876 , \8875 );
nand \U$58 ( \8877 , \8873 , \8876 );
not \U$59 ( \8878 , \8877 );
not \U$60 ( \8879 , \8878 );
or \U$61 ( \8880 , \8869 , \8879 );
buf \U$62 ( \8881 , RIe00b330_4420);
not \U$63 ( \8882 , \8881 );
or \U$64 ( \8883 , RIe5319e0_6884, RIe549770_6843);
not \U$65 ( \8884 , \8883 );
nand \U$66 ( \8885 , \8884 , \8846 );
not \U$67 ( \8886 , \8885 );
not \U$68 ( \8887 , \8886 );
or \U$69 ( \8888 , \8882 , \8887 );
nand \U$70 ( \8889 , \8880 , \8888 );
nand \U$71 ( \8890 , \8876 , \8856 );
not \U$72 ( \8891 , \8890 );
not \U$73 ( \8892 , \8891 );
buf \U$74 ( \8893 , RIe160838_5254);
not \U$75 ( \8894 , \8893 );
or \U$76 ( \8895 , \8892 , \8894 );
buf \U$77 ( \8896 , RIe0d49f0_4816);
not \U$78 ( \8897 , \8896 );
nand \U$79 ( \8898 , \8846 , \8873 );
not \U$80 ( \8899 , \8898 );
not \U$81 ( \8900 , \8899 );
or \U$82 ( \8901 , \8897 , \8900 );
nand \U$83 ( \8902 , \8895 , \8901 );
nor \U$84 ( \8903 , \8889 , \8902 );
buf \U$85 ( \8904 , RIda11c00_2446);
not \U$86 ( \8905 , \8829 );
not \U$87 ( \8906 , RIe548ff0_6844);
not \U$88 ( \8907 , \8906 );
or \U$89 ( \8908 , \8905 , \8907 );
not \U$90 ( \8909 , \8908 );
and \U$91 ( \8910 , \8909 , \8839 );
not \U$92 ( \8911 , \8910 );
not \U$93 ( \8912 , \8911 );
buf \U$94 ( \8913 , \8912 );
nand \U$95 ( \8914 , \8904 , \8913 );
buf \U$96 ( \8915 , RIe269120_5609);
nand \U$97 ( \8916 , \8839 , \8876 );
not \U$98 ( \8917 , \8916 );
not \U$99 ( \8918 , \8917 );
not \U$100 ( \8919 , \8918 );
nand \U$101 ( \8920 , \8915 , \8919 );
buf \U$102 ( \8921 , RId958f08_2058);
nand \U$103 ( \8922 , \8909 , \8856 );
not \U$104 ( \8923 , \8922 );
not \U$105 ( \8924 , \8923 );
not \U$106 ( \8925 , \8924 );
and \U$107 ( \8926 , \8921 , \8925 );
buf \U$108 ( \8927 , RId888d80_1669);
and \U$109 ( \8928 , \8833 , \8873 );
not \U$110 ( \8929 , \8928 );
not \U$111 ( \8930 , \8929 );
and \U$112 ( \8931 , \8927 , \8930 );
nor \U$113 ( \8932 , \8926 , \8931 );
nand \U$114 ( \8933 , \8914 , \8920 , \8932 );
buf \U$115 ( \8934 , RIdc6ed48_3642);
nand \U$116 ( \8935 , \8884 , \8876 );
not \U$117 ( \8936 , \8935 );
not \U$118 ( \8937 , \8936 );
not \U$119 ( \8938 , \8937 );
and \U$120 ( \8939 , \8934 , \8938 );
buf \U$121 ( \8940 , RIe5c2e08_6791);
nand \U$122 ( \8941 , \8909 , \8884 );
not \U$123 ( \8942 , \8941 );
not \U$124 ( \8943 , \8942 );
not \U$125 ( \8944 , \8943 );
and \U$126 ( \8945 , \8940 , \8944 );
nor \U$127 ( \8946 , \8939 , \8945 );
buf \U$128 ( \8947 , RId6f3a80_883);
nand \U$129 ( \8948 , \8909 , \8873 );
not \U$130 ( \8949 , \8948 );
not \U$131 ( \8950 , \8949 );
not \U$132 ( \8951 , \8950 );
and \U$133 ( \8952 , \8947 , \8951 );
buf \U$134 ( \8953 , RId7bf4e0_1272);
nand \U$135 ( \8954 , \8833 , \8884 );
not \U$136 ( \8955 , \8954 );
not \U$137 ( \8956 , \8955 );
not \U$138 ( \8957 , \8956 );
and \U$139 ( \8958 , \8953 , \8957 );
nor \U$140 ( \8959 , \8952 , \8958 );
nand \U$141 ( \8960 , \8946 , \8959 );
nor \U$142 ( \8961 , \8933 , \8960 );
nand \U$143 ( \8962 , \8867 , \8903 , \8961 );
not \U$144 ( \8963 , \8962 );
not \U$145 ( \8964 , RIb7b93b0_251);
xnor \U$146 ( \8965 , \8963 , \8964 );
buf \U$147 ( \8966 , RIdba4548_3251);
not \U$148 ( \8967 , \8966 );
not \U$149 ( \8968 , \8840 );
or \U$150 ( \8969 , \8967 , \8968 );
buf \U$151 ( \8970 , RIe4fa198_6396);
not \U$152 ( \8971 , \8970 );
not \U$153 ( \8972 , \8847 );
not \U$154 ( \8973 , \8972 );
or \U$155 ( \8974 , \8971 , \8973 );
nand \U$156 ( \8975 , \8969 , \8974 );
buf \U$157 ( \8976 , RIdaebc88_2833);
not \U$158 ( \8977 , \8976 );
or \U$159 ( \8978 , \8977 , \8858 );
buf \U$160 ( \8979 , RIe431ac8_5998);
not \U$161 ( \8980 , \8979 );
not \U$162 ( \8981 , \8862 );
not \U$163 ( \8982 , \8981 );
or \U$164 ( \8983 , \8980 , \8982 );
nand \U$165 ( \8984 , \8978 , \8983 );
nor \U$166 ( \8985 , \8975 , \8984 );
buf \U$167 ( \8986 , RIde3ed88_4025);
not \U$168 ( \8987 , \8986 );
not \U$169 ( \8988 , \8878 );
or \U$170 ( \8989 , \8987 , \8988 );
buf \U$171 ( \8990 , RIe00ce60_4418);
not \U$172 ( \8991 , \8990 );
not \U$173 ( \8992 , \8886 );
or \U$174 ( \8993 , \8991 , \8992 );
nand \U$175 ( \8994 , \8989 , \8993 );
not \U$176 ( \8995 , \8891 );
buf \U$177 ( \8996 , RIe1615d0_5253);
not \U$178 ( \8997 , \8996 );
or \U$179 ( \8998 , \8995 , \8997 );
buf \U$180 ( \8999 , RIe0d62c8_4814);
not \U$181 ( \9000 , \8999 );
not \U$182 ( \9001 , \8898 );
not \U$183 ( \9002 , \9001 );
or \U$184 ( \9003 , \9000 , \9002 );
nand \U$185 ( \9004 , \8998 , \9003 );
nor \U$186 ( \9005 , \8994 , \9004 );
buf \U$187 ( \9006 , RIda13640_2444);
buf \U$188 ( \9007 , \8912 );
nand \U$189 ( \9008 , \9006 , \9007 );
buf \U$190 ( \9009 , RIe26a7a0_5607);
nand \U$191 ( \9010 , \9009 , \8919 );
buf \U$192 ( \9011 , RId95a600_2056);
not \U$193 ( \9012 , \8924 );
and \U$194 ( \9013 , \9011 , \9012 );
buf \U$195 ( \9014 , RId88a478_1667);
not \U$196 ( \9015 , \8928 );
not \U$197 ( \9016 , \9015 );
and \U$198 ( \9017 , \9014 , \9016 );
nor \U$199 ( \9018 , \9013 , \9017 );
nand \U$200 ( \9019 , \9008 , \9010 , \9018 );
buf \U$201 ( \9020 , RIdc70800_3640);
not \U$202 ( \9021 , \8935 );
not \U$203 ( \9022 , \9021 );
not \U$204 ( \9023 , \9022 );
and \U$205 ( \9024 , \9020 , \9023 );
buf \U$206 ( \9025 , RIe5c4500_6789);
not \U$207 ( \9026 , \8942 );
not \U$208 ( \9027 , \9026 );
and \U$209 ( \9028 , \9025 , \9027 );
nor \U$210 ( \9029 , \9024 , \9028 );
buf \U$211 ( \9030 , RId6f5100_881);
not \U$212 ( \9031 , \8949 );
not \U$213 ( \9032 , \9031 );
and \U$214 ( \9033 , \9030 , \9032 );
buf \U$215 ( \9034 , RId7c0e30_1270);
not \U$216 ( \9035 , \8954 );
not \U$217 ( \9036 , \9035 );
not \U$218 ( \9037 , \9036 );
and \U$219 ( \9038 , \9034 , \9037 );
nor \U$220 ( \9039 , \9033 , \9038 );
nand \U$221 ( \9040 , \9029 , \9039 );
nor \U$222 ( \9041 , \9019 , \9040 );
nand \U$223 ( \9042 , \8985 , \9005 , \9041 );
not \U$224 ( \9043 , \9042 );
not \U$225 ( \9044 , RIb7b94a0_249);
xnor \U$226 ( \9045 , \9043 , \9044 );
buf \U$227 ( \9046 , RIdbb7328_3228);
not \U$228 ( \9047 , \9046 );
or \U$229 ( \9048 , \9047 , \8841 );
buf \U$230 ( \9049 , RIe4f7a38_6399);
not \U$231 ( \9050 , \9049 );
not \U$232 ( \9051 , \8972 );
or \U$233 ( \9052 , \9050 , \9051 );
nand \U$234 ( \9053 , \9048 , \9052 );
buf \U$235 ( \9054 , RIdae97f8_2836);
not \U$236 ( \9055 , \9054 );
or \U$237 ( \9056 , \9055 , \8858 );
buf \U$238 ( \9057 , RIe42f4d0_6001);
not \U$239 ( \9058 , \9057 );
not \U$240 ( \9059 , \8863 );
or \U$241 ( \9060 , \9058 , \9059 );
nand \U$242 ( \9061 , \9056 , \9060 );
nor \U$243 ( \9062 , \9053 , \9061 );
buf \U$244 ( \9063 , RIde3c448_4028);
not \U$245 ( \9064 , \9063 );
not \U$246 ( \9065 , \8878 );
or \U$247 ( \9066 , \9064 , \9065 );
buf \U$248 ( \9067 , RIe00a598_4421);
not \U$249 ( \9068 , \9067 );
or \U$250 ( \9069 , \9068 , \8887 );
nand \U$251 ( \9070 , \9066 , \9069 );
not \U$252 ( \9071 , \8891 );
buf \U$253 ( \9072 , RIe172718_5244);
not \U$254 ( \9073 , \9072 );
or \U$255 ( \9074 , \9071 , \9073 );
buf \U$256 ( \9075 , RIe0d3dc0_4817);
not \U$257 ( \9076 , \9075 );
not \U$258 ( \9077 , \8899 );
or \U$259 ( \9078 , \9076 , \9077 );
nand \U$260 ( \9079 , \9074 , \9078 );
nor \U$261 ( \9080 , \9070 , \9079 );
buf \U$262 ( \9081 , RIda10df0_2447);
not \U$263 ( \9082 , \9081 );
not \U$264 ( \9083 , \8913 );
or \U$265 ( \9084 , \9082 , \9083 );
buf \U$266 ( \9085 , RIe268568_5610);
not \U$267 ( \9086 , \9085 );
not \U$268 ( \9087 , \8919 );
or \U$269 ( \9088 , \9086 , \9087 );
buf \U$270 ( \9089 , RId9582d8_2059);
not \U$271 ( \9090 , \8923 );
not \U$272 ( \9091 , \9090 );
and \U$273 ( \9092 , \9089 , \9091 );
buf \U$274 ( \9093 , RId888240_1670);
not \U$275 ( \9094 , \9015 );
and \U$276 ( \9095 , \9093 , \9094 );
nor \U$277 ( \9096 , \9092 , \9095 );
nand \U$278 ( \9097 , \9084 , \9088 , \9096 );
buf \U$279 ( \9098 , RIdc6e280_3643);
not \U$280 ( \9099 , \8936 );
not \U$281 ( \9100 , \9099 );
and \U$282 ( \9101 , \9098 , \9100 );
buf \U$283 ( \9102 , RIe5c22c8_6792);
not \U$284 ( \9103 , \8942 );
not \U$285 ( \9104 , \9103 );
and \U$286 ( \9105 , \9102 , \9104 );
nor \U$287 ( \9106 , \9101 , \9105 );
buf \U$288 ( \9107 , RId7064a0_859);
not \U$289 ( \9108 , \8948 );
not \U$290 ( \9109 , \9108 );
not \U$291 ( \9110 , \9109 );
and \U$292 ( \9111 , \9107 , \9110 );
buf \U$293 ( \9112 , RId7be838_1273);
not \U$294 ( \9113 , \9036 );
and \U$295 ( \9114 , \9112 , \9113 );
nor \U$296 ( \9115 , \9111 , \9114 );
nand \U$297 ( \9116 , \9106 , \9115 );
nor \U$298 ( \9117 , \9097 , \9116 );
nand \U$299 ( \9118 , \9062 , \9080 , \9117 );
not \U$300 ( \9119 , RIb7af720_252);
xnor \U$301 ( \9120 , \9118 , \9119 );
buf \U$302 ( \9121 , RIdbb6518_3229);
not \U$303 ( \9122 , \9121 );
or \U$304 ( \9123 , \9122 , \8841 );
buf \U$305 ( \9124 , RIe4f6ef8_6400);
not \U$306 ( \9125 , \9124 );
not \U$307 ( \9126 , \8972 );
or \U$308 ( \9127 , \9125 , \9126 );
nand \U$309 ( \9128 , \9123 , \9127 );
buf \U$310 ( \9129 , RIdae8a60_2837);
not \U$311 ( \9130 , \9129 );
or \U$312 ( \9131 , \9130 , \8858 );
buf \U$313 ( \9132 , RIe42e8a0_6002);
not \U$314 ( \9133 , \9132 );
or \U$315 ( \9134 , \9133 , \9059 );
nand \U$316 ( \9135 , \9131 , \9134 );
nor \U$317 ( \9136 , \9128 , \9135 );
buf \U$318 ( \9137 , RIde3b728_4029);
not \U$319 ( \9138 , \9137 );
not \U$320 ( \9139 , \8877 );
not \U$321 ( \9140 , \9139 );
or \U$322 ( \9141 , \9138 , \9140 );
buf \U$323 ( \9142 , RIe009710_4422);
not \U$324 ( \9143 , \9142 );
or \U$325 ( \9144 , \9143 , \8992 );
nand \U$326 ( \9145 , \9141 , \9144 );
not \U$327 ( \9146 , \8891 );
buf \U$328 ( \9147 , RIe163e20_5250);
not \U$329 ( \9148 , \9147 );
or \U$330 ( \9149 , \9146 , \9148 );
buf \U$331 ( \9150 , RIe0d2e48_4818);
not \U$332 ( \9151 , \9150 );
or \U$333 ( \9152 , \9151 , \8900 );
nand \U$334 ( \9153 , \9149 , \9152 );
nor \U$335 ( \9154 , \9145 , \9153 );
buf \U$336 ( \9155 , RIda101c0_2448);
nand \U$337 ( \9156 , \9155 , \8913 );
buf \U$338 ( \9157 , RIe2679b0_5611);
nand \U$339 ( \9158 , \9157 , \8919 );
buf \U$340 ( \9159 , RId957720_2060);
not \U$341 ( \9160 , \8923 );
not \U$342 ( \9161 , \9160 );
and \U$343 ( \9162 , \9159 , \9161 );
buf \U$344 ( \9163 , RId89b638_1645);
not \U$345 ( \9164 , \9015 );
and \U$346 ( \9165 , \9163 , \9164 );
nor \U$347 ( \9166 , \9162 , \9165 );
nand \U$348 ( \9167 , \9156 , \9158 , \9166 );
buf \U$349 ( \9168 , RIdc6d740_3644);
not \U$350 ( \9169 , \8936 );
not \U$351 ( \9170 , \9169 );
and \U$352 ( \9171 , \9168 , \9170 );
buf \U$353 ( \9172 , RIe5c1710_6793);
not \U$354 ( \9173 , \9103 );
and \U$355 ( \9174 , \9172 , \9173 );
nor \U$356 ( \9175 , \9171 , \9174 );
buf \U$357 ( \9176 , RId705780_860);
not \U$358 ( \9177 , \9108 );
not \U$359 ( \9178 , \9177 );
and \U$360 ( \9179 , \9176 , \9178 );
buf \U$361 ( \9180 , RId7d2338_1248);
not \U$362 ( \9181 , \9035 );
not \U$363 ( \9182 , \9181 );
and \U$364 ( \9183 , \9180 , \9182 );
nor \U$365 ( \9184 , \9179 , \9183 );
nand \U$366 ( \9185 , \9175 , \9184 );
nor \U$367 ( \9186 , \9167 , \9185 );
nand \U$368 ( \9187 , \9136 , \9154 , \9186 );
not \U$369 ( \9188 , RIb7af6a8_253);
xnor \U$370 ( \9189 , \9187 , \9188 );
nor \U$371 ( \9190 , \9120 , \9189 );
nand \U$372 ( \9191 , \8965 , \9045 , \9190 );
not \U$373 ( \9192 , \9191 );
buf \U$374 ( \9193 , RIe4faf30_6395);
not \U$375 ( \9194 , \9193 );
or \U$376 ( \9195 , \9194 , \8973 );
buf \U$377 ( \9196 , RIdba51f0_3250);
not \U$378 ( \9197 , \9196 );
or \U$379 ( \9198 , \9197 , \8968 );
nand \U$380 ( \9199 , \9195 , \9198 );
buf \U$381 ( \9200 , RIe4326f8_5997);
not \U$382 ( \9201 , \9200 );
not \U$383 ( \9202 , \8863 );
or \U$384 ( \9203 , \9201 , \9202 );
buf \U$385 ( \9204 , RIdad5d70_2860);
not \U$386 ( \9205 , \9204 );
not \U$387 ( \9206 , \8857 );
or \U$388 ( \9207 , \9205 , \9206 );
nand \U$389 ( \9208 , \9203 , \9207 );
nor \U$390 ( \9209 , \9199 , \9208 );
buf \U$391 ( \9210 , RIde3fb20_4024);
and \U$392 ( \9211 , \9210 , \9139 );
buf \U$393 ( \9212 , RIe00db80_4417);
not \U$394 ( \9213 , \8885 );
and \U$395 ( \9214 , \9212 , \9213 );
or \U$396 ( \9215 , \9211 , \9214 );
buf \U$397 ( \9216 , RIe164b40_5249);
not \U$398 ( \9217 , \9216 );
or \U$399 ( \9218 , \9071 , \9217 );
buf \U$400 ( \9219 , RIe0d6fe8_4813);
not \U$401 ( \9220 , \9219 );
not \U$402 ( \9221 , \9001 );
or \U$403 ( \9222 , \9220 , \9221 );
nand \U$404 ( \9223 , \9218 , \9222 );
nor \U$405 ( \9224 , \9215 , \9223 );
buf \U$406 ( \9225 , RIda143d8_2443);
not \U$407 ( \9226 , \9225 );
or \U$408 ( \9227 , \9226 , \8911 );
buf \U$409 ( \9228 , RIe26b2e0_5606);
nand \U$410 ( \9229 , \9228 , \8919 );
buf \U$411 ( \9230 , RId95b1b8_2055);
not \U$412 ( \9231 , \8924 );
and \U$413 ( \9232 , \9230 , \9231 );
buf \U$414 ( \9233 , RId88b030_1666);
not \U$415 ( \9234 , \8928 );
not \U$416 ( \9235 , \9234 );
and \U$417 ( \9236 , \9233 , \9235 );
nor \U$418 ( \9237 , \9232 , \9236 );
nand \U$419 ( \9238 , \9227 , \9229 , \9237 );
buf \U$420 ( \9239 , RIdc71610_3639);
not \U$421 ( \9240 , \9099 );
and \U$422 ( \9241 , \9239 , \9240 );
buf \U$423 ( \9242 , RIe5c4fc8_6788);
not \U$424 ( \9243 , \8942 );
not \U$425 ( \9244 , \9243 );
and \U$426 ( \9245 , \9242 , \9244 );
nor \U$427 ( \9246 , \9241 , \9245 );
buf \U$428 ( \9247 , RId6f5cb8_880);
not \U$429 ( \9248 , \9108 );
not \U$430 ( \9249 , \9248 );
and \U$431 ( \9250 , \9247 , \9249 );
buf \U$432 ( \9251 , RId7c1b50_1269);
not \U$433 ( \9252 , \8955 );
not \U$434 ( \9253 , \9252 );
and \U$435 ( \9254 , \9251 , \9253 );
nor \U$436 ( \9255 , \9250 , \9254 );
nand \U$437 ( \9256 , \9246 , \9255 );
nor \U$438 ( \9257 , \9238 , \9256 );
nand \U$439 ( \9258 , \9209 , \9224 , \9257 );
not \U$440 ( \9259 , \9258 );
not \U$441 ( \9260 , RIb7b9518_248);
xnor \U$442 ( \9261 , \9259 , \9260 );
buf \U$443 ( \9262 , RIdba3828_3252);
not \U$444 ( \9263 , \9262 );
or \U$445 ( \9264 , \9263 , \8968 );
buf \U$446 ( \9265 , RIe4f9388_6397);
not \U$447 ( \9266 , \9265 );
or \U$448 ( \9267 , \9266 , \8973 );
nand \U$449 ( \9268 , \9264 , \9267 );
buf \U$450 ( \9269 , RIdaeb0d0_2834);
not \U$451 ( \9270 , \9269 );
or \U$452 ( \9271 , \9270 , \9206 );
buf \U$453 ( \9272 , RIe430e20_5999);
not \U$454 ( \9273 , \9272 );
or \U$455 ( \9274 , \9273 , \8982 );
nand \U$456 ( \9275 , \9271 , \9274 );
nor \U$457 ( \9276 , \9268 , \9275 );
buf \U$458 ( \9277 , RIde3df00_4026);
not \U$459 ( \9278 , \9277 );
not \U$460 ( \9279 , \9139 );
or \U$461 ( \9280 , \9278 , \9279 );
buf \U$462 ( \9281 , RIe00c0c8_4419);
not \U$463 ( \9282 , \9281 );
or \U$464 ( \9283 , \9282 , \8887 );
nand \U$465 ( \9284 , \9280 , \9283 );
not \U$466 ( \9285 , \8891 );
buf \U$467 ( \9286 , RIe163088_5251);
not \U$468 ( \9287 , \9286 );
or \U$469 ( \9288 , \9285 , \9287 );
buf \U$470 ( \9289 , RIe0d55a8_4815);
not \U$471 ( \9290 , \9289 );
not \U$472 ( \9291 , \9001 );
or \U$473 ( \9292 , \9290 , \9291 );
nand \U$474 ( \9293 , \9288 , \9292 );
nor \U$475 ( \9294 , \9284 , \9293 );
buf \U$476 ( \9295 , RIda12920_2445);
nand \U$477 ( \9296 , \9295 , \8913 );
buf \U$478 ( \9297 , RIe269c60_5608);
nand \U$479 ( \9298 , \9297 , \8919 );
buf \U$480 ( \9299 , RId959a48_2057);
not \U$481 ( \9300 , \9160 );
and \U$482 ( \9301 , \9299 , \9300 );
buf \U$483 ( \9302 , RId889938_1668);
not \U$484 ( \9303 , \9234 );
and \U$485 ( \9304 , \9302 , \9303 );
nor \U$486 ( \9305 , \9301 , \9304 );
nand \U$487 ( \9306 , \9296 , \9298 , \9305 );
buf \U$488 ( \9307 , RIdc6f9f0_3641);
not \U$489 ( \9308 , \9022 );
and \U$490 ( \9309 , \9307 , \9308 );
buf \U$491 ( \9310 , RIe5c3948_6790);
not \U$492 ( \9311 , \8942 );
not \U$493 ( \9312 , \9311 );
and \U$494 ( \9313 , \9310 , \9312 );
nor \U$495 ( \9314 , \9309 , \9313 );
buf \U$496 ( \9315 , RId6f4638_882);
not \U$497 ( \9316 , \8949 );
not \U$498 ( \9317 , \9316 );
and \U$499 ( \9318 , \9315 , \9317 );
buf \U$500 ( \9319 , RId7c0110_1271);
not \U$501 ( \9320 , \9181 );
and \U$502 ( \9321 , \9319 , \9320 );
nor \U$503 ( \9322 , \9318 , \9321 );
nand \U$504 ( \9323 , \9314 , \9322 );
nor \U$505 ( \9324 , \9306 , \9323 );
nand \U$506 ( \9325 , \9276 , \9294 , \9324 );
not \U$507 ( \9326 , \9325 );
not \U$508 ( \9327 , RIb7b9428_250);
xnor \U$509 ( \9328 , \9326 , \9327 );
nand \U$510 ( \9329 , \9261 , \9328 );
not \U$511 ( \9330 , \9329 );
buf \U$512 ( \9331 , RIdba6bb8_3248);
not \U$513 ( \9332 , \9331 );
or \U$514 ( \9333 , \9332 , \8968 );
buf \U$515 ( \9334 , RIe4fc9e8_6393);
not \U$516 ( \9335 , \9334 );
or \U$517 ( \9336 , \9335 , \8973 );
nand \U$518 ( \9337 , \9333 , \9336 );
buf \U$519 ( \9338 , RIdad7918_2858);
not \U$520 ( \9339 , \9338 );
or \U$521 ( \9340 , \9339 , \9206 );
buf \U$522 ( \9341 , RIe4340c0_5995);
not \U$523 ( \9342 , \9341 );
or \U$524 ( \9343 , \9342 , \8982 );
nand \U$525 ( \9344 , \9340 , \9343 );
nor \U$526 ( \9345 , \9337 , \9344 );
buf \U$527 ( \9346 , RIde415d8_4022);
and \U$528 ( \9347 , \9346 , \9139 );
buf \U$529 ( \9348 , RIe00f6b0_4415);
and \U$530 ( \9349 , \9348 , \9213 );
or \U$531 ( \9350 , \9347 , \9349 );
not \U$532 ( \9351 , \8892 );
not \U$533 ( \9352 , \9351 );
buf \U$534 ( \9353 , RIe162368_5252);
not \U$535 ( \9354 , \9353 );
or \U$536 ( \9355 , \9352 , \9354 );
buf \U$537 ( \9356 , RIe0d89b0_4811);
not \U$538 ( \9357 , \9356 );
or \U$539 ( \9358 , \9357 , \9002 );
nand \U$540 ( \9359 , \9355 , \9358 );
nor \U$541 ( \9360 , \9350 , \9359 );
buf \U$542 ( \9361 , RIda15da0_2441);
buf \U$543 ( \9362 , \8912 );
nand \U$544 ( \9363 , \9361 , \9362 );
buf \U$545 ( \9364 , RIe26ce10_5604);
nand \U$546 ( \9365 , \9364 , \8919 );
buf \U$547 ( \9366 , RId95c8b0_2053);
not \U$548 ( \9367 , \8924 );
and \U$549 ( \9368 , \9366 , \9367 );
buf \U$550 ( \9369 , RId88c728_1664);
not \U$551 ( \9370 , \9234 );
and \U$552 ( \9371 , \9369 , \9370 );
nor \U$553 ( \9372 , \9368 , \9371 );
nand \U$554 ( \9373 , \9363 , \9365 , \9372 );
buf \U$555 ( \9374 , RIdd731d8_3637);
buf \U$556 ( \9375 , \9021 );
nand \U$557 ( \9376 , \9374 , \9375 );
buf \U$558 ( \9377 , RId7c3590_1267);
not \U$559 ( \9378 , \8956 );
nand \U$560 ( \9379 , \9377 , \9378 );
buf \U$561 ( \9380 , RIe5c6738_6786);
not \U$562 ( \9381 , \8941 );
not \U$563 ( \9382 , \9381 );
not \U$564 ( \9383 , \9382 );
and \U$565 ( \9384 , \9380 , \9383 );
buf \U$566 ( \9385 , RId6f73b0_878);
and \U$567 ( \9386 , \9385 , \9108 );
nor \U$568 ( \9387 , \9384 , \9386 );
nand \U$569 ( \9388 , \9376 , \9379 , \9387 );
nor \U$570 ( \9389 , \9373 , \9388 );
nand \U$571 ( \9390 , \9345 , \9360 , \9389 );
not \U$572 ( \9391 , \9390 );
not \U$573 ( \9392 , RIb7b9608_246);
xnor \U$574 ( \9393 , \9391 , \9392 );
buf \U$575 ( \9394 , RIdba5e98_3249);
not \U$576 ( \9395 , \9394 );
or \U$577 ( \9396 , \9395 , \8968 );
buf \U$578 ( \9397 , RIe4fbcc8_6394);
not \U$579 ( \9398 , \9397 );
or \U$580 ( \9399 , \9398 , \8847 );
nand \U$581 ( \9400 , \9396 , \9399 );
buf \U$582 ( \9401 , RIdad6b80_2859);
not \U$583 ( \9402 , \9401 );
or \U$584 ( \9403 , \9402 , \9206 );
buf \U$585 ( \9404 , RIe4333a0_5996);
not \U$586 ( \9405 , \9404 );
or \U$587 ( \9406 , \9405 , \9202 );
nand \U$588 ( \9407 , \9403 , \9406 );
nor \U$589 ( \9408 , \9400 , \9407 );
buf \U$590 ( \9409 , RIde408b8_4023);
not \U$591 ( \9410 , \9409 );
not \U$592 ( \9411 , \8877 );
not \U$593 ( \9412 , \9411 );
or \U$594 ( \9413 , \9410 , \9412 );
buf \U$595 ( \9414 , RIe00e918_4416);
not \U$596 ( \9415 , \9414 );
or \U$597 ( \9416 , \9415 , \8992 );
nand \U$598 ( \9417 , \9413 , \9416 );
buf \U$599 ( \9418 , RIe1658d8_5248);
not \U$600 ( \9419 , \9418 );
or \U$601 ( \9420 , \9146 , \9419 );
buf \U$602 ( \9421 , RIe0d7d08_4812);
not \U$603 ( \9422 , \9421 );
not \U$604 ( \9423 , \9001 );
or \U$605 ( \9424 , \9422 , \9423 );
nand \U$606 ( \9425 , \9420 , \9424 );
nor \U$607 ( \9426 , \9417 , \9425 );
buf \U$608 ( \9427 , RIda150f8_2442);
buf \U$609 ( \9428 , \8912 );
nand \U$610 ( \9429 , \9427 , \9428 );
buf \U$611 ( \9430 , RIe26c000_5605);
nand \U$612 ( \9431 , \9430 , \8919 );
buf \U$613 ( \9432 , RId95bcf8_2054);
not \U$614 ( \9433 , \8924 );
and \U$615 ( \9434 , \9432 , \9433 );
buf \U$616 ( \9435 , RId88bbe8_1665);
not \U$617 ( \9436 , \8929 );
and \U$618 ( \9437 , \9435 , \9436 );
nor \U$619 ( \9438 , \9434 , \9437 );
nand \U$620 ( \9439 , \9429 , \9431 , \9438 );
buf \U$621 ( \9440 , RIdc72420_3638);
not \U$622 ( \9441 , \8936 );
not \U$623 ( \9442 , \9441 );
and \U$624 ( \9443 , \9440 , \9442 );
buf \U$625 ( \9444 , RIe5c5bf8_6787);
not \U$626 ( \9445 , \9381 );
not \U$627 ( \9446 , \9445 );
and \U$628 ( \9447 , \9444 , \9446 );
nor \U$629 ( \9448 , \9443 , \9447 );
buf \U$630 ( \9449 , RId6f68e8_879);
not \U$631 ( \9450 , \8949 );
not \U$632 ( \9451 , \9450 );
and \U$633 ( \9452 , \9449 , \9451 );
buf \U$634 ( \9453 , RId7c2870_1268);
and \U$635 ( \9454 , \9453 , \8955 );
nor \U$636 ( \9455 , \9452 , \9454 );
nand \U$637 ( \9456 , \9448 , \9455 );
nor \U$638 ( \9457 , \9439 , \9456 );
nand \U$639 ( \9458 , \9408 , \9426 , \9457 );
not \U$640 ( \9459 , \9458 );
not \U$641 ( \9460 , RIb7b9590_247);
xnor \U$642 ( \9461 , \9459 , \9460 );
and \U$643 ( \9462 , \9330 , \9393 , \9461 );
not \U$644 ( \9463 , RIe5349b0_6879);
not \U$645 ( \9464 , \9463 );
and \U$646 ( \9465 , \9464 , \9411 );
not \U$647 ( \9466 , \8885 );
not \U$648 ( \9467 , RIe5341b8_6880);
not \U$649 ( \9468 , \9467 );
and \U$650 ( \9469 , \9466 , \9468 );
nor \U$651 ( \9470 , \9465 , \9469 );
not \U$652 ( \9471 , RIe5339c0_6881);
not \U$653 ( \9472 , \9471 );
not \U$654 ( \9473 , \8892 );
and \U$655 ( \9474 , \9472 , \9473 );
not \U$656 ( \9475 , RIe5331c8_6882);
not \U$657 ( \9476 , \9475 );
and \U$658 ( \9477 , \8919 , \9476 );
nor \U$659 ( \9478 , \9474 , \9477 );
not \U$660 ( \9479 , RIe5329d0_6883);
buf \U$661 ( \9480 , \9479 );
or \U$662 ( \9481 , \9480 , \9026 );
not \U$663 ( \9482 , RIeb72150_6905);
or \U$664 ( \9483 , \9482 , \8973 );
nand \U$665 ( \9484 , \9481 , \9483 );
not \U$666 ( \9485 , RIe5359a0_6877);
or \U$667 ( \9486 , \9485 , \8858 );
not \U$668 ( \9487 , RIe5351a8_6878);
or \U$669 ( \9488 , \9487 , \8968 );
nand \U$670 ( \9489 , \9486 , \9488 );
nor \U$671 ( \9490 , \9484 , \9489 );
nand \U$672 ( \9491 , \9470 , \9478 , \9490 );
not \U$673 ( \9492 , RIeab7d00_6896);
or \U$674 ( \9493 , \9492 , \9160 );
not \U$675 ( \9494 , RIeab78c8_6895);
not \U$676 ( \9495 , \8910 );
or \U$677 ( \9496 , \9494 , \9495 );
nand \U$678 ( \9497 , \9493 , \9496 );
not \U$679 ( \9498 , RIeab6518_6891);
or \U$680 ( \9499 , \9498 , \9252 );
not \U$681 ( \9500 , RIeacfa18_6902);
or \U$682 ( \9501 , \9500 , \8929 );
nand \U$683 ( \9502 , \9499 , \9501 );
nor \U$684 ( \9503 , \9497 , \9502 );
not \U$685 ( \9504 , RIeab80c0_6897);
or \U$686 ( \9505 , \9504 , \8864 );
not \U$687 ( \9506 , RIeb352c8_6904);
or \U$688 ( \9507 , \9506 , \9031 );
nand \U$689 ( \9508 , \9505 , \9507 );
not \U$690 ( \9509 , RIea94af8_6890);
or \U$691 ( \9510 , \9509 , \9169 );
not \U$692 ( \9511 , RIeab87c8_6898);
or \U$693 ( \9512 , \9511 , \9077 );
nand \U$694 ( \9513 , \9510 , \9512 );
nor \U$695 ( \9514 , \9508 , \9513 );
nand \U$696 ( \9515 , \9503 , \9514 );
nor \U$697 ( \9516 , \9491 , \9515 );
not \U$698 ( \9517 , \9516 );
buf \U$699 ( \9518 , RIe15c260_5259);
not \U$700 ( \9519 , \9518 );
not \U$701 ( \9520 , \9519 );
and \U$702 ( \9521 , \9520 , \9473 );
buf \U$703 ( \9522 , RIe0f3878_4787);
buf \U$704 ( \9523 , \9522 );
and \U$705 ( \9524 , \9001 , \9523 );
nor \U$706 ( \9525 , \9521 , \9524 );
buf \U$707 ( \9526 , RIde5d760_3998);
not \U$708 ( \9527 , \9526 );
not \U$709 ( \9528 , \9527 );
and \U$710 ( \9529 , \9528 , \9139 );
buf \U$711 ( \9530 , RIdfce700_4467);
and \U$712 ( \9531 , \9213 , \9530 );
nor \U$713 ( \9532 , \9529 , \9531 );
buf \U$714 ( \9533 , RIe3f7760_6049);
not \U$715 ( \9534 , \9533 );
or \U$716 ( \9535 , \9534 , \8864 );
buf \U$717 ( \9536 , RIe3887c0_5578);
not \U$718 ( \9537 , \9536 );
not \U$719 ( \9538 , \8916 );
not \U$720 ( \9539 , \9538 );
or \U$721 ( \9540 , \9537 , \9539 );
nand \U$722 ( \9541 , \9535 , \9540 );
buf \U$723 ( \9542 , RIe5e3568_6762);
not \U$724 ( \9543 , \9542 );
or \U$725 ( \9544 , \9543 , \8943 );
buf \U$726 ( \9545 , RIe51acb8_6366);
not \U$727 ( \9546 , \9545 );
or \U$728 ( \9547 , \9546 , \8849 );
nand \U$729 ( \9548 , \9544 , \9547 );
nor \U$730 ( \9549 , \9541 , \9548 );
nand \U$731 ( \9550 , \9525 , \9532 , \9549 );
buf \U$732 ( \9551 , RId7e6f90_1232);
not \U$733 ( \9552 , \9551 );
or \U$734 ( \9553 , \9552 , \9181 );
buf \U$735 ( \9554 , RId71e398_838);
not \U$736 ( \9555 , \9554 );
not \U$737 ( \9556 , \9555 );
not \U$738 ( \9557 , \9556 );
or \U$739 ( \9558 , \9557 , \9316 );
nand \U$740 ( \9559 , \9553 , \9558 );
buf \U$741 ( \9560 , RId8ac078_1630);
not \U$742 ( \9561 , \9560 );
or \U$743 ( \9562 , \9561 , \9234 );
buf \U$744 ( \9563 , RId97ab20_2022);
not \U$745 ( \9564 , \9563 );
or \U$746 ( \9565 , \9564 , \9090 );
nand \U$747 ( \9566 , \9562 , \9565 );
nor \U$748 ( \9567 , \9559 , \9566 );
buf \U$749 ( \9568 , RIdb01d80_2813);
not \U$750 ( \9569 , \9568 );
or \U$751 ( \9570 , \9569 , \8858 );
buf \U$752 ( \9571 , RIda2def0_2418);
not \U$753 ( \9572 , \9571 );
or \U$754 ( \9573 , \9572 , \9495 );
nand \U$755 ( \9574 , \9570 , \9573 );
buf \U$756 ( \9575 , RIdbcc7f0_3208);
not \U$757 ( \9576 , \9575 );
or \U$758 ( \9577 , \9576 , \8841 );
buf \U$759 ( \9578 , RIdd963e0_3603);
not \U$760 ( \9579 , \9578 );
or \U$761 ( \9580 , \9579 , \9022 );
nand \U$762 ( \9581 , \9577 , \9580 );
nor \U$763 ( \9582 , \9574 , \9581 );
nand \U$764 ( \9583 , \9567 , \9582 );
nor \U$765 ( \9584 , \9550 , \9583 );
not \U$766 ( \9585 , RIb7af3d8_259);
xnor \U$767 ( \9586 , \9584 , \9585 );
buf \U$768 ( \9587 , RIe182a68_5243);
not \U$769 ( \9588 , \9587 );
not \U$770 ( \9589 , \9588 );
not \U$771 ( \9590 , \8892 );
and \U$772 ( \9591 , \9589 , \9590 );
buf \U$773 ( \9592 , RIe0f3008_4788);
buf \U$774 ( \9593 , \9592 );
and \U$775 ( \9594 , \9001 , \9593 );
nor \U$776 ( \9595 , \9591 , \9594 );
buf \U$777 ( \9596 , RIde5ad30_4003);
not \U$778 ( \9597 , \9596 );
not \U$779 ( \9598 , \9597 );
and \U$780 ( \9599 , \9598 , \9411 );
buf \U$781 ( \9600 , RIdfc11b8_4469);
and \U$782 ( \9601 , \9466 , \9600 );
nor \U$783 ( \9602 , \9599 , \9601 );
buf \U$784 ( \9603 , RIe3f8a98_6047);
not \U$785 ( \9604 , \9603 );
or \U$786 ( \9605 , \9604 , \8864 );
buf \U$787 ( \9606 , RIe385d90_5583);
not \U$788 ( \9607 , \9606 );
or \U$789 ( \9608 , \9607 , \8918 );
nand \U$790 ( \9609 , \9605 , \9608 );
buf \U$791 ( \9610 , RIe5e09d0_6767);
not \U$792 ( \9611 , \9610 );
or \U$793 ( \9612 , \9611 , \9382 );
buf \U$794 ( \9613 , RIe4af828_6445);
not \U$795 ( \9614 , \9613 );
or \U$796 ( \9615 , \9614 , \9126 );
nand \U$797 ( \9616 , \9612 , \9615 );
nor \U$798 ( \9617 , \9609 , \9616 );
nand \U$799 ( \9618 , \9595 , \9602 , \9617 );
buf \U$800 ( \9619 , RId7e5f28_1234);
not \U$801 ( \9620 , \9619 );
or \U$802 ( \9621 , \9620 , \8956 );
buf \U$803 ( \9622 , RId71bad0_843);
not \U$804 ( \9623 , \9622 );
not \U$805 ( \9624 , \9623 );
not \U$806 ( \9625 , \9624 );
or \U$807 ( \9626 , \9625 , \9316 );
nand \U$808 ( \9627 , \9621 , \9626 );
buf \U$809 ( \9628 , RId8ab538_1631);
not \U$810 ( \9629 , \9628 );
or \U$811 ( \9630 , \9629 , \9234 );
buf \U$812 ( \9631 , RId977f88_2027);
not \U$813 ( \9632 , \9631 );
or \U$814 ( \9633 , \9632 , \9160 );
nand \U$815 ( \9634 , \9630 , \9633 );
nor \U$816 ( \9635 , \9627 , \9634 );
buf \U$817 ( \9636 , RIdaff2d8_2817);
not \U$818 ( \9637 , \9636 );
or \U$819 ( \9638 , \9637 , \9206 );
buf \U$820 ( \9639 , RIda2b970_2422);
not \U$821 ( \9640 , \9639 );
or \U$822 ( \9641 , \9640 , \9495 );
nand \U$823 ( \9642 , \9638 , \9641 );
buf \U$824 ( \9643 , RIdbcac48_3211);
not \U$825 ( \9644 , \9643 );
or \U$826 ( \9645 , \9644 , \8841 );
buf \U$827 ( \9646 , RIdd93500_3608);
not \U$828 ( \9647 , \9646 );
or \U$829 ( \9648 , \9647 , \8937 );
nand \U$830 ( \9649 , \9645 , \9648 );
nor \U$831 ( \9650 , \9642 , \9649 );
nand \U$832 ( \9651 , \9635 , \9650 );
nor \U$833 ( \9652 , \9618 , \9651 );
not \U$834 ( \9653 , RIb7af630_254);
xnor \U$835 ( \9654 , \9652 , \9653 );
buf \U$836 ( \9655 , RIdaffda0_2816);
buf \U$837 ( \9656 , \9655 );
not \U$838 ( \9657 , \9656 );
buf \U$839 ( \9658 , \9657 );
or \U$840 ( \9659 , \9658 , \9206 );
buf \U$841 ( \9660 , RIda2c258_2421);
not \U$842 ( \9661 , \9660 );
or \U$843 ( \9662 , \9661 , \8911 );
nand \U$844 ( \9663 , \9659 , \9662 );
buf \U$845 ( \9664 , RIdb62338_3285);
not \U$846 ( \9665 , \9664 );
or \U$847 ( \9666 , \9665 , \8841 );
buf \U$848 ( \9667 , RIdd93ed8_3607);
not \U$849 ( \9668 , \9667 );
or \U$850 ( \9669 , \9668 , \9022 );
nand \U$851 ( \9670 , \9666 , \9669 );
nor \U$852 ( \9671 , \9663 , \9670 );
buf \U$853 ( \9672 , RIde5b618_4002);
not \U$854 ( \9673 , \9672 );
or \U$855 ( \9674 , \9673 , \8879 );
buf \U$856 ( \9675 , RIdfc07e0_4470);
not \U$857 ( \9676 , \9675 );
or \U$858 ( \9677 , \9676 , \8887 );
nand \U$859 ( \9678 , \9674 , \9677 );
buf \U$860 ( \9679 , RIe1bcc68_5184);
not \U$861 ( \9680 , \9679 );
or \U$862 ( \9681 , \8995 , \9680 );
buf \U$863 ( \9682 , RIe088e38_4865);
not \U$864 ( \9683 , \9682 );
or \U$865 ( \9684 , \9683 , \9291 );
nand \U$866 ( \9685 , \9681 , \9684 );
nor \U$867 ( \9686 , \9678 , \9685 );
buf \U$868 ( \9687 , RId978960_2026);
buf \U$869 ( \9688 , \8923 );
nand \U$870 ( \9689 , \9687 , \9688 );
buf \U$871 ( \9690 , RId8ae508_1629);
nand \U$872 ( \9691 , \9690 , \8928 );
buf \U$873 ( \9692 , RId71c2c8_842);
not \U$874 ( \9693 , \9316 );
and \U$875 ( \9694 , \9692 , \9693 );
buf \U$876 ( \9695 , RId7827c0_1310);
not \U$877 ( \9696 , \9036 );
and \U$878 ( \9697 , \9695 , \9696 );
nor \U$879 ( \9698 , \9694 , \9697 );
nand \U$880 ( \9699 , \9689 , \9691 , \9698 );
not \U$881 ( \9700 , \9699 );
buf \U$882 ( \9701 , RIe386678_5582);
not \U$883 ( \9702 , \9538 );
not \U$884 ( \9703 , \9702 );
and \U$885 ( \9704 , \9701 , \9703 );
buf \U$886 ( \9705 , RIe450d88_5972);
buf \U$887 ( \9706 , \9705 );
not \U$888 ( \9707 , \8864 );
and \U$889 ( \9708 , \9706 , \9707 );
nor \U$890 ( \9709 , \9704 , \9708 );
buf \U$891 ( \9710 , RIe519818_6368);
not \U$892 ( \9711 , \9126 );
and \U$893 ( \9712 , \9710 , \9711 );
buf \U$894 ( \9713 , RIe5e1330_6766);
not \U$895 ( \9714 , \9382 );
and \U$896 ( \9715 , \9713 , \9714 );
nor \U$897 ( \9716 , \9712 , \9715 );
and \U$898 ( \9717 , \9700 , \9709 , \9716 );
nand \U$899 ( \9718 , \9671 , \9686 , \9717 );
not \U$900 ( \9719 , RIb7af5b8_255);
xnor \U$901 ( \9720 , \9718 , \9719 );
buf \U$902 ( \9721 , RIdabee68_2890);
not \U$903 ( \9722 , \9721 );
or \U$904 ( \9723 , \9722 , \9206 );
buf \U$905 ( \9724 , RIda2cbb8_2420);
not \U$906 ( \9725 , \9724 );
or \U$907 ( \9726 , \9725 , \9495 );
nand \U$908 ( \9727 , \9723 , \9726 );
buf \U$909 ( \9728 , RIdb8a760_3284);
not \U$910 ( \9729 , \9728 );
or \U$911 ( \9730 , \9729 , \8841 );
buf \U$912 ( \9731 , RIdd95288_3605);
not \U$913 ( \9732 , \9731 );
or \U$914 ( \9733 , \9732 , \8937 );
nand \U$915 ( \9734 , \9730 , \9733 );
nor \U$916 ( \9735 , \9727 , \9734 );
buf \U$917 ( \9736 , RIde5c6f8_4000);
not \U$918 ( \9737 , \9736 );
or \U$919 ( \9738 , \9737 , \9065 );
buf \U$920 ( \9739 , RIe02a8c0_4391);
not \U$921 ( \9740 , \9739 );
not \U$922 ( \9741 , \9466 );
or \U$923 ( \9742 , \9740 , \9741 );
nand \U$924 ( \9743 , \9738 , \9742 );
buf \U$925 ( \9744 , RIe1bdd48_5182);
not \U$926 ( \9745 , \9744 );
or \U$927 ( \9746 , \8995 , \9745 );
buf \U$928 ( \9747 , RIe0aeb60_4864);
not \U$929 ( \9748 , \9747 );
or \U$930 ( \9749 , \9748 , \9291 );
nand \U$931 ( \9750 , \9746 , \9749 );
nor \U$932 ( \9751 , \9743 , \9750 );
buf \U$933 ( \9752 , RId9799c8_2024);
buf \U$934 ( \9753 , \8923 );
nand \U$935 ( \9754 , \9752 , \9753 );
buf \U$936 ( \9755 , RId8aed00_1628);
not \U$937 ( \9756 , \9015 );
buf \U$938 ( \9757 , \9756 );
nand \U$939 ( \9758 , \9755 , \9757 );
buf \U$940 ( \9759 , RId71d330_840);
not \U$941 ( \9760 , \8949 );
not \U$942 ( \9761 , \9760 );
and \U$943 ( \9762 , \9759 , \9761 );
buf \U$944 ( \9763 , RId790848_1309);
not \U$945 ( \9764 , \9181 );
and \U$946 ( \9765 , \9763 , \9764 );
nor \U$947 ( \9766 , \9762 , \9765 );
nand \U$948 ( \9767 , \9754 , \9758 , \9766 );
not \U$949 ( \9768 , \9767 );
buf \U$950 ( \9769 , RIe3876e0_5580);
not \U$951 ( \9770 , \9539 );
and \U$952 ( \9771 , \9769 , \9770 );
buf \U$953 ( \9772 , RIe3e5628_6050);
not \U$954 ( \9773 , \8982 );
and \U$955 ( \9774 , \9772 , \9773 );
nor \U$956 ( \9775 , \9771 , \9774 );
buf \U$957 ( \9776 , RIe51a2e0_6367);
not \U$958 ( \9777 , \8849 );
and \U$959 ( \9778 , \9776 , \9777 );
buf \U$960 ( \9779 , RIe5e2488_6764);
not \U$961 ( \9780 , \8942 );
not \U$962 ( \9781 , \9780 );
and \U$963 ( \9782 , \9779 , \9781 );
nor \U$964 ( \9783 , \9778 , \9782 );
and \U$965 ( \9784 , \9768 , \9775 , \9783 );
nand \U$966 ( \9785 , \9735 , \9751 , \9784 );
not \U$967 ( \9786 , RIb7af4c8_257);
xnor \U$968 ( \9787 , \9785 , \9786 );
nor \U$969 ( \9788 , \9720 , \9787 );
nand \U$970 ( \9789 , \9586 , \9654 , \9788 );
buf \U$971 ( \9790 , RIe1be5b8_5181);
not \U$972 ( \9791 , \9790 );
not \U$973 ( \9792 , \9791 );
and \U$974 ( \9793 , \9792 , \9473 );
buf \U$975 ( \9794 , RIe0b0870_4861);
and \U$976 ( \9795 , \9001 , \9794 );
nor \U$977 ( \9796 , \9793 , \9795 );
buf \U$978 ( \9797 , RIde5dfd0_3997);
not \U$979 ( \9798 , \9797 );
not \U$980 ( \9799 , \9798 );
and \U$981 ( \9800 , \9799 , \8878 );
buf \U$982 ( \9801 , RIdfcf2b8_4466);
and \U$983 ( \9802 , \8886 , \9801 );
nor \U$984 ( \9803 , \9800 , \9802 );
buf \U$985 ( \9804 , RIe451670_5971);
buf \U$986 ( \9805 , \9804 );
not \U$987 ( \9806 , \9805 );
or \U$988 ( \9807 , \9806 , \9202 );
buf \U$989 ( \9808 , RIe388fb8_5577);
not \U$990 ( \9809 , \9808 );
not \U$991 ( \9810 , \9538 );
or \U$992 ( \9811 , \9809 , \9810 );
nand \U$993 ( \9812 , \9807 , \9811 );
buf \U$994 ( \9813 , RIe588848_6840);
not \U$995 ( \9814 , \9813 );
or \U$996 ( \9815 , \9814 , \8943 );
buf \U$997 ( \9816 , RIe4bd310_6442);
not \U$998 ( \9817 , \9816 );
or \U$999 ( \9818 , \9817 , \9051 );
nand \U$1000 ( \9819 , \9815 , \9818 );
nor \U$1001 ( \9820 , \9812 , \9819 );
nand \U$1002 ( \9821 , \9796 , \9803 , \9820 );
buf \U$1003 ( \9822 , RId7a4bb8_1307);
not \U$1004 ( \9823 , \9822 );
nand \U$1005 ( \9824 , \8833 , \8884 );
or \U$1006 ( \9825 , \9823 , \9824 );
buf \U$1007 ( \9826 , RId71ec08_837);
not \U$1008 ( \9827 , \9826 );
or \U$1009 ( \9828 , \9827 , \8950 );
nand \U$1010 ( \9829 , \9825 , \9828 );
buf \U$1011 ( \9830 , RId86c4d8_1705);
not \U$1012 ( \9831 , \9830 );
or \U$1013 ( \9832 , \9831 , \8929 );
buf \U$1014 ( \9833 , RId97b318_2021);
not \U$1015 ( \9834 , \9833 );
or \U$1016 ( \9835 , \9834 , \9090 );
nand \U$1017 ( \9836 , \9832 , \9835 );
nor \U$1018 ( \9837 , \9829 , \9836 );
buf \U$1019 ( \9838 , RIdb02668_2812);
buf \U$1020 ( \9839 , \9838 );
not \U$1021 ( \9840 , \9839 );
or \U$1022 ( \9841 , \9840 , \9206 );
buf \U$1023 ( \9842 , RIda2e760_2417);
not \U$1024 ( \9843 , \9842 );
not \U$1025 ( \9844 , \8910 );
or \U$1026 ( \9845 , \9843 , \9844 );
nand \U$1027 ( \9846 , \9841 , \9845 );
buf \U$1028 ( \9847 , RIdbcd0d8_3207);
not \U$1029 ( \9848 , \9847 );
or \U$1030 ( \9849 , \9848 , \8841 );
buf \U$1031 ( \9850 , RIdd96cc8_3602);
not \U$1032 ( \9851 , \9850 );
or \U$1033 ( \9852 , \9851 , \9441 );
nand \U$1034 ( \9853 , \9849 , \9852 );
nor \U$1035 ( \9854 , \9846 , \9853 );
nand \U$1036 ( \9855 , \9837 , \9854 );
nor \U$1037 ( \9856 , \9821 , \9855 );
not \U$1038 ( \9857 , RIb7a5bf8_260);
xnor \U$1039 ( \9858 , \9856 , \9857 );
buf \U$1040 ( \9859 , RIe15b900_5260);
not \U$1041 ( \9860 , \9859 );
not \U$1042 ( \9861 , \9860 );
and \U$1043 ( \9862 , \9861 , \9590 );
buf \U$1044 ( \9863 , RIe0f4070_4786);
buf \U$1045 ( \9864 , \9863 );
and \U$1046 ( \9865 , \9001 , \9864 );
nor \U$1047 ( \9866 , \9862 , \9865 );
buf \U$1048 ( \9867 , RIde5e840_3996);
not \U$1049 ( \9868 , \9867 );
not \U$1050 ( \9869 , \9868 );
and \U$1051 ( \9870 , \9869 , \9139 );
buf \U$1052 ( \9871 , RIdfcfc90_4465);
and \U$1053 ( \9872 , \9213 , \9871 );
nor \U$1054 ( \9873 , \9870 , \9872 );
buf \U$1055 ( \9874 , RIe3f9470_6046);
not \U$1056 ( \9875 , \9874 );
or \U$1057 ( \9876 , \9875 , \9202 );
buf \U$1058 ( \9877 , RIe3898a0_5576);
not \U$1059 ( \9878 , \9877 );
or \U$1060 ( \9879 , \9878 , \8918 );
nand \U$1061 ( \9880 , \9876 , \9879 );
buf \U$1062 ( \9881 , RIe5e3e50_6761);
not \U$1063 ( \9882 , \9881 );
not \U$1064 ( \9883 , \9882 );
not \U$1065 ( \9884 , \9883 );
or \U$1066 ( \9885 , \9884 , \9311 );
buf \U$1067 ( \9886 , RIe4b0a70_6443);
not \U$1068 ( \9887 , \9886 );
or \U$1069 ( \9888 , \9887 , \8973 );
nand \U$1070 ( \9889 , \9885 , \9888 );
nor \U$1071 ( \9890 , \9880 , \9889 );
nand \U$1072 ( \9891 , \9866 , \9873 , \9890 );
buf \U$1073 ( \9892 , RId7e7800_1231);
not \U$1074 ( \9893 , \9892 );
not \U$1075 ( \9894 , \9893 );
not \U$1076 ( \9895 , \9894 );
or \U$1077 ( \9896 , \9895 , \9181 );
buf \U$1078 ( \9897 , RId71f400_836);
not \U$1079 ( \9898 , \9897 );
or \U$1080 ( \9899 , \9898 , \9109 );
nand \U$1081 ( \9900 , \9896 , \9899 );
buf \U$1082 ( \9901 , RId8b0290_1626);
buf \U$1083 ( \9902 , \9901 );
not \U$1084 ( \9903 , \9902 );
or \U$1085 ( \9904 , \9903 , \9015 );
buf \U$1086 ( \9905 , RId97bc00_2020);
not \U$1087 ( \9906 , \9905 );
or \U$1088 ( \9907 , \9906 , \8924 );
nand \U$1089 ( \9908 , \9904 , \9907 );
nor \U$1090 ( \9909 , \9900 , \9908 );
buf \U$1091 ( \9910 , RIdb02f50_2811);
not \U$1092 ( \9911 , \9910 );
or \U$1093 ( \9912 , \9911 , \9206 );
buf \U$1094 ( \9913 , RIda2f0c0_2416);
not \U$1095 ( \9914 , \9913 );
or \U$1096 ( \9915 , \9914 , \8911 );
nand \U$1097 ( \9916 , \9912 , \9915 );
buf \U$1098 ( \9917 , RIdbcd9c0_3206);
not \U$1099 ( \9918 , \9917 );
or \U$1100 ( \9919 , \9918 , \8841 );
buf \U$1101 ( \9920 , RIdd97538_3601);
not \U$1102 ( \9921 , \9920 );
or \U$1103 ( \9922 , \9921 , \9099 );
nand \U$1104 ( \9923 , \9919 , \9922 );
nor \U$1105 ( \9924 , \9916 , \9923 );
nand \U$1106 ( \9925 , \9909 , \9924 );
nor \U$1107 ( \9926 , \9891 , \9925 );
not \U$1108 ( \9927 , RIb7a0c48_261);
xnor \U$1109 ( \9928 , \9926 , \9927 );
buf \U$1110 ( \9929 , RIe3f9e48_6045);
not \U$1111 ( \9930 , \9929 );
or \U$1112 ( \9931 , \9930 , \9059 );
buf \U$1113 ( \9932 , RIe387ed8_5579);
not \U$1114 ( \9933 , \9932 );
or \U$1115 ( \9934 , \9933 , \8918 );
nand \U$1116 ( \9935 , \9931 , \9934 );
buf \U$1117 ( \9936 , RIe5e2d70_6763);
not \U$1118 ( \9937 , \9936 );
or \U$1119 ( \9938 , \9937 , \8943 );
buf \U$1120 ( \9939 , RIe4bdce8_6441);
not \U$1121 ( \9940 , \9939 );
or \U$1122 ( \9941 , \9940 , \9126 );
nand \U$1123 ( \9942 , \9938 , \9941 );
nor \U$1124 ( \9943 , \9935 , \9942 );
buf \U$1125 ( \9944 , RIde5cf68_3999);
not \U$1126 ( \9945 , \9944 );
or \U$1127 ( \9946 , \9945 , \9140 );
buf \U$1128 ( \9947 , RIdfcdc38_4468);
not \U$1129 ( \9948 , \9947 );
or \U$1130 ( \9949 , \9948 , \9741 );
nand \U$1131 ( \9950 , \9946 , \9949 );
buf \U$1132 ( \9951 , RIe183440_5242);
not \U$1133 ( \9952 , \9951 );
or \U$1134 ( \9953 , \8892 , \9952 );
buf \U$1135 ( \9954 , RIe0aff10_4862);
not \U$1136 ( \9955 , \9954 );
or \U$1137 ( \9956 , \9955 , \9423 );
nand \U$1138 ( \9957 , \9953 , \9956 );
nor \U$1139 ( \9958 , \9950 , \9957 );
buf \U$1140 ( \9959 , RId97a238_2023);
buf \U$1141 ( \9960 , \8923 );
nand \U$1142 ( \9961 , \9959 , \9960 );
buf \U$1143 ( \9962 , RId8af7c8_1627);
buf \U$1144 ( \9963 , \9756 );
nand \U$1145 ( \9964 , \9962 , \9963 );
buf \U$1146 ( \9965 , RId71dba0_839);
not \U$1147 ( \9966 , \9031 );
and \U$1148 ( \9967 , \9965 , \9966 );
buf \U$1149 ( \9968 , RId7a41e0_1308);
not \U$1150 ( \9969 , \9035 );
not \U$1151 ( \9970 , \9969 );
and \U$1152 ( \9971 , \9968 , \9970 );
nor \U$1153 ( \9972 , \9967 , \9971 );
nand \U$1154 ( \9973 , \9961 , \9964 , \9972 );
not \U$1155 ( \9974 , \9973 );
buf \U$1156 ( \9975 , RIda2d4a0_2419);
and \U$1157 ( \9976 , \8913 , \9975 );
buf \U$1158 ( \9977 , RIdb01498_2814);
buf \U$1159 ( \9978 , \8857 );
and \U$1160 ( \9979 , \9977 , \9978 );
nor \U$1161 ( \9980 , \9976 , \9979 );
buf \U$1162 ( \9981 , \8840 );
buf \U$1163 ( \9982 , RIdbcbe18_3209);
and \U$1164 ( \9983 , \9981 , \9982 );
buf \U$1165 ( \9984 , RIdd95b70_3604);
buf \U$1166 ( \9985 , \8936 );
and \U$1167 ( \9986 , \9984 , \9985 );
nor \U$1168 ( \9987 , \9983 , \9986 );
and \U$1169 ( \9988 , \9974 , \9980 , \9987 );
nand \U$1170 ( \9989 , \9943 , \9958 , \9988 );
not \U$1171 ( \9990 , RIb7af450_258);
xnor \U$1172 ( \9991 , \9989 , \9990 );
buf \U$1173 ( \9992 , RIde5be10_4001);
not \U$1174 ( \9993 , \9992 );
not \U$1175 ( \9994 , \9139 );
or \U$1176 ( \9995 , \9993 , \9994 );
buf \U$1177 ( \9996 , RIe02a050_4392);
not \U$1178 ( \9997 , \9996 );
not \U$1179 ( \9998 , \9466 );
or \U$1180 ( \9999 , \9997 , \9998 );
nand \U$1181 ( \10000 , \9995 , \9999 );
buf \U$1182 ( \10001 , RIe1bd4d8_5183);
not \U$1183 ( \10002 , \10001 );
or \U$1184 ( \10003 , \9285 , \10002 );
buf \U$1185 ( \10004 , RIe0af538_4863);
not \U$1186 ( \10005 , \10004 );
or \U$1187 ( \10006 , \10005 , \9291 );
nand \U$1188 ( \10007 , \10003 , \10006 );
nor \U$1189 ( \10008 , \10000 , \10007 );
buf \U$1190 ( \10009 , RIe3f8048_6048);
not \U$1191 ( \10010 , \10009 );
or \U$1192 ( \10011 , \10010 , \9059 );
buf \U$1193 ( \10012 , RIe386e70_5581);
not \U$1194 ( \10013 , \10012 );
not \U$1195 ( \10014 , \9538 );
or \U$1196 ( \10015 , \10013 , \10014 );
nand \U$1197 ( \10016 , \10011 , \10015 );
buf \U$1198 ( \10017 , RIe5e1ba0_6765);
not \U$1199 ( \10018 , \10017 );
or \U$1200 ( \10019 , \10018 , \9382 );
buf \U$1201 ( \10020 , RIe4b0200_6444);
not \U$1202 ( \10021 , \10020 );
or \U$1203 ( \10022 , \10021 , \8849 );
nand \U$1204 ( \10023 , \10019 , \10022 );
nor \U$1205 ( \10024 , \10016 , \10023 );
buf \U$1206 ( \10025 , RId9791d0_2025);
nand \U$1207 ( \10026 , \10025 , \9688 );
buf \U$1208 ( \10027 , RId86cf28_1704);
buf \U$1209 ( \10028 , \9756 );
nand \U$1210 ( \10029 , \10027 , \10028 );
buf \U$1211 ( \10030 , RId71cb38_841);
not \U$1212 ( \10031 , \9108 );
not \U$1213 ( \10032 , \10031 );
and \U$1214 ( \10033 , \10030 , \10032 );
buf \U$1215 ( \10034 , RId7e6798_1233);
buf \U$1216 ( \10035 , \10034 );
not \U$1217 ( \10036 , \9969 );
and \U$1218 ( \10037 , \10035 , \10036 );
nor \U$1219 ( \10038 , \10033 , \10037 );
nand \U$1220 ( \10039 , \10026 , \10029 , \10038 );
not \U$1221 ( \10040 , \10039 );
buf \U$1222 ( \10041 , RId9cdfc8_2495);
and \U$1223 ( \10042 , \8913 , \10041 );
buf \U$1224 ( \10043 , RIdb00bb0_2815);
and \U$1225 ( \10044 , \10043 , \9978 );
nor \U$1226 ( \10045 , \10042 , \10044 );
buf \U$1227 ( \10046 , \8840 );
buf \U$1228 ( \10047 , RIdbcb530_3210);
and \U$1229 ( \10048 , \10046 , \10047 );
buf \U$1230 ( \10049 , RIdd94928_3606);
buf \U$1231 ( \10050 , \8936 );
and \U$1232 ( \10051 , \10049 , \10050 );
nor \U$1233 ( \10052 , \10048 , \10051 );
and \U$1234 ( \10053 , \10040 , \10045 , \10052 );
nand \U$1235 ( \10054 , \10008 , \10024 , \10053 );
not \U$1236 ( \10055 , RIb7af540_256);
xnor \U$1237 ( \10056 , \10054 , \10055 );
nor \U$1238 ( \10057 , \9991 , \10056 );
nand \U$1239 ( \10058 , \9858 , \9928 , \10057 );
nor \U$1240 ( \10059 , \9517 , \9789 , \10058 );
nand \U$1241 ( \10060 , \9192 , \9462 , \10059 );
not \U$1242 ( \10061 , \10060 );
not \U$1243 ( \10062 , \9494 );
not \U$1244 ( \10063 , \10062 );
not \U$1245 ( \10064 , RIe548ff0_6844);
not \U$1246 ( \10065 , \10064 );
xor \U$1247 ( \10066 , \8837 , \10065 );
not \U$1248 ( \10067 , \8830 );
not \U$1249 ( \10068 , \10067 );
or \U$1250 ( \10069 , \10066 , \10068 );
not \U$1251 ( \10070 , \10069 );
not \U$1252 ( \10071 , \10070 );
or \U$1253 ( \10072 , \8872 , \10071 );
not \U$1254 ( \10073 , \10072 );
not \U$1255 ( \10074 , \10073 );
or \U$1256 ( \10075 , \10063 , \10074 );
not \U$1257 ( \10076 , \8884 );
or \U$1258 ( \10077 , \8830 , \10076 );
not \U$1259 ( \10078 , \10077 );
not \U$1260 ( \10079 , \10078 );
or \U$1261 ( \10080 , \10066 , \10079 );
not \U$1262 ( \10081 , \10080 );
not \U$1263 ( \10082 , \10081 );
or \U$1264 ( \10083 , \9492 , \10082 );
nand \U$1265 ( \10084 , \10075 , \10083 );
not \U$1266 ( \10085 , \9498 );
not \U$1267 ( \10086 , \10085 );
not \U$1268 ( \10087 , \8830 );
or \U$1269 ( \10088 , \10066 , \10087 );
not \U$1270 ( \10089 , \10088 );
not \U$1271 ( \10090 , \10089 );
or \U$1272 ( \10091 , \8855 , \10090 );
not \U$1273 ( \10092 , \10091 );
not \U$1274 ( \10093 , \10092 );
or \U$1275 ( \10094 , \10086 , \10093 );
not \U$1276 ( \10095 , \8839 );
or \U$1277 ( \10096 , \10067 , \10095 );
not \U$1278 ( \10097 , \10096 );
not \U$1279 ( \10098 , \10097 );
or \U$1280 ( \10099 , \10066 , \10098 );
not \U$1281 ( \10100 , \10099 );
not \U$1282 ( \10101 , \10100 );
or \U$1283 ( \10102 , \9500 , \10101 );
nand \U$1284 ( \10103 , \10094 , \10102 );
nor \U$1285 ( \10104 , \10084 , \10103 );
not \U$1286 ( \10105 , \10066 );
or \U$1287 ( \10106 , \10067 , \10105 );
not \U$1288 ( \10107 , \10106 );
not \U$1289 ( \10108 , \10107 );
or \U$1290 ( \10109 , \8883 , \10108 );
or \U$1291 ( \10110 , \9504 , \10109 );
not \U$1292 ( \10111 , \10070 );
or \U$1293 ( \10112 , \8838 , \10111 );
not \U$1294 ( \10113 , \10112 );
not \U$1295 ( \10114 , \10113 );
or \U$1296 ( \10115 , \9506 , \10114 );
nand \U$1297 ( \10116 , \10110 , \10115 );
not \U$1298 ( \10117 , \10116 );
nand \U$1299 ( \10118 , \10066 , \10097 );
not \U$1300 ( \10119 , \10118 );
not \U$1301 ( \10120 , \9511 );
nand \U$1302 ( \10121 , \10119 , \10120 );
not \U$1303 ( \10122 , \10066 );
or \U$1304 ( \10123 , \8830 , \10122 );
not \U$1305 ( \10124 , \10123 );
not \U$1306 ( \10125 , \10124 );
or \U$1307 ( \10126 , \8855 , \10125 );
not \U$1308 ( \10127 , \10126 );
not \U$1309 ( \10128 , \10127 );
or \U$1310 ( \10129 , \9509 , \10128 );
and \U$1311 ( \10130 , \10117 , \10121 , \10129 );
not \U$1312 ( \10131 , \10107 );
or \U$1313 ( \10132 , \8855 , \10131 );
not \U$1314 ( \10133 , \10132 );
not \U$1315 ( \10134 , \10133 );
or \U$1316 ( \10135 , \9467 , \10134 );
not \U$1317 ( \10136 , \10124 );
or \U$1318 ( \10137 , \8838 , \10136 );
not \U$1319 ( \10138 , \10137 );
not \U$1320 ( \10139 , \10138 );
or \U$1321 ( \10140 , \9463 , \10139 );
not \U$1322 ( \10141 , \10124 );
or \U$1323 ( \10142 , \8872 , \10141 );
not \U$1324 ( \10143 , \10142 );
and \U$1325 ( \10144 , \10143 , \9476 );
nand \U$1326 ( \10145 , \10078 , \10066 );
not \U$1327 ( \10146 , \10145 );
not \U$1328 ( \10147 , \10146 );
not \U$1329 ( \10148 , \10147 );
and \U$1330 ( \10149 , \9472 , \10148 );
nor \U$1331 ( \10150 , \10144 , \10149 );
nand \U$1332 ( \10151 , \10135 , \10140 , \10150 );
not \U$1333 ( \10152 , \9480 );
not \U$1334 ( \10153 , \10070 );
or \U$1335 ( \10154 , \8855 , \10153 );
not \U$1336 ( \10155 , \10154 );
and \U$1337 ( \10156 , \10152 , \10155 );
not \U$1338 ( \10157 , \10156 );
not \U$1339 ( \10158 , \10107 );
or \U$1340 ( \10159 , \8872 , \10158 );
not \U$1341 ( \10160 , \10159 );
not \U$1342 ( \10161 , \10160 );
or \U$1343 ( \10162 , \9482 , \10161 );
not \U$1344 ( \10163 , \9487 );
not \U$1345 ( \10164 , \10089 );
or \U$1346 ( \10165 , \8872 , \10164 );
not \U$1347 ( \10166 , \10165 );
and \U$1348 ( \10167 , \10163 , \10166 );
not \U$1349 ( \10168 , \9485 );
not \U$1350 ( \10169 , \10089 );
or \U$1351 ( \10170 , \8883 , \10169 );
not \U$1352 ( \10171 , \10170 );
and \U$1353 ( \10172 , \10168 , \10171 );
nor \U$1354 ( \10173 , \10167 , \10172 );
nand \U$1355 ( \10174 , \10157 , \10162 , \10173 );
nor \U$1356 ( \10175 , \10151 , \10174 );
nand \U$1357 ( \10176 , \10104 , \10130 , \10175 );
not \U$1358 ( \10177 , \10176 );
not \U$1359 ( \10178 , \9772 );
not \U$1360 ( \10179 , \10109 );
not \U$1361 ( \10180 , \10179 );
or \U$1362 ( \10181 , \10178 , \10180 );
not \U$1363 ( \10182 , \9769 );
not \U$1364 ( \10183 , \10143 );
or \U$1365 ( \10184 , \10182 , \10183 );
nand \U$1366 ( \10185 , \10181 , \10184 );
not \U$1367 ( \10186 , \9776 );
or \U$1368 ( \10187 , \10186 , \10159 );
not \U$1369 ( \10188 , \9779 );
not \U$1370 ( \10189 , \10070 );
or \U$1371 ( \10190 , \8855 , \10189 );
or \U$1372 ( \10191 , \10188 , \10190 );
nand \U$1373 ( \10192 , \10187 , \10191 );
nor \U$1374 ( \10193 , \10185 , \10192 );
not \U$1375 ( \10194 , \9763 );
not \U$1376 ( \10195 , \10092 );
or \U$1377 ( \10196 , \10194 , \10195 );
not \U$1378 ( \10197 , \9759 );
not \U$1379 ( \10198 , \10113 );
or \U$1380 ( \10199 , \10197 , \10198 );
nand \U$1381 ( \10200 , \10196 , \10199 );
not \U$1382 ( \10201 , \10200 );
nand \U$1383 ( \10202 , \9755 , \10100 );
nand \U$1384 ( \10203 , \9752 , \10081 );
and \U$1385 ( \10204 , \10201 , \10202 , \10203 );
not \U$1386 ( \10205 , \10145 );
and \U$1387 ( \10206 , \9744 , \10205 );
not \U$1388 ( \10207 , \10206 );
nand \U$1389 ( \10208 , \10066 , \10097 );
not \U$1390 ( \10209 , \10208 );
and \U$1391 ( \10210 , \9747 , \10209 );
not \U$1392 ( \10211 , \10210 );
not \U$1393 ( \10212 , \10132 );
and \U$1394 ( \10213 , \10212 , \9739 );
and \U$1395 ( \10214 , \9736 , \10138 );
nor \U$1396 ( \10215 , \10213 , \10214 );
and \U$1397 ( \10216 , \10207 , \10211 , \10215 );
not \U$1398 ( \10217 , \10216 );
nand \U$1399 ( \10218 , \9731 , \10127 );
not \U$1400 ( \10219 , \10089 );
or \U$1401 ( \10220 , \8872 , \10219 );
not \U$1402 ( \10221 , \10220 );
and \U$1403 ( \10222 , \9728 , \10221 );
not \U$1404 ( \10223 , \10222 );
not \U$1405 ( \10224 , \10073 );
not \U$1406 ( \10225 , \10224 );
and \U$1407 ( \10226 , \9724 , \10225 );
not \U$1408 ( \10227 , \10089 );
or \U$1409 ( \10228 , \8883 , \10227 );
not \U$1410 ( \10229 , \10228 );
and \U$1411 ( \10230 , \9721 , \10229 );
nor \U$1412 ( \10231 , \10226 , \10230 );
nand \U$1413 ( \10232 , \10218 , \10223 , \10231 );
nor \U$1414 ( \10233 , \10217 , \10232 );
nand \U$1415 ( \10234 , \10193 , \10204 , \10233 );
xnor \U$1416 ( \10235 , RIb7af4c8_257, \10234 );
not \U$1417 ( \10236 , \10109 );
nand \U$1418 ( \10237 , \9705 , \10236 );
nand \U$1419 ( \10238 , \9701 , \10143 );
nand \U$1420 ( \10239 , \10237 , \10238 );
not \U$1421 ( \10240 , \9710 );
not \U$1422 ( \10241 , \10107 );
or \U$1423 ( \10242 , \8872 , \10241 );
or \U$1424 ( \10243 , \10240 , \10242 );
not \U$1425 ( \10244 , \9713 );
or \U$1426 ( \10245 , \10244 , \10154 );
nand \U$1427 ( \10246 , \10243 , \10245 );
nor \U$1428 ( \10247 , \10239 , \10246 );
not \U$1429 ( \10248 , \9695 );
or \U$1430 ( \10249 , \10248 , \10195 );
not \U$1431 ( \10250 , \9692 );
or \U$1432 ( \10251 , \10250 , \10198 );
nand \U$1433 ( \10252 , \10249 , \10251 );
not \U$1434 ( \10253 , \10252 );
nand \U$1435 ( \10254 , \9690 , \10100 );
nand \U$1436 ( \10255 , \9687 , \10081 );
and \U$1437 ( \10256 , \10253 , \10254 , \10255 );
not \U$1438 ( \10257 , \10145 );
and \U$1439 ( \10258 , \9679 , \10257 );
not \U$1440 ( \10259 , \10258 );
nand \U$1441 ( \10260 , \10066 , \10097 );
not \U$1442 ( \10261 , \10260 );
and \U$1443 ( \10262 , \9682 , \10261 );
not \U$1444 ( \10263 , \10262 );
and \U$1445 ( \10264 , \10133 , \9675 );
and \U$1446 ( \10265 , \9672 , \10138 );
nor \U$1447 ( \10266 , \10264 , \10265 );
and \U$1448 ( \10267 , \10259 , \10263 , \10266 );
not \U$1449 ( \10268 , \10267 );
nand \U$1450 ( \10269 , \9667 , \10127 );
not \U$1451 ( \10270 , \10089 );
or \U$1452 ( \10271 , \8872 , \10270 );
not \U$1453 ( \10272 , \10271 );
and \U$1454 ( \10273 , \9664 , \10272 );
not \U$1455 ( \10274 , \10273 );
not \U$1456 ( \10275 , \10073 );
not \U$1457 ( \10276 , \10275 );
and \U$1458 ( \10277 , \9660 , \10276 );
not \U$1459 ( \10278 , \10089 );
or \U$1460 ( \10279 , \8883 , \10278 );
not \U$1461 ( \10280 , \10279 );
and \U$1462 ( \10281 , \9656 , \10280 );
nor \U$1463 ( \10282 , \10277 , \10281 );
nand \U$1464 ( \10283 , \10269 , \10274 , \10282 );
nor \U$1465 ( \10284 , \10268 , \10283 );
nand \U$1466 ( \10285 , \10247 , \10256 , \10284 );
xnor \U$1467 ( \10286 , RIb7af5b8_255, \10285 );
not \U$1468 ( \10287 , \10165 );
and \U$1469 ( \10288 , \9196 , \10287 );
not \U$1470 ( \10289 , \10288 );
not \U$1471 ( \10290 , \10126 );
nand \U$1472 ( \10291 , \9239 , \10290 );
not \U$1473 ( \10292 , \10170 );
and \U$1474 ( \10293 , \9204 , \10292 );
not \U$1475 ( \10294 , \10224 );
and \U$1476 ( \10295 , \9225 , \10294 );
nor \U$1477 ( \10296 , \10293 , \10295 );
nand \U$1478 ( \10297 , \10289 , \10291 , \10296 );
not \U$1479 ( \10298 , \10097 );
or \U$1480 ( \10299 , \10066 , \10298 );
not \U$1481 ( \10300 , \10299 );
and \U$1482 ( \10301 , \9233 , \10300 );
not \U$1483 ( \10302 , \10301 );
nand \U$1484 ( \10303 , \9230 , \10081 );
not \U$1485 ( \10304 , \10114 );
and \U$1486 ( \10305 , \9247 , \10304 );
not \U$1487 ( \10306 , \10093 );
and \U$1488 ( \10307 , \9251 , \10306 );
nor \U$1489 ( \10308 , \10305 , \10307 );
nand \U$1490 ( \10309 , \10302 , \10303 , \10308 );
nor \U$1491 ( \10310 , \10297 , \10309 );
not \U$1492 ( \10311 , \10147 );
and \U$1493 ( \10312 , \9216 , \10311 );
not \U$1494 ( \10313 , \10312 );
not \U$1495 ( \10314 , \10118 );
and \U$1496 ( \10315 , \9219 , \10314 );
not \U$1497 ( \10316 , \10315 );
and \U$1498 ( \10317 , \10212 , \9212 );
not \U$1499 ( \10318 , \10137 );
and \U$1500 ( \10319 , \9210 , \10318 );
nor \U$1501 ( \10320 , \10317 , \10319 );
and \U$1502 ( \10321 , \10313 , \10316 , \10320 );
not \U$1503 ( \10322 , \10321 );
not \U$1504 ( \10323 , \9242 );
or \U$1505 ( \10324 , \10323 , \10154 );
not \U$1506 ( \10325 , \10142 );
nand \U$1507 ( \10326 , \9228 , \10325 );
nand \U$1508 ( \10327 , \9200 , \10179 );
nand \U$1509 ( \10328 , \9193 , \10160 );
and \U$1510 ( \10329 , \10324 , \10326 , \10327 , \10328 );
not \U$1511 ( \10330 , \10329 );
nor \U$1512 ( \10331 , \10322 , \10330 );
nand \U$1513 ( \10332 , \10310 , \10331 );
xnor \U$1514 ( \10333 , \10332 , \9260 );
not \U$1515 ( \10334 , \10271 );
and \U$1516 ( \10335 , \8966 , \10334 );
not \U$1517 ( \10336 , \10335 );
nand \U$1518 ( \10337 , \9020 , \10127 );
not \U$1519 ( \10338 , \10279 );
and \U$1520 ( \10339 , \8976 , \10338 );
not \U$1521 ( \10340 , \10073 );
not \U$1522 ( \10341 , \10340 );
and \U$1523 ( \10342 , \9006 , \10341 );
nor \U$1524 ( \10343 , \10339 , \10342 );
nand \U$1525 ( \10344 , \10336 , \10337 , \10343 );
not \U$1526 ( \10345 , \10097 );
or \U$1527 ( \10346 , \10066 , \10345 );
not \U$1528 ( \10347 , \10346 );
and \U$1529 ( \10348 , \9014 , \10347 );
not \U$1530 ( \10349 , \10348 );
nand \U$1531 ( \10350 , \9011 , \10081 );
not \U$1532 ( \10351 , \10114 );
and \U$1533 ( \10352 , \9030 , \10351 );
not \U$1534 ( \10353 , \10093 );
and \U$1535 ( \10354 , \9034 , \10353 );
nor \U$1536 ( \10355 , \10352 , \10354 );
nand \U$1537 ( \10356 , \10349 , \10350 , \10355 );
nor \U$1538 ( \10357 , \10344 , \10356 );
not \U$1539 ( \10358 , \10146 );
not \U$1540 ( \10359 , \10358 );
and \U$1541 ( \10360 , \8996 , \10359 );
not \U$1542 ( \10361 , \10360 );
not \U$1543 ( \10362 , \10260 );
and \U$1544 ( \10363 , \8999 , \10362 );
not \U$1545 ( \10364 , \10363 );
and \U$1546 ( \10365 , \10212 , \8990 );
and \U$1547 ( \10366 , \8986 , \10138 );
nor \U$1548 ( \10367 , \10365 , \10366 );
and \U$1549 ( \10368 , \10361 , \10364 , \10367 );
not \U$1550 ( \10369 , \10368 );
not \U$1551 ( \10370 , \9025 );
or \U$1552 ( \10371 , \10370 , \10190 );
nand \U$1553 ( \10372 , \9009 , \10325 );
nand \U$1554 ( \10373 , \8979 , \10179 );
nand \U$1555 ( \10374 , \8970 , \10160 );
and \U$1556 ( \10375 , \10371 , \10372 , \10373 , \10374 );
not \U$1557 ( \10376 , \10375 );
nor \U$1558 ( \10377 , \10369 , \10376 );
nand \U$1559 ( \10378 , \10357 , \10377 );
xnor \U$1560 ( \10379 , \10378 , \9044 );
nor \U$1561 ( \10380 , \10333 , \10379 );
nand \U$1562 ( \10381 , \10235 , \10286 , \10380 );
not \U$1563 ( \10382 , \10381 );
not \U$1564 ( \10383 , \10220 );
and \U$1565 ( \10384 , \9262 , \10383 );
not \U$1566 ( \10385 , \10384 );
nand \U$1567 ( \10386 , \9307 , \10127 );
not \U$1568 ( \10387 , \10228 );
and \U$1569 ( \10388 , \9269 , \10387 );
not \U$1570 ( \10389 , \10340 );
and \U$1571 ( \10390 , \9295 , \10389 );
nor \U$1572 ( \10391 , \10388 , \10390 );
nand \U$1573 ( \10392 , \10385 , \10386 , \10391 );
not \U$1574 ( \10393 , \10099 );
and \U$1575 ( \10394 , \9302 , \10393 );
not \U$1576 ( \10395 , \10394 );
nand \U$1577 ( \10396 , \9299 , \10081 );
not \U$1578 ( \10397 , \10114 );
and \U$1579 ( \10398 , \9315 , \10397 );
not \U$1580 ( \10399 , \10093 );
and \U$1581 ( \10400 , \9319 , \10399 );
nor \U$1582 ( \10401 , \10398 , \10400 );
nand \U$1583 ( \10402 , \10395 , \10396 , \10401 );
nor \U$1584 ( \10403 , \10392 , \10402 );
not \U$1585 ( \10404 , \10145 );
and \U$1586 ( \10405 , \9286 , \10404 );
not \U$1587 ( \10406 , \10405 );
not \U$1588 ( \10407 , \10208 );
and \U$1589 ( \10408 , \9289 , \10407 );
not \U$1590 ( \10409 , \10408 );
and \U$1591 ( \10410 , \10212 , \9281 );
and \U$1592 ( \10411 , \9277 , \10138 );
nor \U$1593 ( \10412 , \10410 , \10411 );
and \U$1594 ( \10413 , \10406 , \10409 , \10412 );
not \U$1595 ( \10414 , \10413 );
not \U$1596 ( \10415 , \9310 );
not \U$1597 ( \10416 , \10070 );
or \U$1598 ( \10417 , \8855 , \10416 );
or \U$1599 ( \10418 , \10415 , \10417 );
nand \U$1600 ( \10419 , \9297 , \10325 );
nand \U$1601 ( \10420 , \9272 , \10236 );
not \U$1602 ( \10421 , \10160 );
or \U$1603 ( \10422 , \9266 , \10421 );
and \U$1604 ( \10423 , \10418 , \10419 , \10420 , \10422 );
not \U$1605 ( \10424 , \10423 );
nor \U$1606 ( \10425 , \10414 , \10424 );
nand \U$1607 ( \10426 , \10403 , \10425 );
xnor \U$1608 ( \10427 , \10426 , \9327 );
not \U$1609 ( \10428 , \10165 );
and \U$1610 ( \10429 , \9394 , \10428 );
not \U$1611 ( \10430 , \10429 );
nand \U$1612 ( \10431 , \9440 , \10127 );
not \U$1613 ( \10432 , \10170 );
and \U$1614 ( \10433 , \9401 , \10432 );
not \U$1615 ( \10434 , \10275 );
and \U$1616 ( \10435 , \9427 , \10434 );
nor \U$1617 ( \10436 , \10433 , \10435 );
nand \U$1618 ( \10437 , \10430 , \10431 , \10436 );
not \U$1619 ( \10438 , \10299 );
and \U$1620 ( \10439 , \9435 , \10438 );
not \U$1621 ( \10440 , \10439 );
nand \U$1622 ( \10441 , \9432 , \10081 );
not \U$1623 ( \10442 , \10114 );
and \U$1624 ( \10443 , \9449 , \10442 );
not \U$1625 ( \10444 , \10093 );
and \U$1626 ( \10445 , \9453 , \10444 );
nor \U$1627 ( \10446 , \10443 , \10445 );
nand \U$1628 ( \10447 , \10440 , \10441 , \10446 );
nor \U$1629 ( \10448 , \10437 , \10447 );
not \U$1630 ( \10449 , \10358 );
and \U$1631 ( \10450 , \9418 , \10449 );
not \U$1632 ( \10451 , \10450 );
not \U$1633 ( \10452 , \10118 );
and \U$1634 ( \10453 , \9421 , \10452 );
not \U$1635 ( \10454 , \10453 );
not \U$1636 ( \10455 , \9409 );
not \U$1637 ( \10456 , \10455 );
and \U$1638 ( \10457 , \10456 , \10138 );
and \U$1639 ( \10458 , \10133 , \9414 );
nor \U$1640 ( \10459 , \10457 , \10458 );
and \U$1641 ( \10460 , \10451 , \10454 , \10459 );
not \U$1642 ( \10461 , \10460 );
not \U$1643 ( \10462 , \9444 );
or \U$1644 ( \10463 , \10462 , \10154 );
not \U$1645 ( \10464 , \9430 );
not \U$1646 ( \10465 , \10143 );
or \U$1647 ( \10466 , \10464 , \10465 );
not \U$1648 ( \10467 , \10236 );
or \U$1649 ( \10468 , \9405 , \10467 );
not \U$1650 ( \10469 , \10160 );
or \U$1651 ( \10470 , \9398 , \10469 );
and \U$1652 ( \10471 , \10463 , \10466 , \10468 , \10470 );
not \U$1653 ( \10472 , \10471 );
nor \U$1654 ( \10473 , \10461 , \10472 );
nand \U$1655 ( \10474 , \10448 , \10473 );
xnor \U$1656 ( \10475 , \10474 , \9460 );
nor \U$1657 ( \10476 , \10427 , \10475 );
nand \U$1658 ( \10477 , \9646 , \10290 );
not \U$1659 ( \10478 , \10271 );
and \U$1660 ( \10479 , \9643 , \10478 );
not \U$1661 ( \10480 , \10479 );
not \U$1662 ( \10481 , \10340 );
and \U$1663 ( \10482 , \9639 , \10481 );
not \U$1664 ( \10483 , \10279 );
and \U$1665 ( \10484 , \9636 , \10483 );
nor \U$1666 ( \10485 , \10482 , \10484 );
nand \U$1667 ( \10486 , \10477 , \10480 , \10485 );
not \U$1668 ( \10487 , \10080 );
and \U$1669 ( \10488 , \9631 , \10487 );
not \U$1670 ( \10489 , \10488 );
not \U$1671 ( \10490 , \10346 );
and \U$1672 ( \10491 , \9628 , \10490 );
not \U$1673 ( \10492 , \10491 );
not \U$1674 ( \10493 , \10114 );
and \U$1675 ( \10494 , \9622 , \10493 );
not \U$1676 ( \10495 , \10093 );
and \U$1677 ( \10496 , \9619 , \10495 );
nor \U$1678 ( \10497 , \10494 , \10496 );
and \U$1679 ( \10498 , \10489 , \10492 , \10497 );
not \U$1680 ( \10499 , \10498 );
nor \U$1681 ( \10500 , \10486 , \10499 );
not \U$1682 ( \10501 , \10145 );
and \U$1683 ( \10502 , \9587 , \10501 );
not \U$1684 ( \10503 , \10502 );
not \U$1685 ( \10504 , \10260 );
and \U$1686 ( \10505 , \9593 , \10504 );
not \U$1687 ( \10506 , \10505 );
and \U$1688 ( \10507 , \10133 , \9600 );
and \U$1689 ( \10508 , \9596 , \10138 );
nor \U$1690 ( \10509 , \10507 , \10508 );
and \U$1691 ( \10510 , \10503 , \10506 , \10509 );
not \U$1692 ( \10511 , \10510 );
or \U$1693 ( \10512 , \9611 , \10190 );
nand \U$1694 ( \10513 , \9603 , \10179 );
nand \U$1695 ( \10514 , \9606 , \10143 );
nand \U$1696 ( \10515 , \9613 , \10160 );
and \U$1697 ( \10516 , \10512 , \10513 , \10514 , \10515 );
not \U$1698 ( \10517 , \10516 );
nor \U$1699 ( \10518 , \10511 , \10517 );
nand \U$1700 ( \10519 , \10500 , \10518 );
xnor \U$1701 ( \10520 , \10519 , \9653 );
not \U$1702 ( \10521 , \10220 );
and \U$1703 ( \10522 , \9331 , \10521 );
not \U$1704 ( \10523 , \10522 );
nand \U$1705 ( \10524 , \9374 , \10127 );
not \U$1706 ( \10525 , \10228 );
and \U$1707 ( \10526 , \9338 , \10525 );
not \U$1708 ( \10527 , \10074 );
and \U$1709 ( \10528 , \9361 , \10527 );
nor \U$1710 ( \10529 , \10526 , \10528 );
nand \U$1711 ( \10530 , \10523 , \10524 , \10529 );
not \U$1712 ( \10531 , \10099 );
and \U$1713 ( \10532 , \9369 , \10531 );
not \U$1714 ( \10533 , \10532 );
nand \U$1715 ( \10534 , \9366 , \10081 );
not \U$1716 ( \10535 , \10093 );
and \U$1717 ( \10536 , \9377 , \10535 );
not \U$1718 ( \10537 , \10114 );
and \U$1719 ( \10538 , \9385 , \10537 );
nor \U$1720 ( \10539 , \10536 , \10538 );
nand \U$1721 ( \10540 , \10533 , \10534 , \10539 );
nor \U$1722 ( \10541 , \10530 , \10540 );
not \U$1723 ( \10542 , \10145 );
and \U$1724 ( \10543 , \9353 , \10542 );
not \U$1725 ( \10544 , \10543 );
not \U$1726 ( \10545 , \10208 );
and \U$1727 ( \10546 , \9356 , \10545 );
not \U$1728 ( \10547 , \10546 );
and \U$1729 ( \10548 , \10212 , \9348 );
and \U$1730 ( \10549 , \9346 , \10138 );
nor \U$1731 ( \10550 , \10548 , \10549 );
and \U$1732 ( \10551 , \10544 , \10547 , \10550 );
not \U$1733 ( \10552 , \10551 );
not \U$1734 ( \10553 , \9380 );
or \U$1735 ( \10554 , \10553 , \10417 );
nand \U$1736 ( \10555 , \9364 , \10143 );
nand \U$1737 ( \10556 , \9341 , \10236 );
nand \U$1738 ( \10557 , \9334 , \10160 );
and \U$1739 ( \10558 , \10554 , \10555 , \10556 , \10557 );
not \U$1740 ( \10559 , \10558 );
nor \U$1741 ( \10560 , \10552 , \10559 );
nand \U$1742 ( \10561 , \10541 , \10560 );
xnor \U$1743 ( \10562 , \10561 , \9392 );
nor \U$1744 ( \10563 , \10520 , \10562 );
and \U$1745 ( \10564 , \10382 , \10476 , \10563 );
nand \U$1746 ( \10565 , \9920 , \10127 );
not \U$1747 ( \10566 , \10165 );
and \U$1748 ( \10567 , \9917 , \10566 );
not \U$1749 ( \10568 , \10567 );
not \U$1750 ( \10569 , \10340 );
and \U$1751 ( \10570 , \9913 , \10569 );
not \U$1752 ( \10571 , \10170 );
and \U$1753 ( \10572 , \9910 , \10571 );
nor \U$1754 ( \10573 , \10570 , \10572 );
nand \U$1755 ( \10574 , \10565 , \10568 , \10573 );
not \U$1756 ( \10575 , \10080 );
and \U$1757 ( \10576 , \9905 , \10575 );
not \U$1758 ( \10577 , \10576 );
not \U$1759 ( \10578 , \10299 );
and \U$1760 ( \10579 , \9902 , \10578 );
not \U$1761 ( \10580 , \10579 );
not \U$1762 ( \10581 , \10198 );
and \U$1763 ( \10582 , \9897 , \10581 );
not \U$1764 ( \10583 , \10195 );
and \U$1765 ( \10584 , \9892 , \10583 );
nor \U$1766 ( \10585 , \10582 , \10584 );
and \U$1767 ( \10586 , \10577 , \10580 , \10585 );
not \U$1768 ( \10587 , \10586 );
nor \U$1769 ( \10588 , \10574 , \10587 );
not \U$1770 ( \10589 , \10145 );
and \U$1771 ( \10590 , \9859 , \10589 );
not \U$1772 ( \10591 , \10590 );
not \U$1773 ( \10592 , \10208 );
and \U$1774 ( \10593 , \9864 , \10592 );
not \U$1775 ( \10594 , \10593 );
and \U$1776 ( \10595 , \10133 , \9871 );
and \U$1777 ( \10596 , \9867 , \10138 );
nor \U$1778 ( \10597 , \10595 , \10596 );
and \U$1779 ( \10598 , \10591 , \10594 , \10597 );
not \U$1780 ( \10599 , \10598 );
or \U$1781 ( \10600 , \9884 , \10417 );
nand \U$1782 ( \10601 , \9874 , \10179 );
nand \U$1783 ( \10602 , \9877 , \10143 );
nand \U$1784 ( \10603 , \9886 , \10160 );
and \U$1785 ( \10604 , \10600 , \10601 , \10602 , \10603 );
not \U$1786 ( \10605 , \10604 );
nor \U$1787 ( \10606 , \10599 , \10605 );
nand \U$1788 ( \10607 , \10588 , \10606 );
xnor \U$1789 ( \10608 , RIb7a0c48_261, \10607 );
nand \U$1790 ( \10609 , \9996 , \10133 );
nand \U$1791 ( \10610 , \9992 , \10138 );
nand \U$1792 ( \10611 , \10609 , \10610 );
not \U$1793 ( \10612 , \10611 );
nand \U$1794 ( \10613 , \10119 , \10004 );
nand \U$1795 ( \10614 , \10001 , \10146 );
and \U$1796 ( \10615 , \10612 , \10613 , \10614 );
nand \U$1797 ( \10616 , \10009 , \10236 );
nand \U$1798 ( \10617 , \10012 , \10143 );
nand \U$1799 ( \10618 , \10616 , \10617 );
not \U$1800 ( \10619 , \10020 );
not \U$1801 ( \10620 , \10107 );
or \U$1802 ( \10621 , \8872 , \10620 );
or \U$1803 ( \10622 , \10619 , \10621 );
or \U$1804 ( \10623 , \10018 , \10417 );
nand \U$1805 ( \10624 , \10622 , \10623 );
nor \U$1806 ( \10625 , \10618 , \10624 );
nand \U$1807 ( \10626 , \10049 , \10127 );
not \U$1808 ( \10627 , \10220 );
and \U$1809 ( \10628 , \10047 , \10627 );
not \U$1810 ( \10629 , \10628 );
not \U$1811 ( \10630 , \10224 );
and \U$1812 ( \10631 , \10041 , \10630 );
not \U$1813 ( \10632 , \10228 );
and \U$1814 ( \10633 , \10043 , \10632 );
nor \U$1815 ( \10634 , \10631 , \10633 );
nand \U$1816 ( \10635 , \10626 , \10629 , \10634 );
not \U$1817 ( \10636 , \10080 );
and \U$1818 ( \10637 , \10025 , \10636 );
not \U$1819 ( \10638 , \10637 );
not \U$1820 ( \10639 , \10099 );
and \U$1821 ( \10640 , \10027 , \10639 );
not \U$1822 ( \10641 , \10640 );
not \U$1823 ( \10642 , \10198 );
and \U$1824 ( \10643 , \10030 , \10642 );
not \U$1825 ( \10644 , \10195 );
and \U$1826 ( \10645 , \10035 , \10644 );
nor \U$1827 ( \10646 , \10643 , \10645 );
and \U$1828 ( \10647 , \10638 , \10641 , \10646 );
not \U$1829 ( \10648 , \10647 );
nor \U$1830 ( \10649 , \10635 , \10648 );
nand \U$1831 ( \10650 , \10615 , \10625 , \10649 );
xnor \U$1832 ( \10651 , RIb7af540_256, \10650 );
nand \U$1833 ( \10652 , \9578 , \10290 );
not \U$1834 ( \10653 , \10165 );
and \U$1835 ( \10654 , \9575 , \10653 );
not \U$1836 ( \10655 , \10654 );
not \U$1837 ( \10656 , \10275 );
and \U$1838 ( \10657 , \9571 , \10656 );
not \U$1839 ( \10658 , \10170 );
and \U$1840 ( \10659 , \9568 , \10658 );
nor \U$1841 ( \10660 , \10657 , \10659 );
nand \U$1842 ( \10661 , \10652 , \10655 , \10660 );
not \U$1843 ( \10662 , \10080 );
and \U$1844 ( \10663 , \9563 , \10662 );
not \U$1845 ( \10664 , \10663 );
not \U$1846 ( \10665 , \10299 );
and \U$1847 ( \10666 , \9560 , \10665 );
not \U$1848 ( \10667 , \10666 );
not \U$1849 ( \10668 , \10114 );
and \U$1850 ( \10669 , \9554 , \10668 );
not \U$1851 ( \10670 , \10093 );
and \U$1852 ( \10671 , \9551 , \10670 );
nor \U$1853 ( \10672 , \10669 , \10671 );
and \U$1854 ( \10673 , \10664 , \10667 , \10672 );
not \U$1855 ( \10674 , \10673 );
nor \U$1856 ( \10675 , \10661 , \10674 );
not \U$1857 ( \10676 , \10358 );
and \U$1858 ( \10677 , \9518 , \10676 );
not \U$1859 ( \10678 , \10677 );
not \U$1860 ( \10679 , \10118 );
and \U$1861 ( \10680 , \9523 , \10679 );
not \U$1862 ( \10681 , \10680 );
and \U$1863 ( \10682 , \10133 , \9530 );
and \U$1864 ( \10683 , \9526 , \10138 );
nor \U$1865 ( \10684 , \10682 , \10683 );
and \U$1866 ( \10685 , \10678 , \10681 , \10684 );
not \U$1867 ( \10686 , \10685 );
or \U$1868 ( \10687 , \9543 , \10154 );
nand \U$1869 ( \10688 , \9533 , \10179 );
nand \U$1870 ( \10689 , \9536 , \10325 );
nand \U$1871 ( \10690 , \9545 , \10160 );
and \U$1872 ( \10691 , \10687 , \10688 , \10689 , \10690 );
not \U$1873 ( \10692 , \10691 );
nor \U$1874 ( \10693 , \10686 , \10692 );
nand \U$1875 ( \10694 , \10675 , \10693 );
xnor \U$1876 ( \10695 , \10694 , \9585 );
nand \U$1877 ( \10696 , \9984 , \10290 );
not \U$1878 ( \10697 , \10271 );
and \U$1879 ( \10698 , \9982 , \10697 );
not \U$1880 ( \10699 , \10698 );
not \U$1881 ( \10700 , \10275 );
and \U$1882 ( \10701 , \9975 , \10700 );
not \U$1883 ( \10702 , \10279 );
and \U$1884 ( \10703 , \9977 , \10702 );
nor \U$1885 ( \10704 , \10701 , \10703 );
nand \U$1886 ( \10705 , \10696 , \10699 , \10704 );
not \U$1887 ( \10706 , \10080 );
and \U$1888 ( \10707 , \9959 , \10706 );
not \U$1889 ( \10708 , \10707 );
buf \U$1890 ( \10709 , \9962 );
not \U$1891 ( \10710 , \10346 );
and \U$1892 ( \10711 , \10709 , \10710 );
not \U$1893 ( \10712 , \10711 );
not \U$1894 ( \10713 , \10198 );
and \U$1895 ( \10714 , \9965 , \10713 );
not \U$1896 ( \10715 , \10195 );
and \U$1897 ( \10716 , \9968 , \10715 );
nor \U$1898 ( \10717 , \10714 , \10716 );
and \U$1899 ( \10718 , \10708 , \10712 , \10717 );
not \U$1900 ( \10719 , \10718 );
nor \U$1901 ( \10720 , \10705 , \10719 );
not \U$1902 ( \10721 , \10145 );
and \U$1903 ( \10722 , \9951 , \10721 );
not \U$1904 ( \10723 , \10722 );
not \U$1905 ( \10724 , \10260 );
and \U$1906 ( \10725 , \9954 , \10724 );
not \U$1907 ( \10726 , \10725 );
and \U$1908 ( \10727 , \10133 , \9947 );
and \U$1909 ( \10728 , \9944 , \10138 );
nor \U$1910 ( \10729 , \10727 , \10728 );
and \U$1911 ( \10730 , \10723 , \10726 , \10729 );
not \U$1912 ( \10731 , \10730 );
or \U$1913 ( \10732 , \9937 , \10190 );
nand \U$1914 ( \10733 , \9929 , \10179 );
nand \U$1915 ( \10734 , \9932 , \10143 );
nand \U$1916 ( \10735 , \9939 , \10160 );
and \U$1917 ( \10736 , \10732 , \10733 , \10734 , \10735 );
not \U$1918 ( \10737 , \10736 );
nor \U$1919 ( \10738 , \10731 , \10737 );
nand \U$1920 ( \10739 , \10720 , \10738 );
xnor \U$1921 ( \10740 , \10739 , \9990 );
nor \U$1922 ( \10741 , \10695 , \10740 );
nand \U$1923 ( \10742 , \10608 , \10651 , \10741 );
not \U$1924 ( \10743 , \10220 );
and \U$1925 ( \10744 , \8827 , \10743 );
not \U$1926 ( \10745 , \10744 );
nand \U$1927 ( \10746 , \8934 , \10127 );
not \U$1928 ( \10747 , \10228 );
and \U$1929 ( \10748 , \8852 , \10747 );
not \U$1930 ( \10749 , \10340 );
and \U$1931 ( \10750 , \8904 , \10749 );
nor \U$1932 ( \10751 , \10748 , \10750 );
nand \U$1933 ( \10752 , \10745 , \10746 , \10751 );
not \U$1934 ( \10753 , \10099 );
and \U$1935 ( \10754 , \8927 , \10753 );
not \U$1936 ( \10755 , \10754 );
nand \U$1937 ( \10756 , \8921 , \10081 );
not \U$1938 ( \10757 , \10198 );
and \U$1939 ( \10758 , \8947 , \10757 );
not \U$1940 ( \10759 , \10093 );
and \U$1941 ( \10760 , \8953 , \10759 );
nor \U$1942 ( \10761 , \10758 , \10760 );
nand \U$1943 ( \10762 , \10755 , \10756 , \10761 );
nor \U$1944 ( \10763 , \10752 , \10762 );
not \U$1945 ( \10764 , \10358 );
and \U$1946 ( \10765 , \8893 , \10764 );
not \U$1947 ( \10766 , \10765 );
not \U$1948 ( \10767 , \10118 );
and \U$1949 ( \10768 , \8896 , \10767 );
not \U$1950 ( \10769 , \10768 );
and \U$1951 ( \10770 , \10133 , \8881 );
and \U$1952 ( \10771 , \8868 , \10138 );
nor \U$1953 ( \10772 , \10770 , \10771 );
and \U$1954 ( \10773 , \10766 , \10769 , \10772 );
not \U$1955 ( \10774 , \10773 );
not \U$1956 ( \10775 , \8940 );
or \U$1957 ( \10776 , \10775 , \10154 );
nand \U$1958 ( \10777 , \8915 , \10143 );
nand \U$1959 ( \10778 , \8860 , \10236 );
nand \U$1960 ( \10779 , \8843 , \10160 );
and \U$1961 ( \10780 , \10776 , \10777 , \10778 , \10779 );
not \U$1962 ( \10781 , \10780 );
nor \U$1963 ( \10782 , \10774 , \10781 );
nand \U$1964 ( \10783 , \10763 , \10782 );
xnor \U$1965 ( \10784 , RIb7b93b0_251, \10783 );
nand \U$1966 ( \10785 , \9801 , \10133 );
nand \U$1967 ( \10786 , \9797 , \10138 );
nand \U$1968 ( \10787 , \10785 , \10786 );
not \U$1969 ( \10788 , \10787 );
nand \U$1970 ( \10789 , \10119 , \9794 );
nand \U$1971 ( \10790 , \9790 , \10146 );
and \U$1972 ( \10791 , \10788 , \10789 , \10790 );
nand \U$1973 ( \10792 , \9804 , \10236 );
nand \U$1974 ( \10793 , \9808 , \10143 );
nand \U$1975 ( \10794 , \10792 , \10793 );
not \U$1976 ( \10795 , \9816 );
or \U$1977 ( \10796 , \10795 , \10242 );
or \U$1978 ( \10797 , \9814 , \10154 );
nand \U$1979 ( \10798 , \10796 , \10797 );
nor \U$1980 ( \10799 , \10794 , \10798 );
nand \U$1981 ( \10800 , \9850 , \10127 );
not \U$1982 ( \10801 , \10271 );
and \U$1983 ( \10802 , \9847 , \10801 );
not \U$1984 ( \10803 , \10802 );
not \U$1985 ( \10804 , \10074 );
and \U$1986 ( \10805 , \9842 , \10804 );
not \U$1987 ( \10806 , \10279 );
and \U$1988 ( \10807 , \9839 , \10806 );
nor \U$1989 ( \10808 , \10805 , \10807 );
nand \U$1990 ( \10809 , \10800 , \10803 , \10808 );
not \U$1991 ( \10810 , \10080 );
and \U$1992 ( \10811 , \9833 , \10810 );
not \U$1993 ( \10812 , \10811 );
not \U$1994 ( \10813 , \10346 );
and \U$1995 ( \10814 , \9830 , \10813 );
not \U$1996 ( \10815 , \10814 );
not \U$1997 ( \10816 , \10198 );
and \U$1998 ( \10817 , \9826 , \10816 );
not \U$1999 ( \10818 , \10195 );
and \U$2000 ( \10819 , \9822 , \10818 );
nor \U$2001 ( \10820 , \10817 , \10819 );
and \U$2002 ( \10821 , \10812 , \10815 , \10820 );
not \U$2003 ( \10822 , \10821 );
nor \U$2004 ( \10823 , \10809 , \10822 );
nand \U$2005 ( \10824 , \10791 , \10799 , \10823 );
xnor \U$2006 ( \10825 , RIb7a5bf8_260, \10824 );
not \U$2007 ( \10826 , \10165 );
and \U$2008 ( \10827 , \9046 , \10826 );
not \U$2009 ( \10828 , \10827 );
nand \U$2010 ( \10829 , \9098 , \10127 );
not \U$2011 ( \10830 , \10170 );
and \U$2012 ( \10831 , \9054 , \10830 );
not \U$2013 ( \10832 , \10224 );
and \U$2014 ( \10833 , \9081 , \10832 );
nor \U$2015 ( \10834 , \10831 , \10833 );
nand \U$2016 ( \10835 , \10828 , \10829 , \10834 );
not \U$2017 ( \10836 , \10299 );
and \U$2018 ( \10837 , \9093 , \10836 );
not \U$2019 ( \10838 , \10837 );
nand \U$2020 ( \10839 , \9089 , \10081 );
not \U$2021 ( \10840 , \10114 );
and \U$2022 ( \10841 , \9107 , \10840 );
not \U$2023 ( \10842 , \10092 );
not \U$2024 ( \10843 , \10842 );
and \U$2025 ( \10844 , \9112 , \10843 );
nor \U$2026 ( \10845 , \10841 , \10844 );
nand \U$2027 ( \10846 , \10838 , \10839 , \10845 );
nor \U$2028 ( \10847 , \10835 , \10846 );
not \U$2029 ( \10848 , \10145 );
and \U$2030 ( \10849 , \9072 , \10848 );
not \U$2031 ( \10850 , \10849 );
not \U$2032 ( \10851 , \10260 );
and \U$2033 ( \10852 , \9075 , \10851 );
not \U$2034 ( \10853 , \10852 );
and \U$2035 ( \10854 , \10212 , \9067 );
and \U$2036 ( \10855 , \9063 , \10138 );
nor \U$2037 ( \10856 , \10854 , \10855 );
and \U$2038 ( \10857 , \10850 , \10853 , \10856 );
not \U$2039 ( \10858 , \10857 );
not \U$2040 ( \10859 , \9102 );
or \U$2041 ( \10860 , \10859 , \10190 );
nand \U$2042 ( \10861 , \9085 , \10325 );
nand \U$2043 ( \10862 , \9057 , \10236 );
nand \U$2044 ( \10863 , \9049 , \10160 );
and \U$2045 ( \10864 , \10860 , \10861 , \10862 , \10863 );
not \U$2046 ( \10865 , \10864 );
nor \U$2047 ( \10866 , \10858 , \10865 );
nand \U$2048 ( \10867 , \10847 , \10866 );
xnor \U$2049 ( \10868 , \10867 , \9119 );
not \U$2050 ( \10869 , \10271 );
and \U$2051 ( \10870 , \9121 , \10869 );
not \U$2052 ( \10871 , \10870 );
nand \U$2053 ( \10872 , \9168 , \10127 );
not \U$2054 ( \10873 , \10279 );
and \U$2055 ( \10874 , \9129 , \10873 );
not \U$2056 ( \10875 , \10275 );
and \U$2057 ( \10876 , \9155 , \10875 );
nor \U$2058 ( \10877 , \10874 , \10876 );
nand \U$2059 ( \10878 , \10871 , \10872 , \10877 );
not \U$2060 ( \10879 , \10346 );
and \U$2061 ( \10880 , \9163 , \10879 );
not \U$2062 ( \10881 , \10880 );
nand \U$2063 ( \10882 , \9159 , \10081 );
not \U$2064 ( \10883 , \10114 );
and \U$2065 ( \10884 , \9176 , \10883 );
not \U$2066 ( \10885 , \10842 );
and \U$2067 ( \10886 , \9180 , \10885 );
nor \U$2068 ( \10887 , \10884 , \10886 );
nand \U$2069 ( \10888 , \10881 , \10882 , \10887 );
nor \U$2070 ( \10889 , \10878 , \10888 );
not \U$2071 ( \10890 , \10147 );
and \U$2072 ( \10891 , \9147 , \10890 );
not \U$2073 ( \10892 , \10891 );
not \U$2074 ( \10893 , \10208 );
and \U$2075 ( \10894 , \9150 , \10893 );
not \U$2076 ( \10895 , \10894 );
and \U$2077 ( \10896 , \10133 , \9142 );
and \U$2078 ( \10897 , \9137 , \10138 );
nor \U$2079 ( \10898 , \10896 , \10897 );
and \U$2080 ( \10899 , \10892 , \10895 , \10898 );
not \U$2081 ( \10900 , \10899 );
not \U$2082 ( \10901 , \9172 );
or \U$2083 ( \10902 , \10901 , \10417 );
nand \U$2084 ( \10903 , \9157 , \10143 );
nand \U$2085 ( \10904 , \9132 , \10236 );
nand \U$2086 ( \10905 , \9124 , \10160 );
and \U$2087 ( \10906 , \10902 , \10903 , \10904 , \10905 );
not \U$2088 ( \10907 , \10906 );
nor \U$2089 ( \10908 , \10900 , \10907 );
nand \U$2090 ( \10909 , \10889 , \10908 );
xnor \U$2091 ( \10910 , \10909 , \9188 );
nor \U$2092 ( \10911 , \10868 , \10910 );
nand \U$2093 ( \10912 , \10784 , \10825 , \10911 );
nor \U$2094 ( \10913 , \10742 , \10912 );
nand \U$2095 ( \10914 , \10177 , \10564 , \10913 );
not \U$2096 ( \10915 , \10914 );
not \U$2097 ( \10916 , \10915 );
nand \U$2098 ( \10917 , \8905 , \8870 );
xor \U$2099 ( \10918 , \8837 , \10917 );
not \U$2100 ( \10919 , \8834 );
not \U$2101 ( \10920 , \10919 );
not \U$2102 ( \10921 , \10067 );
or \U$2103 ( \10922 , \10919 , \10921 );
nand \U$2104 ( \10923 , \10917 , \10922 );
not \U$2105 ( \10924 , \10923 );
or \U$2106 ( \10925 , \10920 , \10924 );
not \U$2107 ( \10926 , \10925 );
and \U$2108 ( \10927 , \10918 , \10926 );
not \U$2109 ( \10928 , \8836 );
not \U$2110 ( \10929 , \10917 );
or \U$2111 ( \10930 , \10928 , \10929 );
xor \U$2112 ( \10931 , \10065 , \10930 );
not \U$2113 ( \10932 , \10931 );
nand \U$2114 ( \10933 , \10927 , \10932 );
not \U$2115 ( \10934 , \10933 );
not \U$2116 ( \10935 , \10934 );
or \U$2117 ( \10936 , \9492 , \10935 );
not \U$2118 ( \10937 , \8834 );
not \U$2119 ( \10938 , \10923 );
or \U$2120 ( \10939 , \10937 , \10938 );
not \U$2121 ( \10940 , \10939 );
and \U$2122 ( \10941 , \10918 , \10940 );
nand \U$2123 ( \10942 , \10941 , \10932 );
not \U$2124 ( \10943 , \10942 );
not \U$2125 ( \10944 , \10943 );
or \U$2126 ( \10945 , \9494 , \10944 );
nand \U$2127 ( \10946 , \10936 , \10945 );
not \U$2128 ( \10947 , \10923 );
not \U$2129 ( \10948 , \10947 );
or \U$2130 ( \10949 , \10920 , \10948 );
not \U$2131 ( \10950 , \10949 );
not \U$2132 ( \10951 , \10918 );
and \U$2133 ( \10952 , \10950 , \10951 );
nand \U$2134 ( \10953 , \10952 , \10932 );
not \U$2135 ( \10954 , \10953 );
not \U$2136 ( \10955 , \10954 );
or \U$2137 ( \10956 , \9498 , \10955 );
not \U$2138 ( \10957 , \10947 );
or \U$2139 ( \10958 , \8870 , \10957 );
not \U$2140 ( \10959 , \10958 );
and \U$2141 ( \10960 , \10959 , \10951 );
nand \U$2142 ( \10961 , \10960 , \10932 );
not \U$2143 ( \10962 , \10961 );
not \U$2144 ( \10963 , \10962 );
or \U$2145 ( \10964 , \9500 , \10963 );
nand \U$2146 ( \10965 , \10956 , \10964 );
nor \U$2147 ( \10966 , \10946 , \10965 );
nand \U$2148 ( \10967 , \10940 , \10951 );
not \U$2149 ( \10968 , \10967 );
and \U$2150 ( \10969 , \10968 , \10932 );
not \U$2151 ( \10970 , \10969 );
or \U$2152 ( \10971 , \9506 , \10970 );
and \U$2153 ( \10972 , \10926 , \10951 );
nand \U$2154 ( \10973 , \10931 , \10972 );
or \U$2155 ( \10974 , \9509 , \10973 );
nand \U$2156 ( \10975 , \10971 , \10974 );
not \U$2157 ( \10976 , \9504 );
not \U$2158 ( \10977 , \10976 );
and \U$2159 ( \10978 , \10950 , \10918 );
nand \U$2160 ( \10979 , \10931 , \10978 );
or \U$2161 ( \10980 , \10977 , \10979 );
and \U$2162 ( \10981 , \10931 , \10960 );
not \U$2163 ( \10982 , \10981 );
or \U$2164 ( \10983 , \9511 , \10982 );
nand \U$2165 ( \10984 , \10980 , \10983 );
nor \U$2166 ( \10985 , \10975 , \10984 );
not \U$2167 ( \10986 , \9463 );
nand \U$2168 ( \10987 , \10931 , \10968 );
not \U$2169 ( \10988 , \10987 );
and \U$2170 ( \10989 , \10986 , \10988 );
nand \U$2171 ( \10990 , \10931 , \10952 );
buf \U$2172 ( \10991 , \10990 );
not \U$2173 ( \10992 , \10991 );
and \U$2174 ( \10993 , \9468 , \10992 );
nor \U$2175 ( \10994 , \10989 , \10993 );
nand \U$2176 ( \10995 , \10931 , \10927 );
buf \U$2177 ( \10996 , \10995 );
not \U$2178 ( \10997 , \10996 );
and \U$2179 ( \10998 , \9472 , \10997 );
nand \U$2180 ( \10999 , \10931 , \10941 );
buf \U$2181 ( \11000 , \10999 );
not \U$2182 ( \11001 , \11000 );
and \U$2183 ( \11002 , \9476 , \11001 );
nor \U$2184 ( \11003 , \10998 , \11002 );
nand \U$2185 ( \11004 , \10994 , \11003 );
not \U$2186 ( \11005 , \9487 );
and \U$2187 ( \11006 , \10959 , \10918 );
nand \U$2188 ( \11007 , \11006 , \10932 );
not \U$2189 ( \11008 , \11007 );
not \U$2190 ( \11009 , \11008 );
not \U$2191 ( \11010 , \11009 );
and \U$2192 ( \11011 , \11005 , \11010 );
nand \U$2193 ( \11012 , \10978 , \10932 );
not \U$2194 ( \11013 , \11012 );
not \U$2195 ( \11014 , \11013 );
not \U$2196 ( \11015 , \11014 );
and \U$2197 ( \11016 , \11015 , \10168 );
nor \U$2198 ( \11017 , \11011 , \11016 );
not \U$2199 ( \11018 , \9482 );
nand \U$2200 ( \11019 , \10931 , \11006 );
not \U$2201 ( \11020 , \11019 );
and \U$2202 ( \11021 , \11018 , \11020 );
nand \U$2203 ( \11022 , \10972 , \10932 );
not \U$2204 ( \11023 , \11022 );
and \U$2205 ( \11024 , \11023 , \10152 );
nor \U$2206 ( \11025 , \11021 , \11024 );
nand \U$2207 ( \11026 , \11017 , \11025 );
nor \U$2208 ( \11027 , \11004 , \11026 );
nand \U$2209 ( \11028 , \10966 , \10985 , \11027 );
not \U$2210 ( \11029 , \11028 );
not \U$2211 ( \11030 , \8971 );
and \U$2212 ( \11031 , \11030 , \11020 );
nand \U$2213 ( \11032 , \10931 , \10978 );
not \U$2214 ( \11033 , \11032 );
and \U$2215 ( \11034 , \11033 , \8979 );
nor \U$2216 ( \11035 , \11031 , \11034 );
not \U$2217 ( \11036 , \9020 );
not \U$2218 ( \11037 , \11036 );
nand \U$2219 ( \11038 , \10931 , \10972 );
not \U$2220 ( \11039 , \11038 );
and \U$2221 ( \11040 , \11037 , \11039 );
and \U$2222 ( \11041 , \11023 , \9025 );
nor \U$2223 ( \11042 , \11040 , \11041 );
nand \U$2224 ( \11043 , \10931 , \10952 );
buf \U$2225 ( \11044 , \11043 );
or \U$2226 ( \11045 , \8991 , \11044 );
not \U$2227 ( \11046 , \8986 );
nand \U$2228 ( \11047 , \10931 , \10968 );
or \U$2229 ( \11048 , \11046 , \11047 );
nand \U$2230 ( \11049 , \11045 , \11048 );
nand \U$2231 ( \11050 , \10931 , \10927 );
buf \U$2232 ( \11051 , \11050 );
or \U$2233 ( \11052 , \8997 , \11051 );
not \U$2234 ( \11053 , \10981 );
or \U$2235 ( \11054 , \9000 , \11053 );
nand \U$2236 ( \11055 , \11052 , \11054 );
nor \U$2237 ( \11056 , \11049 , \11055 );
nand \U$2238 ( \11057 , \11035 , \11042 , \11056 );
not \U$2239 ( \11058 , \9014 );
or \U$2240 ( \11059 , \11058 , \10963 );
not \U$2241 ( \11060 , \9011 );
not \U$2242 ( \11061 , \10934 );
or \U$2243 ( \11062 , \11060 , \11061 );
nand \U$2244 ( \11063 , \11059 , \11062 );
not \U$2245 ( \11064 , \9034 );
not \U$2246 ( \11065 , \10954 );
or \U$2247 ( \11066 , \11064 , \11065 );
not \U$2248 ( \11067 , \9030 );
not \U$2249 ( \11068 , \10969 );
or \U$2250 ( \11069 , \11067 , \11068 );
nand \U$2251 ( \11070 , \11066 , \11069 );
nor \U$2252 ( \11071 , \11063 , \11070 );
or \U$2253 ( \11072 , \8967 , \11009 );
not \U$2254 ( \11073 , \9009 );
nand \U$2255 ( \11074 , \10931 , \10941 );
buf \U$2256 ( \11075 , \11074 );
or \U$2257 ( \11076 , \11073 , \11075 );
nand \U$2258 ( \11077 , \11072 , \11076 );
not \U$2259 ( \11078 , \8976 );
or \U$2260 ( \11079 , \11078 , \11014 );
not \U$2261 ( \11080 , \9006 );
not \U$2262 ( \11081 , \10943 );
or \U$2263 ( \11082 , \11080 , \11081 );
nand \U$2264 ( \11083 , \11079 , \11082 );
nor \U$2265 ( \11084 , \11077 , \11083 );
nand \U$2266 ( \11085 , \11071 , \11084 );
nor \U$2267 ( \11086 , \11057 , \11085 );
xnor \U$2268 ( \11087 , \11086 , \9044 );
not \U$2269 ( \11088 , \9193 );
not \U$2270 ( \11089 , \11088 );
and \U$2271 ( \11090 , \11089 , \11020 );
and \U$2272 ( \11091 , \11033 , \9200 );
nor \U$2273 ( \11092 , \11090 , \11091 );
not \U$2274 ( \11093 , \9239 );
not \U$2275 ( \11094 , \11093 );
and \U$2276 ( \11095 , \11094 , \11039 );
and \U$2277 ( \11096 , \11023 , \9242 );
nor \U$2278 ( \11097 , \11095 , \11096 );
not \U$2279 ( \11098 , \9212 );
buf \U$2280 ( \11099 , \11043 );
or \U$2281 ( \11100 , \11098 , \11099 );
not \U$2282 ( \11101 , \9210 );
nand \U$2283 ( \11102 , \10931 , \10968 );
or \U$2284 ( \11103 , \11101 , \11102 );
nand \U$2285 ( \11104 , \11100 , \11103 );
buf \U$2286 ( \11105 , \11050 );
or \U$2287 ( \11106 , \9217 , \11105 );
or \U$2288 ( \11107 , \9220 , \10982 );
nand \U$2289 ( \11108 , \11106 , \11107 );
nor \U$2290 ( \11109 , \11104 , \11108 );
nand \U$2291 ( \11110 , \11092 , \11097 , \11109 );
not \U$2292 ( \11111 , \9233 );
or \U$2293 ( \11112 , \11111 , \10963 );
not \U$2294 ( \11113 , \9230 );
not \U$2295 ( \11114 , \10934 );
or \U$2296 ( \11115 , \11113 , \11114 );
nand \U$2297 ( \11116 , \11112 , \11115 );
not \U$2298 ( \11117 , \9251 );
not \U$2299 ( \11118 , \10954 );
or \U$2300 ( \11119 , \11117 , \11118 );
not \U$2301 ( \11120 , \9247 );
or \U$2302 ( \11121 , \11120 , \11068 );
nand \U$2303 ( \11122 , \11119 , \11121 );
nor \U$2304 ( \11123 , \11116 , \11122 );
or \U$2305 ( \11124 , \9197 , \11009 );
not \U$2306 ( \11125 , \9228 );
buf \U$2307 ( \11126 , \11074 );
or \U$2308 ( \11127 , \11125 , \11126 );
nand \U$2309 ( \11128 , \11124 , \11127 );
not \U$2310 ( \11129 , \9204 );
or \U$2311 ( \11130 , \11129 , \11014 );
not \U$2312 ( \11131 , \10943 );
or \U$2313 ( \11132 , \9226 , \11131 );
nand \U$2314 ( \11133 , \11130 , \11132 );
nor \U$2315 ( \11134 , \11128 , \11133 );
nand \U$2316 ( \11135 , \11123 , \11134 );
nor \U$2317 ( \11136 , \11110 , \11135 );
xnor \U$2318 ( \11137 , \11136 , \9260 );
not \U$2319 ( \11138 , \9706 );
or \U$2320 ( \11139 , \11138 , \10979 );
not \U$2321 ( \11140 , \9701 );
or \U$2322 ( \11141 , \11140 , \11126 );
nand \U$2323 ( \11142 , \11139 , \11141 );
nand \U$2324 ( \11143 , \10972 , \10932 );
or \U$2325 ( \11144 , \10244 , \11143 );
not \U$2326 ( \11145 , \9710 );
or \U$2327 ( \11146 , \11145 , \11019 );
nand \U$2328 ( \11147 , \11144 , \11146 );
nor \U$2329 ( \11148 , \11142 , \11147 );
or \U$2330 ( \11149 , \10248 , \10955 );
or \U$2331 ( \11150 , \10250 , \11068 );
nand \U$2332 ( \11151 , \11149 , \11150 );
not \U$2333 ( \11152 , \9687 );
or \U$2334 ( \11153 , \11152 , \11061 );
not \U$2335 ( \11154 , \9690 );
or \U$2336 ( \11155 , \11154 , \10963 );
nand \U$2337 ( \11156 , \11153 , \11155 );
nor \U$2338 ( \11157 , \11151 , \11156 );
not \U$2339 ( \11158 , \11053 );
and \U$2340 ( \11159 , \9682 , \11158 );
buf \U$2341 ( \11160 , \10995 );
not \U$2342 ( \11161 , \11160 );
and \U$2343 ( \11162 , \9679 , \11161 );
nor \U$2344 ( \11163 , \11159 , \11162 );
not \U$2345 ( \11164 , \11047 );
and \U$2346 ( \11165 , \9672 , \11164 );
not \U$2347 ( \11166 , \11044 );
and \U$2348 ( \11167 , \9675 , \11166 );
nor \U$2349 ( \11168 , \11165 , \11167 );
nand \U$2350 ( \11169 , \11163 , \11168 );
and \U$2351 ( \11170 , \11010 , \9664 );
and \U$2352 ( \11171 , \9667 , \11039 );
nor \U$2353 ( \11172 , \11170 , \11171 );
and \U$2354 ( \11173 , \11015 , \9656 );
not \U$2355 ( \11174 , \11081 );
and \U$2356 ( \11175 , \9660 , \11174 );
nor \U$2357 ( \11176 , \11173 , \11175 );
nand \U$2358 ( \11177 , \11172 , \11176 );
nor \U$2359 ( \11178 , \11169 , \11177 );
nand \U$2360 ( \11179 , \11148 , \11157 , \11178 );
xnor \U$2361 ( \11180 , \11179 , \9719 );
or \U$2362 ( \11181 , \10178 , \11032 );
buf \U$2363 ( \11182 , \10999 );
or \U$2364 ( \11183 , \10182 , \11182 );
nand \U$2365 ( \11184 , \11181 , \11183 );
or \U$2366 ( \11185 , \10188 , \11022 );
not \U$2367 ( \11186 , \9776 );
or \U$2368 ( \11187 , \11186 , \11019 );
nand \U$2369 ( \11188 , \11185 , \11187 );
nor \U$2370 ( \11189 , \11184 , \11188 );
or \U$2371 ( \11190 , \10194 , \10955 );
or \U$2372 ( \11191 , \10197 , \10970 );
nand \U$2373 ( \11192 , \11190 , \11191 );
not \U$2374 ( \11193 , \9752 );
or \U$2375 ( \11194 , \11193 , \10935 );
not \U$2376 ( \11195 , \9755 );
or \U$2377 ( \11196 , \11195 , \10963 );
nand \U$2378 ( \11197 , \11194 , \11196 );
nor \U$2379 ( \11198 , \11192 , \11197 );
not \U$2380 ( \11199 , \10981 );
not \U$2381 ( \11200 , \11199 );
and \U$2382 ( \11201 , \9747 , \11200 );
nand \U$2383 ( \11202 , \10931 , \10927 );
buf \U$2384 ( \11203 , \11202 );
not \U$2385 ( \11204 , \11203 );
and \U$2386 ( \11205 , \9744 , \11204 );
nor \U$2387 ( \11206 , \11201 , \11205 );
not \U$2388 ( \11207 , \11102 );
and \U$2389 ( \11208 , \9736 , \11207 );
buf \U$2390 ( \11209 , \10990 );
not \U$2391 ( \11210 , \11209 );
and \U$2392 ( \11211 , \9739 , \11210 );
nor \U$2393 ( \11212 , \11208 , \11211 );
nand \U$2394 ( \11213 , \11206 , \11212 );
and \U$2395 ( \11214 , \11010 , \9728 );
and \U$2396 ( \11215 , \9731 , \11039 );
nor \U$2397 ( \11216 , \11214 , \11215 );
and \U$2398 ( \11217 , \11015 , \9721 );
and \U$2399 ( \11218 , \9724 , \11174 );
nor \U$2400 ( \11219 , \11217 , \11218 );
nand \U$2401 ( \11220 , \11216 , \11219 );
nor \U$2402 ( \11221 , \11213 , \11220 );
nand \U$2403 ( \11222 , \11189 , \11198 , \11221 );
xnor \U$2404 ( \11223 , \11222 , \9786 );
nor \U$2405 ( \11224 , \11180 , \11223 );
nand \U$2406 ( \11225 , \11087 , \11137 , \11224 );
not \U$2407 ( \11226 , \9398 );
and \U$2408 ( \11227 , \11226 , \11020 );
and \U$2409 ( \11228 , \11033 , \9404 );
nor \U$2410 ( \11229 , \11227 , \11228 );
not \U$2411 ( \11230 , \9440 );
not \U$2412 ( \11231 , \11230 );
and \U$2413 ( \11232 , \11231 , \11039 );
and \U$2414 ( \11233 , \11023 , \9444 );
nor \U$2415 ( \11234 , \11232 , \11233 );
or \U$2416 ( \11235 , \9415 , \10991 );
or \U$2417 ( \11236 , \10455 , \11102 );
nand \U$2418 ( \11237 , \11235 , \11236 );
or \U$2419 ( \11238 , \9419 , \11203 );
or \U$2420 ( \11239 , \9422 , \10982 );
nand \U$2421 ( \11240 , \11238 , \11239 );
nor \U$2422 ( \11241 , \11237 , \11240 );
nand \U$2423 ( \11242 , \11229 , \11234 , \11241 );
not \U$2424 ( \11243 , \9435 );
or \U$2425 ( \11244 , \11243 , \10963 );
not \U$2426 ( \11245 , \9432 );
or \U$2427 ( \11246 , \11245 , \11114 );
nand \U$2428 ( \11247 , \11244 , \11246 );
not \U$2429 ( \11248 , \9453 );
or \U$2430 ( \11249 , \11248 , \11118 );
not \U$2431 ( \11250 , \9449 );
or \U$2432 ( \11251 , \11250 , \10970 );
nand \U$2433 ( \11252 , \11249 , \11251 );
nor \U$2434 ( \11253 , \11247 , \11252 );
or \U$2435 ( \11254 , \9395 , \11009 );
or \U$2436 ( \11255 , \10464 , \11075 );
nand \U$2437 ( \11256 , \11254 , \11255 );
not \U$2438 ( \11257 , \9401 );
or \U$2439 ( \11258 , \11257 , \11014 );
not \U$2440 ( \11259 , \9427 );
or \U$2441 ( \11260 , \11259 , \11131 );
nand \U$2442 ( \11261 , \11258 , \11260 );
nor \U$2443 ( \11262 , \11256 , \11261 );
nand \U$2444 ( \11263 , \11253 , \11262 );
nor \U$2445 ( \11264 , \11242 , \11263 );
xnor \U$2446 ( \11265 , \11264 , \9460 );
not \U$2447 ( \11266 , \9266 );
and \U$2448 ( \11267 , \11266 , \11020 );
and \U$2449 ( \11268 , \11033 , \9272 );
nor \U$2450 ( \11269 , \11267 , \11268 );
not \U$2451 ( \11270 , \9307 );
not \U$2452 ( \11271 , \11270 );
and \U$2453 ( \11272 , \11271 , \11039 );
and \U$2454 ( \11273 , \11023 , \9310 );
nor \U$2455 ( \11274 , \11272 , \11273 );
or \U$2456 ( \11275 , \9282 , \11044 );
not \U$2457 ( \11276 , \9277 );
or \U$2458 ( \11277 , \11276 , \10987 );
nand \U$2459 ( \11278 , \11275 , \11277 );
buf \U$2460 ( \11279 , \11202 );
or \U$2461 ( \11280 , \9287 , \11279 );
not \U$2462 ( \11281 , \10981 );
or \U$2463 ( \11282 , \9290 , \11281 );
nand \U$2464 ( \11283 , \11280 , \11282 );
nor \U$2465 ( \11284 , \11278 , \11283 );
nand \U$2466 ( \11285 , \11269 , \11274 , \11284 );
not \U$2467 ( \11286 , \9302 );
or \U$2468 ( \11287 , \11286 , \10963 );
not \U$2469 ( \11288 , \9299 );
or \U$2470 ( \11289 , \11288 , \11061 );
nand \U$2471 ( \11290 , \11287 , \11289 );
not \U$2472 ( \11291 , \9319 );
or \U$2473 ( \11292 , \11291 , \11065 );
not \U$2474 ( \11293 , \9315 );
or \U$2475 ( \11294 , \11293 , \11068 );
nand \U$2476 ( \11295 , \11292 , \11294 );
nor \U$2477 ( \11296 , \11290 , \11295 );
or \U$2478 ( \11297 , \9263 , \11009 );
not \U$2479 ( \11298 , \9297 );
or \U$2480 ( \11299 , \11298 , \11000 );
nand \U$2481 ( \11300 , \11297 , \11299 );
not \U$2482 ( \11301 , \9269 );
or \U$2483 ( \11302 , \11301 , \11014 );
not \U$2484 ( \11303 , \9295 );
or \U$2485 ( \11304 , \11303 , \11131 );
nand \U$2486 ( \11305 , \11302 , \11304 );
nor \U$2487 ( \11306 , \11300 , \11305 );
nand \U$2488 ( \11307 , \11296 , \11306 );
nor \U$2489 ( \11308 , \11285 , \11307 );
xnor \U$2490 ( \11309 , \11308 , \9327 );
or \U$2491 ( \11310 , \9620 , \11065 );
or \U$2492 ( \11311 , \9625 , \11068 );
nand \U$2493 ( \11312 , \11310 , \11311 );
or \U$2494 ( \11313 , \9632 , \11061 );
not \U$2495 ( \11314 , \9628 );
or \U$2496 ( \11315 , \11314 , \10963 );
nand \U$2497 ( \11316 , \11313 , \11315 );
nor \U$2498 ( \11317 , \11312 , \11316 );
or \U$2499 ( \11318 , \9640 , \11081 );
nand \U$2500 ( \11319 , \10972 , \10932 );
or \U$2501 ( \11320 , \9611 , \11319 );
nand \U$2502 ( \11321 , \11318 , \11320 );
not \U$2503 ( \11322 , \9643 );
or \U$2504 ( \11323 , \11322 , \11009 );
or \U$2505 ( \11324 , \9637 , \11014 );
nand \U$2506 ( \11325 , \11323 , \11324 );
nor \U$2507 ( \11326 , \11321 , \11325 );
not \U$2508 ( \11327 , \10981 );
not \U$2509 ( \11328 , \11327 );
and \U$2510 ( \11329 , \9593 , \11328 );
not \U$2511 ( \11330 , \11279 );
and \U$2512 ( \11331 , \9587 , \11330 );
nor \U$2513 ( \11332 , \11329 , \11331 );
not \U$2514 ( \11333 , \10987 );
and \U$2515 ( \11334 , \9596 , \11333 );
not \U$2516 ( \11335 , \10991 );
and \U$2517 ( \11336 , \9600 , \11335 );
nor \U$2518 ( \11337 , \11334 , \11336 );
nand \U$2519 ( \11338 , \11332 , \11337 );
not \U$2520 ( \11339 , \11020 );
or \U$2521 ( \11340 , \9614 , \11339 );
not \U$2522 ( \11341 , \11033 );
or \U$2523 ( \11342 , \9604 , \11341 );
not \U$2524 ( \11343 , \11038 );
and \U$2525 ( \11344 , \9646 , \11343 );
not \U$2526 ( \11345 , \11075 );
and \U$2527 ( \11346 , \9606 , \11345 );
nor \U$2528 ( \11347 , \11344 , \11346 );
nand \U$2529 ( \11348 , \11340 , \11342 , \11347 );
nor \U$2530 ( \11349 , \11338 , \11348 );
nand \U$2531 ( \11350 , \11317 , \11326 , \11349 );
xnor \U$2532 ( \11351 , \11350 , \9653 );
not \U$2533 ( \11352 , \9361 );
not \U$2534 ( \11353 , \11352 );
and \U$2535 ( \11354 , \11353 , \11174 );
and \U$2536 ( \11355 , \11015 , \9338 );
nor \U$2537 ( \11356 , \11354 , \11355 );
not \U$2538 ( \11357 , \9364 );
not \U$2539 ( \11358 , \11357 );
not \U$2540 ( \11359 , \11075 );
and \U$2541 ( \11360 , \11358 , \11359 );
and \U$2542 ( \11361 , \11010 , \9331 );
nor \U$2543 ( \11362 , \11360 , \11361 );
nand \U$2544 ( \11363 , \11356 , \11362 );
not \U$2545 ( \11364 , \11363 );
not \U$2546 ( \11365 , \9366 );
not \U$2547 ( \11366 , \11365 );
not \U$2548 ( \11367 , \11061 );
and \U$2549 ( \11368 , \11366 , \11367 );
and \U$2550 ( \11369 , \10962 , \9369 );
nor \U$2551 ( \11370 , \11368 , \11369 );
not \U$2552 ( \11371 , \9377 );
not \U$2553 ( \11372 , \11371 );
and \U$2554 ( \11373 , \11372 , \10954 );
not \U$2555 ( \11374 , \10970 );
and \U$2556 ( \11375 , \11374 , \9385 );
nor \U$2557 ( \11376 , \11373 , \11375 );
and \U$2558 ( \11377 , \11364 , \11370 , \11376 );
not \U$2559 ( \11378 , \11053 );
and \U$2560 ( \11379 , \9356 , \11378 );
not \U$2561 ( \11380 , \11203 );
and \U$2562 ( \11381 , \9353 , \11380 );
nor \U$2563 ( \11382 , \11379 , \11381 );
not \U$2564 ( \11383 , \11047 );
and \U$2565 ( \11384 , \9346 , \11383 );
not \U$2566 ( \11385 , \11099 );
and \U$2567 ( \11386 , \9348 , \11385 );
nor \U$2568 ( \11387 , \11384 , \11386 );
nand \U$2569 ( \11388 , \11382 , \11387 );
nand \U$2570 ( \11389 , \10931 , \10978 );
or \U$2571 ( \11390 , \9342 , \11389 );
not \U$2572 ( \11391 , \11023 );
or \U$2573 ( \11392 , \10553 , \11391 );
not \U$2574 ( \11393 , \9374 );
not \U$2575 ( \11394 , \11039 );
or \U$2576 ( \11395 , \11393 , \11394 );
not \U$2577 ( \11396 , \11020 );
or \U$2578 ( \11397 , \9335 , \11396 );
and \U$2579 ( \11398 , \11390 , \11392 , \11395 , \11397 );
not \U$2580 ( \11399 , \11398 );
nor \U$2581 ( \11400 , \11388 , \11399 );
nand \U$2582 ( \11401 , \11377 , \11400 );
xnor \U$2583 ( \11402 , \11401 , \9392 );
nor \U$2584 ( \11403 , \11351 , \11402 );
nand \U$2585 ( \11404 , \11265 , \11309 , \11403 );
nor \U$2586 ( \11405 , \11225 , \11404 );
not \U$2587 ( \11406 , \9125 );
and \U$2588 ( \11407 , \11406 , \11020 );
and \U$2589 ( \11408 , \11033 , \9132 );
nor \U$2590 ( \11409 , \11407 , \11408 );
not \U$2591 ( \11410 , \9168 );
not \U$2592 ( \11411 , \11410 );
and \U$2593 ( \11412 , \11411 , \11039 );
and \U$2594 ( \11413 , \11023 , \9172 );
nor \U$2595 ( \11414 , \11412 , \11413 );
or \U$2596 ( \11415 , \9143 , \11209 );
not \U$2597 ( \11416 , \9137 );
or \U$2598 ( \11417 , \11416 , \10987 );
nand \U$2599 ( \11418 , \11415 , \11417 );
or \U$2600 ( \11419 , \9148 , \11051 );
or \U$2601 ( \11420 , \9151 , \11281 );
nand \U$2602 ( \11421 , \11419 , \11420 );
nor \U$2603 ( \11422 , \11418 , \11421 );
nand \U$2604 ( \11423 , \11409 , \11414 , \11422 );
not \U$2605 ( \11424 , \9163 );
or \U$2606 ( \11425 , \11424 , \10963 );
not \U$2607 ( \11426 , \9159 );
or \U$2608 ( \11427 , \11426 , \11061 );
nand \U$2609 ( \11428 , \11425 , \11427 );
not \U$2610 ( \11429 , \9180 );
or \U$2611 ( \11430 , \11429 , \11118 );
not \U$2612 ( \11431 , \9176 );
or \U$2613 ( \11432 , \11431 , \11068 );
nand \U$2614 ( \11433 , \11430 , \11432 );
nor \U$2615 ( \11434 , \11428 , \11433 );
or \U$2616 ( \11435 , \9122 , \11009 );
not \U$2617 ( \11436 , \9157 );
or \U$2618 ( \11437 , \11436 , \11126 );
nand \U$2619 ( \11438 , \11435 , \11437 );
not \U$2620 ( \11439 , \9129 );
or \U$2621 ( \11440 , \11439 , \11014 );
not \U$2622 ( \11441 , \9155 );
or \U$2623 ( \11442 , \11441 , \11081 );
nand \U$2624 ( \11443 , \11440 , \11442 );
nor \U$2625 ( \11444 , \11438 , \11443 );
nand \U$2626 ( \11445 , \11434 , \11444 );
nor \U$2627 ( \11446 , \11423 , \11445 );
xnor \U$2628 ( \11447 , \11446 , \9188 );
not \U$2629 ( \11448 , \9050 );
and \U$2630 ( \11449 , \11448 , \11020 );
and \U$2631 ( \11450 , \11033 , \9057 );
nor \U$2632 ( \11451 , \11449 , \11450 );
not \U$2633 ( \11452 , \9098 );
not \U$2634 ( \11453 , \11452 );
and \U$2635 ( \11454 , \11453 , \11039 );
and \U$2636 ( \11455 , \11023 , \9102 );
nor \U$2637 ( \11456 , \11454 , \11455 );
or \U$2638 ( \11457 , \9068 , \10991 );
not \U$2639 ( \11458 , \9063 );
or \U$2640 ( \11459 , \11458 , \11047 );
nand \U$2641 ( \11460 , \11457 , \11459 );
or \U$2642 ( \11461 , \9073 , \11105 );
or \U$2643 ( \11462 , \9076 , \11281 );
nand \U$2644 ( \11463 , \11461 , \11462 );
nor \U$2645 ( \11464 , \11460 , \11463 );
nand \U$2646 ( \11465 , \11451 , \11456 , \11464 );
not \U$2647 ( \11466 , \9093 );
or \U$2648 ( \11467 , \11466 , \10963 );
not \U$2649 ( \11468 , \9089 );
or \U$2650 ( \11469 , \11468 , \11114 );
nand \U$2651 ( \11470 , \11467 , \11469 );
not \U$2652 ( \11471 , \9112 );
or \U$2653 ( \11472 , \11471 , \10955 );
not \U$2654 ( \11473 , \9107 );
or \U$2655 ( \11474 , \11473 , \11068 );
nand \U$2656 ( \11475 , \11472 , \11474 );
nor \U$2657 ( \11476 , \11470 , \11475 );
or \U$2658 ( \11477 , \9047 , \11009 );
or \U$2659 ( \11478 , \9086 , \11182 );
nand \U$2660 ( \11479 , \11477 , \11478 );
not \U$2661 ( \11480 , \9054 );
or \U$2662 ( \11481 , \11480 , \11014 );
or \U$2663 ( \11482 , \9082 , \11081 );
nand \U$2664 ( \11483 , \11481 , \11482 );
nor \U$2665 ( \11484 , \11479 , \11483 );
nand \U$2666 ( \11485 , \11476 , \11484 );
nor \U$2667 ( \11486 , \11465 , \11485 );
xnor \U$2668 ( \11487 , \11486 , \9119 );
not \U$2669 ( \11488 , \9813 );
or \U$2670 ( \11489 , \11488 , \11022 );
or \U$2671 ( \11490 , \9798 , \10987 );
nand \U$2672 ( \11491 , \11489 , \11490 );
not \U$2673 ( \11492 , \9794 );
or \U$2674 ( \11493 , \11492 , \10982 );
not \U$2675 ( \11494 , \9801 );
or \U$2676 ( \11495 , \11494 , \11099 );
nand \U$2677 ( \11496 , \11493 , \11495 );
nor \U$2678 ( \11497 , \11491 , \11496 );
or \U$2679 ( \11498 , \9809 , \11000 );
or \U$2680 ( \11499 , \9851 , \11038 );
nand \U$2681 ( \11500 , \11498 , \11499 );
or \U$2682 ( \11501 , \9817 , \11019 );
or \U$2683 ( \11502 , \9806 , \11389 );
nand \U$2684 ( \11503 , \11501 , \11502 );
nor \U$2685 ( \11504 , \11500 , \11503 );
not \U$2686 ( \11505 , \9847 );
not \U$2687 ( \11506 , \11010 );
or \U$2688 ( \11507 , \11505 , \11506 );
not \U$2689 ( \11508 , \11015 );
or \U$2690 ( \11509 , \9840 , \11508 );
not \U$2691 ( \11510 , \11160 );
and \U$2692 ( \11511 , \9790 , \11510 );
not \U$2693 ( \11512 , \10944 );
and \U$2694 ( \11513 , \9842 , \11512 );
nor \U$2695 ( \11514 , \11511 , \11513 );
nand \U$2696 ( \11515 , \11507 , \11509 , \11514 );
not \U$2697 ( \11516 , \9834 );
and \U$2698 ( \11517 , \11516 , \11367 );
and \U$2699 ( \11518 , \10962 , \9830 );
nor \U$2700 ( \11519 , \11517 , \11518 );
not \U$2701 ( \11520 , \9827 );
and \U$2702 ( \11521 , \11520 , \11374 );
and \U$2703 ( \11522 , \10954 , \9822 );
nor \U$2704 ( \11523 , \11521 , \11522 );
nand \U$2705 ( \11524 , \11519 , \11523 );
nor \U$2706 ( \11525 , \11515 , \11524 );
nand \U$2707 ( \11526 , \11497 , \11504 , \11525 );
xnor \U$2708 ( \11527 , \11526 , \9857 );
not \U$2709 ( \11528 , \8904 );
not \U$2710 ( \11529 , \11528 );
and \U$2711 ( \11530 , \11529 , \11174 );
and \U$2712 ( \11531 , \11015 , \8852 );
nor \U$2713 ( \11532 , \11530 , \11531 );
not \U$2714 ( \11533 , \8915 );
not \U$2715 ( \11534 , \11533 );
and \U$2716 ( \11535 , \11534 , \11359 );
and \U$2717 ( \11536 , \11010 , \8827 );
nor \U$2718 ( \11537 , \11535 , \11536 );
nand \U$2719 ( \11538 , \11532 , \11537 );
not \U$2720 ( \11539 , \11538 );
not \U$2721 ( \11540 , \8921 );
not \U$2722 ( \11541 , \11540 );
and \U$2723 ( \11542 , \11541 , \11367 );
and \U$2724 ( \11543 , \10962 , \8927 );
nor \U$2725 ( \11544 , \11542 , \11543 );
not \U$2726 ( \11545 , \8947 );
not \U$2727 ( \11546 , \11545 );
and \U$2728 ( \11547 , \11546 , \11374 );
and \U$2729 ( \11548 , \10954 , \8953 );
nor \U$2730 ( \11549 , \11547 , \11548 );
and \U$2731 ( \11550 , \11539 , \11544 , \11549 );
not \U$2732 ( \11551 , \11053 );
and \U$2733 ( \11552 , \8896 , \11551 );
not \U$2734 ( \11553 , \11051 );
and \U$2735 ( \11554 , \8893 , \11553 );
nor \U$2736 ( \11555 , \11552 , \11554 );
not \U$2737 ( \11556 , \11102 );
and \U$2738 ( \11557 , \8868 , \11556 );
not \U$2739 ( \11558 , \10991 );
and \U$2740 ( \11559 , \8881 , \11558 );
nor \U$2741 ( \11560 , \11557 , \11559 );
nand \U$2742 ( \11561 , \11555 , \11560 );
or \U$2743 ( \11562 , \8861 , \10979 );
not \U$2744 ( \11563 , \11023 );
or \U$2745 ( \11564 , \10775 , \11563 );
not \U$2746 ( \11565 , \8934 );
not \U$2747 ( \11566 , \11039 );
or \U$2748 ( \11567 , \11565 , \11566 );
not \U$2749 ( \11568 , \11020 );
or \U$2750 ( \11569 , \8844 , \11568 );
and \U$2751 ( \11570 , \11562 , \11564 , \11567 , \11569 );
not \U$2752 ( \11571 , \11570 );
nor \U$2753 ( \11572 , \11561 , \11571 );
nand \U$2754 ( \11573 , \11550 , \11572 );
xnor \U$2755 ( \11574 , \11573 , \8964 );
nor \U$2756 ( \11575 , \11527 , \11574 );
nand \U$2757 ( \11576 , \11447 , \11487 , \11575 );
not \U$2758 ( \11577 , \11576 );
or \U$2759 ( \11578 , \9552 , \10955 );
or \U$2760 ( \11579 , \9557 , \11068 );
nand \U$2761 ( \11580 , \11578 , \11579 );
or \U$2762 ( \11581 , \9564 , \10935 );
not \U$2763 ( \11582 , \9560 );
or \U$2764 ( \11583 , \11582 , \10963 );
nand \U$2765 ( \11584 , \11581 , \11583 );
nor \U$2766 ( \11585 , \11580 , \11584 );
or \U$2767 ( \11586 , \9572 , \11081 );
or \U$2768 ( \11587 , \9543 , \11143 );
nand \U$2769 ( \11588 , \11586 , \11587 );
not \U$2770 ( \11589 , \9575 );
or \U$2771 ( \11590 , \11589 , \11009 );
or \U$2772 ( \11591 , \9569 , \11014 );
nand \U$2773 ( \11592 , \11590 , \11591 );
nor \U$2774 ( \11593 , \11588 , \11592 );
not \U$2775 ( \11594 , \11199 );
and \U$2776 ( \11595 , \9523 , \11594 );
not \U$2777 ( \11596 , \11279 );
and \U$2778 ( \11597 , \9518 , \11596 );
nor \U$2779 ( \11598 , \11595 , \11597 );
not \U$2780 ( \11599 , \11102 );
and \U$2781 ( \11600 , \9526 , \11599 );
not \U$2782 ( \11601 , \11209 );
and \U$2783 ( \11602 , \9530 , \11601 );
nor \U$2784 ( \11603 , \11600 , \11602 );
nand \U$2785 ( \11604 , \11598 , \11603 );
not \U$2786 ( \11605 , \11020 );
or \U$2787 ( \11606 , \9546 , \11605 );
not \U$2788 ( \11607 , \11033 );
or \U$2789 ( \11608 , \9534 , \11607 );
not \U$2790 ( \11609 , \10973 );
and \U$2791 ( \11610 , \9578 , \11609 );
not \U$2792 ( \11611 , \11075 );
and \U$2793 ( \11612 , \9536 , \11611 );
nor \U$2794 ( \11613 , \11610 , \11612 );
nand \U$2795 ( \11614 , \11606 , \11608 , \11613 );
nor \U$2796 ( \11615 , \11604 , \11614 );
nand \U$2797 ( \11616 , \11585 , \11593 , \11615 );
xnor \U$2798 ( \11617 , \11616 , \9585 );
not \U$2799 ( \11618 , \9968 );
or \U$2800 ( \11619 , \11618 , \11118 );
not \U$2801 ( \11620 , \9965 );
or \U$2802 ( \11621 , \11620 , \11068 );
nand \U$2803 ( \11622 , \11619 , \11621 );
not \U$2804 ( \11623 , \9959 );
or \U$2805 ( \11624 , \11623 , \11061 );
not \U$2806 ( \11625 , \10709 );
or \U$2807 ( \11626 , \11625 , \10963 );
nand \U$2808 ( \11627 , \11624 , \11626 );
nor \U$2809 ( \11628 , \11622 , \11627 );
not \U$2810 ( \11629 , \9975 );
or \U$2811 ( \11630 , \11629 , \11081 );
or \U$2812 ( \11631 , \9937 , \11319 );
nand \U$2813 ( \11632 , \11630 , \11631 );
not \U$2814 ( \11633 , \9982 );
or \U$2815 ( \11634 , \11633 , \11009 );
not \U$2816 ( \11635 , \9977 );
or \U$2817 ( \11636 , \11635 , \11014 );
nand \U$2818 ( \11637 , \11634 , \11636 );
nor \U$2819 ( \11638 , \11632 , \11637 );
not \U$2820 ( \11639 , \10982 );
and \U$2821 ( \11640 , \9954 , \11639 );
not \U$2822 ( \11641 , \11051 );
and \U$2823 ( \11642 , \9951 , \11641 );
nor \U$2824 ( \11643 , \11640 , \11642 );
not \U$2825 ( \11644 , \10987 );
and \U$2826 ( \11645 , \9944 , \11644 );
not \U$2827 ( \11646 , \11044 );
and \U$2828 ( \11647 , \9947 , \11646 );
nor \U$2829 ( \11648 , \11645 , \11647 );
nand \U$2830 ( \11649 , \11643 , \11648 );
not \U$2831 ( \11650 , \11020 );
or \U$2832 ( \11651 , \9940 , \11650 );
not \U$2833 ( \11652 , \11033 );
or \U$2834 ( \11653 , \9930 , \11652 );
not \U$2835 ( \11654 , \11038 );
and \U$2836 ( \11655 , \9984 , \11654 );
not \U$2837 ( \11656 , \11000 );
and \U$2838 ( \11657 , \9932 , \11656 );
nor \U$2839 ( \11658 , \11655 , \11657 );
nand \U$2840 ( \11659 , \11651 , \11653 , \11658 );
nor \U$2841 ( \11660 , \11649 , \11659 );
nand \U$2842 ( \11661 , \11628 , \11638 , \11660 );
xnor \U$2843 ( \11662 , \11661 , \9990 );
nor \U$2844 ( \11663 , \11617 , \11662 );
not \U$2845 ( \11664 , \10017 );
or \U$2846 ( \11665 , \11664 , \11143 );
not \U$2847 ( \11666 , \9992 );
or \U$2848 ( \11667 , \11666 , \11047 );
nand \U$2849 ( \11668 , \11665 , \11667 );
or \U$2850 ( \11669 , \10005 , \11199 );
or \U$2851 ( \11670 , \9997 , \11209 );
nand \U$2852 ( \11671 , \11669 , \11670 );
nor \U$2853 ( \11672 , \11668 , \11671 );
or \U$2854 ( \11673 , \10013 , \11075 );
not \U$2855 ( \11674 , \10049 );
or \U$2856 ( \11675 , \11674 , \10973 );
nand \U$2857 ( \11676 , \11673 , \11675 );
or \U$2858 ( \11677 , \10021 , \11019 );
or \U$2859 ( \11678 , \10010 , \11032 );
nand \U$2860 ( \11679 , \11677 , \11678 );
nor \U$2861 ( \11680 , \11676 , \11679 );
not \U$2862 ( \11681 , \10047 );
not \U$2863 ( \11682 , \11010 );
or \U$2864 ( \11683 , \11681 , \11682 );
not \U$2865 ( \11684 , \10043 );
not \U$2866 ( \11685 , \11015 );
or \U$2867 ( \11686 , \11684 , \11685 );
not \U$2868 ( \11687 , \11105 );
and \U$2869 ( \11688 , \10001 , \11687 );
not \U$2870 ( \11689 , \10944 );
and \U$2871 ( \11690 , \11689 , \10041 );
nor \U$2872 ( \11691 , \11688 , \11690 );
nand \U$2873 ( \11692 , \11683 , \11686 , \11691 );
not \U$2874 ( \11693 , \10025 );
not \U$2875 ( \11694 , \11693 );
and \U$2876 ( \11695 , \11694 , \11367 );
and \U$2877 ( \11696 , \10962 , \10027 );
nor \U$2878 ( \11697 , \11695 , \11696 );
not \U$2879 ( \11698 , \10030 );
not \U$2880 ( \11699 , \11698 );
and \U$2881 ( \11700 , \11699 , \11374 );
and \U$2882 ( \11701 , \10954 , \10035 );
nor \U$2883 ( \11702 , \11700 , \11701 );
nand \U$2884 ( \11703 , \11697 , \11702 );
nor \U$2885 ( \11704 , \11692 , \11703 );
nand \U$2886 ( \11705 , \11672 , \11680 , \11704 );
xnor \U$2887 ( \11706 , \11705 , \10055 );
or \U$2888 ( \11707 , \9895 , \11065 );
or \U$2889 ( \11708 , \9898 , \11068 );
nand \U$2890 ( \11709 , \11707 , \11708 );
or \U$2891 ( \11710 , \9906 , \11061 );
not \U$2892 ( \11711 , \9902 );
or \U$2893 ( \11712 , \11711 , \10963 );
nand \U$2894 ( \11713 , \11710 , \11712 );
nor \U$2895 ( \11714 , \11709 , \11713 );
or \U$2896 ( \11715 , \9914 , \11131 );
or \U$2897 ( \11716 , \9884 , \11319 );
nand \U$2898 ( \11717 , \11715 , \11716 );
not \U$2899 ( \11718 , \9917 );
or \U$2900 ( \11719 , \11718 , \11009 );
or \U$2901 ( \11720 , \9911 , \11014 );
nand \U$2902 ( \11721 , \11719 , \11720 );
nor \U$2903 ( \11722 , \11717 , \11721 );
not \U$2904 ( \11723 , \11281 );
and \U$2905 ( \11724 , \9864 , \11723 );
not \U$2906 ( \11725 , \10996 );
and \U$2907 ( \11726 , \9859 , \11725 );
nor \U$2908 ( \11727 , \11724 , \11726 );
not \U$2909 ( \11728 , \11047 );
and \U$2910 ( \11729 , \9867 , \11728 );
not \U$2911 ( \11730 , \11099 );
and \U$2912 ( \11731 , \9871 , \11730 );
nor \U$2913 ( \11732 , \11729 , \11731 );
nand \U$2914 ( \11733 , \11727 , \11732 );
not \U$2915 ( \11734 , \11020 );
or \U$2916 ( \11735 , \9887 , \11734 );
not \U$2917 ( \11736 , \11033 );
or \U$2918 ( \11737 , \9875 , \11736 );
not \U$2919 ( \11738 , \10973 );
and \U$2920 ( \11739 , \9920 , \11738 );
not \U$2921 ( \11740 , \11182 );
and \U$2922 ( \11741 , \9877 , \11740 );
nor \U$2923 ( \11742 , \11739 , \11741 );
nand \U$2924 ( \11743 , \11735 , \11737 , \11742 );
nor \U$2925 ( \11744 , \11733 , \11743 );
nand \U$2926 ( \11745 , \11714 , \11722 , \11744 );
xnor \U$2927 ( \11746 , \11745 , \9927 );
nor \U$2928 ( \11747 , \11706 , \11746 );
and \U$2929 ( \11748 , \11577 , \11663 , \11747 );
nand \U$2930 ( \11749 , \11029 , \11405 , \11748 );
not \U$2931 ( \11750 , \11749 );
not \U$2932 ( \11751 , \11750 );
xor \U$2933 ( \11752 , \10928 , \10922 );
not \U$2934 ( \11753 , \11752 );
not \U$2935 ( \11754 , \10928 );
not \U$2936 ( \11755 , \10922 );
or \U$2937 ( \11756 , \11754 , \11755 );
xor \U$2938 ( \11757 , RIe548ff0_6844, \11756 );
not \U$2939 ( \11758 , \11757 );
or \U$2940 ( \11759 , \11753 , \11758 );
not \U$2941 ( \11760 , \11759 );
not \U$2942 ( \11761 , \11760 );
or \U$2943 ( \11762 , \10949 , \11761 );
or \U$2944 ( \11763 , \9492 , \11762 );
not \U$2945 ( \11764 , \11760 );
or \U$2946 ( \11765 , \10958 , \11764 );
not \U$2947 ( \11766 , \11765 );
not \U$2948 ( \11767 , \11766 );
or \U$2949 ( \11768 , \9494 , \11767 );
nand \U$2950 ( \11769 , \11763 , \11768 );
not \U$2951 ( \11770 , \11757 );
or \U$2952 ( \11771 , \11752 , \11770 );
not \U$2953 ( \11772 , \11771 );
not \U$2954 ( \11773 , \11772 );
or \U$2955 ( \11774 , \10925 , \11773 );
or \U$2956 ( \11775 , \9498 , \11774 );
not \U$2957 ( \11776 , \11772 );
or \U$2958 ( \11777 , \10939 , \11776 );
or \U$2959 ( \11778 , \9500 , \11777 );
nand \U$2960 ( \11779 , \11775 , \11778 );
nor \U$2961 ( \11780 , \11769 , \11779 );
not \U$2962 ( \11781 , \11757 );
not \U$2963 ( \11782 , \11781 );
or \U$2964 ( \11783 , \11753 , \11782 );
not \U$2965 ( \11784 , \11783 );
not \U$2966 ( \11785 , \11784 );
or \U$2967 ( \11786 , \10925 , \11785 );
not \U$2968 ( \11787 , \11786 );
not \U$2969 ( \11788 , \11787 );
or \U$2970 ( \11789 , \9504 , \11788 );
not \U$2971 ( \11790 , \11772 );
or \U$2972 ( \11791 , \10958 , \11790 );
or \U$2973 ( \11792 , \9506 , \11791 );
nand \U$2974 ( \11793 , \11789 , \11792 );
not \U$2975 ( \11794 , \11781 );
or \U$2976 ( \11795 , \11752 , \11794 );
not \U$2977 ( \11796 , \11795 );
not \U$2978 ( \11797 , \11796 );
or \U$2979 ( \11798 , \10949 , \11797 );
not \U$2980 ( \11799 , \11798 );
not \U$2981 ( \11800 , \11799 );
or \U$2982 ( \11801 , \9509 , \11800 );
not \U$2983 ( \11802 , \11796 );
or \U$2984 ( \11803 , \10939 , \11802 );
not \U$2985 ( \11804 , \11803 );
not \U$2986 ( \11805 , \11804 );
or \U$2987 ( \11806 , \9511 , \11805 );
nand \U$2988 ( \11807 , \11801 , \11806 );
nor \U$2989 ( \11808 , \11793 , \11807 );
not \U$2990 ( \11809 , \9487 );
not \U$2991 ( \11810 , \11760 );
or \U$2992 ( \11811 , \10939 , \11810 );
not \U$2993 ( \11812 , \11811 );
not \U$2994 ( \11813 , \11812 );
not \U$2995 ( \11814 , \11813 );
and \U$2996 ( \11815 , \11809 , \11814 );
not \U$2997 ( \11816 , \11760 );
or \U$2998 ( \11817 , \10925 , \11816 );
not \U$2999 ( \11818 , \11817 );
and \U$3000 ( \11819 , \11818 , \10168 );
nor \U$3001 ( \11820 , \11815 , \11819 );
not \U$3002 ( \11821 , \9482 );
not \U$3003 ( \11822 , \11784 );
or \U$3004 ( \11823 , \10939 , \11822 );
not \U$3005 ( \11824 , \11823 );
not \U$3006 ( \11825 , \11824 );
not \U$3007 ( \11826 , \11825 );
and \U$3008 ( \11827 , \11821 , \11826 );
not \U$3009 ( \11828 , \11772 );
or \U$3010 ( \11829 , \10949 , \11828 );
not \U$3011 ( \11830 , \11829 );
not \U$3012 ( \11831 , \11830 );
not \U$3013 ( \11832 , \11831 );
and \U$3014 ( \11833 , \11832 , \10152 );
nor \U$3015 ( \11834 , \11827 , \11833 );
nand \U$3016 ( \11835 , \11820 , \11834 );
not \U$3017 ( \11836 , \11835 );
not \U$3018 ( \11837 , \9471 );
not \U$3019 ( \11838 , \11784 );
or \U$3020 ( \11839 , \11838 , \10949 );
not \U$3021 ( \11840 , \11839 );
and \U$3022 ( \11841 , \11837 , \11840 );
not \U$3023 ( \11842 , \11784 );
or \U$3024 ( \11843 , \10958 , \11842 );
not \U$3025 ( \11844 , \11843 );
not \U$3026 ( \11845 , \11844 );
not \U$3027 ( \11846 , \11845 );
and \U$3028 ( \11847 , \11846 , \9476 );
nor \U$3029 ( \11848 , \11841 , \11847 );
not \U$3030 ( \11849 , \9463 );
not \U$3031 ( \11850 , \11796 );
or \U$3032 ( \11851 , \11850 , \10958 );
not \U$3033 ( \11852 , \11851 );
and \U$3034 ( \11853 , \11849 , \11852 );
not \U$3035 ( \11854 , \11796 );
or \U$3036 ( \11855 , \11854 , \10925 );
not \U$3037 ( \11856 , \11855 );
and \U$3038 ( \11857 , \11856 , \9468 );
nor \U$3039 ( \11858 , \11853 , \11857 );
and \U$3040 ( \11859 , \11836 , \11848 , \11858 );
nand \U$3041 ( \11860 , \11780 , \11808 , \11859 );
not \U$3042 ( \11861 , \11860 );
not \U$3043 ( \11862 , \9732 );
not \U$3044 ( \11863 , \11799 );
not \U$3045 ( \11864 , \11863 );
and \U$3046 ( \11865 , \11862 , \11864 );
and \U$3047 ( \11866 , \11814 , \9728 );
nor \U$3048 ( \11867 , \11865 , \11866 );
not \U$3049 ( \11868 , \9725 );
not \U$3050 ( \11869 , \11765 );
and \U$3051 ( \11870 , \11868 , \11869 );
and \U$3052 ( \11871 , \11818 , \9721 );
nor \U$3053 ( \11872 , \11870 , \11871 );
not \U$3054 ( \11873 , \11796 );
or \U$3055 ( \11874 , \10925 , \11873 );
or \U$3056 ( \11875 , \9740 , \11874 );
not \U$3057 ( \11876 , \9736 );
not \U$3058 ( \11877 , \11796 );
or \U$3059 ( \11878 , \10958 , \11877 );
or \U$3060 ( \11879 , \11876 , \11878 );
nand \U$3061 ( \11880 , \11875 , \11879 );
not \U$3062 ( \11881 , \11784 );
or \U$3063 ( \11882 , \10949 , \11881 );
or \U$3064 ( \11883 , \9745 , \11882 );
not \U$3065 ( \11884 , \11804 );
or \U$3066 ( \11885 , \9748 , \11884 );
nand \U$3067 ( \11886 , \11883 , \11885 );
nor \U$3068 ( \11887 , \11880 , \11886 );
nand \U$3069 ( \11888 , \11867 , \11872 , \11887 );
not \U$3070 ( \11889 , \11195 );
not \U$3071 ( \11890 , \11777 );
and \U$3072 ( \11891 , \11889 , \11890 );
not \U$3073 ( \11892 , \11762 );
and \U$3074 ( \11893 , \11892 , \9752 );
nor \U$3075 ( \11894 , \11891 , \11893 );
not \U$3076 ( \11895 , \10197 );
not \U$3077 ( \11896 , \11791 );
and \U$3078 ( \11897 , \11895 , \11896 );
not \U$3079 ( \11898 , \11774 );
and \U$3080 ( \11899 , \11898 , \9763 );
nor \U$3081 ( \11900 , \11897 , \11899 );
not \U$3082 ( \11901 , \11787 );
or \U$3083 ( \11902 , \10178 , \11901 );
not \U$3084 ( \11903 , \11844 );
or \U$3085 ( \11904 , \10182 , \11903 );
nand \U$3086 ( \11905 , \11902 , \11904 );
or \U$3087 ( \11906 , \10188 , \11831 );
not \U$3088 ( \11907 , \11824 );
or \U$3089 ( \11908 , \11186 , \11907 );
nand \U$3090 ( \11909 , \11906 , \11908 );
nor \U$3091 ( \11910 , \11905 , \11909 );
nand \U$3092 ( \11911 , \11894 , \11900 , \11910 );
nor \U$3093 ( \11912 , \11888 , \11911 );
xnor \U$3094 ( \11913 , \11912 , \9786 );
not \U$3095 ( \11914 , \9668 );
and \U$3096 ( \11915 , \11914 , \11864 );
and \U$3097 ( \11916 , \11814 , \9664 );
nor \U$3098 ( \11917 , \11915 , \11916 );
not \U$3099 ( \11918 , \9661 );
and \U$3100 ( \11919 , \11918 , \11869 );
and \U$3101 ( \11920 , \11818 , \9656 );
nor \U$3102 ( \11921 , \11919 , \11920 );
or \U$3103 ( \11922 , \9676 , \11855 );
not \U$3104 ( \11923 , \9672 );
or \U$3105 ( \11924 , \11923 , \11851 );
nand \U$3106 ( \11925 , \11922 , \11924 );
or \U$3107 ( \11926 , \9680 , \11839 );
or \U$3108 ( \11927 , \9683 , \11805 );
nand \U$3109 ( \11928 , \11926 , \11927 );
nor \U$3110 ( \11929 , \11925 , \11928 );
nand \U$3111 ( \11930 , \11917 , \11921 , \11929 );
and \U$3112 ( \11931 , \11892 , \9687 );
and \U$3113 ( \11932 , \9690 , \11890 );
nor \U$3114 ( \11933 , \11931 , \11932 );
not \U$3115 ( \11934 , \11774 );
and \U$3116 ( \11935 , \11934 , \9695 );
not \U$3117 ( \11936 , \11791 );
and \U$3118 ( \11937 , \9692 , \11936 );
nor \U$3119 ( \11938 , \11935 , \11937 );
or \U$3120 ( \11939 , \11138 , \11901 );
or \U$3121 ( \11940 , \11140 , \11845 );
nand \U$3122 ( \11941 , \11939 , \11940 );
or \U$3123 ( \11942 , \10244 , \11831 );
or \U$3124 ( \11943 , \11145 , \11907 );
nand \U$3125 ( \11944 , \11942 , \11943 );
nor \U$3126 ( \11945 , \11941 , \11944 );
nand \U$3127 ( \11946 , \11933 , \11938 , \11945 );
nor \U$3128 ( \11947 , \11930 , \11946 );
xnor \U$3129 ( \11948 , \11947 , \9719 );
or \U$3130 ( \11949 , \11088 , \11825 );
not \U$3131 ( \11950 , \11830 );
or \U$3132 ( \11951 , \10323 , \11950 );
nand \U$3133 ( \11952 , \11949 , \11951 );
or \U$3134 ( \11953 , \11125 , \11845 );
not \U$3135 ( \11954 , \9200 );
or \U$3136 ( \11955 , \11954 , \11901 );
nand \U$3137 ( \11956 , \11953 , \11955 );
nor \U$3138 ( \11957 , \11952 , \11956 );
not \U$3139 ( \11958 , \11796 );
or \U$3140 ( \11959 , \10925 , \11958 );
or \U$3141 ( \11960 , \11098 , \11959 );
not \U$3142 ( \11961 , \11796 );
or \U$3143 ( \11962 , \10958 , \11961 );
or \U$3144 ( \11963 , \11101 , \11962 );
nand \U$3145 ( \11964 , \11960 , \11963 );
not \U$3146 ( \11965 , \11784 );
or \U$3147 ( \11966 , \10949 , \11965 );
or \U$3148 ( \11967 , \9217 , \11966 );
or \U$3149 ( \11968 , \9220 , \11884 );
nand \U$3150 ( \11969 , \11967 , \11968 );
nor \U$3151 ( \11970 , \11964 , \11969 );
and \U$3152 ( \11971 , \11869 , \9225 );
and \U$3153 ( \11972 , \9204 , \11818 );
nor \U$3154 ( \11973 , \11971 , \11972 );
and \U$3155 ( \11974 , \11814 , \9196 );
and \U$3156 ( \11975 , \9239 , \11864 );
nor \U$3157 ( \11976 , \11974 , \11975 );
nand \U$3158 ( \11977 , \11973 , \11976 );
not \U$3159 ( \11978 , \11977 );
not \U$3160 ( \11979 , \11777 );
and \U$3161 ( \11980 , \11979 , \9233 );
and \U$3162 ( \11981 , \9230 , \11892 );
nor \U$3163 ( \11982 , \11980 , \11981 );
and \U$3164 ( \11983 , \11934 , \9251 );
and \U$3165 ( \11984 , \9247 , \11936 );
nor \U$3166 ( \11985 , \11983 , \11984 );
and \U$3167 ( \11986 , \11978 , \11982 , \11985 );
nand \U$3168 ( \11987 , \11957 , \11970 , \11986 );
xnor \U$3169 ( \11988 , \11987 , \9260 );
or \U$3170 ( \11989 , \8971 , \11907 );
or \U$3171 ( \11990 , \10370 , \11950 );
nand \U$3172 ( \11991 , \11989 , \11990 );
or \U$3173 ( \11992 , \11073 , \11903 );
or \U$3174 ( \11993 , \8980 , \11788 );
nand \U$3175 ( \11994 , \11992 , \11993 );
nor \U$3176 ( \11995 , \11991 , \11994 );
or \U$3177 ( \11996 , \8991 , \11855 );
or \U$3178 ( \11997 , \11046 , \11851 );
nand \U$3179 ( \11998 , \11996 , \11997 );
or \U$3180 ( \11999 , \8997 , \11839 );
or \U$3181 ( \12000 , \9000 , \11805 );
nand \U$3182 ( \12001 , \11999 , \12000 );
nor \U$3183 ( \12002 , \11998 , \12001 );
and \U$3184 ( \12003 , \11869 , \9006 );
and \U$3185 ( \12004 , \8976 , \11818 );
nor \U$3186 ( \12005 , \12003 , \12004 );
and \U$3187 ( \12006 , \11814 , \8966 );
and \U$3188 ( \12007 , \9020 , \11864 );
nor \U$3189 ( \12008 , \12006 , \12007 );
nand \U$3190 ( \12009 , \12005 , \12008 );
not \U$3191 ( \12010 , \12009 );
and \U$3192 ( \12011 , \11979 , \9014 );
and \U$3193 ( \12012 , \9011 , \11892 );
nor \U$3194 ( \12013 , \12011 , \12012 );
and \U$3195 ( \12014 , \11898 , \9034 );
and \U$3196 ( \12015 , \9030 , \11896 );
nor \U$3197 ( \12016 , \12014 , \12015 );
and \U$3198 ( \12017 , \12010 , \12013 , \12016 );
nand \U$3199 ( \12018 , \11995 , \12002 , \12017 );
xnor \U$3200 ( \12019 , \12018 , \9044 );
nor \U$3201 ( \12020 , \11988 , \12019 );
nand \U$3202 ( \12021 , \11913 , \11948 , \12020 );
not \U$3203 ( \12022 , \12021 );
or \U$3204 ( \12023 , \9266 , \11825 );
or \U$3205 ( \12024 , \10415 , \11831 );
nand \U$3206 ( \12025 , \12023 , \12024 );
or \U$3207 ( \12026 , \11298 , \11903 );
or \U$3208 ( \12027 , \9273 , \11788 );
nand \U$3209 ( \12028 , \12026 , \12027 );
nor \U$3210 ( \12029 , \12025 , \12028 );
or \U$3211 ( \12030 , \9282 , \11874 );
or \U$3212 ( \12031 , \11276 , \11878 );
nand \U$3213 ( \12032 , \12030 , \12031 );
or \U$3214 ( \12033 , \9287 , \11882 );
or \U$3215 ( \12034 , \9290 , \11805 );
nand \U$3216 ( \12035 , \12033 , \12034 );
nor \U$3217 ( \12036 , \12032 , \12035 );
not \U$3218 ( \12037 , \9270 );
and \U$3219 ( \12038 , \12037 , \11818 );
and \U$3220 ( \12039 , \11869 , \9295 );
nor \U$3221 ( \12040 , \12038 , \12039 );
not \U$3222 ( \12041 , \11270 );
and \U$3223 ( \12042 , \12041 , \11864 );
and \U$3224 ( \12043 , \11814 , \9262 );
nor \U$3225 ( \12044 , \12042 , \12043 );
nand \U$3226 ( \12045 , \12040 , \12044 );
not \U$3227 ( \12046 , \12045 );
not \U$3228 ( \12047 , \11288 );
and \U$3229 ( \12048 , \12047 , \11892 );
and \U$3230 ( \12049 , \11979 , \9302 );
nor \U$3231 ( \12050 , \12048 , \12049 );
not \U$3232 ( \12051 , \11293 );
and \U$3233 ( \12052 , \12051 , \11896 );
and \U$3234 ( \12053 , \11898 , \9319 );
nor \U$3235 ( \12054 , \12052 , \12053 );
and \U$3236 ( \12055 , \12046 , \12050 , \12054 );
nand \U$3237 ( \12056 , \12029 , \12036 , \12055 );
xnor \U$3238 ( \12057 , \12056 , \9327 );
or \U$3239 ( \12058 , \9398 , \11825 );
or \U$3240 ( \12059 , \10462 , \11831 );
nand \U$3241 ( \12060 , \12058 , \12059 );
or \U$3242 ( \12061 , \10464 , \11903 );
or \U$3243 ( \12062 , \9405 , \11788 );
nand \U$3244 ( \12063 , \12061 , \12062 );
nor \U$3245 ( \12064 , \12060 , \12063 );
or \U$3246 ( \12065 , \9415 , \11959 );
or \U$3247 ( \12066 , \10455 , \11962 );
nand \U$3248 ( \12067 , \12065 , \12066 );
or \U$3249 ( \12068 , \9419 , \11966 );
or \U$3250 ( \12069 , \9422 , \11805 );
nand \U$3251 ( \12070 , \12068 , \12069 );
nor \U$3252 ( \12071 , \12067 , \12070 );
not \U$3253 ( \12072 , \9402 );
and \U$3254 ( \12073 , \12072 , \11818 );
and \U$3255 ( \12074 , \11869 , \9427 );
nor \U$3256 ( \12075 , \12073 , \12074 );
not \U$3257 ( \12076 , \11230 );
and \U$3258 ( \12077 , \12076 , \11864 );
and \U$3259 ( \12078 , \11814 , \9394 );
nor \U$3260 ( \12079 , \12077 , \12078 );
nand \U$3261 ( \12080 , \12075 , \12079 );
not \U$3262 ( \12081 , \12080 );
not \U$3263 ( \12082 , \11245 );
and \U$3264 ( \12083 , \12082 , \11892 );
and \U$3265 ( \12084 , \11979 , \9435 );
nor \U$3266 ( \12085 , \12083 , \12084 );
not \U$3267 ( \12086 , \11250 );
and \U$3268 ( \12087 , \12086 , \11896 );
and \U$3269 ( \12088 , \11898 , \9453 );
nor \U$3270 ( \12089 , \12087 , \12088 );
and \U$3271 ( \12090 , \12081 , \12085 , \12089 );
nand \U$3272 ( \12091 , \12064 , \12071 , \12090 );
xnor \U$3273 ( \12092 , \12091 , \9460 );
nor \U$3274 ( \12093 , \12057 , \12092 );
or \U$3275 ( \12094 , \9620 , \11774 );
or \U$3276 ( \12095 , \9625 , \11791 );
nand \U$3277 ( \12096 , \12094 , \12095 );
or \U$3278 ( \12097 , \9632 , \11762 );
or \U$3279 ( \12098 , \11314 , \11777 );
nand \U$3280 ( \12099 , \12097 , \12098 );
nor \U$3281 ( \12100 , \12096 , \12099 );
or \U$3282 ( \12101 , \9637 , \11817 );
or \U$3283 ( \12102 , \9640 , \11767 );
nand \U$3284 ( \12103 , \12101 , \12102 );
or \U$3285 ( \12104 , \9647 , \11800 );
or \U$3286 ( \12105 , \11322 , \11813 );
nand \U$3287 ( \12106 , \12104 , \12105 );
nor \U$3288 ( \12107 , \12103 , \12106 );
not \U$3289 ( \12108 , \9593 );
not \U$3290 ( \12109 , \12108 );
not \U$3291 ( \12110 , \11884 );
and \U$3292 ( \12111 , \12109 , \12110 );
and \U$3293 ( \12112 , \11840 , \9587 );
nor \U$3294 ( \12113 , \12111 , \12112 );
not \U$3295 ( \12114 , \9597 );
and \U$3296 ( \12115 , \12114 , \11852 );
and \U$3297 ( \12116 , \11856 , \9600 );
nor \U$3298 ( \12117 , \12115 , \12116 );
nand \U$3299 ( \12118 , \12113 , \12117 );
not \U$3300 ( \12119 , \12118 );
not \U$3301 ( \12120 , \9607 );
and \U$3302 ( \12121 , \12120 , \11846 );
not \U$3303 ( \12122 , \11901 );
and \U$3304 ( \12123 , \12122 , \9603 );
nor \U$3305 ( \12124 , \12121 , \12123 );
not \U$3306 ( \12125 , \9614 );
and \U$3307 ( \12126 , \12125 , \11826 );
and \U$3308 ( \12127 , \11832 , \9610 );
nor \U$3309 ( \12128 , \12126 , \12127 );
and \U$3310 ( \12129 , \12119 , \12124 , \12128 );
nand \U$3311 ( \12130 , \12100 , \12107 , \12129 );
xnor \U$3312 ( \12131 , \12130 , \9653 );
or \U$3313 ( \12132 , \9335 , \11825 );
or \U$3314 ( \12133 , \10553 , \11831 );
nand \U$3315 ( \12134 , \12132 , \12133 );
or \U$3316 ( \12135 , \11357 , \11845 );
or \U$3317 ( \12136 , \9342 , \11788 );
nand \U$3318 ( \12137 , \12135 , \12136 );
nor \U$3319 ( \12138 , \12134 , \12137 );
not \U$3320 ( \12139 , \9348 );
or \U$3321 ( \12140 , \12139 , \11855 );
not \U$3322 ( \12141 , \9346 );
or \U$3323 ( \12142 , \12141 , \11851 );
nand \U$3324 ( \12143 , \12140 , \12142 );
or \U$3325 ( \12144 , \9354 , \11839 );
or \U$3326 ( \12145 , \9357 , \11805 );
nand \U$3327 ( \12146 , \12144 , \12145 );
nor \U$3328 ( \12147 , \12143 , \12146 );
not \U$3329 ( \12148 , \9339 );
and \U$3330 ( \12149 , \12148 , \11818 );
and \U$3331 ( \12150 , \11869 , \9361 );
nor \U$3332 ( \12151 , \12149 , \12150 );
not \U$3333 ( \12152 , \11393 );
and \U$3334 ( \12153 , \12152 , \11864 );
and \U$3335 ( \12154 , \11814 , \9331 );
nor \U$3336 ( \12155 , \12153 , \12154 );
nand \U$3337 ( \12156 , \12151 , \12155 );
not \U$3338 ( \12157 , \12156 );
not \U$3339 ( \12158 , \11365 );
and \U$3340 ( \12159 , \12158 , \11892 );
and \U$3341 ( \12160 , \11979 , \9369 );
nor \U$3342 ( \12161 , \12159 , \12160 );
not \U$3343 ( \12162 , \11371 );
and \U$3344 ( \12163 , \12162 , \11934 );
and \U$3345 ( \12164 , \11896 , \9385 );
nor \U$3346 ( \12165 , \12163 , \12164 );
and \U$3347 ( \12166 , \12157 , \12161 , \12165 );
nand \U$3348 ( \12167 , \12138 , \12147 , \12166 );
xnor \U$3349 ( \12168 , \12167 , \9392 );
nor \U$3350 ( \12169 , \12131 , \12168 );
and \U$3351 ( \12170 , \12022 , \12093 , \12169 );
not \U$3352 ( \12171 , \9887 );
and \U$3353 ( \12172 , \12171 , \11826 );
and \U$3354 ( \12173 , \11832 , \9881 );
nor \U$3355 ( \12174 , \12172 , \12173 );
and \U$3356 ( \12175 , \12122 , \9874 );
and \U$3357 ( \12176 , \9877 , \11846 );
nor \U$3358 ( \12177 , \12175 , \12176 );
not \U$3359 ( \12178 , \9871 );
or \U$3360 ( \12179 , \12178 , \11959 );
or \U$3361 ( \12180 , \9868 , \11962 );
nand \U$3362 ( \12181 , \12179 , \12180 );
or \U$3363 ( \12182 , \9860 , \11966 );
not \U$3364 ( \12183 , \9864 );
or \U$3365 ( \12184 , \12183 , \11805 );
nand \U$3366 ( \12185 , \12182 , \12184 );
nor \U$3367 ( \12186 , \12181 , \12185 );
nand \U$3368 ( \12187 , \12174 , \12177 , \12186 );
not \U$3369 ( \12188 , \12187 );
or \U$3370 ( \12189 , \9911 , \11817 );
or \U$3371 ( \12190 , \9914 , \11767 );
nand \U$3372 ( \12191 , \12189 , \12190 );
or \U$3373 ( \12192 , \9921 , \11800 );
not \U$3374 ( \12193 , \11812 );
or \U$3375 ( \12194 , \11718 , \12193 );
nand \U$3376 ( \12195 , \12192 , \12194 );
nor \U$3377 ( \12196 , \12191 , \12195 );
or \U$3378 ( \12197 , \9895 , \11774 );
or \U$3379 ( \12198 , \9898 , \11791 );
nand \U$3380 ( \12199 , \12197 , \12198 );
or \U$3381 ( \12200 , \9906 , \11762 );
or \U$3382 ( \12201 , \11711 , \11777 );
nand \U$3383 ( \12202 , \12200 , \12201 );
nor \U$3384 ( \12203 , \12199 , \12202 );
and \U$3385 ( \12204 , \12188 , \12196 , \12203 );
xnor \U$3386 ( \12205 , \12204 , \9927 );
and \U$3387 ( \12206 , \11832 , \10017 );
and \U$3388 ( \12207 , \10020 , \11826 );
nor \U$3389 ( \12208 , \12206 , \12207 );
and \U$3390 ( \12209 , \12122 , \10009 );
and \U$3391 ( \12210 , \10012 , \11846 );
nor \U$3392 ( \12211 , \12209 , \12210 );
or \U$3393 ( \12212 , \9997 , \11874 );
or \U$3394 ( \12213 , \11666 , \11878 );
nand \U$3395 ( \12214 , \12212 , \12213 );
or \U$3396 ( \12215 , \10002 , \11882 );
or \U$3397 ( \12216 , \10005 , \11805 );
nand \U$3398 ( \12217 , \12215 , \12216 );
nor \U$3399 ( \12218 , \12214 , \12217 );
nand \U$3400 ( \12219 , \12208 , \12211 , \12218 );
not \U$3401 ( \12220 , \12219 );
or \U$3402 ( \12221 , \11684 , \11817 );
not \U$3403 ( \12222 , \10041 );
or \U$3404 ( \12223 , \12222 , \11767 );
nand \U$3405 ( \12224 , \12221 , \12223 );
or \U$3406 ( \12225 , \11674 , \11800 );
or \U$3407 ( \12226 , \11681 , \12193 );
nand \U$3408 ( \12227 , \12225 , \12226 );
nor \U$3409 ( \12228 , \12224 , \12227 );
not \U$3410 ( \12229 , \10035 );
buf \U$3411 ( \12230 , \12229 );
or \U$3412 ( \12231 , \12230 , \11774 );
or \U$3413 ( \12232 , \11698 , \11791 );
nand \U$3414 ( \12233 , \12231 , \12232 );
or \U$3415 ( \12234 , \11693 , \11762 );
not \U$3416 ( \12235 , \10027 );
or \U$3417 ( \12236 , \12235 , \11777 );
nand \U$3418 ( \12237 , \12234 , \12236 );
nor \U$3419 ( \12238 , \12233 , \12237 );
and \U$3420 ( \12239 , \12220 , \12228 , \12238 );
xnor \U$3421 ( \12240 , \12239 , \10055 );
or \U$3422 ( \12241 , \9552 , \11774 );
or \U$3423 ( \12242 , \9557 , \11791 );
nand \U$3424 ( \12243 , \12241 , \12242 );
or \U$3425 ( \12244 , \9564 , \11762 );
or \U$3426 ( \12245 , \11582 , \11777 );
nand \U$3427 ( \12246 , \12244 , \12245 );
nor \U$3428 ( \12247 , \12243 , \12246 );
or \U$3429 ( \12248 , \9569 , \11817 );
or \U$3430 ( \12249 , \9572 , \11767 );
nand \U$3431 ( \12250 , \12248 , \12249 );
or \U$3432 ( \12251 , \9579 , \11800 );
or \U$3433 ( \12252 , \11589 , \12193 );
nand \U$3434 ( \12253 , \12251 , \12252 );
nor \U$3435 ( \12254 , \12250 , \12253 );
and \U$3436 ( \12255 , \11840 , \9518 );
and \U$3437 ( \12256 , \9522 , \12110 );
nor \U$3438 ( \12257 , \12255 , \12256 );
and \U$3439 ( \12258 , \11856 , \9530 );
and \U$3440 ( \12259 , \9526 , \11852 );
nor \U$3441 ( \12260 , \12258 , \12259 );
nand \U$3442 ( \12261 , \12257 , \12260 );
not \U$3443 ( \12262 , \12261 );
and \U$3444 ( \12263 , \12122 , \9533 );
and \U$3445 ( \12264 , \9536 , \11846 );
nor \U$3446 ( \12265 , \12263 , \12264 );
and \U$3447 ( \12266 , \11832 , \9542 );
and \U$3448 ( \12267 , \9545 , \11826 );
nor \U$3449 ( \12268 , \12266 , \12267 );
and \U$3450 ( \12269 , \12262 , \12265 , \12268 );
nand \U$3451 ( \12270 , \12247 , \12254 , \12269 );
xnor \U$3452 ( \12271 , \12270 , \9585 );
or \U$3453 ( \12272 , \11618 , \11774 );
or \U$3454 ( \12273 , \11620 , \11791 );
nand \U$3455 ( \12274 , \12272 , \12273 );
or \U$3456 ( \12275 , \11623 , \11762 );
or \U$3457 ( \12276 , \11625 , \11777 );
nand \U$3458 ( \12277 , \12275 , \12276 );
nor \U$3459 ( \12278 , \12274 , \12277 );
or \U$3460 ( \12279 , \11635 , \11817 );
or \U$3461 ( \12280 , \11629 , \11767 );
nand \U$3462 ( \12281 , \12279 , \12280 );
not \U$3463 ( \12282 , \9984 );
or \U$3464 ( \12283 , \12282 , \11800 );
or \U$3465 ( \12284 , \11633 , \11813 );
nand \U$3466 ( \12285 , \12283 , \12284 );
nor \U$3467 ( \12286 , \12281 , \12285 );
and \U$3468 ( \12287 , \11840 , \9951 );
and \U$3469 ( \12288 , \9954 , \12110 );
nor \U$3470 ( \12289 , \12287 , \12288 );
and \U$3471 ( \12290 , \11856 , \9947 );
and \U$3472 ( \12291 , \9944 , \11852 );
nor \U$3473 ( \12292 , \12290 , \12291 );
nand \U$3474 ( \12293 , \12289 , \12292 );
not \U$3475 ( \12294 , \12293 );
and \U$3476 ( \12295 , \12122 , \9929 );
and \U$3477 ( \12296 , \9932 , \11846 );
nor \U$3478 ( \12297 , \12295 , \12296 );
and \U$3479 ( \12298 , \11832 , \9936 );
and \U$3480 ( \12299 , \9939 , \11826 );
nor \U$3481 ( \12300 , \12298 , \12299 );
and \U$3482 ( \12301 , \12294 , \12297 , \12300 );
nand \U$3483 ( \12302 , \12278 , \12286 , \12301 );
xnor \U$3484 ( \12303 , \12302 , \9990 );
nor \U$3485 ( \12304 , \12271 , \12303 );
nand \U$3486 ( \12305 , \12205 , \12240 , \12304 );
not \U$3487 ( \12306 , \12305 );
or \U$3488 ( \12307 , \9823 , \11774 );
or \U$3489 ( \12308 , \9827 , \11791 );
nand \U$3490 ( \12309 , \12307 , \12308 );
or \U$3491 ( \12310 , \9834 , \11762 );
not \U$3492 ( \12311 , \9830 );
or \U$3493 ( \12312 , \12311 , \11777 );
nand \U$3494 ( \12313 , \12310 , \12312 );
nor \U$3495 ( \12314 , \12309 , \12313 );
or \U$3496 ( \12315 , \9840 , \11817 );
or \U$3497 ( \12316 , \9843 , \11767 );
nand \U$3498 ( \12317 , \12315 , \12316 );
or \U$3499 ( \12318 , \9851 , \11800 );
or \U$3500 ( \12319 , \11505 , \11813 );
nand \U$3501 ( \12320 , \12318 , \12319 );
nor \U$3502 ( \12321 , \12317 , \12320 );
not \U$3503 ( \12322 , \11492 );
and \U$3504 ( \12323 , \12322 , \12110 );
and \U$3505 ( \12324 , \11840 , \9790 );
nor \U$3506 ( \12325 , \12323 , \12324 );
not \U$3507 ( \12326 , \9798 );
and \U$3508 ( \12327 , \12326 , \11852 );
and \U$3509 ( \12328 , \11856 , \9801 );
nor \U$3510 ( \12329 , \12327 , \12328 );
nand \U$3511 ( \12330 , \12325 , \12329 );
not \U$3512 ( \12331 , \12330 );
not \U$3513 ( \12332 , \9809 );
and \U$3514 ( \12333 , \12332 , \11846 );
and \U$3515 ( \12334 , \12122 , \9805 );
nor \U$3516 ( \12335 , \12333 , \12334 );
not \U$3517 ( \12336 , \9817 );
and \U$3518 ( \12337 , \12336 , \11826 );
and \U$3519 ( \12338 , \11832 , \9813 );
nor \U$3520 ( \12339 , \12337 , \12338 );
and \U$3521 ( \12340 , \12331 , \12335 , \12339 );
nand \U$3522 ( \12341 , \12314 , \12321 , \12340 );
xnor \U$3523 ( \12342 , \12341 , \9857 );
or \U$3524 ( \12343 , \8844 , \11825 );
or \U$3525 ( \12344 , \10775 , \11950 );
nand \U$3526 ( \12345 , \12343 , \12344 );
or \U$3527 ( \12346 , \11533 , \11845 );
or \U$3528 ( \12347 , \8861 , \11901 );
nand \U$3529 ( \12348 , \12346 , \12347 );
nor \U$3530 ( \12349 , \12345 , \12348 );
or \U$3531 ( \12350 , \8882 , \11855 );
not \U$3532 ( \12351 , \8868 );
or \U$3533 ( \12352 , \12351 , \11851 );
nand \U$3534 ( \12353 , \12350 , \12352 );
or \U$3535 ( \12354 , \8894 , \11839 );
or \U$3536 ( \12355 , \8897 , \11805 );
nand \U$3537 ( \12356 , \12354 , \12355 );
nor \U$3538 ( \12357 , \12353 , \12356 );
not \U$3539 ( \12358 , \8853 );
and \U$3540 ( \12359 , \12358 , \11818 );
and \U$3541 ( \12360 , \11869 , \8904 );
nor \U$3542 ( \12361 , \12359 , \12360 );
not \U$3543 ( \12362 , \11565 );
and \U$3544 ( \12363 , \12362 , \11864 );
and \U$3545 ( \12364 , \11814 , \8827 );
nor \U$3546 ( \12365 , \12363 , \12364 );
nand \U$3547 ( \12366 , \12361 , \12365 );
not \U$3548 ( \12367 , \12366 );
not \U$3549 ( \12368 , \11540 );
and \U$3550 ( \12369 , \12368 , \11892 );
and \U$3551 ( \12370 , \11979 , \8927 );
nor \U$3552 ( \12371 , \12369 , \12370 );
not \U$3553 ( \12372 , \11545 );
and \U$3554 ( \12373 , \12372 , \11936 );
and \U$3555 ( \12374 , \11934 , \8953 );
nor \U$3556 ( \12375 , \12373 , \12374 );
and \U$3557 ( \12376 , \12367 , \12371 , \12375 );
nand \U$3558 ( \12377 , \12349 , \12357 , \12376 );
xnor \U$3559 ( \12378 , \12377 , \8964 );
nor \U$3560 ( \12379 , \12342 , \12378 );
or \U$3561 ( \12380 , \9050 , \11825 );
or \U$3562 ( \12381 , \10859 , \11831 );
nand \U$3563 ( \12382 , \12380 , \12381 );
or \U$3564 ( \12383 , \9086 , \11903 );
or \U$3565 ( \12384 , \9058 , \11901 );
nand \U$3566 ( \12385 , \12383 , \12384 );
nor \U$3567 ( \12386 , \12382 , \12385 );
or \U$3568 ( \12387 , \9068 , \11874 );
or \U$3569 ( \12388 , \11458 , \11878 );
nand \U$3570 ( \12389 , \12387 , \12388 );
or \U$3571 ( \12390 , \9073 , \11882 );
or \U$3572 ( \12391 , \9076 , \11805 );
nand \U$3573 ( \12392 , \12390 , \12391 );
nor \U$3574 ( \12393 , \12389 , \12392 );
not \U$3575 ( \12394 , \9055 );
and \U$3576 ( \12395 , \12394 , \11818 );
and \U$3577 ( \12396 , \11869 , \9081 );
nor \U$3578 ( \12397 , \12395 , \12396 );
not \U$3579 ( \12398 , \11452 );
and \U$3580 ( \12399 , \12398 , \11864 );
and \U$3581 ( \12400 , \11814 , \9046 );
nor \U$3582 ( \12401 , \12399 , \12400 );
nand \U$3583 ( \12402 , \12397 , \12401 );
not \U$3584 ( \12403 , \12402 );
and \U$3585 ( \12404 , \11979 , \9093 );
and \U$3586 ( \12405 , \9089 , \11892 );
nor \U$3587 ( \12406 , \12404 , \12405 );
and \U$3588 ( \12407 , \11898 , \9112 );
and \U$3589 ( \12408 , \9107 , \11896 );
nor \U$3590 ( \12409 , \12407 , \12408 );
and \U$3591 ( \12410 , \12403 , \12406 , \12409 );
nand \U$3592 ( \12411 , \12386 , \12393 , \12410 );
xnor \U$3593 ( \12412 , \12411 , \9119 );
or \U$3594 ( \12413 , \9125 , \11825 );
or \U$3595 ( \12414 , \10901 , \11950 );
nand \U$3596 ( \12415 , \12413 , \12414 );
or \U$3597 ( \12416 , \11436 , \11845 );
or \U$3598 ( \12417 , \9133 , \11901 );
nand \U$3599 ( \12418 , \12416 , \12417 );
nor \U$3600 ( \12419 , \12415 , \12418 );
or \U$3601 ( \12420 , \9143 , \11959 );
or \U$3602 ( \12421 , \11416 , \11962 );
nand \U$3603 ( \12422 , \12420 , \12421 );
or \U$3604 ( \12423 , \9148 , \11966 );
or \U$3605 ( \12424 , \9151 , \11805 );
nand \U$3606 ( \12425 , \12423 , \12424 );
nor \U$3607 ( \12426 , \12422 , \12425 );
not \U$3608 ( \12427 , \9130 );
and \U$3609 ( \12428 , \12427 , \11818 );
and \U$3610 ( \12429 , \11869 , \9155 );
nor \U$3611 ( \12430 , \12428 , \12429 );
not \U$3612 ( \12431 , \11410 );
and \U$3613 ( \12432 , \12431 , \11864 );
and \U$3614 ( \12433 , \11814 , \9121 );
nor \U$3615 ( \12434 , \12432 , \12433 );
nand \U$3616 ( \12435 , \12430 , \12434 );
not \U$3617 ( \12436 , \12435 );
not \U$3618 ( \12437 , \11426 );
and \U$3619 ( \12438 , \12437 , \11892 );
and \U$3620 ( \12439 , \11979 , \9163 );
nor \U$3621 ( \12440 , \12438 , \12439 );
and \U$3622 ( \12441 , \11934 , \9180 );
and \U$3623 ( \12442 , \9176 , \11936 );
nor \U$3624 ( \12443 , \12441 , \12442 );
and \U$3625 ( \12444 , \12436 , \12440 , \12443 );
nand \U$3626 ( \12445 , \12419 , \12426 , \12444 );
xnor \U$3627 ( \12446 , \12445 , \9188 );
nor \U$3628 ( \12447 , \12412 , \12446 );
and \U$3629 ( \12448 , \12306 , \12379 , \12447 );
nand \U$3630 ( \12449 , \11861 , \12170 , \12448 );
and \U$3631 ( \12450 , \10916 , \11751 , \12449 );
not \U$3632 ( \12451 , \12450 );
buf \U$3633 ( \12452 , RIea91330_6888);
not \U$3634 ( \12453 , \10065 );
not \U$3635 ( \12454 , \12453 );
buf \U$3636 ( \12455 , \12454 );
not \U$3637 ( \12456 , \8836 );
buf \U$3638 ( \12457 , \12456 );
not \U$3639 ( \12458 , \8829 );
buf \U$3640 ( \12459 , \12458 );
buf \U$3641 ( \12460 , \8835 );
and \U$3642 ( \12461 , \12459 , \12460 );
and \U$3643 ( \12462 , \12457 , \12461 );
or \U$3644 ( \12463 , \12455 , \12462 );
and \U$3645 ( \12464 , \12452 , \12463 );
buf \U$3646 ( \12465 , \12464 );
not \U$3647 ( \12466 , \12460 );
buf \U$3648 ( \12467 , \12466 );
not \U$3649 ( \12468 , \12467 );
xor \U$3650 ( \12469 , \12459 , \12460 );
buf \U$3651 ( \12470 , \12469 );
not \U$3652 ( \12471 , \12470 );
nand \U$3653 ( \12472 , \12468 , \12471 );
xor \U$3654 ( \12473 , \12457 , \12461 );
buf \U$3655 ( \12474 , \12473 );
not \U$3656 ( \12475 , \12474 );
xnor \U$3657 ( \12476 , \12455 , \12462 );
buf \U$3658 ( \12477 , \12476 );
not \U$3659 ( \12478 , \12477 );
nand \U$3660 ( \12479 , \12475 , \12478 );
or \U$3661 ( \12480 , \12472 , \12479 );
xor \U$3662 ( \12481 , \12452 , \12463 );
buf \U$3663 ( \12482 , \12481 );
nand \U$3664 ( \12483 , \12480 , \12482 );
not \U$3665 ( \12484 , \12483 );
or \U$3666 ( \12485 , \12465 , \12484 );
not \U$3667 ( \12486 , \12485 );
not \U$3668 ( \12487 , \9500 );
not \U$3669 ( \12488 , \10097 );
or \U$3670 ( \12489 , \10065 , \12488 );
not \U$3671 ( \12490 , \12489 );
not \U$3672 ( \12491 , \12490 );
not \U$3673 ( \12492 , \10096 );
or \U$3674 ( \12493 , \8906 , \12492 );
nand \U$3675 ( \12494 , \12491 , \12493 );
not \U$3676 ( \12495 , \12494 );
not \U$3677 ( \12496 , \11006 );
or \U$3678 ( \12497 , \12495 , \12496 );
not \U$3679 ( \12498 , \12497 );
and \U$3680 ( \12499 , \12487 , \12498 );
not \U$3681 ( \12500 , \10978 );
or \U$3682 ( \12501 , \12495 , \12500 );
not \U$3683 ( \12502 , \12501 );
and \U$3684 ( \12503 , \12502 , \10085 );
nor \U$3685 ( \12504 , \12499 , \12503 );
not \U$3686 ( \12505 , \9494 );
not \U$3687 ( \12506 , \10968 );
or \U$3688 ( \12507 , \12495 , \12506 );
not \U$3689 ( \12508 , \12507 );
and \U$3690 ( \12509 , \12505 , \12508 );
not \U$3691 ( \12510 , \10972 );
or \U$3692 ( \12511 , \12495 , \12510 );
not \U$3693 ( \12512 , \12511 );
not \U$3694 ( \12513 , \9492 );
and \U$3695 ( \12514 , \12512 , \12513 );
nor \U$3696 ( \12515 , \12509 , \12514 );
nand \U$3697 ( \12516 , \12504 , \12515 );
not \U$3698 ( \12517 , \12516 );
not \U$3699 ( \12518 , \9506 );
not \U$3700 ( \12519 , \10941 );
or \U$3701 ( \12520 , \12495 , \12519 );
not \U$3702 ( \12521 , \12520 );
and \U$3703 ( \12522 , \12518 , \12521 );
not \U$3704 ( \12523 , \10952 );
or \U$3705 ( \12524 , \12494 , \12523 );
not \U$3706 ( \12525 , \12524 );
and \U$3707 ( \12526 , \12525 , \10976 );
nor \U$3708 ( \12527 , \12522 , \12526 );
not \U$3709 ( \12528 , \9509 );
not \U$3710 ( \12529 , \10927 );
or \U$3711 ( \12530 , \12494 , \12529 );
not \U$3712 ( \12531 , \12530 );
and \U$3713 ( \12532 , \12528 , \12531 );
not \U$3714 ( \12533 , \11006 );
or \U$3715 ( \12534 , \12494 , \12533 );
not \U$3716 ( \12535 , \12534 );
and \U$3717 ( \12536 , \12535 , \10120 );
nor \U$3718 ( \12537 , \12532 , \12536 );
and \U$3719 ( \12538 , \12517 , \12527 , \12537 );
not \U$3720 ( \12539 , \9487 );
not \U$3721 ( \12540 , \10960 );
or \U$3722 ( \12541 , \12495 , \12540 );
not \U$3723 ( \12542 , \12541 );
and \U$3724 ( \12543 , \12539 , \12542 );
not \U$3725 ( \12544 , \10952 );
or \U$3726 ( \12545 , \12495 , \12544 );
not \U$3727 ( \12546 , \12545 );
and \U$3728 ( \12547 , \12546 , \10168 );
nor \U$3729 ( \12548 , \12543 , \12547 );
not \U$3730 ( \12549 , \9480 );
not \U$3731 ( \12550 , \10927 );
or \U$3732 ( \12551 , \12495 , \12550 );
not \U$3733 ( \12552 , \12551 );
and \U$3734 ( \12553 , \12549 , \12552 );
not \U$3735 ( \12554 , \10960 );
or \U$3736 ( \12555 , \12494 , \12554 );
not \U$3737 ( \12556 , \12555 );
not \U$3738 ( \12557 , \9482 );
and \U$3739 ( \12558 , \12556 , \12557 );
nor \U$3740 ( \12559 , \12553 , \12558 );
nand \U$3741 ( \12560 , \12548 , \12559 );
not \U$3742 ( \12561 , \12560 );
not \U$3743 ( \12562 , \9471 );
not \U$3744 ( \12563 , \10972 );
or \U$3745 ( \12564 , \12494 , \12563 );
not \U$3746 ( \12565 , \12564 );
and \U$3747 ( \12566 , \12562 , \12565 );
not \U$3748 ( \12567 , \10968 );
or \U$3749 ( \12568 , \12494 , \12567 );
not \U$3750 ( \12569 , \12568 );
and \U$3751 ( \12570 , \12569 , \9476 );
nor \U$3752 ( \12571 , \12566 , \12570 );
not \U$3753 ( \12572 , \9463 );
not \U$3754 ( \12573 , \10941 );
or \U$3755 ( \12574 , \12494 , \12573 );
not \U$3756 ( \12575 , \12574 );
and \U$3757 ( \12576 , \12572 , \12575 );
not \U$3758 ( \12577 , \10978 );
or \U$3759 ( \12578 , \12494 , \12577 );
not \U$3760 ( \12579 , \12578 );
and \U$3761 ( \12580 , \12579 , \9468 );
nor \U$3762 ( \12581 , \12576 , \12580 );
and \U$3763 ( \12582 , \12561 , \12571 , \12581 );
nand \U$3764 ( \12583 , \12538 , \12582 );
not \U$3765 ( \12584 , \12583 );
not \U$3766 ( \12585 , \11067 );
and \U$3767 ( \12586 , \12585 , \12521 );
and \U$3768 ( \12587 , \12502 , \9034 );
nor \U$3769 ( \12588 , \12586 , \12587 );
not \U$3770 ( \12589 , \11060 );
not \U$3771 ( \12590 , \12511 );
and \U$3772 ( \12591 , \12589 , \12590 );
and \U$3773 ( \12592 , \12498 , \9014 );
nor \U$3774 ( \12593 , \12591 , \12592 );
nand \U$3775 ( \12594 , \12588 , \12593 );
not \U$3776 ( \12595 , \12594 );
not \U$3777 ( \12596 , \10370 );
not \U$3778 ( \12597 , \12551 );
and \U$3779 ( \12598 , \12596 , \12597 );
and \U$3780 ( \12599 , \12556 , \8970 );
nor \U$3781 ( \12600 , \12598 , \12599 );
not \U$3782 ( \12601 , \8980 );
and \U$3783 ( \12602 , \12601 , \12525 );
and \U$3784 ( \12603 , \12569 , \9009 );
nor \U$3785 ( \12604 , \12602 , \12603 );
and \U$3786 ( \12605 , \12595 , \12600 , \12604 );
not \U$3787 ( \12606 , \8977 );
and \U$3788 ( \12607 , \12606 , \12546 );
and \U$3789 ( \12608 , \12508 , \9006 );
nor \U$3790 ( \12609 , \12607 , \12608 );
not \U$3791 ( \12610 , \11036 );
not \U$3792 ( \12611 , \12530 );
and \U$3793 ( \12612 , \12610 , \12611 );
and \U$3794 ( \12613 , \12542 , \8966 );
nor \U$3795 ( \12614 , \12612 , \12613 );
nand \U$3796 ( \12615 , \12609 , \12614 );
not \U$3797 ( \12616 , \12615 );
not \U$3798 ( \12617 , \11046 );
not \U$3799 ( \12618 , \12574 );
and \U$3800 ( \12619 , \12617 , \12618 );
and \U$3801 ( \12620 , \12579 , \8990 );
nor \U$3802 ( \12621 , \12619 , \12620 );
not \U$3803 ( \12622 , \8997 );
and \U$3804 ( \12623 , \12622 , \12565 );
and \U$3805 ( \12624 , \12535 , \8999 );
nor \U$3806 ( \12625 , \12623 , \12624 );
and \U$3807 ( \12626 , \12616 , \12621 , \12625 );
nand \U$3808 ( \12627 , \12605 , \12626 );
xnor \U$3809 ( \12628 , RIb7b94a0_249, \12627 );
not \U$3810 ( \12629 , \11120 );
and \U$3811 ( \12630 , \12629 , \12521 );
and \U$3812 ( \12631 , \12502 , \9251 );
nor \U$3813 ( \12632 , \12630 , \12631 );
not \U$3814 ( \12633 , \11113 );
and \U$3815 ( \12634 , \12633 , \12590 );
and \U$3816 ( \12635 , \12498 , \9233 );
nor \U$3817 ( \12636 , \12634 , \12635 );
nand \U$3818 ( \12637 , \12632 , \12636 );
not \U$3819 ( \12638 , \12637 );
not \U$3820 ( \12639 , \10323 );
and \U$3821 ( \12640 , \12639 , \12597 );
and \U$3822 ( \12641 , \12556 , \9193 );
nor \U$3823 ( \12642 , \12640 , \12641 );
not \U$3824 ( \12643 , \11954 );
and \U$3825 ( \12644 , \12643 , \12525 );
and \U$3826 ( \12645 , \12569 , \9228 );
nor \U$3827 ( \12646 , \12644 , \12645 );
and \U$3828 ( \12647 , \12638 , \12642 , \12646 );
not \U$3829 ( \12648 , \9205 );
and \U$3830 ( \12649 , \12648 , \12546 );
and \U$3831 ( \12650 , \12508 , \9225 );
nor \U$3832 ( \12651 , \12649 , \12650 );
not \U$3833 ( \12652 , \11093 );
and \U$3834 ( \12653 , \12652 , \12611 );
and \U$3835 ( \12654 , \12542 , \9196 );
nor \U$3836 ( \12655 , \12653 , \12654 );
nand \U$3837 ( \12656 , \12651 , \12655 );
not \U$3838 ( \12657 , \12656 );
not \U$3839 ( \12658 , \11101 );
and \U$3840 ( \12659 , \12658 , \12618 );
and \U$3841 ( \12660 , \12579 , \9212 );
nor \U$3842 ( \12661 , \12659 , \12660 );
not \U$3843 ( \12662 , \9217 );
and \U$3844 ( \12663 , \12662 , \12565 );
and \U$3845 ( \12664 , \12535 , \9219 );
nor \U$3846 ( \12665 , \12663 , \12664 );
and \U$3847 ( \12666 , \12657 , \12661 , \12665 );
nand \U$3848 ( \12667 , \12647 , \12666 );
xnor \U$3849 ( \12668 , RIb7b9518_248, \12667 );
not \U$3850 ( \12669 , \11152 );
and \U$3851 ( \12670 , \12669 , \12590 );
and \U$3852 ( \12671 , \12498 , \9690 );
nor \U$3853 ( \12672 , \12670 , \12671 );
not \U$3854 ( \12673 , \10250 );
and \U$3855 ( \12674 , \12673 , \12521 );
and \U$3856 ( \12675 , \12502 , \9695 );
nor \U$3857 ( \12676 , \12674 , \12675 );
nand \U$3858 ( \12677 , \12672 , \12676 );
not \U$3859 ( \12678 , \12677 );
not \U$3860 ( \12679 , \11140 );
and \U$3861 ( \12680 , \12679 , \12569 );
and \U$3862 ( \12681 , \12525 , \9706 );
nor \U$3863 ( \12682 , \12680 , \12681 );
not \U$3864 ( \12683 , \10244 );
not \U$3865 ( \12684 , \12551 );
and \U$3866 ( \12685 , \12683 , \12684 );
and \U$3867 ( \12686 , \12556 , \9710 );
nor \U$3868 ( \12687 , \12685 , \12686 );
and \U$3869 ( \12688 , \12678 , \12682 , \12687 );
not \U$3870 ( \12689 , \9668 );
and \U$3871 ( \12690 , \12689 , \12611 );
and \U$3872 ( \12691 , \12542 , \9664 );
nor \U$3873 ( \12692 , \12690 , \12691 );
not \U$3874 ( \12693 , \9661 );
and \U$3875 ( \12694 , \12693 , \12508 );
and \U$3876 ( \12695 , \12546 , \9656 );
nor \U$3877 ( \12696 , \12694 , \12695 );
nand \U$3878 ( \12697 , \12692 , \12696 );
not \U$3879 ( \12698 , \12697 );
not \U$3880 ( \12699 , \11923 );
and \U$3881 ( \12700 , \12699 , \12618 );
and \U$3882 ( \12701 , \12579 , \9675 );
nor \U$3883 ( \12702 , \12700 , \12701 );
not \U$3884 ( \12703 , \9680 );
and \U$3885 ( \12704 , \12703 , \12565 );
and \U$3886 ( \12705 , \12535 , \9682 );
nor \U$3887 ( \12706 , \12704 , \12705 );
and \U$3888 ( \12707 , \12698 , \12702 , \12706 );
nand \U$3889 ( \12708 , \12688 , \12707 );
xnor \U$3890 ( \12709 , \12708 , \9719 );
not \U$3891 ( \12710 , \11193 );
and \U$3892 ( \12711 , \12710 , \12590 );
and \U$3893 ( \12712 , \12498 , \9755 );
nor \U$3894 ( \12713 , \12711 , \12712 );
not \U$3895 ( \12714 , \10197 );
and \U$3896 ( \12715 , \12714 , \12521 );
and \U$3897 ( \12716 , \12502 , \9763 );
nor \U$3898 ( \12717 , \12715 , \12716 );
nand \U$3899 ( \12718 , \12713 , \12717 );
not \U$3900 ( \12719 , \12718 );
not \U$3901 ( \12720 , \10182 );
and \U$3902 ( \12721 , \12720 , \12569 );
and \U$3903 ( \12722 , \12525 , \9772 );
nor \U$3904 ( \12723 , \12721 , \12722 );
not \U$3905 ( \12724 , \10188 );
and \U$3906 ( \12725 , \12724 , \12684 );
and \U$3907 ( \12726 , \12556 , \9776 );
nor \U$3908 ( \12727 , \12725 , \12726 );
and \U$3909 ( \12728 , \12719 , \12723 , \12727 );
not \U$3910 ( \12729 , \9732 );
and \U$3911 ( \12730 , \12729 , \12611 );
and \U$3912 ( \12731 , \12542 , \9728 );
nor \U$3913 ( \12732 , \12730 , \12731 );
not \U$3914 ( \12733 , \9725 );
and \U$3915 ( \12734 , \12733 , \12508 );
and \U$3916 ( \12735 , \12546 , \9721 );
nor \U$3917 ( \12736 , \12734 , \12735 );
nand \U$3918 ( \12737 , \12732 , \12736 );
not \U$3919 ( \12738 , \12737 );
not \U$3920 ( \12739 , \11876 );
and \U$3921 ( \12740 , \12739 , \12618 );
and \U$3922 ( \12741 , \12579 , \9739 );
nor \U$3923 ( \12742 , \12740 , \12741 );
not \U$3924 ( \12743 , \9745 );
and \U$3925 ( \12744 , \12743 , \12565 );
and \U$3926 ( \12745 , \12535 , \9747 );
nor \U$3927 ( \12746 , \12744 , \12745 );
and \U$3928 ( \12747 , \12738 , \12742 , \12746 );
nand \U$3929 ( \12748 , \12728 , \12747 );
xnor \U$3930 ( \12749 , \12748 , \9786 );
nor \U$3931 ( \12750 , \12709 , \12749 );
nand \U$3932 ( \12751 , \12628 , \12668 , \12750 );
not \U$3933 ( \12752 , \12751 );
not \U$3934 ( \12753 , \11293 );
and \U$3935 ( \12754 , \12753 , \12521 );
and \U$3936 ( \12755 , \12502 , \9319 );
nor \U$3937 ( \12756 , \12754 , \12755 );
not \U$3938 ( \12757 , \11288 );
and \U$3939 ( \12758 , \12757 , \12590 );
and \U$3940 ( \12759 , \12498 , \9302 );
nor \U$3941 ( \12760 , \12758 , \12759 );
nand \U$3942 ( \12761 , \12756 , \12760 );
not \U$3943 ( \12762 , \12761 );
not \U$3944 ( \12763 , \10415 );
and \U$3945 ( \12764 , \12763 , \12552 );
and \U$3946 ( \12765 , \12556 , \9265 );
nor \U$3947 ( \12766 , \12764 , \12765 );
not \U$3948 ( \12767 , \9273 );
and \U$3949 ( \12768 , \12767 , \12525 );
and \U$3950 ( \12769 , \12569 , \9297 );
nor \U$3951 ( \12770 , \12768 , \12769 );
and \U$3952 ( \12771 , \12762 , \12766 , \12770 );
not \U$3953 ( \12772 , \9270 );
and \U$3954 ( \12773 , \12772 , \12546 );
and \U$3955 ( \12774 , \12508 , \9295 );
nor \U$3956 ( \12775 , \12773 , \12774 );
not \U$3957 ( \12776 , \11270 );
and \U$3958 ( \12777 , \12776 , \12611 );
and \U$3959 ( \12778 , \12542 , \9262 );
nor \U$3960 ( \12779 , \12777 , \12778 );
nand \U$3961 ( \12780 , \12775 , \12779 );
not \U$3962 ( \12781 , \12780 );
not \U$3963 ( \12782 , \11276 );
and \U$3964 ( \12783 , \12782 , \12618 );
and \U$3965 ( \12784 , \12579 , \9281 );
nor \U$3966 ( \12785 , \12783 , \12784 );
not \U$3967 ( \12786 , \9287 );
and \U$3968 ( \12787 , \12786 , \12565 );
and \U$3969 ( \12788 , \12535 , \9289 );
nor \U$3970 ( \12789 , \12787 , \12788 );
and \U$3971 ( \12790 , \12781 , \12785 , \12789 );
nand \U$3972 ( \12791 , \12771 , \12790 );
xnor \U$3973 ( \12792 , \12791 , \9327 );
not \U$3974 ( \12793 , \11250 );
and \U$3975 ( \12794 , \12793 , \12521 );
and \U$3976 ( \12795 , \12502 , \9453 );
nor \U$3977 ( \12796 , \12794 , \12795 );
not \U$3978 ( \12797 , \11245 );
and \U$3979 ( \12798 , \12797 , \12590 );
and \U$3980 ( \12799 , \12498 , \9435 );
nor \U$3981 ( \12800 , \12798 , \12799 );
nand \U$3982 ( \12801 , \12796 , \12800 );
not \U$3983 ( \12802 , \12801 );
not \U$3984 ( \12803 , \10462 );
and \U$3985 ( \12804 , \12803 , \12597 );
and \U$3986 ( \12805 , \12556 , \9397 );
nor \U$3987 ( \12806 , \12804 , \12805 );
not \U$3988 ( \12807 , \9405 );
and \U$3989 ( \12808 , \12807 , \12525 );
and \U$3990 ( \12809 , \12569 , \9430 );
nor \U$3991 ( \12810 , \12808 , \12809 );
and \U$3992 ( \12811 , \12802 , \12806 , \12810 );
not \U$3993 ( \12812 , \9402 );
and \U$3994 ( \12813 , \12812 , \12546 );
and \U$3995 ( \12814 , \12508 , \9427 );
nor \U$3996 ( \12815 , \12813 , \12814 );
not \U$3997 ( \12816 , \11230 );
and \U$3998 ( \12817 , \12816 , \12611 );
and \U$3999 ( \12818 , \12542 , \9394 );
nor \U$4000 ( \12819 , \12817 , \12818 );
nand \U$4001 ( \12820 , \12815 , \12819 );
not \U$4002 ( \12821 , \12820 );
not \U$4003 ( \12822 , \10455 );
and \U$4004 ( \12823 , \12822 , \12618 );
and \U$4005 ( \12824 , \12579 , \9414 );
nor \U$4006 ( \12825 , \12823 , \12824 );
not \U$4007 ( \12826 , \9419 );
and \U$4008 ( \12827 , \12826 , \12565 );
and \U$4009 ( \12828 , \12535 , \9421 );
nor \U$4010 ( \12829 , \12827 , \12828 );
and \U$4011 ( \12830 , \12821 , \12825 , \12829 );
nand \U$4012 ( \12831 , \12811 , \12830 );
xnor \U$4013 ( \12832 , \12831 , \9460 );
nor \U$4014 ( \12833 , \12792 , \12832 );
not \U$4015 ( \12834 , \9647 );
and \U$4016 ( \12835 , \12834 , \12611 );
and \U$4017 ( \12836 , \12542 , \9643 );
nor \U$4018 ( \12837 , \12835 , \12836 );
not \U$4019 ( \12838 , \9640 );
and \U$4020 ( \12839 , \12838 , \12508 );
and \U$4021 ( \12840 , \12546 , \9636 );
nor \U$4022 ( \12841 , \12839 , \12840 );
nand \U$4023 ( \12842 , \12837 , \12841 );
not \U$4024 ( \12843 , \12842 );
not \U$4025 ( \12844 , \9625 );
and \U$4026 ( \12845 , \12844 , \12521 );
and \U$4027 ( \12846 , \12502 , \9619 );
nor \U$4028 ( \12847 , \12845 , \12846 );
not \U$4029 ( \12848 , \9632 );
and \U$4030 ( \12849 , \12848 , \12590 );
and \U$4031 ( \12850 , \12498 , \9628 );
nor \U$4032 ( \12851 , \12849 , \12850 );
and \U$4033 ( \12852 , \12843 , \12847 , \12851 );
not \U$4034 ( \12853 , \9588 );
and \U$4035 ( \12854 , \12853 , \12565 );
and \U$4036 ( \12855 , \12535 , \9593 );
nor \U$4037 ( \12856 , \12854 , \12855 );
not \U$4038 ( \12857 , \9597 );
and \U$4039 ( \12858 , \12857 , \12618 );
and \U$4040 ( \12859 , \12579 , \9600 );
nor \U$4041 ( \12860 , \12858 , \12859 );
nand \U$4042 ( \12861 , \12856 , \12860 );
not \U$4043 ( \12862 , \12861 );
not \U$4044 ( \12863 , \9607 );
and \U$4045 ( \12864 , \12863 , \12569 );
and \U$4046 ( \12865 , \12525 , \9603 );
nor \U$4047 ( \12866 , \12864 , \12865 );
not \U$4048 ( \12867 , \9611 );
and \U$4049 ( \12868 , \12867 , \12597 );
and \U$4050 ( \12869 , \12556 , \9613 );
nor \U$4051 ( \12870 , \12868 , \12869 );
and \U$4052 ( \12871 , \12862 , \12866 , \12870 );
nand \U$4053 ( \12872 , \12852 , \12871 );
xnor \U$4054 ( \12873 , \12872 , \9653 );
not \U$4055 ( \12874 , \9385 );
not \U$4056 ( \12875 , \12874 );
and \U$4057 ( \12876 , \12875 , \12521 );
and \U$4058 ( \12877 , \12502 , \9377 );
nor \U$4059 ( \12878 , \12876 , \12877 );
not \U$4060 ( \12879 , \11365 );
and \U$4061 ( \12880 , \12879 , \12590 );
and \U$4062 ( \12881 , \12498 , \9369 );
nor \U$4063 ( \12882 , \12880 , \12881 );
nand \U$4064 ( \12883 , \12878 , \12882 );
not \U$4065 ( \12884 , \12883 );
not \U$4066 ( \12885 , \10553 );
and \U$4067 ( \12886 , \12885 , \12552 );
and \U$4068 ( \12887 , \12556 , \9334 );
nor \U$4069 ( \12888 , \12886 , \12887 );
not \U$4070 ( \12889 , \9342 );
and \U$4071 ( \12890 , \12889 , \12525 );
and \U$4072 ( \12891 , \12569 , \9364 );
nor \U$4073 ( \12892 , \12890 , \12891 );
and \U$4074 ( \12893 , \12884 , \12888 , \12892 );
not \U$4075 ( \12894 , \9339 );
and \U$4076 ( \12895 , \12894 , \12546 );
and \U$4077 ( \12896 , \12508 , \9361 );
nor \U$4078 ( \12897 , \12895 , \12896 );
not \U$4079 ( \12898 , \11393 );
and \U$4080 ( \12899 , \12898 , \12611 );
and \U$4081 ( \12900 , \12542 , \9331 );
nor \U$4082 ( \12901 , \12899 , \12900 );
nand \U$4083 ( \12902 , \12897 , \12901 );
not \U$4084 ( \12903 , \12902 );
not \U$4085 ( \12904 , \12141 );
and \U$4086 ( \12905 , \12904 , \12618 );
and \U$4087 ( \12906 , \12579 , \9348 );
nor \U$4088 ( \12907 , \12905 , \12906 );
not \U$4089 ( \12908 , \9354 );
and \U$4090 ( \12909 , \12908 , \12565 );
and \U$4091 ( \12910 , \12535 , \9356 );
nor \U$4092 ( \12911 , \12909 , \12910 );
and \U$4093 ( \12912 , \12903 , \12907 , \12911 );
nand \U$4094 ( \12913 , \12893 , \12912 );
xnor \U$4095 ( \12914 , \12913 , \9392 );
nor \U$4096 ( \12915 , \12873 , \12914 );
and \U$4097 ( \12916 , \12752 , \12833 , \12915 );
not \U$4098 ( \12917 , \11431 );
and \U$4099 ( \12918 , \12917 , \12521 );
and \U$4100 ( \12919 , \12502 , \9180 );
nor \U$4101 ( \12920 , \12918 , \12919 );
not \U$4102 ( \12921 , \11426 );
and \U$4103 ( \12922 , \12921 , \12590 );
and \U$4104 ( \12923 , \12498 , \9163 );
nor \U$4105 ( \12924 , \12922 , \12923 );
nand \U$4106 ( \12925 , \12920 , \12924 );
not \U$4107 ( \12926 , \12925 );
not \U$4108 ( \12927 , \10901 );
and \U$4109 ( \12928 , \12927 , \12552 );
and \U$4110 ( \12929 , \12556 , \9124 );
nor \U$4111 ( \12930 , \12928 , \12929 );
not \U$4112 ( \12931 , \9133 );
and \U$4113 ( \12932 , \12931 , \12525 );
and \U$4114 ( \12933 , \12569 , \9157 );
nor \U$4115 ( \12934 , \12932 , \12933 );
and \U$4116 ( \12935 , \12926 , \12930 , \12934 );
not \U$4117 ( \12936 , \9130 );
and \U$4118 ( \12937 , \12936 , \12546 );
and \U$4119 ( \12938 , \12508 , \9155 );
nor \U$4120 ( \12939 , \12937 , \12938 );
not \U$4121 ( \12940 , \11410 );
and \U$4122 ( \12941 , \12940 , \12531 );
and \U$4123 ( \12942 , \12542 , \9121 );
nor \U$4124 ( \12943 , \12941 , \12942 );
nand \U$4125 ( \12944 , \12939 , \12943 );
not \U$4126 ( \12945 , \12944 );
not \U$4127 ( \12946 , \11416 );
and \U$4128 ( \12947 , \12946 , \12575 );
and \U$4129 ( \12948 , \12579 , \9142 );
nor \U$4130 ( \12949 , \12947 , \12948 );
not \U$4131 ( \12950 , \9148 );
and \U$4132 ( \12951 , \12950 , \12565 );
and \U$4133 ( \12952 , \12535 , \9150 );
nor \U$4134 ( \12953 , \12951 , \12952 );
and \U$4135 ( \12954 , \12945 , \12949 , \12953 );
nand \U$4136 ( \12955 , \12935 , \12954 );
xnor \U$4137 ( \12956 , RIb7af6a8_253, \12955 );
not \U$4138 ( \12957 , \11473 );
and \U$4139 ( \12958 , \12957 , \12521 );
and \U$4140 ( \12959 , \12502 , \9112 );
nor \U$4141 ( \12960 , \12958 , \12959 );
not \U$4142 ( \12961 , \11468 );
and \U$4143 ( \12962 , \12961 , \12590 );
and \U$4144 ( \12963 , \12498 , \9093 );
nor \U$4145 ( \12964 , \12962 , \12963 );
nand \U$4146 ( \12965 , \12960 , \12964 );
not \U$4147 ( \12966 , \12965 );
not \U$4148 ( \12967 , \10859 );
and \U$4149 ( \12968 , \12967 , \12597 );
and \U$4150 ( \12969 , \12556 , \9049 );
nor \U$4151 ( \12970 , \12968 , \12969 );
not \U$4152 ( \12971 , \9058 );
and \U$4153 ( \12972 , \12971 , \12525 );
and \U$4154 ( \12973 , \12569 , \9085 );
nor \U$4155 ( \12974 , \12972 , \12973 );
and \U$4156 ( \12975 , \12966 , \12970 , \12974 );
not \U$4157 ( \12976 , \9055 );
and \U$4158 ( \12977 , \12976 , \12546 );
and \U$4159 ( \12978 , \12508 , \9081 );
nor \U$4160 ( \12979 , \12977 , \12978 );
not \U$4161 ( \12980 , \11452 );
and \U$4162 ( \12981 , \12980 , \12531 );
and \U$4163 ( \12982 , \12542 , \9046 );
nor \U$4164 ( \12983 , \12981 , \12982 );
nand \U$4165 ( \12984 , \12979 , \12983 );
not \U$4166 ( \12985 , \12984 );
not \U$4167 ( \12986 , \11458 );
and \U$4168 ( \12987 , \12986 , \12575 );
and \U$4169 ( \12988 , \12579 , \9067 );
nor \U$4170 ( \12989 , \12987 , \12988 );
not \U$4171 ( \12990 , \9073 );
and \U$4172 ( \12991 , \12990 , \12565 );
and \U$4173 ( \12992 , \12535 , \9075 );
nor \U$4174 ( \12993 , \12991 , \12992 );
and \U$4175 ( \12994 , \12985 , \12989 , \12993 );
nand \U$4176 ( \12995 , \12975 , \12994 );
xnor \U$4177 ( \12996 , RIb7af720_252, \12995 );
not \U$4178 ( \12997 , \9851 );
and \U$4179 ( \12998 , \12997 , \12611 );
and \U$4180 ( \12999 , \12542 , \9847 );
nor \U$4181 ( \13000 , \12998 , \12999 );
not \U$4182 ( \13001 , \9843 );
and \U$4183 ( \13002 , \13001 , \12508 );
and \U$4184 ( \13003 , \12546 , \9839 );
nor \U$4185 ( \13004 , \13002 , \13003 );
nand \U$4186 ( \13005 , \13000 , \13004 );
not \U$4187 ( \13006 , \13005 );
not \U$4188 ( \13007 , \9827 );
and \U$4189 ( \13008 , \13007 , \12521 );
and \U$4190 ( \13009 , \12502 , \9822 );
nor \U$4191 ( \13010 , \13008 , \13009 );
not \U$4192 ( \13011 , \9834 );
and \U$4193 ( \13012 , \13011 , \12590 );
and \U$4194 ( \13013 , \12498 , \9830 );
nor \U$4195 ( \13014 , \13012 , \13013 );
and \U$4196 ( \13015 , \13006 , \13010 , \13014 );
not \U$4197 ( \13016 , \9791 );
and \U$4198 ( \13017 , \13016 , \12565 );
and \U$4199 ( \13018 , \12535 , \9794 );
nor \U$4200 ( \13019 , \13017 , \13018 );
not \U$4201 ( \13020 , \9798 );
and \U$4202 ( \13021 , \13020 , \12618 );
and \U$4203 ( \13022 , \12579 , \9801 );
nor \U$4204 ( \13023 , \13021 , \13022 );
nand \U$4205 ( \13024 , \13019 , \13023 );
not \U$4206 ( \13025 , \13024 );
not \U$4207 ( \13026 , \9809 );
and \U$4208 ( \13027 , \13026 , \12569 );
and \U$4209 ( \13028 , \12525 , \9805 );
nor \U$4210 ( \13029 , \13027 , \13028 );
not \U$4211 ( \13030 , \9814 );
and \U$4212 ( \13031 , \13030 , \12597 );
and \U$4213 ( \13032 , \12556 , \9816 );
nor \U$4214 ( \13033 , \13031 , \13032 );
and \U$4215 ( \13034 , \13025 , \13029 , \13033 );
nand \U$4216 ( \13035 , \13015 , \13034 );
xnor \U$4217 ( \13036 , \13035 , \9857 );
not \U$4218 ( \13037 , \11545 );
and \U$4219 ( \13038 , \13037 , \12521 );
and \U$4220 ( \13039 , \12502 , \8953 );
nor \U$4221 ( \13040 , \13038 , \13039 );
not \U$4222 ( \13041 , \11540 );
and \U$4223 ( \13042 , \13041 , \12590 );
and \U$4224 ( \13043 , \12498 , \8927 );
nor \U$4225 ( \13044 , \13042 , \13043 );
nand \U$4226 ( \13045 , \13040 , \13044 );
not \U$4227 ( \13046 , \13045 );
not \U$4228 ( \13047 , \10775 );
and \U$4229 ( \13048 , \13047 , \12597 );
and \U$4230 ( \13049 , \12556 , \8843 );
nor \U$4231 ( \13050 , \13048 , \13049 );
not \U$4232 ( \13051 , \8861 );
and \U$4233 ( \13052 , \13051 , \12525 );
and \U$4234 ( \13053 , \12569 , \8915 );
nor \U$4235 ( \13054 , \13052 , \13053 );
and \U$4236 ( \13055 , \13046 , \13050 , \13054 );
not \U$4237 ( \13056 , \8853 );
and \U$4238 ( \13057 , \13056 , \12546 );
and \U$4239 ( \13058 , \12508 , \8904 );
nor \U$4240 ( \13059 , \13057 , \13058 );
not \U$4241 ( \13060 , \11565 );
and \U$4242 ( \13061 , \13060 , \12611 );
and \U$4243 ( \13062 , \12542 , \8827 );
nor \U$4244 ( \13063 , \13061 , \13062 );
nand \U$4245 ( \13064 , \13059 , \13063 );
not \U$4246 ( \13065 , \13064 );
not \U$4247 ( \13066 , \12351 );
and \U$4248 ( \13067 , \13066 , \12618 );
and \U$4249 ( \13068 , \12579 , \8881 );
nor \U$4250 ( \13069 , \13067 , \13068 );
not \U$4251 ( \13070 , \8894 );
and \U$4252 ( \13071 , \13070 , \12565 );
and \U$4253 ( \13072 , \12535 , \8896 );
nor \U$4254 ( \13073 , \13071 , \13072 );
and \U$4255 ( \13074 , \13065 , \13069 , \13073 );
nand \U$4256 ( \13075 , \13055 , \13074 );
xnor \U$4257 ( \13076 , \13075 , \8964 );
nor \U$4258 ( \13077 , \13036 , \13076 );
nand \U$4259 ( \13078 , \12956 , \12996 , \13077 );
not \U$4260 ( \13079 , \13078 );
not \U$4261 ( \13080 , \9579 );
and \U$4262 ( \13081 , \13080 , \12611 );
and \U$4263 ( \13082 , \12542 , \9575 );
nor \U$4264 ( \13083 , \13081 , \13082 );
not \U$4265 ( \13084 , \9572 );
and \U$4266 ( \13085 , \13084 , \12508 );
and \U$4267 ( \13086 , \12546 , \9568 );
nor \U$4268 ( \13087 , \13085 , \13086 );
nand \U$4269 ( \13088 , \13083 , \13087 );
not \U$4270 ( \13089 , \13088 );
not \U$4271 ( \13090 , \9557 );
and \U$4272 ( \13091 , \13090 , \12521 );
and \U$4273 ( \13092 , \12502 , \9551 );
nor \U$4274 ( \13093 , \13091 , \13092 );
not \U$4275 ( \13094 , \9564 );
and \U$4276 ( \13095 , \13094 , \12590 );
and \U$4277 ( \13096 , \12498 , \9560 );
nor \U$4278 ( \13097 , \13095 , \13096 );
and \U$4279 ( \13098 , \13089 , \13093 , \13097 );
not \U$4280 ( \13099 , \9519 );
and \U$4281 ( \13100 , \13099 , \12565 );
and \U$4282 ( \13101 , \12535 , \9523 );
nor \U$4283 ( \13102 , \13100 , \13101 );
not \U$4284 ( \13103 , \9527 );
and \U$4285 ( \13104 , \13103 , \12618 );
and \U$4286 ( \13105 , \12579 , \9530 );
nor \U$4287 ( \13106 , \13104 , \13105 );
nand \U$4288 ( \13107 , \13102 , \13106 );
not \U$4289 ( \13108 , \13107 );
not \U$4290 ( \13109 , \9537 );
and \U$4291 ( \13110 , \13109 , \12569 );
and \U$4292 ( \13111 , \12525 , \9533 );
nor \U$4293 ( \13112 , \13110 , \13111 );
not \U$4294 ( \13113 , \9543 );
and \U$4295 ( \13114 , \13113 , \12552 );
and \U$4296 ( \13115 , \12556 , \9545 );
nor \U$4297 ( \13116 , \13114 , \13115 );
and \U$4298 ( \13117 , \13108 , \13112 , \13116 );
nand \U$4299 ( \13118 , \13098 , \13117 );
xnor \U$4300 ( \13119 , \13118 , \9585 );
not \U$4301 ( \13120 , \11635 );
and \U$4302 ( \13121 , \13120 , \12546 );
and \U$4303 ( \13122 , \12508 , \9975 );
nor \U$4304 ( \13123 , \13121 , \13122 );
not \U$4305 ( \13124 , \12282 );
and \U$4306 ( \13125 , \13124 , \12611 );
and \U$4307 ( \13126 , \12542 , \9982 );
nor \U$4308 ( \13127 , \13125 , \13126 );
nand \U$4309 ( \13128 , \13123 , \13127 );
not \U$4310 ( \13129 , \13128 );
not \U$4311 ( \13130 , \11623 );
and \U$4312 ( \13131 , \13130 , \12512 );
and \U$4313 ( \13132 , \12498 , \10709 );
nor \U$4314 ( \13133 , \13131 , \13132 );
not \U$4315 ( \13134 , \11620 );
and \U$4316 ( \13135 , \13134 , \12521 );
and \U$4317 ( \13136 , \12502 , \9968 );
nor \U$4318 ( \13137 , \13135 , \13136 );
and \U$4319 ( \13138 , \13129 , \13133 , \13137 );
not \U$4320 ( \13139 , \9952 );
and \U$4321 ( \13140 , \13139 , \12565 );
and \U$4322 ( \13141 , \12535 , \9954 );
nor \U$4323 ( \13142 , \13140 , \13141 );
not \U$4324 ( \13143 , \9944 );
not \U$4325 ( \13144 , \13143 );
and \U$4326 ( \13145 , \13144 , \12618 );
and \U$4327 ( \13146 , \12579 , \9947 );
nor \U$4328 ( \13147 , \13145 , \13146 );
nand \U$4329 ( \13148 , \13142 , \13147 );
not \U$4330 ( \13149 , \13148 );
not \U$4331 ( \13150 , \9933 );
and \U$4332 ( \13151 , \13150 , \12569 );
and \U$4333 ( \13152 , \12525 , \9929 );
nor \U$4334 ( \13153 , \13151 , \13152 );
not \U$4335 ( \13154 , \9937 );
and \U$4336 ( \13155 , \13154 , \12597 );
and \U$4337 ( \13156 , \12556 , \9939 );
nor \U$4338 ( \13157 , \13155 , \13156 );
and \U$4339 ( \13158 , \13149 , \13153 , \13157 );
nand \U$4340 ( \13159 , \13138 , \13158 );
xnor \U$4341 ( \13160 , \13159 , \9990 );
nor \U$4342 ( \13161 , \13119 , \13160 );
not \U$4343 ( \13162 , \11674 );
and \U$4344 ( \13163 , \13162 , \12611 );
and \U$4345 ( \13164 , \12542 , \10047 );
nor \U$4346 ( \13165 , \13163 , \13164 );
not \U$4347 ( \13166 , \12222 );
and \U$4348 ( \13167 , \13166 , \12508 );
and \U$4349 ( \13168 , \12546 , \10043 );
nor \U$4350 ( \13169 , \13167 , \13168 );
nand \U$4351 ( \13170 , \13165 , \13169 );
not \U$4352 ( \13171 , \13170 );
not \U$4353 ( \13172 , \11698 );
and \U$4354 ( \13173 , \13172 , \12521 );
and \U$4355 ( \13174 , \12502 , \10035 );
nor \U$4356 ( \13175 , \13173 , \13174 );
not \U$4357 ( \13176 , \11693 );
and \U$4358 ( \13177 , \13176 , \12590 );
and \U$4359 ( \13178 , \12498 , \10027 );
nor \U$4360 ( \13179 , \13177 , \13178 );
and \U$4361 ( \13180 , \13171 , \13175 , \13179 );
not \U$4362 ( \13181 , \10002 );
and \U$4363 ( \13182 , \13181 , \12565 );
and \U$4364 ( \13183 , \12535 , \10004 );
nor \U$4365 ( \13184 , \13182 , \13183 );
not \U$4366 ( \13185 , \11666 );
and \U$4367 ( \13186 , \13185 , \12618 );
and \U$4368 ( \13187 , \12579 , \9996 );
nor \U$4369 ( \13188 , \13186 , \13187 );
nand \U$4370 ( \13189 , \13184 , \13188 );
not \U$4371 ( \13190 , \13189 );
not \U$4372 ( \13191 , \10013 );
and \U$4373 ( \13192 , \13191 , \12569 );
and \U$4374 ( \13193 , \12525 , \10009 );
nor \U$4375 ( \13194 , \13192 , \13193 );
not \U$4376 ( \13195 , \10018 );
and \U$4377 ( \13196 , \13195 , \12552 );
and \U$4378 ( \13197 , \12556 , \10020 );
nor \U$4379 ( \13198 , \13196 , \13197 );
and \U$4380 ( \13199 , \13190 , \13194 , \13198 );
nand \U$4381 ( \13200 , \13180 , \13199 );
xnor \U$4382 ( \13201 , \13200 , \10055 );
not \U$4383 ( \13202 , \9921 );
and \U$4384 ( \13203 , \13202 , \12611 );
and \U$4385 ( \13204 , \12542 , \9917 );
nor \U$4386 ( \13205 , \13203 , \13204 );
not \U$4387 ( \13206 , \9914 );
and \U$4388 ( \13207 , \13206 , \12508 );
and \U$4389 ( \13208 , \12546 , \9910 );
nor \U$4390 ( \13209 , \13207 , \13208 );
nand \U$4391 ( \13210 , \13205 , \13209 );
not \U$4392 ( \13211 , \13210 );
not \U$4393 ( \13212 , \9898 );
and \U$4394 ( \13213 , \13212 , \12521 );
and \U$4395 ( \13214 , \12502 , \9892 );
nor \U$4396 ( \13215 , \13213 , \13214 );
not \U$4397 ( \13216 , \9906 );
and \U$4398 ( \13217 , \13216 , \12512 );
and \U$4399 ( \13218 , \12498 , \9902 );
nor \U$4400 ( \13219 , \13217 , \13218 );
and \U$4401 ( \13220 , \13211 , \13215 , \13219 );
not \U$4402 ( \13221 , \9860 );
and \U$4403 ( \13222 , \13221 , \12565 );
and \U$4404 ( \13223 , \12535 , \9864 );
nor \U$4405 ( \13224 , \13222 , \13223 );
not \U$4406 ( \13225 , \9868 );
and \U$4407 ( \13226 , \13225 , \12618 );
and \U$4408 ( \13227 , \12579 , \9871 );
nor \U$4409 ( \13228 , \13226 , \13227 );
nand \U$4410 ( \13229 , \13224 , \13228 );
not \U$4411 ( \13230 , \13229 );
not \U$4412 ( \13231 , \9878 );
and \U$4413 ( \13232 , \13231 , \12569 );
and \U$4414 ( \13233 , \12525 , \9874 );
nor \U$4415 ( \13234 , \13232 , \13233 );
not \U$4416 ( \13235 , \9884 );
and \U$4417 ( \13236 , \13235 , \12552 );
and \U$4418 ( \13237 , \12556 , \9886 );
nor \U$4419 ( \13238 , \13236 , \13237 );
and \U$4420 ( \13239 , \13230 , \13234 , \13238 );
nand \U$4421 ( \13240 , \13220 , \13239 );
xnor \U$4422 ( \13241 , \13240 , \9927 );
nor \U$4423 ( \13242 , \13201 , \13241 );
and \U$4424 ( \13243 , \13079 , \13161 , \13242 );
nand \U$4425 ( \13244 , \12584 , \12916 , \13243 );
not \U$4426 ( \13245 , \13244 );
not \U$4427 ( \13246 , \13245 );
or \U$4428 ( \13247 , \12486 , \13246 );
not \U$4429 ( \13248 , \11754 );
or \U$4430 ( \13249 , \10065 , \13248 );
nand \U$4431 ( \13250 , \8906 , \10917 );
nand \U$4432 ( \13251 , \13249 , \13250 );
not \U$4433 ( \13252 , \13251 );
not \U$4434 ( \13253 , \12453 );
nand \U$4435 ( \13254 , \8837 , \13253 );
not \U$4436 ( \13255 , \13254 );
not \U$4437 ( \13256 , \10917 );
nand \U$4438 ( \13257 , \13255 , \13256 );
nand \U$4439 ( \13258 , \13252 , \13257 );
or \U$4440 ( \13259 , \9285 , \9492 );
or \U$4441 ( \13260 , \9494 , \9539 );
nand \U$4442 ( \13261 , \13259 , \13260 );
not \U$4443 ( \13262 , \9500 );
not \U$4444 ( \13263 , \13262 );
or \U$4445 ( \13264 , \13263 , \9002 );
or \U$4446 ( \13265 , \9498 , \9998 );
nand \U$4447 ( \13266 , \13264 , \13265 );
nor \U$4448 ( \13267 , \13261 , \13266 );
nand \U$4449 ( \13268 , \12453 , \10078 );
not \U$4450 ( \13269 , \13268 );
not \U$4451 ( \13270 , \9509 );
and \U$4452 ( \13271 , \13269 , \13270 );
or \U$4453 ( \13272 , \9504 , \9206 );
or \U$4454 ( \13273 , \9506 , \8879 );
nand \U$4455 ( \13274 , \13272 , \13273 );
not \U$4456 ( \13275 , \9015 );
and \U$4457 ( \13276 , \10120 , \13275 );
nor \U$4458 ( \13277 , \13271 , \13274 , \13276 );
not \U$4459 ( \13278 , \10078 );
or \U$4460 ( \13279 , \13278 , \8906 );
or \U$4461 ( \13280 , \9480 , \13279 );
not \U$4462 ( \13281 , \12490 );
or \U$4463 ( \13282 , \9482 , \13281 );
nand \U$4464 ( \13283 , \13280 , \13282 );
not \U$4465 ( \13284 , \10031 );
and \U$4466 ( \13285 , \10986 , \13284 );
not \U$4467 ( \13286 , \8955 );
not \U$4468 ( \13287 , \13286 );
and \U$4469 ( \13288 , \9468 , \13287 );
nor \U$4470 ( \13289 , \13285 , \13288 );
not \U$4471 ( \13290 , \9471 );
and \U$4472 ( \13291 , \13290 , \9753 );
and \U$4473 ( \13292 , \8913 , \9476 );
nor \U$4474 ( \13293 , \13291 , \13292 );
not \U$4475 ( \13294 , \10097 );
or \U$4476 ( \13295 , \8906 , \13294 );
not \U$4477 ( \13296 , \13295 );
and \U$4478 ( \13297 , \13296 , \10163 );
not \U$4479 ( \13298 , \8862 );
and \U$4480 ( \13299 , \13298 , \10168 );
nor \U$4481 ( \13300 , \13297 , \13299 );
nand \U$4482 ( \13301 , \13289 , \13293 , \13300 );
nor \U$4483 ( \13302 , \13283 , \13301 );
nand \U$4484 ( \13303 , \13267 , \13277 , \13302 );
not \U$4485 ( \13304 , \13303 );
not \U$4486 ( \13305 , \9728 );
or \U$4487 ( \13306 , \13305 , \13295 );
nand \U$4488 ( \13307 , \9731 , \13269 );
not \U$4489 ( \13308 , \9539 );
and \U$4490 ( \13309 , \9724 , \13308 );
not \U$4491 ( \13310 , \9202 );
and \U$4492 ( \13311 , \9721 , \13310 );
nor \U$4493 ( \13312 , \13309 , \13311 );
or \U$4494 ( \13313 , \9740 , \8956 );
or \U$4495 ( \13314 , \11876 , \10031 );
nand \U$4496 ( \13315 , \13313 , \13314 );
not \U$4497 ( \13316 , \9747 );
or \U$4498 ( \13317 , \13316 , \9015 );
or \U$4499 ( \13318 , \9745 , \9160 );
nand \U$4500 ( \13319 , \13317 , \13318 );
nor \U$4501 ( \13320 , \13315 , \13319 );
and \U$4502 ( \13321 , \13306 , \13307 , \13312 , \13320 );
not \U$4503 ( \13322 , \13321 );
not \U$4504 ( \13323 , \13322 );
not \U$4505 ( \13324 , \9759 );
not \U$4506 ( \13325 , \9411 );
or \U$4507 ( \13326 , \13324 , \13325 );
or \U$4508 ( \13327 , \10194 , \9998 );
nand \U$4509 ( \13328 , \13326 , \13327 );
or \U$4510 ( \13329 , \9285 , \11193 );
or \U$4511 ( \13330 , \11195 , \9423 );
nand \U$4512 ( \13331 , \13329 , \13330 );
nor \U$4513 ( \13332 , \13328 , \13331 );
not \U$4514 ( \13333 , \10188 );
not \U$4515 ( \13334 , \13279 );
and \U$4516 ( \13335 , \13333 , \13334 );
not \U$4517 ( \13336 , \13281 );
and \U$4518 ( \13337 , \9776 , \13336 );
or \U$4519 ( \13338 , \10178 , \9206 );
or \U$4520 ( \13339 , \10182 , \9844 );
nand \U$4521 ( \13340 , \13338 , \13339 );
nor \U$4522 ( \13341 , \13335 , \13337 , \13340 );
and \U$4523 ( \13342 , \13323 , \13332 , \13341 );
xnor \U$4524 ( \13343 , \13342 , \9786 );
not \U$4525 ( \13344 , \9664 );
or \U$4526 ( \13345 , \13344 , \13295 );
not \U$4527 ( \13346 , \13269 );
or \U$4528 ( \13347 , \9668 , \13346 );
not \U$4529 ( \13348 , \9702 );
and \U$4530 ( \13349 , \9660 , \13348 );
not \U$4531 ( \13350 , \9202 );
and \U$4532 ( \13351 , \9656 , \13350 );
nor \U$4533 ( \13352 , \13349 , \13351 );
not \U$4534 ( \13353 , \8955 );
or \U$4535 ( \13354 , \9676 , \13353 );
or \U$4536 ( \13355 , \11923 , \9248 );
nand \U$4537 ( \13356 , \13354 , \13355 );
not \U$4538 ( \13357 , \9682 );
or \U$4539 ( \13358 , \13357 , \8929 );
or \U$4540 ( \13359 , \9680 , \8924 );
nand \U$4541 ( \13360 , \13358 , \13359 );
nor \U$4542 ( \13361 , \13356 , \13360 );
and \U$4543 ( \13362 , \13345 , \13347 , \13352 , \13361 );
not \U$4544 ( \13363 , \13362 );
not \U$4545 ( \13364 , \13363 );
not \U$4546 ( \13365 , \9692 );
not \U$4547 ( \13366 , \9139 );
or \U$4548 ( \13367 , \13365 , \13366 );
or \U$4549 ( \13368 , \10248 , \9998 );
nand \U$4550 ( \13369 , \13367 , \13368 );
or \U$4551 ( \13370 , \9146 , \11152 );
or \U$4552 ( \13371 , \11154 , \9002 );
nand \U$4553 ( \13372 , \13370 , \13371 );
nor \U$4554 ( \13373 , \13369 , \13372 );
not \U$4555 ( \13374 , \10244 );
and \U$4556 ( \13375 , \13374 , \13334 );
not \U$4557 ( \13376 , \13281 );
and \U$4558 ( \13377 , \9710 , \13376 );
or \U$4559 ( \13378 , \11138 , \8858 );
or \U$4560 ( \13379 , \11140 , \8911 );
nand \U$4561 ( \13380 , \13378 , \13379 );
nor \U$4562 ( \13381 , \13375 , \13377 , \13380 );
and \U$4563 ( \13382 , \13364 , \13373 , \13381 );
xnor \U$4564 ( \13383 , \13382 , \9719 );
not \U$4565 ( \13384 , \9242 );
or \U$4566 ( \13385 , \13384 , \13279 );
or \U$4567 ( \13386 , \11088 , \12491 );
nand \U$4568 ( \13387 , \13385 , \13386 );
not \U$4569 ( \13388 , \13387 );
nand \U$4570 ( \13389 , \9204 , \13298 );
buf \U$4571 ( \13390 , \8857 );
nand \U$4572 ( \13391 , \9200 , \13390 );
not \U$4573 ( \13392 , \9844 );
and \U$4574 ( \13393 , \9228 , \13392 );
not \U$4575 ( \13394 , \8918 );
and \U$4576 ( \13395 , \9225 , \13394 );
nor \U$4577 ( \13396 , \13393 , \13395 );
nand \U$4578 ( \13397 , \13389 , \13391 , \13396 );
or \U$4579 ( \13398 , \11111 , \9221 );
nand \U$4580 ( \13399 , \9251 , \8886 );
nand \U$4581 ( \13400 , \9247 , \8878 );
nand \U$4582 ( \13401 , \9230 , \9351 );
and \U$4583 ( \13402 , \13398 , \13399 , \13400 , \13401 );
not \U$4584 ( \13403 , \13402 );
nor \U$4585 ( \13404 , \13397 , \13403 );
buf \U$4586 ( \13405 , \8923 );
nand \U$4587 ( \13406 , \9216 , \13405 );
nand \U$4588 ( \13407 , \9219 , \9757 );
not \U$4589 ( \13408 , \9760 );
and \U$4590 ( \13409 , \9210 , \13408 );
not \U$4591 ( \13410 , \8956 );
and \U$4592 ( \13411 , \9212 , \13410 );
nor \U$4593 ( \13412 , \13409 , \13411 );
nand \U$4594 ( \13413 , \13406 , \13407 , \13412 );
not \U$4595 ( \13414 , \9239 );
or \U$4596 ( \13415 , \13414 , \13268 );
or \U$4597 ( \13416 , \9197 , \13295 );
nand \U$4598 ( \13417 , \13415 , \13416 );
nor \U$4599 ( \13418 , \13413 , \13417 );
nand \U$4600 ( \13419 , \13388 , \13404 , \13418 );
xnor \U$4601 ( \13420 , \13419 , \9260 );
not \U$4602 ( \13421 , \9025 );
or \U$4603 ( \13422 , \13421 , \13279 );
or \U$4604 ( \13423 , \8971 , \12491 );
nand \U$4605 ( \13424 , \13422 , \13423 );
not \U$4606 ( \13425 , \13424 );
nand \U$4607 ( \13426 , \8976 , \8981 );
buf \U$4608 ( \13427 , \8857 );
nand \U$4609 ( \13428 , \8979 , \13427 );
not \U$4610 ( \13429 , \8911 );
and \U$4611 ( \13430 , \9009 , \13429 );
not \U$4612 ( \13431 , \9702 );
and \U$4613 ( \13432 , \9006 , \13431 );
nor \U$4614 ( \13433 , \13430 , \13432 );
nand \U$4615 ( \13434 , \13426 , \13428 , \13433 );
or \U$4616 ( \13435 , \11058 , \9291 );
nand \U$4617 ( \13436 , \9034 , \9213 );
nand \U$4618 ( \13437 , \9030 , \9411 );
nand \U$4619 ( \13438 , \9011 , \9351 );
and \U$4620 ( \13439 , \13435 , \13436 , \13437 , \13438 );
not \U$4621 ( \13440 , \13439 );
nor \U$4622 ( \13441 , \13434 , \13440 );
nand \U$4623 ( \13442 , \8996 , \9960 );
nand \U$4624 ( \13443 , \8999 , \9963 );
not \U$4625 ( \13444 , \8950 );
and \U$4626 ( \13445 , \8986 , \13444 );
not \U$4627 ( \13446 , \13353 );
and \U$4628 ( \13447 , \8990 , \13446 );
nor \U$4629 ( \13448 , \13445 , \13447 );
nand \U$4630 ( \13449 , \13442 , \13443 , \13448 );
not \U$4631 ( \13450 , \9020 );
or \U$4632 ( \13451 , \13450 , \13268 );
or \U$4633 ( \13452 , \8967 , \13295 );
nand \U$4634 ( \13453 , \13451 , \13452 );
nor \U$4635 ( \13454 , \13449 , \13453 );
nand \U$4636 ( \13455 , \13425 , \13441 , \13454 );
xnor \U$4637 ( \13456 , \13455 , \9044 );
nor \U$4638 ( \13457 , \13420 , \13456 );
nand \U$4639 ( \13458 , \13343 , \13383 , \13457 );
not \U$4640 ( \13459 , \13458 );
not \U$4641 ( \13460 , \9310 );
or \U$4642 ( \13461 , \13460 , \13279 );
or \U$4643 ( \13462 , \9266 , \12491 );
nand \U$4644 ( \13463 , \13461 , \13462 );
not \U$4645 ( \13464 , \13463 );
not \U$4646 ( \13465 , \8863 );
or \U$4647 ( \13466 , \9270 , \13465 );
buf \U$4648 ( \13467 , \8857 );
not \U$4649 ( \13468 , \13467 );
or \U$4650 ( \13469 , \9273 , \13468 );
not \U$4651 ( \13470 , \9495 );
and \U$4652 ( \13471 , \9297 , \13470 );
not \U$4653 ( \13472 , \10014 );
and \U$4654 ( \13473 , \9295 , \13472 );
nor \U$4655 ( \13474 , \13471 , \13473 );
nand \U$4656 ( \13475 , \13466 , \13469 , \13474 );
or \U$4657 ( \13476 , \11286 , \9002 );
not \U$4658 ( \13477 , \9213 );
or \U$4659 ( \13478 , \11291 , \13477 );
not \U$4660 ( \13479 , \9139 );
or \U$4661 ( \13480 , \11293 , \13479 );
nand \U$4662 ( \13481 , \9299 , \9351 );
and \U$4663 ( \13482 , \13476 , \13478 , \13480 , \13481 );
not \U$4664 ( \13483 , \13482 );
nor \U$4665 ( \13484 , \13475 , \13483 );
not \U$4666 ( \13485 , \9753 );
or \U$4667 ( \13486 , \9287 , \13485 );
not \U$4668 ( \13487 , \8928 );
or \U$4669 ( \13488 , \9290 , \13487 );
not \U$4670 ( \13489 , \9109 );
and \U$4671 ( \13490 , \9277 , \13489 );
not \U$4672 ( \13491 , \13286 );
and \U$4673 ( \13492 , \9281 , \13491 );
nor \U$4674 ( \13493 , \13490 , \13492 );
nand \U$4675 ( \13494 , \13486 , \13488 , \13493 );
not \U$4676 ( \13495 , \9307 );
or \U$4677 ( \13496 , \13495 , \13268 );
or \U$4678 ( \13497 , \9263 , \13295 );
nand \U$4679 ( \13498 , \13496 , \13497 );
nor \U$4680 ( \13499 , \13494 , \13498 );
nand \U$4681 ( \13500 , \13464 , \13484 , \13499 );
xnor \U$4682 ( \13501 , \13500 , \9327 );
not \U$4683 ( \13502 , \9444 );
or \U$4684 ( \13503 , \13502 , \13279 );
or \U$4685 ( \13504 , \9398 , \12491 );
nand \U$4686 ( \13505 , \13503 , \13504 );
not \U$4687 ( \13506 , \13505 );
nand \U$4688 ( \13507 , \9401 , \8981 );
nand \U$4689 ( \13508 , \9404 , \9978 );
not \U$4690 ( \13509 , \9844 );
and \U$4691 ( \13510 , \9430 , \13509 );
not \U$4692 ( \13511 , \9810 );
and \U$4693 ( \13512 , \9427 , \13511 );
nor \U$4694 ( \13513 , \13510 , \13512 );
nand \U$4695 ( \13514 , \13507 , \13508 , \13513 );
or \U$4696 ( \13515 , \11243 , \9423 );
nand \U$4697 ( \13516 , \9453 , \8886 );
nand \U$4698 ( \13517 , \9449 , \9411 );
nand \U$4699 ( \13518 , \9432 , \9351 );
and \U$4700 ( \13519 , \13515 , \13516 , \13517 , \13518 );
not \U$4701 ( \13520 , \13519 );
nor \U$4702 ( \13521 , \13514 , \13520 );
nand \U$4703 ( \13522 , \9418 , \9960 );
or \U$4704 ( \13523 , \9422 , \8929 );
not \U$4705 ( \13524 , \9177 );
and \U$4706 ( \13525 , \9409 , \13524 );
not \U$4707 ( \13526 , \9252 );
and \U$4708 ( \13527 , \9414 , \13526 );
nor \U$4709 ( \13528 , \13525 , \13527 );
nand \U$4710 ( \13529 , \13522 , \13523 , \13528 );
not \U$4711 ( \13530 , \9440 );
or \U$4712 ( \13531 , \13530 , \13268 );
or \U$4713 ( \13532 , \9395 , \13295 );
nand \U$4714 ( \13533 , \13531 , \13532 );
nor \U$4715 ( \13534 , \13529 , \13533 );
nand \U$4716 ( \13535 , \13506 , \13521 , \13534 );
xnor \U$4717 ( \13536 , \13535 , \9460 );
nor \U$4718 ( \13537 , \13501 , \13536 );
not \U$4719 ( \13538 , \9600 );
or \U$4720 ( \13539 , \13538 , \9252 );
not \U$4721 ( \13540 , \9108 );
or \U$4722 ( \13541 , \9597 , \13540 );
nand \U$4723 ( \13542 , \13539 , \13541 );
not \U$4724 ( \13543 , \13542 );
not \U$4725 ( \13544 , \9593 );
or \U$4726 ( \13545 , \13544 , \9015 );
or \U$4727 ( \13546 , \9588 , \9090 );
nand \U$4728 ( \13547 , \13545 , \13546 );
not \U$4729 ( \13548 , \13547 );
not \U$4730 ( \13549 , \9611 );
and \U$4731 ( \13550 , \13549 , \13334 );
not \U$4732 ( \13551 , \13281 );
and \U$4733 ( \13552 , \9613 , \13551 );
or \U$4734 ( \13553 , \9604 , \9206 );
or \U$4735 ( \13554 , \9607 , \8911 );
nand \U$4736 ( \13555 , \13553 , \13554 );
nor \U$4737 ( \13556 , \13550 , \13552 , \13555 );
and \U$4738 ( \13557 , \13543 , \13548 , \13556 );
not \U$4739 ( \13558 , \13557 );
and \U$4740 ( \13559 , \9622 , \8878 );
and \U$4741 ( \13560 , \9619 , \9213 );
or \U$4742 ( \13561 , \13559 , \13560 );
or \U$4743 ( \13562 , \9071 , \9632 );
or \U$4744 ( \13563 , \11314 , \8900 );
nand \U$4745 ( \13564 , \13562 , \13563 );
nor \U$4746 ( \13565 , \13561 , \13564 );
not \U$4747 ( \13566 , \9647 );
and \U$4748 ( \13567 , \13566 , \13269 );
not \U$4749 ( \13568 , \13295 );
and \U$4750 ( \13569 , \9643 , \13568 );
or \U$4751 ( \13570 , \9637 , \8864 );
or \U$4752 ( \13571 , \9640 , \10014 );
nand \U$4753 ( \13572 , \13570 , \13571 );
nor \U$4754 ( \13573 , \13567 , \13569 , \13572 );
nand \U$4755 ( \13574 , \13565 , \13573 );
nor \U$4756 ( \13575 , \13558 , \13574 );
xnor \U$4757 ( \13576 , RIb7af630_254, \13575 );
not \U$4758 ( \13577 , \9380 );
or \U$4759 ( \13578 , \13577 , \13279 );
or \U$4760 ( \13579 , \9335 , \13281 );
nand \U$4761 ( \13580 , \13578 , \13579 );
not \U$4762 ( \13581 , \13580 );
not \U$4763 ( \13582 , \8981 );
or \U$4764 ( \13583 , \9339 , \13582 );
buf \U$4765 ( \13584 , \8857 );
not \U$4766 ( \13585 , \13584 );
or \U$4767 ( \13586 , \9342 , \13585 );
not \U$4768 ( \13587 , \8911 );
and \U$4769 ( \13588 , \9364 , \13587 );
not \U$4770 ( \13589 , \9810 );
and \U$4771 ( \13590 , \9361 , \13589 );
nor \U$4772 ( \13591 , \13588 , \13590 );
nand \U$4773 ( \13592 , \13583 , \13586 , \13591 );
not \U$4774 ( \13593 , \9369 );
not \U$4775 ( \13594 , \9001 );
or \U$4776 ( \13595 , \13593 , \13594 );
nand \U$4777 ( \13596 , \9366 , \9351 );
not \U$4778 ( \13597 , \12874 );
and \U$4779 ( \13598 , \13597 , \9411 );
and \U$4780 ( \13599 , \9466 , \9377 );
nor \U$4781 ( \13600 , \13598 , \13599 );
nand \U$4782 ( \13601 , \13595 , \13596 , \13600 );
nor \U$4783 ( \13602 , \13592 , \13601 );
not \U$4784 ( \13603 , \9753 );
or \U$4785 ( \13604 , \9354 , \13603 );
not \U$4786 ( \13605 , \10028 );
or \U$4787 ( \13606 , \9357 , \13605 );
not \U$4788 ( \13607 , \13540 );
and \U$4789 ( \13608 , \9346 , \13607 );
not \U$4790 ( \13609 , \9036 );
and \U$4791 ( \13610 , \9348 , \13609 );
nor \U$4792 ( \13611 , \13608 , \13610 );
nand \U$4793 ( \13612 , \13604 , \13606 , \13611 );
not \U$4794 ( \13613 , \9374 );
or \U$4795 ( \13614 , \13613 , \13268 );
or \U$4796 ( \13615 , \9332 , \13295 );
nand \U$4797 ( \13616 , \13614 , \13615 );
nor \U$4798 ( \13617 , \13612 , \13616 );
nand \U$4799 ( \13618 , \13581 , \13602 , \13617 );
xnor \U$4800 ( \13619 , \13618 , \9392 );
nor \U$4801 ( \13620 , \13576 , \13619 );
and \U$4802 ( \13621 , \13459 , \13537 , \13620 );
or \U$4803 ( \13622 , \9948 , \9181 );
or \U$4804 ( \13623 , \13143 , \9109 );
nand \U$4805 ( \13624 , \13622 , \13623 );
not \U$4806 ( \13625 , \13624 );
not \U$4807 ( \13626 , \9954 );
or \U$4808 ( \13627 , \13626 , \9015 );
or \U$4809 ( \13628 , \9952 , \9090 );
nand \U$4810 ( \13629 , \13627 , \13628 );
not \U$4811 ( \13630 , \13629 );
and \U$4812 ( \13631 , \9936 , \13334 );
not \U$4813 ( \13632 , \13281 );
and \U$4814 ( \13633 , \9939 , \13632 );
or \U$4815 ( \13634 , \9930 , \9206 );
or \U$4816 ( \13635 , \9933 , \9495 );
nand \U$4817 ( \13636 , \13634 , \13635 );
nor \U$4818 ( \13637 , \13631 , \13633 , \13636 );
and \U$4819 ( \13638 , \13625 , \13630 , \13637 );
not \U$4820 ( \13639 , \13638 );
not \U$4821 ( \13640 , \9965 );
or \U$4822 ( \13641 , \13640 , \13325 );
or \U$4823 ( \13642 , \11618 , \9741 );
nand \U$4824 ( \13643 , \13641 , \13642 );
or \U$4825 ( \13644 , \9285 , \11623 );
or \U$4826 ( \13645 , \11625 , \8900 );
nand \U$4827 ( \13646 , \13644 , \13645 );
nor \U$4828 ( \13647 , \13643 , \13646 );
and \U$4829 ( \13648 , \9984 , \13269 );
not \U$4830 ( \13649 , \13295 );
and \U$4831 ( \13650 , \9982 , \13649 );
or \U$4832 ( \13651 , \11635 , \8864 );
or \U$4833 ( \13652 , \11629 , \8918 );
nand \U$4834 ( \13653 , \13651 , \13652 );
nor \U$4835 ( \13654 , \13648 , \13650 , \13653 );
nand \U$4836 ( \13655 , \13647 , \13654 );
nor \U$4837 ( \13656 , \13639 , \13655 );
xnor \U$4838 ( \13657 , \13656 , \9990 );
not \U$4839 ( \13658 , \9530 );
or \U$4840 ( \13659 , \13658 , \9824 );
or \U$4841 ( \13660 , \9527 , \9177 );
nand \U$4842 ( \13661 , \13659 , \13660 );
not \U$4843 ( \13662 , \13661 );
not \U$4844 ( \13663 , \9523 );
or \U$4845 ( \13664 , \13663 , \9234 );
or \U$4846 ( \13665 , \9519 , \9160 );
nand \U$4847 ( \13666 , \13664 , \13665 );
not \U$4848 ( \13667 , \13666 );
and \U$4849 ( \13668 , \9542 , \13334 );
not \U$4850 ( \13669 , \13281 );
and \U$4851 ( \13670 , \9545 , \13669 );
or \U$4852 ( \13671 , \9534 , \9206 );
or \U$4853 ( \13672 , \9537 , \9495 );
nand \U$4854 ( \13673 , \13671 , \13672 );
nor \U$4855 ( \13674 , \13668 , \13670 , \13673 );
and \U$4856 ( \13675 , \13662 , \13667 , \13674 );
not \U$4857 ( \13676 , \13675 );
not \U$4858 ( \13677 , \9554 );
or \U$4859 ( \13678 , \13677 , \9994 );
or \U$4860 ( \13679 , \9552 , \9741 );
nand \U$4861 ( \13680 , \13678 , \13679 );
or \U$4862 ( \13681 , \9071 , \9564 );
or \U$4863 ( \13682 , \11582 , \9002 );
nand \U$4864 ( \13683 , \13681 , \13682 );
nor \U$4865 ( \13684 , \13680 , \13683 );
and \U$4866 ( \13685 , \9578 , \13269 );
not \U$4867 ( \13686 , \13295 );
and \U$4868 ( \13687 , \9575 , \13686 );
or \U$4869 ( \13688 , \9569 , \8982 );
or \U$4870 ( \13689 , \9572 , \9702 );
nand \U$4871 ( \13690 , \13688 , \13689 );
nor \U$4872 ( \13691 , \13685 , \13687 , \13690 );
nand \U$4873 ( \13692 , \13684 , \13691 );
nor \U$4874 ( \13693 , \13676 , \13692 );
xnor \U$4875 ( \13694 , \13693 , \9585 );
or \U$4876 ( \13695 , \9997 , \9824 );
or \U$4877 ( \13696 , \11666 , \8950 );
nand \U$4878 ( \13697 , \13695 , \13696 );
not \U$4879 ( \13698 , \10004 );
or \U$4880 ( \13699 , \13698 , \8929 );
or \U$4881 ( \13700 , \10002 , \8924 );
nand \U$4882 ( \13701 , \13699 , \13700 );
nor \U$4883 ( \13702 , \13697 , \13701 );
and \U$4884 ( \13703 , \10017 , \13334 );
not \U$4885 ( \13704 , \13281 );
and \U$4886 ( \13705 , \10020 , \13704 );
or \U$4887 ( \13706 , \10010 , \9206 );
or \U$4888 ( \13707 , \10013 , \8911 );
nand \U$4889 ( \13708 , \13706 , \13707 );
nor \U$4890 ( \13709 , \13703 , \13705 , \13708 );
nand \U$4891 ( \13710 , \13702 , \13709 );
not \U$4892 ( \13711 , \10030 );
or \U$4893 ( \13712 , \13711 , \9412 );
or \U$4894 ( \13713 , \12230 , \9741 );
nand \U$4895 ( \13714 , \13712 , \13713 );
or \U$4896 ( \13715 , \9285 , \11693 );
or \U$4897 ( \13716 , \12235 , \9077 );
nand \U$4898 ( \13717 , \13715 , \13716 );
nor \U$4899 ( \13718 , \13714 , \13717 );
and \U$4900 ( \13719 , \10049 , \13269 );
not \U$4901 ( \13720 , \13295 );
and \U$4902 ( \13721 , \10047 , \13720 );
or \U$4903 ( \13722 , \11684 , \8982 );
or \U$4904 ( \13723 , \12222 , \8918 );
nand \U$4905 ( \13724 , \13722 , \13723 );
nor \U$4906 ( \13725 , \13719 , \13721 , \13724 );
nand \U$4907 ( \13726 , \13718 , \13725 );
nor \U$4908 ( \13727 , \13710 , \13726 );
xnor \U$4909 ( \13728 , RIb7af540_256, \13727 );
or \U$4910 ( \13729 , \12178 , \13286 );
or \U$4911 ( \13730 , \9868 , \9031 );
nand \U$4912 ( \13731 , \13729 , \13730 );
not \U$4913 ( \13732 , \13731 );
not \U$4914 ( \13733 , \9864 );
or \U$4915 ( \13734 , \13733 , \8929 );
or \U$4916 ( \13735 , \9860 , \9090 );
nand \U$4917 ( \13736 , \13734 , \13735 );
not \U$4918 ( \13737 , \13736 );
and \U$4919 ( \13738 , \9881 , \13334 );
not \U$4920 ( \13739 , \12491 );
and \U$4921 ( \13740 , \9886 , \13739 );
or \U$4922 ( \13741 , \9875 , \9206 );
or \U$4923 ( \13742 , \9878 , \8911 );
nand \U$4924 ( \13743 , \13741 , \13742 );
nor \U$4925 ( \13744 , \13738 , \13740 , \13743 );
and \U$4926 ( \13745 , \13732 , \13737 , \13744 );
not \U$4927 ( \13746 , \13745 );
not \U$4928 ( \13747 , \9897 );
not \U$4929 ( \13748 , \8878 );
or \U$4930 ( \13749 , \13747 , \13748 );
not \U$4931 ( \13750 , \8886 );
or \U$4932 ( \13751 , \9895 , \13750 );
nand \U$4933 ( \13752 , \13749 , \13751 );
or \U$4934 ( \13753 , \9071 , \9906 );
or \U$4935 ( \13754 , \11711 , \9221 );
nand \U$4936 ( \13755 , \13753 , \13754 );
nor \U$4937 ( \13756 , \13752 , \13755 );
and \U$4938 ( \13757 , \9920 , \13269 );
not \U$4939 ( \13758 , \13295 );
and \U$4940 ( \13759 , \9917 , \13758 );
or \U$4941 ( \13760 , \9911 , \8982 );
or \U$4942 ( \13761 , \9914 , \8918 );
nand \U$4943 ( \13762 , \13760 , \13761 );
nor \U$4944 ( \13763 , \13757 , \13759 , \13762 );
nand \U$4945 ( \13764 , \13756 , \13763 );
nor \U$4946 ( \13765 , \13746 , \13764 );
xnor \U$4947 ( \13766 , RIb7a0c48_261, \13765 );
nor \U$4948 ( \13767 , \13728 , \13766 );
nand \U$4949 ( \13768 , \13657 , \13694 , \13767 );
not \U$4950 ( \13769 , \9172 );
or \U$4951 ( \13770 , \13769 , \13279 );
or \U$4952 ( \13771 , \9125 , \13281 );
nand \U$4953 ( \13772 , \13770 , \13771 );
not \U$4954 ( \13773 , \13772 );
nand \U$4955 ( \13774 , \9129 , \13298 );
nand \U$4956 ( \13775 , \9132 , \9978 );
not \U$4957 ( \13776 , \9844 );
and \U$4958 ( \13777 , \9157 , \13776 );
not \U$4959 ( \13778 , \9810 );
and \U$4960 ( \13779 , \9155 , \13778 );
nor \U$4961 ( \13780 , \13777 , \13779 );
nand \U$4962 ( \13781 , \13774 , \13775 , \13780 );
or \U$4963 ( \13782 , \11424 , \9077 );
nand \U$4964 ( \13783 , \9180 , \9466 );
nand \U$4965 ( \13784 , \9176 , \8878 );
nand \U$4966 ( \13785 , \9159 , \9351 );
and \U$4967 ( \13786 , \13782 , \13783 , \13784 , \13785 );
not \U$4968 ( \13787 , \13786 );
nor \U$4969 ( \13788 , \13781 , \13787 );
nand \U$4970 ( \13789 , \9147 , \9688 );
or \U$4971 ( \13790 , \9151 , \9234 );
not \U$4972 ( \13791 , \9450 );
and \U$4973 ( \13792 , \9137 , \13791 );
not \U$4974 ( \13793 , \8956 );
and \U$4975 ( \13794 , \9142 , \13793 );
nor \U$4976 ( \13795 , \13792 , \13794 );
nand \U$4977 ( \13796 , \13789 , \13790 , \13795 );
not \U$4978 ( \13797 , \9168 );
or \U$4979 ( \13798 , \13797 , \13268 );
or \U$4980 ( \13799 , \9122 , \13295 );
nand \U$4981 ( \13800 , \13798 , \13799 );
nor \U$4982 ( \13801 , \13796 , \13800 );
nand \U$4983 ( \13802 , \13773 , \13788 , \13801 );
xnor \U$4984 ( \13803 , RIb7af6a8_253, \13802 );
not \U$4985 ( \13804 , \9102 );
or \U$4986 ( \13805 , \13804 , \13279 );
or \U$4987 ( \13806 , \9050 , \13281 );
nand \U$4988 ( \13807 , \13805 , \13806 );
not \U$4989 ( \13808 , \13807 );
not \U$4990 ( \13809 , \8981 );
or \U$4991 ( \13810 , \9055 , \13809 );
not \U$4992 ( \13811 , \13584 );
or \U$4993 ( \13812 , \9058 , \13811 );
not \U$4994 ( \13813 , \8911 );
and \U$4995 ( \13814 , \9085 , \13813 );
not \U$4996 ( \13815 , \10014 );
and \U$4997 ( \13816 , \9081 , \13815 );
nor \U$4998 ( \13817 , \13814 , \13816 );
nand \U$4999 ( \13818 , \13810 , \13812 , \13817 );
or \U$5000 ( \13819 , \11466 , \9077 );
not \U$5001 ( \13820 , \8886 );
or \U$5002 ( \13821 , \11471 , \13820 );
not \U$5003 ( \13822 , \9411 );
or \U$5004 ( \13823 , \11473 , \13822 );
nand \U$5005 ( \13824 , \9089 , \9351 );
and \U$5006 ( \13825 , \13819 , \13821 , \13823 , \13824 );
not \U$5007 ( \13826 , \13825 );
nor \U$5008 ( \13827 , \13818 , \13826 );
not \U$5009 ( \13828 , \9753 );
or \U$5010 ( \13829 , \9073 , \13828 );
not \U$5011 ( \13830 , \9757 );
or \U$5012 ( \13831 , \9076 , \13830 );
not \U$5013 ( \13832 , \9248 );
and \U$5014 ( \13833 , \9063 , \13832 );
not \U$5015 ( \13834 , \9824 );
and \U$5016 ( \13835 , \9067 , \13834 );
nor \U$5017 ( \13836 , \13833 , \13835 );
nand \U$5018 ( \13837 , \13829 , \13831 , \13836 );
not \U$5019 ( \13838 , \9098 );
or \U$5020 ( \13839 , \13838 , \13268 );
or \U$5021 ( \13840 , \9047 , \13295 );
nand \U$5022 ( \13841 , \13839 , \13840 );
nor \U$5023 ( \13842 , \13837 , \13841 );
nand \U$5024 ( \13843 , \13808 , \13827 , \13842 );
xnor \U$5025 ( \13844 , RIb7af720_252, \13843 );
or \U$5026 ( \13845 , \11494 , \13353 );
or \U$5027 ( \13846 , \9798 , \9760 );
nand \U$5028 ( \13847 , \13845 , \13846 );
not \U$5029 ( \13848 , \9794 );
or \U$5030 ( \13849 , \13848 , \9015 );
or \U$5031 ( \13850 , \9791 , \9160 );
nand \U$5032 ( \13851 , \13849 , \13850 );
nor \U$5033 ( \13852 , \13847 , \13851 );
not \U$5034 ( \13853 , \9814 );
and \U$5035 ( \13854 , \13853 , \13334 );
not \U$5036 ( \13855 , \13281 );
and \U$5037 ( \13856 , \9816 , \13855 );
or \U$5038 ( \13857 , \9806 , \9206 );
or \U$5039 ( \13858 , \9809 , \9844 );
nand \U$5040 ( \13859 , \13857 , \13858 );
nor \U$5041 ( \13860 , \13854 , \13856 , \13859 );
nand \U$5042 ( \13861 , \13852 , \13860 );
not \U$5043 ( \13862 , \9826 );
or \U$5044 ( \13863 , \13862 , \9065 );
or \U$5045 ( \13864 , \9823 , \8887 );
nand \U$5046 ( \13865 , \13863 , \13864 );
or \U$5047 ( \13866 , \9352 , \9834 );
or \U$5048 ( \13867 , \12311 , \9423 );
nand \U$5049 ( \13868 , \13866 , \13867 );
nor \U$5050 ( \13869 , \13865 , \13868 );
not \U$5051 ( \13870 , \9851 );
and \U$5052 ( \13871 , \13870 , \13269 );
not \U$5053 ( \13872 , \13295 );
and \U$5054 ( \13873 , \9847 , \13872 );
or \U$5055 ( \13874 , \9840 , \8982 );
or \U$5056 ( \13875 , \9843 , \9702 );
nand \U$5057 ( \13876 , \13874 , \13875 );
nor \U$5058 ( \13877 , \13871 , \13873 , \13876 );
nand \U$5059 ( \13878 , \13869 , \13877 );
nor \U$5060 ( \13879 , \13861 , \13878 );
xnor \U$5061 ( \13880 , RIb7a5bf8_260, \13879 );
not \U$5062 ( \13881 , \8940 );
or \U$5063 ( \13882 , \13881 , \13279 );
or \U$5064 ( \13883 , \8844 , \13281 );
nand \U$5065 ( \13884 , \13882 , \13883 );
not \U$5066 ( \13885 , \13884 );
nand \U$5067 ( \13886 , \8852 , \8863 );
nand \U$5068 ( \13887 , \8860 , \13584 );
not \U$5069 ( \13888 , \9495 );
and \U$5070 ( \13889 , \8915 , \13888 );
not \U$5071 ( \13890 , \9810 );
and \U$5072 ( \13891 , \8904 , \13890 );
nor \U$5073 ( \13892 , \13889 , \13891 );
nand \U$5074 ( \13893 , \13886 , \13887 , \13892 );
not \U$5075 ( \13894 , \8927 );
or \U$5076 ( \13895 , \13894 , \9423 );
nand \U$5077 ( \13896 , \8953 , \9213 );
nand \U$5078 ( \13897 , \8947 , \9139 );
nand \U$5079 ( \13898 , \8921 , \9351 );
and \U$5080 ( \13899 , \13895 , \13896 , \13897 , \13898 );
not \U$5081 ( \13900 , \13899 );
nor \U$5082 ( \13901 , \13893 , \13900 );
nand \U$5083 ( \13902 , \8893 , \9688 );
nand \U$5084 ( \13903 , \8896 , \10028 );
not \U$5085 ( \13904 , \10031 );
and \U$5086 ( \13905 , \8868 , \13904 );
not \U$5087 ( \13906 , \9036 );
and \U$5088 ( \13907 , \8881 , \13906 );
nor \U$5089 ( \13908 , \13905 , \13907 );
nand \U$5090 ( \13909 , \13902 , \13903 , \13908 );
not \U$5091 ( \13910 , \8934 );
or \U$5092 ( \13911 , \13910 , \13268 );
or \U$5093 ( \13912 , \8828 , \13295 );
nand \U$5094 ( \13913 , \13911 , \13912 );
nor \U$5095 ( \13914 , \13909 , \13913 );
nand \U$5096 ( \13915 , \13885 , \13901 , \13914 );
xnor \U$5097 ( \13916 , \13915 , \8964 );
nor \U$5098 ( \13917 , \13880 , \13916 );
nand \U$5099 ( \13918 , \13803 , \13844 , \13917 );
nor \U$5100 ( \13919 , \13768 , \13918 );
nand \U$5101 ( \13920 , \13304 , \13621 , \13919 );
nand \U$5102 ( \13921 , \13258 , \13920 );
or \U$5103 ( \13922 , \13247 , \13921 );
not \U$5104 ( \13923 , RIea91330_6888);
xnor \U$5105 ( \13924 , \13923 , \10065 );
not \U$5106 ( \13925 , \13924 );
not \U$5107 ( \13926 , \8837 );
not \U$5108 ( \13927 , \12453 );
nand \U$5109 ( \13928 , \13926 , \13927 );
nor \U$5110 ( \13929 , \13928 , \10937 , \8905 );
or \U$5111 ( \13930 , \13925 , \13929 );
not \U$5112 ( \13931 , \10065 );
or \U$5113 ( \13932 , \13923 , \13931 );
nand \U$5114 ( \13933 , \13930 , \13932 );
not \U$5115 ( \13934 , \13933 );
not \U$5116 ( \13935 , \13920 );
nand \U$5117 ( \13936 , \13934 , \13935 );
not \U$5118 ( \13937 , \13936 );
not \U$5119 ( \13938 , \13935 );
or \U$5120 ( \13939 , \13934 , \13938 );
not \U$5121 ( \13940 , \13939 );
or \U$5122 ( \13941 , \13937 , \13940 );
not \U$5123 ( \13942 , \13941 );
or \U$5124 ( \13943 , \10065 , \13942 );
not \U$5125 ( \13944 , \13935 );
and \U$5126 ( \13945 , \12495 , \13944 );
not \U$5127 ( \13946 , \13245 );
or \U$5128 ( \13947 , \12485 , \13946 );
not \U$5129 ( \13948 , \13947 );
nand \U$5130 ( \13949 , \13945 , \13948 );
not \U$5131 ( \13950 , RIe548ff0_6844);
not \U$5132 ( \13951 , \10928 );
and \U$5133 ( \13952 , \13950 , \13951 );
not \U$5134 ( \13953 , \8833 );
and \U$5135 ( \13954 , \13953 , \10928 );
or \U$5136 ( \13955 , \13952 , \13954 );
nand \U$5137 ( \13956 , \13955 , \8875 );
not \U$5138 ( \13957 , \13956 );
not \U$5139 ( \13958 , \13244 );
or \U$5140 ( \13959 , \13935 , \13958 );
not \U$5141 ( \13960 , \13959 );
buf \U$5142 ( \13961 , RIea91330_6888);
buf \U$5143 ( \13962 , \13253 );
buf \U$5144 ( \13963 , \12456 );
buf \U$5145 ( \13964 , \12458 );
not \U$5146 ( \13965 , \13964 );
not \U$5147 ( \13966 , \13965 );
and \U$5148 ( \13967 , \13963 , \13966 );
or \U$5149 ( \13968 , \13962 , \13967 );
and \U$5150 ( \13969 , \13961 , \13968 );
buf \U$5151 ( \13970 , \13969 );
not \U$5152 ( \13971 , \13970 );
buf \U$5153 ( \13972 , \10937 );
not \U$5154 ( \13973 , \13972 );
buf \U$5155 ( \13974 , \13965 );
not \U$5156 ( \13975 , \13974 );
nand \U$5157 ( \13976 , \13973 , \13975 );
xor \U$5158 ( \13977 , \13963 , \13966 );
buf \U$5159 ( \13978 , \13977 );
not \U$5160 ( \13979 , \13978 );
xnor \U$5161 ( \13980 , \13962 , \13967 );
buf \U$5162 ( \13981 , \13980 );
not \U$5163 ( \13982 , \13981 );
nand \U$5164 ( \13983 , \13979 , \13982 );
or \U$5165 ( \13984 , \13976 , \13983 );
xor \U$5166 ( \13985 , \13961 , \13968 );
buf \U$5167 ( \13986 , \13985 );
nand \U$5168 ( \13987 , \13984 , \13986 );
nand \U$5169 ( \13988 , \13971 , \13987 );
not \U$5170 ( \13989 , \13988 );
not \U$5171 ( \13990 , \8905 );
or \U$5172 ( \13991 , \10937 , \13990 );
xor \U$5173 ( \13992 , \10928 , \8830 );
and \U$5174 ( \13993 , \13992 , \13956 );
not \U$5175 ( \13994 , \13993 );
or \U$5176 ( \13995 , \13991 , \13994 );
or \U$5177 ( \13996 , \9492 , \13995 );
not \U$5178 ( \13997 , \13993 );
or \U$5179 ( \13998 , \10917 , \13997 );
or \U$5180 ( \13999 , \9494 , \13998 );
nand \U$5181 ( \14000 , \13996 , \13999 );
not \U$5182 ( \14001 , \13956 );
or \U$5183 ( \14002 , \13992 , \14001 );
not \U$5184 ( \14003 , \14002 );
not \U$5185 ( \14004 , \14003 );
or \U$5186 ( \14005 , \10922 , \14004 );
or \U$5187 ( \14006 , \9498 , \14005 );
not \U$5188 ( \14007 , \8835 );
or \U$5189 ( \14008 , \8905 , \14007 );
not \U$5190 ( \14009 , \14003 );
or \U$5191 ( \14010 , \14008 , \14009 );
not \U$5192 ( \14011 , \14010 );
not \U$5193 ( \14012 , \14011 );
or \U$5194 ( \14013 , \9500 , \14012 );
nand \U$5195 ( \14014 , \14006 , \14013 );
nor \U$5196 ( \14015 , \14000 , \14014 );
not \U$5197 ( \14016 , \14003 );
or \U$5198 ( \14017 , \10917 , \14016 );
not \U$5199 ( \14018 , \14017 );
not \U$5200 ( \14019 , \9506 );
and \U$5201 ( \14020 , \14018 , \14019 );
not \U$5202 ( \14021 , \13956 );
and \U$5203 ( \14022 , \14021 , \13992 );
not \U$5204 ( \14023 , \14022 );
or \U$5205 ( \14024 , \10922 , \14023 );
not \U$5206 ( \14025 , \14024 );
nand \U$5207 ( \14026 , \14025 , \10976 );
not \U$5208 ( \14027 , \14026 );
not \U$5209 ( \14028 , \14021 );
or \U$5210 ( \14029 , \13992 , \14028 );
not \U$5211 ( \14030 , \14029 );
not \U$5212 ( \14031 , \14030 );
or \U$5213 ( \14032 , \13991 , \14031 );
not \U$5214 ( \14033 , \14032 );
not \U$5215 ( \14034 , \14033 );
or \U$5216 ( \14035 , \9509 , \14034 );
not \U$5217 ( \14036 , \14030 );
or \U$5218 ( \14037 , \14008 , \14036 );
not \U$5219 ( \14038 , \14037 );
not \U$5220 ( \14039 , \14038 );
or \U$5221 ( \14040 , \9511 , \14039 );
nand \U$5222 ( \14041 , \14035 , \14040 );
nor \U$5223 ( \14042 , \14020 , \14027 , \14041 );
not \U$5224 ( \14043 , \14022 );
or \U$5225 ( \14044 , \10917 , \14043 );
not \U$5226 ( \14045 , \14044 );
nand \U$5227 ( \14046 , \14045 , \9476 );
not \U$5228 ( \14047 , \14022 );
or \U$5229 ( \14048 , \13991 , \14047 );
not \U$5230 ( \14049 , \14048 );
nand \U$5231 ( \14050 , \14049 , \9472 );
not \U$5232 ( \14051 , \9467 );
not \U$5233 ( \14052 , \14030 );
or \U$5234 ( \14053 , \10922 , \14052 );
not \U$5235 ( \14054 , \14053 );
and \U$5236 ( \14055 , \14051 , \14054 );
not \U$5237 ( \14056 , \14030 );
or \U$5238 ( \14057 , \10917 , \14056 );
not \U$5239 ( \14058 , \14057 );
and \U$5240 ( \14059 , \14058 , \10986 );
nor \U$5241 ( \14060 , \14055 , \14059 );
nand \U$5242 ( \14061 , \14046 , \14050 , \14060 );
not \U$5243 ( \14062 , \13993 );
or \U$5244 ( \14063 , \14008 , \14062 );
not \U$5245 ( \14064 , \14063 );
not \U$5246 ( \14065 , \14064 );
not \U$5247 ( \14066 , \14065 );
and \U$5248 ( \14067 , \10163 , \14066 );
not \U$5249 ( \14068 , \13993 );
or \U$5250 ( \14069 , \10922 , \14068 );
not \U$5251 ( \14070 , \14069 );
and \U$5252 ( \14071 , \10168 , \14070 );
nor \U$5253 ( \14072 , \14067 , \14071 );
not \U$5254 ( \14073 , \9480 );
not \U$5255 ( \14074 , \14003 );
or \U$5256 ( \14075 , \13991 , \14074 );
not \U$5257 ( \14076 , \14075 );
and \U$5258 ( \14077 , \14073 , \14076 );
not \U$5259 ( \14078 , \14022 );
or \U$5260 ( \14079 , \14078 , \14008 );
not \U$5261 ( \14080 , \14079 );
and \U$5262 ( \14081 , \14080 , \12557 );
nor \U$5263 ( \14082 , \14077 , \14081 );
nand \U$5264 ( \14083 , \14072 , \14082 );
nor \U$5265 ( \14084 , \14061 , \14083 );
nand \U$5266 ( \14085 , \14015 , \14042 , \14084 );
not \U$5267 ( \14086 , \14085 );
nand \U$5268 ( \14087 , \14045 , \9364 );
nand \U$5269 ( \14088 , \14025 , \9341 );
nand \U$5270 ( \14089 , \14087 , \14088 );
not \U$5271 ( \14090 , \14089 );
not \U$5272 ( \14091 , \14075 );
nand \U$5273 ( \14092 , \9380 , \14091 );
nand \U$5274 ( \14093 , \14080 , \9334 );
and \U$5275 ( \14094 , \14090 , \14092 , \14093 );
or \U$5276 ( \14095 , \13593 , \14012 );
not \U$5277 ( \14096 , \13993 );
or \U$5278 ( \14097 , \13991 , \14096 );
or \U$5279 ( \14098 , \11365 , \14097 );
nand \U$5280 ( \14099 , \14095 , \14098 );
not \U$5281 ( \14100 , \14003 );
or \U$5282 ( \14101 , \10917 , \14100 );
or \U$5283 ( \14102 , \12874 , \14101 );
not \U$5284 ( \14103 , \14003 );
or \U$5285 ( \14104 , \10922 , \14103 );
or \U$5286 ( \14105 , \11371 , \14104 );
nand \U$5287 ( \14106 , \14102 , \14105 );
nor \U$5288 ( \14107 , \14099 , \14106 );
not \U$5289 ( \14108 , \14048 );
nand \U$5290 ( \14109 , \14108 , \9353 );
nand \U$5291 ( \14110 , \9356 , \14038 );
and \U$5292 ( \14111 , \14058 , \9346 );
not \U$5293 ( \14112 , \14053 );
and \U$5294 ( \14113 , \9348 , \14112 );
nor \U$5295 ( \14114 , \14111 , \14113 );
nand \U$5296 ( \14115 , \14109 , \14110 , \14114 );
not \U$5297 ( \14116 , \13993 );
or \U$5298 ( \14117 , \10922 , \14116 );
not \U$5299 ( \14118 , \14117 );
and \U$5300 ( \14119 , \9338 , \14118 );
not \U$5301 ( \14120 , \13993 );
or \U$5302 ( \14121 , \10917 , \14120 );
not \U$5303 ( \14122 , \14121 );
and \U$5304 ( \14123 , \9361 , \14122 );
nor \U$5305 ( \14124 , \14119 , \14123 );
not \U$5306 ( \14125 , \14032 );
and \U$5307 ( \14126 , \9374 , \14125 );
not \U$5308 ( \14127 , \14063 );
and \U$5309 ( \14128 , \9331 , \14127 );
nor \U$5310 ( \14129 , \14126 , \14128 );
nand \U$5311 ( \14130 , \14124 , \14129 );
nor \U$5312 ( \14131 , \14115 , \14130 );
nand \U$5313 ( \14132 , \14094 , \14107 , \14131 );
xnor \U$5314 ( \14133 , RIb7b9608_246, \14132 );
not \U$5315 ( \14134 , \14003 );
or \U$5316 ( \14135 , \10922 , \14134 );
or \U$5317 ( \14136 , \9620 , \14135 );
not \U$5318 ( \14137 , \14003 );
or \U$5319 ( \14138 , \10917 , \14137 );
or \U$5320 ( \14139 , \9625 , \14138 );
nand \U$5321 ( \14140 , \14136 , \14139 );
not \U$5322 ( \14141 , \9628 );
or \U$5323 ( \14142 , \14141 , \14012 );
or \U$5324 ( \14143 , \9632 , \13995 );
nand \U$5325 ( \14144 , \14142 , \14143 );
nor \U$5326 ( \14145 , \14140 , \14144 );
or \U$5327 ( \14146 , \9637 , \14069 );
or \U$5328 ( \14147 , \9640 , \13998 );
nand \U$5329 ( \14148 , \14146 , \14147 );
or \U$5330 ( \14149 , \9647 , \14032 );
or \U$5331 ( \14150 , \11322 , \14065 );
nand \U$5332 ( \14151 , \14149 , \14150 );
nor \U$5333 ( \14152 , \14148 , \14151 );
nand \U$5334 ( \14153 , \14108 , \9587 );
not \U$5335 ( \14154 , \14038 );
or \U$5336 ( \14155 , \12108 , \14154 );
not \U$5337 ( \14156 , \13538 );
and \U$5338 ( \14157 , \14156 , \14112 );
and \U$5339 ( \14158 , \14058 , \9596 );
nor \U$5340 ( \14159 , \14157 , \14158 );
nand \U$5341 ( \14160 , \14153 , \14155 , \14159 );
not \U$5342 ( \14161 , \14080 );
or \U$5343 ( \14162 , \9614 , \14161 );
nand \U$5344 ( \14163 , \14025 , \9603 );
nand \U$5345 ( \14164 , \14045 , \9606 );
not \U$5346 ( \14165 , \14091 );
or \U$5347 ( \14166 , \9611 , \14165 );
and \U$5348 ( \14167 , \14162 , \14163 , \14164 , \14166 );
not \U$5349 ( \14168 , \14167 );
nor \U$5350 ( \14169 , \14160 , \14168 );
nand \U$5351 ( \14170 , \14145 , \14152 , \14169 );
xnor \U$5352 ( \14171 , RIb7af630_254, \14170 );
nand \U$5353 ( \14172 , \14045 , \9297 );
nand \U$5354 ( \14173 , \14025 , \9272 );
nand \U$5355 ( \14174 , \14172 , \14173 );
not \U$5356 ( \14175 , \14174 );
not \U$5357 ( \14176 , \14076 );
or \U$5358 ( \14177 , \10415 , \14176 );
nand \U$5359 ( \14178 , \14080 , \9265 );
and \U$5360 ( \14179 , \14175 , \14177 , \14178 );
not \U$5361 ( \14180 , \14011 );
or \U$5362 ( \14181 , \11286 , \14180 );
not \U$5363 ( \14182 , \13993 );
or \U$5364 ( \14183 , \13991 , \14182 );
or \U$5365 ( \14184 , \11288 , \14183 );
nand \U$5366 ( \14185 , \14181 , \14184 );
or \U$5367 ( \14186 , \11293 , \14017 );
or \U$5368 ( \14187 , \11291 , \14135 );
nand \U$5369 ( \14188 , \14186 , \14187 );
nor \U$5370 ( \14189 , \14185 , \14188 );
nand \U$5371 ( \14190 , \14108 , \9286 );
nand \U$5372 ( \14191 , \9289 , \14038 );
and \U$5373 ( \14192 , \14058 , \9277 );
and \U$5374 ( \14193 , \9281 , \14112 );
nor \U$5375 ( \14194 , \14192 , \14193 );
nand \U$5376 ( \14195 , \14190 , \14191 , \14194 );
not \U$5377 ( \14196 , \13993 );
or \U$5378 ( \14197 , \10922 , \14196 );
not \U$5379 ( \14198 , \14197 );
and \U$5380 ( \14199 , \9269 , \14198 );
not \U$5381 ( \14200 , \13993 );
or \U$5382 ( \14201 , \10917 , \14200 );
not \U$5383 ( \14202 , \14201 );
and \U$5384 ( \14203 , \9295 , \14202 );
nor \U$5385 ( \14204 , \14199 , \14203 );
and \U$5386 ( \14205 , \9307 , \14125 );
not \U$5387 ( \14206 , \14065 );
and \U$5388 ( \14207 , \9262 , \14206 );
nor \U$5389 ( \14208 , \14205 , \14207 );
nand \U$5390 ( \14209 , \14204 , \14208 );
nor \U$5391 ( \14210 , \14195 , \14209 );
nand \U$5392 ( \14211 , \14179 , \14189 , \14210 );
xnor \U$5393 ( \14212 , \14211 , \9327 );
nand \U$5394 ( \14213 , \14045 , \9430 );
nand \U$5395 ( \14214 , \14025 , \9404 );
nand \U$5396 ( \14215 , \14213 , \14214 );
not \U$5397 ( \14216 , \14215 );
not \U$5398 ( \14217 , \14091 );
or \U$5399 ( \14218 , \10462 , \14217 );
nand \U$5400 ( \14219 , \14080 , \9397 );
and \U$5401 ( \14220 , \14216 , \14218 , \14219 );
or \U$5402 ( \14221 , \11243 , \14012 );
or \U$5403 ( \14222 , \11245 , \13995 );
nand \U$5404 ( \14223 , \14221 , \14222 );
or \U$5405 ( \14224 , \11250 , \14138 );
or \U$5406 ( \14225 , \11248 , \14005 );
nand \U$5407 ( \14226 , \14224 , \14225 );
nor \U$5408 ( \14227 , \14223 , \14226 );
nand \U$5409 ( \14228 , \14108 , \9418 );
nand \U$5410 ( \14229 , \9421 , \14038 );
and \U$5411 ( \14230 , \14058 , \9409 );
and \U$5412 ( \14231 , \9414 , \14112 );
nor \U$5413 ( \14232 , \14230 , \14231 );
nand \U$5414 ( \14233 , \14228 , \14229 , \14232 );
not \U$5415 ( \14234 , \14069 );
and \U$5416 ( \14235 , \9401 , \14234 );
not \U$5417 ( \14236 , \13998 );
and \U$5418 ( \14237 , \9427 , \14236 );
nor \U$5419 ( \14238 , \14235 , \14237 );
and \U$5420 ( \14239 , \9440 , \14033 );
not \U$5421 ( \14240 , \14065 );
and \U$5422 ( \14241 , \9394 , \14240 );
nor \U$5423 ( \14242 , \14239 , \14241 );
nand \U$5424 ( \14243 , \14238 , \14242 );
nor \U$5425 ( \14244 , \14233 , \14243 );
nand \U$5426 ( \14245 , \14220 , \14227 , \14244 );
xnor \U$5427 ( \14246 , \14245 , \9460 );
nor \U$5428 ( \14247 , \14212 , \14246 );
nand \U$5429 ( \14248 , \14133 , \14171 , \14247 );
not \U$5430 ( \14249 , \14248 );
or \U$5431 ( \14250 , \10244 , \14075 );
or \U$5432 ( \14251 , \11145 , \14079 );
nand \U$5433 ( \14252 , \14250 , \14251 );
not \U$5434 ( \14253 , \14252 );
nand \U$5435 ( \14254 , \14045 , \9701 );
nand \U$5436 ( \14255 , \14025 , \9706 );
and \U$5437 ( \14256 , \14253 , \14254 , \14255 );
or \U$5438 ( \14257 , \10248 , \14005 );
or \U$5439 ( \14258 , \10250 , \14101 );
nand \U$5440 ( \14259 , \14257 , \14258 );
not \U$5441 ( \14260 , \9690 );
or \U$5442 ( \14261 , \14260 , \14180 );
or \U$5443 ( \14262 , \11152 , \14097 );
nand \U$5444 ( \14263 , \14261 , \14262 );
nor \U$5445 ( \14264 , \14259 , \14263 );
nand \U$5446 ( \14265 , \14108 , \9679 );
nand \U$5447 ( \14266 , \9682 , \14038 );
and \U$5448 ( \14267 , \14058 , \9672 );
and \U$5449 ( \14268 , \9675 , \14112 );
nor \U$5450 ( \14269 , \14267 , \14268 );
nand \U$5451 ( \14270 , \14265 , \14266 , \14269 );
nand \U$5452 ( \14271 , \9667 , \14033 );
not \U$5453 ( \14272 , \14065 );
nand \U$5454 ( \14273 , \9664 , \14272 );
not \U$5455 ( \14274 , \14121 );
and \U$5456 ( \14275 , \9660 , \14274 );
not \U$5457 ( \14276 , \14117 );
and \U$5458 ( \14277 , \9656 , \14276 );
nor \U$5459 ( \14278 , \14275 , \14277 );
nand \U$5460 ( \14279 , \14271 , \14273 , \14278 );
nor \U$5461 ( \14280 , \14270 , \14279 );
nand \U$5462 ( \14281 , \14256 , \14264 , \14280 );
xnor \U$5463 ( \14282 , \14281 , \9719 );
or \U$5464 ( \14283 , \10188 , \14075 );
or \U$5465 ( \14284 , \11186 , \14079 );
nand \U$5466 ( \14285 , \14283 , \14284 );
not \U$5467 ( \14286 , \14285 );
nand \U$5468 ( \14287 , \14045 , \9769 );
nand \U$5469 ( \14288 , \14025 , \9772 );
and \U$5470 ( \14289 , \14286 , \14287 , \14288 );
or \U$5471 ( \14290 , \10194 , \14104 );
or \U$5472 ( \14291 , \10197 , \14017 );
nand \U$5473 ( \14292 , \14290 , \14291 );
not \U$5474 ( \14293 , \9755 );
or \U$5475 ( \14294 , \14293 , \14180 );
or \U$5476 ( \14295 , \11193 , \14183 );
nand \U$5477 ( \14296 , \14294 , \14295 );
nor \U$5478 ( \14297 , \14292 , \14296 );
nand \U$5479 ( \14298 , \14108 , \9744 );
nand \U$5480 ( \14299 , \9747 , \14038 );
and \U$5481 ( \14300 , \14058 , \9736 );
and \U$5482 ( \14301 , \9739 , \14112 );
nor \U$5483 ( \14302 , \14300 , \14301 );
nand \U$5484 ( \14303 , \14298 , \14299 , \14302 );
nand \U$5485 ( \14304 , \9731 , \14125 );
nand \U$5486 ( \14305 , \9728 , \14272 );
not \U$5487 ( \14306 , \14201 );
and \U$5488 ( \14307 , \9724 , \14306 );
not \U$5489 ( \14308 , \14197 );
and \U$5490 ( \14309 , \9721 , \14308 );
nor \U$5491 ( \14310 , \14307 , \14309 );
nand \U$5492 ( \14311 , \14304 , \14305 , \14310 );
nor \U$5493 ( \14312 , \14303 , \14311 );
nand \U$5494 ( \14313 , \14289 , \14297 , \14312 );
xnor \U$5495 ( \14314 , \14313 , \9786 );
nor \U$5496 ( \14315 , \14282 , \14314 );
nand \U$5497 ( \14316 , \14045 , \9228 );
nand \U$5498 ( \14317 , \14025 , \9200 );
nand \U$5499 ( \14318 , \14316 , \14317 );
not \U$5500 ( \14319 , \14318 );
not \U$5501 ( \14320 , \14091 );
or \U$5502 ( \14321 , \10323 , \14320 );
nand \U$5503 ( \14322 , \14080 , \9193 );
and \U$5504 ( \14323 , \14319 , \14321 , \14322 );
or \U$5505 ( \14324 , \11111 , \14180 );
or \U$5506 ( \14325 , \11113 , \13995 );
nand \U$5507 ( \14326 , \14324 , \14325 );
or \U$5508 ( \14327 , \11120 , \14138 );
or \U$5509 ( \14328 , \11117 , \14005 );
nand \U$5510 ( \14329 , \14327 , \14328 );
nor \U$5511 ( \14330 , \14326 , \14329 );
nand \U$5512 ( \14331 , \14108 , \9216 );
nand \U$5513 ( \14332 , \9219 , \14038 );
and \U$5514 ( \14333 , \14058 , \9210 );
and \U$5515 ( \14334 , \9212 , \14112 );
nor \U$5516 ( \14335 , \14333 , \14334 );
nand \U$5517 ( \14336 , \14331 , \14332 , \14335 );
not \U$5518 ( \14337 , \14069 );
and \U$5519 ( \14338 , \9204 , \14337 );
not \U$5520 ( \14339 , \13998 );
and \U$5521 ( \14340 , \9225 , \14339 );
nor \U$5522 ( \14341 , \14338 , \14340 );
and \U$5523 ( \14342 , \9239 , \14033 );
not \U$5524 ( \14343 , \14063 );
and \U$5525 ( \14344 , \9196 , \14343 );
nor \U$5526 ( \14345 , \14342 , \14344 );
nand \U$5527 ( \14346 , \14341 , \14345 );
nor \U$5528 ( \14347 , \14336 , \14346 );
nand \U$5529 ( \14348 , \14323 , \14330 , \14347 );
xnor \U$5530 ( \14349 , \14348 , \9260 );
nand \U$5531 ( \14350 , \14045 , \9009 );
nand \U$5532 ( \14351 , \14025 , \8979 );
nand \U$5533 ( \14352 , \14350 , \14351 );
not \U$5534 ( \14353 , \14352 );
nand \U$5535 ( \14354 , \9025 , \14091 );
nand \U$5536 ( \14355 , \14080 , \8970 );
and \U$5537 ( \14356 , \14353 , \14354 , \14355 );
or \U$5538 ( \14357 , \11058 , \14180 );
or \U$5539 ( \14358 , \11060 , \14097 );
nand \U$5540 ( \14359 , \14357 , \14358 );
or \U$5541 ( \14360 , \11067 , \14101 );
or \U$5542 ( \14361 , \11064 , \14104 );
nand \U$5543 ( \14362 , \14360 , \14361 );
nor \U$5544 ( \14363 , \14359 , \14362 );
nand \U$5545 ( \14364 , \14108 , \8996 );
nand \U$5546 ( \14365 , \8999 , \14038 );
and \U$5547 ( \14366 , \14058 , \8986 );
and \U$5548 ( \14367 , \8990 , \14112 );
nor \U$5549 ( \14368 , \14366 , \14367 );
nand \U$5550 ( \14369 , \14364 , \14365 , \14368 );
not \U$5551 ( \14370 , \14117 );
and \U$5552 ( \14371 , \8976 , \14370 );
not \U$5553 ( \14372 , \14121 );
and \U$5554 ( \14373 , \9006 , \14372 );
nor \U$5555 ( \14374 , \14371 , \14373 );
and \U$5556 ( \14375 , \9020 , \14033 );
not \U$5557 ( \14376 , \14063 );
and \U$5558 ( \14377 , \8966 , \14376 );
nor \U$5559 ( \14378 , \14375 , \14377 );
nand \U$5560 ( \14379 , \14374 , \14378 );
nor \U$5561 ( \14380 , \14369 , \14379 );
nand \U$5562 ( \14381 , \14356 , \14363 , \14380 );
xnor \U$5563 ( \14382 , \14381 , \9044 );
nor \U$5564 ( \14383 , \14349 , \14382 );
and \U$5565 ( \14384 , \14249 , \14315 , \14383 );
or \U$5566 ( \14385 , \11618 , \14104 );
or \U$5567 ( \14386 , \11620 , \14017 );
nand \U$5568 ( \14387 , \14385 , \14386 );
not \U$5569 ( \14388 , \10709 );
or \U$5570 ( \14389 , \14388 , \14012 );
or \U$5571 ( \14390 , \11623 , \14183 );
nand \U$5572 ( \14391 , \14389 , \14390 );
nor \U$5573 ( \14392 , \14387 , \14391 );
or \U$5574 ( \14393 , \11635 , \14117 );
or \U$5575 ( \14394 , \11629 , \14121 );
nand \U$5576 ( \14395 , \14393 , \14394 );
or \U$5577 ( \14396 , \12282 , \14032 );
or \U$5578 ( \14397 , \11633 , \14065 );
nand \U$5579 ( \14398 , \14396 , \14397 );
nor \U$5580 ( \14399 , \14395 , \14398 );
nand \U$5581 ( \14400 , \14049 , \9951 );
not \U$5582 ( \14401 , \14038 );
or \U$5583 ( \14402 , \9955 , \14401 );
not \U$5584 ( \14403 , \9948 );
and \U$5585 ( \14404 , \14403 , \14054 );
and \U$5586 ( \14405 , \14058 , \9944 );
nor \U$5587 ( \14406 , \14404 , \14405 );
nand \U$5588 ( \14407 , \14400 , \14402 , \14406 );
or \U$5589 ( \14408 , \9940 , \14161 );
nand \U$5590 ( \14409 , \14025 , \9929 );
nand \U$5591 ( \14410 , \14045 , \9932 );
not \U$5592 ( \14411 , \14076 );
or \U$5593 ( \14412 , \9937 , \14411 );
and \U$5594 ( \14413 , \14408 , \14409 , \14410 , \14412 );
not \U$5595 ( \14414 , \14413 );
nor \U$5596 ( \14415 , \14407 , \14414 );
nand \U$5597 ( \14416 , \14392 , \14399 , \14415 );
xnor \U$5598 ( \14417 , RIb7af450_258, \14416 );
or \U$5599 ( \14418 , \9552 , \14005 );
or \U$5600 ( \14419 , \9557 , \14101 );
nand \U$5601 ( \14420 , \14418 , \14419 );
not \U$5602 ( \14421 , \9560 );
or \U$5603 ( \14422 , \14421 , \14012 );
or \U$5604 ( \14423 , \9564 , \14097 );
nand \U$5605 ( \14424 , \14422 , \14423 );
nor \U$5606 ( \14425 , \14420 , \14424 );
or \U$5607 ( \14426 , \9569 , \14197 );
or \U$5608 ( \14427 , \9572 , \14201 );
nand \U$5609 ( \14428 , \14426 , \14427 );
or \U$5610 ( \14429 , \9579 , \14032 );
or \U$5611 ( \14430 , \11589 , \14065 );
nand \U$5612 ( \14431 , \14429 , \14430 );
nor \U$5613 ( \14432 , \14428 , \14431 );
nand \U$5614 ( \14433 , \14049 , \9518 );
not \U$5615 ( \14434 , \9523 );
not \U$5616 ( \14435 , \14038 );
or \U$5617 ( \14436 , \14434 , \14435 );
not \U$5618 ( \14437 , \13658 );
and \U$5619 ( \14438 , \14437 , \14054 );
and \U$5620 ( \14439 , \14058 , \9526 );
nor \U$5621 ( \14440 , \14438 , \14439 );
nand \U$5622 ( \14441 , \14433 , \14436 , \14440 );
or \U$5623 ( \14442 , \9546 , \14161 );
nand \U$5624 ( \14443 , \14025 , \9533 );
nand \U$5625 ( \14444 , \14045 , \9536 );
not \U$5626 ( \14445 , \14091 );
or \U$5627 ( \14446 , \9543 , \14445 );
and \U$5628 ( \14447 , \14442 , \14443 , \14444 , \14446 );
not \U$5629 ( \14448 , \14447 );
nor \U$5630 ( \14449 , \14441 , \14448 );
nand \U$5631 ( \14450 , \14425 , \14432 , \14449 );
xnor \U$5632 ( \14451 , RIb7af3d8_259, \14450 );
not \U$5633 ( \14452 , \14125 );
or \U$5634 ( \14453 , \11674 , \14452 );
not \U$5635 ( \14454 , \14272 );
or \U$5636 ( \14455 , \11681 , \14454 );
not \U$5637 ( \14456 , \14201 );
and \U$5638 ( \14457 , \10041 , \14456 );
not \U$5639 ( \14458 , \14197 );
and \U$5640 ( \14459 , \10043 , \14458 );
nor \U$5641 ( \14460 , \14457 , \14459 );
nand \U$5642 ( \14461 , \14453 , \14455 , \14460 );
not \U$5643 ( \14462 , \14461 );
or \U$5644 ( \14463 , \12230 , \14135 );
or \U$5645 ( \14464 , \11698 , \14138 );
nand \U$5646 ( \14465 , \14463 , \14464 );
not \U$5647 ( \14466 , \10027 );
or \U$5648 ( \14467 , \14466 , \14012 );
or \U$5649 ( \14468 , \11693 , \13995 );
nand \U$5650 ( \14469 , \14467 , \14468 );
nor \U$5651 ( \14470 , \14465 , \14469 );
or \U$5652 ( \14471 , \10021 , \14161 );
nand \U$5653 ( \14472 , \14025 , \10009 );
nand \U$5654 ( \14473 , \14045 , \10012 );
nand \U$5655 ( \14474 , \10017 , \14076 );
and \U$5656 ( \14475 , \14471 , \14472 , \14473 , \14474 );
not \U$5657 ( \14476 , \14475 );
not \U$5658 ( \14477 , \14476 );
not \U$5659 ( \14478 , \9997 );
and \U$5660 ( \14479 , \14478 , \14112 );
and \U$5661 ( \14480 , \14058 , \9992 );
nor \U$5662 ( \14481 , \14479 , \14480 );
not \U$5663 ( \14482 , \10002 );
and \U$5664 ( \14483 , \14482 , \14108 );
and \U$5665 ( \14484 , \14038 , \10004 );
nor \U$5666 ( \14485 , \14483 , \14484 );
and \U$5667 ( \14486 , \14477 , \14481 , \14485 );
nand \U$5668 ( \14487 , \14462 , \14470 , \14486 );
xnor \U$5669 ( \14488 , \14487 , \10055 );
or \U$5670 ( \14489 , \9895 , \14005 );
or \U$5671 ( \14490 , \9898 , \14101 );
nand \U$5672 ( \14491 , \14489 , \14490 );
not \U$5673 ( \14492 , \9902 );
or \U$5674 ( \14493 , \14492 , \14012 );
or \U$5675 ( \14494 , \9906 , \14097 );
nand \U$5676 ( \14495 , \14493 , \14494 );
nor \U$5677 ( \14496 , \14491 , \14495 );
or \U$5678 ( \14497 , \9911 , \14069 );
or \U$5679 ( \14498 , \9914 , \13998 );
nand \U$5680 ( \14499 , \14497 , \14498 );
or \U$5681 ( \14500 , \9921 , \14032 );
or \U$5682 ( \14501 , \11718 , \14065 );
nand \U$5683 ( \14502 , \14500 , \14501 );
nor \U$5684 ( \14503 , \14499 , \14502 );
nand \U$5685 ( \14504 , \14108 , \9859 );
not \U$5686 ( \14505 , \14038 );
or \U$5687 ( \14506 , \12183 , \14505 );
not \U$5688 ( \14507 , \12178 );
and \U$5689 ( \14508 , \14507 , \14112 );
and \U$5690 ( \14509 , \14058 , \9867 );
nor \U$5691 ( \14510 , \14508 , \14509 );
nand \U$5692 ( \14511 , \14504 , \14506 , \14510 );
or \U$5693 ( \14512 , \9887 , \14161 );
nand \U$5694 ( \14513 , \14025 , \9874 );
nand \U$5695 ( \14514 , \14045 , \9877 );
not \U$5696 ( \14515 , \14076 );
or \U$5697 ( \14516 , \9884 , \14515 );
and \U$5698 ( \14517 , \14512 , \14513 , \14514 , \14516 );
not \U$5699 ( \14518 , \14517 );
nor \U$5700 ( \14519 , \14511 , \14518 );
nand \U$5701 ( \14520 , \14496 , \14503 , \14519 );
xnor \U$5702 ( \14521 , \14520 , \9927 );
nor \U$5703 ( \14522 , \14488 , \14521 );
nand \U$5704 ( \14523 , \14417 , \14451 , \14522 );
not \U$5705 ( \14524 , \14523 );
nand \U$5706 ( \14525 , \9850 , \14033 );
nand \U$5707 ( \14526 , \9847 , \14272 );
not \U$5708 ( \14527 , \13998 );
and \U$5709 ( \14528 , \9842 , \14527 );
not \U$5710 ( \14529 , \14069 );
and \U$5711 ( \14530 , \9839 , \14529 );
nor \U$5712 ( \14531 , \14528 , \14530 );
nand \U$5713 ( \14532 , \14525 , \14526 , \14531 );
not \U$5714 ( \14533 , \14532 );
or \U$5715 ( \14534 , \9823 , \14104 );
or \U$5716 ( \14535 , \9827 , \14017 );
nand \U$5717 ( \14536 , \14534 , \14535 );
not \U$5718 ( \14537 , \9830 );
or \U$5719 ( \14538 , \14537 , \14012 );
or \U$5720 ( \14539 , \9834 , \14183 );
nand \U$5721 ( \14540 , \14538 , \14539 );
nor \U$5722 ( \14541 , \14536 , \14540 );
or \U$5723 ( \14542 , \9817 , \14161 );
nand \U$5724 ( \14543 , \14025 , \9805 );
nand \U$5725 ( \14544 , \14045 , \9808 );
not \U$5726 ( \14545 , \14091 );
or \U$5727 ( \14546 , \9814 , \14545 );
and \U$5728 ( \14547 , \14542 , \14543 , \14544 , \14546 );
not \U$5729 ( \14548 , \14547 );
not \U$5730 ( \14549 , \14548 );
not \U$5731 ( \14550 , \11494 );
and \U$5732 ( \14551 , \14550 , \14112 );
and \U$5733 ( \14552 , \14058 , \9797 );
nor \U$5734 ( \14553 , \14551 , \14552 );
not \U$5735 ( \14554 , \9791 );
and \U$5736 ( \14555 , \14554 , \14108 );
and \U$5737 ( \14556 , \14038 , \9794 );
nor \U$5738 ( \14557 , \14555 , \14556 );
and \U$5739 ( \14558 , \14549 , \14553 , \14557 );
nand \U$5740 ( \14559 , \14533 , \14541 , \14558 );
xnor \U$5741 ( \14560 , \14559 , \9857 );
nand \U$5742 ( \14561 , \14045 , \8915 );
nand \U$5743 ( \14562 , \14025 , \8860 );
nand \U$5744 ( \14563 , \14561 , \14562 );
not \U$5745 ( \14564 , \14563 );
not \U$5746 ( \14565 , \14076 );
or \U$5747 ( \14566 , \10775 , \14565 );
nand \U$5748 ( \14567 , \14080 , \8843 );
and \U$5749 ( \14568 , \14564 , \14566 , \14567 );
or \U$5750 ( \14569 , \13894 , \14012 );
or \U$5751 ( \14570 , \11540 , \14183 );
nand \U$5752 ( \14571 , \14569 , \14570 );
or \U$5753 ( \14572 , \11545 , \14017 );
not \U$5754 ( \14573 , \8953 );
or \U$5755 ( \14574 , \14573 , \14135 );
nand \U$5756 ( \14575 , \14572 , \14574 );
nor \U$5757 ( \14576 , \14571 , \14575 );
nand \U$5758 ( \14577 , \14108 , \8893 );
not \U$5759 ( \14578 , \14038 );
or \U$5760 ( \14579 , \8897 , \14578 );
not \U$5761 ( \14580 , \8882 );
and \U$5762 ( \14581 , \14580 , \14112 );
and \U$5763 ( \14582 , \14058 , \8868 );
nor \U$5764 ( \14583 , \14581 , \14582 );
nand \U$5765 ( \14584 , \14577 , \14579 , \14583 );
not \U$5766 ( \14585 , \14117 );
and \U$5767 ( \14586 , \8852 , \14585 );
not \U$5768 ( \14587 , \14121 );
and \U$5769 ( \14588 , \8904 , \14587 );
nor \U$5770 ( \14589 , \14586 , \14588 );
not \U$5771 ( \14590 , \11565 );
and \U$5772 ( \14591 , \14590 , \14033 );
not \U$5773 ( \14592 , \14063 );
and \U$5774 ( \14593 , \8827 , \14592 );
nor \U$5775 ( \14594 , \14591 , \14593 );
nand \U$5776 ( \14595 , \14589 , \14594 );
nor \U$5777 ( \14596 , \14584 , \14595 );
nand \U$5778 ( \14597 , \14568 , \14576 , \14596 );
xnor \U$5779 ( \14598 , \14597 , \8964 );
nor \U$5780 ( \14599 , \14560 , \14598 );
nand \U$5781 ( \14600 , \14045 , \9085 );
nand \U$5782 ( \14601 , \14025 , \9057 );
nand \U$5783 ( \14602 , \14600 , \14601 );
not \U$5784 ( \14603 , \14602 );
nand \U$5785 ( \14604 , \9102 , \14076 );
nand \U$5786 ( \14605 , \14080 , \9049 );
and \U$5787 ( \14606 , \14603 , \14604 , \14605 );
or \U$5788 ( \14607 , \11466 , \14012 );
or \U$5789 ( \14608 , \11468 , \13995 );
nand \U$5790 ( \14609 , \14607 , \14608 );
or \U$5791 ( \14610 , \11473 , \14138 );
or \U$5792 ( \14611 , \11471 , \14005 );
nand \U$5793 ( \14612 , \14610 , \14611 );
nor \U$5794 ( \14613 , \14609 , \14612 );
nand \U$5795 ( \14614 , \14108 , \9072 );
nand \U$5796 ( \14615 , \9075 , \14038 );
and \U$5797 ( \14616 , \14058 , \9063 );
and \U$5798 ( \14617 , \9067 , \14112 );
nor \U$5799 ( \14618 , \14616 , \14617 );
nand \U$5800 ( \14619 , \14614 , \14615 , \14618 );
not \U$5801 ( \14620 , \14197 );
and \U$5802 ( \14621 , \9054 , \14620 );
not \U$5803 ( \14622 , \14201 );
and \U$5804 ( \14623 , \9081 , \14622 );
nor \U$5805 ( \14624 , \14621 , \14623 );
and \U$5806 ( \14625 , \9098 , \14125 );
not \U$5807 ( \14626 , \14063 );
and \U$5808 ( \14627 , \9046 , \14626 );
nor \U$5809 ( \14628 , \14625 , \14627 );
nand \U$5810 ( \14629 , \14624 , \14628 );
nor \U$5811 ( \14630 , \14619 , \14629 );
nand \U$5812 ( \14631 , \14606 , \14613 , \14630 );
xnor \U$5813 ( \14632 , \14631 , \9119 );
nand \U$5814 ( \14633 , \14045 , \9157 );
nand \U$5815 ( \14634 , \14025 , \9132 );
nand \U$5816 ( \14635 , \14633 , \14634 );
not \U$5817 ( \14636 , \14635 );
nand \U$5818 ( \14637 , \9172 , \14076 );
nand \U$5819 ( \14638 , \14080 , \9124 );
and \U$5820 ( \14639 , \14636 , \14637 , \14638 );
or \U$5821 ( \14640 , \11424 , \14180 );
or \U$5822 ( \14641 , \11426 , \14097 );
nand \U$5823 ( \14642 , \14640 , \14641 );
or \U$5824 ( \14643 , \11431 , \14101 );
or \U$5825 ( \14644 , \11429 , \14104 );
nand \U$5826 ( \14645 , \14643 , \14644 );
nor \U$5827 ( \14646 , \14642 , \14645 );
nand \U$5828 ( \14647 , \14108 , \9147 );
nand \U$5829 ( \14648 , \9150 , \14038 );
and \U$5830 ( \14649 , \14058 , \9137 );
and \U$5831 ( \14650 , \9142 , \14112 );
nor \U$5832 ( \14651 , \14649 , \14650 );
nand \U$5833 ( \14652 , \14647 , \14648 , \14651 );
not \U$5834 ( \14653 , \14069 );
and \U$5835 ( \14654 , \9129 , \14653 );
not \U$5836 ( \14655 , \13998 );
and \U$5837 ( \14656 , \9155 , \14655 );
nor \U$5838 ( \14657 , \14654 , \14656 );
and \U$5839 ( \14658 , \9168 , \14125 );
not \U$5840 ( \14659 , \14063 );
and \U$5841 ( \14660 , \9121 , \14659 );
nor \U$5842 ( \14661 , \14658 , \14660 );
nand \U$5843 ( \14662 , \14657 , \14661 );
nor \U$5844 ( \14663 , \14652 , \14662 );
nand \U$5845 ( \14664 , \14639 , \14646 , \14663 );
xnor \U$5846 ( \14665 , \14664 , \9188 );
nor \U$5847 ( \14666 , \14632 , \14665 );
and \U$5848 ( \14667 , \14524 , \14599 , \14666 );
nand \U$5849 ( \14668 , \14086 , \14384 , \14667 );
not \U$5850 ( \14669 , \14668 );
not \U$5851 ( \14670 , \14669 );
or \U$5852 ( \14671 , \13989 , \14670 );
not \U$5853 ( \14672 , \14671 );
not \U$5854 ( \14673 , \14669 );
or \U$5855 ( \14674 , \13988 , \14673 );
not \U$5856 ( \14675 , \14674 );
or \U$5857 ( \14676 , \14672 , \14675 );
and \U$5858 ( \14677 , \13957 , \13960 , \14676 );
not \U$5859 ( \14678 , \14677 );
and \U$5860 ( \14679 , \13922 , \13943 , \13949 , \14678 );
not \U$5861 ( \14680 , \14679 );
not \U$5862 ( \14681 , \13245 );
and \U$5863 ( \14682 , \14681 , \13920 , \14668 );
not \U$5864 ( \14683 , \11757 );
buf \U$5865 ( \14684 , RIea91330_6888);
not \U$5866 ( \14685 , \12453 );
buf \U$5867 ( \14686 , \14685 );
buf \U$5868 ( \14687 , \12456 );
buf \U$5869 ( \14688 , \12458 );
buf \U$5870 ( \14689 , \10937 );
or \U$5871 ( \14690 , \14688 , \14689 );
and \U$5872 ( \14691 , \14687 , \14690 );
or \U$5873 ( \14692 , \14686 , \14691 );
and \U$5874 ( \14693 , \14684 , \14692 );
buf \U$5875 ( \14694 , \14693 );
not \U$5876 ( \14695 , \14694 );
not \U$5877 ( \14696 , \14689 );
buf \U$5878 ( \14697 , \14696 );
not \U$5879 ( \14698 , \14697 );
xnor \U$5880 ( \14699 , \14688 , \14689 );
buf \U$5881 ( \14700 , \14699 );
not \U$5882 ( \14701 , \14700 );
nand \U$5883 ( \14702 , \14698 , \14701 );
xor \U$5884 ( \14703 , \14687 , \14690 );
buf \U$5885 ( \14704 , \14703 );
not \U$5886 ( \14705 , \14704 );
xnor \U$5887 ( \14706 , \14686 , \14691 );
buf \U$5888 ( \14707 , \14706 );
not \U$5889 ( \14708 , \14707 );
nand \U$5890 ( \14709 , \14705 , \14708 );
or \U$5891 ( \14710 , \14702 , \14709 );
xor \U$5892 ( \14711 , \14684 , \14692 );
buf \U$5893 ( \14712 , \14711 );
nand \U$5894 ( \14713 , \14710 , \14712 );
and \U$5895 ( \14714 , \14695 , \14713 );
or \U$5896 ( \14715 , \9492 , \11966 );
or \U$5897 ( \14716 , \9494 , \11903 );
nand \U$5898 ( \14717 , \14715 , \14716 );
or \U$5899 ( \14718 , \9498 , \11959 );
or \U$5900 ( \14719 , \9500 , \11884 );
nand \U$5901 ( \14720 , \14718 , \14719 );
nor \U$5902 ( \14721 , \14717 , \14720 );
or \U$5903 ( \14722 , \9504 , \11817 );
or \U$5904 ( \14723 , \9506 , \11962 );
nand \U$5905 ( \14724 , \14722 , \14723 );
or \U$5906 ( \14725 , \9509 , \11950 );
or \U$5907 ( \14726 , \9511 , \11777 );
nand \U$5908 ( \14727 , \14725 , \14726 );
nor \U$5909 ( \14728 , \14724 , \14727 );
not \U$5910 ( \14729 , \9487 );
and \U$5911 ( \14730 , \14729 , \11826 );
and \U$5912 ( \14731 , \12122 , \10168 );
nor \U$5913 ( \14732 , \14730 , \14731 );
not \U$5914 ( \14733 , \9480 );
and \U$5915 ( \14734 , \14733 , \11864 );
and \U$5916 ( \14735 , \11814 , \12557 );
nor \U$5917 ( \14736 , \14734 , \14735 );
nand \U$5918 ( \14737 , \14732 , \14736 );
not \U$5919 ( \14738 , \14737 );
not \U$5920 ( \14739 , \9471 );
and \U$5921 ( \14740 , \14739 , \11892 );
and \U$5922 ( \14741 , \11869 , \9476 );
nor \U$5923 ( \14742 , \14740 , \14741 );
not \U$5924 ( \14743 , \9463 );
and \U$5925 ( \14744 , \14743 , \11936 );
and \U$5926 ( \14745 , \11934 , \9468 );
nor \U$5927 ( \14746 , \14744 , \14745 );
and \U$5928 ( \14747 , \14738 , \14742 , \14746 );
nand \U$5929 ( \14748 , \14721 , \14728 , \14747 );
not \U$5930 ( \14749 , \14748 );
and \U$5931 ( \14750 , \11846 , \9006 );
and \U$5932 ( \14751 , \8976 , \12122 );
nor \U$5933 ( \14752 , \14750 , \14751 );
and \U$5934 ( \14753 , \11832 , \9020 );
and \U$5935 ( \14754 , \8966 , \11826 );
nor \U$5936 ( \14755 , \14753 , \14754 );
or \U$5937 ( \14756 , \8991 , \11774 );
or \U$5938 ( \14757 , \11046 , \11791 );
nand \U$5939 ( \14758 , \14756 , \14757 );
or \U$5940 ( \14759 , \8997 , \11762 );
or \U$5941 ( \14760 , \9000 , \11777 );
nand \U$5942 ( \14761 , \14759 , \14760 );
nor \U$5943 ( \14762 , \14758 , \14761 );
nand \U$5944 ( \14763 , \14752 , \14755 , \14762 );
and \U$5945 ( \14764 , \11852 , \9030 );
and \U$5946 ( \14765 , \9034 , \11856 );
nor \U$5947 ( \14766 , \14764 , \14765 );
and \U$5948 ( \14767 , \12110 , \9014 );
and \U$5949 ( \14768 , \9011 , \11840 );
nor \U$5950 ( \14769 , \14767 , \14768 );
or \U$5951 ( \14770 , \8971 , \12193 );
or \U$5952 ( \14771 , \10370 , \11863 );
nand \U$5953 ( \14772 , \14770 , \14771 );
or \U$5954 ( \14773 , \11073 , \11767 );
or \U$5955 ( \14774 , \8980 , \11817 );
nand \U$5956 ( \14775 , \14773 , \14774 );
nor \U$5957 ( \14776 , \14772 , \14775 );
nand \U$5958 ( \14777 , \14766 , \14769 , \14776 );
nor \U$5959 ( \14778 , \14763 , \14777 );
xnor \U$5960 ( \14779 , \14778 , \9044 );
and \U$5961 ( \14780 , \11846 , \9225 );
and \U$5962 ( \14781 , \9204 , \12122 );
nor \U$5963 ( \14782 , \14780 , \14781 );
and \U$5964 ( \14783 , \11832 , \9239 );
and \U$5965 ( \14784 , \9196 , \11826 );
nor \U$5966 ( \14785 , \14783 , \14784 );
or \U$5967 ( \14786 , \11098 , \11774 );
or \U$5968 ( \14787 , \11101 , \11791 );
nand \U$5969 ( \14788 , \14786 , \14787 );
or \U$5970 ( \14789 , \9217 , \11762 );
or \U$5971 ( \14790 , \9220 , \11777 );
nand \U$5972 ( \14791 , \14789 , \14790 );
nor \U$5973 ( \14792 , \14788 , \14791 );
nand \U$5974 ( \14793 , \14782 , \14785 , \14792 );
and \U$5975 ( \14794 , \11852 , \9247 );
and \U$5976 ( \14795 , \9251 , \11856 );
nor \U$5977 ( \14796 , \14794 , \14795 );
and \U$5978 ( \14797 , \12110 , \9233 );
and \U$5979 ( \14798 , \9230 , \11840 );
nor \U$5980 ( \14799 , \14797 , \14798 );
or \U$5981 ( \14800 , \11088 , \11813 );
or \U$5982 ( \14801 , \10323 , \11863 );
nand \U$5983 ( \14802 , \14800 , \14801 );
or \U$5984 ( \14803 , \11125 , \11767 );
or \U$5985 ( \14804 , \11954 , \11817 );
nand \U$5986 ( \14805 , \14803 , \14804 );
nor \U$5987 ( \14806 , \14802 , \14805 );
nand \U$5988 ( \14807 , \14796 , \14799 , \14806 );
nor \U$5989 ( \14808 , \14793 , \14807 );
xnor \U$5990 ( \14809 , \14808 , \9260 );
or \U$5991 ( \14810 , \9266 , \12193 );
or \U$5992 ( \14811 , \10415 , \11863 );
nand \U$5993 ( \14812 , \14810 , \14811 );
or \U$5994 ( \14813 , \11298 , \11767 );
or \U$5995 ( \14814 , \9273 , \11817 );
nand \U$5996 ( \14815 , \14813 , \14814 );
nor \U$5997 ( \14816 , \14812 , \14815 );
or \U$5998 ( \14817 , \11286 , \11805 );
or \U$5999 ( \14818 , \11288 , \11839 );
nand \U$6000 ( \14819 , \14817 , \14818 );
or \U$6001 ( \14820 , \11293 , \11851 );
or \U$6002 ( \14821 , \11291 , \11855 );
nand \U$6003 ( \14822 , \14820 , \14821 );
nor \U$6004 ( \14823 , \14819 , \14822 );
and \U$6005 ( \14824 , \11846 , \9295 );
and \U$6006 ( \14825 , \9269 , \12122 );
nor \U$6007 ( \14826 , \14824 , \14825 );
and \U$6008 ( \14827 , \11832 , \9307 );
and \U$6009 ( \14828 , \9262 , \11826 );
nor \U$6010 ( \14829 , \14827 , \14828 );
nand \U$6011 ( \14830 , \14826 , \14829 );
not \U$6012 ( \14831 , \14830 );
and \U$6013 ( \14832 , \11898 , \9281 );
and \U$6014 ( \14833 , \9277 , \11896 );
nor \U$6015 ( \14834 , \14832 , \14833 );
not \U$6016 ( \14835 , \11762 );
and \U$6017 ( \14836 , \14835 , \9286 );
and \U$6018 ( \14837 , \9289 , \11979 );
nor \U$6019 ( \14838 , \14836 , \14837 );
and \U$6020 ( \14839 , \14831 , \14834 , \14838 );
nand \U$6021 ( \14840 , \14816 , \14823 , \14839 );
xnor \U$6022 ( \14841 , \14840 , \9327 );
not \U$6023 ( \14842 , \9397 );
not \U$6024 ( \14843 , \11812 );
or \U$6025 ( \14844 , \14842 , \14843 );
or \U$6026 ( \14845 , \10462 , \11863 );
nand \U$6027 ( \14846 , \14844 , \14845 );
or \U$6028 ( \14847 , \10464 , \11767 );
or \U$6029 ( \14848 , \9405 , \11817 );
nand \U$6030 ( \14849 , \14847 , \14848 );
nor \U$6031 ( \14850 , \14846 , \14849 );
or \U$6032 ( \14851 , \11243 , \11805 );
or \U$6033 ( \14852 , \11245 , \11882 );
nand \U$6034 ( \14853 , \14851 , \14852 );
or \U$6035 ( \14854 , \11250 , \11878 );
or \U$6036 ( \14855 , \11248 , \11874 );
nand \U$6037 ( \14856 , \14854 , \14855 );
nor \U$6038 ( \14857 , \14853 , \14856 );
and \U$6039 ( \14858 , \11846 , \9427 );
and \U$6040 ( \14859 , \9401 , \12122 );
nor \U$6041 ( \14860 , \14858 , \14859 );
and \U$6042 ( \14861 , \11832 , \9440 );
and \U$6043 ( \14862 , \9394 , \11826 );
nor \U$6044 ( \14863 , \14861 , \14862 );
nand \U$6045 ( \14864 , \14860 , \14863 );
not \U$6046 ( \14865 , \14864 );
and \U$6047 ( \14866 , \11934 , \9414 );
and \U$6048 ( \14867 , \9409 , \11936 );
nor \U$6049 ( \14868 , \14866 , \14867 );
and \U$6050 ( \14869 , \14835 , \9418 );
and \U$6051 ( \14870 , \9421 , \11979 );
nor \U$6052 ( \14871 , \14869 , \14870 );
and \U$6053 ( \14872 , \14865 , \14868 , \14871 );
nand \U$6054 ( \14873 , \14850 , \14857 , \14872 );
xnor \U$6055 ( \14874 , \14873 , \9460 );
nor \U$6056 ( \14875 , \14841 , \14874 );
nand \U$6057 ( \14876 , \14779 , \14809 , \14875 );
not \U$6058 ( \14877 , \14876 );
or \U$6059 ( \14878 , \8844 , \11813 );
or \U$6060 ( \14879 , \10775 , \11863 );
nand \U$6061 ( \14880 , \14878 , \14879 );
or \U$6062 ( \14881 , \11533 , \11767 );
or \U$6063 ( \14882 , \8861 , \11817 );
nand \U$6064 ( \14883 , \14881 , \14882 );
nor \U$6065 ( \14884 , \14880 , \14883 );
or \U$6066 ( \14885 , \13894 , \11805 );
or \U$6067 ( \14886 , \11540 , \11966 );
nand \U$6068 ( \14887 , \14885 , \14886 );
or \U$6069 ( \14888 , \11545 , \11962 );
or \U$6070 ( \14889 , \14573 , \11959 );
nand \U$6071 ( \14890 , \14888 , \14889 );
nor \U$6072 ( \14891 , \14887 , \14890 );
not \U$6073 ( \14892 , \11843 );
and \U$6074 ( \14893 , \14892 , \8904 );
and \U$6075 ( \14894 , \8852 , \12122 );
nor \U$6076 ( \14895 , \14893 , \14894 );
and \U$6077 ( \14896 , \11832 , \8934 );
and \U$6078 ( \14897 , \8827 , \11826 );
nor \U$6079 ( \14898 , \14896 , \14897 );
nand \U$6080 ( \14899 , \14895 , \14898 );
not \U$6081 ( \14900 , \14899 );
not \U$6082 ( \14901 , \12351 );
and \U$6083 ( \14902 , \14901 , \11936 );
and \U$6084 ( \14903 , \11934 , \8881 );
nor \U$6085 ( \14904 , \14902 , \14903 );
not \U$6086 ( \14905 , \8897 );
and \U$6087 ( \14906 , \14905 , \11979 );
and \U$6088 ( \14907 , \14835 , \8893 );
nor \U$6089 ( \14908 , \14906 , \14907 );
and \U$6090 ( \14909 , \14900 , \14904 , \14908 );
nand \U$6091 ( \14910 , \14884 , \14891 , \14909 );
xnor \U$6092 ( \14911 , \14910 , \8964 );
or \U$6093 ( \14912 , \9050 , \11813 );
or \U$6094 ( \14913 , \10859 , \11863 );
nand \U$6095 ( \14914 , \14912 , \14913 );
or \U$6096 ( \14915 , \9086 , \11767 );
or \U$6097 ( \14916 , \9058 , \11817 );
nand \U$6098 ( \14917 , \14915 , \14916 );
nor \U$6099 ( \14918 , \14914 , \14917 );
or \U$6100 ( \14919 , \11466 , \11805 );
or \U$6101 ( \14920 , \11468 , \11839 );
nand \U$6102 ( \14921 , \14919 , \14920 );
or \U$6103 ( \14922 , \11473 , \11851 );
or \U$6104 ( \14923 , \11471 , \11855 );
nand \U$6105 ( \14924 , \14922 , \14923 );
nor \U$6106 ( \14925 , \14921 , \14924 );
and \U$6107 ( \14926 , \11846 , \9081 );
and \U$6108 ( \14927 , \9054 , \12122 );
nor \U$6109 ( \14928 , \14926 , \14927 );
and \U$6110 ( \14929 , \11832 , \9098 );
and \U$6111 ( \14930 , \9046 , \11826 );
nor \U$6112 ( \14931 , \14929 , \14930 );
nand \U$6113 ( \14932 , \14928 , \14931 );
not \U$6114 ( \14933 , \14932 );
not \U$6115 ( \14934 , \11458 );
and \U$6116 ( \14935 , \14934 , \11896 );
and \U$6117 ( \14936 , \11898 , \9067 );
nor \U$6118 ( \14937 , \14935 , \14936 );
not \U$6119 ( \14938 , \9076 );
and \U$6120 ( \14939 , \14938 , \11979 );
and \U$6121 ( \14940 , \14835 , \9072 );
nor \U$6122 ( \14941 , \14939 , \14940 );
and \U$6123 ( \14942 , \14933 , \14937 , \14941 );
nand \U$6124 ( \14943 , \14918 , \14925 , \14942 );
xnor \U$6125 ( \14944 , \14943 , \9119 );
nor \U$6126 ( \14945 , \14911 , \14944 );
or \U$6127 ( \14946 , \9335 , \11813 );
or \U$6128 ( \14947 , \10553 , \11863 );
nand \U$6129 ( \14948 , \14946 , \14947 );
or \U$6130 ( \14949 , \11357 , \11767 );
or \U$6131 ( \14950 , \9342 , \11817 );
nand \U$6132 ( \14951 , \14949 , \14950 );
nor \U$6133 ( \14952 , \14948 , \14951 );
or \U$6134 ( \14953 , \13593 , \11805 );
or \U$6135 ( \14954 , \11365 , \11882 );
nand \U$6136 ( \14955 , \14953 , \14954 );
or \U$6137 ( \14956 , \12874 , \11878 );
or \U$6138 ( \14957 , \11371 , \11874 );
nand \U$6139 ( \14958 , \14956 , \14957 );
nor \U$6140 ( \14959 , \14955 , \14958 );
not \U$6141 ( \14960 , \9339 );
and \U$6142 ( \14961 , \14960 , \12122 );
and \U$6143 ( \14962 , \11846 , \9361 );
nor \U$6144 ( \14963 , \14961 , \14962 );
not \U$6145 ( \14964 , \9332 );
and \U$6146 ( \14965 , \14964 , \11826 );
and \U$6147 ( \14966 , \11832 , \9374 );
nor \U$6148 ( \14967 , \14965 , \14966 );
nand \U$6149 ( \14968 , \14963 , \14967 );
not \U$6150 ( \14969 , \14968 );
not \U$6151 ( \14970 , \12141 );
and \U$6152 ( \14971 , \14970 , \11936 );
and \U$6153 ( \14972 , \11934 , \9348 );
nor \U$6154 ( \14973 , \14971 , \14972 );
not \U$6155 ( \14974 , \9357 );
and \U$6156 ( \14975 , \14974 , \11979 );
and \U$6157 ( \14976 , \14835 , \9353 );
nor \U$6158 ( \14977 , \14975 , \14976 );
and \U$6159 ( \14978 , \14969 , \14973 , \14977 );
nand \U$6160 ( \14979 , \14952 , \14959 , \14978 );
xnor \U$6161 ( \14980 , \14979 , \9392 );
or \U$6162 ( \14981 , \9125 , \12193 );
or \U$6163 ( \14982 , \10901 , \11863 );
nand \U$6164 ( \14983 , \14981 , \14982 );
or \U$6165 ( \14984 , \11436 , \11767 );
or \U$6166 ( \14985 , \9133 , \11817 );
nand \U$6167 ( \14986 , \14984 , \14985 );
nor \U$6168 ( \14987 , \14983 , \14986 );
or \U$6169 ( \14988 , \11424 , \11884 );
or \U$6170 ( \14989 , \11426 , \11966 );
nand \U$6171 ( \14990 , \14988 , \14989 );
or \U$6172 ( \14991 , \11431 , \11962 );
or \U$6173 ( \14992 , \11429 , \11959 );
nand \U$6174 ( \14993 , \14991 , \14992 );
nor \U$6175 ( \14994 , \14990 , \14993 );
not \U$6176 ( \14995 , \9130 );
and \U$6177 ( \14996 , \14995 , \12122 );
and \U$6178 ( \14997 , \11846 , \9155 );
nor \U$6179 ( \14998 , \14996 , \14997 );
not \U$6180 ( \14999 , \9122 );
and \U$6181 ( \15000 , \14999 , \11826 );
and \U$6182 ( \15001 , \11832 , \9168 );
nor \U$6183 ( \15002 , \15000 , \15001 );
nand \U$6184 ( \15003 , \14998 , \15002 );
not \U$6185 ( \15004 , \15003 );
not \U$6186 ( \15005 , \11416 );
and \U$6187 ( \15006 , \15005 , \11896 );
and \U$6188 ( \15007 , \11898 , \9142 );
nor \U$6189 ( \15008 , \15006 , \15007 );
not \U$6190 ( \15009 , \9151 );
and \U$6191 ( \15010 , \15009 , \11979 );
and \U$6192 ( \15011 , \14835 , \9147 );
nor \U$6193 ( \15012 , \15010 , \15011 );
and \U$6194 ( \15013 , \15004 , \15008 , \15012 );
nand \U$6195 ( \15014 , \14987 , \14994 , \15013 );
xnor \U$6196 ( \15015 , \15014 , \9188 );
nor \U$6197 ( \15016 , \14980 , \15015 );
and \U$6198 ( \15017 , \14877 , \14945 , \15016 );
and \U$6199 ( \15018 , \11814 , \9545 );
and \U$6200 ( \15019 , \9542 , \11864 );
nor \U$6201 ( \15020 , \15018 , \15019 );
and \U$6202 ( \15021 , \11818 , \9533 );
and \U$6203 ( \15022 , \9536 , \11869 );
nor \U$6204 ( \15023 , \15021 , \15022 );
or \U$6205 ( \15024 , \13658 , \11774 );
or \U$6206 ( \15025 , \9527 , \11791 );
nand \U$6207 ( \15026 , \15024 , \15025 );
or \U$6208 ( \15027 , \9519 , \11762 );
or \U$6209 ( \15028 , \14434 , \11777 );
nand \U$6210 ( \15029 , \15027 , \15028 );
nor \U$6211 ( \15030 , \15026 , \15029 );
nand \U$6212 ( \15031 , \15020 , \15023 , \15030 );
and \U$6213 ( \15032 , \11832 , \9578 );
and \U$6214 ( \15033 , \9575 , \11826 );
nor \U$6215 ( \15034 , \15032 , \15033 );
and \U$6216 ( \15035 , \12122 , \9568 );
and \U$6217 ( \15036 , \9571 , \11846 );
nor \U$6218 ( \15037 , \15035 , \15036 );
or \U$6219 ( \15038 , \9552 , \11855 );
or \U$6220 ( \15039 , \9557 , \11851 );
nand \U$6221 ( \15040 , \15038 , \15039 );
or \U$6222 ( \15041 , \9564 , \11839 );
or \U$6223 ( \15042 , \11582 , \11884 );
nand \U$6224 ( \15043 , \15041 , \15042 );
nor \U$6225 ( \15044 , \15040 , \15043 );
nand \U$6226 ( \15045 , \15034 , \15037 , \15044 );
nor \U$6227 ( \15046 , \15031 , \15045 );
xnor \U$6228 ( \15047 , \15046 , \9585 );
and \U$6229 ( \15048 , \11892 , \9744 );
and \U$6230 ( \15049 , \9747 , \11979 );
nor \U$6231 ( \15050 , \15048 , \15049 );
and \U$6232 ( \15051 , \11898 , \9739 );
and \U$6233 ( \15052 , \9736 , \11896 );
nor \U$6234 ( \15053 , \15051 , \15052 );
or \U$6235 ( \15054 , \9722 , \11901 );
or \U$6236 ( \15055 , \9725 , \11845 );
nand \U$6237 ( \15056 , \15054 , \15055 );
or \U$6238 ( \15057 , \9732 , \11950 );
or \U$6239 ( \15058 , \13305 , \11907 );
nand \U$6240 ( \15059 , \15057 , \15058 );
nor \U$6241 ( \15060 , \15056 , \15059 );
nand \U$6242 ( \15061 , \15050 , \15053 , \15060 );
and \U$6243 ( \15062 , \11814 , \9776 );
and \U$6244 ( \15063 , \9779 , \11864 );
nor \U$6245 ( \15064 , \15062 , \15063 );
and \U$6246 ( \15065 , \11818 , \9772 );
and \U$6247 ( \15066 , \9769 , \11869 );
nor \U$6248 ( \15067 , \15065 , \15066 );
or \U$6249 ( \15068 , \10194 , \11959 );
or \U$6250 ( \15069 , \10197 , \11962 );
nand \U$6251 ( \15070 , \15068 , \15069 );
or \U$6252 ( \15071 , \11193 , \11966 );
or \U$6253 ( \15072 , \11195 , \11884 );
nand \U$6254 ( \15073 , \15071 , \15072 );
nor \U$6255 ( \15074 , \15070 , \15073 );
nand \U$6256 ( \15075 , \15064 , \15067 , \15074 );
nor \U$6257 ( \15076 , \15061 , \15075 );
xnor \U$6258 ( \15077 , \15076 , \9786 );
or \U$6259 ( \15078 , \9620 , \11855 );
or \U$6260 ( \15079 , \9625 , \11851 );
nand \U$6261 ( \15080 , \15078 , \15079 );
or \U$6262 ( \15081 , \9632 , \11839 );
or \U$6263 ( \15082 , \11314 , \11805 );
nand \U$6264 ( \15083 , \15081 , \15082 );
nor \U$6265 ( \15084 , \15080 , \15083 );
not \U$6266 ( \15085 , \9639 );
not \U$6267 ( \15086 , \11844 );
or \U$6268 ( \15087 , \15085 , \15086 );
or \U$6269 ( \15088 , \9637 , \11901 );
nand \U$6270 ( \15089 , \15087 , \15088 );
or \U$6271 ( \15090 , \9647 , \11831 );
or \U$6272 ( \15091 , \11322 , \11907 );
nand \U$6273 ( \15092 , \15090 , \15091 );
nor \U$6274 ( \15093 , \15089 , \15092 );
and \U$6275 ( \15094 , \14835 , \9587 );
and \U$6276 ( \15095 , \9592 , \11979 );
nor \U$6277 ( \15096 , \15094 , \15095 );
not \U$6278 ( \15097 , \11774 );
and \U$6279 ( \15098 , \15097 , \9600 );
not \U$6280 ( \15099 , \11791 );
and \U$6281 ( \15100 , \9596 , \15099 );
nor \U$6282 ( \15101 , \15098 , \15100 );
nand \U$6283 ( \15102 , \15096 , \15101 );
not \U$6284 ( \15103 , \15102 );
and \U$6285 ( \15104 , \11818 , \9603 );
and \U$6286 ( \15105 , \9606 , \11869 );
nor \U$6287 ( \15106 , \15104 , \15105 );
and \U$6288 ( \15107 , \11814 , \9613 );
and \U$6289 ( \15108 , \9610 , \11864 );
nor \U$6290 ( \15109 , \15107 , \15108 );
and \U$6291 ( \15110 , \15103 , \15106 , \15109 );
nand \U$6292 ( \15111 , \15084 , \15093 , \15110 );
xnor \U$6293 ( \15112 , \15111 , \9653 );
or \U$6294 ( \15113 , \11138 , \11817 );
or \U$6295 ( \15114 , \11140 , \11767 );
nand \U$6296 ( \15115 , \15113 , \15114 );
or \U$6297 ( \15116 , \10244 , \11800 );
or \U$6298 ( \15117 , \11145 , \12193 );
nand \U$6299 ( \15118 , \15116 , \15117 );
nor \U$6300 ( \15119 , \15115 , \15118 );
or \U$6301 ( \15120 , \10248 , \11874 );
or \U$6302 ( \15121 , \10250 , \11878 );
nand \U$6303 ( \15122 , \15120 , \15121 );
or \U$6304 ( \15123 , \11152 , \11882 );
or \U$6305 ( \15124 , \11154 , \11884 );
nand \U$6306 ( \15125 , \15123 , \15124 );
nor \U$6307 ( \15126 , \15122 , \15125 );
not \U$6308 ( \15127 , \9683 );
and \U$6309 ( \15128 , \15127 , \11890 );
and \U$6310 ( \15129 , \14835 , \9679 );
nor \U$6311 ( \15130 , \15128 , \15129 );
not \U$6312 ( \15131 , \11923 );
and \U$6313 ( \15132 , \15131 , \11936 );
and \U$6314 ( \15133 , \15097 , \9675 );
nor \U$6315 ( \15134 , \15132 , \15133 );
nand \U$6316 ( \15135 , \15130 , \15134 );
not \U$6317 ( \15136 , \15135 );
and \U$6318 ( \15137 , \12122 , \9656 );
and \U$6319 ( \15138 , \9660 , \11846 );
nor \U$6320 ( \15139 , \15137 , \15138 );
and \U$6321 ( \15140 , \11832 , \9667 );
and \U$6322 ( \15141 , \9664 , \11826 );
nor \U$6323 ( \15142 , \15140 , \15141 );
and \U$6324 ( \15143 , \15136 , \15139 , \15142 );
nand \U$6325 ( \15144 , \15119 , \15126 , \15143 );
xnor \U$6326 ( \15145 , \15144 , \9719 );
nor \U$6327 ( \15146 , \15112 , \15145 );
nand \U$6328 ( \15147 , \15047 , \15077 , \15146 );
not \U$6329 ( \15148 , \15147 );
or \U$6330 ( \15149 , \11618 , \11874 );
or \U$6331 ( \15150 , \11620 , \11878 );
nand \U$6332 ( \15151 , \15149 , \15150 );
or \U$6333 ( \15152 , \11623 , \11882 );
or \U$6334 ( \15153 , \11625 , \11884 );
nand \U$6335 ( \15154 , \15152 , \15153 );
nor \U$6336 ( \15155 , \15151 , \15154 );
or \U$6337 ( \15156 , \11635 , \11788 );
or \U$6338 ( \15157 , \11629 , \11845 );
nand \U$6339 ( \15158 , \15156 , \15157 );
not \U$6340 ( \15159 , \9984 );
not \U$6341 ( \15160 , \11830 );
or \U$6342 ( \15161 , \15159 , \15160 );
or \U$6343 ( \15162 , \11633 , \11907 );
nand \U$6344 ( \15163 , \15161 , \15162 );
nor \U$6345 ( \15164 , \15158 , \15163 );
and \U$6346 ( \15165 , \14835 , \9951 );
and \U$6347 ( \15166 , \9954 , \11979 );
nor \U$6348 ( \15167 , \15165 , \15166 );
and \U$6349 ( \15168 , \15097 , \9947 );
and \U$6350 ( \15169 , \9944 , \11896 );
nor \U$6351 ( \15170 , \15168 , \15169 );
nand \U$6352 ( \15171 , \15167 , \15170 );
not \U$6353 ( \15172 , \15171 );
and \U$6354 ( \15173 , \11818 , \9929 );
and \U$6355 ( \15174 , \9932 , \11869 );
nor \U$6356 ( \15175 , \15173 , \15174 );
and \U$6357 ( \15176 , \11814 , \9939 );
and \U$6358 ( \15177 , \9936 , \11864 );
nor \U$6359 ( \15178 , \15176 , \15177 );
and \U$6360 ( \15179 , \15172 , \15175 , \15178 );
nand \U$6361 ( \15180 , \15155 , \15164 , \15179 );
xnor \U$6362 ( \15181 , \15180 , \9990 );
or \U$6363 ( \15182 , \12230 , \11959 );
or \U$6364 ( \15183 , \11698 , \11962 );
nand \U$6365 ( \15184 , \15182 , \15183 );
or \U$6366 ( \15185 , \11693 , \11966 );
or \U$6367 ( \15186 , \12235 , \11884 );
nand \U$6368 ( \15187 , \15185 , \15186 );
nor \U$6369 ( \15188 , \15184 , \15187 );
or \U$6370 ( \15189 , \11684 , \11788 );
or \U$6371 ( \15190 , \12222 , \11845 );
nand \U$6372 ( \15191 , \15189 , \15190 );
or \U$6373 ( \15192 , \11674 , \11950 );
or \U$6374 ( \15193 , \11681 , \11907 );
nand \U$6375 ( \15194 , \15192 , \15193 );
nor \U$6376 ( \15195 , \15191 , \15194 );
and \U$6377 ( \15196 , \11814 , \10020 );
and \U$6378 ( \15197 , \10017 , \11864 );
nor \U$6379 ( \15198 , \15196 , \15197 );
and \U$6380 ( \15199 , \11818 , \10009 );
and \U$6381 ( \15200 , \10012 , \11869 );
nor \U$6382 ( \15201 , \15199 , \15200 );
nand \U$6383 ( \15202 , \15198 , \15201 );
not \U$6384 ( \15203 , \15202 );
and \U$6385 ( \15204 , \11898 , \9996 );
and \U$6386 ( \15205 , \9992 , \11936 );
nor \U$6387 ( \15206 , \15204 , \15205 );
and \U$6388 ( \15207 , \14835 , \10001 );
and \U$6389 ( \15208 , \10004 , \11890 );
nor \U$6390 ( \15209 , \15207 , \15208 );
and \U$6391 ( \15210 , \15203 , \15206 , \15209 );
nand \U$6392 ( \15211 , \15188 , \15195 , \15210 );
xnor \U$6393 ( \15212 , \15211 , \10055 );
nor \U$6394 ( \15213 , \15181 , \15212 );
or \U$6395 ( \15214 , \9895 , \11855 );
or \U$6396 ( \15215 , \9898 , \11851 );
nand \U$6397 ( \15216 , \15214 , \15215 );
or \U$6398 ( \15217 , \9906 , \11839 );
or \U$6399 ( \15218 , \11711 , \11884 );
nand \U$6400 ( \15219 , \15217 , \15218 );
nor \U$6401 ( \15220 , \15216 , \15219 );
or \U$6402 ( \15221 , \9911 , \11788 );
or \U$6403 ( \15222 , \9914 , \11903 );
nand \U$6404 ( \15223 , \15221 , \15222 );
or \U$6405 ( \15224 , \9921 , \11950 );
or \U$6406 ( \15225 , \11718 , \11907 );
nand \U$6407 ( \15226 , \15224 , \15225 );
nor \U$6408 ( \15227 , \15223 , \15226 );
and \U$6409 ( \15228 , \14835 , \9859 );
and \U$6410 ( \15229 , \9863 , \11979 );
nor \U$6411 ( \15230 , \15228 , \15229 );
and \U$6412 ( \15231 , \15097 , \9871 );
and \U$6413 ( \15232 , \9867 , \15099 );
nor \U$6414 ( \15233 , \15231 , \15232 );
nand \U$6415 ( \15234 , \15230 , \15233 );
not \U$6416 ( \15235 , \15234 );
and \U$6417 ( \15236 , \11818 , \9874 );
and \U$6418 ( \15237 , \9877 , \11869 );
nor \U$6419 ( \15238 , \15236 , \15237 );
not \U$6420 ( \15239 , \9884 );
not \U$6421 ( \15240 , \11798 );
and \U$6422 ( \15241 , \15239 , \15240 );
and \U$6423 ( \15242 , \11814 , \9886 );
or \U$6424 ( \15243 , \15241 , \15242 );
not \U$6425 ( \15244 , \15243 );
and \U$6426 ( \15245 , \15235 , \15238 , \15244 );
nand \U$6427 ( \15246 , \15220 , \15227 , \15245 );
xnor \U$6428 ( \15247 , \15246 , \9927 );
or \U$6429 ( \15248 , \9823 , \11874 );
or \U$6430 ( \15249 , \9827 , \11878 );
nand \U$6431 ( \15250 , \15248 , \15249 );
or \U$6432 ( \15251 , \9834 , \11882 );
or \U$6433 ( \15252 , \12311 , \11884 );
nand \U$6434 ( \15253 , \15251 , \15252 );
nor \U$6435 ( \15254 , \15250 , \15253 );
or \U$6436 ( \15255 , \9840 , \11788 );
or \U$6437 ( \15256 , \9843 , \11903 );
nand \U$6438 ( \15257 , \15255 , \15256 );
or \U$6439 ( \15258 , \9851 , \11950 );
or \U$6440 ( \15259 , \11505 , \11907 );
nand \U$6441 ( \15260 , \15258 , \15259 );
nor \U$6442 ( \15261 , \15257 , \15260 );
and \U$6443 ( \15262 , \11814 , \9816 );
and \U$6444 ( \15263 , \9813 , \11864 );
nor \U$6445 ( \15264 , \15262 , \15263 );
and \U$6446 ( \15265 , \11818 , \9805 );
and \U$6447 ( \15266 , \9808 , \11869 );
nor \U$6448 ( \15267 , \15265 , \15266 );
nand \U$6449 ( \15268 , \15264 , \15267 );
not \U$6450 ( \15269 , \15268 );
and \U$6451 ( \15270 , \11934 , \9801 );
and \U$6452 ( \15271 , \9797 , \11936 );
nor \U$6453 ( \15272 , \15270 , \15271 );
and \U$6454 ( \15273 , \14835 , \9790 );
and \U$6455 ( \15274 , \9794 , \11979 );
nor \U$6456 ( \15275 , \15273 , \15274 );
and \U$6457 ( \15276 , \15269 , \15272 , \15275 );
nand \U$6458 ( \15277 , \15254 , \15261 , \15276 );
xnor \U$6459 ( \15278 , \15277 , \9857 );
nor \U$6460 ( \15279 , \15247 , \15278 );
and \U$6461 ( \15280 , \15148 , \15213 , \15279 );
nand \U$6462 ( \15281 , \14749 , \15017 , \15280 );
not \U$6463 ( \15282 , \15281 );
not \U$6464 ( \15283 , \15282 );
or \U$6465 ( \15284 , \14714 , \15283 );
not \U$6466 ( \15285 , \15284 );
nand \U$6467 ( \15286 , \14714 , \15282 );
not \U$6468 ( \15287 , \15286 );
or \U$6469 ( \15288 , \15285 , \15287 );
not \U$6470 ( \15289 , \15288 );
not \U$6471 ( \15290 , \15289 );
and \U$6472 ( \15291 , \14683 , \15290 );
not \U$6473 ( \15292 , \10066 );
buf \U$6474 ( \15293 , RIea91330_6888);
buf \U$6475 ( \15294 , \14685 );
buf \U$6476 ( \15295 , \12456 );
not \U$6477 ( \15296 , \15295 );
not \U$6478 ( \15297 , \15296 );
or \U$6479 ( \15298 , \15294 , \15297 );
and \U$6480 ( \15299 , \15293 , \15298 );
buf \U$6481 ( \15300 , \15299 );
not \U$6482 ( \15301 , \15300 );
buf \U$6483 ( \15302 , \10919 );
not \U$6484 ( \15303 , \15302 );
buf \U$6485 ( \15304 , \12458 );
not \U$6486 ( \15305 , \15304 );
nand \U$6487 ( \15306 , \15303 , \15305 );
buf \U$6488 ( \15307 , \15296 );
not \U$6489 ( \15308 , \15307 );
xnor \U$6490 ( \15309 , \15294 , \15297 );
buf \U$6491 ( \15310 , \15309 );
not \U$6492 ( \15311 , \15310 );
nand \U$6493 ( \15312 , \15308 , \15311 );
or \U$6494 ( \15313 , \15306 , \15312 );
xor \U$6495 ( \15314 , \15293 , \15298 );
buf \U$6496 ( \15315 , \15314 );
nand \U$6497 ( \15316 , \15313 , \15315 );
and \U$6498 ( \15317 , \15301 , \15316 );
not \U$6499 ( \15318 , \10138 );
or \U$6500 ( \15319 , \9506 , \15318 );
not \U$6501 ( \15320 , \10417 );
and \U$6502 ( \15321 , \13270 , \15320 );
not \U$6503 ( \15322 , \10228 );
and \U$6504 ( \15323 , \10976 , \15322 );
nor \U$6505 ( \15324 , \15321 , \15323 );
not \U$6506 ( \15325 , \10100 );
or \U$6507 ( \15326 , \9511 , \15325 );
nand \U$6508 ( \15327 , \15319 , \15324 , \15326 );
not \U$6509 ( \15328 , \15327 );
and \U$6510 ( \15329 , \10143 , \10062 );
not \U$6511 ( \15330 , \10358 );
and \U$6512 ( \15331 , \12513 , \15330 );
nor \U$6513 ( \15332 , \15329 , \15331 );
and \U$6514 ( \15333 , \10133 , \10085 );
not \U$6515 ( \15334 , \10118 );
and \U$6516 ( \15335 , \13262 , \15334 );
nor \U$6517 ( \15336 , \15333 , \15335 );
and \U$6518 ( \15337 , \15328 , \15332 , \15336 );
not \U$6519 ( \15338 , \10080 );
and \U$6520 ( \15339 , \9472 , \15338 );
not \U$6521 ( \15340 , \15339 );
not \U$6522 ( \15341 , \10275 );
and \U$6523 ( \15342 , \9476 , \15341 );
not \U$6524 ( \15343 , \15342 );
not \U$6525 ( \15344 , \10114 );
and \U$6526 ( \15345 , \10986 , \15344 );
not \U$6527 ( \15346 , \10093 );
and \U$6528 ( \15347 , \9468 , \15346 );
nor \U$6529 ( \15348 , \15345 , \15347 );
nand \U$6530 ( \15349 , \15340 , \15343 , \15348 );
or \U$6531 ( \15350 , \9482 , \10220 );
not \U$6532 ( \15351 , \10236 );
or \U$6533 ( \15352 , \9485 , \15351 );
not \U$6534 ( \15353 , \10160 );
or \U$6535 ( \15354 , \9487 , \15353 );
not \U$6536 ( \15355 , \10127 );
or \U$6537 ( \15356 , \9480 , \15355 );
and \U$6538 ( \15357 , \15350 , \15352 , \15354 , \15356 );
not \U$6539 ( \15358 , \15357 );
nor \U$6540 ( \15359 , \15349 , \15358 );
nand \U$6541 ( \15360 , \15337 , \15359 );
not \U$6542 ( \15361 , \15360 );
or \U$6543 ( \15362 , \8967 , \10621 );
or \U$6544 ( \15363 , \11036 , \10417 );
nand \U$6545 ( \15364 , \15362 , \15363 );
not \U$6546 ( \15365 , \15364 );
nand \U$6547 ( \15366 , \8976 , \10236 );
nand \U$6548 ( \15367 , \9006 , \10143 );
and \U$6549 ( \15368 , \15365 , \15366 , \15367 );
or \U$6550 ( \15369 , \8991 , \10842 );
or \U$6551 ( \15370 , \11046 , \10114 );
nand \U$6552 ( \15371 , \15369 , \15370 );
not \U$6553 ( \15372 , \15371 );
nand \U$6554 ( \15373 , \8999 , \10100 );
not \U$6555 ( \15374 , \10080 );
nand \U$6556 ( \15375 , \8996 , \15374 );
and \U$6557 ( \15376 , \15372 , \15373 , \15375 );
not \U$6558 ( \15377 , \10145 );
and \U$6559 ( \15378 , \9011 , \15377 );
not \U$6560 ( \15379 , \15378 );
not \U$6561 ( \15380 , \10260 );
and \U$6562 ( \15381 , \9014 , \15380 );
not \U$6563 ( \15382 , \15381 );
and \U$6564 ( \15383 , \10318 , \9030 );
and \U$6565 ( \15384 , \9034 , \10212 );
nor \U$6566 ( \15385 , \15383 , \15384 );
and \U$6567 ( \15386 , \15379 , \15382 , \15385 );
not \U$6568 ( \15387 , \15386 );
not \U$6569 ( \15388 , \10220 );
and \U$6570 ( \15389 , \8970 , \15388 );
not \U$6571 ( \15390 , \15389 );
nand \U$6572 ( \15391 , \9025 , \10127 );
not \U$6573 ( \15392 , \10170 );
and \U$6574 ( \15393 , \8979 , \15392 );
not \U$6575 ( \15394 , \10224 );
and \U$6576 ( \15395 , \9009 , \15394 );
nor \U$6577 ( \15396 , \15393 , \15395 );
nand \U$6578 ( \15397 , \15390 , \15391 , \15396 );
nor \U$6579 ( \15398 , \15387 , \15397 );
nand \U$6580 ( \15399 , \15368 , \15376 , \15398 );
xnor \U$6581 ( \15400 , RIb7b94a0_249, \15399 );
or \U$6582 ( \15401 , \9197 , \10159 );
or \U$6583 ( \15402 , \11093 , \10190 );
nand \U$6584 ( \15403 , \15401 , \15402 );
not \U$6585 ( \15404 , \15403 );
nand \U$6586 ( \15405 , \9204 , \10236 );
nand \U$6587 ( \15406 , \9225 , \10143 );
and \U$6588 ( \15407 , \15404 , \15405 , \15406 );
or \U$6589 ( \15408 , \11098 , \10842 );
or \U$6590 ( \15409 , \11101 , \10114 );
nand \U$6591 ( \15410 , \15408 , \15409 );
not \U$6592 ( \15411 , \15410 );
nand \U$6593 ( \15412 , \9219 , \10100 );
nand \U$6594 ( \15413 , \9216 , \15374 );
and \U$6595 ( \15414 , \15411 , \15412 , \15413 );
not \U$6596 ( \15415 , \10145 );
and \U$6597 ( \15416 , \9230 , \15415 );
not \U$6598 ( \15417 , \15416 );
not \U$6599 ( \15418 , \10118 );
and \U$6600 ( \15419 , \9233 , \15418 );
not \U$6601 ( \15420 , \15419 );
and \U$6602 ( \15421 , \10318 , \9247 );
and \U$6603 ( \15422 , \9251 , \10212 );
nor \U$6604 ( \15423 , \15421 , \15422 );
and \U$6605 ( \15424 , \15417 , \15420 , \15423 );
not \U$6606 ( \15425 , \15424 );
not \U$6607 ( \15426 , \10271 );
and \U$6608 ( \15427 , \9193 , \15426 );
not \U$6609 ( \15428 , \15427 );
nand \U$6610 ( \15429 , \9242 , \10127 );
not \U$6611 ( \15430 , \10228 );
and \U$6612 ( \15431 , \9200 , \15430 );
not \U$6613 ( \15432 , \10340 );
and \U$6614 ( \15433 , \9228 , \15432 );
nor \U$6615 ( \15434 , \15431 , \15433 );
nand \U$6616 ( \15435 , \15428 , \15429 , \15434 );
nor \U$6617 ( \15436 , \15425 , \15435 );
nand \U$6618 ( \15437 , \15407 , \15414 , \15436 );
xnor \U$6619 ( \15438 , RIb7b9518_248, \15437 );
or \U$6620 ( \15439 , \9263 , \10621 );
or \U$6621 ( \15440 , \11270 , \10417 );
nand \U$6622 ( \15441 , \15439 , \15440 );
not \U$6623 ( \15442 , \15441 );
nand \U$6624 ( \15443 , \9269 , \10179 );
nand \U$6625 ( \15444 , \9295 , \10325 );
and \U$6626 ( \15445 , \15442 , \15443 , \15444 );
or \U$6627 ( \15446 , \9282 , \10842 );
or \U$6628 ( \15447 , \11276 , \10114 );
nand \U$6629 ( \15448 , \15446 , \15447 );
not \U$6630 ( \15449 , \15448 );
nand \U$6631 ( \15450 , \9289 , \10100 );
nand \U$6632 ( \15451 , \9286 , \15374 );
and \U$6633 ( \15452 , \15449 , \15450 , \15451 );
not \U$6634 ( \15453 , \10145 );
and \U$6635 ( \15454 , \9299 , \15453 );
not \U$6636 ( \15455 , \15454 );
not \U$6637 ( \15456 , \10260 );
and \U$6638 ( \15457 , \9302 , \15456 );
not \U$6639 ( \15458 , \15457 );
and \U$6640 ( \15459 , \10318 , \9315 );
and \U$6641 ( \15460 , \9319 , \10212 );
nor \U$6642 ( \15461 , \15459 , \15460 );
and \U$6643 ( \15462 , \15455 , \15458 , \15461 );
not \U$6644 ( \15463 , \15462 );
not \U$6645 ( \15464 , \10220 );
and \U$6646 ( \15465 , \9265 , \15464 );
not \U$6647 ( \15466 , \15465 );
nand \U$6648 ( \15467 , \9310 , \10290 );
not \U$6649 ( \15468 , \10170 );
and \U$6650 ( \15469 , \9272 , \15468 );
not \U$6651 ( \15470 , \10074 );
and \U$6652 ( \15471 , \9297 , \15470 );
nor \U$6653 ( \15472 , \15469 , \15471 );
nand \U$6654 ( \15473 , \15466 , \15467 , \15472 );
nor \U$6655 ( \15474 , \15463 , \15473 );
nand \U$6656 ( \15475 , \15445 , \15452 , \15474 );
xnor \U$6657 ( \15476 , \15475 , \9327 );
or \U$6658 ( \15477 , \9395 , \10242 );
or \U$6659 ( \15478 , \11230 , \10154 );
nand \U$6660 ( \15479 , \15477 , \15478 );
not \U$6661 ( \15480 , \15479 );
nand \U$6662 ( \15481 , \9401 , \10179 );
nand \U$6663 ( \15482 , \9427 , \10325 );
and \U$6664 ( \15483 , \15480 , \15481 , \15482 );
or \U$6665 ( \15484 , \9415 , \10842 );
or \U$6666 ( \15485 , \10455 , \10114 );
nand \U$6667 ( \15486 , \15484 , \15485 );
not \U$6668 ( \15487 , \15486 );
nand \U$6669 ( \15488 , \9421 , \10100 );
nand \U$6670 ( \15489 , \9418 , \15374 );
and \U$6671 ( \15490 , \15487 , \15488 , \15489 );
not \U$6672 ( \15491 , \10145 );
and \U$6673 ( \15492 , \9432 , \15491 );
not \U$6674 ( \15493 , \15492 );
not \U$6675 ( \15494 , \10208 );
and \U$6676 ( \15495 , \9435 , \15494 );
not \U$6677 ( \15496 , \15495 );
and \U$6678 ( \15497 , \10318 , \9449 );
and \U$6679 ( \15498 , \9453 , \10212 );
nor \U$6680 ( \15499 , \15497 , \15498 );
and \U$6681 ( \15500 , \15493 , \15496 , \15499 );
not \U$6682 ( \15501 , \15500 );
not \U$6683 ( \15502 , \10165 );
and \U$6684 ( \15503 , \9397 , \15502 );
not \U$6685 ( \15504 , \15503 );
nand \U$6686 ( \15505 , \9444 , \10290 );
not \U$6687 ( \15506 , \10279 );
and \U$6688 ( \15507 , \9404 , \15506 );
not \U$6689 ( \15508 , \10224 );
and \U$6690 ( \15509 , \9430 , \15508 );
nor \U$6691 ( \15510 , \15507 , \15509 );
nand \U$6692 ( \15511 , \15504 , \15505 , \15510 );
nor \U$6693 ( \15512 , \15501 , \15511 );
nand \U$6694 ( \15513 , \15483 , \15490 , \15512 );
xnor \U$6695 ( \15514 , \15513 , \9460 );
nor \U$6696 ( \15515 , \15476 , \15514 );
nand \U$6697 ( \15516 , \15400 , \15438 , \15515 );
not \U$6698 ( \15517 , \15516 );
or \U$6699 ( \15518 , \8828 , \10242 );
or \U$6700 ( \15519 , \11565 , \10154 );
nand \U$6701 ( \15520 , \15518 , \15519 );
not \U$6702 ( \15521 , \15520 );
nand \U$6703 ( \15522 , \8852 , \10179 );
nand \U$6704 ( \15523 , \8904 , \10325 );
and \U$6705 ( \15524 , \15521 , \15522 , \15523 );
or \U$6706 ( \15525 , \8882 , \10842 );
or \U$6707 ( \15526 , \12351 , \10114 );
nand \U$6708 ( \15527 , \15525 , \15526 );
not \U$6709 ( \15528 , \15527 );
nand \U$6710 ( \15529 , \8896 , \10100 );
nand \U$6711 ( \15530 , \8893 , \15374 );
and \U$6712 ( \15531 , \15528 , \15529 , \15530 );
not \U$6713 ( \15532 , \10145 );
and \U$6714 ( \15533 , \8921 , \15532 );
not \U$6715 ( \15534 , \15533 );
not \U$6716 ( \15535 , \10208 );
and \U$6717 ( \15536 , \8927 , \15535 );
not \U$6718 ( \15537 , \15536 );
and \U$6719 ( \15538 , \10318 , \8947 );
and \U$6720 ( \15539 , \8953 , \10212 );
nor \U$6721 ( \15540 , \15538 , \15539 );
and \U$6722 ( \15541 , \15534 , \15537 , \15540 );
not \U$6723 ( \15542 , \15541 );
not \U$6724 ( \15543 , \10165 );
and \U$6725 ( \15544 , \8843 , \15543 );
not \U$6726 ( \15545 , \15544 );
nand \U$6727 ( \15546 , \8940 , \10290 );
not \U$6728 ( \15547 , \10279 );
and \U$6729 ( \15548 , \8860 , \15547 );
not \U$6730 ( \15549 , \10340 );
and \U$6731 ( \15550 , \8915 , \15549 );
nor \U$6732 ( \15551 , \15548 , \15550 );
nand \U$6733 ( \15552 , \15545 , \15546 , \15551 );
nor \U$6734 ( \15553 , \15542 , \15552 );
nand \U$6735 ( \15554 , \15524 , \15531 , \15553 );
xnor \U$6736 ( \15555 , \15554 , \8964 );
or \U$6737 ( \15556 , \9047 , \10159 );
or \U$6738 ( \15557 , \11452 , \10190 );
nand \U$6739 ( \15558 , \15556 , \15557 );
not \U$6740 ( \15559 , \15558 );
nand \U$6741 ( \15560 , \9054 , \10179 );
nand \U$6742 ( \15561 , \9081 , \10325 );
and \U$6743 ( \15562 , \15559 , \15560 , \15561 );
or \U$6744 ( \15563 , \9068 , \10842 );
or \U$6745 ( \15564 , \11458 , \10114 );
nand \U$6746 ( \15565 , \15563 , \15564 );
not \U$6747 ( \15566 , \15565 );
nand \U$6748 ( \15567 , \9075 , \10100 );
nand \U$6749 ( \15568 , \9072 , \15374 );
and \U$6750 ( \15569 , \15566 , \15567 , \15568 );
not \U$6751 ( \15570 , \10147 );
and \U$6752 ( \15571 , \9089 , \15570 );
not \U$6753 ( \15572 , \15571 );
not \U$6754 ( \15573 , \10118 );
and \U$6755 ( \15574 , \9093 , \15573 );
not \U$6756 ( \15575 , \15574 );
and \U$6757 ( \15576 , \10318 , \9107 );
and \U$6758 ( \15577 , \9112 , \10212 );
nor \U$6759 ( \15578 , \15576 , \15577 );
and \U$6760 ( \15579 , \15572 , \15575 , \15578 );
not \U$6761 ( \15580 , \15579 );
not \U$6762 ( \15581 , \10271 );
and \U$6763 ( \15582 , \9049 , \15581 );
not \U$6764 ( \15583 , \15582 );
nand \U$6765 ( \15584 , \9102 , \10290 );
not \U$6766 ( \15585 , \10228 );
and \U$6767 ( \15586 , \9057 , \15585 );
not \U$6768 ( \15587 , \10224 );
and \U$6769 ( \15588 , \9085 , \15587 );
nor \U$6770 ( \15589 , \15586 , \15588 );
nand \U$6771 ( \15590 , \15583 , \15584 , \15589 );
nor \U$6772 ( \15591 , \15580 , \15590 );
nand \U$6773 ( \15592 , \15562 , \15569 , \15591 );
xnor \U$6774 ( \15593 , \15592 , \9119 );
nor \U$6775 ( \15594 , \15555 , \15593 );
or \U$6776 ( \15595 , \9332 , \10621 );
or \U$6777 ( \15596 , \11393 , \10417 );
nand \U$6778 ( \15597 , \15595 , \15596 );
not \U$6779 ( \15598 , \15597 );
nand \U$6780 ( \15599 , \9338 , \10179 );
nand \U$6781 ( \15600 , \9361 , \10325 );
and \U$6782 ( \15601 , \15598 , \15599 , \15600 );
or \U$6783 ( \15602 , \12139 , \10195 );
or \U$6784 ( \15603 , \12141 , \10198 );
nand \U$6785 ( \15604 , \15602 , \15603 );
not \U$6786 ( \15605 , \15604 );
nand \U$6787 ( \15606 , \9356 , \10100 );
nand \U$6788 ( \15607 , \9353 , \15374 );
and \U$6789 ( \15608 , \15605 , \15606 , \15607 );
not \U$6790 ( \15609 , \10145 );
and \U$6791 ( \15610 , \9366 , \15609 );
not \U$6792 ( \15611 , \15610 );
not \U$6793 ( \15612 , \10260 );
and \U$6794 ( \15613 , \9369 , \15612 );
not \U$6795 ( \15614 , \15613 );
and \U$6796 ( \15615 , \10318 , \9385 );
and \U$6797 ( \15616 , \9377 , \10212 );
nor \U$6798 ( \15617 , \15615 , \15616 );
and \U$6799 ( \15618 , \15611 , \15614 , \15617 );
not \U$6800 ( \15619 , \15618 );
not \U$6801 ( \15620 , \10220 );
and \U$6802 ( \15621 , \9334 , \15620 );
not \U$6803 ( \15622 , \15621 );
nand \U$6804 ( \15623 , \9380 , \10290 );
not \U$6805 ( \15624 , \10170 );
and \U$6806 ( \15625 , \9341 , \15624 );
not \U$6807 ( \15626 , \10275 );
and \U$6808 ( \15627 , \9364 , \15626 );
nor \U$6809 ( \15628 , \15625 , \15627 );
nand \U$6810 ( \15629 , \15622 , \15623 , \15628 );
nor \U$6811 ( \15630 , \15619 , \15629 );
nand \U$6812 ( \15631 , \15601 , \15608 , \15630 );
xnor \U$6813 ( \15632 , \15631 , \9392 );
or \U$6814 ( \15633 , \9122 , \10242 );
or \U$6815 ( \15634 , \11410 , \10154 );
nand \U$6816 ( \15635 , \15633 , \15634 );
not \U$6817 ( \15636 , \15635 );
nand \U$6818 ( \15637 , \9129 , \10179 );
nand \U$6819 ( \15638 , \9155 , \10325 );
and \U$6820 ( \15639 , \15636 , \15637 , \15638 );
or \U$6821 ( \15640 , \9143 , \10195 );
or \U$6822 ( \15641 , \11416 , \10198 );
nand \U$6823 ( \15642 , \15640 , \15641 );
not \U$6824 ( \15643 , \15642 );
nand \U$6825 ( \15644 , \9150 , \10100 );
nand \U$6826 ( \15645 , \9147 , \15374 );
and \U$6827 ( \15646 , \15643 , \15644 , \15645 );
not \U$6828 ( \15647 , \10358 );
and \U$6829 ( \15648 , \9159 , \15647 );
not \U$6830 ( \15649 , \15648 );
not \U$6831 ( \15650 , \10208 );
and \U$6832 ( \15651 , \9163 , \15650 );
not \U$6833 ( \15652 , \15651 );
and \U$6834 ( \15653 , \10318 , \9176 );
and \U$6835 ( \15654 , \9180 , \10212 );
nor \U$6836 ( \15655 , \15653 , \15654 );
and \U$6837 ( \15656 , \15649 , \15652 , \15655 );
not \U$6838 ( \15657 , \15656 );
not \U$6839 ( \15658 , \10165 );
and \U$6840 ( \15659 , \9124 , \15658 );
not \U$6841 ( \15660 , \15659 );
nand \U$6842 ( \15661 , \9172 , \10290 );
not \U$6843 ( \15662 , \10279 );
and \U$6844 ( \15663 , \9132 , \15662 );
not \U$6845 ( \15664 , \10275 );
and \U$6846 ( \15665 , \9157 , \15664 );
nor \U$6847 ( \15666 , \15663 , \15665 );
nand \U$6848 ( \15667 , \15660 , \15661 , \15666 );
nor \U$6849 ( \15668 , \15657 , \15667 );
nand \U$6850 ( \15669 , \15639 , \15646 , \15668 );
xnor \U$6851 ( \15670 , \15669 , \9188 );
nor \U$6852 ( \15671 , \15632 , \15670 );
and \U$6853 ( \15672 , \15517 , \15594 , \15671 );
not \U$6854 ( \15673 , \10165 );
and \U$6855 ( \15674 , \15673 , \9816 );
and \U$6856 ( \15675 , \10290 , \9813 );
nor \U$6857 ( \15676 , \15674 , \15675 );
not \U$6858 ( \15677 , \10074 );
and \U$6859 ( \15678 , \9808 , \15677 );
not \U$6860 ( \15679 , \10170 );
and \U$6861 ( \15680 , \9805 , \15679 );
nor \U$6862 ( \15681 , \15678 , \15680 );
or \U$6863 ( \15682 , \11494 , \10195 );
or \U$6864 ( \15683 , \9798 , \10198 );
nand \U$6865 ( \15684 , \15682 , \15683 );
not \U$6866 ( \15685 , \15684 );
nand \U$6867 ( \15686 , \9794 , \10100 );
nand \U$6868 ( \15687 , \9790 , \15374 );
and \U$6869 ( \15688 , \15685 , \15686 , \15687 );
nand \U$6870 ( \15689 , \15676 , \15681 , \15688 );
and \U$6871 ( \15690 , \9847 , \10160 );
not \U$6872 ( \15691 , \10190 );
and \U$6873 ( \15692 , \9850 , \15691 );
nor \U$6874 ( \15693 , \15690 , \15692 );
and \U$6875 ( \15694 , \10236 , \9839 );
and \U$6876 ( \15695 , \9842 , \10143 );
nor \U$6877 ( \15696 , \15694 , \15695 );
nand \U$6878 ( \15697 , \9822 , \10133 );
nand \U$6879 ( \15698 , \9826 , \10318 );
nand \U$6880 ( \15699 , \15697 , \15698 );
not \U$6881 ( \15700 , \15699 );
nand \U$6882 ( \15701 , \10119 , \9830 );
nand \U$6883 ( \15702 , \9833 , \10146 );
and \U$6884 ( \15703 , \15700 , \15701 , \15702 );
nand \U$6885 ( \15704 , \15693 , \15696 , \15703 );
nor \U$6886 ( \15705 , \15689 , \15704 );
xnor \U$6887 ( \15706 , \15705 , \9857 );
nand \U$6888 ( \15707 , \9892 , \10133 );
nand \U$6889 ( \15708 , \9897 , \10138 );
nand \U$6890 ( \15709 , \15707 , \15708 );
not \U$6891 ( \15710 , \15709 );
nand \U$6892 ( \15711 , \10119 , \9902 );
nand \U$6893 ( \15712 , \9905 , \10146 );
and \U$6894 ( \15713 , \15710 , \15711 , \15712 );
nand \U$6895 ( \15714 , \9910 , \10179 );
nand \U$6896 ( \15715 , \9913 , \10143 );
nand \U$6897 ( \15716 , \15714 , \15715 );
not \U$6898 ( \15717 , \9917 );
or \U$6899 ( \15718 , \15717 , \10159 );
or \U$6900 ( \15719 , \9921 , \10190 );
nand \U$6901 ( \15720 , \15718 , \15719 );
nor \U$6902 ( \15721 , \15716 , \15720 );
not \U$6903 ( \15722 , \10080 );
and \U$6904 ( \15723 , \9859 , \15722 );
not \U$6905 ( \15724 , \15723 );
not \U$6906 ( \15725 , \10299 );
and \U$6907 ( \15726 , \9864 , \15725 );
not \U$6908 ( \15727 , \15726 );
not \U$6909 ( \15728 , \10114 );
and \U$6910 ( \15729 , \9867 , \15728 );
not \U$6911 ( \15730 , \10842 );
and \U$6912 ( \15731 , \9871 , \15730 );
nor \U$6913 ( \15732 , \15729 , \15731 );
and \U$6914 ( \15733 , \15724 , \15727 , \15732 );
not \U$6915 ( \15734 , \15733 );
nand \U$6916 ( \15735 , \9881 , \10127 );
not \U$6917 ( \15736 , \10271 );
and \U$6918 ( \15737 , \9886 , \15736 );
not \U$6919 ( \15738 , \15737 );
not \U$6920 ( \15739 , \10224 );
and \U$6921 ( \15740 , \9877 , \15739 );
not \U$6922 ( \15741 , \10228 );
and \U$6923 ( \15742 , \9874 , \15741 );
nor \U$6924 ( \15743 , \15740 , \15742 );
nand \U$6925 ( \15744 , \15735 , \15738 , \15743 );
nor \U$6926 ( \15745 , \15734 , \15744 );
nand \U$6927 ( \15746 , \15713 , \15721 , \15745 );
xnor \U$6928 ( \15747 , RIb7a0c48_261, \15746 );
nand \U$6929 ( \15748 , \9968 , \10212 );
nand \U$6930 ( \15749 , \9965 , \10318 );
nand \U$6931 ( \15750 , \15748 , \15749 );
not \U$6932 ( \15751 , \15750 );
nand \U$6933 ( \15752 , \10119 , \10709 );
nand \U$6934 ( \15753 , \9959 , \10146 );
and \U$6935 ( \15754 , \15751 , \15752 , \15753 );
nand \U$6936 ( \15755 , \9977 , \10179 );
nand \U$6937 ( \15756 , \9975 , \10325 );
nand \U$6938 ( \15757 , \15755 , \15756 );
not \U$6939 ( \15758 , \9982 );
or \U$6940 ( \15759 , \15758 , \10621 );
or \U$6941 ( \15760 , \12282 , \10417 );
nand \U$6942 ( \15761 , \15759 , \15760 );
nor \U$6943 ( \15762 , \15757 , \15761 );
not \U$6944 ( \15763 , \10080 );
and \U$6945 ( \15764 , \9951 , \15763 );
not \U$6946 ( \15765 , \15764 );
not \U$6947 ( \15766 , \10346 );
and \U$6948 ( \15767 , \9954 , \15766 );
not \U$6949 ( \15768 , \15767 );
not \U$6950 ( \15769 , \10114 );
and \U$6951 ( \15770 , \9944 , \15769 );
not \U$6952 ( \15771 , \10842 );
and \U$6953 ( \15772 , \9947 , \15771 );
nor \U$6954 ( \15773 , \15770 , \15772 );
and \U$6955 ( \15774 , \15765 , \15768 , \15773 );
not \U$6956 ( \15775 , \15774 );
nand \U$6957 ( \15776 , \9936 , \10290 );
not \U$6958 ( \15777 , \10220 );
and \U$6959 ( \15778 , \9939 , \15777 );
not \U$6960 ( \15779 , \15778 );
not \U$6961 ( \15780 , \10275 );
and \U$6962 ( \15781 , \9932 , \15780 );
not \U$6963 ( \15782 , \10170 );
and \U$6964 ( \15783 , \9929 , \15782 );
nor \U$6965 ( \15784 , \15781 , \15783 );
nand \U$6966 ( \15785 , \15776 , \15779 , \15784 );
nor \U$6967 ( \15786 , \15775 , \15785 );
nand \U$6968 ( \15787 , \15754 , \15762 , \15786 );
xnor \U$6969 ( \15788 , \15787 , \9990 );
nand \U$6970 ( \15789 , \10034 , \10133 );
nand \U$6971 ( \15790 , \10030 , \10138 );
nand \U$6972 ( \15791 , \15789 , \15790 );
not \U$6973 ( \15792 , \15791 );
nand \U$6974 ( \15793 , \10119 , \10027 );
nand \U$6975 ( \15794 , \10025 , \10146 );
and \U$6976 ( \15795 , \15792 , \15793 , \15794 );
nand \U$6977 ( \15796 , \10043 , \10179 );
nand \U$6978 ( \15797 , \10041 , \10325 );
nand \U$6979 ( \15798 , \15796 , \15797 );
not \U$6980 ( \15799 , \10047 );
or \U$6981 ( \15800 , \15799 , \10242 );
or \U$6982 ( \15801 , \11674 , \10154 );
nand \U$6983 ( \15802 , \15800 , \15801 );
nor \U$6984 ( \15803 , \15798 , \15802 );
nand \U$6985 ( \15804 , \10017 , \10290 );
not \U$6986 ( \15805 , \10165 );
and \U$6987 ( \15806 , \10020 , \15805 );
not \U$6988 ( \15807 , \15806 );
not \U$6989 ( \15808 , \10074 );
and \U$6990 ( \15809 , \15808 , \10012 );
not \U$6991 ( \15810 , \10279 );
and \U$6992 ( \15811 , \10009 , \15810 );
nor \U$6993 ( \15812 , \15809 , \15811 );
nand \U$6994 ( \15813 , \15804 , \15807 , \15812 );
not \U$6995 ( \15814 , \10080 );
and \U$6996 ( \15815 , \10001 , \15814 );
not \U$6997 ( \15816 , \15815 );
not \U$6998 ( \15817 , \10099 );
and \U$6999 ( \15818 , \10004 , \15817 );
not \U$7000 ( \15819 , \15818 );
not \U$7001 ( \15820 , \10198 );
and \U$7002 ( \15821 , \15820 , \9992 );
not \U$7003 ( \15822 , \10195 );
and \U$7004 ( \15823 , \15822 , \9996 );
nor \U$7005 ( \15824 , \15821 , \15823 );
and \U$7006 ( \15825 , \15816 , \15819 , \15824 );
not \U$7007 ( \15826 , \15825 );
nor \U$7008 ( \15827 , \15813 , \15826 );
nand \U$7009 ( \15828 , \15795 , \15803 , \15827 );
xnor \U$7010 ( \15829 , \15828 , \10055 );
nor \U$7011 ( \15830 , \15788 , \15829 );
nand \U$7012 ( \15831 , \15706 , \15747 , \15830 );
not \U$7013 ( \15832 , \15831 );
nand \U$7014 ( \15833 , \9619 , \10133 );
nand \U$7015 ( \15834 , \9622 , \10318 );
nand \U$7016 ( \15835 , \15833 , \15834 );
not \U$7017 ( \15836 , \15835 );
nand \U$7018 ( \15837 , \10119 , \9628 );
nand \U$7019 ( \15838 , \9631 , \10146 );
and \U$7020 ( \15839 , \15836 , \15837 , \15838 );
nand \U$7021 ( \15840 , \9636 , \10179 );
nand \U$7022 ( \15841 , \9639 , \10325 );
nand \U$7023 ( \15842 , \15840 , \15841 );
not \U$7024 ( \15843 , \9643 );
or \U$7025 ( \15844 , \15843 , \10159 );
or \U$7026 ( \15845 , \9647 , \10190 );
nand \U$7027 ( \15846 , \15844 , \15845 );
nor \U$7028 ( \15847 , \15842 , \15846 );
not \U$7029 ( \15848 , \10080 );
and \U$7030 ( \15849 , \9587 , \15848 );
not \U$7031 ( \15850 , \15849 );
not \U$7032 ( \15851 , \10099 );
and \U$7033 ( \15852 , \9593 , \15851 );
not \U$7034 ( \15853 , \15852 );
not \U$7035 ( \15854 , \10114 );
and \U$7036 ( \15855 , \9596 , \15854 );
not \U$7037 ( \15856 , \10842 );
and \U$7038 ( \15857 , \9600 , \15856 );
nor \U$7039 ( \15858 , \15855 , \15857 );
and \U$7040 ( \15859 , \15850 , \15853 , \15858 );
not \U$7041 ( \15860 , \15859 );
nand \U$7042 ( \15861 , \9610 , \10290 );
not \U$7043 ( \15862 , \10271 );
and \U$7044 ( \15863 , \9613 , \15862 );
not \U$7045 ( \15864 , \15863 );
not \U$7046 ( \15865 , \10224 );
and \U$7047 ( \15866 , \9606 , \15865 );
not \U$7048 ( \15867 , \10228 );
and \U$7049 ( \15868 , \9603 , \15867 );
nor \U$7050 ( \15869 , \15866 , \15868 );
nand \U$7051 ( \15870 , \15861 , \15864 , \15869 );
nor \U$7052 ( \15871 , \15860 , \15870 );
nand \U$7053 ( \15872 , \15839 , \15847 , \15871 );
xnor \U$7054 ( \15873 , \15872 , \9653 );
nand \U$7055 ( \15874 , \9655 , \10179 );
nand \U$7056 ( \15875 , \9660 , \10325 );
nand \U$7057 ( \15876 , \15874 , \15875 );
not \U$7058 ( \15877 , \9664 );
or \U$7059 ( \15878 , \15877 , \10621 );
or \U$7060 ( \15879 , \9668 , \10417 );
nand \U$7061 ( \15880 , \15878 , \15879 );
nor \U$7062 ( \15881 , \15876 , \15880 );
or \U$7063 ( \15882 , \9676 , \10195 );
or \U$7064 ( \15883 , \11923 , \10198 );
nand \U$7065 ( \15884 , \15882 , \15883 );
not \U$7066 ( \15885 , \15884 );
nand \U$7067 ( \15886 , \9682 , \10100 );
nand \U$7068 ( \15887 , \9679 , \15374 );
and \U$7069 ( \15888 , \15885 , \15886 , \15887 );
not \U$7070 ( \15889 , \10145 );
and \U$7071 ( \15890 , \9687 , \15889 );
not \U$7072 ( \15891 , \15890 );
not \U$7073 ( \15892 , \10118 );
and \U$7074 ( \15893 , \9690 , \15892 );
not \U$7075 ( \15894 , \15893 );
and \U$7076 ( \15895 , \10212 , \9695 );
and \U$7077 ( \15896 , \9692 , \10318 );
nor \U$7078 ( \15897 , \15895 , \15896 );
and \U$7079 ( \15898 , \15891 , \15894 , \15897 );
not \U$7080 ( \15899 , \15898 );
nand \U$7081 ( \15900 , \9713 , \10290 );
not \U$7082 ( \15901 , \10220 );
and \U$7083 ( \15902 , \9710 , \15901 );
not \U$7084 ( \15903 , \15902 );
not \U$7085 ( \15904 , \10275 );
and \U$7086 ( \15905 , \9701 , \15904 );
not \U$7087 ( \15906 , \10170 );
and \U$7088 ( \15907 , \9706 , \15906 );
nor \U$7089 ( \15908 , \15905 , \15907 );
nand \U$7090 ( \15909 , \15900 , \15903 , \15908 );
nor \U$7091 ( \15910 , \15899 , \15909 );
nand \U$7092 ( \15911 , \15881 , \15888 , \15910 );
xnor \U$7093 ( \15912 , \15911 , \9719 );
nor \U$7094 ( \15913 , \15873 , \15912 );
nand \U$7095 ( \15914 , \9721 , \10179 );
nand \U$7096 ( \15915 , \9724 , \10325 );
nand \U$7097 ( \15916 , \15914 , \15915 );
not \U$7098 ( \15917 , \9728 );
or \U$7099 ( \15918 , \15917 , \10242 );
or \U$7100 ( \15919 , \9732 , \10154 );
nand \U$7101 ( \15920 , \15918 , \15919 );
nor \U$7102 ( \15921 , \15916 , \15920 );
or \U$7103 ( \15922 , \9740 , \10195 );
or \U$7104 ( \15923 , \11876 , \10198 );
nand \U$7105 ( \15924 , \15922 , \15923 );
not \U$7106 ( \15925 , \15924 );
nand \U$7107 ( \15926 , \9747 , \10100 );
nand \U$7108 ( \15927 , \9744 , \15374 );
and \U$7109 ( \15928 , \15925 , \15926 , \15927 );
not \U$7110 ( \15929 , \10145 );
and \U$7111 ( \15930 , \9752 , \15929 );
not \U$7112 ( \15931 , \15930 );
not \U$7113 ( \15932 , \10260 );
and \U$7114 ( \15933 , \9755 , \15932 );
not \U$7115 ( \15934 , \15933 );
and \U$7116 ( \15935 , \10212 , \9763 );
and \U$7117 ( \15936 , \9759 , \10318 );
nor \U$7118 ( \15937 , \15935 , \15936 );
and \U$7119 ( \15938 , \15931 , \15934 , \15937 );
not \U$7120 ( \15939 , \15938 );
nand \U$7121 ( \15940 , \9779 , \10290 );
not \U$7122 ( \15941 , \10165 );
and \U$7123 ( \15942 , \9776 , \15941 );
not \U$7124 ( \15943 , \15942 );
not \U$7125 ( \15944 , \10340 );
and \U$7126 ( \15945 , \9769 , \15944 );
not \U$7127 ( \15946 , \10279 );
and \U$7128 ( \15947 , \9772 , \15946 );
nor \U$7129 ( \15948 , \15945 , \15947 );
nand \U$7130 ( \15949 , \15940 , \15943 , \15948 );
nor \U$7131 ( \15950 , \15939 , \15949 );
nand \U$7132 ( \15951 , \15921 , \15928 , \15950 );
xnor \U$7133 ( \15952 , \15951 , \9786 );
nand \U$7134 ( \15953 , \9551 , \10133 );
nand \U$7135 ( \15954 , \9554 , \10138 );
nand \U$7136 ( \15955 , \15953 , \15954 );
not \U$7137 ( \15956 , \15955 );
nand \U$7138 ( \15957 , \10119 , \9560 );
nand \U$7139 ( \15958 , \9563 , \10146 );
and \U$7140 ( \15959 , \15956 , \15957 , \15958 );
nand \U$7141 ( \15960 , \9568 , \10179 );
nand \U$7142 ( \15961 , \9571 , \10325 );
nand \U$7143 ( \15962 , \15960 , \15961 );
not \U$7144 ( \15963 , \9575 );
or \U$7145 ( \15964 , \15963 , \10159 );
or \U$7146 ( \15965 , \9579 , \10190 );
nand \U$7147 ( \15966 , \15964 , \15965 );
nor \U$7148 ( \15967 , \15962 , \15966 );
not \U$7149 ( \15968 , \10080 );
and \U$7150 ( \15969 , \9518 , \15968 );
not \U$7151 ( \15970 , \15969 );
not \U$7152 ( \15971 , \10299 );
and \U$7153 ( \15972 , \9523 , \15971 );
not \U$7154 ( \15973 , \15972 );
not \U$7155 ( \15974 , \10198 );
and \U$7156 ( \15975 , \9526 , \15974 );
not \U$7157 ( \15976 , \10093 );
and \U$7158 ( \15977 , \9530 , \15976 );
nor \U$7159 ( \15978 , \15975 , \15977 );
and \U$7160 ( \15979 , \15970 , \15973 , \15978 );
not \U$7161 ( \15980 , \15979 );
nand \U$7162 ( \15981 , \9542 , \10290 );
not \U$7163 ( \15982 , \10271 );
and \U$7164 ( \15983 , \9545 , \15982 );
not \U$7165 ( \15984 , \15983 );
not \U$7166 ( \15985 , \10340 );
and \U$7167 ( \15986 , \9536 , \15985 );
not \U$7168 ( \15987 , \10228 );
and \U$7169 ( \15988 , \9533 , \15987 );
nor \U$7170 ( \15989 , \15986 , \15988 );
nand \U$7171 ( \15990 , \15981 , \15984 , \15989 );
nor \U$7172 ( \15991 , \15980 , \15990 );
nand \U$7173 ( \15992 , \15959 , \15967 , \15991 );
xnor \U$7174 ( \15993 , \15992 , \9585 );
nor \U$7175 ( \15994 , \15952 , \15993 );
and \U$7176 ( \15995 , \15832 , \15913 , \15994 );
nand \U$7177 ( \15996 , \15361 , \15672 , \15995 );
not \U$7178 ( \15997 , \15996 );
not \U$7179 ( \15998 , \15997 );
or \U$7180 ( \15999 , \15317 , \15998 );
not \U$7181 ( \16000 , \15999 );
nand \U$7182 ( \16001 , \15317 , \15997 );
not \U$7183 ( \16002 , \16001 );
or \U$7184 ( \16003 , \16000 , \16002 );
not \U$7185 ( \16004 , \16003 );
not \U$7186 ( \16005 , \16004 );
and \U$7187 ( \16006 , \15292 , \16005 );
not \U$7188 ( \16007 , \10931 );
buf \U$7189 ( \16008 , \12454 );
buf \U$7190 ( \16009 , \12456 );
buf \U$7191 ( \16010 , \12458 );
buf \U$7192 ( \16011 , \8835 );
and \U$7193 ( \16012 , \16010 , \16011 );
or \U$7194 ( \16013 , \16009 , \16012 );
xnor \U$7195 ( \16014 , \16008 , \16013 );
buf \U$7196 ( \16015 , \16014 );
not \U$7197 ( \16016 , \16015 );
xnor \U$7198 ( \16017 , \16009 , \16012 );
buf \U$7199 ( \16018 , \16017 );
xor \U$7200 ( \16019 , \16010 , \16011 );
buf \U$7201 ( \16020 , \16019 );
not \U$7202 ( \16021 , \16011 );
buf \U$7203 ( \16022 , \16021 );
nor \U$7204 ( \16023 , \16018 , \16020 , \16022 );
and \U$7205 ( \16024 , \16016 , \16023 );
buf \U$7206 ( \16025 , RIea91330_6888);
or \U$7207 ( \16026 , \16008 , \16013 );
xor \U$7208 ( \16027 , \16025 , \16026 );
buf \U$7209 ( \16028 , \16027 );
not \U$7210 ( \16029 , \16028 );
or \U$7211 ( \16030 , \16024 , \16029 );
and \U$7212 ( \16031 , \16025 , \16026 );
buf \U$7213 ( \16032 , \16031 );
not \U$7214 ( \16033 , \16032 );
nand \U$7215 ( \16034 , \16030 , \16033 );
or \U$7216 ( \16035 , \9492 , \11051 );
or \U$7217 ( \16036 , \9494 , \11075 );
nand \U$7218 ( \16037 , \16035 , \16036 );
or \U$7219 ( \16038 , \9498 , \11044 );
or \U$7220 ( \16039 , \9500 , \11327 );
nand \U$7221 ( \16040 , \16038 , \16039 );
nor \U$7222 ( \16041 , \16037 , \16040 );
or \U$7223 ( \16042 , \9504 , \11014 );
or \U$7224 ( \16043 , \9506 , \11102 );
nand \U$7225 ( \16044 , \16042 , \16043 );
or \U$7226 ( \16045 , \9509 , \11143 );
not \U$7227 ( \16046 , \10962 );
or \U$7228 ( \16047 , \9511 , \16046 );
nand \U$7229 ( \16048 , \16045 , \16047 );
nor \U$7230 ( \16049 , \16044 , \16048 );
not \U$7231 ( \16050 , \10954 );
or \U$7232 ( \16051 , \9467 , \16050 );
not \U$7233 ( \16052 , \11374 );
or \U$7234 ( \16053 , \9463 , \16052 );
not \U$7235 ( \16054 , \10935 );
and \U$7236 ( \16055 , \9472 , \16054 );
not \U$7237 ( \16056 , \10944 );
and \U$7238 ( \16057 , \9476 , \16056 );
nor \U$7239 ( \16058 , \16055 , \16057 );
nand \U$7240 ( \16059 , \16051 , \16053 , \16058 );
not \U$7241 ( \16060 , \11033 );
or \U$7242 ( \16061 , \9485 , \16060 );
not \U$7243 ( \16062 , \11020 );
or \U$7244 ( \16063 , \9487 , \16062 );
not \U$7245 ( \16064 , \9480 );
and \U$7246 ( \16065 , \16064 , \11039 );
and \U$7247 ( \16066 , \11010 , \12557 );
nor \U$7248 ( \16067 , \16065 , \16066 );
nand \U$7249 ( \16068 , \16061 , \16063 , \16067 );
nor \U$7250 ( \16069 , \16059 , \16068 );
nand \U$7251 ( \16070 , \16041 , \16049 , \16069 );
not \U$7252 ( \16071 , \16070 );
or \U$7253 ( \16072 , \9537 , \11131 );
or \U$7254 ( \16073 , \9543 , \11038 );
nand \U$7255 ( \16074 , \16072 , \16073 );
or \U$7256 ( \16075 , \9546 , \11009 );
or \U$7257 ( \16076 , \9534 , \11014 );
nand \U$7258 ( \16077 , \16075 , \16076 );
nor \U$7259 ( \16078 , \16074 , \16077 );
or \U$7260 ( \16079 , \13658 , \11065 );
or \U$7261 ( \16080 , \9527 , \10970 );
nand \U$7262 ( \16081 , \16079 , \16080 );
or \U$7263 ( \16082 , \9519 , \11114 );
or \U$7264 ( \16083 , \14434 , \16046 );
nand \U$7265 ( \16084 , \16082 , \16083 );
nor \U$7266 ( \16085 , \16081 , \16084 );
nand \U$7267 ( \16086 , \16078 , \16085 );
not \U$7268 ( \16087 , \16086 );
or \U$7269 ( \16088 , \9569 , \10979 );
or \U$7270 ( \16089 , \9572 , \11182 );
nand \U$7271 ( \16090 , \16088 , \16089 );
or \U$7272 ( \16091 , \9579 , \11143 );
or \U$7273 ( \16092 , \11589 , \11019 );
nand \U$7274 ( \16093 , \16091 , \16092 );
nor \U$7275 ( \16094 , \16090 , \16093 );
or \U$7276 ( \16095 , \9552 , \11099 );
or \U$7277 ( \16096 , \9557 , \11047 );
nand \U$7278 ( \16097 , \16095 , \16096 );
or \U$7279 ( \16098 , \9564 , \10996 );
or \U$7280 ( \16099 , \11582 , \11327 );
nand \U$7281 ( \16100 , \16098 , \16099 );
nor \U$7282 ( \16101 , \16097 , \16100 );
and \U$7283 ( \16102 , \16087 , \16094 , \16101 );
xnor \U$7284 ( \16103 , \16102 , \9585 );
or \U$7285 ( \16104 , \9607 , \11131 );
or \U$7286 ( \16105 , \9611 , \10973 );
nand \U$7287 ( \16106 , \16104 , \16105 );
or \U$7288 ( \16107 , \9614 , \11009 );
or \U$7289 ( \16108 , \9604 , \11014 );
nand \U$7290 ( \16109 , \16107 , \16108 );
nor \U$7291 ( \16110 , \16106 , \16109 );
or \U$7292 ( \16111 , \13538 , \10955 );
or \U$7293 ( \16112 , \9597 , \10970 );
nand \U$7294 ( \16113 , \16111 , \16112 );
or \U$7295 ( \16114 , \9588 , \10935 );
or \U$7296 ( \16115 , \12108 , \16046 );
nand \U$7297 ( \16116 , \16114 , \16115 );
nor \U$7298 ( \16117 , \16113 , \16116 );
nand \U$7299 ( \16118 , \16110 , \16117 );
not \U$7300 ( \16119 , \16118 );
or \U$7301 ( \16120 , \9637 , \11389 );
or \U$7302 ( \16121 , \9640 , \11126 );
nand \U$7303 ( \16122 , \16120 , \16121 );
or \U$7304 ( \16123 , \9647 , \11319 );
or \U$7305 ( \16124 , \11322 , \11019 );
nand \U$7306 ( \16125 , \16123 , \16124 );
nor \U$7307 ( \16126 , \16122 , \16125 );
or \U$7308 ( \16127 , \9620 , \11209 );
or \U$7309 ( \16128 , \9625 , \11102 );
nand \U$7310 ( \16129 , \16127 , \16128 );
or \U$7311 ( \16130 , \9632 , \11160 );
or \U$7312 ( \16131 , \11314 , \11327 );
nand \U$7313 ( \16132 , \16130 , \16131 );
nor \U$7314 ( \16133 , \16129 , \16132 );
and \U$7315 ( \16134 , \16119 , \16126 , \16133 );
xnor \U$7316 ( \16135 , \16134 , \9653 );
or \U$7317 ( \16136 , \11393 , \11143 );
or \U$7318 ( \16137 , \10553 , \10973 );
nand \U$7319 ( \16138 , \16136 , \16137 );
or \U$7320 ( \16139 , \9339 , \10979 );
or \U$7321 ( \16140 , \9332 , \11019 );
nand \U$7322 ( \16141 , \16139 , \16140 );
nor \U$7323 ( \16142 , \16138 , \16141 );
or \U$7324 ( \16143 , \12139 , \11065 );
or \U$7325 ( \16144 , \12141 , \11068 );
nand \U$7326 ( \16145 , \16143 , \16144 );
or \U$7327 ( \16146 , \9354 , \11061 );
or \U$7328 ( \16147 , \9357 , \10963 );
nand \U$7329 ( \16148 , \16146 , \16147 );
nor \U$7330 ( \16149 , \16145 , \16148 );
not \U$7331 ( \16150 , \11199 );
and \U$7332 ( \16151 , \9369 , \16150 );
not \U$7333 ( \16152 , \11209 );
and \U$7334 ( \16153 , \9377 , \16152 );
nor \U$7335 ( \16154 , \16151 , \16153 );
not \U$7336 ( \16155 , \11182 );
and \U$7337 ( \16156 , \9361 , \16155 );
not \U$7338 ( \16157 , \11105 );
and \U$7339 ( \16158 , \9366 , \16157 );
nor \U$7340 ( \16159 , \16156 , \16158 );
nand \U$7341 ( \16160 , \16154 , \16159 );
not \U$7342 ( \16161 , \11357 );
and \U$7343 ( \16162 , \16161 , \11174 );
and \U$7344 ( \16163 , \11015 , \9341 );
nor \U$7345 ( \16164 , \16162 , \16163 );
not \U$7346 ( \16165 , \12874 );
not \U$7347 ( \16166 , \11102 );
and \U$7348 ( \16167 , \16165 , \16166 );
and \U$7349 ( \16168 , \11010 , \9334 );
nor \U$7350 ( \16169 , \16167 , \16168 );
nand \U$7351 ( \16170 , \16164 , \16169 );
nor \U$7352 ( \16171 , \16160 , \16170 );
nand \U$7353 ( \16172 , \16142 , \16149 , \16171 );
xnor \U$7354 ( \16173 , \16172 , \9392 );
or \U$7355 ( \16174 , \11410 , \11022 );
or \U$7356 ( \16175 , \10901 , \11038 );
nand \U$7357 ( \16176 , \16174 , \16175 );
or \U$7358 ( \16177 , \9130 , \11032 );
or \U$7359 ( \16178 , \9122 , \11019 );
nand \U$7360 ( \16179 , \16177 , \16178 );
nor \U$7361 ( \16180 , \16176 , \16179 );
or \U$7362 ( \16181 , \9143 , \11118 );
or \U$7363 ( \16182 , \11416 , \11068 );
nand \U$7364 ( \16183 , \16181 , \16182 );
or \U$7365 ( \16184 , \9148 , \10935 );
or \U$7366 ( \16185 , \9151 , \10963 );
nand \U$7367 ( \16186 , \16184 , \16185 );
nor \U$7368 ( \16187 , \16183 , \16186 );
not \U$7369 ( \16188 , \11199 );
and \U$7370 ( \16189 , \9163 , \16188 );
not \U$7371 ( \16190 , \11044 );
and \U$7372 ( \16191 , \9180 , \16190 );
nor \U$7373 ( \16192 , \16189 , \16191 );
not \U$7374 ( \16193 , \11075 );
and \U$7375 ( \16194 , \9155 , \16193 );
not \U$7376 ( \16195 , \10996 );
and \U$7377 ( \16196 , \9159 , \16195 );
nor \U$7378 ( \16197 , \16194 , \16196 );
nand \U$7379 ( \16198 , \16192 , \16197 );
and \U$7380 ( \16199 , \11015 , \9132 );
and \U$7381 ( \16200 , \9157 , \11174 );
nor \U$7382 ( \16201 , \16199 , \16200 );
and \U$7383 ( \16202 , \11010 , \9124 );
and \U$7384 ( \16203 , \9176 , \16166 );
nor \U$7385 ( \16204 , \16202 , \16203 );
nand \U$7386 ( \16205 , \16201 , \16204 );
nor \U$7387 ( \16206 , \16198 , \16205 );
nand \U$7388 ( \16207 , \16180 , \16187 , \16206 );
xnor \U$7389 ( \16208 , \16207 , \9188 );
nor \U$7390 ( \16209 , \16173 , \16208 );
nand \U$7391 ( \16210 , \16103 , \16135 , \16209 );
not \U$7392 ( \16211 , \16210 );
or \U$7393 ( \16212 , \11565 , \11319 );
or \U$7394 ( \16213 , \10775 , \10973 );
nand \U$7395 ( \16214 , \16212 , \16213 );
or \U$7396 ( \16215 , \8853 , \11389 );
or \U$7397 ( \16216 , \8828 , \11019 );
nand \U$7398 ( \16217 , \16215 , \16216 );
nor \U$7399 ( \16218 , \16214 , \16217 );
or \U$7400 ( \16219 , \8882 , \11118 );
or \U$7401 ( \16220 , \12351 , \11068 );
nand \U$7402 ( \16221 , \16219 , \16220 );
or \U$7403 ( \16222 , \8894 , \11061 );
or \U$7404 ( \16223 , \8897 , \10963 );
nand \U$7405 ( \16224 , \16222 , \16223 );
nor \U$7406 ( \16225 , \16221 , \16224 );
not \U$7407 ( \16226 , \10982 );
and \U$7408 ( \16227 , \8927 , \16226 );
not \U$7409 ( \16228 , \11044 );
and \U$7410 ( \16229 , \8953 , \16228 );
nor \U$7411 ( \16230 , \16227 , \16229 );
not \U$7412 ( \16231 , \11000 );
and \U$7413 ( \16232 , \8904 , \16231 );
not \U$7414 ( \16233 , \11105 );
and \U$7415 ( \16234 , \8921 , \16233 );
nor \U$7416 ( \16235 , \16232 , \16234 );
nand \U$7417 ( \16236 , \16230 , \16235 );
not \U$7418 ( \16237 , \11533 );
and \U$7419 ( \16238 , \16237 , \11174 );
and \U$7420 ( \16239 , \11015 , \8860 );
nor \U$7421 ( \16240 , \16238 , \16239 );
not \U$7422 ( \16241 , \11545 );
and \U$7423 ( \16242 , \16241 , \16166 );
and \U$7424 ( \16243 , \11010 , \8843 );
nor \U$7425 ( \16244 , \16242 , \16243 );
nand \U$7426 ( \16245 , \16240 , \16244 );
nor \U$7427 ( \16246 , \16236 , \16245 );
nand \U$7428 ( \16247 , \16218 , \16225 , \16246 );
xnor \U$7429 ( \16248 , \16247 , \8964 );
or \U$7430 ( \16249 , \11452 , \11143 );
or \U$7431 ( \16250 , \10859 , \11038 );
nand \U$7432 ( \16251 , \16249 , \16250 );
or \U$7433 ( \16252 , \9055 , \10979 );
or \U$7434 ( \16253 , \9047 , \11019 );
nand \U$7435 ( \16254 , \16252 , \16253 );
nor \U$7436 ( \16255 , \16251 , \16254 );
or \U$7437 ( \16256 , \9068 , \11065 );
or \U$7438 ( \16257 , \11458 , \11068 );
nand \U$7439 ( \16258 , \16256 , \16257 );
or \U$7440 ( \16259 , \9073 , \10935 );
or \U$7441 ( \16260 , \9076 , \10963 );
nand \U$7442 ( \16261 , \16259 , \16260 );
nor \U$7443 ( \16262 , \16258 , \16261 );
not \U$7444 ( \16263 , \11327 );
and \U$7445 ( \16264 , \9093 , \16263 );
not \U$7446 ( \16265 , \11209 );
and \U$7447 ( \16266 , \9112 , \16265 );
nor \U$7448 ( \16267 , \16264 , \16266 );
not \U$7449 ( \16268 , \11182 );
and \U$7450 ( \16269 , \9081 , \16268 );
not \U$7451 ( \16270 , \11203 );
and \U$7452 ( \16271 , \9089 , \16270 );
nor \U$7453 ( \16272 , \16269 , \16271 );
nand \U$7454 ( \16273 , \16267 , \16272 );
not \U$7455 ( \16274 , \9086 );
and \U$7456 ( \16275 , \16274 , \11174 );
and \U$7457 ( \16276 , \11015 , \9057 );
nor \U$7458 ( \16277 , \16275 , \16276 );
not \U$7459 ( \16278 , \11473 );
and \U$7460 ( \16279 , \16278 , \16166 );
and \U$7461 ( \16280 , \11010 , \9049 );
nor \U$7462 ( \16281 , \16279 , \16280 );
nand \U$7463 ( \16282 , \16277 , \16281 );
nor \U$7464 ( \16283 , \16273 , \16282 );
nand \U$7465 ( \16284 , \16255 , \16262 , \16283 );
xnor \U$7466 ( \16285 , \16284 , \9119 );
nor \U$7467 ( \16286 , \16248 , \16285 );
or \U$7468 ( \16287 , \11270 , \11022 );
or \U$7469 ( \16288 , \10415 , \10973 );
nand \U$7470 ( \16289 , \16287 , \16288 );
or \U$7471 ( \16290 , \9270 , \11032 );
or \U$7472 ( \16291 , \9263 , \11019 );
nand \U$7473 ( \16292 , \16290 , \16291 );
nor \U$7474 ( \16293 , \16289 , \16292 );
or \U$7475 ( \16294 , \9282 , \11118 );
or \U$7476 ( \16295 , \11276 , \11068 );
nand \U$7477 ( \16296 , \16294 , \16295 );
or \U$7478 ( \16297 , \9287 , \10935 );
or \U$7479 ( \16298 , \9290 , \10963 );
nand \U$7480 ( \16299 , \16297 , \16298 );
nor \U$7481 ( \16300 , \16296 , \16299 );
not \U$7482 ( \16301 , \11199 );
and \U$7483 ( \16302 , \16301 , \9302 );
not \U$7484 ( \16303 , \10991 );
and \U$7485 ( \16304 , \9319 , \16303 );
nor \U$7486 ( \16305 , \16302 , \16304 );
not \U$7487 ( \16306 , \11126 );
and \U$7488 ( \16307 , \9295 , \16306 );
not \U$7489 ( \16308 , \11279 );
and \U$7490 ( \16309 , \9299 , \16308 );
nor \U$7491 ( \16310 , \16307 , \16309 );
nand \U$7492 ( \16311 , \16305 , \16310 );
not \U$7493 ( \16312 , \11298 );
and \U$7494 ( \16313 , \16312 , \11174 );
and \U$7495 ( \16314 , \11015 , \9272 );
nor \U$7496 ( \16315 , \16313 , \16314 );
not \U$7497 ( \16316 , \11293 );
and \U$7498 ( \16317 , \16316 , \16166 );
and \U$7499 ( \16318 , \11010 , \9265 );
nor \U$7500 ( \16319 , \16317 , \16318 );
nand \U$7501 ( \16320 , \16315 , \16319 );
nor \U$7502 ( \16321 , \16311 , \16320 );
nand \U$7503 ( \16322 , \16293 , \16300 , \16321 );
xnor \U$7504 ( \16323 , \16322 , \9327 );
or \U$7505 ( \16324 , \11230 , \11319 );
or \U$7506 ( \16325 , \10462 , \11038 );
nand \U$7507 ( \16326 , \16324 , \16325 );
or \U$7508 ( \16327 , \9402 , \11389 );
or \U$7509 ( \16328 , \9395 , \11019 );
nand \U$7510 ( \16329 , \16327 , \16328 );
nor \U$7511 ( \16330 , \16326 , \16329 );
or \U$7512 ( \16331 , \9415 , \10955 );
or \U$7513 ( \16332 , \10455 , \11068 );
nand \U$7514 ( \16333 , \16331 , \16332 );
or \U$7515 ( \16334 , \9419 , \10935 );
or \U$7516 ( \16335 , \9422 , \10963 );
nand \U$7517 ( \16336 , \16334 , \16335 );
nor \U$7518 ( \16337 , \16333 , \16336 );
not \U$7519 ( \16338 , \10982 );
and \U$7520 ( \16339 , \9435 , \16338 );
not \U$7521 ( \16340 , \11099 );
and \U$7522 ( \16341 , \9453 , \16340 );
nor \U$7523 ( \16342 , \16339 , \16341 );
not \U$7524 ( \16343 , \11126 );
and \U$7525 ( \16344 , \9427 , \16343 );
not \U$7526 ( \16345 , \11051 );
and \U$7527 ( \16346 , \9432 , \16345 );
nor \U$7528 ( \16347 , \16344 , \16346 );
nand \U$7529 ( \16348 , \16342 , \16347 );
not \U$7530 ( \16349 , \10464 );
and \U$7531 ( \16350 , \16349 , \11174 );
and \U$7532 ( \16351 , \11015 , \9404 );
nor \U$7533 ( \16352 , \16350 , \16351 );
not \U$7534 ( \16353 , \11250 );
and \U$7535 ( \16354 , \16353 , \16166 );
and \U$7536 ( \16355 , \11010 , \9397 );
nor \U$7537 ( \16356 , \16354 , \16355 );
nand \U$7538 ( \16357 , \16352 , \16356 );
nor \U$7539 ( \16358 , \16348 , \16357 );
nand \U$7540 ( \16359 , \16330 , \16337 , \16358 );
xnor \U$7541 ( \16360 , \16359 , \9460 );
nor \U$7542 ( \16361 , \16323 , \16360 );
and \U$7543 ( \16362 , \16211 , \16286 , \16361 );
not \U$7544 ( \16363 , \11023 );
or \U$7545 ( \16364 , \9851 , \16363 );
not \U$7546 ( \16365 , \11020 );
or \U$7547 ( \16366 , \11505 , \16365 );
not \U$7548 ( \16367 , \11126 );
and \U$7549 ( \16368 , \9842 , \16367 );
not \U$7550 ( \16369 , \10979 );
and \U$7551 ( \16370 , \9839 , \16369 );
nor \U$7552 ( \16371 , \16368 , \16370 );
nand \U$7553 ( \16372 , \16364 , \16366 , \16371 );
not \U$7554 ( \16373 , \16372 );
not \U$7555 ( \16374 , \11102 );
and \U$7556 ( \16375 , \9826 , \16374 );
not \U$7557 ( \16376 , \11209 );
and \U$7558 ( \16377 , \9822 , \16376 );
nor \U$7559 ( \16378 , \16375 , \16377 );
not \U$7560 ( \16379 , \11281 );
and \U$7561 ( \16380 , \9830 , \16379 );
not \U$7562 ( \16381 , \11160 );
and \U$7563 ( \16382 , \9833 , \16381 );
nor \U$7564 ( \16383 , \16380 , \16382 );
and \U$7565 ( \16384 , \16373 , \16378 , \16383 );
not \U$7566 ( \16385 , \11010 );
or \U$7567 ( \16386 , \9817 , \16385 );
not \U$7568 ( \16387 , \11015 );
or \U$7569 ( \16388 , \9806 , \16387 );
not \U$7570 ( \16389 , \10973 );
and \U$7571 ( \16390 , \9813 , \16389 );
not \U$7572 ( \16391 , \10944 );
and \U$7573 ( \16392 , \9808 , \16391 );
nor \U$7574 ( \16393 , \16390 , \16392 );
nand \U$7575 ( \16394 , \16386 , \16388 , \16393 );
not \U$7576 ( \16395 , \9791 );
and \U$7577 ( \16396 , \16395 , \11367 );
and \U$7578 ( \16397 , \10962 , \9794 );
nor \U$7579 ( \16398 , \16396 , \16397 );
not \U$7580 ( \16399 , \9798 );
and \U$7581 ( \16400 , \16399 , \11374 );
and \U$7582 ( \16401 , \10954 , \9801 );
nor \U$7583 ( \16402 , \16400 , \16401 );
nand \U$7584 ( \16403 , \16398 , \16402 );
nor \U$7585 ( \16404 , \16394 , \16403 );
nand \U$7586 ( \16405 , \16384 , \16404 );
xnor \U$7587 ( \16406 , RIb7a5bf8_260, \16405 );
or \U$7588 ( \16407 , \9878 , \11081 );
or \U$7589 ( \16408 , \9884 , \11038 );
nand \U$7590 ( \16409 , \16407 , \16408 );
or \U$7591 ( \16410 , \9887 , \11009 );
or \U$7592 ( \16411 , \9875 , \11014 );
nand \U$7593 ( \16412 , \16410 , \16411 );
nor \U$7594 ( \16413 , \16409 , \16412 );
or \U$7595 ( \16414 , \12178 , \10955 );
or \U$7596 ( \16415 , \9868 , \10970 );
nand \U$7597 ( \16416 , \16414 , \16415 );
or \U$7598 ( \16417 , \9860 , \11114 );
or \U$7599 ( \16418 , \12183 , \16046 );
nand \U$7600 ( \16419 , \16417 , \16418 );
nor \U$7601 ( \16420 , \16416 , \16419 );
nand \U$7602 ( \16421 , \16413 , \16420 );
not \U$7603 ( \16422 , \16421 );
or \U$7604 ( \16423 , \9911 , \11032 );
or \U$7605 ( \16424 , \9914 , \11000 );
nand \U$7606 ( \16425 , \16423 , \16424 );
or \U$7607 ( \16426 , \9921 , \11022 );
or \U$7608 ( \16427 , \11718 , \11019 );
nand \U$7609 ( \16428 , \16426 , \16427 );
nor \U$7610 ( \16429 , \16425 , \16428 );
or \U$7611 ( \16430 , \9895 , \11099 );
or \U$7612 ( \16431 , \9898 , \10987 );
nand \U$7613 ( \16432 , \16430 , \16431 );
or \U$7614 ( \16433 , \9906 , \11105 );
or \U$7615 ( \16434 , \11711 , \11053 );
nand \U$7616 ( \16435 , \16433 , \16434 );
nor \U$7617 ( \16436 , \16432 , \16435 );
and \U$7618 ( \16437 , \16422 , \16429 , \16436 );
xnor \U$7619 ( \16438 , \16437 , \9927 );
or \U$7620 ( \16439 , \9933 , \11131 );
or \U$7621 ( \16440 , \9937 , \10973 );
nand \U$7622 ( \16441 , \16439 , \16440 );
or \U$7623 ( \16442 , \9940 , \11009 );
or \U$7624 ( \16443 , \9930 , \11014 );
nand \U$7625 ( \16444 , \16442 , \16443 );
nor \U$7626 ( \16445 , \16441 , \16444 );
or \U$7627 ( \16446 , \9948 , \11118 );
or \U$7628 ( \16447 , \13143 , \10970 );
nand \U$7629 ( \16448 , \16446 , \16447 );
or \U$7630 ( \16449 , \9952 , \11114 );
or \U$7631 ( \16450 , \9955 , \16046 );
nand \U$7632 ( \16451 , \16449 , \16450 );
nor \U$7633 ( \16452 , \16448 , \16451 );
nand \U$7634 ( \16453 , \9984 , \11023 );
nand \U$7635 ( \16454 , \9982 , \11020 );
not \U$7636 ( \16455 , \11000 );
and \U$7637 ( \16456 , \9975 , \16455 );
not \U$7638 ( \16457 , \11389 );
and \U$7639 ( \16458 , \9977 , \16457 );
nor \U$7640 ( \16459 , \16456 , \16458 );
nand \U$7641 ( \16460 , \16453 , \16454 , \16459 );
not \U$7642 ( \16461 , \16460 );
not \U$7643 ( \16462 , \10987 );
and \U$7644 ( \16463 , \9965 , \16462 );
not \U$7645 ( \16464 , \11099 );
and \U$7646 ( \16465 , \9968 , \16464 );
nor \U$7647 ( \16466 , \16463 , \16465 );
not \U$7648 ( \16467 , \11281 );
and \U$7649 ( \16468 , \10709 , \16467 );
not \U$7650 ( \16469 , \11160 );
and \U$7651 ( \16470 , \9959 , \16469 );
nor \U$7652 ( \16471 , \16468 , \16470 );
and \U$7653 ( \16472 , \16461 , \16466 , \16471 );
nand \U$7654 ( \16473 , \16445 , \16452 , \16472 );
xnor \U$7655 ( \16474 , \16473 , \9990 );
nand \U$7656 ( \16475 , \10049 , \11023 );
nand \U$7657 ( \16476 , \10047 , \11020 );
not \U$7658 ( \16477 , \11075 );
and \U$7659 ( \16478 , \16477 , \10041 );
not \U$7660 ( \16479 , \11032 );
and \U$7661 ( \16480 , \10043 , \16479 );
nor \U$7662 ( \16481 , \16478 , \16480 );
nand \U$7663 ( \16482 , \16475 , \16476 , \16481 );
not \U$7664 ( \16483 , \16482 );
not \U$7665 ( \16484 , \11047 );
and \U$7666 ( \16485 , \10030 , \16484 );
not \U$7667 ( \16486 , \10991 );
and \U$7668 ( \16487 , \10035 , \16486 );
nor \U$7669 ( \16488 , \16485 , \16487 );
not \U$7670 ( \16489 , \11327 );
and \U$7671 ( \16490 , \10027 , \16489 );
not \U$7672 ( \16491 , \10996 );
and \U$7673 ( \16492 , \10025 , \16491 );
nor \U$7674 ( \16493 , \16490 , \16492 );
and \U$7675 ( \16494 , \16483 , \16488 , \16493 );
not \U$7676 ( \16495 , \11010 );
or \U$7677 ( \16496 , \10021 , \16495 );
not \U$7678 ( \16497 , \11015 );
or \U$7679 ( \16498 , \10010 , \16497 );
not \U$7680 ( \16499 , \11038 );
and \U$7681 ( \16500 , \10017 , \16499 );
not \U$7682 ( \16501 , \10944 );
and \U$7683 ( \16502 , \16501 , \10012 );
nor \U$7684 ( \16503 , \16500 , \16502 );
nand \U$7685 ( \16504 , \16496 , \16498 , \16503 );
not \U$7686 ( \16505 , \10002 );
and \U$7687 ( \16506 , \16505 , \11367 );
and \U$7688 ( \16507 , \10962 , \10004 );
nor \U$7689 ( \16508 , \16506 , \16507 );
not \U$7690 ( \16509 , \11666 );
and \U$7691 ( \16510 , \16509 , \11374 );
and \U$7692 ( \16511 , \10954 , \9996 );
nor \U$7693 ( \16512 , \16510 , \16511 );
nand \U$7694 ( \16513 , \16508 , \16512 );
nor \U$7695 ( \16514 , \16504 , \16513 );
nand \U$7696 ( \16515 , \16494 , \16514 );
xnor \U$7697 ( \16516 , \16515 , \10055 );
nor \U$7698 ( \16517 , \16474 , \16516 );
nand \U$7699 ( \16518 , \16406 , \16438 , \16517 );
not \U$7700 ( \16519 , \16518 );
or \U$7701 ( \16520 , \9722 , \11389 );
or \U$7702 ( \16521 , \9725 , \11182 );
nand \U$7703 ( \16522 , \16520 , \16521 );
or \U$7704 ( \16523 , \9732 , \11319 );
or \U$7705 ( \16524 , \13305 , \11019 );
nand \U$7706 ( \16525 , \16523 , \16524 );
nor \U$7707 ( \16526 , \16522 , \16525 );
or \U$7708 ( \16527 , \9740 , \11065 );
or \U$7709 ( \16528 , \11876 , \10970 );
nand \U$7710 ( \16529 , \16527 , \16528 );
or \U$7711 ( \16530 , \9745 , \11114 );
or \U$7712 ( \16531 , \9748 , \16046 );
nand \U$7713 ( \16532 , \16530 , \16531 );
nor \U$7714 ( \16533 , \16529 , \16532 );
not \U$7715 ( \16534 , \11053 );
and \U$7716 ( \16535 , \9755 , \16534 );
not \U$7717 ( \16536 , \11203 );
and \U$7718 ( \16537 , \9752 , \16536 );
nor \U$7719 ( \16538 , \16535 , \16537 );
not \U$7720 ( \16539 , \10987 );
and \U$7721 ( \16540 , \9759 , \16539 );
not \U$7722 ( \16541 , \11209 );
and \U$7723 ( \16542 , \9763 , \16541 );
nor \U$7724 ( \16543 , \16540 , \16542 );
nand \U$7725 ( \16544 , \16538 , \16543 );
not \U$7726 ( \16545 , \11010 );
or \U$7727 ( \16546 , \11186 , \16545 );
not \U$7728 ( \16547 , \11015 );
or \U$7729 ( \16548 , \10178 , \16547 );
not \U$7730 ( \16549 , \11038 );
and \U$7731 ( \16550 , \9779 , \16549 );
not \U$7732 ( \16551 , \10944 );
and \U$7733 ( \16552 , \9769 , \16551 );
nor \U$7734 ( \16553 , \16550 , \16552 );
nand \U$7735 ( \16554 , \16546 , \16548 , \16553 );
nor \U$7736 ( \16555 , \16544 , \16554 );
nand \U$7737 ( \16556 , \16526 , \16533 , \16555 );
xnor \U$7738 ( \16557 , \16556 , \9786 );
or \U$7739 ( \16558 , \9658 , \10979 );
or \U$7740 ( \16559 , \9661 , \11000 );
nand \U$7741 ( \16560 , \16558 , \16559 );
or \U$7742 ( \16561 , \9668 , \11143 );
or \U$7743 ( \16562 , \13344 , \11019 );
nand \U$7744 ( \16563 , \16561 , \16562 );
nor \U$7745 ( \16564 , \16560 , \16563 );
or \U$7746 ( \16565 , \9676 , \11118 );
or \U$7747 ( \16566 , \11923 , \10970 );
nand \U$7748 ( \16567 , \16565 , \16566 );
or \U$7749 ( \16568 , \9680 , \11114 );
or \U$7750 ( \16569 , \9683 , \16046 );
nand \U$7751 ( \16570 , \16568 , \16569 );
nor \U$7752 ( \16571 , \16567 , \16570 );
not \U$7753 ( \16572 , \11327 );
and \U$7754 ( \16573 , \9690 , \16572 );
not \U$7755 ( \16574 , \11279 );
and \U$7756 ( \16575 , \9687 , \16574 );
nor \U$7757 ( \16576 , \16573 , \16575 );
not \U$7758 ( \16577 , \11047 );
and \U$7759 ( \16578 , \9692 , \16577 );
not \U$7760 ( \16579 , \10991 );
and \U$7761 ( \16580 , \9695 , \16579 );
nor \U$7762 ( \16581 , \16578 , \16580 );
nand \U$7763 ( \16582 , \16576 , \16581 );
not \U$7764 ( \16583 , \11010 );
or \U$7765 ( \16584 , \11145 , \16583 );
not \U$7766 ( \16585 , \11015 );
or \U$7767 ( \16586 , \11138 , \16585 );
not \U$7768 ( \16587 , \10973 );
and \U$7769 ( \16588 , \9713 , \16587 );
not \U$7770 ( \16589 , \11131 );
and \U$7771 ( \16590 , \9701 , \16589 );
nor \U$7772 ( \16591 , \16588 , \16590 );
nand \U$7773 ( \16592 , \16584 , \16586 , \16591 );
nor \U$7774 ( \16593 , \16582 , \16592 );
nand \U$7775 ( \16594 , \16564 , \16571 , \16593 );
xnor \U$7776 ( \16595 , \16594 , \9719 );
nor \U$7777 ( \16596 , \16557 , \16595 );
or \U$7778 ( \16597 , \11036 , \11022 );
or \U$7779 ( \16598 , \10370 , \10973 );
nand \U$7780 ( \16599 , \16597 , \16598 );
or \U$7781 ( \16600 , \8977 , \11032 );
or \U$7782 ( \16601 , \8967 , \11019 );
nand \U$7783 ( \16602 , \16600 , \16601 );
nor \U$7784 ( \16603 , \16599 , \16602 );
or \U$7785 ( \16604 , \8991 , \10955 );
or \U$7786 ( \16605 , \11046 , \10970 );
nand \U$7787 ( \16606 , \16604 , \16605 );
or \U$7788 ( \16607 , \8997 , \11114 );
or \U$7789 ( \16608 , \9000 , \16046 );
nand \U$7790 ( \16609 , \16607 , \16608 );
nor \U$7791 ( \16610 , \16606 , \16609 );
not \U$7792 ( \16611 , \11053 );
and \U$7793 ( \16612 , \9014 , \16611 );
not \U$7794 ( \16613 , \10991 );
and \U$7795 ( \16614 , \9034 , \16613 );
nor \U$7796 ( \16615 , \16612 , \16614 );
not \U$7797 ( \16616 , \11182 );
and \U$7798 ( \16617 , \9006 , \16616 );
not \U$7799 ( \16618 , \11203 );
and \U$7800 ( \16619 , \9011 , \16618 );
nor \U$7801 ( \16620 , \16617 , \16619 );
nand \U$7802 ( \16621 , \16615 , \16620 );
not \U$7803 ( \16622 , \11073 );
and \U$7804 ( \16623 , \16622 , \11174 );
and \U$7805 ( \16624 , \11015 , \8979 );
nor \U$7806 ( \16625 , \16623 , \16624 );
not \U$7807 ( \16626 , \11067 );
and \U$7808 ( \16627 , \16626 , \16166 );
and \U$7809 ( \16628 , \11010 , \8970 );
nor \U$7810 ( \16629 , \16627 , \16628 );
nand \U$7811 ( \16630 , \16625 , \16629 );
nor \U$7812 ( \16631 , \16621 , \16630 );
nand \U$7813 ( \16632 , \16603 , \16610 , \16631 );
xnor \U$7814 ( \16633 , \16632 , \9044 );
or \U$7815 ( \16634 , \11093 , \11319 );
or \U$7816 ( \16635 , \10323 , \11038 );
nand \U$7817 ( \16636 , \16634 , \16635 );
or \U$7818 ( \16637 , \9205 , \11389 );
or \U$7819 ( \16638 , \9197 , \11019 );
nand \U$7820 ( \16639 , \16637 , \16638 );
nor \U$7821 ( \16640 , \16636 , \16639 );
or \U$7822 ( \16641 , \11098 , \11065 );
or \U$7823 ( \16642 , \11101 , \10970 );
nand \U$7824 ( \16643 , \16641 , \16642 );
or \U$7825 ( \16644 , \9217 , \11114 );
or \U$7826 ( \16645 , \9220 , \16046 );
nand \U$7827 ( \16646 , \16644 , \16645 );
nor \U$7828 ( \16647 , \16643 , \16646 );
not \U$7829 ( \16648 , \11281 );
and \U$7830 ( \16649 , \9233 , \16648 );
not \U$7831 ( \16650 , \11044 );
and \U$7832 ( \16651 , \9251 , \16650 );
nor \U$7833 ( \16652 , \16649 , \16651 );
not \U$7834 ( \16653 , \11126 );
and \U$7835 ( \16654 , \9225 , \16653 );
not \U$7836 ( \16655 , \11279 );
and \U$7837 ( \16656 , \9230 , \16655 );
nor \U$7838 ( \16657 , \16654 , \16656 );
nand \U$7839 ( \16658 , \16652 , \16657 );
not \U$7840 ( \16659 , \11125 );
and \U$7841 ( \16660 , \16659 , \11174 );
and \U$7842 ( \16661 , \11015 , \9200 );
nor \U$7843 ( \16662 , \16660 , \16661 );
not \U$7844 ( \16663 , \11120 );
and \U$7845 ( \16664 , \16663 , \16166 );
and \U$7846 ( \16665 , \11010 , \9193 );
nor \U$7847 ( \16666 , \16664 , \16665 );
nand \U$7848 ( \16667 , \16662 , \16666 );
nor \U$7849 ( \16668 , \16658 , \16667 );
nand \U$7850 ( \16669 , \16640 , \16647 , \16668 );
xnor \U$7851 ( \16670 , \16669 , \9260 );
nor \U$7852 ( \16671 , \16633 , \16670 );
and \U$7853 ( \16672 , \16519 , \16596 , \16671 );
nand \U$7854 ( \16673 , \16071 , \16362 , \16672 );
not \U$7855 ( \16674 , \16673 );
not \U$7856 ( \16675 , \16674 );
or \U$7857 ( \16676 , \16034 , \16675 );
not \U$7858 ( \16677 , \16676 );
and \U$7859 ( \16678 , \16007 , \16677 );
not \U$7860 ( \16679 , \16034 );
not \U$7861 ( \16680 , \16674 );
or \U$7862 ( \16681 , \16679 , \16680 );
not \U$7863 ( \16682 , \16681 );
not \U$7864 ( \16683 , \13249 );
not \U$7865 ( \16684 , \16683 );
not \U$7866 ( \16685 , \13256 );
and \U$7867 ( \16686 , \16684 , \16685 );
not \U$7868 ( \16687 , \10065 );
and \U$7869 ( \16688 , \16687 , \13256 );
or \U$7870 ( \16689 , \16686 , \16688 );
not \U$7871 ( \16690 , \16689 );
or \U$7872 ( \16691 , \13255 , \16690 );
and \U$7873 ( \16692 , \16682 , \16691 );
nor \U$7874 ( \16693 , \16678 , \16692 );
nand \U$7875 ( \16694 , \16676 , \16681 );
not \U$7876 ( \16695 , \16694 );
not \U$7877 ( \16696 , \8876 );
not \U$7878 ( \16697 , \8837 );
and \U$7879 ( \16698 , \16696 , \16697 );
not \U$7880 ( \16699 , \8906 );
and \U$7881 ( \16700 , \16699 , \8837 );
or \U$7882 ( \16701 , \16698 , \16700 );
nand \U$7883 ( \16702 , \16701 , \8832 );
not \U$7884 ( \16703 , \16702 );
not \U$7885 ( \16704 , \16703 );
buf \U$7886 ( \16705 , \14685 );
buf \U$7887 ( \16706 , \12456 );
buf \U$7888 ( \16707 , \12458 );
not \U$7889 ( \16708 , \16707 );
not \U$7890 ( \16709 , \16708 );
or \U$7891 ( \16710 , \16706 , \16709 );
xnor \U$7892 ( \16711 , \16705 , \16710 );
buf \U$7893 ( \16712 , \16711 );
not \U$7894 ( \16713 , \16712 );
xnor \U$7895 ( \16714 , \16706 , \16709 );
buf \U$7896 ( \16715 , \16714 );
buf \U$7897 ( \16716 , \16708 );
buf \U$7898 ( \16717 , \8835 );
nor \U$7899 ( \16718 , \16715 , \16716 , \16717 );
and \U$7900 ( \16719 , \16713 , \16718 );
buf \U$7901 ( \16720 , RIea91330_6888);
or \U$7902 ( \16721 , \16705 , \16710 );
xor \U$7903 ( \16722 , \16720 , \16721 );
buf \U$7904 ( \16723 , \16722 );
not \U$7905 ( \16724 , \16723 );
or \U$7906 ( \16725 , \16719 , \16724 );
and \U$7907 ( \16726 , \16720 , \16721 );
buf \U$7908 ( \16727 , \16726 );
not \U$7909 ( \16728 , \16727 );
nand \U$7910 ( \16729 , \16725 , \16728 );
not \U$7911 ( \16730 , \16729 );
not \U$7912 ( \16731 , \9492 );
not \U$7913 ( \16732 , \16702 );
or \U$7914 ( \16733 , \13992 , \16732 );
not \U$7915 ( \16734 , \16733 );
not \U$7916 ( \16735 , \16734 );
or \U$7917 ( \16736 , \16735 , \13991 );
not \U$7918 ( \16737 , \16736 );
and \U$7919 ( \16738 , \16731 , \16737 );
and \U$7920 ( \16739 , \13992 , \16702 );
not \U$7921 ( \16740 , \16739 );
or \U$7922 ( \16741 , \10922 , \16740 );
not \U$7923 ( \16742 , \16741 );
not \U$7924 ( \16743 , \16742 );
or \U$7925 ( \16744 , \9498 , \16743 );
not \U$7926 ( \16745 , \16739 );
or \U$7927 ( \16746 , \16745 , \14008 );
or \U$7928 ( \16747 , \9500 , \16746 );
nand \U$7929 ( \16748 , \16744 , \16747 );
not \U$7930 ( \16749 , \16734 );
or \U$7931 ( \16750 , \10917 , \16749 );
not \U$7932 ( \16751 , \16750 );
and \U$7933 ( \16752 , \10062 , \16751 );
nor \U$7934 ( \16753 , \16738 , \16748 , \16752 );
not \U$7935 ( \16754 , \16703 );
or \U$7936 ( \16755 , \13992 , \16754 );
not \U$7937 ( \16756 , \16755 );
not \U$7938 ( \16757 , \16756 );
or \U$7939 ( \16758 , \10922 , \16757 );
or \U$7940 ( \16759 , \9504 , \16758 );
not \U$7941 ( \16760 , \16739 );
or \U$7942 ( \16761 , \10917 , \16760 );
not \U$7943 ( \16762 , \16761 );
not \U$7944 ( \16763 , \16762 );
or \U$7945 ( \16764 , \9506 , \16763 );
nand \U$7946 ( \16765 , \16759 , \16764 );
and \U$7947 ( \16766 , \16703 , \13992 );
not \U$7948 ( \16767 , \16766 );
or \U$7949 ( \16768 , \13991 , \16767 );
not \U$7950 ( \16769 , \16768 );
not \U$7951 ( \16770 , \16769 );
or \U$7952 ( \16771 , \9509 , \16770 );
not \U$7953 ( \16772 , \16766 );
or \U$7954 ( \16773 , \14008 , \16772 );
not \U$7955 ( \16774 , \16773 );
not \U$7956 ( \16775 , \16774 );
or \U$7957 ( \16776 , \9511 , \16775 );
nand \U$7958 ( \16777 , \16771 , \16776 );
nor \U$7959 ( \16778 , \16765 , \16777 );
not \U$7960 ( \16779 , \16766 );
or \U$7961 ( \16780 , \10922 , \16779 );
not \U$7962 ( \16781 , \16780 );
not \U$7963 ( \16782 , \16781 );
or \U$7964 ( \16783 , \9467 , \16782 );
not \U$7965 ( \16784 , \16766 );
or \U$7966 ( \16785 , \10917 , \16784 );
not \U$7967 ( \16786 , \16785 );
not \U$7968 ( \16787 , \16786 );
or \U$7969 ( \16788 , \9463 , \16787 );
not \U$7970 ( \16789 , \9471 );
not \U$7971 ( \16790 , \16756 );
or \U$7972 ( \16791 , \13991 , \16790 );
not \U$7973 ( \16792 , \16791 );
and \U$7974 ( \16793 , \16789 , \16792 );
not \U$7975 ( \16794 , \16756 );
or \U$7976 ( \16795 , \10917 , \16794 );
not \U$7977 ( \16796 , \16795 );
and \U$7978 ( \16797 , \16796 , \9476 );
nor \U$7979 ( \16798 , \16793 , \16797 );
nand \U$7980 ( \16799 , \16783 , \16788 , \16798 );
not \U$7981 ( \16800 , \16734 );
or \U$7982 ( \16801 , \10922 , \16800 );
not \U$7983 ( \16802 , \16801 );
not \U$7984 ( \16803 , \16802 );
or \U$7985 ( \16804 , \9485 , \16803 );
not \U$7986 ( \16805 , \16734 );
or \U$7987 ( \16806 , \14008 , \16805 );
not \U$7988 ( \16807 , \16806 );
not \U$7989 ( \16808 , \16807 );
or \U$7990 ( \16809 , \9487 , \16808 );
not \U$7991 ( \16810 , \9482 );
not \U$7992 ( \16811 , \16756 );
or \U$7993 ( \16812 , \14008 , \16811 );
not \U$7994 ( \16813 , \16812 );
and \U$7995 ( \16814 , \16810 , \16813 );
not \U$7996 ( \16815 , \16739 );
or \U$7997 ( \16816 , \13991 , \16815 );
not \U$7998 ( \16817 , \16816 );
not \U$7999 ( \16818 , \16817 );
not \U$8000 ( \16819 , \16818 );
and \U$8001 ( \16820 , \10152 , \16819 );
nor \U$8002 ( \16821 , \16814 , \16820 );
nand \U$8003 ( \16822 , \16804 , \16809 , \16821 );
nor \U$8004 ( \16823 , \16799 , \16822 );
nand \U$8005 ( \16824 , \16753 , \16778 , \16823 );
not \U$8006 ( \16825 , \16824 );
or \U$8007 ( \16826 , \9398 , \16812 );
or \U$8008 ( \16827 , \10462 , \16818 );
nand \U$8009 ( \16828 , \16826 , \16827 );
not \U$8010 ( \16829 , \16828 );
not \U$8011 ( \16830 , \16758 );
not \U$8012 ( \16831 , \16830 );
or \U$8013 ( \16832 , \9405 , \16831 );
not \U$8014 ( \16833 , \16796 );
or \U$8015 ( \16834 , \10464 , \16833 );
and \U$8016 ( \16835 , \16829 , \16832 , \16834 );
not \U$8017 ( \16836 , \16746 );
and \U$8018 ( \16837 , \16836 , \9435 );
not \U$8019 ( \16838 , \16762 );
or \U$8020 ( \16839 , \11250 , \16838 );
not \U$8021 ( \16840 , \16742 );
or \U$8022 ( \16841 , \11248 , \16840 );
nand \U$8023 ( \16842 , \16839 , \16841 );
not \U$8024 ( \16843 , \16734 );
or \U$8025 ( \16844 , \13991 , \16843 );
not \U$8026 ( \16845 , \16844 );
and \U$8027 ( \16846 , \9432 , \16845 );
nor \U$8028 ( \16847 , \16837 , \16842 , \16846 );
not \U$8029 ( \16848 , \16781 );
or \U$8030 ( \16849 , \9415 , \16848 );
not \U$8031 ( \16850 , \16786 );
or \U$8032 ( \16851 , \10455 , \16850 );
and \U$8033 ( \16852 , \16774 , \9421 );
and \U$8034 ( \16853 , \16792 , \9418 );
nor \U$8035 ( \16854 , \16852 , \16853 );
nand \U$8036 ( \16855 , \16849 , \16851 , \16854 );
not \U$8037 ( \16856 , \16750 );
not \U$8038 ( \16857 , \16856 );
or \U$8039 ( \16858 , \11259 , \16857 );
not \U$8040 ( \16859 , \16801 );
not \U$8041 ( \16860 , \16859 );
or \U$8042 ( \16861 , \9402 , \16860 );
not \U$8043 ( \16862 , \9395 );
and \U$8044 ( \16863 , \16862 , \16807 );
not \U$8045 ( \16864 , \16768 );
and \U$8046 ( \16865 , \16864 , \9440 );
nor \U$8047 ( \16866 , \16863 , \16865 );
nand \U$8048 ( \16867 , \16858 , \16861 , \16866 );
nor \U$8049 ( \16868 , \16855 , \16867 );
nand \U$8050 ( \16869 , \16835 , \16847 , \16868 );
xnor \U$8051 ( \16870 , RIb7b9590_247, \16869 );
or \U$8052 ( \16871 , \9266 , \16812 );
or \U$8053 ( \16872 , \10415 , \16818 );
nand \U$8054 ( \16873 , \16871 , \16872 );
not \U$8055 ( \16874 , \16873 );
not \U$8056 ( \16875 , \16830 );
or \U$8057 ( \16876 , \9273 , \16875 );
not \U$8058 ( \16877 , \16795 );
not \U$8059 ( \16878 , \16877 );
or \U$8060 ( \16879 , \11298 , \16878 );
and \U$8061 ( \16880 , \16874 , \16876 , \16879 );
not \U$8062 ( \16881 , \16739 );
or \U$8063 ( \16882 , \14008 , \16881 );
not \U$8064 ( \16883 , \16882 );
and \U$8065 ( \16884 , \16883 , \9302 );
not \U$8066 ( \16885 , \16762 );
or \U$8067 ( \16886 , \11293 , \16885 );
or \U$8068 ( \16887 , \11291 , \16743 );
nand \U$8069 ( \16888 , \16886 , \16887 );
not \U$8070 ( \16889 , \16736 );
and \U$8071 ( \16890 , \9299 , \16889 );
nor \U$8072 ( \16891 , \16884 , \16888 , \16890 );
not \U$8073 ( \16892 , \16781 );
or \U$8074 ( \16893 , \9282 , \16892 );
not \U$8075 ( \16894 , \16786 );
or \U$8076 ( \16895 , \11276 , \16894 );
not \U$8077 ( \16896 , \16773 );
and \U$8078 ( \16897 , \16896 , \9289 );
not \U$8079 ( \16898 , \16791 );
and \U$8080 ( \16899 , \16898 , \9286 );
nor \U$8081 ( \16900 , \16897 , \16899 );
nand \U$8082 ( \16901 , \16893 , \16895 , \16900 );
not \U$8083 ( \16902 , \16856 );
or \U$8084 ( \16903 , \11303 , \16902 );
not \U$8085 ( \16904 , \16859 );
or \U$8086 ( \16905 , \9270 , \16904 );
not \U$8087 ( \16906 , \9263 );
and \U$8088 ( \16907 , \16906 , \16807 );
and \U$8089 ( \16908 , \16864 , \9307 );
nor \U$8090 ( \16909 , \16907 , \16908 );
nand \U$8091 ( \16910 , \16903 , \16905 , \16909 );
nor \U$8092 ( \16911 , \16901 , \16910 );
nand \U$8093 ( \16912 , \16880 , \16891 , \16911 );
xnor \U$8094 ( \16913 , RIb7b9428_250, \16912 );
or \U$8095 ( \16914 , \9335 , \16812 );
or \U$8096 ( \16915 , \10553 , \16818 );
nand \U$8097 ( \16916 , \16914 , \16915 );
not \U$8098 ( \16917 , \16916 );
not \U$8099 ( \16918 , \16758 );
not \U$8100 ( \16919 , \16918 );
or \U$8101 ( \16920 , \9342 , \16919 );
not \U$8102 ( \16921 , \16877 );
or \U$8103 ( \16922 , \11357 , \16921 );
and \U$8104 ( \16923 , \16917 , \16920 , \16922 );
not \U$8105 ( \16924 , \16882 );
and \U$8106 ( \16925 , \16924 , \9369 );
not \U$8107 ( \16926 , \16762 );
or \U$8108 ( \16927 , \12874 , \16926 );
or \U$8109 ( \16928 , \11371 , \16840 );
nand \U$8110 ( \16929 , \16927 , \16928 );
not \U$8111 ( \16930 , \16844 );
and \U$8112 ( \16931 , \9366 , \16930 );
nor \U$8113 ( \16932 , \16925 , \16929 , \16931 );
not \U$8114 ( \16933 , \16781 );
or \U$8115 ( \16934 , \12139 , \16933 );
not \U$8116 ( \16935 , \16786 );
or \U$8117 ( \16936 , \12141 , \16935 );
and \U$8118 ( \16937 , \16896 , \9356 );
and \U$8119 ( \16938 , \16898 , \9353 );
nor \U$8120 ( \16939 , \16937 , \16938 );
nand \U$8121 ( \16940 , \16934 , \16936 , \16939 );
not \U$8122 ( \16941 , \16856 );
or \U$8123 ( \16942 , \11352 , \16941 );
not \U$8124 ( \16943 , \16859 );
or \U$8125 ( \16944 , \9339 , \16943 );
not \U$8126 ( \16945 , \9332 );
and \U$8127 ( \16946 , \16945 , \16807 );
and \U$8128 ( \16947 , \16864 , \9374 );
nor \U$8129 ( \16948 , \16946 , \16947 );
nand \U$8130 ( \16949 , \16942 , \16944 , \16948 );
nor \U$8131 ( \16950 , \16940 , \16949 );
nand \U$8132 ( \16951 , \16923 , \16932 , \16950 );
xnor \U$8133 ( \16952 , \16951 , \9392 );
or \U$8134 ( \16953 , \9125 , \16812 );
not \U$8135 ( \16954 , \16817 );
or \U$8136 ( \16955 , \10901 , \16954 );
nand \U$8137 ( \16956 , \16953 , \16955 );
not \U$8138 ( \16957 , \16956 );
not \U$8139 ( \16958 , \16918 );
or \U$8140 ( \16959 , \9133 , \16958 );
not \U$8141 ( \16960 , \16877 );
or \U$8142 ( \16961 , \11436 , \16960 );
and \U$8143 ( \16962 , \16957 , \16959 , \16961 );
not \U$8144 ( \16963 , \16746 );
and \U$8145 ( \16964 , \16963 , \9163 );
not \U$8146 ( \16965 , \16762 );
or \U$8147 ( \16966 , \11431 , \16965 );
or \U$8148 ( \16967 , \11429 , \16743 );
nand \U$8149 ( \16968 , \16966 , \16967 );
not \U$8150 ( \16969 , \16734 );
or \U$8151 ( \16970 , \13991 , \16969 );
not \U$8152 ( \16971 , \16970 );
and \U$8153 ( \16972 , \9159 , \16971 );
nor \U$8154 ( \16973 , \16964 , \16968 , \16972 );
not \U$8155 ( \16974 , \16781 );
or \U$8156 ( \16975 , \9143 , \16974 );
not \U$8157 ( \16976 , \16786 );
or \U$8158 ( \16977 , \11416 , \16976 );
and \U$8159 ( \16978 , \16774 , \9150 );
and \U$8160 ( \16979 , \16792 , \9147 );
nor \U$8161 ( \16980 , \16978 , \16979 );
nand \U$8162 ( \16981 , \16975 , \16977 , \16980 );
not \U$8163 ( \16982 , \16856 );
or \U$8164 ( \16983 , \11441 , \16982 );
not \U$8165 ( \16984 , \16859 );
or \U$8166 ( \16985 , \9130 , \16984 );
not \U$8167 ( \16986 , \9122 );
not \U$8168 ( \16987 , \16806 );
and \U$8169 ( \16988 , \16986 , \16987 );
and \U$8170 ( \16989 , \16864 , \9168 );
nor \U$8171 ( \16990 , \16988 , \16989 );
nand \U$8172 ( \16991 , \16983 , \16985 , \16990 );
nor \U$8173 ( \16992 , \16981 , \16991 );
nand \U$8174 ( \16993 , \16962 , \16973 , \16992 );
xnor \U$8175 ( \16994 , \16993 , \9188 );
nor \U$8176 ( \16995 , \16952 , \16994 );
nand \U$8177 ( \16996 , \16870 , \16913 , \16995 );
not \U$8178 ( \16997 , \16996 );
or \U$8179 ( \16998 , \11088 , \16812 );
or \U$8180 ( \16999 , \10323 , \16818 );
nand \U$8181 ( \17000 , \16998 , \16999 );
not \U$8182 ( \17001 , \17000 );
not \U$8183 ( \17002 , \16918 );
or \U$8184 ( \17003 , \11954 , \17002 );
not \U$8185 ( \17004 , \16796 );
or \U$8186 ( \17005 , \11125 , \17004 );
and \U$8187 ( \17006 , \17001 , \17003 , \17005 );
not \U$8188 ( \17007 , \16882 );
and \U$8189 ( \17008 , \17007 , \9233 );
or \U$8190 ( \17009 , \11120 , \16926 );
or \U$8191 ( \17010 , \11117 , \16743 );
nand \U$8192 ( \17011 , \17009 , \17010 );
not \U$8193 ( \17012 , \16970 );
and \U$8194 ( \17013 , \9230 , \17012 );
nor \U$8195 ( \17014 , \17008 , \17011 , \17013 );
not \U$8196 ( \17015 , \16781 );
or \U$8197 ( \17016 , \11098 , \17015 );
not \U$8198 ( \17017 , \16786 );
or \U$8199 ( \17018 , \11101 , \17017 );
and \U$8200 ( \17019 , \16896 , \9219 );
and \U$8201 ( \17020 , \16898 , \9216 );
nor \U$8202 ( \17021 , \17019 , \17020 );
nand \U$8203 ( \17022 , \17016 , \17018 , \17021 );
not \U$8204 ( \17023 , \16856 );
or \U$8205 ( \17024 , \9226 , \17023 );
not \U$8206 ( \17025 , \16859 );
or \U$8207 ( \17026 , \9205 , \17025 );
not \U$8208 ( \17027 , \9197 );
and \U$8209 ( \17028 , \17027 , \16807 );
and \U$8210 ( \17029 , \16864 , \9239 );
nor \U$8211 ( \17030 , \17028 , \17029 );
nand \U$8212 ( \17031 , \17024 , \17026 , \17030 );
nor \U$8213 ( \17032 , \17022 , \17031 );
nand \U$8214 ( \17033 , \17006 , \17014 , \17032 );
xnor \U$8215 ( \17034 , \17033 , \9260 );
or \U$8216 ( \17035 , \8971 , \16812 );
not \U$8217 ( \17036 , \16817 );
or \U$8218 ( \17037 , \10370 , \17036 );
nand \U$8219 ( \17038 , \17035 , \17037 );
not \U$8220 ( \17039 , \17038 );
not \U$8221 ( \17040 , \16830 );
or \U$8222 ( \17041 , \8980 , \17040 );
not \U$8223 ( \17042 , \16796 );
or \U$8224 ( \17043 , \11073 , \17042 );
and \U$8225 ( \17044 , \17039 , \17041 , \17043 );
not \U$8226 ( \17045 , \16746 );
and \U$8227 ( \17046 , \17045 , \9014 );
or \U$8228 ( \17047 , \11067 , \16965 );
or \U$8229 ( \17048 , \11064 , \16840 );
nand \U$8230 ( \17049 , \17047 , \17048 );
not \U$8231 ( \17050 , \16736 );
and \U$8232 ( \17051 , \9011 , \17050 );
nor \U$8233 ( \17052 , \17046 , \17049 , \17051 );
not \U$8234 ( \17053 , \16781 );
or \U$8235 ( \17054 , \8991 , \17053 );
not \U$8236 ( \17055 , \16786 );
or \U$8237 ( \17056 , \11046 , \17055 );
and \U$8238 ( \17057 , \16896 , \8999 );
and \U$8239 ( \17058 , \16898 , \8996 );
nor \U$8240 ( \17059 , \17057 , \17058 );
nand \U$8241 ( \17060 , \17054 , \17056 , \17059 );
not \U$8242 ( \17061 , \16856 );
or \U$8243 ( \17062 , \11080 , \17061 );
not \U$8244 ( \17063 , \16859 );
or \U$8245 ( \17064 , \8977 , \17063 );
not \U$8246 ( \17065 , \8967 );
and \U$8247 ( \17066 , \17065 , \16807 );
and \U$8248 ( \17067 , \16864 , \9020 );
nor \U$8249 ( \17068 , \17066 , \17067 );
nand \U$8250 ( \17069 , \17062 , \17064 , \17068 );
nor \U$8251 ( \17070 , \17060 , \17069 );
nand \U$8252 ( \17071 , \17044 , \17052 , \17070 );
xnor \U$8253 ( \17072 , \17071 , \9044 );
nor \U$8254 ( \17073 , \17034 , \17072 );
or \U$8255 ( \17074 , \8844 , \16812 );
or \U$8256 ( \17075 , \10775 , \17036 );
nand \U$8257 ( \17076 , \17074 , \17075 );
not \U$8258 ( \17077 , \17076 );
not \U$8259 ( \17078 , \16918 );
or \U$8260 ( \17079 , \8861 , \17078 );
not \U$8261 ( \17080 , \16796 );
or \U$8262 ( \17081 , \11533 , \17080 );
and \U$8263 ( \17082 , \17077 , \17079 , \17081 );
not \U$8264 ( \17083 , \16882 );
and \U$8265 ( \17084 , \17083 , \8927 );
not \U$8266 ( \17085 , \16762 );
or \U$8267 ( \17086 , \11545 , \17085 );
or \U$8268 ( \17087 , \14573 , \16840 );
nand \U$8269 ( \17088 , \17086 , \17087 );
not \U$8270 ( \17089 , \16844 );
and \U$8271 ( \17090 , \8921 , \17089 );
nor \U$8272 ( \17091 , \17084 , \17088 , \17090 );
not \U$8273 ( \17092 , \16781 );
or \U$8274 ( \17093 , \8882 , \17092 );
not \U$8275 ( \17094 , \16786 );
or \U$8276 ( \17095 , \12351 , \17094 );
and \U$8277 ( \17096 , \16774 , \8896 );
and \U$8278 ( \17097 , \16792 , \8893 );
nor \U$8279 ( \17098 , \17096 , \17097 );
nand \U$8280 ( \17099 , \17093 , \17095 , \17098 );
not \U$8281 ( \17100 , \16856 );
or \U$8282 ( \17101 , \11528 , \17100 );
not \U$8283 ( \17102 , \16859 );
or \U$8284 ( \17103 , \8853 , \17102 );
not \U$8285 ( \17104 , \8828 );
and \U$8286 ( \17105 , \17104 , \16807 );
and \U$8287 ( \17106 , \16864 , \8934 );
nor \U$8288 ( \17107 , \17105 , \17106 );
nand \U$8289 ( \17108 , \17101 , \17103 , \17107 );
nor \U$8290 ( \17109 , \17099 , \17108 );
nand \U$8291 ( \17110 , \17082 , \17091 , \17109 );
xnor \U$8292 ( \17111 , \17110 , \8964 );
or \U$8293 ( \17112 , \9050 , \16812 );
or \U$8294 ( \17113 , \10859 , \16818 );
nand \U$8295 ( \17114 , \17112 , \17113 );
not \U$8296 ( \17115 , \17114 );
not \U$8297 ( \17116 , \16918 );
or \U$8298 ( \17117 , \9058 , \17116 );
not \U$8299 ( \17118 , \16877 );
or \U$8300 ( \17119 , \9086 , \17118 );
and \U$8301 ( \17120 , \17115 , \17117 , \17119 );
not \U$8302 ( \17121 , \16746 );
and \U$8303 ( \17122 , \17121 , \9093 );
not \U$8304 ( \17123 , \16739 );
or \U$8305 ( \17124 , \10917 , \17123 );
or \U$8306 ( \17125 , \11473 , \17124 );
or \U$8307 ( \17126 , \11471 , \16743 );
nand \U$8308 ( \17127 , \17125 , \17126 );
not \U$8309 ( \17128 , \16970 );
and \U$8310 ( \17129 , \9089 , \17128 );
nor \U$8311 ( \17130 , \17122 , \17127 , \17129 );
not \U$8312 ( \17131 , \16781 );
or \U$8313 ( \17132 , \9068 , \17131 );
not \U$8314 ( \17133 , \16786 );
or \U$8315 ( \17134 , \11458 , \17133 );
and \U$8316 ( \17135 , \16774 , \9075 );
and \U$8317 ( \17136 , \16792 , \9072 );
nor \U$8318 ( \17137 , \17135 , \17136 );
nand \U$8319 ( \17138 , \17132 , \17134 , \17137 );
not \U$8320 ( \17139 , \16856 );
or \U$8321 ( \17140 , \9082 , \17139 );
not \U$8322 ( \17141 , \16859 );
or \U$8323 ( \17142 , \9055 , \17141 );
not \U$8324 ( \17143 , \9047 );
and \U$8325 ( \17144 , \17143 , \16987 );
and \U$8326 ( \17145 , \16864 , \9098 );
nor \U$8327 ( \17146 , \17144 , \17145 );
nand \U$8328 ( \17147 , \17140 , \17142 , \17146 );
nor \U$8329 ( \17148 , \17138 , \17147 );
nand \U$8330 ( \17149 , \17120 , \17130 , \17148 );
xnor \U$8331 ( \17150 , \17149 , \9119 );
nor \U$8332 ( \17151 , \17111 , \17150 );
and \U$8333 ( \17152 , \16997 , \17073 , \17151 );
or \U$8334 ( \17153 , \9722 , \16801 );
or \U$8335 ( \17154 , \9725 , \16750 );
nand \U$8336 ( \17155 , \17153 , \17154 );
or \U$8337 ( \17156 , \13305 , \16806 );
not \U$8338 ( \17157 , \16864 );
or \U$8339 ( \17158 , \9732 , \17157 );
nand \U$8340 ( \17159 , \17156 , \17158 );
nor \U$8341 ( \17160 , \17155 , \17159 );
not \U$8342 ( \17161 , \16781 );
or \U$8343 ( \17162 , \9740 , \17161 );
not \U$8344 ( \17163 , \16786 );
or \U$8345 ( \17164 , \11876 , \17163 );
nand \U$8346 ( \17165 , \17162 , \17164 );
not \U$8347 ( \17166 , \16792 );
or \U$8348 ( \17167 , \9745 , \17166 );
not \U$8349 ( \17168 , \16774 );
or \U$8350 ( \17169 , \9748 , \17168 );
nand \U$8351 ( \17170 , \17167 , \17169 );
nor \U$8352 ( \17171 , \17165 , \17170 );
not \U$8353 ( \17172 , \16737 );
or \U$8354 ( \17173 , \11193 , \17172 );
not \U$8355 ( \17174 , \16746 );
not \U$8356 ( \17175 , \17174 );
or \U$8357 ( \17176 , \11195 , \17175 );
not \U$8358 ( \17177 , \16763 );
and \U$8359 ( \17178 , \17177 , \9759 );
not \U$8360 ( \17179 , \16742 );
not \U$8361 ( \17180 , \17179 );
and \U$8362 ( \17181 , \9763 , \17180 );
nor \U$8363 ( \17182 , \17178 , \17181 );
nand \U$8364 ( \17183 , \17173 , \17176 , \17182 );
or \U$8365 ( \17184 , \10188 , \16954 );
not \U$8366 ( \17185 , \16918 );
or \U$8367 ( \17186 , \10178 , \17185 );
not \U$8368 ( \17187 , \16796 );
or \U$8369 ( \17188 , \10182 , \17187 );
not \U$8370 ( \17189 , \16813 );
or \U$8371 ( \17190 , \11186 , \17189 );
and \U$8372 ( \17191 , \17184 , \17186 , \17188 , \17190 );
not \U$8373 ( \17192 , \17191 );
nor \U$8374 ( \17193 , \17183 , \17192 );
nand \U$8375 ( \17194 , \17160 , \17171 , \17193 );
xnor \U$8376 ( \17195 , RIb7af4c8_257, \17194 );
or \U$8377 ( \17196 , \9658 , \16801 );
or \U$8378 ( \17197 , \9661 , \16750 );
nand \U$8379 ( \17198 , \17196 , \17197 );
or \U$8380 ( \17199 , \13344 , \16806 );
not \U$8381 ( \17200 , \16864 );
or \U$8382 ( \17201 , \9668 , \17200 );
nand \U$8383 ( \17202 , \17199 , \17201 );
nor \U$8384 ( \17203 , \17198 , \17202 );
not \U$8385 ( \17204 , \16781 );
or \U$8386 ( \17205 , \9676 , \17204 );
not \U$8387 ( \17206 , \16786 );
or \U$8388 ( \17207 , \11923 , \17206 );
nand \U$8389 ( \17208 , \17205 , \17207 );
not \U$8390 ( \17209 , \16898 );
or \U$8391 ( \17210 , \9680 , \17209 );
not \U$8392 ( \17211 , \16896 );
or \U$8393 ( \17212 , \9683 , \17211 );
nand \U$8394 ( \17213 , \17210 , \17212 );
nor \U$8395 ( \17214 , \17208 , \17213 );
not \U$8396 ( \17215 , \16737 );
or \U$8397 ( \17216 , \11152 , \17215 );
not \U$8398 ( \17217 , \17174 );
or \U$8399 ( \17218 , \11154 , \17217 );
not \U$8400 ( \17219 , \16762 );
not \U$8401 ( \17220 , \17219 );
and \U$8402 ( \17221 , \17220 , \9692 );
not \U$8403 ( \17222 , \17179 );
and \U$8404 ( \17223 , \9695 , \17222 );
nor \U$8405 ( \17224 , \17221 , \17223 );
nand \U$8406 ( \17225 , \17216 , \17218 , \17224 );
or \U$8407 ( \17226 , \10244 , \16954 );
not \U$8408 ( \17227 , \16918 );
or \U$8409 ( \17228 , \11138 , \17227 );
not \U$8410 ( \17229 , \16877 );
or \U$8411 ( \17230 , \11140 , \17229 );
not \U$8412 ( \17231 , \16812 );
not \U$8413 ( \17232 , \17231 );
or \U$8414 ( \17233 , \11145 , \17232 );
and \U$8415 ( \17234 , \17226 , \17228 , \17230 , \17233 );
not \U$8416 ( \17235 , \17234 );
nor \U$8417 ( \17236 , \17225 , \17235 );
nand \U$8418 ( \17237 , \17203 , \17214 , \17236 );
xnor \U$8419 ( \17238 , RIb7af5b8_255, \17237 );
or \U$8420 ( \17239 , \9552 , \16840 );
not \U$8421 ( \17240 , \16762 );
or \U$8422 ( \17241 , \9557 , \17240 );
nand \U$8423 ( \17242 , \17239 , \17241 );
or \U$8424 ( \17243 , \9564 , \16844 );
or \U$8425 ( \17244 , \11582 , \16882 );
nand \U$8426 ( \17245 , \17243 , \17244 );
nor \U$8427 ( \17246 , \17242 , \17245 );
or \U$8428 ( \17247 , \9569 , \16801 );
or \U$8429 ( \17248 , \9572 , \16750 );
nand \U$8430 ( \17249 , \17247 , \17248 );
or \U$8431 ( \17250 , \11589 , \16806 );
not \U$8432 ( \17251 , \16864 );
or \U$8433 ( \17252 , \9579 , \17251 );
nand \U$8434 ( \17253 , \17250 , \17252 );
nor \U$8435 ( \17254 , \17249 , \17253 );
not \U$8436 ( \17255 , \16781 );
or \U$8437 ( \17256 , \13658 , \17255 );
not \U$8438 ( \17257 , \16786 );
or \U$8439 ( \17258 , \9527 , \17257 );
and \U$8440 ( \17259 , \16896 , \9523 );
and \U$8441 ( \17260 , \16898 , \9518 );
nor \U$8442 ( \17261 , \17259 , \17260 );
nand \U$8443 ( \17262 , \17256 , \17258 , \17261 );
or \U$8444 ( \17263 , \9543 , \16954 );
not \U$8445 ( \17264 , \16918 );
or \U$8446 ( \17265 , \9534 , \17264 );
not \U$8447 ( \17266 , \16877 );
or \U$8448 ( \17267 , \9537 , \17266 );
not \U$8449 ( \17268 , \16813 );
or \U$8450 ( \17269 , \9546 , \17268 );
and \U$8451 ( \17270 , \17263 , \17265 , \17267 , \17269 );
not \U$8452 ( \17271 , \17270 );
nor \U$8453 ( \17272 , \17262 , \17271 );
nand \U$8454 ( \17273 , \17246 , \17254 , \17272 );
xnor \U$8455 ( \17274 , \17273 , \9585 );
or \U$8456 ( \17275 , \11618 , \16840 );
not \U$8457 ( \17276 , \16762 );
or \U$8458 ( \17277 , \11620 , \17276 );
nand \U$8459 ( \17278 , \17275 , \17277 );
or \U$8460 ( \17279 , \11623 , \16736 );
or \U$8461 ( \17280 , \11625 , \16746 );
nand \U$8462 ( \17281 , \17279 , \17280 );
nor \U$8463 ( \17282 , \17278 , \17281 );
or \U$8464 ( \17283 , \11635 , \16801 );
or \U$8465 ( \17284 , \11629 , \16750 );
nand \U$8466 ( \17285 , \17283 , \17284 );
or \U$8467 ( \17286 , \11633 , \16806 );
not \U$8468 ( \17287 , \16864 );
or \U$8469 ( \17288 , \12282 , \17287 );
nand \U$8470 ( \17289 , \17286 , \17288 );
nor \U$8471 ( \17290 , \17285 , \17289 );
not \U$8472 ( \17291 , \16781 );
or \U$8473 ( \17292 , \9948 , \17291 );
not \U$8474 ( \17293 , \16786 );
or \U$8475 ( \17294 , \13143 , \17293 );
and \U$8476 ( \17295 , \16896 , \9954 );
and \U$8477 ( \17296 , \16898 , \9951 );
nor \U$8478 ( \17297 , \17295 , \17296 );
nand \U$8479 ( \17298 , \17292 , \17294 , \17297 );
or \U$8480 ( \17299 , \9937 , \16954 );
not \U$8481 ( \17300 , \16918 );
or \U$8482 ( \17301 , \9930 , \17300 );
not \U$8483 ( \17302 , \16877 );
or \U$8484 ( \17303 , \9933 , \17302 );
not \U$8485 ( \17304 , \16813 );
or \U$8486 ( \17305 , \9940 , \17304 );
and \U$8487 ( \17306 , \17299 , \17301 , \17303 , \17305 );
not \U$8488 ( \17307 , \17306 );
nor \U$8489 ( \17308 , \17298 , \17307 );
nand \U$8490 ( \17309 , \17282 , \17290 , \17308 );
xnor \U$8491 ( \17310 , \17309 , \9990 );
nor \U$8492 ( \17311 , \17274 , \17310 );
nand \U$8493 ( \17312 , \17195 , \17238 , \17311 );
or \U$8494 ( \17313 , \9620 , \16840 );
not \U$8495 ( \17314 , \16762 );
or \U$8496 ( \17315 , \9625 , \17314 );
nand \U$8497 ( \17316 , \17313 , \17315 );
or \U$8498 ( \17317 , \9632 , \16736 );
or \U$8499 ( \17318 , \11314 , \16882 );
nand \U$8500 ( \17319 , \17317 , \17318 );
nor \U$8501 ( \17320 , \17316 , \17319 );
or \U$8502 ( \17321 , \9637 , \16801 );
or \U$8503 ( \17322 , \9640 , \16750 );
nand \U$8504 ( \17323 , \17321 , \17322 );
or \U$8505 ( \17324 , \11322 , \16806 );
not \U$8506 ( \17325 , \16769 );
or \U$8507 ( \17326 , \9647 , \17325 );
nand \U$8508 ( \17327 , \17324 , \17326 );
nor \U$8509 ( \17328 , \17323 , \17327 );
not \U$8510 ( \17329 , \16781 );
or \U$8511 ( \17330 , \13538 , \17329 );
not \U$8512 ( \17331 , \16786 );
or \U$8513 ( \17332 , \9597 , \17331 );
and \U$8514 ( \17333 , \16774 , \9593 );
and \U$8515 ( \17334 , \16792 , \9587 );
nor \U$8516 ( \17335 , \17333 , \17334 );
nand \U$8517 ( \17336 , \17330 , \17332 , \17335 );
or \U$8518 ( \17337 , \9611 , \16954 );
not \U$8519 ( \17338 , \16918 );
or \U$8520 ( \17339 , \9604 , \17338 );
not \U$8521 ( \17340 , \16796 );
or \U$8522 ( \17341 , \9607 , \17340 );
not \U$8523 ( \17342 , \17231 );
or \U$8524 ( \17343 , \9614 , \17342 );
and \U$8525 ( \17344 , \17337 , \17339 , \17341 , \17343 );
not \U$8526 ( \17345 , \17344 );
nor \U$8527 ( \17346 , \17336 , \17345 );
nand \U$8528 ( \17347 , \17320 , \17328 , \17346 );
xnor \U$8529 ( \17348 , RIb7af630_254, \17347 );
not \U$8530 ( \17349 , \16781 );
or \U$8531 ( \17350 , \11494 , \17349 );
not \U$8532 ( \17351 , \16786 );
or \U$8533 ( \17352 , \9798 , \17351 );
nand \U$8534 ( \17353 , \17350 , \17352 );
not \U$8535 ( \17354 , \16898 );
or \U$8536 ( \17355 , \9791 , \17354 );
not \U$8537 ( \17356 , \16896 );
or \U$8538 ( \17357 , \11492 , \17356 );
nand \U$8539 ( \17358 , \17355 , \17357 );
nor \U$8540 ( \17359 , \17353 , \17358 );
not \U$8541 ( \17360 , \17231 );
or \U$8542 ( \17361 , \17360 , \9817 );
or \U$8543 ( \17362 , \9814 , \16954 );
nand \U$8544 ( \17363 , \17361 , \17362 );
not \U$8545 ( \17364 , \17363 );
not \U$8546 ( \17365 , \16877 );
or \U$8547 ( \17366 , \9809 , \17365 );
not \U$8548 ( \17367 , \16918 );
or \U$8549 ( \17368 , \9806 , \17367 );
and \U$8550 ( \17369 , \17364 , \17366 , \17368 );
nand \U$8551 ( \17370 , \17359 , \17369 );
not \U$8552 ( \17371 , \11505 );
and \U$8553 ( \17372 , \17371 , \16807 );
and \U$8554 ( \17373 , \16769 , \9850 );
nor \U$8555 ( \17374 , \17372 , \17373 );
not \U$8556 ( \17375 , \9843 );
and \U$8557 ( \17376 , \17375 , \16856 );
and \U$8558 ( \17377 , \16859 , \9839 );
nor \U$8559 ( \17378 , \17376 , \17377 );
or \U$8560 ( \17379 , \9823 , \16840 );
not \U$8561 ( \17380 , \16762 );
or \U$8562 ( \17381 , \9827 , \17380 );
nand \U$8563 ( \17382 , \17379 , \17381 );
or \U$8564 ( \17383 , \9834 , \16844 );
or \U$8565 ( \17384 , \12311 , \16746 );
nand \U$8566 ( \17385 , \17383 , \17384 );
nor \U$8567 ( \17386 , \17382 , \17385 );
nand \U$8568 ( \17387 , \17374 , \17378 , \17386 );
nor \U$8569 ( \17388 , \17370 , \17387 );
xnor \U$8570 ( \17389 , \17388 , \9857 );
not \U$8571 ( \17390 , \16737 );
or \U$8572 ( \17391 , \11693 , \17390 );
not \U$8573 ( \17392 , \17174 );
or \U$8574 ( \17393 , \12235 , \17392 );
not \U$8575 ( \17394 , \17314 );
and \U$8576 ( \17395 , \17394 , \10030 );
not \U$8577 ( \17396 , \17179 );
and \U$8578 ( \17397 , \17396 , \10035 );
nor \U$8579 ( \17398 , \17395 , \17397 );
nand \U$8580 ( \17399 , \17391 , \17393 , \17398 );
not \U$8581 ( \17400 , \17399 );
or \U$8582 ( \17401 , \11684 , \16801 );
or \U$8583 ( \17402 , \12222 , \16750 );
nand \U$8584 ( \17403 , \17401 , \17402 );
or \U$8585 ( \17404 , \11681 , \16806 );
not \U$8586 ( \17405 , \16864 );
or \U$8587 ( \17406 , \11674 , \17405 );
nand \U$8588 ( \17407 , \17404 , \17406 );
nor \U$8589 ( \17408 , \17403 , \17407 );
or \U$8590 ( \17409 , \10018 , \16954 );
not \U$8591 ( \17410 , \16918 );
or \U$8592 ( \17411 , \10010 , \17410 );
not \U$8593 ( \17412 , \16796 );
or \U$8594 ( \17413 , \10013 , \17412 );
not \U$8595 ( \17414 , \16813 );
or \U$8596 ( \17415 , \10021 , \17414 );
and \U$8597 ( \17416 , \17409 , \17411 , \17413 , \17415 );
not \U$8598 ( \17417 , \17416 );
not \U$8599 ( \17418 , \16781 );
or \U$8600 ( \17419 , \9997 , \17418 );
not \U$8601 ( \17420 , \16786 );
or \U$8602 ( \17421 , \11666 , \17420 );
not \U$8603 ( \17422 , \16773 );
and \U$8604 ( \17423 , \17422 , \10004 );
not \U$8605 ( \17424 , \16791 );
and \U$8606 ( \17425 , \17424 , \10001 );
nor \U$8607 ( \17426 , \17423 , \17425 );
nand \U$8608 ( \17427 , \17419 , \17421 , \17426 );
nor \U$8609 ( \17428 , \17417 , \17427 );
nand \U$8610 ( \17429 , \17400 , \17408 , \17428 );
xnor \U$8611 ( \17430 , \17429 , \10055 );
or \U$8612 ( \17431 , \9895 , \16840 );
not \U$8613 ( \17432 , \16762 );
or \U$8614 ( \17433 , \9898 , \17432 );
nand \U$8615 ( \17434 , \17431 , \17433 );
or \U$8616 ( \17435 , \9906 , \16970 );
or \U$8617 ( \17436 , \11711 , \16882 );
nand \U$8618 ( \17437 , \17435 , \17436 );
nor \U$8619 ( \17438 , \17434 , \17437 );
or \U$8620 ( \17439 , \9911 , \16801 );
or \U$8621 ( \17440 , \9914 , \16750 );
nand \U$8622 ( \17441 , \17439 , \17440 );
or \U$8623 ( \17442 , \11718 , \16806 );
nand \U$8624 ( \17443 , \9920 , \16864 );
nand \U$8625 ( \17444 , \17442 , \17443 );
nor \U$8626 ( \17445 , \17441 , \17444 );
nand \U$8627 ( \17446 , \9871 , \16781 );
nand \U$8628 ( \17447 , \9867 , \16786 );
and \U$8629 ( \17448 , \16774 , \9864 );
and \U$8630 ( \17449 , \16792 , \9859 );
nor \U$8631 ( \17450 , \17448 , \17449 );
nand \U$8632 ( \17451 , \17446 , \17447 , \17450 );
or \U$8633 ( \17452 , \9884 , \16954 );
nand \U$8634 ( \17453 , \9874 , \16918 );
nand \U$8635 ( \17454 , \9877 , \16877 );
nand \U$8636 ( \17455 , \9886 , \17231 );
and \U$8637 ( \17456 , \17452 , \17453 , \17454 , \17455 );
not \U$8638 ( \17457 , \17456 );
nor \U$8639 ( \17458 , \17451 , \17457 );
nand \U$8640 ( \17459 , \17438 , \17445 , \17458 );
xnor \U$8641 ( \17460 , \17459 , \9927 );
nor \U$8642 ( \17461 , \17430 , \17460 );
nand \U$8643 ( \17462 , \17348 , \17389 , \17461 );
nor \U$8644 ( \17463 , \17312 , \17462 );
nand \U$8645 ( \17464 , \16825 , \17152 , \17463 );
not \U$8646 ( \17465 , \17464 );
not \U$8647 ( \17466 , \17465 );
or \U$8648 ( \17467 , \16730 , \17466 );
not \U$8649 ( \17468 , \17467 );
nand \U$8650 ( \17469 , \16730 , \17465 );
not \U$8651 ( \17470 , \17469 );
or \U$8652 ( \17471 , \17468 , \17470 );
not \U$8653 ( \17472 , \17471 );
not \U$8654 ( \17473 , \17472 );
and \U$8655 ( \17474 , \16704 , \17473 );
buf \U$8656 ( \17475 , \13253 );
buf \U$8657 ( \17476 , \12456 );
buf \U$8658 ( \17477 , \12458 );
buf \U$8659 ( \17478 , \10919 );
or \U$8660 ( \17479 , \17477 , \17478 );
or \U$8661 ( \17480 , \17476 , \17479 );
xnor \U$8662 ( \17481 , \17475 , \17480 );
buf \U$8663 ( \17482 , \17481 );
not \U$8664 ( \17483 , \17482 );
xnor \U$8665 ( \17484 , \17476 , \17479 );
buf \U$8666 ( \17485 , \17484 );
xnor \U$8667 ( \17486 , \17477 , \17478 );
buf \U$8668 ( \17487 , \17486 );
not \U$8669 ( \17488 , \17478 );
buf \U$8670 ( \17489 , \17488 );
nor \U$8671 ( \17490 , \17485 , \17487 , \17489 );
and \U$8672 ( \17491 , \17483 , \17490 );
buf \U$8673 ( \17492 , RIea91330_6888);
or \U$8674 ( \17493 , \17475 , \17480 );
xor \U$8675 ( \17494 , \17492 , \17493 );
buf \U$8676 ( \17495 , \17494 );
not \U$8677 ( \17496 , \17495 );
or \U$8678 ( \17497 , \17491 , \17496 );
and \U$8679 ( \17498 , \17492 , \17493 );
buf \U$8680 ( \17499 , \17498 );
not \U$8681 ( \17500 , \17499 );
nand \U$8682 ( \17501 , \17497 , \17500 );
not \U$8683 ( \17502 , \17501 );
not \U$8684 ( \17503 , \9482 );
nand \U$8685 ( \17504 , \8906 , \10077 );
not \U$8686 ( \17505 , \10078 );
or \U$8687 ( \17506 , \8906 , \17505 );
nand \U$8688 ( \17507 , \17504 , \17506 );
not \U$8689 ( \17508 , \17507 );
and \U$8690 ( \17509 , \17508 , \11753 );
not \U$8691 ( \17510 , \17509 );
or \U$8692 ( \17511 , \10939 , \17510 );
not \U$8693 ( \17512 , \17511 );
and \U$8694 ( \17513 , \17503 , \17512 );
nand \U$8695 ( \17514 , \11753 , \17507 );
not \U$8696 ( \17515 , \17514 );
not \U$8697 ( \17516 , \17515 );
or \U$8698 ( \17517 , \10925 , \17516 );
not \U$8699 ( \17518 , \17517 );
not \U$8700 ( \17519 , \17518 );
or \U$8701 ( \17520 , \9485 , \17519 );
not \U$8702 ( \17521 , \17515 );
or \U$8703 ( \17522 , \17521 , \10939 );
or \U$8704 ( \17523 , \9487 , \17522 );
nand \U$8705 ( \17524 , \17520 , \17523 );
and \U$8706 ( \17525 , \17508 , \11752 );
not \U$8707 ( \17526 , \17525 );
or \U$8708 ( \17527 , \10925 , \17526 );
not \U$8709 ( \17528 , \17527 );
and \U$8710 ( \17529 , \9468 , \17528 );
or \U$8711 ( \17530 , \17513 , \17524 , \17529 );
not \U$8712 ( \17531 , \17530 );
not \U$8713 ( \17532 , \17509 );
or \U$8714 ( \17533 , \10958 , \17532 );
or \U$8715 ( \17534 , \9475 , \17533 );
not \U$8716 ( \17535 , \17509 );
or \U$8717 ( \17536 , \10949 , \17535 );
or \U$8718 ( \17537 , \9471 , \17536 );
nand \U$8719 ( \17538 , \17534 , \17537 );
not \U$8720 ( \17539 , \17525 );
or \U$8721 ( \17540 , \10958 , \17539 );
or \U$8722 ( \17541 , \9463 , \17540 );
and \U$8723 ( \17542 , \11752 , \17507 );
not \U$8724 ( \17543 , \17542 );
or \U$8725 ( \17544 , \10949 , \17543 );
or \U$8726 ( \17545 , \9480 , \17544 );
nand \U$8727 ( \17546 , \17541 , \17545 );
nor \U$8728 ( \17547 , \17538 , \17546 );
not \U$8729 ( \17548 , \17542 );
or \U$8730 ( \17549 , \17548 , \10925 );
not \U$8731 ( \17550 , \17549 );
not \U$8732 ( \17551 , \17550 );
or \U$8733 ( \17552 , \9498 , \17551 );
not \U$8734 ( \17553 , \17542 );
or \U$8735 ( \17554 , \10939 , \17553 );
not \U$8736 ( \17555 , \17554 );
not \U$8737 ( \17556 , \17555 );
or \U$8738 ( \17557 , \17556 , \9500 );
not \U$8739 ( \17558 , \17515 );
or \U$8740 ( \17559 , \17558 , \10958 );
not \U$8741 ( \17560 , \17559 );
and \U$8742 ( \17561 , \17560 , \10062 );
not \U$8743 ( \17562 , \17515 );
or \U$8744 ( \17563 , \10949 , \17562 );
not \U$8745 ( \17564 , \17563 );
and \U$8746 ( \17565 , \12513 , \17564 );
nor \U$8747 ( \17566 , \17561 , \17565 );
nand \U$8748 ( \17567 , \17552 , \17557 , \17566 );
not \U$8749 ( \17568 , \17567 );
not \U$8750 ( \17569 , \9506 );
not \U$8751 ( \17570 , \17542 );
or \U$8752 ( \17571 , \10958 , \17570 );
not \U$8753 ( \17572 , \17571 );
and \U$8754 ( \17573 , \17569 , \17572 );
not \U$8755 ( \17574 , \17509 );
or \U$8756 ( \17575 , \10925 , \17574 );
not \U$8757 ( \17576 , \17575 );
and \U$8758 ( \17577 , \17576 , \10976 );
nor \U$8759 ( \17578 , \17573 , \17577 );
not \U$8760 ( \17579 , \9511 );
not \U$8761 ( \17580 , \17525 );
or \U$8762 ( \17581 , \10939 , \17580 );
not \U$8763 ( \17582 , \17581 );
not \U$8764 ( \17583 , \17582 );
not \U$8765 ( \17584 , \17583 );
and \U$8766 ( \17585 , \17579 , \17584 );
not \U$8767 ( \17586 , \17525 );
or \U$8768 ( \17587 , \10949 , \17586 );
not \U$8769 ( \17588 , \17587 );
and \U$8770 ( \17589 , \17588 , \13270 );
nor \U$8771 ( \17590 , \17585 , \17589 );
and \U$8772 ( \17591 , \17568 , \17578 , \17590 );
nand \U$8773 ( \17592 , \17531 , \17547 , \17591 );
not \U$8774 ( \17593 , \17592 );
not \U$8775 ( \17594 , \9107 );
or \U$8776 ( \17595 , \17594 , \17571 );
not \U$8777 ( \17596 , \17509 );
or \U$8778 ( \17597 , \17596 , \10939 );
or \U$8779 ( \17598 , \9050 , \17597 );
nand \U$8780 ( \17599 , \17595 , \17598 );
not \U$8781 ( \17600 , \17509 );
or \U$8782 ( \17601 , \10958 , \17600 );
or \U$8783 ( \17602 , \9086 , \17601 );
not \U$8784 ( \17603 , \17576 );
or \U$8785 ( \17604 , \9058 , \17603 );
nand \U$8786 ( \17605 , \17602 , \17604 );
nor \U$8787 ( \17606 , \17599 , \17605 );
or \U$8788 ( \17607 , \11468 , \17563 );
or \U$8789 ( \17608 , \9082 , \17559 );
nand \U$8790 ( \17609 , \17607 , \17608 );
or \U$8791 ( \17610 , \11471 , \17549 );
not \U$8792 ( \17611 , \17542 );
or \U$8793 ( \17612 , \17611 , \10939 );
or \U$8794 ( \17613 , \11466 , \17612 );
nand \U$8795 ( \17614 , \17610 , \17613 );
nor \U$8796 ( \17615 , \17609 , \17614 );
not \U$8797 ( \17616 , \9068 );
not \U$8798 ( \17617 , \17527 );
and \U$8799 ( \17618 , \17616 , \17617 );
and \U$8800 ( \17619 , \17582 , \9075 );
nor \U$8801 ( \17620 , \17618 , \17619 );
not \U$8802 ( \17621 , \10859 );
not \U$8803 ( \17622 , \17542 );
or \U$8804 ( \17623 , \17622 , \10949 );
not \U$8805 ( \17624 , \17623 );
and \U$8806 ( \17625 , \17621 , \17624 );
not \U$8807 ( \17626 , \17540 );
and \U$8808 ( \17627 , \17626 , \9063 );
nor \U$8809 ( \17628 , \17625 , \17627 );
nand \U$8810 ( \17629 , \17620 , \17628 );
not \U$8811 ( \17630 , \17629 );
not \U$8812 ( \17631 , \9073 );
not \U$8813 ( \17632 , \17536 );
and \U$8814 ( \17633 , \17631 , \17632 );
and \U$8815 ( \17634 , \17588 , \9098 );
nor \U$8816 ( \17635 , \17633 , \17634 );
not \U$8817 ( \17636 , \17522 );
and \U$8818 ( \17637 , \9046 , \17636 );
not \U$8819 ( \17638 , \17518 );
not \U$8820 ( \17639 , \17638 );
and \U$8821 ( \17640 , \17639 , \9054 );
nor \U$8822 ( \17641 , \17637 , \17640 );
and \U$8823 ( \17642 , \17630 , \17635 , \17641 );
nand \U$8824 ( \17643 , \17606 , \17615 , \17642 );
xnor \U$8825 ( \17644 , RIb7af720_252, \17643 );
not \U$8826 ( \17645 , \8947 );
not \U$8827 ( \17646 , \17542 );
or \U$8828 ( \17647 , \10958 , \17646 );
or \U$8829 ( \17648 , \17645 , \17647 );
or \U$8830 ( \17649 , \8844 , \17511 );
nand \U$8831 ( \17650 , \17648 , \17649 );
or \U$8832 ( \17651 , \11533 , \17533 );
or \U$8833 ( \17652 , \8861 , \17603 );
nand \U$8834 ( \17653 , \17651 , \17652 );
nor \U$8835 ( \17654 , \17650 , \17653 );
not \U$8836 ( \17655 , \17515 );
or \U$8837 ( \17656 , \10949 , \17655 );
or \U$8838 ( \17657 , \11540 , \17656 );
not \U$8839 ( \17658 , \17515 );
or \U$8840 ( \17659 , \17658 , \10958 );
or \U$8841 ( \17660 , \11528 , \17659 );
nand \U$8842 ( \17661 , \17657 , \17660 );
not \U$8843 ( \17662 , \17542 );
or \U$8844 ( \17663 , \10925 , \17662 );
or \U$8845 ( \17664 , \14573 , \17663 );
or \U$8846 ( \17665 , \13894 , \17554 );
nand \U$8847 ( \17666 , \17664 , \17665 );
nor \U$8848 ( \17667 , \17661 , \17666 );
not \U$8849 ( \17668 , \8882 );
and \U$8850 ( \17669 , \17668 , \17617 );
and \U$8851 ( \17670 , \17582 , \8896 );
nor \U$8852 ( \17671 , \17669 , \17670 );
not \U$8853 ( \17672 , \10775 );
and \U$8854 ( \17673 , \17672 , \17624 );
not \U$8855 ( \17674 , \17540 );
and \U$8856 ( \17675 , \17674 , \8868 );
nor \U$8857 ( \17676 , \17673 , \17675 );
nand \U$8858 ( \17677 , \17671 , \17676 );
not \U$8859 ( \17678 , \17677 );
not \U$8860 ( \17679 , \8894 );
not \U$8861 ( \17680 , \17536 );
and \U$8862 ( \17681 , \17679 , \17680 );
and \U$8863 ( \17682 , \17588 , \8934 );
nor \U$8864 ( \17683 , \17681 , \17682 );
not \U$8865 ( \17684 , \17515 );
or \U$8866 ( \17685 , \17684 , \10939 );
not \U$8867 ( \17686 , \17685 );
and \U$8868 ( \17687 , \8827 , \17686 );
not \U$8869 ( \17688 , \17638 );
and \U$8870 ( \17689 , \17688 , \8852 );
nor \U$8871 ( \17690 , \17687 , \17689 );
and \U$8872 ( \17691 , \17678 , \17683 , \17690 );
nand \U$8873 ( \17692 , \17654 , \17667 , \17691 );
xnor \U$8874 ( \17693 , RIb7b93b0_251, \17692 );
not \U$8875 ( \17694 , \9247 );
or \U$8876 ( \17695 , \17694 , \17571 );
or \U$8877 ( \17696 , \11088 , \17597 );
nand \U$8878 ( \17697 , \17695 , \17696 );
or \U$8879 ( \17698 , \11125 , \17533 );
or \U$8880 ( \17699 , \11954 , \17603 );
nand \U$8881 ( \17700 , \17698 , \17699 );
nor \U$8882 ( \17701 , \17697 , \17700 );
or \U$8883 ( \17702 , \11113 , \17563 );
or \U$8884 ( \17703 , \9226 , \17559 );
nand \U$8885 ( \17704 , \17702 , \17703 );
or \U$8886 ( \17705 , \11117 , \17549 );
or \U$8887 ( \17706 , \11111 , \17554 );
nand \U$8888 ( \17707 , \17705 , \17706 );
nor \U$8889 ( \17708 , \17704 , \17707 );
not \U$8890 ( \17709 , \11098 );
and \U$8891 ( \17710 , \17709 , \17617 );
and \U$8892 ( \17711 , \17582 , \9219 );
nor \U$8893 ( \17712 , \17710 , \17711 );
not \U$8894 ( \17713 , \10323 );
and \U$8895 ( \17714 , \17713 , \17624 );
and \U$8896 ( \17715 , \17626 , \9210 );
nor \U$8897 ( \17716 , \17714 , \17715 );
nand \U$8898 ( \17717 , \17712 , \17716 );
not \U$8899 ( \17718 , \17717 );
not \U$8900 ( \17719 , \9217 );
and \U$8901 ( \17720 , \17719 , \17680 );
and \U$8902 ( \17721 , \17588 , \9239 );
nor \U$8903 ( \17722 , \17720 , \17721 );
not \U$8904 ( \17723 , \17522 );
and \U$8905 ( \17724 , \9196 , \17723 );
not \U$8906 ( \17725 , \17638 );
and \U$8907 ( \17726 , \17725 , \9204 );
nor \U$8908 ( \17727 , \17724 , \17726 );
and \U$8909 ( \17728 , \17718 , \17722 , \17727 );
nand \U$8910 ( \17729 , \17701 , \17708 , \17728 );
xnor \U$8911 ( \17730 , \17729 , \9260 );
not \U$8912 ( \17731 , \9030 );
not \U$8913 ( \17732 , \17542 );
or \U$8914 ( \17733 , \10958 , \17732 );
or \U$8915 ( \17734 , \17731 , \17733 );
not \U$8916 ( \17735 , \17509 );
or \U$8917 ( \17736 , \17735 , \10939 );
or \U$8918 ( \17737 , \8971 , \17736 );
nand \U$8919 ( \17738 , \17734 , \17737 );
or \U$8920 ( \17739 , \11073 , \17601 );
or \U$8921 ( \17740 , \8980 , \17603 );
nand \U$8922 ( \17741 , \17739 , \17740 );
nor \U$8923 ( \17742 , \17738 , \17741 );
not \U$8924 ( \17743 , \17515 );
or \U$8925 ( \17744 , \17743 , \10949 );
or \U$8926 ( \17745 , \11060 , \17744 );
not \U$8927 ( \17746 , \17515 );
or \U$8928 ( \17747 , \17746 , \10958 );
or \U$8929 ( \17748 , \11080 , \17747 );
nand \U$8930 ( \17749 , \17745 , \17748 );
not \U$8931 ( \17750 , \17542 );
or \U$8932 ( \17751 , \10925 , \17750 );
or \U$8933 ( \17752 , \11064 , \17751 );
or \U$8934 ( \17753 , \11058 , \17612 );
nand \U$8935 ( \17754 , \17752 , \17753 );
nor \U$8936 ( \17755 , \17749 , \17754 );
not \U$8937 ( \17756 , \8991 );
and \U$8938 ( \17757 , \17756 , \17617 );
and \U$8939 ( \17758 , \17582 , \8999 );
nor \U$8940 ( \17759 , \17757 , \17758 );
not \U$8941 ( \17760 , \10370 );
and \U$8942 ( \17761 , \17760 , \17624 );
and \U$8943 ( \17762 , \17674 , \8986 );
nor \U$8944 ( \17763 , \17761 , \17762 );
nand \U$8945 ( \17764 , \17759 , \17763 );
not \U$8946 ( \17765 , \17764 );
not \U$8947 ( \17766 , \8997 );
and \U$8948 ( \17767 , \17766 , \17680 );
and \U$8949 ( \17768 , \17588 , \9020 );
nor \U$8950 ( \17769 , \17767 , \17768 );
not \U$8951 ( \17770 , \17515 );
or \U$8952 ( \17771 , \17770 , \10939 );
not \U$8953 ( \17772 , \17771 );
and \U$8954 ( \17773 , \8966 , \17772 );
not \U$8955 ( \17774 , \17638 );
and \U$8956 ( \17775 , \17774 , \8976 );
nor \U$8957 ( \17776 , \17773 , \17775 );
and \U$8958 ( \17777 , \17765 , \17769 , \17776 );
nand \U$8959 ( \17778 , \17742 , \17755 , \17777 );
xnor \U$8960 ( \17779 , \17778 , \9044 );
nor \U$8961 ( \17780 , \17730 , \17779 );
nand \U$8962 ( \17781 , \17644 , \17693 , \17780 );
not \U$8963 ( \17782 , \17781 );
not \U$8964 ( \17783 , \9315 );
or \U$8965 ( \17784 , \17783 , \17733 );
or \U$8966 ( \17785 , \9266 , \17736 );
nand \U$8967 ( \17786 , \17784 , \17785 );
or \U$8968 ( \17787 , \11298 , \17533 );
or \U$8969 ( \17788 , \9273 , \17603 );
nand \U$8970 ( \17789 , \17787 , \17788 );
nor \U$8971 ( \17790 , \17786 , \17789 );
or \U$8972 ( \17791 , \11288 , \17744 );
or \U$8973 ( \17792 , \11303 , \17747 );
nand \U$8974 ( \17793 , \17791 , \17792 );
or \U$8975 ( \17794 , \11291 , \17751 );
or \U$8976 ( \17795 , \11286 , \17554 );
nand \U$8977 ( \17796 , \17794 , \17795 );
nor \U$8978 ( \17797 , \17793 , \17796 );
not \U$8979 ( \17798 , \9282 );
and \U$8980 ( \17799 , \17798 , \17617 );
and \U$8981 ( \17800 , \17582 , \9289 );
nor \U$8982 ( \17801 , \17799 , \17800 );
not \U$8983 ( \17802 , \10415 );
and \U$8984 ( \17803 , \17802 , \17624 );
and \U$8985 ( \17804 , \17674 , \9277 );
nor \U$8986 ( \17805 , \17803 , \17804 );
nand \U$8987 ( \17806 , \17801 , \17805 );
not \U$8988 ( \17807 , \17806 );
not \U$8989 ( \17808 , \9287 );
and \U$8990 ( \17809 , \17808 , \17680 );
and \U$8991 ( \17810 , \17588 , \9307 );
nor \U$8992 ( \17811 , \17809 , \17810 );
not \U$8993 ( \17812 , \17771 );
and \U$8994 ( \17813 , \9262 , \17812 );
not \U$8995 ( \17814 , \17638 );
and \U$8996 ( \17815 , \17814 , \9269 );
nor \U$8997 ( \17816 , \17813 , \17815 );
and \U$8998 ( \17817 , \17807 , \17811 , \17816 );
nand \U$8999 ( \17818 , \17790 , \17797 , \17817 );
xnor \U$9000 ( \17819 , \17818 , \9327 );
not \U$9001 ( \17820 , \9449 );
or \U$9002 ( \17821 , \17820 , \17647 );
or \U$9003 ( \17822 , \9398 , \17511 );
nand \U$9004 ( \17823 , \17821 , \17822 );
or \U$9005 ( \17824 , \10464 , \17601 );
not \U$9006 ( \17825 , \17576 );
or \U$9007 ( \17826 , \9405 , \17825 );
nand \U$9008 ( \17827 , \17824 , \17826 );
nor \U$9009 ( \17828 , \17823 , \17827 );
or \U$9010 ( \17829 , \11245 , \17656 );
or \U$9011 ( \17830 , \11259 , \17659 );
nand \U$9012 ( \17831 , \17829 , \17830 );
or \U$9013 ( \17832 , \11248 , \17663 );
or \U$9014 ( \17833 , \11243 , \17612 );
nand \U$9015 ( \17834 , \17832 , \17833 );
nor \U$9016 ( \17835 , \17831 , \17834 );
not \U$9017 ( \17836 , \9415 );
and \U$9018 ( \17837 , \17836 , \17617 );
and \U$9019 ( \17838 , \17582 , \9421 );
nor \U$9020 ( \17839 , \17837 , \17838 );
not \U$9021 ( \17840 , \10462 );
and \U$9022 ( \17841 , \17840 , \17624 );
and \U$9023 ( \17842 , \17626 , \9409 );
nor \U$9024 ( \17843 , \17841 , \17842 );
nand \U$9025 ( \17844 , \17839 , \17843 );
not \U$9026 ( \17845 , \17844 );
not \U$9027 ( \17846 , \9419 );
and \U$9028 ( \17847 , \17846 , \17680 );
and \U$9029 ( \17848 , \17588 , \9440 );
nor \U$9030 ( \17849 , \17847 , \17848 );
not \U$9031 ( \17850 , \17685 );
and \U$9032 ( \17851 , \9394 , \17850 );
not \U$9033 ( \17852 , \17519 );
and \U$9034 ( \17853 , \9401 , \17852 );
nor \U$9035 ( \17854 , \17851 , \17853 );
and \U$9036 ( \17855 , \17845 , \17849 , \17854 );
nand \U$9037 ( \17856 , \17828 , \17835 , \17855 );
xnor \U$9038 ( \17857 , \17856 , \9460 );
nor \U$9039 ( \17858 , \17819 , \17857 );
not \U$9040 ( \17859 , \9385 );
or \U$9041 ( \17860 , \17859 , \17571 );
or \U$9042 ( \17861 , \9335 , \17597 );
nand \U$9043 ( \17862 , \17860 , \17861 );
or \U$9044 ( \17863 , \11357 , \17533 );
or \U$9045 ( \17864 , \9342 , \17603 );
nand \U$9046 ( \17865 , \17863 , \17864 );
nor \U$9047 ( \17866 , \17862 , \17865 );
or \U$9048 ( \17867 , \11365 , \17563 );
or \U$9049 ( \17868 , \11352 , \17559 );
nand \U$9050 ( \17869 , \17867 , \17868 );
or \U$9051 ( \17870 , \11371 , \17549 );
or \U$9052 ( \17871 , \13593 , \17554 );
nand \U$9053 ( \17872 , \17870 , \17871 );
nor \U$9054 ( \17873 , \17869 , \17872 );
not \U$9055 ( \17874 , \12139 );
and \U$9056 ( \17875 , \17874 , \17617 );
and \U$9057 ( \17876 , \17582 , \9356 );
nor \U$9058 ( \17877 , \17875 , \17876 );
not \U$9059 ( \17878 , \10553 );
and \U$9060 ( \17879 , \17878 , \17624 );
not \U$9061 ( \17880 , \17540 );
and \U$9062 ( \17881 , \17880 , \9346 );
nor \U$9063 ( \17882 , \17879 , \17881 );
nand \U$9064 ( \17883 , \17877 , \17882 );
not \U$9065 ( \17884 , \17883 );
not \U$9066 ( \17885 , \9354 );
and \U$9067 ( \17886 , \17885 , \17680 );
and \U$9068 ( \17887 , \17588 , \9374 );
nor \U$9069 ( \17888 , \17886 , \17887 );
not \U$9070 ( \17889 , \17522 );
and \U$9071 ( \17890 , \9331 , \17889 );
not \U$9072 ( \17891 , \17519 );
and \U$9073 ( \17892 , \17891 , \9338 );
nor \U$9074 ( \17893 , \17890 , \17892 );
and \U$9075 ( \17894 , \17884 , \17888 , \17893 );
nand \U$9076 ( \17895 , \17866 , \17873 , \17894 );
xnor \U$9077 ( \17896 , \17895 , \9392 );
not \U$9078 ( \17897 , \9176 );
or \U$9079 ( \17898 , \17897 , \17733 );
or \U$9080 ( \17899 , \9125 , \17736 );
nand \U$9081 ( \17900 , \17898 , \17899 );
or \U$9082 ( \17901 , \11436 , \17601 );
or \U$9083 ( \17902 , \9133 , \17825 );
nand \U$9084 ( \17903 , \17901 , \17902 );
nor \U$9085 ( \17904 , \17900 , \17903 );
or \U$9086 ( \17905 , \11426 , \17744 );
or \U$9087 ( \17906 , \11441 , \17747 );
nand \U$9088 ( \17907 , \17905 , \17906 );
or \U$9089 ( \17908 , \11429 , \17751 );
or \U$9090 ( \17909 , \11424 , \17612 );
nand \U$9091 ( \17910 , \17908 , \17909 );
nor \U$9092 ( \17911 , \17907 , \17910 );
not \U$9093 ( \17912 , \9143 );
and \U$9094 ( \17913 , \17912 , \17617 );
and \U$9095 ( \17914 , \17582 , \9150 );
nor \U$9096 ( \17915 , \17913 , \17914 );
not \U$9097 ( \17916 , \10901 );
and \U$9098 ( \17917 , \17916 , \17624 );
and \U$9099 ( \17918 , \17674 , \9137 );
nor \U$9100 ( \17919 , \17917 , \17918 );
nand \U$9101 ( \17920 , \17915 , \17919 );
not \U$9102 ( \17921 , \17920 );
not \U$9103 ( \17922 , \9148 );
and \U$9104 ( \17923 , \17922 , \17632 );
and \U$9105 ( \17924 , \17588 , \9168 );
nor \U$9106 ( \17925 , \17923 , \17924 );
not \U$9107 ( \17926 , \17771 );
and \U$9108 ( \17927 , \9121 , \17926 );
not \U$9109 ( \17928 , \17518 );
not \U$9110 ( \17929 , \17928 );
and \U$9111 ( \17930 , \17929 , \9129 );
nor \U$9112 ( \17931 , \17927 , \17930 );
and \U$9113 ( \17932 , \17921 , \17925 , \17931 );
nand \U$9114 ( \17933 , \17904 , \17911 , \17932 );
xnor \U$9115 ( \17934 , \17933 , \9188 );
nor \U$9116 ( \17935 , \17896 , \17934 );
and \U$9117 ( \17936 , \17782 , \17858 , \17935 );
not \U$9118 ( \17937 , \17555 );
or \U$9119 ( \17938 , \11195 , \17937 );
not \U$9120 ( \17939 , \17550 );
or \U$9121 ( \17940 , \10194 , \17939 );
not \U$9122 ( \17941 , \10197 );
and \U$9123 ( \17942 , \17941 , \17572 );
and \U$9124 ( \17943 , \17588 , \9731 );
nor \U$9125 ( \17944 , \17942 , \17943 );
nand \U$9126 ( \17945 , \17938 , \17940 , \17944 );
not \U$9127 ( \17946 , \17597 );
not \U$9128 ( \17947 , \17946 );
or \U$9129 ( \17948 , \11186 , \17947 );
not \U$9130 ( \17949 , \17576 );
or \U$9131 ( \17950 , \10178 , \17949 );
not \U$9132 ( \17951 , \17656 );
and \U$9133 ( \17952 , \17951 , \9752 );
not \U$9134 ( \17953 , \17601 );
and \U$9135 ( \17954 , \17953 , \9769 );
nor \U$9136 ( \17955 , \17952 , \17954 );
nand \U$9137 ( \17956 , \17948 , \17950 , \17955 );
nor \U$9138 ( \17957 , \17945 , \17956 );
not \U$9139 ( \17958 , \9740 );
and \U$9140 ( \17959 , \17958 , \17617 );
and \U$9141 ( \17960 , \17582 , \9747 );
nor \U$9142 ( \17961 , \17959 , \17960 );
not \U$9143 ( \17962 , \10188 );
and \U$9144 ( \17963 , \17962 , \17624 );
and \U$9145 ( \17964 , \17626 , \9736 );
nor \U$9146 ( \17965 , \17963 , \17964 );
nand \U$9147 ( \17966 , \17961 , \17965 );
not \U$9148 ( \17967 , \17966 );
not \U$9149 ( \17968 , \9725 );
not \U$9150 ( \17969 , \17559 );
and \U$9151 ( \17970 , \17968 , \17969 );
and \U$9152 ( \17971 , \17680 , \9744 );
nor \U$9153 ( \17972 , \17970 , \17971 );
not \U$9154 ( \17973 , \17519 );
and \U$9155 ( \17974 , \9721 , \17973 );
not \U$9156 ( \17975 , \17685 );
and \U$9157 ( \17976 , \9728 , \17975 );
nor \U$9158 ( \17977 , \17974 , \17976 );
and \U$9159 ( \17978 , \17967 , \17972 , \17977 );
nand \U$9160 ( \17979 , \17957 , \17978 );
xnor \U$9161 ( \17980 , RIb7af4c8_257, \17979 );
or \U$9162 ( \17981 , \9658 , \17519 );
or \U$9163 ( \17982 , \9661 , \17659 );
nand \U$9164 ( \17983 , \17981 , \17982 );
or \U$9165 ( \17984 , \9668 , \17587 );
or \U$9166 ( \17985 , \13344 , \17771 );
nand \U$9167 ( \17986 , \17984 , \17985 );
nor \U$9168 ( \17987 , \17983 , \17986 );
not \U$9169 ( \17988 , \17617 );
or \U$9170 ( \17989 , \9676 , \17988 );
not \U$9171 ( \17990 , \17880 );
or \U$9172 ( \17991 , \11923 , \17990 );
nand \U$9173 ( \17992 , \17989 , \17991 );
not \U$9174 ( \17993 , \17632 );
or \U$9175 ( \17994 , \9680 , \17993 );
not \U$9176 ( \17995 , \17582 );
or \U$9177 ( \17996 , \9683 , \17995 );
nand \U$9178 ( \17997 , \17994 , \17996 );
nor \U$9179 ( \17998 , \17992 , \17997 );
nand \U$9180 ( \17999 , \17987 , \17998 );
not \U$9181 ( \18000 , \11138 );
and \U$9182 ( \18001 , \18000 , \17576 );
and \U$9183 ( \18002 , \17946 , \9710 );
nor \U$9184 ( \18003 , \18001 , \18002 );
not \U$9185 ( \18004 , \10244 );
and \U$9186 ( \18005 , \18004 , \17624 );
not \U$9187 ( \18006 , \17601 );
and \U$9188 ( \18007 , \18006 , \9701 );
nor \U$9189 ( \18008 , \18005 , \18007 );
or \U$9190 ( \18009 , \10248 , \17663 );
or \U$9191 ( \18010 , \10250 , \17647 );
nand \U$9192 ( \18011 , \18009 , \18010 );
not \U$9193 ( \18012 , \9690 );
or \U$9194 ( \18013 , \18012 , \17612 );
or \U$9195 ( \18014 , \11152 , \17744 );
nand \U$9196 ( \18015 , \18013 , \18014 );
nor \U$9197 ( \18016 , \18011 , \18015 );
nand \U$9198 ( \18017 , \18003 , \18008 , \18016 );
nor \U$9199 ( \18018 , \17999 , \18017 );
xnor \U$9200 ( \18019 , \18018 , \9719 );
or \U$9201 ( \18020 , \9537 , \17533 );
or \U$9202 ( \18021 , \9519 , \17536 );
nand \U$9203 ( \18022 , \18020 , \18021 );
or \U$9204 ( \18023 , \9546 , \17736 );
or \U$9205 ( \18024 , \9534 , \17825 );
nand \U$9206 ( \18025 , \18023 , \18024 );
nor \U$9207 ( \18026 , \18022 , \18025 );
or \U$9208 ( \18027 , \9527 , \17540 );
or \U$9209 ( \18028 , \9543 , \17623 );
nand \U$9210 ( \18029 , \18027 , \18028 );
not \U$9211 ( \18030 , \17582 );
or \U$9212 ( \18031 , \14434 , \18030 );
not \U$9213 ( \18032 , \17617 );
or \U$9214 ( \18033 , \13658 , \18032 );
nand \U$9215 ( \18034 , \18031 , \18033 );
nor \U$9216 ( \18035 , \18029 , \18034 );
not \U$9217 ( \18036 , \17587 );
not \U$9218 ( \18037 , \18036 );
or \U$9219 ( \18038 , \9579 , \18037 );
not \U$9220 ( \18039 , \17685 );
not \U$9221 ( \18040 , \18039 );
or \U$9222 ( \18041 , \11589 , \18040 );
not \U$9223 ( \18042 , \17659 );
and \U$9224 ( \18043 , \18042 , \9571 );
not \U$9225 ( \18044 , \17928 );
and \U$9226 ( \18045 , \18044 , \9568 );
nor \U$9227 ( \18046 , \18043 , \18045 );
nand \U$9228 ( \18047 , \18038 , \18041 , \18046 );
not \U$9229 ( \18048 , \9564 );
not \U$9230 ( \18049 , \17744 );
and \U$9231 ( \18050 , \18048 , \18049 );
and \U$9232 ( \18051 , \17555 , \9560 );
nor \U$9233 ( \18052 , \18050 , \18051 );
not \U$9234 ( \18053 , \9557 );
and \U$9235 ( \18054 , \18053 , \17572 );
and \U$9236 ( \18055 , \17550 , \9551 );
nor \U$9237 ( \18056 , \18054 , \18055 );
nand \U$9238 ( \18057 , \18052 , \18056 );
nor \U$9239 ( \18058 , \18047 , \18057 );
nand \U$9240 ( \18059 , \18026 , \18035 , \18058 );
xnor \U$9241 ( \18060 , \18059 , \9585 );
or \U$9242 ( \18061 , \9933 , \17601 );
or \U$9243 ( \18062 , \9952 , \17536 );
nand \U$9244 ( \18063 , \18061 , \18062 );
or \U$9245 ( \18064 , \9940 , \17511 );
or \U$9246 ( \18065 , \9930 , \17825 );
nand \U$9247 ( \18066 , \18064 , \18065 );
nor \U$9248 ( \18067 , \18063 , \18066 );
or \U$9249 ( \18068 , \13143 , \17540 );
or \U$9250 ( \18069 , \9937 , \17544 );
nand \U$9251 ( \18070 , \18068 , \18069 );
not \U$9252 ( \18071 , \17582 );
or \U$9253 ( \18072 , \9955 , \18071 );
not \U$9254 ( \18073 , \17617 );
or \U$9255 ( \18074 , \9948 , \18073 );
nand \U$9256 ( \18075 , \18072 , \18074 );
nor \U$9257 ( \18076 , \18070 , \18075 );
not \U$9258 ( \18077 , \17588 );
or \U$9259 ( \18078 , \12282 , \18077 );
not \U$9260 ( \18079 , \18039 );
or \U$9261 ( \18080 , \11633 , \18079 );
not \U$9262 ( \18081 , \17747 );
and \U$9263 ( \18082 , \9975 , \18081 );
not \U$9264 ( \18083 , \17519 );
and \U$9265 ( \18084 , \18083 , \9977 );
nor \U$9266 ( \18085 , \18082 , \18084 );
nand \U$9267 ( \18086 , \18078 , \18080 , \18085 );
not \U$9268 ( \18087 , \11623 );
and \U$9269 ( \18088 , \18087 , \18049 );
and \U$9270 ( \18089 , \17555 , \10709 );
nor \U$9271 ( \18090 , \18088 , \18089 );
not \U$9272 ( \18091 , \11620 );
and \U$9273 ( \18092 , \18091 , \17572 );
and \U$9274 ( \18093 , \17550 , \9968 );
nor \U$9275 ( \18094 , \18092 , \18093 );
nand \U$9276 ( \18095 , \18090 , \18094 );
nor \U$9277 ( \18096 , \18086 , \18095 );
nand \U$9278 ( \18097 , \18067 , \18076 , \18096 );
xnor \U$9279 ( \18098 , \18097 , \9990 );
nor \U$9280 ( \18099 , \18060 , \18098 );
nand \U$9281 ( \18100 , \17980 , \18019 , \18099 );
not \U$9282 ( \18101 , \18100 );
not \U$9283 ( \18102 , \17617 );
or \U$9284 ( \18103 , \9997 , \18102 );
not \U$9285 ( \18104 , \17674 );
or \U$9286 ( \18105 , \11666 , \18104 );
nand \U$9287 ( \18106 , \18103 , \18105 );
not \U$9288 ( \18107 , \17632 );
or \U$9289 ( \18108 , \10002 , \18107 );
not \U$9290 ( \18109 , \17582 );
or \U$9291 ( \18110 , \10005 , \18109 );
nand \U$9292 ( \18111 , \18108 , \18110 );
nor \U$9293 ( \18112 , \18106 , \18111 );
not \U$9294 ( \18113 , \10017 );
or \U$9295 ( \18114 , \18113 , \17544 );
or \U$9296 ( \18115 , \10013 , \17533 );
nand \U$9297 ( \18116 , \18114 , \18115 );
or \U$9298 ( \18117 , \10021 , \17597 );
or \U$9299 ( \18118 , \10010 , \17825 );
nand \U$9300 ( \18119 , \18117 , \18118 );
nor \U$9301 ( \18120 , \18116 , \18119 );
not \U$9302 ( \18121 , \18036 );
or \U$9303 ( \18122 , \11674 , \18121 );
not \U$9304 ( \18123 , \18039 );
or \U$9305 ( \18124 , \11681 , \18123 );
not \U$9306 ( \18125 , \17559 );
and \U$9307 ( \18126 , \10041 , \18125 );
not \U$9308 ( \18127 , \17928 );
and \U$9309 ( \18128 , \10043 , \18127 );
nor \U$9310 ( \18129 , \18126 , \18128 );
nand \U$9311 ( \18130 , \18122 , \18124 , \18129 );
not \U$9312 ( \18131 , \11693 );
and \U$9313 ( \18132 , \18131 , \18049 );
and \U$9314 ( \18133 , \17555 , \10027 );
nor \U$9315 ( \18134 , \18132 , \18133 );
not \U$9316 ( \18135 , \11698 );
and \U$9317 ( \18136 , \18135 , \17572 );
and \U$9318 ( \18137 , \17550 , \10035 );
nor \U$9319 ( \18138 , \18136 , \18137 );
nand \U$9320 ( \18139 , \18134 , \18138 );
nor \U$9321 ( \18140 , \18130 , \18139 );
nand \U$9322 ( \18141 , \18112 , \18120 , \18140 );
xnor \U$9323 ( \18142 , \18141 , \10055 );
or \U$9324 ( \18143 , \9878 , \17533 );
or \U$9325 ( \18144 , \9860 , \17536 );
nand \U$9326 ( \18145 , \18143 , \18144 );
or \U$9327 ( \18146 , \9887 , \17736 );
or \U$9328 ( \18147 , \9875 , \17825 );
nand \U$9329 ( \18148 , \18146 , \18147 );
nor \U$9330 ( \18149 , \18145 , \18148 );
or \U$9331 ( \18150 , \9868 , \17540 );
not \U$9332 ( \18151 , \17542 );
or \U$9333 ( \18152 , \10949 , \18151 );
or \U$9334 ( \18153 , \9884 , \18152 );
nand \U$9335 ( \18154 , \18150 , \18153 );
not \U$9336 ( \18155 , \17582 );
or \U$9337 ( \18156 , \12183 , \18155 );
not \U$9338 ( \18157 , \17617 );
or \U$9339 ( \18158 , \12178 , \18157 );
nand \U$9340 ( \18159 , \18156 , \18158 );
nor \U$9341 ( \18160 , \18154 , \18159 );
not \U$9342 ( \18161 , \18036 );
or \U$9343 ( \18162 , \9921 , \18161 );
not \U$9344 ( \18163 , \18039 );
or \U$9345 ( \18164 , \11718 , \18163 );
not \U$9346 ( \18165 , \17659 );
and \U$9347 ( \18166 , \18165 , \9913 );
not \U$9348 ( \18167 , \17519 );
and \U$9349 ( \18168 , \18167 , \9910 );
nor \U$9350 ( \18169 , \18166 , \18168 );
nand \U$9351 ( \18170 , \18162 , \18164 , \18169 );
not \U$9352 ( \18171 , \9906 );
and \U$9353 ( \18172 , \18171 , \18049 );
and \U$9354 ( \18173 , \17555 , \9902 );
nor \U$9355 ( \18174 , \18172 , \18173 );
not \U$9356 ( \18175 , \9898 );
and \U$9357 ( \18176 , \18175 , \17572 );
and \U$9358 ( \18177 , \17550 , \9892 );
nor \U$9359 ( \18178 , \18176 , \18177 );
nand \U$9360 ( \18179 , \18174 , \18178 );
nor \U$9361 ( \18180 , \18170 , \18179 );
nand \U$9362 ( \18181 , \18149 , \18160 , \18180 );
xnor \U$9363 ( \18182 , \18181 , \9927 );
nor \U$9364 ( \18183 , \18142 , \18182 );
not \U$9365 ( \18184 , \17617 );
or \U$9366 ( \18185 , \11494 , \18184 );
not \U$9367 ( \18186 , \17880 );
or \U$9368 ( \18187 , \9798 , \18186 );
nand \U$9369 ( \18188 , \18185 , \18187 );
not \U$9370 ( \18189 , \17632 );
or \U$9371 ( \18190 , \9791 , \18189 );
not \U$9372 ( \18191 , \17582 );
or \U$9373 ( \18192 , \11492 , \18191 );
nand \U$9374 ( \18193 , \18190 , \18192 );
nor \U$9375 ( \18194 , \18188 , \18193 );
not \U$9376 ( \18195 , \9813 );
or \U$9377 ( \18196 , \18195 , \18152 );
or \U$9378 ( \18197 , \9809 , \17601 );
nand \U$9379 ( \18198 , \18196 , \18197 );
or \U$9380 ( \18199 , \9817 , \17511 );
or \U$9381 ( \18200 , \9806 , \17825 );
nand \U$9382 ( \18201 , \18199 , \18200 );
nor \U$9383 ( \18202 , \18198 , \18201 );
not \U$9384 ( \18203 , \18036 );
or \U$9385 ( \18204 , \9851 , \18203 );
not \U$9386 ( \18205 , \18039 );
or \U$9387 ( \18206 , \11505 , \18205 );
not \U$9388 ( \18207 , \17747 );
and \U$9389 ( \18208 , \9842 , \18207 );
not \U$9390 ( \18209 , \17928 );
and \U$9391 ( \18210 , \9839 , \18209 );
nor \U$9392 ( \18211 , \18208 , \18210 );
nand \U$9393 ( \18212 , \18204 , \18206 , \18211 );
not \U$9394 ( \18213 , \9834 );
and \U$9395 ( \18214 , \18213 , \18049 );
and \U$9396 ( \18215 , \17555 , \9830 );
nor \U$9397 ( \18216 , \18214 , \18215 );
not \U$9398 ( \18217 , \9827 );
and \U$9399 ( \18218 , \18217 , \17572 );
and \U$9400 ( \18219 , \17550 , \9822 );
nor \U$9401 ( \18220 , \18218 , \18219 );
nand \U$9402 ( \18221 , \18216 , \18220 );
nor \U$9403 ( \18222 , \18212 , \18221 );
nand \U$9404 ( \18223 , \18194 , \18202 , \18222 );
xnor \U$9405 ( \18224 , \18223 , \9857 );
or \U$9406 ( \18225 , \9607 , \17601 );
or \U$9407 ( \18226 , \9588 , \17536 );
nand \U$9408 ( \18227 , \18225 , \18226 );
or \U$9409 ( \18228 , \9614 , \17597 );
or \U$9410 ( \18229 , \9604 , \17825 );
nand \U$9411 ( \18230 , \18228 , \18229 );
nor \U$9412 ( \18231 , \18227 , \18230 );
or \U$9413 ( \18232 , \9597 , \17540 );
or \U$9414 ( \18233 , \9611 , \17623 );
nand \U$9415 ( \18234 , \18232 , \18233 );
not \U$9416 ( \18235 , \17582 );
or \U$9417 ( \18236 , \12108 , \18235 );
not \U$9418 ( \18237 , \17617 );
or \U$9419 ( \18238 , \13538 , \18237 );
nand \U$9420 ( \18239 , \18236 , \18238 );
nor \U$9421 ( \18240 , \18234 , \18239 );
not \U$9422 ( \18241 , \18036 );
or \U$9423 ( \18242 , \9647 , \18241 );
not \U$9424 ( \18243 , \18039 );
or \U$9425 ( \18244 , \11322 , \18243 );
not \U$9426 ( \18245 , \17559 );
and \U$9427 ( \18246 , \9639 , \18245 );
not \U$9428 ( \18247 , \17519 );
and \U$9429 ( \18248 , \9636 , \18247 );
nor \U$9430 ( \18249 , \18246 , \18248 );
nand \U$9431 ( \18250 , \18242 , \18244 , \18249 );
not \U$9432 ( \18251 , \9632 );
and \U$9433 ( \18252 , \18251 , \18049 );
and \U$9434 ( \18253 , \17555 , \9628 );
nor \U$9435 ( \18254 , \18252 , \18253 );
not \U$9436 ( \18255 , \9625 );
and \U$9437 ( \18256 , \18255 , \17572 );
and \U$9438 ( \18257 , \17550 , \9619 );
nor \U$9439 ( \18258 , \18256 , \18257 );
nand \U$9440 ( \18259 , \18254 , \18258 );
nor \U$9441 ( \18260 , \18250 , \18259 );
nand \U$9442 ( \18261 , \18231 , \18240 , \18260 );
xnor \U$9443 ( \18262 , \18261 , \9653 );
nor \U$9444 ( \18263 , \18224 , \18262 );
and \U$9445 ( \18264 , \18101 , \18183 , \18263 );
nand \U$9446 ( \18265 , \17593 , \17936 , \18264 );
not \U$9447 ( \18266 , \18265 );
not \U$9448 ( \18267 , \18266 );
or \U$9449 ( \18268 , \17502 , \18267 );
not \U$9450 ( \18269 , \18268 );
not \U$9451 ( \18270 , \18266 );
or \U$9452 ( \18271 , \17501 , \18270 );
not \U$9453 ( \18272 , \18271 );
or \U$9454 ( \18273 , \18269 , \18272 );
or \U$9455 ( \18274 , \8906 , \18273 );
not \U$9456 ( \18275 , \10077 );
or \U$9457 ( \18276 , \8906 , \18275 );
not \U$9458 ( \18277 , \18276 );
nor \U$9459 ( \18278 , \13269 , \18277 );
not \U$9460 ( \18279 , \18278 );
not \U$9461 ( \18280 , \18271 );
and \U$9462 ( \18281 , \18279 , \18280 );
and \U$9463 ( \18282 , \18269 , \17508 );
nor \U$9464 ( \18283 , \18281 , \18282 );
nand \U$9465 ( \18284 , \18274 , \18283 );
not \U$9466 ( \18285 , \18284 );
and \U$9467 ( \18286 , \18285 , \17472 );
or \U$9468 ( \18287 , \17474 , \18286 );
not \U$9469 ( \18288 , \18287 );
and \U$9470 ( \18289 , \16695 , \18288 );
not \U$9471 ( \18290 , \18289 );
and \U$9472 ( \18291 , \16693 , \18290 );
not \U$9473 ( \18292 , \18291 );
and \U$9474 ( \18293 , \18292 , \16004 );
or \U$9475 ( \18294 , \16006 , \18293 );
not \U$9476 ( \18295 , \18294 );
and \U$9477 ( \18296 , \18295 , \15289 );
or \U$9478 ( \18297 , \15291 , \18296 );
not \U$9479 ( \18298 , \18297 );
and \U$9480 ( \18299 , \14682 , \18298 );
or \U$9481 ( \18300 , \14680 , \18299 );
not \U$9482 ( \18301 , \16882 );
and \U$9483 ( \18302 , \10120 , \18301 );
not \U$9484 ( \18303 , \16818 );
and \U$9485 ( \18304 , \13270 , \18303 );
nor \U$9486 ( \18305 , \18302 , \18304 );
not \U$9487 ( \18306 , \9504 );
and \U$9488 ( \18307 , \18306 , \16802 );
buf \U$9489 ( \18308 , \16786 );
and \U$9490 ( \18309 , \18308 , \14019 );
nor \U$9491 ( \18310 , \18307 , \18309 );
nand \U$9492 ( \18311 , \18305 , \18310 );
buf \U$9493 ( \18312 , \16781 );
not \U$9494 ( \18313 , \18312 );
or \U$9495 ( \18314 , \9498 , \18313 );
not \U$9496 ( \18315 , \16774 );
or \U$9497 ( \18316 , \9500 , \18315 );
not \U$9498 ( \18317 , \9492 );
and \U$9499 ( \18318 , \18317 , \16792 );
and \U$9500 ( \18319 , \16877 , \10062 );
nor \U$9501 ( \18320 , \18318 , \18319 );
nand \U$9502 ( \18321 , \18314 , \18316 , \18320 );
nor \U$9503 ( \18322 , \18311 , \18321 );
not \U$9504 ( \18323 , \16750 );
not \U$9505 ( \18324 , \18323 );
or \U$9506 ( \18325 , \9475 , \18324 );
not \U$9507 ( \18326 , \16737 );
or \U$9508 ( \18327 , \9471 , \18326 );
not \U$9509 ( \18328 , \17380 );
and \U$9510 ( \18329 , \10986 , \18328 );
not \U$9511 ( \18330 , \16840 );
and \U$9512 ( \18331 , \9468 , \18330 );
nor \U$9513 ( \18332 , \18329 , \18331 );
nand \U$9514 ( \18333 , \18325 , \18327 , \18332 );
or \U$9515 ( \18334 , \9482 , \16806 );
not \U$9516 ( \18335 , \16830 );
or \U$9517 ( \18336 , \9485 , \18335 );
not \U$9518 ( \18337 , \16813 );
or \U$9519 ( \18338 , \18337 , \9487 );
not \U$9520 ( \18339 , \16769 );
or \U$9521 ( \18340 , \9480 , \18339 );
and \U$9522 ( \18341 , \18334 , \18336 , \18338 , \18340 );
not \U$9523 ( \18342 , \18341 );
nor \U$9524 ( \18343 , \18333 , \18342 );
nand \U$9525 ( \18344 , \18322 , \18343 );
not \U$9526 ( \18345 , \18344 );
not \U$9527 ( \18346 , \13305 );
and \U$9528 ( \18347 , \18346 , \16813 );
not \U$9529 ( \18348 , \16818 );
and \U$9530 ( \18349 , \18348 , \9731 );
nor \U$9531 ( \18350 , \18347 , \18349 );
not \U$9532 ( \18351 , \9722 );
and \U$9533 ( \18352 , \18351 , \16830 );
and \U$9534 ( \18353 , \16877 , \9724 );
nor \U$9535 ( \18354 , \18352 , \18353 );
or \U$9536 ( \18355 , \9740 , \16840 );
not \U$9537 ( \18356 , \16762 );
or \U$9538 ( \18357 , \11876 , \18356 );
nand \U$9539 ( \18358 , \18355 , \18357 );
or \U$9540 ( \18359 , \9745 , \16736 );
or \U$9541 ( \18360 , \9748 , \16746 );
nand \U$9542 ( \18361 , \18359 , \18360 );
nor \U$9543 ( \18362 , \18358 , \18361 );
nand \U$9544 ( \18363 , \18350 , \18354 , \18362 );
not \U$9545 ( \18364 , \11186 );
and \U$9546 ( \18365 , \18364 , \16807 );
and \U$9547 ( \18366 , \16769 , \9779 );
nor \U$9548 ( \18367 , \18365 , \18366 );
not \U$9549 ( \18368 , \10182 );
and \U$9550 ( \18369 , \18368 , \18323 );
and \U$9551 ( \18370 , \16859 , \9772 );
nor \U$9552 ( \18371 , \18369 , \18370 );
not \U$9553 ( \18372 , \18312 );
or \U$9554 ( \18373 , \10194 , \18372 );
not \U$9555 ( \18374 , \18308 );
or \U$9556 ( \18375 , \10197 , \18374 );
nand \U$9557 ( \18376 , \18373 , \18375 );
not \U$9558 ( \18377 , \16792 );
or \U$9559 ( \18378 , \11193 , \18377 );
not \U$9560 ( \18379 , \16774 );
or \U$9561 ( \18380 , \11195 , \18379 );
nand \U$9562 ( \18381 , \18378 , \18380 );
nor \U$9563 ( \18382 , \18376 , \18381 );
nand \U$9564 ( \18383 , \18367 , \18371 , \18382 );
nor \U$9565 ( \18384 , \18363 , \18383 );
xnor \U$9566 ( \18385 , \18384 , \9786 );
not \U$9567 ( \18386 , \13344 );
and \U$9568 ( \18387 , \18386 , \17231 );
not \U$9569 ( \18388 , \16818 );
and \U$9570 ( \18389 , \18388 , \9667 );
nor \U$9571 ( \18390 , \18387 , \18389 );
not \U$9572 ( \18391 , \9658 );
and \U$9573 ( \18392 , \18391 , \16830 );
and \U$9574 ( \18393 , \16796 , \9660 );
nor \U$9575 ( \18394 , \18392 , \18393 );
or \U$9576 ( \18395 , \9676 , \16743 );
or \U$9577 ( \18396 , \11923 , \17219 );
nand \U$9578 ( \18397 , \18395 , \18396 );
or \U$9579 ( \18398 , \9680 , \16844 );
or \U$9580 ( \18399 , \9683 , \16882 );
nand \U$9581 ( \18400 , \18398 , \18399 );
nor \U$9582 ( \18401 , \18397 , \18400 );
nand \U$9583 ( \18402 , \18390 , \18394 , \18401 );
not \U$9584 ( \18403 , \11145 );
and \U$9585 ( \18404 , \18403 , \16807 );
and \U$9586 ( \18405 , \16769 , \9713 );
nor \U$9587 ( \18406 , \18404 , \18405 );
not \U$9588 ( \18407 , \11140 );
and \U$9589 ( \18408 , \18407 , \18323 );
and \U$9590 ( \18409 , \16859 , \9706 );
nor \U$9591 ( \18410 , \18408 , \18409 );
not \U$9592 ( \18411 , \18312 );
or \U$9593 ( \18412 , \10248 , \18411 );
not \U$9594 ( \18413 , \18308 );
or \U$9595 ( \18414 , \10250 , \18413 );
nand \U$9596 ( \18415 , \18412 , \18414 );
not \U$9597 ( \18416 , \16898 );
or \U$9598 ( \18417 , \11152 , \18416 );
not \U$9599 ( \18418 , \16774 );
or \U$9600 ( \18419 , \11154 , \18418 );
nand \U$9601 ( \18420 , \18417 , \18419 );
nor \U$9602 ( \18421 , \18415 , \18420 );
nand \U$9603 ( \18422 , \18406 , \18410 , \18421 );
nor \U$9604 ( \18423 , \18402 , \18422 );
xnor \U$9605 ( \18424 , \18423 , \9719 );
or \U$9606 ( \18425 , \11093 , \17036 );
not \U$9607 ( \18426 , \16877 );
or \U$9608 ( \18427 , \9226 , \18426 );
not \U$9609 ( \18428 , \16830 );
or \U$9610 ( \18429 , \9205 , \18428 );
not \U$9611 ( \18430 , \16813 );
or \U$9612 ( \18431 , \18430 , \9197 );
and \U$9613 ( \18432 , \18425 , \18427 , \18429 , \18431 );
not \U$9614 ( \18433 , \18432 );
not \U$9615 ( \18434 , \18312 );
or \U$9616 ( \18435 , \11117 , \18434 );
not \U$9617 ( \18436 , \18308 );
or \U$9618 ( \18437 , \11120 , \18436 );
not \U$9619 ( \18438 , \11111 );
and \U$9620 ( \18439 , \18438 , \16896 );
and \U$9621 ( \18440 , \16898 , \9230 );
nor \U$9622 ( \18441 , \18439 , \18440 );
nand \U$9623 ( \18442 , \18435 , \18437 , \18441 );
nor \U$9624 ( \18443 , \18433 , \18442 );
nand \U$9625 ( \18444 , \9216 , \16737 );
nand \U$9626 ( \18445 , \9219 , \17174 );
not \U$9627 ( \18446 , \17432 );
and \U$9628 ( \18447 , \9210 , \18446 );
not \U$9629 ( \18448 , \16840 );
and \U$9630 ( \18449 , \9212 , \18448 );
nor \U$9631 ( \18450 , \18447 , \18449 );
nand \U$9632 ( \18451 , \18444 , \18445 , \18450 );
nand \U$9633 ( \18452 , \9228 , \16856 );
nand \U$9634 ( \18453 , \9200 , \16859 );
and \U$9635 ( \18454 , \16769 , \9242 );
and \U$9636 ( \18455 , \9193 , \16807 );
nor \U$9637 ( \18456 , \18454 , \18455 );
nand \U$9638 ( \18457 , \18452 , \18453 , \18456 );
nor \U$9639 ( \18458 , \18451 , \18457 );
nand \U$9640 ( \18459 , \18443 , \18458 );
xnor \U$9641 ( \18460 , \18459 , \9260 );
or \U$9642 ( \18461 , \11036 , \17036 );
nand \U$9643 ( \18462 , \9006 , \16796 );
nand \U$9644 ( \18463 , \8976 , \16830 );
nand \U$9645 ( \18464 , \8966 , \17231 );
and \U$9646 ( \18465 , \18461 , \18462 , \18463 , \18464 );
not \U$9647 ( \18466 , \18465 );
nand \U$9648 ( \18467 , \9034 , \18312 );
nand \U$9649 ( \18468 , \9030 , \18308 );
and \U$9650 ( \18469 , \16792 , \9011 );
and \U$9651 ( \18470 , \9014 , \16774 );
nor \U$9652 ( \18471 , \18469 , \18470 );
nand \U$9653 ( \18472 , \18467 , \18468 , \18471 );
nor \U$9654 ( \18473 , \18466 , \18472 );
not \U$9655 ( \18474 , \16737 );
or \U$9656 ( \18475 , \8997 , \18474 );
not \U$9657 ( \18476 , \17174 );
or \U$9658 ( \18477 , \9000 , \18476 );
not \U$9659 ( \18478 , \17276 );
and \U$9660 ( \18479 , \8986 , \18478 );
not \U$9661 ( \18480 , \17179 );
and \U$9662 ( \18481 , \8990 , \18480 );
nor \U$9663 ( \18482 , \18479 , \18481 );
nand \U$9664 ( \18483 , \18475 , \18477 , \18482 );
not \U$9665 ( \18484 , \16856 );
or \U$9666 ( \18485 , \11073 , \18484 );
not \U$9667 ( \18486 , \16859 );
or \U$9668 ( \18487 , \8980 , \18486 );
not \U$9669 ( \18488 , \8971 );
and \U$9670 ( \18489 , \18488 , \16807 );
and \U$9671 ( \18490 , \16769 , \9025 );
nor \U$9672 ( \18491 , \18489 , \18490 );
nand \U$9673 ( \18492 , \18485 , \18487 , \18491 );
nor \U$9674 ( \18493 , \18483 , \18492 );
nand \U$9675 ( \18494 , \18473 , \18493 );
xnor \U$9676 ( \18495 , \18494 , \9044 );
nor \U$9677 ( \18496 , \18460 , \18495 );
nand \U$9678 ( \18497 , \18385 , \18424 , \18496 );
not \U$9679 ( \18498 , \18497 );
or \U$9680 ( \18499 , \11270 , \17036 );
not \U$9681 ( \18500 , \16796 );
or \U$9682 ( \18501 , \11303 , \18500 );
not \U$9683 ( \18502 , \16830 );
or \U$9684 ( \18503 , \9270 , \18502 );
not \U$9685 ( \18504 , \17231 );
or \U$9686 ( \18505 , \18504 , \9263 );
and \U$9687 ( \18506 , \18499 , \18501 , \18503 , \18505 );
not \U$9688 ( \18507 , \18506 );
not \U$9689 ( \18508 , \18312 );
or \U$9690 ( \18509 , \11291 , \18508 );
not \U$9691 ( \18510 , \18308 );
or \U$9692 ( \18511 , \11293 , \18510 );
not \U$9693 ( \18512 , \11286 );
and \U$9694 ( \18513 , \18512 , \16774 );
and \U$9695 ( \18514 , \16898 , \9299 );
nor \U$9696 ( \18515 , \18513 , \18514 );
nand \U$9697 ( \18516 , \18509 , \18511 , \18515 );
nor \U$9698 ( \18517 , \18507 , \18516 );
not \U$9699 ( \18518 , \16737 );
or \U$9700 ( \18519 , \9287 , \18518 );
not \U$9701 ( \18520 , \17174 );
or \U$9702 ( \18521 , \9290 , \18520 );
not \U$9703 ( \18522 , \17240 );
and \U$9704 ( \18523 , \18522 , \9277 );
not \U$9705 ( \18524 , \17179 );
and \U$9706 ( \18525 , \18524 , \9281 );
nor \U$9707 ( \18526 , \18523 , \18525 );
nand \U$9708 ( \18527 , \18519 , \18521 , \18526 );
nand \U$9709 ( \18528 , \9297 , \16856 );
nand \U$9710 ( \18529 , \9272 , \16802 );
and \U$9711 ( \18530 , \16769 , \9310 );
and \U$9712 ( \18531 , \9265 , \16807 );
nor \U$9713 ( \18532 , \18530 , \18531 );
nand \U$9714 ( \18533 , \18528 , \18529 , \18532 );
nor \U$9715 ( \18534 , \18527 , \18533 );
nand \U$9716 ( \18535 , \18517 , \18534 );
xnor \U$9717 ( \18536 , \18535 , \9327 );
or \U$9718 ( \18537 , \11230 , \17036 );
nand \U$9719 ( \18538 , \9427 , \16796 );
nand \U$9720 ( \18539 , \9401 , \16830 );
nand \U$9721 ( \18540 , \9394 , \16813 );
and \U$9722 ( \18541 , \18537 , \18538 , \18539 , \18540 );
not \U$9723 ( \18542 , \18541 );
nand \U$9724 ( \18543 , \9453 , \18312 );
nand \U$9725 ( \18544 , \9449 , \18308 );
and \U$9726 ( \18545 , \16898 , \9432 );
and \U$9727 ( \18546 , \9435 , \16896 );
nor \U$9728 ( \18547 , \18545 , \18546 );
nand \U$9729 ( \18548 , \18543 , \18544 , \18547 );
nor \U$9730 ( \18549 , \18542 , \18548 );
nand \U$9731 ( \18550 , \9418 , \16737 );
nand \U$9732 ( \18551 , \9421 , \17174 );
not \U$9733 ( \18552 , \18356 );
and \U$9734 ( \18553 , \9409 , \18552 );
not \U$9735 ( \18554 , \17179 );
and \U$9736 ( \18555 , \9414 , \18554 );
nor \U$9737 ( \18556 , \18553 , \18555 );
nand \U$9738 ( \18557 , \18550 , \18551 , \18556 );
nand \U$9739 ( \18558 , \9430 , \18323 );
nand \U$9740 ( \18559 , \9404 , \16802 );
and \U$9741 ( \18560 , \16769 , \9444 );
and \U$9742 ( \18561 , \9397 , \16807 );
nor \U$9743 ( \18562 , \18560 , \18561 );
nand \U$9744 ( \18563 , \18558 , \18559 , \18562 );
nor \U$9745 ( \18564 , \18557 , \18563 );
nand \U$9746 ( \18565 , \18549 , \18564 );
xnor \U$9747 ( \18566 , \18565 , \9460 );
nor \U$9748 ( \18567 , \18536 , \18566 );
or \U$9749 ( \18568 , \9647 , \17036 );
not \U$9750 ( \18569 , \16830 );
or \U$9751 ( \18570 , \9637 , \18569 );
not \U$9752 ( \18571 , \16877 );
or \U$9753 ( \18572 , \9640 , \18571 );
not \U$9754 ( \18573 , \17231 );
or \U$9755 ( \18574 , \18573 , \11322 );
and \U$9756 ( \18575 , \18568 , \18570 , \18572 , \18574 );
not \U$9757 ( \18576 , \18575 );
not \U$9758 ( \18577 , \18312 );
or \U$9759 ( \18578 , \9620 , \18577 );
not \U$9760 ( \18579 , \18308 );
or \U$9761 ( \18580 , \9625 , \18579 );
and \U$9762 ( \18581 , \16774 , \9628 );
and \U$9763 ( \18582 , \16898 , \9631 );
nor \U$9764 ( \18583 , \18581 , \18582 );
nand \U$9765 ( \18584 , \18578 , \18580 , \18583 );
nor \U$9766 ( \18585 , \18576 , \18584 );
not \U$9767 ( \18586 , \16737 );
or \U$9768 ( \18587 , \9588 , \18586 );
not \U$9769 ( \18588 , \17174 );
or \U$9770 ( \18589 , \12108 , \18588 );
not \U$9771 ( \18590 , \18356 );
and \U$9772 ( \18591 , \18590 , \9596 );
not \U$9773 ( \18592 , \17179 );
and \U$9774 ( \18593 , \9600 , \18592 );
nor \U$9775 ( \18594 , \18591 , \18593 );
nand \U$9776 ( \18595 , \18587 , \18589 , \18594 );
or \U$9777 ( \18596 , \9604 , \16801 );
not \U$9778 ( \18597 , \16769 );
or \U$9779 ( \18598 , \9611 , \18597 );
not \U$9780 ( \18599 , \16987 );
or \U$9781 ( \18600 , \9614 , \18599 );
not \U$9782 ( \18601 , \16856 );
or \U$9783 ( \18602 , \9607 , \18601 );
and \U$9784 ( \18603 , \18596 , \18598 , \18600 , \18602 );
not \U$9785 ( \18604 , \18603 );
nor \U$9786 ( \18605 , \18595 , \18604 );
nand \U$9787 ( \18606 , \18585 , \18605 );
xnor \U$9788 ( \18607 , \18606 , \9653 );
or \U$9789 ( \18608 , \11393 , \17036 );
not \U$9790 ( \18609 , \16877 );
or \U$9791 ( \18610 , \11352 , \18609 );
not \U$9792 ( \18611 , \16830 );
or \U$9793 ( \18612 , \9339 , \18611 );
not \U$9794 ( \18613 , \16813 );
or \U$9795 ( \18614 , \18613 , \9332 );
and \U$9796 ( \18615 , \18608 , \18610 , \18612 , \18614 );
not \U$9797 ( \18616 , \18615 );
not \U$9798 ( \18617 , \18308 );
or \U$9799 ( \18618 , \12874 , \18617 );
not \U$9800 ( \18619 , \18312 );
or \U$9801 ( \18620 , \11371 , \18619 );
not \U$9802 ( \18621 , \13593 );
and \U$9803 ( \18622 , \18621 , \16896 );
and \U$9804 ( \18623 , \16792 , \9366 );
nor \U$9805 ( \18624 , \18622 , \18623 );
nand \U$9806 ( \18625 , \18618 , \18620 , \18624 );
nor \U$9807 ( \18626 , \18616 , \18625 );
not \U$9808 ( \18627 , \16737 );
or \U$9809 ( \18628 , \9354 , \18627 );
not \U$9810 ( \18629 , \17174 );
or \U$9811 ( \18630 , \9357 , \18629 );
not \U$9812 ( \18631 , \18356 );
and \U$9813 ( \18632 , \18631 , \9346 );
not \U$9814 ( \18633 , \17179 );
and \U$9815 ( \18634 , \18633 , \9348 );
nor \U$9816 ( \18635 , \18632 , \18634 );
nand \U$9817 ( \18636 , \18628 , \18630 , \18635 );
not \U$9818 ( \18637 , \16856 );
or \U$9819 ( \18638 , \11357 , \18637 );
not \U$9820 ( \18639 , \16802 );
or \U$9821 ( \18640 , \9342 , \18639 );
not \U$9822 ( \18641 , \9335 );
and \U$9823 ( \18642 , \18641 , \16807 );
and \U$9824 ( \18643 , \16769 , \9380 );
nor \U$9825 ( \18644 , \18642 , \18643 );
nand \U$9826 ( \18645 , \18638 , \18640 , \18644 );
nor \U$9827 ( \18646 , \18636 , \18645 );
nand \U$9828 ( \18647 , \18626 , \18646 );
xnor \U$9829 ( \18648 , \18647 , \9392 );
nor \U$9830 ( \18649 , \18607 , \18648 );
and \U$9831 ( \18650 , \18498 , \18567 , \18649 );
not \U$9832 ( \18651 , \9887 );
and \U$9833 ( \18652 , \18651 , \16807 );
and \U$9834 ( \18653 , \16769 , \9881 );
nor \U$9835 ( \18654 , \18652 , \18653 );
not \U$9836 ( \18655 , \9878 );
and \U$9837 ( \18656 , \18655 , \16856 );
and \U$9838 ( \18657 , \16859 , \9874 );
nor \U$9839 ( \18658 , \18656 , \18657 );
or \U$9840 ( \18659 , \12178 , \16743 );
or \U$9841 ( \18660 , \9868 , \16965 );
nand \U$9842 ( \18661 , \18659 , \18660 );
or \U$9843 ( \18662 , \9860 , \16844 );
or \U$9844 ( \18663 , \12183 , \16746 );
nand \U$9845 ( \18664 , \18662 , \18663 );
nor \U$9846 ( \18665 , \18661 , \18664 );
nand \U$9847 ( \18666 , \18654 , \18658 , \18665 );
or \U$9848 ( \18667 , \9895 , \16780 );
not \U$9849 ( \18668 , \18308 );
or \U$9850 ( \18669 , \9898 , \18668 );
nand \U$9851 ( \18670 , \18667 , \18669 );
not \U$9852 ( \18671 , \16792 );
or \U$9853 ( \18672 , \9906 , \18671 );
not \U$9854 ( \18673 , \16896 );
or \U$9855 ( \18674 , \11711 , \18673 );
nand \U$9856 ( \18675 , \18672 , \18674 );
nor \U$9857 ( \18676 , \18670 , \18675 );
not \U$9858 ( \18677 , \16813 );
or \U$9859 ( \18678 , \18677 , \11718 );
or \U$9860 ( \18679 , \9921 , \16954 );
nand \U$9861 ( \18680 , \18678 , \18679 );
not \U$9862 ( \18681 , \18680 );
not \U$9863 ( \18682 , \16877 );
or \U$9864 ( \18683 , \9914 , \18682 );
not \U$9865 ( \18684 , \16830 );
or \U$9866 ( \18685 , \9911 , \18684 );
and \U$9867 ( \18686 , \18681 , \18683 , \18685 );
nand \U$9868 ( \18687 , \18676 , \18686 );
nor \U$9869 ( \18688 , \18666 , \18687 );
xnor \U$9870 ( \18689 , \18688 , \9927 );
not \U$9871 ( \18690 , \10021 );
and \U$9872 ( \18691 , \18690 , \16807 );
and \U$9873 ( \18692 , \16769 , \10017 );
nor \U$9874 ( \18693 , \18691 , \18692 );
not \U$9875 ( \18694 , \10013 );
and \U$9876 ( \18695 , \18694 , \16856 );
and \U$9877 ( \18696 , \16859 , \10009 );
nor \U$9878 ( \18697 , \18695 , \18696 );
or \U$9879 ( \18698 , \9997 , \16743 );
or \U$9880 ( \18699 , \11666 , \16926 );
nand \U$9881 ( \18700 , \18698 , \18699 );
or \U$9882 ( \18701 , \10002 , \16970 );
or \U$9883 ( \18702 , \10005 , \16882 );
nand \U$9884 ( \18703 , \18701 , \18702 );
nor \U$9885 ( \18704 , \18700 , \18703 );
nand \U$9886 ( \18705 , \18693 , \18697 , \18704 );
not \U$9887 ( \18706 , \18312 );
or \U$9888 ( \18707 , \12230 , \18706 );
not \U$9889 ( \18708 , \18308 );
or \U$9890 ( \18709 , \11698 , \18708 );
nand \U$9891 ( \18710 , \18707 , \18709 );
not \U$9892 ( \18711 , \16792 );
or \U$9893 ( \18712 , \11693 , \18711 );
not \U$9894 ( \18713 , \16774 );
or \U$9895 ( \18714 , \12235 , \18713 );
nand \U$9896 ( \18715 , \18712 , \18714 );
nor \U$9897 ( \18716 , \18710 , \18715 );
not \U$9898 ( \18717 , \17231 );
or \U$9899 ( \18718 , \18717 , \11681 );
or \U$9900 ( \18719 , \11674 , \17036 );
nand \U$9901 ( \18720 , \18718 , \18719 );
not \U$9902 ( \18721 , \18720 );
not \U$9903 ( \18722 , \16796 );
or \U$9904 ( \18723 , \12222 , \18722 );
not \U$9905 ( \18724 , \16830 );
or \U$9906 ( \18725 , \11684 , \18724 );
and \U$9907 ( \18726 , \18721 , \18723 , \18725 );
nand \U$9908 ( \18727 , \18716 , \18726 );
nor \U$9909 ( \18728 , \18705 , \18727 );
xnor \U$9910 ( \18729 , \18728 , \10055 );
or \U$9911 ( \18730 , \9579 , \17036 );
not \U$9912 ( \18731 , \16830 );
or \U$9913 ( \18732 , \9569 , \18731 );
not \U$9914 ( \18733 , \16796 );
or \U$9915 ( \18734 , \9572 , \18733 );
not \U$9916 ( \18735 , \17231 );
or \U$9917 ( \18736 , \11589 , \18735 );
and \U$9918 ( \18737 , \18730 , \18732 , \18734 , \18736 );
not \U$9919 ( \18738 , \18737 );
not \U$9920 ( \18739 , \18312 );
or \U$9921 ( \18740 , \9552 , \18739 );
not \U$9922 ( \18741 , \18308 );
or \U$9923 ( \18742 , \9557 , \18741 );
and \U$9924 ( \18743 , \16774 , \9560 );
and \U$9925 ( \18744 , \16792 , \9563 );
nor \U$9926 ( \18745 , \18743 , \18744 );
nand \U$9927 ( \18746 , \18740 , \18742 , \18745 );
nor \U$9928 ( \18747 , \18738 , \18746 );
not \U$9929 ( \18748 , \16737 );
or \U$9930 ( \18749 , \9519 , \18748 );
not \U$9931 ( \18750 , \17174 );
or \U$9932 ( \18751 , \14434 , \18750 );
not \U$9933 ( \18752 , \18356 );
and \U$9934 ( \18753 , \9526 , \18752 );
not \U$9935 ( \18754 , \17179 );
and \U$9936 ( \18755 , \9530 , \18754 );
nor \U$9937 ( \18756 , \18753 , \18755 );
nand \U$9938 ( \18757 , \18749 , \18751 , \18756 );
or \U$9939 ( \18758 , \9534 , \16801 );
not \U$9940 ( \18759 , \16769 );
or \U$9941 ( \18760 , \9543 , \18759 );
not \U$9942 ( \18761 , \16987 );
or \U$9943 ( \18762 , \9546 , \18761 );
not \U$9944 ( \18763 , \16856 );
or \U$9945 ( \18764 , \9537 , \18763 );
and \U$9946 ( \18765 , \18758 , \18760 , \18762 , \18764 );
not \U$9947 ( \18766 , \18765 );
nor \U$9948 ( \18767 , \18757 , \18766 );
nand \U$9949 ( \18768 , \18747 , \18767 );
xnor \U$9950 ( \18769 , \18768 , \9585 );
or \U$9951 ( \18770 , \12282 , \17036 );
not \U$9952 ( \18771 , \16830 );
or \U$9953 ( \18772 , \11635 , \18771 );
not \U$9954 ( \18773 , \16796 );
or \U$9955 ( \18774 , \11629 , \18773 );
not \U$9956 ( \18775 , \16813 );
or \U$9957 ( \18776 , \11633 , \18775 );
and \U$9958 ( \18777 , \18770 , \18772 , \18774 , \18776 );
not \U$9959 ( \18778 , \18777 );
nand \U$9960 ( \18779 , \9968 , \18312 );
nand \U$9961 ( \18780 , \9965 , \18308 );
and \U$9962 ( \18781 , \16896 , \10709 );
and \U$9963 ( \18782 , \16792 , \9959 );
nor \U$9964 ( \18783 , \18781 , \18782 );
nand \U$9965 ( \18784 , \18779 , \18780 , \18783 );
nor \U$9966 ( \18785 , \18778 , \18784 );
nand \U$9967 ( \18786 , \9951 , \16737 );
nand \U$9968 ( \18787 , \9954 , \17174 );
not \U$9969 ( \18788 , \18356 );
and \U$9970 ( \18789 , \9944 , \18788 );
not \U$9971 ( \18790 , \17179 );
and \U$9972 ( \18791 , \9947 , \18790 );
nor \U$9973 ( \18792 , \18789 , \18791 );
nand \U$9974 ( \18793 , \18786 , \18787 , \18792 );
or \U$9975 ( \18794 , \9930 , \16801 );
nand \U$9976 ( \18795 , \9936 , \16769 );
nand \U$9977 ( \18796 , \9939 , \16987 );
nand \U$9978 ( \18797 , \9932 , \16856 );
and \U$9979 ( \18798 , \18794 , \18795 , \18796 , \18797 );
not \U$9980 ( \18799 , \18798 );
nor \U$9981 ( \18800 , \18793 , \18799 );
nand \U$9982 ( \18801 , \18785 , \18800 );
xnor \U$9983 ( \18802 , \18801 , \9990 );
nor \U$9984 ( \18803 , \18769 , \18802 );
nand \U$9985 ( \18804 , \18689 , \18729 , \18803 );
not \U$9986 ( \18805 , \8861 );
and \U$9987 ( \18806 , \18805 , \16802 );
and \U$9988 ( \18807 , \18323 , \8915 );
nor \U$9989 ( \18808 , \18806 , \18807 );
not \U$9990 ( \18809 , \8844 );
and \U$9991 ( \18810 , \18809 , \16807 );
and \U$9992 ( \18811 , \16769 , \8940 );
nor \U$9993 ( \18812 , \18810 , \18811 );
or \U$9994 ( \18813 , \8882 , \16743 );
or \U$9995 ( \18814 , \12351 , \16838 );
nand \U$9996 ( \18815 , \18813 , \18814 );
or \U$9997 ( \18816 , \8894 , \16970 );
or \U$9998 ( \18817 , \8897 , \16746 );
nand \U$9999 ( \18818 , \18816 , \18817 );
nor \U$10000 ( \18819 , \18815 , \18818 );
nand \U$10001 ( \18820 , \18808 , \18812 , \18819 );
nand \U$10002 ( \18821 , \8927 , \16896 );
nand \U$10003 ( \18822 , \8921 , \16898 );
nand \U$10004 ( \18823 , \18821 , \18822 );
nand \U$10005 ( \18824 , \8953 , \18312 );
nand \U$10006 ( \18825 , \8947 , \18308 );
nand \U$10007 ( \18826 , \18824 , \18825 );
nor \U$10008 ( \18827 , \18823 , \18826 );
or \U$10009 ( \18828 , \8828 , \16812 );
or \U$10010 ( \18829 , \11565 , \16954 );
nand \U$10011 ( \18830 , \18828 , \18829 );
not \U$10012 ( \18831 , \18830 );
not \U$10013 ( \18832 , \16830 );
or \U$10014 ( \18833 , \8853 , \18832 );
not \U$10015 ( \18834 , \16877 );
or \U$10016 ( \18835 , \11528 , \18834 );
and \U$10017 ( \18836 , \18831 , \18833 , \18835 );
nand \U$10018 ( \18837 , \18827 , \18836 );
nor \U$10019 ( \18838 , \18820 , \18837 );
xnor \U$10020 ( \18839 , \18838 , \8964 );
not \U$10021 ( \18840 , \9817 );
and \U$10022 ( \18841 , \18840 , \16987 );
and \U$10023 ( \18842 , \16769 , \9813 );
nor \U$10024 ( \18843 , \18841 , \18842 );
not \U$10025 ( \18844 , \9809 );
and \U$10026 ( \18845 , \18844 , \18323 );
and \U$10027 ( \18846 , \16859 , \9805 );
nor \U$10028 ( \18847 , \18845 , \18846 );
or \U$10029 ( \18848 , \11494 , \16743 );
or \U$10030 ( \18849 , \9798 , \16885 );
nand \U$10031 ( \18850 , \18848 , \18849 );
or \U$10032 ( \18851 , \9791 , \16736 );
or \U$10033 ( \18852 , \11492 , \16882 );
nand \U$10034 ( \18853 , \18851 , \18852 );
nor \U$10035 ( \18854 , \18850 , \18853 );
nand \U$10036 ( \18855 , \18843 , \18847 , \18854 );
nand \U$10037 ( \18856 , \9822 , \18312 );
nand \U$10038 ( \18857 , \9826 , \18308 );
nand \U$10039 ( \18858 , \18856 , \18857 );
nand \U$10040 ( \18859 , \9833 , \16898 );
nand \U$10041 ( \18860 , \9830 , \16896 );
nand \U$10042 ( \18861 , \18859 , \18860 );
nor \U$10043 ( \18862 , \18858 , \18861 );
not \U$10044 ( \18863 , \17231 );
or \U$10045 ( \18864 , \18863 , \11505 );
or \U$10046 ( \18865 , \9851 , \17036 );
nand \U$10047 ( \18866 , \18864 , \18865 );
not \U$10048 ( \18867 , \18866 );
not \U$10049 ( \18868 , \16796 );
or \U$10050 ( \18869 , \9843 , \18868 );
not \U$10051 ( \18870 , \16830 );
or \U$10052 ( \18871 , \9840 , \18870 );
and \U$10053 ( \18872 , \18867 , \18869 , \18871 );
nand \U$10054 ( \18873 , \18862 , \18872 );
nor \U$10055 ( \18874 , \18855 , \18873 );
xnor \U$10056 ( \18875 , \18874 , \9857 );
or \U$10057 ( \18876 , \11452 , \16954 );
nand \U$10058 ( \18877 , \9081 , \16877 );
nand \U$10059 ( \18878 , \9054 , \16830 );
nand \U$10060 ( \18879 , \9046 , \16813 );
and \U$10061 ( \18880 , \18876 , \18877 , \18878 , \18879 );
not \U$10062 ( \18881 , \18880 );
nand \U$10063 ( \18882 , \9112 , \18312 );
nand \U$10064 ( \18883 , \9107 , \18308 );
and \U$10065 ( \18884 , \16898 , \9089 );
and \U$10066 ( \18885 , \9093 , \16896 );
nor \U$10067 ( \18886 , \18884 , \18885 );
nand \U$10068 ( \18887 , \18882 , \18883 , \18886 );
nor \U$10069 ( \18888 , \18881 , \18887 );
nand \U$10070 ( \18889 , \9072 , \16737 );
nand \U$10071 ( \18890 , \9075 , \17174 );
not \U$10072 ( \18891 , \17085 );
and \U$10073 ( \18892 , \9063 , \18891 );
not \U$10074 ( \18893 , \16743 );
and \U$10075 ( \18894 , \9067 , \18893 );
nor \U$10076 ( \18895 , \18892 , \18894 );
nand \U$10077 ( \18896 , \18889 , \18890 , \18895 );
nand \U$10078 ( \18897 , \9085 , \16856 );
nand \U$10079 ( \18898 , \9057 , \16859 );
and \U$10080 ( \18899 , \16769 , \9102 );
and \U$10081 ( \18900 , \9049 , \16807 );
nor \U$10082 ( \18901 , \18899 , \18900 );
nand \U$10083 ( \18902 , \18897 , \18898 , \18901 );
nor \U$10084 ( \18903 , \18896 , \18902 );
nand \U$10085 ( \18904 , \18888 , \18903 );
xnor \U$10086 ( \18905 , \18904 , \9119 );
or \U$10087 ( \18906 , \11410 , \16954 );
nand \U$10088 ( \18907 , \9155 , \16877 );
nand \U$10089 ( \18908 , \9129 , \16830 );
nand \U$10090 ( \18909 , \9121 , \17231 );
and \U$10091 ( \18910 , \18906 , \18907 , \18908 , \18909 );
not \U$10092 ( \18911 , \18910 );
nand \U$10093 ( \18912 , \9180 , \18312 );
nand \U$10094 ( \18913 , \9176 , \18308 );
and \U$10095 ( \18914 , \16898 , \9159 );
and \U$10096 ( \18915 , \9163 , \16896 );
nor \U$10097 ( \18916 , \18914 , \18915 );
nand \U$10098 ( \18917 , \18912 , \18913 , \18916 );
nor \U$10099 ( \18918 , \18911 , \18917 );
nand \U$10100 ( \18919 , \9147 , \16737 );
nand \U$10101 ( \18920 , \9150 , \17174 );
not \U$10102 ( \18921 , \18356 );
and \U$10103 ( \18922 , \9137 , \18921 );
not \U$10104 ( \18923 , \17179 );
and \U$10105 ( \18924 , \9142 , \18923 );
nor \U$10106 ( \18925 , \18922 , \18924 );
nand \U$10107 ( \18926 , \18919 , \18920 , \18925 );
nand \U$10108 ( \18927 , \9157 , \16856 );
nand \U$10109 ( \18928 , \9132 , \16802 );
and \U$10110 ( \18929 , \16769 , \9172 );
and \U$10111 ( \18930 , \9124 , \16807 );
nor \U$10112 ( \18931 , \18929 , \18930 );
nand \U$10113 ( \18932 , \18927 , \18928 , \18931 );
nor \U$10114 ( \18933 , \18926 , \18932 );
nand \U$10115 ( \18934 , \18918 , \18933 );
xnor \U$10116 ( \18935 , \18934 , \9188 );
nor \U$10117 ( \18936 , \18905 , \18935 );
nand \U$10118 ( \18937 , \18839 , \18875 , \18936 );
nor \U$10119 ( \18938 , \18804 , \18937 );
nand \U$10120 ( \18939 , \18345 , \18650 , \18938 );
not \U$10121 ( \18940 , \18939 );
or \U$10122 ( \18941 , \9492 , \17536 );
or \U$10123 ( \18942 , \9494 , \17533 );
nand \U$10124 ( \18943 , \18941 , \18942 );
not \U$10125 ( \18944 , \17617 );
not \U$10126 ( \18945 , \18944 );
not \U$10127 ( \18946 , \18945 );
or \U$10128 ( \18947 , \9498 , \18946 );
not \U$10129 ( \18948 , \17584 );
or \U$10130 ( \18949 , \9500 , \18948 );
nand \U$10131 ( \18950 , \18947 , \18949 );
nor \U$10132 ( \18951 , \18943 , \18950 );
or \U$10133 ( \18952 , \9506 , \17540 );
or \U$10134 ( \18953 , \9485 , \17603 );
nand \U$10135 ( \18954 , \18952 , \18953 );
or \U$10136 ( \18955 , \9511 , \17554 );
or \U$10137 ( \18956 , \9504 , \17928 );
nand \U$10138 ( \18957 , \18955 , \18956 );
nor \U$10139 ( \18958 , \18954 , \18957 );
not \U$10140 ( \18959 , \17572 );
or \U$10141 ( \18960 , \9463 , \18959 );
not \U$10142 ( \18961 , \17624 );
or \U$10143 ( \18962 , \9509 , \18961 );
not \U$10144 ( \18963 , \17744 );
and \U$10145 ( \18964 , \9472 , \18963 );
not \U$10146 ( \18965 , \17747 );
and \U$10147 ( \18966 , \9476 , \18965 );
nor \U$10148 ( \18967 , \18964 , \18966 );
nand \U$10149 ( \18968 , \18960 , \18962 , \18967 );
not \U$10150 ( \18969 , \9487 );
and \U$10151 ( \18970 , \18969 , \17946 );
and \U$10152 ( \18971 , \17588 , \10152 );
nor \U$10153 ( \18972 , \18970 , \18971 );
not \U$10154 ( \18973 , \9482 );
and \U$10155 ( \18974 , \18973 , \18039 );
and \U$10156 ( \18975 , \17550 , \9468 );
nor \U$10157 ( \18976 , \18974 , \18975 );
nand \U$10158 ( \18977 , \18972 , \18976 );
nor \U$10159 ( \18978 , \18968 , \18977 );
nand \U$10160 ( \18979 , \18951 , \18958 , \18978 );
not \U$10161 ( \18980 , \18979 );
not \U$10162 ( \18981 , \9740 );
and \U$10163 ( \18982 , \18981 , \17550 );
and \U$10164 ( \18983 , \17555 , \9747 );
nor \U$10165 ( \18984 , \18982 , \18983 );
not \U$10166 ( \18985 , \9732 );
and \U$10167 ( \18986 , \18985 , \17624 );
and \U$10168 ( \18987 , \17572 , \9736 );
nor \U$10169 ( \18988 , \18986 , \18987 );
or \U$10170 ( \18989 , \9725 , \17601 );
or \U$10171 ( \18990 , \9745 , \17656 );
nand \U$10172 ( \18991 , \18989 , \18990 );
or \U$10173 ( \18992 , \13305 , \17597 );
or \U$10174 ( \18993 , \9722 , \17603 );
nand \U$10175 ( \18994 , \18992 , \18993 );
nor \U$10176 ( \18995 , \18991 , \18994 );
nand \U$10177 ( \18996 , \18984 , \18988 , \18995 );
or \U$10178 ( \18997 , \10178 , \17519 );
or \U$10179 ( \18998 , \10182 , \17659 );
nand \U$10180 ( \18999 , \18997 , \18998 );
or \U$10181 ( \19000 , \10188 , \17587 );
or \U$10182 ( \19001 , \11186 , \17771 );
nand \U$10183 ( \19002 , \19000 , \19001 );
nor \U$10184 ( \19003 , \18999 , \19002 );
not \U$10185 ( \19004 , \18945 );
or \U$10186 ( \19005 , \10194 , \19004 );
not \U$10187 ( \19006 , \17674 );
or \U$10188 ( \19007 , \10197 , \19006 );
nand \U$10189 ( \19008 , \19005 , \19007 );
not \U$10190 ( \19009 , \17632 );
or \U$10191 ( \19010 , \19009 , \11193 );
not \U$10192 ( \19011 , \17584 );
or \U$10193 ( \19012 , \11195 , \19011 );
nand \U$10194 ( \19013 , \19010 , \19012 );
nor \U$10195 ( \19014 , \19008 , \19013 );
nand \U$10196 ( \19015 , \19003 , \19014 );
nor \U$10197 ( \19016 , \18996 , \19015 );
xnor \U$10198 ( \19017 , \19016 , \9786 );
not \U$10199 ( \19018 , \9680 );
and \U$10200 ( \19019 , \19018 , \18049 );
and \U$10201 ( \19020 , \17555 , \9682 );
nor \U$10202 ( \19021 , \19019 , \19020 );
not \U$10203 ( \19022 , \11923 );
and \U$10204 ( \19023 , \19022 , \17572 );
and \U$10205 ( \19024 , \17550 , \9675 );
nor \U$10206 ( \19025 , \19023 , \19024 );
or \U$10207 ( \19026 , \9658 , \17603 );
or \U$10208 ( \19027 , \9661 , \17533 );
nand \U$10209 ( \19028 , \19026 , \19027 );
or \U$10210 ( \19029 , \9668 , \18152 );
or \U$10211 ( \19030 , \13344 , \17511 );
nand \U$10212 ( \19031 , \19029 , \19030 );
nor \U$10213 ( \19032 , \19028 , \19031 );
nand \U$10214 ( \19033 , \19021 , \19025 , \19032 );
or \U$10215 ( \19034 , \11138 , \17638 );
or \U$10216 ( \19035 , \11140 , \17747 );
nand \U$10217 ( \19036 , \19034 , \19035 );
or \U$10218 ( \19037 , \10244 , \17587 );
or \U$10219 ( \19038 , \11145 , \17685 );
nand \U$10220 ( \19039 , \19037 , \19038 );
nor \U$10221 ( \19040 , \19036 , \19039 );
not \U$10222 ( \19041 , \18945 );
or \U$10223 ( \19042 , \10248 , \19041 );
not \U$10224 ( \19043 , \17626 );
or \U$10225 ( \19044 , \10250 , \19043 );
nand \U$10226 ( \19045 , \19042 , \19044 );
not \U$10227 ( \19046 , \17632 );
or \U$10228 ( \19047 , \19046 , \11152 );
not \U$10229 ( \19048 , \17584 );
or \U$10230 ( \19049 , \11154 , \19048 );
nand \U$10231 ( \19050 , \19047 , \19049 );
nor \U$10232 ( \19051 , \19045 , \19050 );
nand \U$10233 ( \19052 , \19040 , \19051 );
nor \U$10234 ( \19053 , \19033 , \19052 );
xnor \U$10235 ( \19054 , \19053 , \9719 );
not \U$10236 ( \19055 , \9217 );
not \U$10237 ( \19056 , \17656 );
and \U$10238 ( \19057 , \19055 , \19056 );
or \U$10239 ( \19058 , \11954 , \17638 );
or \U$10240 ( \19059 , \11088 , \17522 );
nand \U$10241 ( \19060 , \19058 , \19059 );
not \U$10242 ( \19061 , \17587 );
and \U$10243 ( \19062 , \19061 , \9242 );
or \U$10244 ( \19063 , \19057 , \19060 , \19062 );
not \U$10245 ( \19064 , \19063 );
or \U$10246 ( \19065 , \11101 , \17571 );
or \U$10247 ( \19066 , \11093 , \17623 );
nand \U$10248 ( \19067 , \19065 , \19066 );
or \U$10249 ( \19068 , \9220 , \17554 );
or \U$10250 ( \19069 , \11098 , \17549 );
nand \U$10251 ( \19070 , \19068 , \19069 );
nor \U$10252 ( \19071 , \19067 , \19070 );
not \U$10253 ( \19072 , \18006 );
or \U$10254 ( \19073 , \9226 , \19072 );
not \U$10255 ( \19074 , \17576 );
or \U$10256 ( \19075 , \9205 , \19074 );
not \U$10257 ( \19076 , \17559 );
and \U$10258 ( \19077 , \19076 , \9228 );
not \U$10259 ( \19078 , \17511 );
and \U$10260 ( \19079 , \9196 , \19078 );
nor \U$10261 ( \19080 , \19077 , \19079 );
nand \U$10262 ( \19081 , \19073 , \19075 , \19080 );
not \U$10263 ( \19082 , \11120 );
and \U$10264 ( \19083 , \19082 , \17880 );
and \U$10265 ( \19084 , \18945 , \9251 );
nor \U$10266 ( \19085 , \19083 , \19084 );
not \U$10267 ( \19086 , \11113 );
and \U$10268 ( \19087 , \19086 , \17680 );
and \U$10269 ( \19088 , \17584 , \9233 );
nor \U$10270 ( \19089 , \19087 , \19088 );
nand \U$10271 ( \19090 , \19085 , \19089 );
nor \U$10272 ( \19091 , \19081 , \19090 );
nand \U$10273 ( \19092 , \19064 , \19071 , \19091 );
xnor \U$10274 ( \19093 , \19092 , \9260 );
not \U$10275 ( \19094 , \8997 );
not \U$10276 ( \19095 , \17563 );
and \U$10277 ( \19096 , \19094 , \19095 );
or \U$10278 ( \19097 , \8980 , \17638 );
or \U$10279 ( \19098 , \8971 , \17685 );
nand \U$10280 ( \19099 , \19097 , \19098 );
not \U$10281 ( \19100 , \17587 );
and \U$10282 ( \19101 , \19100 , \9025 );
or \U$10283 ( \19102 , \19096 , \19099 , \19101 );
not \U$10284 ( \19103 , \19102 );
or \U$10285 ( \19104 , \11046 , \17733 );
or \U$10286 ( \19105 , \11036 , \17544 );
nand \U$10287 ( \19106 , \19104 , \19105 );
or \U$10288 ( \19107 , \9000 , \17612 );
or \U$10289 ( \19108 , \8991 , \17751 );
nand \U$10290 ( \19109 , \19107 , \19108 );
nor \U$10291 ( \19110 , \19106 , \19109 );
not \U$10292 ( \19111 , \18006 );
or \U$10293 ( \19112 , \11080 , \19111 );
not \U$10294 ( \19113 , \17576 );
or \U$10295 ( \19114 , \8977 , \19113 );
not \U$10296 ( \19115 , \17659 );
and \U$10297 ( \19116 , \9009 , \19115 );
not \U$10298 ( \19117 , \17736 );
and \U$10299 ( \19118 , \8966 , \19117 );
nor \U$10300 ( \19119 , \19116 , \19118 );
nand \U$10301 ( \19120 , \19112 , \19114 , \19119 );
not \U$10302 ( \19121 , \11067 );
and \U$10303 ( \19122 , \19121 , \17626 );
and \U$10304 ( \19123 , \18945 , \9034 );
nor \U$10305 ( \19124 , \19122 , \19123 );
not \U$10306 ( \19125 , \11060 );
and \U$10307 ( \19126 , \19125 , \17680 );
and \U$10308 ( \19127 , \17584 , \9014 );
nor \U$10309 ( \19128 , \19126 , \19127 );
nand \U$10310 ( \19129 , \19124 , \19128 );
nor \U$10311 ( \19130 , \19120 , \19129 );
nand \U$10312 ( \19131 , \19103 , \19110 , \19130 );
xnor \U$10313 ( \19132 , \19131 , \9044 );
nor \U$10314 ( \19133 , \19093 , \19132 );
nand \U$10315 ( \19134 , \19017 , \19054 , \19133 );
not \U$10316 ( \19135 , \19134 );
not \U$10317 ( \19136 , \9287 );
not \U$10318 ( \19137 , \17563 );
and \U$10319 ( \19138 , \19136 , \19137 );
or \U$10320 ( \19139 , \9273 , \17638 );
or \U$10321 ( \19140 , \9266 , \17771 );
nand \U$10322 ( \19141 , \19139 , \19140 );
not \U$10323 ( \19142 , \17587 );
and \U$10324 ( \19143 , \19142 , \9310 );
or \U$10325 ( \19144 , \19138 , \19141 , \19143 );
not \U$10326 ( \19145 , \19144 );
or \U$10327 ( \19146 , \11276 , \17647 );
or \U$10328 ( \19147 , \11270 , \18152 );
nand \U$10329 ( \19148 , \19146 , \19147 );
or \U$10330 ( \19149 , \9290 , \17554 );
or \U$10331 ( \19150 , \9282 , \17663 );
nand \U$10332 ( \19151 , \19149 , \19150 );
nor \U$10333 ( \19152 , \19148 , \19151 );
not \U$10334 ( \19153 , \18006 );
or \U$10335 ( \19154 , \11303 , \19153 );
not \U$10336 ( \19155 , \17576 );
or \U$10337 ( \19156 , \9270 , \19155 );
not \U$10338 ( \19157 , \17747 );
and \U$10339 ( \19158 , \9297 , \19157 );
not \U$10340 ( \19159 , \17597 );
and \U$10341 ( \19160 , \9262 , \19159 );
nor \U$10342 ( \19161 , \19158 , \19160 );
nand \U$10343 ( \19162 , \19154 , \19156 , \19161 );
not \U$10344 ( \19163 , \11293 );
and \U$10345 ( \19164 , \19163 , \17674 );
and \U$10346 ( \19165 , \18945 , \9319 );
nor \U$10347 ( \19166 , \19164 , \19165 );
not \U$10348 ( \19167 , \11288 );
and \U$10349 ( \19168 , \19167 , \17680 );
and \U$10350 ( \19169 , \17584 , \9302 );
nor \U$10351 ( \19170 , \19168 , \19169 );
nand \U$10352 ( \19171 , \19166 , \19170 );
nor \U$10353 ( \19172 , \19162 , \19171 );
nand \U$10354 ( \19173 , \19145 , \19152 , \19172 );
xnor \U$10355 ( \19174 , \19173 , \9327 );
not \U$10356 ( \19175 , \9419 );
not \U$10357 ( \19176 , \17744 );
and \U$10358 ( \19177 , \19175 , \19176 );
or \U$10359 ( \19178 , \9405 , \17638 );
or \U$10360 ( \19179 , \9398 , \17522 );
nand \U$10361 ( \19180 , \19178 , \19179 );
not \U$10362 ( \19181 , \17587 );
and \U$10363 ( \19182 , \19181 , \9444 );
or \U$10364 ( \19183 , \19177 , \19180 , \19182 );
not \U$10365 ( \19184 , \19183 );
or \U$10366 ( \19185 , \10455 , \17571 );
or \U$10367 ( \19186 , \11230 , \17623 );
nand \U$10368 ( \19187 , \19185 , \19186 );
or \U$10369 ( \19188 , \9422 , \17612 );
or \U$10370 ( \19189 , \9415 , \17549 );
nand \U$10371 ( \19190 , \19188 , \19189 );
nor \U$10372 ( \19191 , \19187 , \19190 );
not \U$10373 ( \19192 , \18006 );
or \U$10374 ( \19193 , \11259 , \19192 );
not \U$10375 ( \19194 , \17576 );
or \U$10376 ( \19195 , \9402 , \19194 );
not \U$10377 ( \19196 , \17559 );
and \U$10378 ( \19197 , \19196 , \9430 );
not \U$10379 ( \19198 , \17511 );
and \U$10380 ( \19199 , \9394 , \19198 );
nor \U$10381 ( \19200 , \19197 , \19199 );
nand \U$10382 ( \19201 , \19193 , \19195 , \19200 );
not \U$10383 ( \19202 , \11250 );
and \U$10384 ( \19203 , \19202 , \17674 );
and \U$10385 ( \19204 , \18945 , \9453 );
nor \U$10386 ( \19205 , \19203 , \19204 );
not \U$10387 ( \19206 , \11245 );
and \U$10388 ( \19207 , \19206 , \17680 );
and \U$10389 ( \19208 , \17584 , \9435 );
nor \U$10390 ( \19209 , \19207 , \19208 );
nand \U$10391 ( \19210 , \19205 , \19209 );
nor \U$10392 ( \19211 , \19201 , \19210 );
nand \U$10393 ( \19212 , \19184 , \19191 , \19211 );
xnor \U$10394 ( \19213 , \19212 , \9460 );
nor \U$10395 ( \19214 , \19174 , \19213 );
not \U$10396 ( \19215 , \17928 );
and \U$10397 ( \19216 , \9603 , \19215 );
not \U$10398 ( \19217 , \17522 );
and \U$10399 ( \19218 , \9613 , \19217 );
nor \U$10400 ( \19219 , \19216 , \19218 );
not \U$10401 ( \19220 , \17563 );
and \U$10402 ( \19221 , \9587 , \19220 );
not \U$10403 ( \19222 , \17659 );
and \U$10404 ( \19223 , \9606 , \19222 );
nor \U$10405 ( \19224 , \19221 , \19223 );
nand \U$10406 ( \19225 , \19219 , \19224 );
not \U$10407 ( \19226 , \19225 );
or \U$10408 ( \19227 , \9597 , \17733 );
or \U$10409 ( \19228 , \9647 , \17544 );
nand \U$10410 ( \19229 , \19227 , \19228 );
or \U$10411 ( \19230 , \12108 , \17554 );
or \U$10412 ( \19231 , \13538 , \17751 );
nand \U$10413 ( \19232 , \19230 , \19231 );
nor \U$10414 ( \19233 , \19229 , \19232 );
not \U$10415 ( \19234 , \17946 );
or \U$10416 ( \19235 , \11322 , \19234 );
not \U$10417 ( \19236 , \17576 );
or \U$10418 ( \19237 , \9637 , \19236 );
not \U$10419 ( \19238 , \9640 );
and \U$10420 ( \19239 , \19238 , \18006 );
and \U$10421 ( \19240 , \17588 , \9610 );
nor \U$10422 ( \19241 , \19239 , \19240 );
nand \U$10423 ( \19242 , \19235 , \19237 , \19241 );
not \U$10424 ( \19243 , \9632 );
and \U$10425 ( \19244 , \19243 , \17632 );
and \U$10426 ( \19245 , \17582 , \9628 );
nor \U$10427 ( \19246 , \19244 , \19245 );
not \U$10428 ( \19247 , \9625 );
and \U$10429 ( \19248 , \19247 , \17626 );
and \U$10430 ( \19249 , \18945 , \9619 );
nor \U$10431 ( \19250 , \19248 , \19249 );
nand \U$10432 ( \19251 , \19246 , \19250 );
nor \U$10433 ( \19252 , \19242 , \19251 );
nand \U$10434 ( \19253 , \19226 , \19233 , \19252 );
xnor \U$10435 ( \19254 , \19253 , \9653 );
not \U$10436 ( \19255 , \9354 );
not \U$10437 ( \19256 , \17656 );
and \U$10438 ( \19257 , \19255 , \19256 );
or \U$10439 ( \19258 , \9342 , \17638 );
or \U$10440 ( \19259 , \9335 , \17685 );
nand \U$10441 ( \19260 , \19258 , \19259 );
not \U$10442 ( \19261 , \17587 );
and \U$10443 ( \19262 , \19261 , \9380 );
or \U$10444 ( \19263 , \19257 , \19260 , \19262 );
not \U$10445 ( \19264 , \19263 );
or \U$10446 ( \19265 , \12141 , \17647 );
or \U$10447 ( \19266 , \11393 , \18152 );
nand \U$10448 ( \19267 , \19265 , \19266 );
or \U$10449 ( \19268 , \9357 , \17612 );
or \U$10450 ( \19269 , \12139 , \17663 );
nand \U$10451 ( \19270 , \19268 , \19269 );
nor \U$10452 ( \19271 , \19267 , \19270 );
not \U$10453 ( \19272 , \18006 );
or \U$10454 ( \19273 , \11352 , \19272 );
not \U$10455 ( \19274 , \17576 );
or \U$10456 ( \19275 , \9339 , \19274 );
not \U$10457 ( \19276 , \17747 );
and \U$10458 ( \19277 , \9364 , \19276 );
not \U$10459 ( \19278 , \17736 );
and \U$10460 ( \19279 , \9331 , \19278 );
nor \U$10461 ( \19280 , \19277 , \19279 );
nand \U$10462 ( \19281 , \19273 , \19275 , \19280 );
not \U$10463 ( \19282 , \11371 );
and \U$10464 ( \19283 , \19282 , \18945 );
and \U$10465 ( \19284 , \17674 , \9385 );
nor \U$10466 ( \19285 , \19283 , \19284 );
not \U$10467 ( \19286 , \11365 );
and \U$10468 ( \19287 , \19286 , \17680 );
and \U$10469 ( \19288 , \17584 , \9369 );
nor \U$10470 ( \19289 , \19287 , \19288 );
nand \U$10471 ( \19290 , \19285 , \19289 );
nor \U$10472 ( \19291 , \19281 , \19290 );
nand \U$10473 ( \19292 , \19264 , \19271 , \19291 );
xnor \U$10474 ( \19293 , \19292 , \9392 );
nor \U$10475 ( \19294 , \19254 , \19293 );
and \U$10476 ( \19295 , \19135 , \19214 , \19294 );
not \U$10477 ( \19296 , \17928 );
and \U$10478 ( \19297 , \9929 , \19296 );
not \U$10479 ( \19298 , \17685 );
and \U$10480 ( \19299 , \9939 , \19298 );
nor \U$10481 ( \19300 , \19297 , \19299 );
not \U$10482 ( \19301 , \17744 );
and \U$10483 ( \19302 , \9951 , \19301 );
not \U$10484 ( \19303 , \17659 );
and \U$10485 ( \19304 , \9932 , \19303 );
nor \U$10486 ( \19305 , \19302 , \19304 );
nand \U$10487 ( \19306 , \19300 , \19305 );
not \U$10488 ( \19307 , \19306 );
or \U$10489 ( \19308 , \13143 , \17733 );
or \U$10490 ( \19309 , \12282 , \17544 );
nand \U$10491 ( \19310 , \19308 , \19309 );
or \U$10492 ( \19311 , \9955 , \17612 );
or \U$10493 ( \19312 , \9948 , \17751 );
nand \U$10494 ( \19313 , \19311 , \19312 );
nor \U$10495 ( \19314 , \19310 , \19313 );
not \U$10496 ( \19315 , \17946 );
or \U$10497 ( \19316 , \11633 , \19315 );
not \U$10498 ( \19317 , \17576 );
or \U$10499 ( \19318 , \11635 , \19317 );
not \U$10500 ( \19319 , \11629 );
and \U$10501 ( \19320 , \19319 , \18006 );
and \U$10502 ( \19321 , \17588 , \9936 );
nor \U$10503 ( \19322 , \19320 , \19321 );
nand \U$10504 ( \19323 , \19316 , \19318 , \19322 );
not \U$10505 ( \19324 , \11623 );
and \U$10506 ( \19325 , \19324 , \17632 );
and \U$10507 ( \19326 , \17584 , \10709 );
nor \U$10508 ( \19327 , \19325 , \19326 );
not \U$10509 ( \19328 , \11620 );
and \U$10510 ( \19329 , \19328 , \17880 );
and \U$10511 ( \19330 , \18945 , \9968 );
nor \U$10512 ( \19331 , \19329 , \19330 );
nand \U$10513 ( \19332 , \19327 , \19331 );
nor \U$10514 ( \19333 , \19323 , \19332 );
nand \U$10515 ( \19334 , \19307 , \19314 , \19333 );
xnor \U$10516 ( \19335 , RIb7af450_258, \19334 );
not \U$10517 ( \19336 , \17928 );
and \U$10518 ( \19337 , \9533 , \19336 );
not \U$10519 ( \19338 , \17771 );
and \U$10520 ( \19339 , \19338 , \9545 );
nor \U$10521 ( \19340 , \19337 , \19339 );
not \U$10522 ( \19341 , \17656 );
and \U$10523 ( \19342 , \9518 , \19341 );
not \U$10524 ( \19343 , \17559 );
and \U$10525 ( \19344 , \19343 , \9536 );
nor \U$10526 ( \19345 , \19342 , \19344 );
nand \U$10527 ( \19346 , \19340 , \19345 );
not \U$10528 ( \19347 , \19346 );
or \U$10529 ( \19348 , \9527 , \17571 );
or \U$10530 ( \19349 , \9579 , \17623 );
nand \U$10531 ( \19350 , \19348 , \19349 );
or \U$10532 ( \19351 , \14434 , \17554 );
or \U$10533 ( \19352 , \13658 , \17549 );
nand \U$10534 ( \19353 , \19351 , \19352 );
nor \U$10535 ( \19354 , \19350 , \19353 );
not \U$10536 ( \19355 , \17946 );
or \U$10537 ( \19356 , \11589 , \19355 );
not \U$10538 ( \19357 , \17576 );
or \U$10539 ( \19358 , \9569 , \19357 );
not \U$10540 ( \19359 , \9572 );
and \U$10541 ( \19360 , \19359 , \18006 );
and \U$10542 ( \19361 , \17588 , \9542 );
nor \U$10543 ( \19362 , \19360 , \19361 );
nand \U$10544 ( \19363 , \19356 , \19358 , \19362 );
not \U$10545 ( \19364 , \9564 );
and \U$10546 ( \19365 , \19364 , \17632 );
and \U$10547 ( \19366 , \17584 , \9560 );
nor \U$10548 ( \19367 , \19365 , \19366 );
not \U$10549 ( \19368 , \9557 );
and \U$10550 ( \19369 , \19368 , \17880 );
and \U$10551 ( \19370 , \18945 , \9551 );
nor \U$10552 ( \19371 , \19369 , \19370 );
nand \U$10553 ( \19372 , \19367 , \19371 );
nor \U$10554 ( \19373 , \19363 , \19372 );
nand \U$10555 ( \19374 , \19347 , \19354 , \19373 );
xnor \U$10556 ( \19375 , RIb7af3d8_259, \19374 );
not \U$10557 ( \19376 , \17946 );
or \U$10558 ( \19377 , \11681 , \19376 );
not \U$10559 ( \19378 , \17576 );
or \U$10560 ( \19379 , \11684 , \19378 );
not \U$10561 ( \19380 , \17563 );
and \U$10562 ( \19381 , \10001 , \19380 );
not \U$10563 ( \19382 , \17601 );
and \U$10564 ( \19383 , \10041 , \19382 );
nor \U$10565 ( \19384 , \19381 , \19383 );
nand \U$10566 ( \19385 , \19377 , \19379 , \19384 );
not \U$10567 ( \19386 , \11693 );
and \U$10568 ( \19387 , \19386 , \17632 );
and \U$10569 ( \19388 , \17584 , \10027 );
nor \U$10570 ( \19389 , \19387 , \19388 );
not \U$10571 ( \19390 , \11698 );
and \U$10572 ( \19391 , \19390 , \17880 );
and \U$10573 ( \19392 , \18945 , \10035 );
nor \U$10574 ( \19393 , \19391 , \19392 );
nand \U$10575 ( \19394 , \19389 , \19393 );
nor \U$10576 ( \19395 , \19385 , \19394 );
not \U$10577 ( \19396 , \17969 );
or \U$10578 ( \19397 , \10013 , \19396 );
not \U$10579 ( \19398 , \17624 );
or \U$10580 ( \19399 , \11674 , \19398 );
not \U$10581 ( \19400 , \17928 );
and \U$10582 ( \19401 , \10009 , \19400 );
not \U$10583 ( \19402 , \17522 );
and \U$10584 ( \19403 , \10020 , \19402 );
nor \U$10585 ( \19404 , \19401 , \19403 );
nand \U$10586 ( \19405 , \19397 , \19399 , \19404 );
not \U$10587 ( \19406 , \17555 );
or \U$10588 ( \19407 , \10005 , \19406 );
not \U$10589 ( \19408 , \17550 );
or \U$10590 ( \19409 , \9997 , \19408 );
not \U$10591 ( \19410 , \11666 );
and \U$10592 ( \19411 , \19410 , \17572 );
and \U$10593 ( \19412 , \17588 , \10017 );
nor \U$10594 ( \19413 , \19411 , \19412 );
nand \U$10595 ( \19414 , \19407 , \19409 , \19413 );
nor \U$10596 ( \19415 , \19405 , \19414 );
nand \U$10597 ( \19416 , \19395 , \19415 );
xnor \U$10598 ( \19417 , \19416 , \10055 );
not \U$10599 ( \19418 , \17928 );
and \U$10600 ( \19419 , \9874 , \19418 );
not \U$10601 ( \19420 , \17771 );
and \U$10602 ( \19421 , \9886 , \19420 );
nor \U$10603 ( \19422 , \19419 , \19421 );
not \U$10604 ( \19423 , \17656 );
and \U$10605 ( \19424 , \9859 , \19423 );
not \U$10606 ( \19425 , \17747 );
and \U$10607 ( \19426 , \9877 , \19425 );
nor \U$10608 ( \19427 , \19424 , \19426 );
nand \U$10609 ( \19428 , \19422 , \19427 );
not \U$10610 ( \19429 , \19428 );
or \U$10611 ( \19430 , \9868 , \17647 );
or \U$10612 ( \19431 , \9921 , \18152 );
nand \U$10613 ( \19432 , \19430 , \19431 );
or \U$10614 ( \19433 , \12183 , \17554 );
or \U$10615 ( \19434 , \12178 , \17663 );
nand \U$10616 ( \19435 , \19433 , \19434 );
nor \U$10617 ( \19436 , \19432 , \19435 );
not \U$10618 ( \19437 , \17946 );
or \U$10619 ( \19438 , \11718 , \19437 );
not \U$10620 ( \19439 , \17576 );
or \U$10621 ( \19440 , \9911 , \19439 );
not \U$10622 ( \19441 , \9914 );
and \U$10623 ( \19442 , \19441 , \18006 );
and \U$10624 ( \19443 , \17588 , \9881 );
nor \U$10625 ( \19444 , \19442 , \19443 );
nand \U$10626 ( \19445 , \19438 , \19440 , \19444 );
not \U$10627 ( \19446 , \9906 );
and \U$10628 ( \19447 , \19446 , \17632 );
and \U$10629 ( \19448 , \17584 , \9902 );
nor \U$10630 ( \19449 , \19447 , \19448 );
not \U$10631 ( \19450 , \9898 );
and \U$10632 ( \19451 , \19450 , \17880 );
and \U$10633 ( \19452 , \18945 , \9892 );
nor \U$10634 ( \19453 , \19451 , \19452 );
nand \U$10635 ( \19454 , \19449 , \19453 );
nor \U$10636 ( \19455 , \19445 , \19454 );
nand \U$10637 ( \19456 , \19429 , \19436 , \19455 );
xnor \U$10638 ( \19457 , \19456 , \9927 );
nor \U$10639 ( \19458 , \19417 , \19457 );
nand \U$10640 ( \19459 , \19335 , \19375 , \19458 );
not \U$10641 ( \19460 , \9148 );
not \U$10642 ( \19461 , \17656 );
and \U$10643 ( \19462 , \19460 , \19461 );
or \U$10644 ( \19463 , \9133 , \17519 );
or \U$10645 ( \19464 , \9125 , \17685 );
nand \U$10646 ( \19465 , \19463 , \19464 );
not \U$10647 ( \19466 , \17587 );
and \U$10648 ( \19467 , \19466 , \9172 );
or \U$10649 ( \19468 , \19462 , \19465 , \19467 );
not \U$10650 ( \19469 , \19468 );
or \U$10651 ( \19470 , \11416 , \17647 );
or \U$10652 ( \19471 , \11410 , \18152 );
nand \U$10653 ( \19472 , \19470 , \19471 );
or \U$10654 ( \19473 , \9151 , \17612 );
or \U$10655 ( \19474 , \9143 , \17663 );
nand \U$10656 ( \19475 , \19473 , \19474 );
nor \U$10657 ( \19476 , \19472 , \19475 );
not \U$10658 ( \19477 , \18006 );
or \U$10659 ( \19478 , \11441 , \19477 );
nand \U$10660 ( \19479 , \9129 , \17576 );
not \U$10661 ( \19480 , \17747 );
and \U$10662 ( \19481 , \9157 , \19480 );
not \U$10663 ( \19482 , \17736 );
and \U$10664 ( \19483 , \9121 , \19482 );
nor \U$10665 ( \19484 , \19481 , \19483 );
nand \U$10666 ( \19485 , \19478 , \19479 , \19484 );
and \U$10667 ( \19486 , \18945 , \9180 );
and \U$10668 ( \19487 , \9176 , \17674 );
nor \U$10669 ( \19488 , \19486 , \19487 );
and \U$10670 ( \19489 , \17584 , \9163 );
and \U$10671 ( \19490 , \9159 , \17680 );
nor \U$10672 ( \19491 , \19489 , \19490 );
nand \U$10673 ( \19492 , \19488 , \19491 );
nor \U$10674 ( \19493 , \19485 , \19492 );
nand \U$10675 ( \19494 , \19469 , \19476 , \19493 );
xnor \U$10676 ( \19495 , RIb7af6a8_253, \19494 );
not \U$10677 ( \19496 , \9073 );
not \U$10678 ( \19497 , \17563 );
and \U$10679 ( \19498 , \19496 , \19497 );
or \U$10680 ( \19499 , \9058 , \17519 );
or \U$10681 ( \19500 , \9050 , \17522 );
nand \U$10682 ( \19501 , \19499 , \19500 );
not \U$10683 ( \19502 , \17587 );
and \U$10684 ( \19503 , \19502 , \9102 );
or \U$10685 ( \19504 , \19498 , \19501 , \19503 );
not \U$10686 ( \19505 , \19504 );
or \U$10687 ( \19506 , \11458 , \17733 );
or \U$10688 ( \19507 , \11452 , \17544 );
nand \U$10689 ( \19508 , \19506 , \19507 );
or \U$10690 ( \19509 , \9076 , \17554 );
or \U$10691 ( \19510 , \9068 , \17751 );
nand \U$10692 ( \19511 , \19509 , \19510 );
nor \U$10693 ( \19512 , \19508 , \19511 );
nand \U$10694 ( \19513 , \9081 , \18006 );
nand \U$10695 ( \19514 , \9054 , \17576 );
not \U$10696 ( \19515 , \17659 );
and \U$10697 ( \19516 , \9085 , \19515 );
not \U$10698 ( \19517 , \17511 );
and \U$10699 ( \19518 , \9046 , \19517 );
nor \U$10700 ( \19519 , \19516 , \19518 );
nand \U$10701 ( \19520 , \19513 , \19514 , \19519 );
and \U$10702 ( \19521 , \18945 , \9112 );
and \U$10703 ( \19522 , \9107 , \17880 );
nor \U$10704 ( \19523 , \19521 , \19522 );
and \U$10705 ( \19524 , \17584 , \9093 );
and \U$10706 ( \19525 , \9089 , \17680 );
nor \U$10707 ( \19526 , \19524 , \19525 );
nand \U$10708 ( \19527 , \19523 , \19526 );
nor \U$10709 ( \19528 , \19520 , \19527 );
nand \U$10710 ( \19529 , \19505 , \19512 , \19528 );
xnor \U$10711 ( \19530 , RIb7af720_252, \19529 );
nand \U$10712 ( \19531 , \9847 , \17946 );
nand \U$10713 ( \19532 , \9838 , \17576 );
not \U$10714 ( \19533 , \17744 );
and \U$10715 ( \19534 , \9790 , \19533 );
not \U$10716 ( \19535 , \17533 );
and \U$10717 ( \19536 , \19535 , \9842 );
nor \U$10718 ( \19537 , \19534 , \19536 );
nand \U$10719 ( \19538 , \19531 , \19532 , \19537 );
and \U$10720 ( \19539 , \17584 , \9830 );
and \U$10721 ( \19540 , \9833 , \17632 );
nor \U$10722 ( \19541 , \19539 , \19540 );
and \U$10723 ( \19542 , \18945 , \9822 );
and \U$10724 ( \19543 , \9826 , \17626 );
nor \U$10725 ( \19544 , \19542 , \19543 );
nand \U$10726 ( \19545 , \19541 , \19544 );
nor \U$10727 ( \19546 , \19538 , \19545 );
nand \U$10728 ( \19547 , \9808 , \17969 );
nand \U$10729 ( \19548 , \9850 , \17624 );
not \U$10730 ( \19549 , \17928 );
and \U$10731 ( \19550 , \9805 , \19549 );
not \U$10732 ( \19551 , \17685 );
and \U$10733 ( \19552 , \9816 , \19551 );
nor \U$10734 ( \19553 , \19550 , \19552 );
nand \U$10735 ( \19554 , \19547 , \19548 , \19553 );
nand \U$10736 ( \19555 , \9794 , \17555 );
nand \U$10737 ( \19556 , \9801 , \17550 );
and \U$10738 ( \19557 , \17588 , \9813 );
and \U$10739 ( \19558 , \9797 , \17572 );
nor \U$10740 ( \19559 , \19557 , \19558 );
nand \U$10741 ( \19560 , \19555 , \19556 , \19559 );
nor \U$10742 ( \19561 , \19554 , \19560 );
nand \U$10743 ( \19562 , \19546 , \19561 );
xnor \U$10744 ( \19563 , \19562 , \9857 );
not \U$10745 ( \19564 , \8894 );
not \U$10746 ( \19565 , \17744 );
and \U$10747 ( \19566 , \19564 , \19565 );
or \U$10748 ( \19567 , \8861 , \17519 );
or \U$10749 ( \19568 , \8844 , \17771 );
nand \U$10750 ( \19569 , \19567 , \19568 );
not \U$10751 ( \19570 , \17587 );
and \U$10752 ( \19571 , \8940 , \19570 );
or \U$10753 ( \19572 , \19566 , \19569 , \19571 );
not \U$10754 ( \19573 , \19572 );
or \U$10755 ( \19574 , \12351 , \17571 );
or \U$10756 ( \19575 , \11565 , \17623 );
nand \U$10757 ( \19576 , \19574 , \19575 );
or \U$10758 ( \19577 , \8897 , \17612 );
or \U$10759 ( \19578 , \8882 , \17549 );
nand \U$10760 ( \19579 , \19577 , \19578 );
nor \U$10761 ( \19580 , \19576 , \19579 );
nand \U$10762 ( \19581 , \8904 , \18006 );
nand \U$10763 ( \19582 , \8852 , \17576 );
not \U$10764 ( \19583 , \17559 );
and \U$10765 ( \19584 , \19583 , \8915 );
not \U$10766 ( \19585 , \17597 );
and \U$10767 ( \19586 , \8827 , \19585 );
nor \U$10768 ( \19587 , \19584 , \19586 );
nand \U$10769 ( \19588 , \19581 , \19582 , \19587 );
and \U$10770 ( \19589 , \18945 , \8953 );
and \U$10771 ( \19590 , \8947 , \17626 );
nor \U$10772 ( \19591 , \19589 , \19590 );
and \U$10773 ( \19592 , \17584 , \8927 );
and \U$10774 ( \19593 , \8921 , \17680 );
nor \U$10775 ( \19594 , \19592 , \19593 );
nand \U$10776 ( \19595 , \19591 , \19594 );
nor \U$10777 ( \19596 , \19588 , \19595 );
nand \U$10778 ( \19597 , \19573 , \19580 , \19596 );
xnor \U$10779 ( \19598 , \19597 , \8964 );
nor \U$10780 ( \19599 , \19563 , \19598 );
nand \U$10781 ( \19600 , \19495 , \19530 , \19599 );
nor \U$10782 ( \19601 , \19459 , \19600 );
nand \U$10783 ( \19602 , \18980 , \19295 , \19601 );
not \U$10784 ( \19603 , \19602 );
nor \U$10785 ( \19604 , \18940 , \19603 );
and \U$10786 ( \19605 , \18300 , \19604 );
not \U$10787 ( \19606 , \17507 );
buf \U$10788 ( \19607 , RIea91330_6888);
buf \U$10789 ( \19608 , \13927 );
buf \U$10790 ( \19609 , \12456 );
buf \U$10791 ( \19610 , \12458 );
buf \U$10792 ( \19611 , \8870 );
or \U$10793 ( \19612 , \19610 , \19611 );
or \U$10794 ( \19613 , \19609 , \19612 );
and \U$10795 ( \19614 , \19608 , \19613 );
and \U$10796 ( \19615 , \19607 , \19614 );
buf \U$10797 ( \19616 , \19615 );
not \U$10798 ( \19617 , \19616 );
not \U$10799 ( \19618 , \19611 );
buf \U$10800 ( \19619 , \19618 );
not \U$10801 ( \19620 , \19619 );
xnor \U$10802 ( \19621 , \19610 , \19611 );
buf \U$10803 ( \19622 , \19621 );
not \U$10804 ( \19623 , \19622 );
nand \U$10805 ( \19624 , \19620 , \19623 );
xnor \U$10806 ( \19625 , \19609 , \19612 );
buf \U$10807 ( \19626 , \19625 );
not \U$10808 ( \19627 , \19626 );
xor \U$10809 ( \19628 , \19608 , \19613 );
buf \U$10810 ( \19629 , \19628 );
not \U$10811 ( \19630 , \19629 );
nand \U$10812 ( \19631 , \19627 , \19630 );
or \U$10813 ( \19632 , \19624 , \19631 );
xor \U$10814 ( \19633 , \19607 , \19614 );
buf \U$10815 ( \19634 , \19633 );
nand \U$10816 ( \19635 , \19632 , \19634 );
nand \U$10817 ( \19636 , \19617 , \19635 );
not \U$10818 ( \19637 , \19636 );
not \U$10819 ( \19638 , \19603 );
or \U$10820 ( \19639 , \19637 , \19638 );
not \U$10821 ( \19640 , \19639 );
not \U$10822 ( \19641 , \19603 );
or \U$10823 ( \19642 , \19636 , \19641 );
not \U$10824 ( \19643 , \19642 );
or \U$10825 ( \19644 , \19640 , \19643 );
not \U$10826 ( \19645 , \19644 );
or \U$10827 ( \19646 , \18940 , \19645 );
or \U$10828 ( \19647 , \19606 , \19646 );
buf \U$10829 ( \19648 , RIea91330_6888);
buf \U$10830 ( \19649 , \13253 );
buf \U$10831 ( \19650 , \12456 );
buf \U$10832 ( \19651 , \12458 );
or \U$10833 ( \19652 , \19650 , \19651 );
and \U$10834 ( \19653 , \19649 , \19652 );
and \U$10835 ( \19654 , \19648 , \19653 );
buf \U$10836 ( \19655 , \19654 );
not \U$10837 ( \19656 , \19655 );
buf \U$10838 ( \19657 , \8835 );
not \U$10839 ( \19658 , \19657 );
not \U$10840 ( \19659 , \19651 );
buf \U$10841 ( \19660 , \19659 );
not \U$10842 ( \19661 , \19660 );
nand \U$10843 ( \19662 , \19658 , \19661 );
xnor \U$10844 ( \19663 , \19650 , \19651 );
buf \U$10845 ( \19664 , \19663 );
not \U$10846 ( \19665 , \19664 );
xor \U$10847 ( \19666 , \19649 , \19652 );
buf \U$10848 ( \19667 , \19666 );
not \U$10849 ( \19668 , \19667 );
nand \U$10850 ( \19669 , \19665 , \19668 );
or \U$10851 ( \19670 , \19662 , \19669 );
xor \U$10852 ( \19671 , \19648 , \19653 );
buf \U$10853 ( \19672 , \19671 );
nand \U$10854 ( \19673 , \19670 , \19672 );
and \U$10855 ( \19674 , \19656 , \19673 );
not \U$10856 ( \19675 , \18940 );
or \U$10857 ( \19676 , \19674 , \19675 );
not \U$10858 ( \19677 , \19676 );
nand \U$10859 ( \19678 , \19674 , \18940 );
not \U$10860 ( \19679 , \19678 );
or \U$10861 ( \19680 , \19677 , \19679 );
not \U$10862 ( \19681 , \19680 );
or \U$10863 ( \19682 , \16703 , \19681 );
nand \U$10864 ( \19683 , \19647 , \19682 );
nor \U$10865 ( \19684 , \19605 , \19683 );
or \U$10866 ( \19685 , \12451 , \19684 );
buf \U$10867 ( \19686 , RIea91330_6888);
buf \U$10868 ( \19687 , \13927 );
buf \U$10869 ( \19688 , \12456 );
buf \U$10870 ( \19689 , \12458 );
buf \U$10871 ( \19690 , \10937 );
and \U$10872 ( \19691 , \19689 , \19690 );
or \U$10873 ( \19692 , \19688 , \19691 );
and \U$10874 ( \19693 , \19687 , \19692 );
and \U$10875 ( \19694 , \19686 , \19693 );
buf \U$10876 ( \19695 , \19694 );
not \U$10877 ( \19696 , \19690 );
buf \U$10878 ( \19697 , \19696 );
not \U$10879 ( \19698 , \19697 );
xor \U$10880 ( \19699 , \19689 , \19690 );
buf \U$10881 ( \19700 , \19699 );
not \U$10882 ( \19701 , \19700 );
nand \U$10883 ( \19702 , \19698 , \19701 );
xnor \U$10884 ( \19703 , \19688 , \19691 );
buf \U$10885 ( \19704 , \19703 );
not \U$10886 ( \19705 , \19704 );
xor \U$10887 ( \19706 , \19687 , \19692 );
buf \U$10888 ( \19707 , \19706 );
not \U$10889 ( \19708 , \19707 );
nand \U$10890 ( \19709 , \19705 , \19708 );
or \U$10891 ( \19710 , \19702 , \19709 );
xor \U$10892 ( \19711 , \19686 , \19693 );
buf \U$10893 ( \19712 , \19711 );
nand \U$10894 ( \19713 , \19710 , \19712 );
not \U$10895 ( \19714 , \19713 );
or \U$10896 ( \19715 , \19695 , \19714 );
not \U$10897 ( \19716 , \11750 );
or \U$10898 ( \19717 , \19715 , \19716 );
not \U$10899 ( \19718 , \19717 );
not \U$10900 ( \19719 , \19715 );
not \U$10901 ( \19720 , \11750 );
or \U$10902 ( \19721 , \19719 , \19720 );
not \U$10903 ( \19722 , \19721 );
or \U$10904 ( \19723 , \19718 , \19722 );
not \U$10905 ( \19724 , \19723 );
or \U$10906 ( \19725 , \10915 , \19724 );
not \U$10907 ( \19726 , \19725 );
and \U$10908 ( \19727 , \19726 , \12449 , \10931 );
not \U$10909 ( \19728 , \12449 );
not \U$10910 ( \19729 , \19728 );
buf \U$10911 ( \19730 , RIea91330_6888);
buf \U$10912 ( \19731 , \13253 );
buf \U$10913 ( \19732 , \12456 );
not \U$10914 ( \19733 , \19732 );
not \U$10915 ( \19734 , \19733 );
and \U$10916 ( \19735 , \19731 , \19734 );
and \U$10917 ( \19736 , \19730 , \19735 );
buf \U$10918 ( \19737 , \19736 );
not \U$10919 ( \19738 , \19737 );
buf \U$10920 ( \19739 , \10919 );
buf \U$10921 ( \19740 , \12458 );
or \U$10922 ( \19741 , \19739 , \19740 );
buf \U$10923 ( \19742 , \19733 );
xor \U$10924 ( \19743 , \19734 , \19731 );
buf \U$10925 ( \19744 , \19743 );
or \U$10926 ( \19745 , \19742 , \19744 );
or \U$10927 ( \19746 , \19741 , \19745 );
xor \U$10928 ( \19747 , \19730 , \19735 );
buf \U$10929 ( \19748 , \19747 );
nand \U$10930 ( \19749 , \19746 , \19748 );
nand \U$10931 ( \19750 , \19738 , \19749 );
not \U$10932 ( \19751 , \10915 );
or \U$10933 ( \19752 , \19750 , \19751 );
not \U$10934 ( \19753 , \19752 );
not \U$10935 ( \19754 , \19750 );
not \U$10936 ( \19755 , \10915 );
or \U$10937 ( \19756 , \19754 , \19755 );
not \U$10938 ( \19757 , \19756 );
or \U$10939 ( \19758 , \19753 , \19757 );
and \U$10940 ( \19759 , \19729 , \19758 , \10066 );
buf \U$10941 ( \19760 , RIea91330_6888);
buf \U$10942 ( \19761 , \12454 );
buf \U$10943 ( \19762 , \12456 );
buf \U$10944 ( \19763 , \12458 );
buf \U$10945 ( \19764 , \10919 );
or \U$10946 ( \19765 , \19763 , \19764 );
and \U$10947 ( \19766 , \19762 , \19765 );
and \U$10948 ( \19767 , \19761 , \19766 );
and \U$10949 ( \19768 , \19760 , \19767 );
buf \U$10950 ( \19769 , \19768 );
not \U$10951 ( \19770 , \19769 );
not \U$10952 ( \19771 , \19764 );
buf \U$10953 ( \19772 , \19771 );
not \U$10954 ( \19773 , \19772 );
xnor \U$10955 ( \19774 , \19763 , \19764 );
buf \U$10956 ( \19775 , \19774 );
not \U$10957 ( \19776 , \19775 );
nand \U$10958 ( \19777 , \19773 , \19776 );
xor \U$10959 ( \19778 , \19762 , \19765 );
buf \U$10960 ( \19779 , \19778 );
not \U$10961 ( \19780 , \19779 );
xor \U$10962 ( \19781 , \19761 , \19766 );
buf \U$10963 ( \19782 , \19781 );
not \U$10964 ( \19783 , \19782 );
nand \U$10965 ( \19784 , \19780 , \19783 );
or \U$10966 ( \19785 , \19777 , \19784 );
xor \U$10967 ( \19786 , \19760 , \19767 );
buf \U$10968 ( \19787 , \19786 );
nand \U$10969 ( \19788 , \19785 , \19787 );
nand \U$10970 ( \19789 , \19770 , \19788 );
not \U$10971 ( \19790 , \19728 );
or \U$10972 ( \19791 , \19789 , \19790 );
not \U$10973 ( \19792 , \19791 );
not \U$10974 ( \19793 , \19789 );
not \U$10975 ( \19794 , \19728 );
or \U$10976 ( \19795 , \19793 , \19794 );
not \U$10977 ( \19796 , \19795 );
or \U$10978 ( \19797 , \19792 , \19796 );
not \U$10979 ( \19798 , \19797 );
not \U$10980 ( \19799 , \19798 );
and \U$10981 ( \19800 , \11781 , \19799 );
nor \U$10982 ( \19801 , \19727 , \19759 , \19800 );
and \U$10983 ( \19802 , \19685 , \19801 );
nand \U$10984 ( \19803 , \14049 , \12513 );
not \U$10985 ( \19804 , \14044 );
nand \U$10986 ( \19805 , \19804 , \10062 );
nand \U$10987 ( \19806 , \19803 , \19805 );
not \U$10988 ( \19807 , \19806 );
not \U$10989 ( \19808 , \14037 );
not \U$10990 ( \19809 , \19808 );
or \U$10991 ( \19810 , \9500 , \19809 );
not \U$10992 ( \19811 , \14054 );
or \U$10993 ( \19812 , \9498 , \19811 );
and \U$10994 ( \19813 , \19807 , \19810 , \19812 );
not \U$10995 ( \19814 , \14057 );
not \U$10996 ( \19815 , \19814 );
or \U$10997 ( \19816 , \19815 , \9506 );
or \U$10998 ( \19817 , \9504 , \14197 );
nand \U$10999 ( \19818 , \19816 , \19817 );
or \U$11000 ( \19819 , \9509 , \14075 );
or \U$11001 ( \19820 , \9511 , \14180 );
nand \U$11002 ( \19821 , \19819 , \19820 );
nor \U$11003 ( \19822 , \19818 , \19821 );
not \U$11004 ( \19823 , \14135 );
not \U$11005 ( \19824 , \19823 );
or \U$11006 ( \19825 , \9467 , \19824 );
not \U$11007 ( \19826 , \14018 );
or \U$11008 ( \19827 , \9463 , \19826 );
not \U$11009 ( \19828 , \14183 );
and \U$11010 ( \19829 , \9472 , \19828 );
not \U$11011 ( \19830 , \14121 );
and \U$11012 ( \19831 , \9476 , \19830 );
nor \U$11013 ( \19832 , \19829 , \19831 );
nand \U$11014 ( \19833 , \19825 , \19827 , \19832 );
or \U$11015 ( \19834 , \9482 , \14065 );
not \U$11016 ( \19835 , \14024 );
nand \U$11017 ( \19836 , \19835 , \10168 );
nand \U$11018 ( \19837 , \14080 , \10163 );
not \U$11019 ( \19838 , \14125 );
or \U$11020 ( \19839 , \9480 , \19838 );
and \U$11021 ( \19840 , \19834 , \19836 , \19837 , \19839 );
not \U$11022 ( \19841 , \19840 );
nor \U$11023 ( \19842 , \19833 , \19841 );
nand \U$11024 ( \19843 , \19813 , \19822 , \19842 );
not \U$11025 ( \19844 , \19843 );
and \U$11026 ( \19845 , \14272 , \8970 );
not \U$11027 ( \19846 , \14125 );
or \U$11028 ( \19847 , \10370 , \19846 );
not \U$11029 ( \19848 , \19847 );
or \U$11030 ( \19849 , \11073 , \14121 );
or \U$11031 ( \19850 , \8980 , \14069 );
nand \U$11032 ( \19851 , \19849 , \19850 );
nor \U$11033 ( \19852 , \19845 , \19848 , \19851 );
or \U$11034 ( \19853 , \8991 , \14135 );
or \U$11035 ( \19854 , \11046 , \14138 );
nand \U$11036 ( \19855 , \19853 , \19854 );
not \U$11037 ( \19856 , \8999 );
or \U$11038 ( \19857 , \19856 , \14180 );
or \U$11039 ( \19858 , \8997 , \13995 );
nand \U$11040 ( \19859 , \19857 , \19858 );
nor \U$11041 ( \19860 , \19855 , \19859 );
or \U$11042 ( \19861 , \8967 , \14079 );
nand \U$11043 ( \19862 , \19804 , \9006 );
nand \U$11044 ( \19863 , \19835 , \8976 );
nand \U$11045 ( \19864 , \9020 , \14076 );
and \U$11046 ( \19865 , \19861 , \19862 , \19863 , \19864 );
not \U$11047 ( \19866 , \19865 );
not \U$11048 ( \19867 , \19866 );
and \U$11049 ( \19868 , \14049 , \9011 );
and \U$11050 ( \19869 , \19808 , \9014 );
nor \U$11051 ( \19870 , \19868 , \19869 );
not \U$11052 ( \19871 , \11064 );
and \U$11053 ( \19872 , \19871 , \14054 );
and \U$11054 ( \19873 , \19814 , \9030 );
nor \U$11055 ( \19874 , \19872 , \19873 );
and \U$11056 ( \19875 , \19867 , \19870 , \19874 );
nand \U$11057 ( \19876 , \19852 , \19860 , \19875 );
xnor \U$11058 ( \19877 , RIb7b94a0_249, \19876 );
and \U$11059 ( \19878 , \14272 , \9193 );
not \U$11060 ( \19879 , \14033 );
or \U$11061 ( \19880 , \10323 , \19879 );
not \U$11062 ( \19881 , \19880 );
or \U$11063 ( \19882 , \11125 , \14201 );
or \U$11064 ( \19883 , \11954 , \14197 );
nand \U$11065 ( \19884 , \19882 , \19883 );
nor \U$11066 ( \19885 , \19878 , \19881 , \19884 );
or \U$11067 ( \19886 , \11098 , \14104 );
or \U$11068 ( \19887 , \11101 , \14017 );
nand \U$11069 ( \19888 , \19886 , \19887 );
not \U$11070 ( \19889 , \9219 );
or \U$11071 ( \19890 , \19889 , \14180 );
or \U$11072 ( \19891 , \9217 , \14183 );
nand \U$11073 ( \19892 , \19890 , \19891 );
nor \U$11074 ( \19893 , \19888 , \19892 );
or \U$11075 ( \19894 , \9197 , \14161 );
nand \U$11076 ( \19895 , \19804 , \9225 );
nand \U$11077 ( \19896 , \19835 , \9204 );
nand \U$11078 ( \19897 , \9239 , \14091 );
and \U$11079 ( \19898 , \19894 , \19895 , \19896 , \19897 );
not \U$11080 ( \19899 , \19898 );
not \U$11081 ( \19900 , \19899 );
and \U$11082 ( \19901 , \14049 , \9230 );
and \U$11083 ( \19902 , \19808 , \9233 );
nor \U$11084 ( \19903 , \19901 , \19902 );
not \U$11085 ( \19904 , \11117 );
and \U$11086 ( \19905 , \19904 , \14054 );
and \U$11087 ( \19906 , \19814 , \9247 );
nor \U$11088 ( \19907 , \19905 , \19906 );
and \U$11089 ( \19908 , \19900 , \19903 , \19907 );
nand \U$11090 ( \19909 , \19885 , \19893 , \19908 );
xnor \U$11091 ( \19910 , RIb7b9518_248, \19909 );
or \U$11092 ( \19911 , \9668 , \14075 );
or \U$11093 ( \19912 , \13344 , \14079 );
nand \U$11094 ( \19913 , \19911 , \19912 );
not \U$11095 ( \19914 , \19913 );
nand \U$11096 ( \19915 , \19804 , \9660 );
nand \U$11097 ( \19916 , \19835 , \9656 );
and \U$11098 ( \19917 , \19914 , \19915 , \19916 );
or \U$11099 ( \19918 , \9676 , \14135 );
or \U$11100 ( \19919 , \11923 , \14138 );
nand \U$11101 ( \19920 , \19918 , \19919 );
not \U$11102 ( \19921 , \9682 );
or \U$11103 ( \19922 , \19921 , \14180 );
or \U$11104 ( \19923 , \9680 , \13995 );
nand \U$11105 ( \19924 , \19922 , \19923 );
nor \U$11106 ( \19925 , \19920 , \19924 );
nand \U$11107 ( \19926 , \14049 , \9687 );
nand \U$11108 ( \19927 , \9690 , \19808 );
and \U$11109 ( \19928 , \19814 , \9692 );
and \U$11110 ( \19929 , \9695 , \14054 );
nor \U$11111 ( \19930 , \19928 , \19929 );
nand \U$11112 ( \19931 , \19926 , \19927 , \19930 );
nand \U$11113 ( \19932 , \9713 , \14125 );
nand \U$11114 ( \19933 , \9710 , \14272 );
not \U$11115 ( \19934 , \14201 );
and \U$11116 ( \19935 , \9701 , \19934 );
not \U$11117 ( \19936 , \14117 );
and \U$11118 ( \19937 , \9706 , \19936 );
nor \U$11119 ( \19938 , \19935 , \19937 );
nand \U$11120 ( \19939 , \19932 , \19933 , \19938 );
nor \U$11121 ( \19940 , \19931 , \19939 );
nand \U$11122 ( \19941 , \19917 , \19925 , \19940 );
xnor \U$11123 ( \19942 , \19941 , \9719 );
or \U$11124 ( \19943 , \9732 , \14075 );
or \U$11125 ( \19944 , \13305 , \14079 );
nand \U$11126 ( \19945 , \19943 , \19944 );
not \U$11127 ( \19946 , \19945 );
nand \U$11128 ( \19947 , \19804 , \9724 );
nand \U$11129 ( \19948 , \19835 , \9721 );
and \U$11130 ( \19949 , \19946 , \19947 , \19948 );
or \U$11131 ( \19950 , \9740 , \14005 );
or \U$11132 ( \19951 , \11876 , \14101 );
nand \U$11133 ( \19952 , \19950 , \19951 );
not \U$11134 ( \19953 , \9747 );
or \U$11135 ( \19954 , \19953 , \14180 );
or \U$11136 ( \19955 , \9745 , \14097 );
nand \U$11137 ( \19956 , \19954 , \19955 );
nor \U$11138 ( \19957 , \19952 , \19956 );
nand \U$11139 ( \19958 , \14049 , \9752 );
nand \U$11140 ( \19959 , \9755 , \19808 );
and \U$11141 ( \19960 , \19814 , \9759 );
and \U$11142 ( \19961 , \9763 , \14054 );
nor \U$11143 ( \19962 , \19960 , \19961 );
nand \U$11144 ( \19963 , \19958 , \19959 , \19962 );
nand \U$11145 ( \19964 , \9779 , \14125 );
nand \U$11146 ( \19965 , \9776 , \14272 );
not \U$11147 ( \19966 , \13998 );
and \U$11148 ( \19967 , \9769 , \19966 );
not \U$11149 ( \19968 , \14117 );
and \U$11150 ( \19969 , \9772 , \19968 );
nor \U$11151 ( \19970 , \19967 , \19969 );
nand \U$11152 ( \19971 , \19964 , \19965 , \19970 );
nor \U$11153 ( \19972 , \19963 , \19971 );
nand \U$11154 ( \19973 , \19949 , \19957 , \19972 );
xnor \U$11155 ( \19974 , \19973 , \9786 );
nor \U$11156 ( \19975 , \19942 , \19974 );
nand \U$11157 ( \19976 , \19877 , \19910 , \19975 );
and \U$11158 ( \19977 , \14272 , \9334 );
not \U$11159 ( \19978 , \14033 );
or \U$11160 ( \19979 , \10553 , \19978 );
not \U$11161 ( \19980 , \19979 );
or \U$11162 ( \19981 , \11357 , \14121 );
or \U$11163 ( \19982 , \9342 , \14117 );
nand \U$11164 ( \19983 , \19981 , \19982 );
nor \U$11165 ( \19984 , \19977 , \19980 , \19983 );
or \U$11166 ( \19985 , \12139 , \14005 );
or \U$11167 ( \19986 , \12141 , \14101 );
nand \U$11168 ( \19987 , \19985 , \19986 );
not \U$11169 ( \19988 , \9356 );
or \U$11170 ( \19989 , \19988 , \14012 );
or \U$11171 ( \19990 , \9354 , \14097 );
nand \U$11172 ( \19991 , \19989 , \19990 );
nor \U$11173 ( \19992 , \19987 , \19991 );
or \U$11174 ( \19993 , \9332 , \14161 );
nand \U$11175 ( \19994 , \19804 , \9361 );
nand \U$11176 ( \19995 , \19835 , \9338 );
nand \U$11177 ( \19996 , \9374 , \14076 );
and \U$11178 ( \19997 , \19993 , \19994 , \19995 , \19996 );
not \U$11179 ( \19998 , \19997 );
not \U$11180 ( \19999 , \19998 );
and \U$11181 ( \20000 , \14049 , \9366 );
and \U$11182 ( \20001 , \19808 , \9369 );
nor \U$11183 ( \20002 , \20000 , \20001 );
not \U$11184 ( \20003 , \11371 );
and \U$11185 ( \20004 , \20003 , \14054 );
and \U$11186 ( \20005 , \19814 , \9385 );
nor \U$11187 ( \20006 , \20004 , \20005 );
and \U$11188 ( \20007 , \19999 , \20002 , \20006 );
nand \U$11189 ( \20008 , \19984 , \19992 , \20007 );
xnor \U$11190 ( \20009 , RIb7b9608_246, \20008 );
not \U$11191 ( \20010 , \14125 );
or \U$11192 ( \20011 , \9611 , \20010 );
not \U$11193 ( \20012 , \14272 );
or \U$11194 ( \20013 , \9614 , \20012 );
not \U$11195 ( \20014 , \14121 );
and \U$11196 ( \20015 , \9606 , \20014 );
not \U$11197 ( \20016 , \14069 );
and \U$11198 ( \20017 , \9603 , \20016 );
nor \U$11199 ( \20018 , \20015 , \20017 );
nand \U$11200 ( \20019 , \20011 , \20013 , \20018 );
not \U$11201 ( \20020 , \20019 );
or \U$11202 ( \20021 , \13538 , \14135 );
or \U$11203 ( \20022 , \9597 , \14138 );
nand \U$11204 ( \20023 , \20021 , \20022 );
not \U$11205 ( \20024 , \9593 );
or \U$11206 ( \20025 , \20024 , \14012 );
or \U$11207 ( \20026 , \9588 , \13995 );
nand \U$11208 ( \20027 , \20025 , \20026 );
nor \U$11209 ( \20028 , \20023 , \20027 );
or \U$11210 ( \20029 , \11322 , \14079 );
nand \U$11211 ( \20030 , \19835 , \9636 );
nand \U$11212 ( \20031 , \19804 , \9639 );
nand \U$11213 ( \20032 , \9646 , \14076 );
and \U$11214 ( \20033 , \20029 , \20030 , \20031 , \20032 );
not \U$11215 ( \20034 , \20033 );
not \U$11216 ( \20035 , \20034 );
not \U$11217 ( \20036 , \9620 );
and \U$11218 ( \20037 , \20036 , \14054 );
and \U$11219 ( \20038 , \19814 , \9622 );
nor \U$11220 ( \20039 , \20037 , \20038 );
not \U$11221 ( \20040 , \9632 );
and \U$11222 ( \20041 , \20040 , \14049 );
and \U$11223 ( \20042 , \19808 , \9628 );
nor \U$11224 ( \20043 , \20041 , \20042 );
and \U$11225 ( \20044 , \20035 , \20039 , \20043 );
nand \U$11226 ( \20045 , \20020 , \20028 , \20044 );
xnor \U$11227 ( \20046 , RIb7af630_254, \20045 );
and \U$11228 ( \20047 , \14272 , \9265 );
not \U$11229 ( \20048 , \14033 );
or \U$11230 ( \20049 , \10415 , \20048 );
not \U$11231 ( \20050 , \20049 );
or \U$11232 ( \20051 , \11298 , \13998 );
or \U$11233 ( \20052 , \9273 , \14069 );
nand \U$11234 ( \20053 , \20051 , \20052 );
nor \U$11235 ( \20054 , \20047 , \20050 , \20053 );
or \U$11236 ( \20055 , \9282 , \14005 );
or \U$11237 ( \20056 , \11276 , \14101 );
nand \U$11238 ( \20057 , \20055 , \20056 );
not \U$11239 ( \20058 , \9289 );
or \U$11240 ( \20059 , \20058 , \14012 );
or \U$11241 ( \20060 , \9287 , \14097 );
nand \U$11242 ( \20061 , \20059 , \20060 );
nor \U$11243 ( \20062 , \20057 , \20061 );
or \U$11244 ( \20063 , \9263 , \14079 );
nand \U$11245 ( \20064 , \19804 , \9295 );
nand \U$11246 ( \20065 , \19835 , \9269 );
nand \U$11247 ( \20066 , \9307 , \14076 );
and \U$11248 ( \20067 , \20063 , \20064 , \20065 , \20066 );
not \U$11249 ( \20068 , \20067 );
not \U$11250 ( \20069 , \20068 );
and \U$11251 ( \20070 , \14049 , \9299 );
and \U$11252 ( \20071 , \19808 , \9302 );
nor \U$11253 ( \20072 , \20070 , \20071 );
and \U$11254 ( \20073 , \19814 , \9315 );
and \U$11255 ( \20074 , \9319 , \14054 );
nor \U$11256 ( \20075 , \20073 , \20074 );
and \U$11257 ( \20076 , \20069 , \20072 , \20075 );
nand \U$11258 ( \20077 , \20054 , \20062 , \20076 );
xnor \U$11259 ( \20078 , \20077 , \9327 );
and \U$11260 ( \20079 , \14272 , \9397 );
nand \U$11261 ( \20080 , \9444 , \14033 );
not \U$11262 ( \20081 , \20080 );
or \U$11263 ( \20082 , \10464 , \14201 );
or \U$11264 ( \20083 , \9405 , \14197 );
nand \U$11265 ( \20084 , \20082 , \20083 );
nor \U$11266 ( \20085 , \20079 , \20081 , \20084 );
or \U$11267 ( \20086 , \9415 , \14104 );
or \U$11268 ( \20087 , \10455 , \14017 );
nand \U$11269 ( \20088 , \20086 , \20087 );
not \U$11270 ( \20089 , \9421 );
or \U$11271 ( \20090 , \20089 , \14012 );
or \U$11272 ( \20091 , \9419 , \14183 );
nand \U$11273 ( \20092 , \20090 , \20091 );
nor \U$11274 ( \20093 , \20088 , \20092 );
or \U$11275 ( \20094 , \9395 , \14161 );
nand \U$11276 ( \20095 , \19804 , \9427 );
nand \U$11277 ( \20096 , \19835 , \9401 );
nand \U$11278 ( \20097 , \9440 , \14076 );
and \U$11279 ( \20098 , \20094 , \20095 , \20096 , \20097 );
not \U$11280 ( \20099 , \20098 );
not \U$11281 ( \20100 , \20099 );
and \U$11282 ( \20101 , \14049 , \9432 );
and \U$11283 ( \20102 , \19808 , \9435 );
nor \U$11284 ( \20103 , \20101 , \20102 );
and \U$11285 ( \20104 , \19814 , \9449 );
and \U$11286 ( \20105 , \9453 , \14054 );
nor \U$11287 ( \20106 , \20104 , \20105 );
and \U$11288 ( \20107 , \20100 , \20103 , \20106 );
nand \U$11289 ( \20108 , \20085 , \20093 , \20107 );
xnor \U$11290 ( \20109 , \20108 , \9460 );
nor \U$11291 ( \20110 , \20078 , \20109 );
nand \U$11292 ( \20111 , \20009 , \20046 , \20110 );
nor \U$11293 ( \20112 , \19976 , \20111 );
not \U$11294 ( \20113 , \14033 );
or \U$11295 ( \20114 , \9884 , \20113 );
not \U$11296 ( \20115 , \14272 );
or \U$11297 ( \20116 , \9887 , \20115 );
not \U$11298 ( \20117 , \14201 );
and \U$11299 ( \20118 , \9877 , \20117 );
not \U$11300 ( \20119 , \14117 );
and \U$11301 ( \20120 , \9874 , \20119 );
nor \U$11302 ( \20121 , \20118 , \20120 );
nand \U$11303 ( \20122 , \20114 , \20116 , \20121 );
not \U$11304 ( \20123 , \20122 );
or \U$11305 ( \20124 , \12178 , \14104 );
or \U$11306 ( \20125 , \9868 , \14017 );
nand \U$11307 ( \20126 , \20124 , \20125 );
not \U$11308 ( \20127 , \9864 );
or \U$11309 ( \20128 , \20127 , \14180 );
or \U$11310 ( \20129 , \9860 , \14183 );
nand \U$11311 ( \20130 , \20128 , \20129 );
nor \U$11312 ( \20131 , \20126 , \20130 );
or \U$11313 ( \20132 , \11718 , \14161 );
nand \U$11314 ( \20133 , \19835 , \9910 );
nand \U$11315 ( \20134 , \19804 , \9913 );
nand \U$11316 ( \20135 , \9920 , \14076 );
and \U$11317 ( \20136 , \20132 , \20133 , \20134 , \20135 );
not \U$11318 ( \20137 , \20136 );
not \U$11319 ( \20138 , \20137 );
not \U$11320 ( \20139 , \9895 );
and \U$11321 ( \20140 , \20139 , \14054 );
and \U$11322 ( \20141 , \19814 , \9897 );
nor \U$11323 ( \20142 , \20140 , \20141 );
not \U$11324 ( \20143 , \9906 );
and \U$11325 ( \20144 , \20143 , \14049 );
and \U$11326 ( \20145 , \19808 , \9902 );
nor \U$11327 ( \20146 , \20144 , \20145 );
and \U$11328 ( \20147 , \20138 , \20142 , \20146 );
nand \U$11329 ( \20148 , \20123 , \20131 , \20147 );
xnor \U$11330 ( \20149 , RIb7a0c48_261, \20148 );
not \U$11331 ( \20150 , \14033 );
or \U$11332 ( \20151 , \10018 , \20150 );
not \U$11333 ( \20152 , \14272 );
or \U$11334 ( \20153 , \10021 , \20152 );
not \U$11335 ( \20154 , \14121 );
and \U$11336 ( \20155 , \10012 , \20154 );
not \U$11337 ( \20156 , \14069 );
and \U$11338 ( \20157 , \10009 , \20156 );
nor \U$11339 ( \20158 , \20155 , \20157 );
nand \U$11340 ( \20159 , \20151 , \20153 , \20158 );
not \U$11341 ( \20160 , \20159 );
or \U$11342 ( \20161 , \9997 , \14005 );
or \U$11343 ( \20162 , \11666 , \14101 );
nand \U$11344 ( \20163 , \20161 , \20162 );
not \U$11345 ( \20164 , \10004 );
or \U$11346 ( \20165 , \20164 , \14012 );
or \U$11347 ( \20166 , \10002 , \14097 );
nand \U$11348 ( \20167 , \20165 , \20166 );
nor \U$11349 ( \20168 , \20163 , \20167 );
or \U$11350 ( \20169 , \11681 , \14079 );
nand \U$11351 ( \20170 , \19835 , \10043 );
nand \U$11352 ( \20171 , \19804 , \10041 );
nand \U$11353 ( \20172 , \10049 , \14091 );
and \U$11354 ( \20173 , \20169 , \20170 , \20171 , \20172 );
not \U$11355 ( \20174 , \20173 );
not \U$11356 ( \20175 , \20174 );
not \U$11357 ( \20176 , \12230 );
and \U$11358 ( \20177 , \20176 , \14054 );
and \U$11359 ( \20178 , \19814 , \10030 );
nor \U$11360 ( \20179 , \20177 , \20178 );
not \U$11361 ( \20180 , \11693 );
and \U$11362 ( \20181 , \20180 , \14049 );
and \U$11363 ( \20182 , \19808 , \10027 );
nor \U$11364 ( \20183 , \20181 , \20182 );
and \U$11365 ( \20184 , \20175 , \20179 , \20183 );
nand \U$11366 ( \20185 , \20160 , \20168 , \20184 );
xnor \U$11367 ( \20186 , RIb7af540_256, \20185 );
nand \U$11368 ( \20187 , \9542 , \14125 );
nand \U$11369 ( \20188 , \9545 , \14272 );
not \U$11370 ( \20189 , \14201 );
and \U$11371 ( \20190 , \9536 , \20189 );
not \U$11372 ( \20191 , \14117 );
and \U$11373 ( \20192 , \9533 , \20191 );
nor \U$11374 ( \20193 , \20190 , \20192 );
nand \U$11375 ( \20194 , \20187 , \20188 , \20193 );
not \U$11376 ( \20195 , \20194 );
or \U$11377 ( \20196 , \13658 , \14104 );
or \U$11378 ( \20197 , \9527 , \14017 );
nand \U$11379 ( \20198 , \20196 , \20197 );
not \U$11380 ( \20199 , \9523 );
or \U$11381 ( \20200 , \20199 , \14012 );
or \U$11382 ( \20201 , \9519 , \14183 );
nand \U$11383 ( \20202 , \20200 , \20201 );
nor \U$11384 ( \20203 , \20198 , \20202 );
or \U$11385 ( \20204 , \11589 , \14079 );
nand \U$11386 ( \20205 , \19835 , \9568 );
nand \U$11387 ( \20206 , \19804 , \9571 );
nand \U$11388 ( \20207 , \9578 , \14091 );
and \U$11389 ( \20208 , \20204 , \20205 , \20206 , \20207 );
not \U$11390 ( \20209 , \20208 );
not \U$11391 ( \20210 , \20209 );
and \U$11392 ( \20211 , \19814 , \9554 );
and \U$11393 ( \20212 , \9551 , \14054 );
nor \U$11394 ( \20213 , \20211 , \20212 );
and \U$11395 ( \20214 , \19808 , \9560 );
and \U$11396 ( \20215 , \9563 , \14049 );
nor \U$11397 ( \20216 , \20214 , \20215 );
and \U$11398 ( \20217 , \20210 , \20213 , \20216 );
nand \U$11399 ( \20218 , \20195 , \20203 , \20217 );
xnor \U$11400 ( \20219 , \20218 , \9585 );
nand \U$11401 ( \20220 , \9936 , \14033 );
nand \U$11402 ( \20221 , \9939 , \14272 );
not \U$11403 ( \20222 , \13998 );
and \U$11404 ( \20223 , \9932 , \20222 );
not \U$11405 ( \20224 , \14197 );
and \U$11406 ( \20225 , \9929 , \20224 );
nor \U$11407 ( \20226 , \20223 , \20225 );
nand \U$11408 ( \20227 , \20220 , \20221 , \20226 );
not \U$11409 ( \20228 , \20227 );
or \U$11410 ( \20229 , \9948 , \14135 );
or \U$11411 ( \20230 , \13143 , \14138 );
nand \U$11412 ( \20231 , \20229 , \20230 );
not \U$11413 ( \20232 , \9954 );
or \U$11414 ( \20233 , \20232 , \14180 );
or \U$11415 ( \20234 , \9952 , \13995 );
nand \U$11416 ( \20235 , \20233 , \20234 );
nor \U$11417 ( \20236 , \20231 , \20235 );
or \U$11418 ( \20237 , \11633 , \14161 );
nand \U$11419 ( \20238 , \19835 , \9977 );
nand \U$11420 ( \20239 , \19804 , \9975 );
nand \U$11421 ( \20240 , \9984 , \14091 );
and \U$11422 ( \20241 , \20237 , \20238 , \20239 , \20240 );
not \U$11423 ( \20242 , \20241 );
not \U$11424 ( \20243 , \20242 );
and \U$11425 ( \20244 , \19814 , \9965 );
and \U$11426 ( \20245 , \9968 , \14054 );
nor \U$11427 ( \20246 , \20244 , \20245 );
and \U$11428 ( \20247 , \19808 , \10709 );
and \U$11429 ( \20248 , \9959 , \14049 );
nor \U$11430 ( \20249 , \20247 , \20248 );
and \U$11431 ( \20250 , \20243 , \20246 , \20249 );
nand \U$11432 ( \20251 , \20228 , \20236 , \20250 );
xnor \U$11433 ( \20252 , \20251 , \9990 );
nor \U$11434 ( \20253 , \20219 , \20252 );
nand \U$11435 ( \20254 , \20149 , \20186 , \20253 );
not \U$11436 ( \20255 , \20254 );
not \U$11437 ( \20256 , \14125 );
or \U$11438 ( \20257 , \9814 , \20256 );
not \U$11439 ( \20258 , \14272 );
or \U$11440 ( \20259 , \9817 , \20258 );
not \U$11441 ( \20260 , \13998 );
and \U$11442 ( \20261 , \9808 , \20260 );
not \U$11443 ( \20262 , \14197 );
and \U$11444 ( \20263 , \9805 , \20262 );
nor \U$11445 ( \20264 , \20261 , \20263 );
nand \U$11446 ( \20265 , \20257 , \20259 , \20264 );
not \U$11447 ( \20266 , \20265 );
or \U$11448 ( \20267 , \11494 , \14135 );
or \U$11449 ( \20268 , \9798 , \14138 );
nand \U$11450 ( \20269 , \20267 , \20268 );
not \U$11451 ( \20270 , \9794 );
or \U$11452 ( \20271 , \20270 , \14180 );
or \U$11453 ( \20272 , \9791 , \13995 );
nand \U$11454 ( \20273 , \20271 , \20272 );
nor \U$11455 ( \20274 , \20269 , \20273 );
or \U$11456 ( \20275 , \11505 , \14079 );
nand \U$11457 ( \20276 , \19835 , \9839 );
nand \U$11458 ( \20277 , \19804 , \9842 );
nand \U$11459 ( \20278 , \9850 , \14091 );
and \U$11460 ( \20279 , \20275 , \20276 , \20277 , \20278 );
not \U$11461 ( \20280 , \20279 );
not \U$11462 ( \20281 , \20280 );
not \U$11463 ( \20282 , \9823 );
and \U$11464 ( \20283 , \20282 , \14054 );
and \U$11465 ( \20284 , \19814 , \9826 );
nor \U$11466 ( \20285 , \20283 , \20284 );
not \U$11467 ( \20286 , \9834 );
and \U$11468 ( \20287 , \20286 , \14049 );
and \U$11469 ( \20288 , \19808 , \9830 );
nor \U$11470 ( \20289 , \20287 , \20288 );
and \U$11471 ( \20290 , \20281 , \20285 , \20289 );
nand \U$11472 ( \20291 , \20266 , \20274 , \20290 );
xnor \U$11473 ( \20292 , \20291 , \9857 );
and \U$11474 ( \20293 , \14272 , \8843 );
not \U$11475 ( \20294 , \14033 );
or \U$11476 ( \20295 , \10775 , \20294 );
not \U$11477 ( \20296 , \20295 );
or \U$11478 ( \20297 , \11533 , \13998 );
or \U$11479 ( \20298 , \8861 , \14069 );
nand \U$11480 ( \20299 , \20297 , \20298 );
nor \U$11481 ( \20300 , \20293 , \20296 , \20299 );
or \U$11482 ( \20301 , \8882 , \14005 );
or \U$11483 ( \20302 , \12351 , \14101 );
nand \U$11484 ( \20303 , \20301 , \20302 );
not \U$11485 ( \20304 , \8896 );
or \U$11486 ( \20305 , \20304 , \14180 );
or \U$11487 ( \20306 , \8894 , \14097 );
nand \U$11488 ( \20307 , \20305 , \20306 );
nor \U$11489 ( \20308 , \20303 , \20307 );
or \U$11490 ( \20309 , \8828 , \14161 );
nand \U$11491 ( \20310 , \19804 , \8904 );
nand \U$11492 ( \20311 , \19835 , \8852 );
not \U$11493 ( \20312 , \14091 );
or \U$11494 ( \20313 , \11565 , \20312 );
and \U$11495 ( \20314 , \20309 , \20310 , \20311 , \20313 );
not \U$11496 ( \20315 , \20314 );
not \U$11497 ( \20316 , \20315 );
and \U$11498 ( \20317 , \14049 , \8921 );
and \U$11499 ( \20318 , \19808 , \8927 );
nor \U$11500 ( \20319 , \20317 , \20318 );
not \U$11501 ( \20320 , \14573 );
and \U$11502 ( \20321 , \20320 , \14054 );
and \U$11503 ( \20322 , \19814 , \8947 );
nor \U$11504 ( \20323 , \20321 , \20322 );
and \U$11505 ( \20324 , \20316 , \20319 , \20323 );
nand \U$11506 ( \20325 , \20300 , \20308 , \20324 );
xnor \U$11507 ( \20326 , \20325 , \8964 );
nor \U$11508 ( \20327 , \20292 , \20326 );
and \U$11509 ( \20328 , \14272 , \9049 );
not \U$11510 ( \20329 , \14125 );
or \U$11511 ( \20330 , \10859 , \20329 );
not \U$11512 ( \20331 , \20330 );
or \U$11513 ( \20332 , \9086 , \14201 );
or \U$11514 ( \20333 , \9058 , \14197 );
nand \U$11515 ( \20334 , \20332 , \20333 );
nor \U$11516 ( \20335 , \20328 , \20331 , \20334 );
or \U$11517 ( \20336 , \9068 , \14104 );
or \U$11518 ( \20337 , \11458 , \14017 );
nand \U$11519 ( \20338 , \20336 , \20337 );
not \U$11520 ( \20339 , \9075 );
or \U$11521 ( \20340 , \20339 , \14180 );
or \U$11522 ( \20341 , \9073 , \14183 );
nand \U$11523 ( \20342 , \20340 , \20341 );
nor \U$11524 ( \20343 , \20338 , \20342 );
or \U$11525 ( \20344 , \9047 , \14161 );
nand \U$11526 ( \20345 , \19804 , \9081 );
nand \U$11527 ( \20346 , \19835 , \9054 );
nand \U$11528 ( \20347 , \9098 , \14091 );
and \U$11529 ( \20348 , \20344 , \20345 , \20346 , \20347 );
not \U$11530 ( \20349 , \20348 );
not \U$11531 ( \20350 , \20349 );
and \U$11532 ( \20351 , \14049 , \9089 );
and \U$11533 ( \20352 , \19808 , \9093 );
nor \U$11534 ( \20353 , \20351 , \20352 );
not \U$11535 ( \20354 , \11471 );
and \U$11536 ( \20355 , \20354 , \14054 );
and \U$11537 ( \20356 , \19814 , \9107 );
nor \U$11538 ( \20357 , \20355 , \20356 );
and \U$11539 ( \20358 , \20350 , \20353 , \20357 );
nand \U$11540 ( \20359 , \20335 , \20343 , \20358 );
xnor \U$11541 ( \20360 , \20359 , \9119 );
and \U$11542 ( \20361 , \14272 , \9124 );
not \U$11543 ( \20362 , \14125 );
or \U$11544 ( \20363 , \10901 , \20362 );
not \U$11545 ( \20364 , \20363 );
or \U$11546 ( \20365 , \11436 , \14121 );
or \U$11547 ( \20366 , \9133 , \14117 );
nand \U$11548 ( \20367 , \20365 , \20366 );
nor \U$11549 ( \20368 , \20361 , \20364 , \20367 );
or \U$11550 ( \20369 , \9143 , \14135 );
or \U$11551 ( \20370 , \11416 , \14138 );
nand \U$11552 ( \20371 , \20369 , \20370 );
not \U$11553 ( \20372 , \9150 );
or \U$11554 ( \20373 , \20372 , \14180 );
or \U$11555 ( \20374 , \9148 , \13995 );
nand \U$11556 ( \20375 , \20373 , \20374 );
nor \U$11557 ( \20376 , \20371 , \20375 );
or \U$11558 ( \20377 , \9122 , \14079 );
nand \U$11559 ( \20378 , \19804 , \9155 );
nand \U$11560 ( \20379 , \19835 , \9129 );
nand \U$11561 ( \20380 , \9168 , \14076 );
and \U$11562 ( \20381 , \20377 , \20378 , \20379 , \20380 );
not \U$11563 ( \20382 , \20381 );
not \U$11564 ( \20383 , \20382 );
and \U$11565 ( \20384 , \14049 , \9159 );
and \U$11566 ( \20385 , \19808 , \9163 );
nor \U$11567 ( \20386 , \20384 , \20385 );
not \U$11568 ( \20387 , \11429 );
and \U$11569 ( \20388 , \20387 , \14054 );
and \U$11570 ( \20389 , \19814 , \9176 );
nor \U$11571 ( \20390 , \20388 , \20389 );
and \U$11572 ( \20391 , \20383 , \20386 , \20390 );
nand \U$11573 ( \20392 , \20368 , \20376 , \20391 );
xnor \U$11574 ( \20393 , \20392 , \9188 );
nor \U$11575 ( \20394 , \20360 , \20393 );
and \U$11576 ( \20395 , \20255 , \20327 , \20394 );
nand \U$11577 ( \20396 , \19844 , \20112 , \20395 );
not \U$11578 ( \20397 , \20396 );
nor \U$11579 ( \20398 , \19802 , \20397 );
buf \U$11580 ( \20399 , RIea91330_6888);
buf \U$11581 ( \20400 , \13927 );
buf \U$11582 ( \20401 , \12456 );
buf \U$11583 ( \20402 , \12458 );
not \U$11584 ( \20403 , \20402 );
not \U$11585 ( \20404 , \20403 );
and \U$11586 ( \20405 , \20401 , \20404 );
and \U$11587 ( \20406 , \20400 , \20405 );
and \U$11588 ( \20407 , \20399 , \20406 );
buf \U$11589 ( \20408 , \20407 );
not \U$11590 ( \20409 , \20408 );
buf \U$11591 ( \20410 , \8835 );
buf \U$11592 ( \20411 , \20403 );
or \U$11593 ( \20412 , \20410 , \20411 );
xor \U$11594 ( \20413 , \20401 , \20404 );
buf \U$11595 ( \20414 , \20413 );
xor \U$11596 ( \20415 , \20400 , \20405 );
buf \U$11597 ( \20416 , \20415 );
or \U$11598 ( \20417 , \20414 , \20416 );
or \U$11599 ( \20418 , \20412 , \20417 );
xor \U$11600 ( \20419 , \20399 , \20406 );
buf \U$11601 ( \20420 , \20419 );
nand \U$11602 ( \20421 , \20418 , \20420 );
nand \U$11603 ( \20422 , \20409 , \20421 );
not \U$11604 ( \20423 , \20397 );
or \U$11605 ( \20424 , \20422 , \20423 );
not \U$11606 ( \20425 , \20424 );
not \U$11607 ( \20426 , \20422 );
not \U$11608 ( \20427 , \20397 );
or \U$11609 ( \20428 , \20426 , \20427 );
not \U$11610 ( \20429 , \20428 );
or \U$11611 ( \20430 , \20425 , \20429 );
not \U$11612 ( \20431 , \20430 );
not \U$11613 ( \20432 , \20431 );
and \U$11614 ( \20433 , \13956 , \20432 );
or \U$11615 ( \20434 , \20398 , \20433 );
not \U$11616 ( \20435 , \9509 );
and \U$11617 ( \20436 , \20435 , \12552 );
not \U$11618 ( \20437 , \12498 );
not \U$11619 ( \20438 , \20437 );
and \U$11620 ( \20439 , \20438 , \10120 );
nor \U$11621 ( \20440 , \20436 , \20439 );
not \U$11622 ( \20441 , \9506 );
and \U$11623 ( \20442 , \20441 , \12575 );
buf \U$11624 ( \20443 , \12546 );
and \U$11625 ( \20444 , \20443 , \10976 );
nor \U$11626 ( \20445 , \20442 , \20444 );
nand \U$11627 ( \20446 , \20440 , \20445 );
not \U$11628 ( \20447 , \20446 );
not \U$11629 ( \20448 , \9494 );
buf \U$11630 ( \20449 , \12569 );
and \U$11631 ( \20450 , \20448 , \20449 );
not \U$11632 ( \20451 , \12565 );
not \U$11633 ( \20452 , \20451 );
and \U$11634 ( \20453 , \20452 , \12513 );
nor \U$11635 ( \20454 , \20450 , \20453 );
not \U$11636 ( \20455 , \9500 );
buf \U$11637 ( \20456 , \12535 );
and \U$11638 ( \20457 , \20455 , \20456 );
buf \U$11639 ( \20458 , \12579 );
and \U$11640 ( \20459 , \20458 , \10085 );
nor \U$11641 ( \20460 , \20457 , \20459 );
and \U$11642 ( \20461 , \20447 , \20454 , \20460 );
not \U$11643 ( \20462 , \9463 );
buf \U$11644 ( \20463 , \12521 );
and \U$11645 ( \20464 , \20462 , \20463 );
buf \U$11646 ( \20465 , \12502 );
and \U$11647 ( \20466 , \20465 , \9468 );
nor \U$11648 ( \20467 , \20464 , \20466 );
not \U$11649 ( \20468 , \9471 );
and \U$11650 ( \20469 , \20468 , \12512 );
buf \U$11651 ( \20470 , \12508 );
and \U$11652 ( \20471 , \20470 , \9476 );
nor \U$11653 ( \20472 , \20469 , \20471 );
nand \U$11654 ( \20473 , \20467 , \20472 );
not \U$11655 ( \20474 , \20473 );
not \U$11656 ( \20475 , \9480 );
and \U$11657 ( \20476 , \20475 , \12531 );
buf \U$11658 ( \20477 , \12542 );
and \U$11659 ( \20478 , \20477 , \12557 );
nor \U$11660 ( \20479 , \20476 , \20478 );
not \U$11661 ( \20480 , \9487 );
buf \U$11662 ( \20481 , \12556 );
and \U$11663 ( \20482 , \20480 , \20481 );
buf \U$11664 ( \20483 , \12525 );
and \U$11665 ( \20484 , \20483 , \10168 );
nor \U$11666 ( \20485 , \20482 , \20484 );
and \U$11667 ( \20486 , \20474 , \20479 , \20485 );
nand \U$11668 ( \20487 , \20461 , \20486 );
not \U$11669 ( \20488 , \20487 );
not \U$11670 ( \20489 , \11067 );
and \U$11671 ( \20490 , \20489 , \12575 );
and \U$11672 ( \20491 , \20458 , \9034 );
nor \U$11673 ( \20492 , \20490 , \20491 );
not \U$11674 ( \20493 , \11060 );
and \U$11675 ( \20494 , \20493 , \20452 );
and \U$11676 ( \20495 , \20456 , \9014 );
nor \U$11677 ( \20496 , \20494 , \20495 );
nand \U$11678 ( \20497 , \20492 , \20496 );
not \U$11679 ( \20498 , \20497 );
not \U$11680 ( \20499 , \11036 );
and \U$11681 ( \20500 , \20499 , \12597 );
and \U$11682 ( \20501 , \20481 , \8966 );
nor \U$11683 ( \20502 , \20500 , \20501 );
not \U$11684 ( \20503 , \8977 );
and \U$11685 ( \20504 , \20503 , \20483 );
and \U$11686 ( \20505 , \20449 , \9006 );
nor \U$11687 ( \20506 , \20504 , \20505 );
and \U$11688 ( \20507 , \20498 , \20502 , \20506 );
and \U$11689 ( \20508 , \20470 , \9009 );
and \U$11690 ( \20509 , \8979 , \20443 );
nor \U$11691 ( \20510 , \20508 , \20509 );
and \U$11692 ( \20511 , \20477 , \8970 );
and \U$11693 ( \20512 , \9025 , \12531 );
nor \U$11694 ( \20513 , \20511 , \20512 );
nand \U$11695 ( \20514 , \20510 , \20513 );
not \U$11696 ( \20515 , \20514 );
not \U$11697 ( \20516 , \11046 );
and \U$11698 ( \20517 , \20516 , \20463 );
and \U$11699 ( \20518 , \20465 , \8990 );
nor \U$11700 ( \20519 , \20517 , \20518 );
not \U$11701 ( \20520 , \8997 );
and \U$11702 ( \20521 , \20520 , \12512 );
and \U$11703 ( \20522 , \20438 , \8999 );
nor \U$11704 ( \20523 , \20521 , \20522 );
and \U$11705 ( \20524 , \20515 , \20519 , \20523 );
nand \U$11706 ( \20525 , \20507 , \20524 );
xnor \U$11707 ( \20526 , RIb7b94a0_249, \20525 );
and \U$11708 ( \20527 , \20458 , \9251 );
and \U$11709 ( \20528 , \9247 , \12575 );
nor \U$11710 ( \20529 , \20527 , \20528 );
and \U$11711 ( \20530 , \20456 , \9233 );
and \U$11712 ( \20531 , \9230 , \20452 );
nor \U$11713 ( \20532 , \20530 , \20531 );
nand \U$11714 ( \20533 , \20529 , \20532 );
not \U$11715 ( \20534 , \20533 );
not \U$11716 ( \20535 , \11093 );
and \U$11717 ( \20536 , \20535 , \12597 );
and \U$11718 ( \20537 , \20481 , \9196 );
nor \U$11719 ( \20538 , \20536 , \20537 );
not \U$11720 ( \20539 , \9205 );
and \U$11721 ( \20540 , \20539 , \20483 );
and \U$11722 ( \20541 , \20449 , \9225 );
nor \U$11723 ( \20542 , \20540 , \20541 );
and \U$11724 ( \20543 , \20534 , \20538 , \20542 );
and \U$11725 ( \20544 , \20470 , \9228 );
and \U$11726 ( \20545 , \9200 , \20443 );
nor \U$11727 ( \20546 , \20544 , \20545 );
and \U$11728 ( \20547 , \20477 , \9193 );
and \U$11729 ( \20548 , \9242 , \12531 );
nor \U$11730 ( \20549 , \20547 , \20548 );
nand \U$11731 ( \20550 , \20546 , \20549 );
not \U$11732 ( \20551 , \20550 );
not \U$11733 ( \20552 , \11101 );
and \U$11734 ( \20553 , \20552 , \20463 );
and \U$11735 ( \20554 , \20465 , \9212 );
nor \U$11736 ( \20555 , \20553 , \20554 );
not \U$11737 ( \20556 , \9217 );
and \U$11738 ( \20557 , \20556 , \12512 );
and \U$11739 ( \20558 , \20438 , \9219 );
nor \U$11740 ( \20559 , \20557 , \20558 );
and \U$11741 ( \20560 , \20551 , \20555 , \20559 );
nand \U$11742 ( \20561 , \20543 , \20560 );
xnor \U$11743 ( \20562 , RIb7b9518_248, \20561 );
and \U$11744 ( \20563 , \20477 , \9710 );
and \U$11745 ( \20564 , \9713 , \12531 );
nor \U$11746 ( \20565 , \20563 , \20564 );
and \U$11747 ( \20566 , \20443 , \9706 );
and \U$11748 ( \20567 , \9701 , \20470 );
nor \U$11749 ( \20568 , \20566 , \20567 );
nand \U$11750 ( \20569 , \20565 , \20568 );
not \U$11751 ( \20570 , \20569 );
and \U$11752 ( \20571 , \20458 , \9695 );
and \U$11753 ( \20572 , \9692 , \12575 );
nor \U$11754 ( \20573 , \20571 , \20572 );
and \U$11755 ( \20574 , \20456 , \9690 );
and \U$11756 ( \20575 , \9687 , \20452 );
nor \U$11757 ( \20576 , \20574 , \20575 );
and \U$11758 ( \20577 , \20570 , \20573 , \20576 );
and \U$11759 ( \20578 , \20438 , \9682 );
and \U$11760 ( \20579 , \9679 , \12512 );
nor \U$11761 ( \20580 , \20578 , \20579 );
and \U$11762 ( \20581 , \20465 , \9675 );
and \U$11763 ( \20582 , \9672 , \20463 );
nor \U$11764 ( \20583 , \20581 , \20582 );
nand \U$11765 ( \20584 , \20580 , \20583 );
not \U$11766 ( \20585 , \20584 );
and \U$11767 ( \20586 , \20483 , \9656 );
and \U$11768 ( \20587 , \9660 , \20449 );
nor \U$11769 ( \20588 , \20586 , \20587 );
and \U$11770 ( \20589 , \20481 , \9664 );
and \U$11771 ( \20590 , \9667 , \12597 );
nor \U$11772 ( \20591 , \20589 , \20590 );
and \U$11773 ( \20592 , \20585 , \20588 , \20591 );
nand \U$11774 ( \20593 , \20577 , \20592 );
xnor \U$11775 ( \20594 , \20593 , \9719 );
and \U$11776 ( \20595 , \20477 , \9776 );
and \U$11777 ( \20596 , \9779 , \12531 );
nor \U$11778 ( \20597 , \20595 , \20596 );
and \U$11779 ( \20598 , \20443 , \9772 );
and \U$11780 ( \20599 , \9769 , \20470 );
nor \U$11781 ( \20600 , \20598 , \20599 );
nand \U$11782 ( \20601 , \20597 , \20600 );
not \U$11783 ( \20602 , \20601 );
and \U$11784 ( \20603 , \20458 , \9763 );
and \U$11785 ( \20604 , \9759 , \12575 );
nor \U$11786 ( \20605 , \20603 , \20604 );
and \U$11787 ( \20606 , \20456 , \9755 );
and \U$11788 ( \20607 , \9752 , \20452 );
nor \U$11789 ( \20608 , \20606 , \20607 );
and \U$11790 ( \20609 , \20602 , \20605 , \20608 );
not \U$11791 ( \20610 , \9745 );
and \U$11792 ( \20611 , \20610 , \12512 );
and \U$11793 ( \20612 , \20438 , \9747 );
nor \U$11794 ( \20613 , \20611 , \20612 );
not \U$11795 ( \20614 , \11876 );
and \U$11796 ( \20615 , \20614 , \20463 );
and \U$11797 ( \20616 , \20465 , \9739 );
nor \U$11798 ( \20617 , \20615 , \20616 );
nand \U$11799 ( \20618 , \20613 , \20617 );
not \U$11800 ( \20619 , \20618 );
not \U$11801 ( \20620 , \9725 );
and \U$11802 ( \20621 , \20620 , \20449 );
and \U$11803 ( \20622 , \20483 , \9721 );
nor \U$11804 ( \20623 , \20621 , \20622 );
not \U$11805 ( \20624 , \9732 );
and \U$11806 ( \20625 , \20624 , \12552 );
and \U$11807 ( \20626 , \20481 , \9728 );
nor \U$11808 ( \20627 , \20625 , \20626 );
and \U$11809 ( \20628 , \20619 , \20623 , \20627 );
nand \U$11810 ( \20629 , \20609 , \20628 );
xnor \U$11811 ( \20630 , \20629 , \9786 );
nor \U$11812 ( \20631 , \20594 , \20630 );
nand \U$11813 ( \20632 , \20526 , \20562 , \20631 );
not \U$11814 ( \20633 , \20632 );
not \U$11815 ( \20634 , \11293 );
and \U$11816 ( \20635 , \20634 , \12575 );
and \U$11817 ( \20636 , \20458 , \9319 );
nor \U$11818 ( \20637 , \20635 , \20636 );
not \U$11819 ( \20638 , \11288 );
and \U$11820 ( \20639 , \20638 , \20452 );
and \U$11821 ( \20640 , \20456 , \9302 );
nor \U$11822 ( \20641 , \20639 , \20640 );
nand \U$11823 ( \20642 , \20637 , \20641 );
not \U$11824 ( \20643 , \20642 );
not \U$11825 ( \20644 , \11270 );
and \U$11826 ( \20645 , \20644 , \12597 );
and \U$11827 ( \20646 , \20481 , \9262 );
nor \U$11828 ( \20647 , \20645 , \20646 );
not \U$11829 ( \20648 , \9270 );
and \U$11830 ( \20649 , \20648 , \20483 );
and \U$11831 ( \20650 , \20449 , \9295 );
nor \U$11832 ( \20651 , \20649 , \20650 );
and \U$11833 ( \20652 , \20643 , \20647 , \20651 );
not \U$11834 ( \20653 , \9273 );
and \U$11835 ( \20654 , \20653 , \20443 );
and \U$11836 ( \20655 , \20470 , \9297 );
nor \U$11837 ( \20656 , \20654 , \20655 );
not \U$11838 ( \20657 , \10415 );
and \U$11839 ( \20658 , \20657 , \12531 );
and \U$11840 ( \20659 , \20477 , \9265 );
nor \U$11841 ( \20660 , \20658 , \20659 );
nand \U$11842 ( \20661 , \20656 , \20660 );
not \U$11843 ( \20662 , \20661 );
not \U$11844 ( \20663 , \11276 );
and \U$11845 ( \20664 , \20663 , \20463 );
and \U$11846 ( \20665 , \20465 , \9281 );
nor \U$11847 ( \20666 , \20664 , \20665 );
not \U$11848 ( \20667 , \9287 );
and \U$11849 ( \20668 , \20667 , \12512 );
and \U$11850 ( \20669 , \20438 , \9289 );
nor \U$11851 ( \20670 , \20668 , \20669 );
and \U$11852 ( \20671 , \20662 , \20666 , \20670 );
nand \U$11853 ( \20672 , \20652 , \20671 );
xnor \U$11854 ( \20673 , \20672 , \9327 );
not \U$11855 ( \20674 , \11250 );
and \U$11856 ( \20675 , \20674 , \12575 );
and \U$11857 ( \20676 , \20458 , \9453 );
nor \U$11858 ( \20677 , \20675 , \20676 );
not \U$11859 ( \20678 , \11245 );
and \U$11860 ( \20679 , \20678 , \20452 );
and \U$11861 ( \20680 , \20456 , \9435 );
nor \U$11862 ( \20681 , \20679 , \20680 );
nand \U$11863 ( \20682 , \20677 , \20681 );
not \U$11864 ( \20683 , \20682 );
not \U$11865 ( \20684 , \11230 );
and \U$11866 ( \20685 , \20684 , \12597 );
and \U$11867 ( \20686 , \20481 , \9394 );
nor \U$11868 ( \20687 , \20685 , \20686 );
not \U$11869 ( \20688 , \9402 );
and \U$11870 ( \20689 , \20688 , \20483 );
and \U$11871 ( \20690 , \20449 , \9427 );
nor \U$11872 ( \20691 , \20689 , \20690 );
and \U$11873 ( \20692 , \20683 , \20687 , \20691 );
not \U$11874 ( \20693 , \9405 );
and \U$11875 ( \20694 , \20693 , \20443 );
and \U$11876 ( \20695 , \20470 , \9430 );
nor \U$11877 ( \20696 , \20694 , \20695 );
not \U$11878 ( \20697 , \10462 );
and \U$11879 ( \20698 , \20697 , \12531 );
and \U$11880 ( \20699 , \20477 , \9397 );
nor \U$11881 ( \20700 , \20698 , \20699 );
nand \U$11882 ( \20701 , \20696 , \20700 );
not \U$11883 ( \20702 , \20701 );
not \U$11884 ( \20703 , \10455 );
and \U$11885 ( \20704 , \20703 , \20463 );
and \U$11886 ( \20705 , \20465 , \9414 );
nor \U$11887 ( \20706 , \20704 , \20705 );
not \U$11888 ( \20707 , \9419 );
and \U$11889 ( \20708 , \20707 , \12512 );
and \U$11890 ( \20709 , \20438 , \9421 );
nor \U$11891 ( \20710 , \20708 , \20709 );
and \U$11892 ( \20711 , \20702 , \20706 , \20710 );
nand \U$11893 ( \20712 , \20692 , \20711 );
xnor \U$11894 ( \20713 , \20712 , \9460 );
nor \U$11895 ( \20714 , \20673 , \20713 );
not \U$11896 ( \20715 , \9632 );
and \U$11897 ( \20716 , \20715 , \20452 );
and \U$11898 ( \20717 , \20456 , \9628 );
nor \U$11899 ( \20718 , \20716 , \20717 );
not \U$11900 ( \20719 , \9625 );
and \U$11901 ( \20720 , \20719 , \12575 );
and \U$11902 ( \20721 , \20458 , \9619 );
nor \U$11903 ( \20722 , \20720 , \20721 );
nand \U$11904 ( \20723 , \20718 , \20722 );
not \U$11905 ( \20724 , \20723 );
not \U$11906 ( \20725 , \9640 );
and \U$11907 ( \20726 , \20725 , \20449 );
and \U$11908 ( \20727 , \20483 , \9636 );
nor \U$11909 ( \20728 , \20726 , \20727 );
not \U$11910 ( \20729 , \9647 );
and \U$11911 ( \20730 , \20729 , \12552 );
and \U$11912 ( \20731 , \20481 , \9643 );
nor \U$11913 ( \20732 , \20730 , \20731 );
and \U$11914 ( \20733 , \20724 , \20728 , \20732 );
not \U$11915 ( \20734 , \9611 );
and \U$11916 ( \20735 , \20734 , \12531 );
and \U$11917 ( \20736 , \20477 , \9613 );
nor \U$11918 ( \20737 , \20735 , \20736 );
not \U$11919 ( \20738 , \9607 );
and \U$11920 ( \20739 , \20738 , \20470 );
and \U$11921 ( \20740 , \20443 , \9603 );
nor \U$11922 ( \20741 , \20739 , \20740 );
nand \U$11923 ( \20742 , \20737 , \20741 );
not \U$11924 ( \20743 , \20742 );
not \U$11925 ( \20744 , \9597 );
and \U$11926 ( \20745 , \20744 , \20463 );
and \U$11927 ( \20746 , \20465 , \9600 );
nor \U$11928 ( \20747 , \20745 , \20746 );
not \U$11929 ( \20748 , \9588 );
and \U$11930 ( \20749 , \20748 , \12512 );
and \U$11931 ( \20750 , \20438 , \9593 );
nor \U$11932 ( \20751 , \20749 , \20750 );
and \U$11933 ( \20752 , \20743 , \20747 , \20751 );
nand \U$11934 ( \20753 , \20733 , \20752 );
xnor \U$11935 ( \20754 , \20753 , \9653 );
not \U$11936 ( \20755 , \12874 );
and \U$11937 ( \20756 , \20755 , \12575 );
and \U$11938 ( \20757 , \20458 , \9377 );
nor \U$11939 ( \20758 , \20756 , \20757 );
not \U$11940 ( \20759 , \11365 );
and \U$11941 ( \20760 , \20759 , \20452 );
and \U$11942 ( \20761 , \20456 , \9369 );
nor \U$11943 ( \20762 , \20760 , \20761 );
nand \U$11944 ( \20763 , \20758 , \20762 );
not \U$11945 ( \20764 , \20763 );
not \U$11946 ( \20765 , \11393 );
and \U$11947 ( \20766 , \20765 , \12552 );
and \U$11948 ( \20767 , \20481 , \9331 );
nor \U$11949 ( \20768 , \20766 , \20767 );
not \U$11950 ( \20769 , \9339 );
and \U$11951 ( \20770 , \20769 , \20483 );
and \U$11952 ( \20771 , \20449 , \9361 );
nor \U$11953 ( \20772 , \20770 , \20771 );
and \U$11954 ( \20773 , \20764 , \20768 , \20772 );
not \U$11955 ( \20774 , \9342 );
and \U$11956 ( \20775 , \20774 , \20443 );
and \U$11957 ( \20776 , \20470 , \9364 );
nor \U$11958 ( \20777 , \20775 , \20776 );
not \U$11959 ( \20778 , \10553 );
and \U$11960 ( \20779 , \20778 , \12531 );
and \U$11961 ( \20780 , \20477 , \9334 );
nor \U$11962 ( \20781 , \20779 , \20780 );
nand \U$11963 ( \20782 , \20777 , \20781 );
not \U$11964 ( \20783 , \20782 );
not \U$11965 ( \20784 , \12141 );
and \U$11966 ( \20785 , \20784 , \20463 );
and \U$11967 ( \20786 , \20465 , \9348 );
nor \U$11968 ( \20787 , \20785 , \20786 );
not \U$11969 ( \20788 , \9354 );
and \U$11970 ( \20789 , \20788 , \12512 );
and \U$11971 ( \20790 , \20438 , \9356 );
nor \U$11972 ( \20791 , \20789 , \20790 );
and \U$11973 ( \20792 , \20783 , \20787 , \20791 );
nand \U$11974 ( \20793 , \20773 , \20792 );
xnor \U$11975 ( \20794 , \20793 , \9392 );
nor \U$11976 ( \20795 , \20754 , \20794 );
and \U$11977 ( \20796 , \20633 , \20714 , \20795 );
not \U$11978 ( \20797 , \9906 );
and \U$11979 ( \20798 , \20797 , \20452 );
and \U$11980 ( \20799 , \20456 , \9902 );
nor \U$11981 ( \20800 , \20798 , \20799 );
not \U$11982 ( \20801 , \9898 );
and \U$11983 ( \20802 , \20801 , \12575 );
and \U$11984 ( \20803 , \20458 , \9892 );
nor \U$11985 ( \20804 , \20802 , \20803 );
nand \U$11986 ( \20805 , \20800 , \20804 );
not \U$11987 ( \20806 , \20805 );
not \U$11988 ( \20807 , \9914 );
and \U$11989 ( \20808 , \20807 , \20449 );
and \U$11990 ( \20809 , \20483 , \9910 );
nor \U$11991 ( \20810 , \20808 , \20809 );
not \U$11992 ( \20811 , \9921 );
and \U$11993 ( \20812 , \20811 , \12552 );
and \U$11994 ( \20813 , \20481 , \9917 );
nor \U$11995 ( \20814 , \20812 , \20813 );
and \U$11996 ( \20815 , \20806 , \20810 , \20814 );
not \U$11997 ( \20816 , \9884 );
and \U$11998 ( \20817 , \20816 , \12531 );
and \U$11999 ( \20818 , \20477 , \9886 );
nor \U$12000 ( \20819 , \20817 , \20818 );
not \U$12001 ( \20820 , \9878 );
and \U$12002 ( \20821 , \20820 , \20470 );
and \U$12003 ( \20822 , \20443 , \9874 );
nor \U$12004 ( \20823 , \20821 , \20822 );
nand \U$12005 ( \20824 , \20819 , \20823 );
not \U$12006 ( \20825 , \20824 );
not \U$12007 ( \20826 , \9868 );
and \U$12008 ( \20827 , \20826 , \20463 );
and \U$12009 ( \20828 , \20465 , \9871 );
nor \U$12010 ( \20829 , \20827 , \20828 );
not \U$12011 ( \20830 , \9860 );
and \U$12012 ( \20831 , \20830 , \12512 );
and \U$12013 ( \20832 , \20438 , \9864 );
nor \U$12014 ( \20833 , \20831 , \20832 );
and \U$12015 ( \20834 , \20825 , \20829 , \20833 );
nand \U$12016 ( \20835 , \20815 , \20834 );
xnor \U$12017 ( \20836 , RIb7a0c48_261, \20835 );
not \U$12018 ( \20837 , \11693 );
and \U$12019 ( \20838 , \20837 , \20452 );
and \U$12020 ( \20839 , \20456 , \10027 );
nor \U$12021 ( \20840 , \20838 , \20839 );
not \U$12022 ( \20841 , \11698 );
and \U$12023 ( \20842 , \20841 , \12575 );
and \U$12024 ( \20843 , \20458 , \10035 );
nor \U$12025 ( \20844 , \20842 , \20843 );
nand \U$12026 ( \20845 , \20840 , \20844 );
not \U$12027 ( \20846 , \20845 );
not \U$12028 ( \20847 , \12222 );
and \U$12029 ( \20848 , \20847 , \20449 );
and \U$12030 ( \20849 , \20483 , \10043 );
nor \U$12031 ( \20850 , \20848 , \20849 );
not \U$12032 ( \20851 , \11674 );
and \U$12033 ( \20852 , \20851 , \12597 );
and \U$12034 ( \20853 , \20481 , \10047 );
nor \U$12035 ( \20854 , \20852 , \20853 );
and \U$12036 ( \20855 , \20846 , \20850 , \20854 );
not \U$12037 ( \20856 , \10018 );
and \U$12038 ( \20857 , \20856 , \12531 );
and \U$12039 ( \20858 , \20477 , \10020 );
nor \U$12040 ( \20859 , \20857 , \20858 );
not \U$12041 ( \20860 , \10013 );
and \U$12042 ( \20861 , \20860 , \20470 );
and \U$12043 ( \20862 , \20443 , \10009 );
nor \U$12044 ( \20863 , \20861 , \20862 );
nand \U$12045 ( \20864 , \20859 , \20863 );
not \U$12046 ( \20865 , \20864 );
not \U$12047 ( \20866 , \11666 );
and \U$12048 ( \20867 , \20866 , \20463 );
and \U$12049 ( \20868 , \20465 , \9996 );
nor \U$12050 ( \20869 , \20867 , \20868 );
not \U$12051 ( \20870 , \10002 );
and \U$12052 ( \20871 , \20870 , \12512 );
and \U$12053 ( \20872 , \20438 , \10004 );
nor \U$12054 ( \20873 , \20871 , \20872 );
and \U$12055 ( \20874 , \20865 , \20869 , \20873 );
nand \U$12056 ( \20875 , \20855 , \20874 );
xnor \U$12057 ( \20876 , RIb7af540_256, \20875 );
not \U$12058 ( \20877 , \9564 );
and \U$12059 ( \20878 , \20877 , \20452 );
and \U$12060 ( \20879 , \20456 , \9560 );
nor \U$12061 ( \20880 , \20878 , \20879 );
not \U$12062 ( \20881 , \9557 );
and \U$12063 ( \20882 , \20881 , \12575 );
and \U$12064 ( \20883 , \20458 , \9551 );
nor \U$12065 ( \20884 , \20882 , \20883 );
nand \U$12066 ( \20885 , \20880 , \20884 );
not \U$12067 ( \20886 , \20885 );
not \U$12068 ( \20887 , \9572 );
and \U$12069 ( \20888 , \20887 , \20449 );
and \U$12070 ( \20889 , \20483 , \9568 );
nor \U$12071 ( \20890 , \20888 , \20889 );
not \U$12072 ( \20891 , \9579 );
and \U$12073 ( \20892 , \20891 , \12597 );
and \U$12074 ( \20893 , \20481 , \9575 );
nor \U$12075 ( \20894 , \20892 , \20893 );
and \U$12076 ( \20895 , \20886 , \20890 , \20894 );
not \U$12077 ( \20896 , \9543 );
and \U$12078 ( \20897 , \20896 , \12531 );
and \U$12079 ( \20898 , \20477 , \9545 );
nor \U$12080 ( \20899 , \20897 , \20898 );
not \U$12081 ( \20900 , \9537 );
and \U$12082 ( \20901 , \20900 , \20470 );
and \U$12083 ( \20902 , \20443 , \9533 );
nor \U$12084 ( \20903 , \20901 , \20902 );
nand \U$12085 ( \20904 , \20899 , \20903 );
not \U$12086 ( \20905 , \20904 );
not \U$12087 ( \20906 , \9527 );
and \U$12088 ( \20907 , \20906 , \20463 );
and \U$12089 ( \20908 , \20465 , \9530 );
nor \U$12090 ( \20909 , \20907 , \20908 );
not \U$12091 ( \20910 , \9519 );
and \U$12092 ( \20911 , \20910 , \12512 );
and \U$12093 ( \20912 , \20438 , \9523 );
nor \U$12094 ( \20913 , \20911 , \20912 );
and \U$12095 ( \20914 , \20905 , \20909 , \20913 );
nand \U$12096 ( \20915 , \20895 , \20914 );
xnor \U$12097 ( \20916 , \20915 , \9585 );
not \U$12098 ( \20917 , \11623 );
and \U$12099 ( \20918 , \20917 , \20452 );
and \U$12100 ( \20919 , \20456 , \10709 );
nor \U$12101 ( \20920 , \20918 , \20919 );
not \U$12102 ( \20921 , \11620 );
and \U$12103 ( \20922 , \20921 , \12575 );
and \U$12104 ( \20923 , \20458 , \9968 );
nor \U$12105 ( \20924 , \20922 , \20923 );
nand \U$12106 ( \20925 , \20920 , \20924 );
not \U$12107 ( \20926 , \20925 );
not \U$12108 ( \20927 , \11629 );
and \U$12109 ( \20928 , \20927 , \20449 );
and \U$12110 ( \20929 , \20483 , \9977 );
nor \U$12111 ( \20930 , \20928 , \20929 );
not \U$12112 ( \20931 , \12282 );
and \U$12113 ( \20932 , \20931 , \12597 );
and \U$12114 ( \20933 , \20481 , \9982 );
nor \U$12115 ( \20934 , \20932 , \20933 );
and \U$12116 ( \20935 , \20926 , \20930 , \20934 );
not \U$12117 ( \20936 , \9937 );
and \U$12118 ( \20937 , \20936 , \12531 );
and \U$12119 ( \20938 , \20477 , \9939 );
nor \U$12120 ( \20939 , \20937 , \20938 );
not \U$12121 ( \20940 , \9933 );
and \U$12122 ( \20941 , \20940 , \20470 );
and \U$12123 ( \20942 , \20443 , \9929 );
nor \U$12124 ( \20943 , \20941 , \20942 );
nand \U$12125 ( \20944 , \20939 , \20943 );
not \U$12126 ( \20945 , \20944 );
not \U$12127 ( \20946 , \13143 );
and \U$12128 ( \20947 , \20946 , \20463 );
and \U$12129 ( \20948 , \20465 , \9947 );
nor \U$12130 ( \20949 , \20947 , \20948 );
not \U$12131 ( \20950 , \9952 );
and \U$12132 ( \20951 , \20950 , \12512 );
and \U$12133 ( \20952 , \20438 , \9954 );
nor \U$12134 ( \20953 , \20951 , \20952 );
and \U$12135 ( \20954 , \20945 , \20949 , \20953 );
nand \U$12136 ( \20955 , \20935 , \20954 );
xnor \U$12137 ( \20956 , \20955 , \9990 );
nor \U$12138 ( \20957 , \20916 , \20956 );
nand \U$12139 ( \20958 , \20836 , \20876 , \20957 );
not \U$12140 ( \20959 , \20958 );
not \U$12141 ( \20960 , \9834 );
and \U$12142 ( \20961 , \20960 , \20452 );
and \U$12143 ( \20962 , \20456 , \9830 );
nor \U$12144 ( \20963 , \20961 , \20962 );
not \U$12145 ( \20964 , \9827 );
and \U$12146 ( \20965 , \20964 , \12575 );
and \U$12147 ( \20966 , \20458 , \9822 );
nor \U$12148 ( \20967 , \20965 , \20966 );
nand \U$12149 ( \20968 , \20963 , \20967 );
not \U$12150 ( \20969 , \20968 );
not \U$12151 ( \20970 , \9843 );
and \U$12152 ( \20971 , \20970 , \20449 );
and \U$12153 ( \20972 , \20483 , \9839 );
nor \U$12154 ( \20973 , \20971 , \20972 );
not \U$12155 ( \20974 , \9851 );
and \U$12156 ( \20975 , \20974 , \12552 );
and \U$12157 ( \20976 , \20481 , \9847 );
nor \U$12158 ( \20977 , \20975 , \20976 );
and \U$12159 ( \20978 , \20969 , \20973 , \20977 );
not \U$12160 ( \20979 , \9814 );
and \U$12161 ( \20980 , \20979 , \12531 );
and \U$12162 ( \20981 , \20477 , \9816 );
nor \U$12163 ( \20982 , \20980 , \20981 );
not \U$12164 ( \20983 , \9809 );
and \U$12165 ( \20984 , \20983 , \20470 );
and \U$12166 ( \20985 , \20443 , \9805 );
nor \U$12167 ( \20986 , \20984 , \20985 );
nand \U$12168 ( \20987 , \20982 , \20986 );
not \U$12169 ( \20988 , \20987 );
not \U$12170 ( \20989 , \9798 );
and \U$12171 ( \20990 , \20989 , \20463 );
and \U$12172 ( \20991 , \20465 , \9801 );
nor \U$12173 ( \20992 , \20990 , \20991 );
not \U$12174 ( \20993 , \9791 );
and \U$12175 ( \20994 , \20993 , \12512 );
and \U$12176 ( \20995 , \20438 , \9794 );
nor \U$12177 ( \20996 , \20994 , \20995 );
and \U$12178 ( \20997 , \20988 , \20992 , \20996 );
nand \U$12179 ( \20998 , \20978 , \20997 );
xnor \U$12180 ( \20999 , \20998 , \9857 );
not \U$12181 ( \21000 , \11545 );
and \U$12182 ( \21001 , \21000 , \12575 );
and \U$12183 ( \21002 , \20458 , \8953 );
nor \U$12184 ( \21003 , \21001 , \21002 );
not \U$12185 ( \21004 , \11540 );
and \U$12186 ( \21005 , \21004 , \20452 );
and \U$12187 ( \21006 , \20456 , \8927 );
nor \U$12188 ( \21007 , \21005 , \21006 );
nand \U$12189 ( \21008 , \21003 , \21007 );
not \U$12190 ( \21009 , \21008 );
not \U$12191 ( \21010 , \11565 );
and \U$12192 ( \21011 , \21010 , \12552 );
and \U$12193 ( \21012 , \20481 , \8827 );
nor \U$12194 ( \21013 , \21011 , \21012 );
not \U$12195 ( \21014 , \8853 );
and \U$12196 ( \21015 , \21014 , \20483 );
and \U$12197 ( \21016 , \20449 , \8904 );
nor \U$12198 ( \21017 , \21015 , \21016 );
and \U$12199 ( \21018 , \21009 , \21013 , \21017 );
not \U$12200 ( \21019 , \8861 );
and \U$12201 ( \21020 , \21019 , \20443 );
and \U$12202 ( \21021 , \20470 , \8915 );
nor \U$12203 ( \21022 , \21020 , \21021 );
not \U$12204 ( \21023 , \10775 );
and \U$12205 ( \21024 , \21023 , \12531 );
and \U$12206 ( \21025 , \20477 , \8843 );
nor \U$12207 ( \21026 , \21024 , \21025 );
nand \U$12208 ( \21027 , \21022 , \21026 );
not \U$12209 ( \21028 , \21027 );
not \U$12210 ( \21029 , \12351 );
and \U$12211 ( \21030 , \21029 , \20463 );
and \U$12212 ( \21031 , \20465 , \8881 );
nor \U$12213 ( \21032 , \21030 , \21031 );
not \U$12214 ( \21033 , \8894 );
and \U$12215 ( \21034 , \21033 , \12512 );
and \U$12216 ( \21035 , \20438 , \8896 );
nor \U$12217 ( \21036 , \21034 , \21035 );
and \U$12218 ( \21037 , \21028 , \21032 , \21036 );
nand \U$12219 ( \21038 , \21018 , \21037 );
xnor \U$12220 ( \21039 , \21038 , \8964 );
nor \U$12221 ( \21040 , \20999 , \21039 );
not \U$12222 ( \21041 , \11473 );
and \U$12223 ( \21042 , \21041 , \12575 );
and \U$12224 ( \21043 , \20458 , \9112 );
nor \U$12225 ( \21044 , \21042 , \21043 );
not \U$12226 ( \21045 , \11468 );
and \U$12227 ( \21046 , \21045 , \20452 );
and \U$12228 ( \21047 , \20456 , \9093 );
nor \U$12229 ( \21048 , \21046 , \21047 );
nand \U$12230 ( \21049 , \21044 , \21048 );
not \U$12231 ( \21050 , \21049 );
not \U$12232 ( \21051 , \11452 );
and \U$12233 ( \21052 , \21051 , \12597 );
and \U$12234 ( \21053 , \20481 , \9046 );
nor \U$12235 ( \21054 , \21052 , \21053 );
not \U$12236 ( \21055 , \9055 );
and \U$12237 ( \21056 , \21055 , \20483 );
and \U$12238 ( \21057 , \20449 , \9081 );
nor \U$12239 ( \21058 , \21056 , \21057 );
and \U$12240 ( \21059 , \21050 , \21054 , \21058 );
not \U$12241 ( \21060 , \9058 );
and \U$12242 ( \21061 , \21060 , \20443 );
and \U$12243 ( \21062 , \20470 , \9085 );
nor \U$12244 ( \21063 , \21061 , \21062 );
not \U$12245 ( \21064 , \10859 );
and \U$12246 ( \21065 , \21064 , \12531 );
and \U$12247 ( \21066 , \20477 , \9049 );
nor \U$12248 ( \21067 , \21065 , \21066 );
nand \U$12249 ( \21068 , \21063 , \21067 );
not \U$12250 ( \21069 , \21068 );
not \U$12251 ( \21070 , \11458 );
and \U$12252 ( \21071 , \21070 , \20463 );
and \U$12253 ( \21072 , \20465 , \9067 );
nor \U$12254 ( \21073 , \21071 , \21072 );
not \U$12255 ( \21074 , \9073 );
and \U$12256 ( \21075 , \21074 , \12512 );
and \U$12257 ( \21076 , \20438 , \9075 );
nor \U$12258 ( \21077 , \21075 , \21076 );
and \U$12259 ( \21078 , \21069 , \21073 , \21077 );
nand \U$12260 ( \21079 , \21059 , \21078 );
xnor \U$12261 ( \21080 , \21079 , \9119 );
not \U$12262 ( \21081 , \11431 );
and \U$12263 ( \21082 , \21081 , \12575 );
and \U$12264 ( \21083 , \20458 , \9180 );
nor \U$12265 ( \21084 , \21082 , \21083 );
not \U$12266 ( \21085 , \11426 );
and \U$12267 ( \21086 , \21085 , \20452 );
and \U$12268 ( \21087 , \20456 , \9163 );
nor \U$12269 ( \21088 , \21086 , \21087 );
nand \U$12270 ( \21089 , \21084 , \21088 );
not \U$12271 ( \21090 , \21089 );
not \U$12272 ( \21091 , \11410 );
and \U$12273 ( \21092 , \21091 , \12552 );
and \U$12274 ( \21093 , \20481 , \9121 );
nor \U$12275 ( \21094 , \21092 , \21093 );
not \U$12276 ( \21095 , \9130 );
and \U$12277 ( \21096 , \21095 , \20483 );
and \U$12278 ( \21097 , \20449 , \9155 );
nor \U$12279 ( \21098 , \21096 , \21097 );
and \U$12280 ( \21099 , \21090 , \21094 , \21098 );
not \U$12281 ( \21100 , \9133 );
and \U$12282 ( \21101 , \21100 , \20443 );
and \U$12283 ( \21102 , \20470 , \9157 );
nor \U$12284 ( \21103 , \21101 , \21102 );
not \U$12285 ( \21104 , \10901 );
and \U$12286 ( \21105 , \21104 , \12531 );
and \U$12287 ( \21106 , \20477 , \9124 );
nor \U$12288 ( \21107 , \21105 , \21106 );
nand \U$12289 ( \21108 , \21103 , \21107 );
not \U$12290 ( \21109 , \21108 );
not \U$12291 ( \21110 , \11416 );
and \U$12292 ( \21111 , \21110 , \20463 );
and \U$12293 ( \21112 , \20465 , \9142 );
nor \U$12294 ( \21113 , \21111 , \21112 );
not \U$12295 ( \21114 , \9148 );
and \U$12296 ( \21115 , \21114 , \12512 );
and \U$12297 ( \21116 , \20438 , \9150 );
nor \U$12298 ( \21117 , \21115 , \21116 );
and \U$12299 ( \21118 , \21109 , \21113 , \21117 );
nand \U$12300 ( \21119 , \21099 , \21118 );
xnor \U$12301 ( \21120 , \21119 , \9188 );
nor \U$12302 ( \21121 , \21080 , \21120 );
and \U$12303 ( \21122 , \20959 , \21040 , \21121 );
nand \U$12304 ( \21123 , \20488 , \20796 , \21122 );
not \U$12305 ( \21124 , \21123 );
not \U$12306 ( \21125 , \21124 );
and \U$12307 ( \21126 , \20434 , \21125 );
buf \U$12308 ( \21127 , RIea91330_6888);
buf \U$12309 ( \21128 , \14685 );
buf \U$12310 ( \21129 , \12456 );
buf \U$12311 ( \21130 , \12458 );
buf \U$12312 ( \21131 , \8870 );
and \U$12313 ( \21132 , \21130 , \21131 );
and \U$12314 ( \21133 , \21129 , \21132 );
and \U$12315 ( \21134 , \21128 , \21133 );
and \U$12316 ( \21135 , \21127 , \21134 );
buf \U$12317 ( \21136 , \21135 );
not \U$12318 ( \21137 , \21136 );
not \U$12319 ( \21138 , \21131 );
buf \U$12320 ( \21139 , \21138 );
not \U$12321 ( \21140 , \21139 );
xor \U$12322 ( \21141 , \21130 , \21131 );
buf \U$12323 ( \21142 , \21141 );
not \U$12324 ( \21143 , \21142 );
nand \U$12325 ( \21144 , \21140 , \21143 );
xor \U$12326 ( \21145 , \21129 , \21132 );
buf \U$12327 ( \21146 , \21145 );
not \U$12328 ( \21147 , \21146 );
xor \U$12329 ( \21148 , \21128 , \21133 );
buf \U$12330 ( \21149 , \21148 );
not \U$12331 ( \21150 , \21149 );
nand \U$12332 ( \21151 , \21147 , \21150 );
or \U$12333 ( \21152 , \21144 , \21151 );
xor \U$12334 ( \21153 , \21127 , \21134 );
buf \U$12335 ( \21154 , \21153 );
nand \U$12336 ( \21155 , \21152 , \21154 );
nand \U$12337 ( \21156 , \21137 , \21155 );
not \U$12338 ( \21157 , \21124 );
or \U$12339 ( \21158 , \21156 , \21157 );
not \U$12340 ( \21159 , \21158 );
not \U$12341 ( \21160 , \21156 );
not \U$12342 ( \21161 , \21124 );
or \U$12343 ( \21162 , \21160 , \21161 );
not \U$12344 ( \21163 , \21162 );
or \U$12345 ( \21164 , \21159 , \21163 );
not \U$12346 ( \21165 , \21164 );
not \U$12347 ( \21166 , \21165 );
and \U$12348 ( \21167 , \21166 , \12494 );
nor \U$12349 ( \21168 , \21126 , \21167 );
or \U$12350 ( \21169 , \10061 , \21168 );
not \U$12351 ( \21170 , \10060 );
nand \U$12352 ( \21171 , \12454 , \21170 );
nand \U$12353 ( \21172 , \21169 , \21171 );
not \U$12354 ( \21173 , \21172 );
not \U$12355 ( \21174 , \21123 );
not \U$12356 ( \21175 , \13245 );
and \U$12357 ( \21176 , \21175 , \13920 , \14668 );
not \U$12358 ( \21177 , \11753 );
not \U$12359 ( \21178 , \15289 );
and \U$12360 ( \21179 , \21177 , \21178 );
not \U$12361 ( \21180 , \11754 );
not \U$12362 ( \21181 , \16004 );
and \U$12363 ( \21182 , \21180 , \21181 );
not \U$12364 ( \21183 , \10951 );
not \U$12365 ( \21184 , \16695 );
and \U$12366 ( \21185 , \21183 , \21184 );
not \U$12367 ( \21186 , \17471 );
or \U$12368 ( \21187 , \13992 , \21186 );
not \U$12369 ( \21188 , \21187 );
not \U$12370 ( \21189 , \18273 );
not \U$12371 ( \21190 , \21189 );
or \U$12372 ( \21191 , \17471 , \21190 );
not \U$12373 ( \21192 , \21191 );
and \U$12374 ( \21193 , \10928 , \21192 );
not \U$12375 ( \21194 , \18273 );
or \U$12376 ( \21195 , \17471 , \21194 );
not \U$12377 ( \21196 , \21195 );
and \U$12378 ( \21197 , \11753 , \21196 );
nor \U$12379 ( \21198 , \21188 , \21193 , \21197 );
not \U$12380 ( \21199 , \21198 );
and \U$12381 ( \21200 , \21199 , \16695 );
or \U$12382 ( \21201 , \21185 , \21200 );
not \U$12383 ( \21202 , \21201 );
and \U$12384 ( \21203 , \21202 , \16004 );
or \U$12385 ( \21204 , \21182 , \21203 );
not \U$12386 ( \21205 , \21204 );
and \U$12387 ( \21206 , \21205 , \15289 );
or \U$12388 ( \21207 , \21179 , \21206 );
and \U$12389 ( \21208 , \21176 , \21207 );
not \U$12390 ( \21209 , \13992 );
not \U$12391 ( \21210 , \13244 );
or \U$12392 ( \21211 , \13935 , \21210 );
not \U$12393 ( \21212 , \14676 );
or \U$12394 ( \21213 , \21209 , \21211 , \21212 );
not \U$12395 ( \21214 , \13941 );
or \U$12396 ( \21215 , \11754 , \21214 );
nand \U$12397 ( \21216 , \21213 , \21215 );
not \U$12398 ( \21217 , \13247 );
not \U$12399 ( \21218 , \13947 );
or \U$12400 ( \21219 , \21217 , \21218 );
not \U$12401 ( \21220 , \21219 );
not \U$12402 ( \21221 , \21220 );
not \U$12403 ( \21222 , \13935 );
and \U$12404 ( \21223 , \21222 , \10951 );
and \U$12405 ( \21224 , \21221 , \21223 );
nor \U$12406 ( \21225 , \21216 , \21224 );
not \U$12407 ( \21226 , \21225 );
nor \U$12408 ( \21227 , \21208 , \21226 );
not \U$12409 ( \21228 , \11750 );
and \U$12410 ( \21229 , \21228 , \18939 );
nand \U$12411 ( \21230 , \10914 , \19602 , \21229 );
or \U$12412 ( \21231 , \21227 , \21230 );
nor \U$12413 ( \21232 , \11752 , \10915 );
not \U$12414 ( \21233 , \11750 );
and \U$12415 ( \21234 , \21232 , \21233 );
not \U$12416 ( \21235 , \21234 );
or \U$12417 ( \21236 , \21235 , \19646 );
not \U$12418 ( \21237 , \19758 );
or \U$12419 ( \21238 , \10928 , \21237 );
not \U$12420 ( \21239 , \21238 );
not \U$12421 ( \21240 , \10915 );
not \U$12422 ( \21241 , \13992 );
and \U$12423 ( \21242 , \21240 , \21241 , \11749 );
not \U$12424 ( \21243 , \21242 );
not \U$12425 ( \21244 , \19680 );
nor \U$12426 ( \21245 , \21243 , \21244 );
not \U$12427 ( \21246 , \19723 );
not \U$12428 ( \21247 , \21246 );
not \U$12429 ( \21248 , \10915 );
and \U$12430 ( \21249 , \10918 , \21248 );
and \U$12431 ( \21250 , \21247 , \21249 );
nor \U$12432 ( \21251 , \21239 , \21245 , \21250 );
nand \U$12433 ( \21252 , \21236 , \21251 );
not \U$12434 ( \21253 , \21252 );
and \U$12435 ( \21254 , \21231 , \21253 );
nor \U$12436 ( \21255 , \21254 , \19728 );
not \U$12437 ( \21256 , \19798 );
and \U$12438 ( \21257 , \21256 , \11752 );
or \U$12439 ( \21258 , \21255 , \21257 );
not \U$12440 ( \21259 , \20397 );
and \U$12441 ( \21260 , \21258 , \21259 );
not \U$12442 ( \21261 , \20431 );
and \U$12443 ( \21262 , \21261 , \13992 );
nor \U$12444 ( \21263 , \21260 , \21262 );
or \U$12445 ( \21264 , \21174 , \21263 );
not \U$12446 ( \21265 , \21164 );
or \U$12447 ( \21266 , \10918 , \21265 );
nand \U$12448 ( \21267 , \21264 , \21266 );
not \U$12449 ( \21268 , \21267 );
not \U$12450 ( \21269 , \21170 );
and \U$12451 ( \21270 , \21268 , \21269 );
not \U$12452 ( \21271 , \8837 );
and \U$12453 ( \21272 , \21271 , \21170 );
or \U$12454 ( \21273 , \21270 , \21272 );
not \U$12455 ( \21274 , \21273 );
or \U$12456 ( \21275 , \21173 , \21274 );
not \U$12457 ( \21276 , \21123 );
not \U$12458 ( \21277 , \19798 );
and \U$12459 ( \21278 , \10920 , \21277 );
not \U$12460 ( \21279 , \13245 );
and \U$12461 ( \21280 , \21279 , \13920 , \14668 );
not \U$12462 ( \21281 , \10920 );
not \U$12463 ( \21282 , \15289 );
and \U$12464 ( \21283 , \21281 , \21282 );
not \U$12465 ( \21284 , \10920 );
not \U$12466 ( \21285 , \16004 );
and \U$12467 ( \21286 , \21284 , \21285 );
not \U$12468 ( \21287 , \10920 );
not \U$12469 ( \21288 , \16695 );
and \U$12470 ( \21289 , \21287 , \21288 );
not \U$12471 ( \21290 , \21195 );
not \U$12472 ( \21291 , \8870 );
and \U$12473 ( \21292 , \21290 , \21291 );
not \U$12474 ( \21293 , \21191 );
not \U$12475 ( \21294 , \21293 );
and \U$12476 ( \21295 , \17472 , \21294 );
not \U$12477 ( \21296 , \21295 );
and \U$12478 ( \21297 , \21296 , \8870 );
or \U$12479 ( \21298 , \21292 , \21297 );
not \U$12480 ( \21299 , \21298 );
and \U$12481 ( \21300 , \21299 , \16695 );
or \U$12482 ( \21301 , \21289 , \21300 );
not \U$12483 ( \21302 , \21301 );
and \U$12484 ( \21303 , \21302 , \16004 );
or \U$12485 ( \21304 , \21286 , \21303 );
not \U$12486 ( \21305 , \21304 );
and \U$12487 ( \21306 , \21305 , \15289 );
or \U$12488 ( \21307 , \21283 , \21306 );
not \U$12489 ( \21308 , \21307 );
and \U$12490 ( \21309 , \21280 , \21308 );
not \U$12491 ( \21310 , \13941 );
or \U$12492 ( \21311 , \10920 , \21310 );
not \U$12493 ( \21312 , \21220 );
and \U$12494 ( \21313 , \21312 , \13920 );
not \U$12495 ( \21314 , \21313 );
not \U$12496 ( \21315 , \10919 );
and \U$12497 ( \21316 , \21314 , \21315 );
not \U$12498 ( \21317 , \21212 );
and \U$12499 ( \21318 , \13244 , \21317 );
not \U$12500 ( \21319 , \21318 );
and \U$12501 ( \21320 , \21319 , \10919 );
or \U$12502 ( \21321 , \21316 , \21320 );
nand \U$12503 ( \21322 , \21311 , \21321 );
or \U$12504 ( \21323 , \21309 , \21322 );
nand \U$12505 ( \21324 , \18939 , \19602 );
not \U$12506 ( \21325 , \21324 );
and \U$12507 ( \21326 , \21323 , \21325 );
not \U$12508 ( \21327 , \19646 );
not \U$12509 ( \21328 , \10937 );
and \U$12510 ( \21329 , \21327 , \21328 );
not \U$12511 ( \21330 , \21244 );
and \U$12512 ( \21331 , \21330 , \10937 );
or \U$12513 ( \21332 , \21329 , \21331 );
nor \U$12514 ( \21333 , \21326 , \21332 );
nand \U$12515 ( \21334 , \10914 , \11749 );
or \U$12516 ( \21335 , \21333 , \21334 );
not \U$12517 ( \21336 , \19725 );
not \U$12518 ( \21337 , \10919 );
and \U$12519 ( \21338 , \21336 , \21337 );
not \U$12520 ( \21339 , \19758 );
not \U$12521 ( \21340 , \21339 );
and \U$12522 ( \21341 , \21340 , \10919 );
or \U$12523 ( \21342 , \21338 , \21341 );
not \U$12524 ( \21343 , \21342 );
and \U$12525 ( \21344 , \21335 , \21343 );
nor \U$12526 ( \21345 , \21344 , \19728 );
or \U$12527 ( \21346 , \21278 , \21345 );
and \U$12528 ( \21347 , \21346 , \20396 );
not \U$12529 ( \21348 , \20431 );
and \U$12530 ( \21349 , \21348 , \10937 );
nor \U$12531 ( \21350 , \21347 , \21349 );
or \U$12532 ( \21351 , \21276 , \21350 );
not \U$12533 ( \21352 , \21164 );
or \U$12534 ( \21353 , \8835 , \21352 );
nand \U$12535 ( \21354 , \21351 , \21353 );
not \U$12536 ( \21355 , \21354 );
not \U$12537 ( \21356 , \21170 );
and \U$12538 ( \21357 , \21355 , \21356 );
not \U$12539 ( \21358 , \8870 );
and \U$12540 ( \21359 , \21358 , \21170 );
or \U$12541 ( \21360 , \21357 , \21359 );
not \U$12542 ( \21361 , \21360 );
not \U$12543 ( \21362 , \21123 );
not \U$12544 ( \21363 , \19798 );
and \U$12545 ( \21364 , \21363 , \10923 );
nor \U$12546 ( \21365 , \13935 , \14669 );
nand \U$12547 ( \21366 , \21365 , \19602 );
not \U$12548 ( \21367 , \21366 );
and \U$12549 ( \21368 , \21367 , \13244 );
not \U$12550 ( \21369 , \16695 );
and \U$12551 ( \21370 , \10923 , \21369 );
not \U$12552 ( \21371 , \21195 );
and \U$12553 ( \21372 , \10923 , \21371 );
not \U$12554 ( \21373 , \17472 );
not \U$12555 ( \21374 , \8830 );
and \U$12556 ( \21375 , \21373 , \21374 );
not \U$12557 ( \21376 , \21191 );
and \U$12558 ( \21377 , \21376 , \8830 );
or \U$12559 ( \21378 , \21375 , \21377 );
nor \U$12560 ( \21379 , \21372 , \21378 );
and \U$12561 ( \21380 , \21379 , \16695 );
or \U$12562 ( \21381 , \21370 , \21380 );
not \U$12563 ( \21382 , \21381 );
nand \U$12564 ( \21383 , \15289 , \16004 );
not \U$12565 ( \21384 , \21383 );
and \U$12566 ( \21385 , \21382 , \21384 );
not \U$12567 ( \21386 , \10947 );
not \U$12568 ( \21387 , \21386 );
not \U$12569 ( \21388 , \15289 );
and \U$12570 ( \21389 , \21387 , \21388 );
not \U$12571 ( \21390 , \8830 );
and \U$12572 ( \21391 , \21390 , \15289 );
or \U$12573 ( \21392 , \21389 , \21391 );
not \U$12574 ( \21393 , \21392 );
and \U$12575 ( \21394 , \21393 , \21383 );
or \U$12576 ( \21395 , \21385 , \21394 );
and \U$12577 ( \21396 , \21368 , \21395 );
not \U$12578 ( \21397 , \19680 );
or \U$12579 ( \21398 , \8905 , \21397 );
not \U$12580 ( \21399 , \21398 );
not \U$12581 ( \21400 , \19644 );
not \U$12582 ( \21401 , \21400 );
not \U$12583 ( \21402 , \10947 );
and \U$12584 ( \21403 , \21401 , \21402 );
not \U$12585 ( \21404 , \13935 );
not \U$12586 ( \21405 , \19603 );
and \U$12587 ( \21406 , \21404 , \21405 , \21219 );
not \U$12588 ( \21407 , \21406 );
not \U$12589 ( \21408 , \21407 );
and \U$12590 ( \21409 , \21408 , \10947 );
or \U$12591 ( \21410 , \21403 , \21409 );
not \U$12592 ( \21411 , \19603 );
nor \U$12593 ( \21412 , \13935 , \13245 );
nand \U$12594 ( \21413 , \21411 , \14676 , \21412 );
not \U$12595 ( \21414 , \21413 );
not \U$12596 ( \21415 , \8905 );
and \U$12597 ( \21416 , \21414 , \21415 );
not \U$12598 ( \21417 , \19602 );
not \U$12599 ( \21418 , \13941 );
or \U$12600 ( \21419 , \21417 , \21418 );
not \U$12601 ( \21420 , \21419 );
and \U$12602 ( \21421 , \21420 , \8905 );
or \U$12603 ( \21422 , \21416 , \21421 );
nor \U$12604 ( \21423 , \21399 , \21410 , \21422 );
not \U$12605 ( \21424 , \21423 );
nor \U$12606 ( \21425 , \21396 , \21424 );
not \U$12607 ( \21426 , \18940 );
not \U$12608 ( \21427 , \21398 );
or \U$12609 ( \21428 , \21426 , \21427 );
not \U$12610 ( \21429 , \11750 );
and \U$12611 ( \21430 , \21429 , \10914 );
nand \U$12612 ( \21431 , \21428 , \21430 );
or \U$12613 ( \21432 , \21425 , \21431 );
not \U$12614 ( \21433 , \10947 );
or \U$12615 ( \21434 , \21433 , \19725 );
not \U$12616 ( \21435 , \19758 );
or \U$12617 ( \21436 , \10067 , \21435 );
nand \U$12618 ( \21437 , \21434 , \21436 );
not \U$12619 ( \21438 , \21437 );
and \U$12620 ( \21439 , \21432 , \21438 );
nor \U$12621 ( \21440 , \21439 , \19728 );
or \U$12622 ( \21441 , \21364 , \21440 );
and \U$12623 ( \21442 , \21441 , \20396 );
not \U$12624 ( \21443 , \20431 );
and \U$12625 ( \21444 , \10067 , \21443 );
nor \U$12626 ( \21445 , \21442 , \21444 );
or \U$12627 ( \21446 , \21362 , \21445 );
not \U$12628 ( \21447 , \21164 );
or \U$12629 ( \21448 , \10923 , \21447 );
nand \U$12630 ( \21449 , \21446 , \21448 );
not \U$12631 ( \21450 , \21449 );
not \U$12632 ( \21451 , \21170 );
and \U$12633 ( \21452 , \21450 , \21451 );
not \U$12634 ( \21453 , \8905 );
and \U$12635 ( \21454 , \21453 , \21170 );
or \U$12636 ( \21455 , \21452 , \21454 );
and \U$12637 ( \21456 , \21361 , \21455 );
not \U$12638 ( \21457 , \21456 );
or \U$12639 ( \21458 , \21275 , \21457 );
not \U$12640 ( \21459 , \21458 );
not \U$12641 ( \21460 , \16694 );
and \U$12642 ( \21461 , \21460 , \17472 , \16004 );
not \U$12643 ( \21462 , \18269 );
not \U$12644 ( \21463 , \13269 );
and \U$12645 ( \21464 , \21462 , \21463 );
not \U$12646 ( \21465 , \18280 );
and \U$12647 ( \21466 , \21465 , \13269 );
or \U$12648 ( \21467 , \21464 , \21466 );
nand \U$12649 ( \21468 , \21467 , \18273 );
not \U$12650 ( \21469 , \21468 );
not \U$12651 ( \21470 , \13923 );
not \U$12652 ( \21471 , \21470 );
not \U$12653 ( \21472 , \21471 );
and \U$12654 ( \21473 , \21469 , \21472 );
not \U$12655 ( \21474 , \13269 );
and \U$12656 ( \21475 , \18280 , \21474 );
and \U$12657 ( \21476 , \18269 , \13269 );
or \U$12658 ( \21477 , \21475 , \21476 );
not \U$12659 ( \21478 , \21477 );
and \U$12660 ( \21479 , \21478 , \21471 );
or \U$12661 ( \21480 , \21473 , \21479 );
not \U$12662 ( \21481 , \21480 );
and \U$12663 ( \21482 , \21461 , \21481 );
not \U$12664 ( \21483 , \21482 );
not \U$12665 ( \21484 , \11756 );
or \U$12666 ( \21485 , \10065 , \21484 );
xnor \U$12667 ( \21486 , \21471 , \21485 );
not \U$12668 ( \21487 , \21486 );
and \U$12669 ( \21488 , \15285 , \21487 );
not \U$12670 ( \21489 , \15286 );
and \U$12671 ( \21490 , \21489 , \21486 );
or \U$12672 ( \21491 , \21488 , \21490 );
not \U$12673 ( \21492 , \21491 );
not \U$12674 ( \21493 , \21470 );
not \U$12675 ( \21494 , \8909 );
or \U$12676 ( \21495 , \8837 , \21494 );
xnor \U$12677 ( \21496 , \21493 , \21495 );
not \U$12678 ( \21497 , \21496 );
and \U$12679 ( \21498 , \17468 , \21497 );
not \U$12680 ( \21499 , \17469 );
and \U$12681 ( \21500 , \21499 , \21496 );
or \U$12682 ( \21501 , \21498 , \21500 );
nand \U$12683 ( \21502 , \16004 , \21501 , \16695 );
not \U$12684 ( \21503 , \16000 );
xnor \U$12685 ( \21504 , \21493 , \13249 );
not \U$12686 ( \21505 , \21504 );
and \U$12687 ( \21506 , \21503 , \21505 );
not \U$12688 ( \21507 , \16001 );
not \U$12689 ( \21508 , \21507 );
and \U$12690 ( \21509 , \21508 , \21504 );
or \U$12691 ( \21510 , \21506 , \21509 );
and \U$12692 ( \21511 , \21492 , \21502 , \21510 );
not \U$12693 ( \21512 , \13256 );
nand \U$12694 ( \21513 , \16683 , \21512 );
xnor \U$12695 ( \21514 , \21513 , \21470 );
not \U$12696 ( \21515 , \16003 );
and \U$12697 ( \21516 , \21514 , \21515 );
and \U$12698 ( \21517 , \21516 , \16682 );
nand \U$12699 ( \21518 , \21471 , \10065 );
not \U$12700 ( \21519 , \21518 );
not \U$12701 ( \21520 , \21493 );
not \U$12702 ( \21521 , \10930 );
not \U$12703 ( \21522 , \21521 );
and \U$12704 ( \21523 , \21520 , \21522 );
not \U$12705 ( \21524 , \21470 );
or \U$12706 ( \21525 , \12454 , \21524 );
not \U$12707 ( \21526 , \21525 );
not \U$12708 ( \21527 , \21526 );
and \U$12709 ( \21528 , \21527 , \21521 );
or \U$12710 ( \21529 , \21523 , \21528 );
not \U$12711 ( \21530 , \21529 );
or \U$12712 ( \21531 , \21519 , \21530 );
not \U$12713 ( \21532 , \16003 );
and \U$12714 ( \21533 , \21531 , \21532 );
and \U$12715 ( \21534 , \21533 , \16677 );
nor \U$12716 ( \21535 , \21517 , \21534 );
and \U$12717 ( \21536 , \21483 , \21511 , \21535 );
or \U$12718 ( \21537 , \15289 , \21491 );
nand \U$12719 ( \21538 , \13244 , \14668 );
not \U$12720 ( \21539 , \21538 );
nand \U$12721 ( \21540 , \21537 , \21539 );
or \U$12722 ( \21541 , \21536 , \21540 );
and \U$12723 ( \21542 , \8908 , \13249 );
not \U$12725 ( \21543 , \14671 );
not \U$12726 ( \21544 , \21493 );
or \U$12727 ( \21545 , \21544 , \21542 );
nand \U$12728 ( \21546 , \21545 , \13932 );
and \U$12729 ( \21547 , \21543 , \13244 , \21546 );
nor \U$12730 ( \21548 , 1'b0 , \21547 );
not \U$12731 ( \21549 , \10067 );
nand \U$12732 ( \21550 , \10928 , \13244 );
not \U$12733 ( \21551 , \21550 );
not \U$12734 ( \21552 , \21493 );
and \U$12735 ( \21553 , \14672 , \21552 );
not \U$12736 ( \21554 , \14674 );
and \U$12737 ( \21555 , \21554 , \21493 );
or \U$12738 ( \21556 , \21553 , \21555 );
and \U$12739 ( \21557 , \21549 , \21551 , \21556 );
not \U$12740 ( \21558 , \21557 );
not \U$12741 ( \21559 , \13932 );
not \U$12742 ( \21560 , \21512 );
and \U$12743 ( \21561 , \8837 , \21560 );
not \U$12744 ( \21562 , \21561 );
not \U$12745 ( \21563 , \21471 );
and \U$12746 ( \21564 , \21562 , \21563 );
not \U$12747 ( \21565 , \13251 );
and \U$12748 ( \21566 , \21565 , \21471 );
or \U$12749 ( \21567 , \21564 , \21566 );
not \U$12750 ( \21568 , \21567 );
or \U$12751 ( \21569 , \21559 , \21568 );
not \U$12752 ( \21570 , \21569 );
not \U$12753 ( \21571 , \21570 );
and \U$12754 ( \21572 , \21571 , \21217 );
not \U$12755 ( \21573 , \21526 );
not \U$12756 ( \21574 , \10097 );
and \U$12757 ( \21575 , \21573 , \21574 );
not \U$12758 ( \21576 , \21493 );
and \U$12759 ( \21577 , \21576 , \10097 );
or \U$12760 ( \21578 , \21575 , \21577 );
not \U$12761 ( \21579 , \21578 );
or \U$12762 ( \21580 , \21519 , \21579 );
and \U$12763 ( \21581 , \13948 , \21580 );
nor \U$12764 ( \21582 , \21572 , \21581 );
nand \U$12765 ( \21583 , \21548 , \21558 , \21582 );
not \U$12766 ( \21584 , \21583 );
and \U$12767 ( \21585 , \21541 , \21584 );
not \U$12768 ( \21586 , \19602 );
or \U$12769 ( \21587 , \13935 , \21586 );
nor \U$12770 ( \21588 , \21585 , \21587 );
not \U$12771 ( \21589 , \19603 );
nand \U$12772 ( \21590 , \21493 , \8906 );
nand \U$12773 ( \21591 , \21590 , \13932 );
not \U$12774 ( \21592 , \13939 );
and \U$12775 ( \21593 , \21591 , \21592 );
and \U$12776 ( \21594 , \21589 , \21593 );
not \U$12777 ( \21595 , \21594 );
not \U$12778 ( \21596 , \19603 );
nand \U$12779 ( \21597 , \21518 , \21525 );
not \U$12780 ( \21598 , \13936 );
and \U$12781 ( \21599 , \21597 , \21598 );
and \U$12782 ( \21600 , \21596 , \21599 );
not \U$12783 ( \21601 , \21600 );
not \U$12784 ( \21602 , \19642 );
not \U$12785 ( \21603 , \21471 );
and \U$12787 ( \21604 , \19640 , \18277 , \21603 );
and \U$12789 ( \21605 , \21602 , \18277 , \21471 );
or \U$12790 ( \21606 , 1'b0 , \21604 , 1'b0 , \21605 );
not \U$12791 ( \21607 , \21606 );
and \U$12792 ( \21608 , \21595 , \21601 , \21607 );
not \U$12793 ( \21609 , \21608 );
or \U$12794 ( \21610 , \21588 , \21609 );
nand \U$12795 ( \21611 , \11749 , \18939 );
not \U$12796 ( \21612 , \21611 );
and \U$12797 ( \21613 , \21610 , \21612 );
not \U$12798 ( \21614 , \19721 );
or \U$12800 ( \21615 , \10928 , \8830 );
and \U$12801 ( \21616 , \21615 , \12454 );
not \U$12802 ( \21617 , \21616 );
not \U$12803 ( \21618 , \21471 );
and \U$12804 ( \21619 , \21617 , \21618 );
and \U$12805 ( \21620 , \8845 , \13254 );
not \U$12806 ( \21621 , \21620 );
and \U$12807 ( \21622 , \21621 , \21471 );
or \U$12808 ( \21623 , \21619 , \21622 );
not \U$12809 ( \21624 , \19678 );
nand \U$12810 ( \21625 , \21623 , \11749 , \21624 );
not \U$12811 ( \21626 , \21620 );
not \U$12812 ( \21627 , \21493 );
and \U$12813 ( \21628 , \21626 , \21627 );
not \U$12814 ( \21629 , \21616 );
and \U$12815 ( \21630 , \21629 , \21493 );
or \U$12816 ( \21631 , \21628 , \21630 );
nand \U$12817 ( \21632 , \21631 , \11749 , \19677 );
and \U$12818 ( \21633 , \21519 , \19718 );
and \U$12819 ( \21634 , \21559 , \21614 );
or \U$12820 ( \21635 , \21633 , \21634 );
nand \U$12821 ( \21636 , \21635 , \10930 );
and \U$12822 ( \21637 , 1'b1 , \21625 , \21632 , \21636 );
not \U$12823 ( \21638 , \21637 );
nor \U$12824 ( \21639 , \21613 , \21638 );
or \U$12825 ( \21640 , \10915 , \21639 );
not \U$12826 ( \21641 , \19753 );
xnor \U$12827 ( \21642 , \13255 , \21470 );
not \U$12828 ( \21643 , \21642 );
and \U$12829 ( \21644 , \21641 , \21643 );
not \U$12830 ( \21645 , \19756 );
not \U$12831 ( \21646 , \21645 );
and \U$12832 ( \21647 , \21646 , \21642 );
or \U$12833 ( \21648 , \21644 , \21647 );
and \U$12834 ( \21649 , \21640 , \21648 );
nor \U$12835 ( \21650 , \21649 , \19728 );
not \U$12836 ( \21651 , \19795 );
not \U$12837 ( \21652 , \11756 );
and \U$12838 ( \21653 , \12454 , \21652 );
not \U$12840 ( \21654 , \21651 );
not \U$12841 ( \21655 , \21493 );
and \U$12842 ( \21656 , \21654 , \21655 );
not \U$12843 ( \21657 , \19792 );
and \U$12844 ( \21658 , \21657 , \21493 );
or \U$12845 ( \21659 , \21656 , \21658 );
not \U$12846 ( \21660 , \21659 );
and \U$12847 ( \21661 , \21660 , \21653 );
or \U$12848 ( \21662 , 1'b0 , \21661 );
or \U$12849 ( \21663 , \21650 , \21662 );
not \U$12850 ( \21664 , \20397 );
and \U$12851 ( \21665 , \21663 , \21664 );
not \U$12852 ( \21666 , \8845 );
and \U$12853 ( \21667 , \8837 , \21666 );
xnor \U$12854 ( \21668 , \21667 , \21470 );
not \U$12855 ( \21669 , \21668 );
and \U$12856 ( \21670 , \20425 , \21669 );
not \U$12857 ( \21671 , \20428 );
and \U$12858 ( \21672 , \21671 , \21668 );
or \U$12859 ( \21673 , \21670 , \21672 );
nor \U$12860 ( \21674 , \21665 , \21673 );
or \U$12861 ( \21675 , \21124 , \21674 );
not \U$12862 ( \21676 , \21162 );
not \U$12864 ( \21677 , \21676 );
not \U$12865 ( \21678 , \21471 );
and \U$12866 ( \21679 , \21677 , \21678 );
not \U$12867 ( \21680 , \21159 );
and \U$12868 ( \21681 , \21680 , \21471 );
or \U$12869 ( \21682 , \21679 , \21681 );
not \U$12870 ( \21683 , \21682 );
and \U$12871 ( \21684 , \21683 , \13296 );
or \U$12872 ( \21685 , 1'b0 , \21684 );
not \U$12873 ( \21686 , \21685 );
nand \U$12874 ( \21687 , \21675 , \21686 );
not \U$12875 ( \21688 , \21170 );
and \U$12876 ( \21689 , \21687 , \21688 );
or \U$12877 ( \21690 , \10922 , \13249 );
nor \U$12878 ( \21691 , \21471 , \21690 );
and \U$12879 ( \21692 , \21691 , \21170 );
or \U$12880 ( \21693 , \21689 , \21692 );
not \U$12881 ( \21694 , \21693 );
and \U$12882 ( \21695 , \21459 , \21694 );
buf \U$12883 ( \21696 , \21695 );
nand \U$12884 ( \21697 , \8826 , \21696 );
not \U$12885 ( \21698 , \21697 );
buf \U$12886 ( \21699 , RIb7b9680_245);
buf \U$12887 ( \21700 , \21699 );
not \U$12888 ( \21701 , RIde4ec88_4006);
or \U$12889 ( \21702 , \21700 , \21701 );
nand \U$12890 ( \21703 , \21702 , \8826 , \21696 );
buf \U$12891 ( \21704 , RIb79b4a0_271);
and \U$12892 ( \21705 , \13923 , \8878 );
buf \U$12893 ( \21706 , \21705 );
nand \U$12894 ( \21707 , \21704 , \21706 );
not \U$12895 ( \21708 , \21707 );
buf \U$12896 ( \21709 , RIb79b338_274);
buf \U$12897 ( \21710 , \21709 );
nand \U$12898 ( \21711 , \21706 , \21710 );
not \U$12899 ( \21712 , \21711 );
nor \U$12900 ( \21713 , \21708 , \21712 );
nand \U$12901 ( \21714 , \21698 , \21703 , \21713 );
or \U$12902 ( \21715 , \8824 , \21714 );
nand \U$12903 ( \21716 , \8826 , \21696 );
not \U$12904 ( \21717 , \21716 );
not \U$12905 ( \21718 , \21717 );
and \U$12906 ( \21719 , \21711 , \21708 );
not \U$12907 ( \21720 , \8822 );
not \U$12908 ( \21721 , \21720 );
or \U$12909 ( \21722 , RIde68f20_3980, \21721 );
nand \U$12910 ( \21723 , \21718 , \21719 , \21722 );
nand \U$12911 ( \21724 , \21715 , \21723 );
not \U$12912 ( \21725 , \21724 );
or \U$12913 ( \21726 , \21717 , \21720 );
not \U$12914 ( \21727 , \8820 );
nand \U$12915 ( \21728 , RIde68638_3981, \21727 );
nand \U$12916 ( \21729 , \21726 , \21728 );
xnor \U$12917 ( \21730 , \21729 , \21716 );
nor \U$12918 ( \21731 , \21725 , \21730 );
not \U$12919 ( \21732 , \21731 );
not \U$12920 ( \21733 , RIde68f20_3980);
and \U$12921 ( \21734 , \21732 , \21733 );
not \U$12922 ( \21735 , \21712 );
not \U$12923 ( \21736 , \21703 );
not \U$12924 ( \21737 , \21736 );
xnor \U$12925 ( \21738 , \21708 , \21717 );
and \U$12926 ( \21739 , \21735 , \21737 , \21738 );
not \U$12927 ( \21740 , \21739 );
not \U$12928 ( \21741 , \21740 );
not \U$12929 ( \21742 , \21741 );
not \U$12930 ( \21743 , \21730 );
and \U$12931 ( \21744 , \21742 , \21743 );
nand \U$12932 ( \21745 , \21714 , \21723 );
nor \U$12933 ( \21746 , \21741 , \21745 );
nor \U$12934 ( \21747 , \21744 , \21746 );
not \U$12935 ( \21748 , \21747 );
and \U$12936 ( \21749 , \21748 , RIde68f20_3980);
or \U$12937 ( \21750 , \21734 , \21749 );
not \U$12938 ( \21751 , RIde612e8_3992);
nand \U$12939 ( \21752 , \21736 , \21711 );
not \U$12940 ( \21753 , \21752 );
not \U$12941 ( \21754 , \21753 );
or \U$12942 ( \21755 , \21751 , \21754 );
not \U$12943 ( \21756 , \21752 );
and \U$12944 ( \21757 , RIde5fec0_3994, \21756 );
not \U$12945 ( \21758 , \21741 );
not \U$12946 ( \21759 , \8820 );
and \U$12947 ( \21760 , \21758 , \21759 );
not \U$12948 ( \21761 , \21724 );
and \U$12949 ( \21762 , \21761 , \8820 );
or \U$12950 ( \21763 , \21760 , \21762 );
not \U$12951 ( \21764 , \21763 );
or \U$12952 ( \21765 , \21757 , \21764 );
nand \U$12953 ( \21766 , \21720 , \21716 );
not \U$12954 ( \21767 , \21717 );
or \U$12955 ( \21768 , \8820 , \21767 );
not \U$12956 ( \21769 , \21768 );
not \U$12957 ( \21770 , RIde68638_3981);
and \U$12958 ( \21771 , \21769 , \21770 );
xnor \U$12959 ( \21772 , \21717 , \21727 );
not \U$12960 ( \21773 , \21772 );
and \U$12961 ( \21774 , \21773 , RIde68638_3981);
or \U$12962 ( \21775 , \21771 , \21774 );
not \U$12963 ( \21776 , \21775 );
and \U$12964 ( \21777 , \21766 , \21776 );
or \U$12965 ( \21778 , \21725 , \21777 );
and \U$12966 ( \21779 , \21741 , RIde68638_3981);
not \U$12967 ( \21780 , \21752 );
and \U$12968 ( \21781 , RIde60988_3993, \21780 );
nor \U$12969 ( \21782 , \21779 , \21781 );
nand \U$12970 ( \21783 , \21778 , \21782 );
nor \U$12971 ( \21784 , \21765 , \21783 );
and \U$12972 ( \21785 , \21750 , \21755 , \21784 );
not \U$12973 ( \21786 , RIde69970_3979);
not \U$12974 ( \21787 , RIde6a2d0_3978);
not \U$12975 ( \21788 , RIde6ad98_3977);
not \U$12976 ( \21789 , \21788 );
nand \U$12977 ( \21790 , \21786 , \21787 , \21789 );
not \U$12978 ( \21791 , \21790 );
not \U$12979 ( \21792 , \21791 );
nor \U$12980 ( \21793 , \21787 , \21786 );
xnor \U$12981 ( \21794 , \21788 , \21793 );
not \U$12982 ( \21795 , \21707 );
and \U$12983 ( \21796 , \21794 , \21795 );
and \U$12984 ( \21797 , \21789 , \21707 );
or \U$12985 ( \21798 , \21796 , \21797 );
not \U$12986 ( \21799 , \21798 );
and \U$12987 ( \21800 , \21792 , \21799 );
nor \U$12988 ( \21801 , \21800 , \21712 );
not \U$12989 ( \21802 , RIde63250_3989);
not \U$12990 ( \21803 , RIde62878_3990);
not \U$12991 ( \21804 , RIde61e28_3991);
nor \U$12992 ( \21805 , \21803 , \21804 );
xnor \U$12993 ( \21806 , \21802 , \21805 );
buf \U$12994 ( \21807 , RIb839848_152);
not \U$12995 ( \21808 , RIe545648_6852);
nand \U$12996 ( \21809 , RIe545dc8_6851, \21808 );
not \U$12997 ( \21810 , RIea90778_6887);
not \U$12998 ( \21811 , \21810 );
not \U$12999 ( \21812 , RIe546890_6849);
not \U$13000 ( \21813 , RIe546098_6850);
nand \U$13001 ( \21814 , \21811 , \21812 , \21813 );
nor \U$13002 ( \21815 , \21809 , \21814 );
buf \U$13003 ( \21816 , \21815 );
and \U$13004 ( \21817 , \21807 , \21816 );
buf \U$13005 ( \21818 , RIb8396e0_155);
nand \U$13006 ( \21819 , \21818 , \21816 );
buf \U$13007 ( \21820 , RIb839668_156);
buf \U$13008 ( \21821 , \21820 );
not \U$13009 ( \21822 , \21821 );
nand \U$13010 ( \21823 , \21819 , \21822 );
not \U$13011 ( \21824 , \21823 );
nand \U$13012 ( \21825 , \21817 , \21824 );
not \U$13013 ( \21826 , \21825 );
not \U$13014 ( \21827 , \21803 );
or \U$13015 ( \21828 , \21802 , \21827 );
not \U$13016 ( \21829 , \21828 );
nand \U$13017 ( \21830 , RIde61e28_3991, \21829 );
nand \U$13018 ( \21831 , \21826 , \21830 );
not \U$13019 ( \21832 , \21831 );
and \U$13020 ( \21833 , \21806 , \21832 );
not \U$13021 ( \21834 , \21830 );
and \U$13022 ( \21835 , \21834 , \21826 );
xnor \U$13023 ( \21836 , \21802 , \21803 );
and \U$13024 ( \21837 , \21828 , \21836 );
nand \U$13025 ( \21838 , \21816 , \21819 , \21821 );
or \U$13026 ( \21839 , \21837 , \21838 );
not \U$13027 ( \21840 , \21822 );
not \U$13028 ( \21841 , \21819 );
or \U$13029 ( \21842 , \21840 , \21817 , \21841 );
nand \U$13030 ( \21843 , \21842 , \21816 );
not \U$13031 ( \21844 , \21843 );
or \U$13032 ( \21845 , \21844 , \21802 );
nand \U$13033 ( \21846 , \21839 , \21845 );
or \U$13034 ( \21847 , \21835 , \21846 );
or \U$13035 ( \21848 , \21833 , \21847 );
not \U$13036 ( \21849 , \21848 );
nor \U$13037 ( \21850 , \21801 , \21849 );
not \U$13038 ( \21851 , \21700 );
buf \U$13039 ( \21852 , RIb79b3b0_273);
nand \U$13040 ( \21853 , \21852 , \21696 );
not \U$13041 ( \21854 , \21853 );
and \U$13042 ( \21855 , \21851 , \21854 );
not \U$13043 ( \21856 , RIde5f3f8_3995);
and \U$13044 ( \21857 , \21856 , \21853 );
or \U$13045 ( \21858 , \21855 , \21857 );
nor \U$13046 ( \21859 , \21850 , \21858 );
or \U$13047 ( \21860 , \21844 , \21804 );
or \U$13048 ( \21861 , \21825 , \21830 );
nand \U$13049 ( \21862 , \21821 , \21816 );
not \U$13050 ( \21863 , \21862 );
nand \U$13051 ( \21864 , \21863 , \21818 );
not \U$13052 ( \21865 , \21864 );
nand \U$13053 ( \21866 , RIde61e28_3991, \21828 );
and \U$13054 ( \21867 , \21830 , \21866 );
or \U$13055 ( \21868 , \21867 , \21862 );
and \U$13056 ( \21869 , \21868 , \21819 );
or \U$13057 ( \21870 , \21865 , \21869 );
or \U$13058 ( \21871 , \21831 , RIde61e28_3991);
nand \U$13059 ( \21872 , \21860 , \21861 , \21870 , \21871 );
not \U$13060 ( \21873 , \21872 );
xor \U$13061 ( \21874 , \21803 , \21804 );
and \U$13062 ( \21875 , \21874 , \21832 );
not \U$13063 ( \21876 , \21803 );
not \U$13064 ( \21877 , \21876 );
not \U$13065 ( \21878 , \21843 );
or \U$13066 ( \21879 , \21877 , \21878 );
not \U$13067 ( \21880 , \21838 );
nand \U$13068 ( \21881 , \21803 , \21828 , \21880 );
nand \U$13069 ( \21882 , \21879 , \21881 , \21864 );
or \U$13070 ( \21883 , \21875 , \21882 );
xor \U$13071 ( \21884 , \21787 , \21786 );
and \U$13072 ( \21885 , \21884 , \21790 , \21719 );
not \U$13073 ( \21886 , \21787 );
and \U$13074 ( \21887 , \21707 , \21886 , \21711 );
or \U$13075 ( \21888 , \21885 , \21887 );
not \U$13076 ( \21889 , \21888 );
or \U$13077 ( \21890 , \21883 , \21889 );
and \U$13078 ( \21891 , \21786 , \21790 , \21719 );
not \U$13079 ( \21892 , \21786 );
and \U$13080 ( \21893 , \21707 , \21892 , \21711 );
nor \U$13081 ( \21894 , \21891 , \21893 );
nand \U$13082 ( \21895 , \21890 , \21894 );
or \U$13083 ( \21896 , \21873 , \21895 );
nand \U$13084 ( \21897 , \21883 , \21889 );
nand \U$13085 ( \21898 , \21896 , \21897 );
nand \U$13086 ( \21899 , \21801 , \21849 );
and \U$13087 ( \21900 , \21898 , \21899 );
nor \U$13088 ( \21901 , \21900 , \21701 );
and \U$13089 ( \21902 , \21859 , \21901 );
nor \U$13090 ( \21903 , \21785 , \21902 );
and \U$13092 ( \21904 , \21903 , 1'b1 );
or \U$13094 ( \21905 , \21904 , 1'b0 );
buf \U$13095 ( \21906 , \21905 );
not \U$13096 ( \21907 , RIe5319e0_6884);
nor \U$13097 ( \21908 , \21907 , RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
not \U$13098 ( \21909 , RIe549ef0_6842);
nor \U$13099 ( \21910 , RIe5319e0_6884, \21909 , RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
or \U$13100 ( \21911 , \21908 , \21910 );
nor \U$13101 ( \21912 , \21907 , \21909 , RIe549770_6843, RIe548ff0_6844, RIea91330_6888);
or \U$13102 ( \21913 , \21911 , \21912 );
not \U$13103 ( \21914 , RIe549770_6843);
nor \U$13104 ( \21915 , RIe5319e0_6884, RIe549ef0_6842, \21914 , RIe548ff0_6844, RIea91330_6888);
or \U$13105 ( \21916 , \21913 , \21915 );
nor \U$13106 ( \21917 , \21907 , RIe549ef0_6842, \21914 , RIe548ff0_6844, RIea91330_6888);
or \U$13107 ( \21918 , \21916 , \21917 );
nor \U$13108 ( \21919 , RIe5319e0_6884, \21909 , \21914 , RIe548ff0_6844, RIea91330_6888);
or \U$13109 ( \21920 , \21918 , \21919 );
nor \U$13110 ( \21921 , \21907 , \21909 , \21914 , RIe548ff0_6844, RIea91330_6888);
or \U$13111 ( \21922 , \21920 , \21921 );
not \U$13112 ( \21923 , RIea91330_6888);
and \U$13113 ( \21924 , \21907 , \21909 , \21914 , RIe548ff0_6844, \21923 );
or \U$13114 ( \21925 , \21922 , \21924 );
and \U$13115 ( \21926 , RIe5319e0_6884, \21909 , \21914 , RIe548ff0_6844, \21923 );
or \U$13116 ( \21927 , \21925 , \21926 );
and \U$13117 ( \21928 , \21907 , RIe549ef0_6842, \21914 , RIe548ff0_6844, \21923 );
or \U$13118 ( \21929 , \21927 , \21928 );
and \U$13119 ( \21930 , RIe5319e0_6884, RIe549ef0_6842, \21914 , RIe548ff0_6844, \21923 );
or \U$13120 ( \21931 , \21929 , \21930 );
and \U$13121 ( \21932 , \21907 , \21909 , RIe549770_6843, RIe548ff0_6844, \21923 );
or \U$13122 ( \21933 , \21931 , \21932 );
and \U$13123 ( \21934 , RIe5319e0_6884, \21909 , RIe549770_6843, RIe548ff0_6844, \21923 );
or \U$13124 ( \21935 , \21933 , \21934 );
and \U$13125 ( \21936 , \21907 , RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \21923 );
or \U$13126 ( \21937 , \21935 , \21936 );
and \U$13127 ( \21938 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \21923 );
or \U$13128 ( \21939 , \21937 , \21938 );
nor \U$13129 ( \21940 , RIe5319e0_6884, RIe549ef0_6842, RIe549770_6843, RIe548ff0_6844, \21923 );
or \U$13130 ( \21941 , \21939 , \21940 );
buf \U$13131 ( \21942 , \21941 );
not \U$13132 ( \21943 , \21942 );
buf \U$13133 ( \21944 , \21943 );
_DC r25610_GF_IsGateDCbyConstraint ( \21945_nR25610 , \21906 , \21944 );
buf \U$13134 ( \21946 , \21945_nR25610 );
and \U$13136 ( \21947 , \21765 , 1'b1 );
or \U$13138 ( \21948 , \21947 , 1'b0 );
buf \U$13139 ( \21949 , \21948 );
_DC r25642_GF_IsGateDCbyConstraint ( \21950_nR25642 , \21949 , \21944 );
buf \U$13140 ( \21951 , \21950_nR25642 );
and \U$13142 ( \21952 , \21783 , 1'b1 );
or \U$13144 ( \21953 , \21952 , 1'b0 );
buf \U$13145 ( \21954 , \21953 );
_DC r25644_GF_IsGateDCbyConstraint ( \21955_nR25644 , \21954 , \21944 );
buf \U$13146 ( \21956 , \21955_nR25644 );
nand \U$13147 ( \21957 , \21755 , \21750 );
and \U$13149 ( \21958 , \21957 , 1'b1 );
or \U$13151 ( \21959 , \21958 , 1'b0 );
buf \U$13152 ( \21960 , \21959 );
_DC r25646_GF_IsGateDCbyConstraint ( \21961_nR25646 , \21960 , \21944 );
buf \U$13153 ( \21962 , \21961_nR25646 );
not \U$13154 ( \21963 , \21858 );
and \U$13156 ( \21964 , \21963 , 1'b1 );
or \U$13158 ( \21965 , \21964 , 1'b0 );
buf \U$13159 ( \21966 , \21965 );
_DC r25614_GF_IsGateDCbyConstraint ( \21967_nR25614 , \21966 , \21944 );
buf \U$13160 ( \21968 , \21967_nR25614 );
not \U$13161 ( \21969 , \21853 );
not \U$13162 ( \21970 , \21969 );
and \U$13163 ( \21971 , RIde4c8e8_4009, \21970 );
buf \U$13164 ( \21972 , RIb7b96f8_244);
and \U$13165 ( \21973 , \21972 , \21969 );
or \U$13166 ( \21974 , \21971 , \21973 );
and \U$13168 ( \21975 , \21974 , 1'b1 );
or \U$13170 ( \21976 , \21975 , 1'b0 );
buf \U$13171 ( \21977 , \21976 );
_DC r25616_GF_IsGateDCbyConstraint ( \21978_nR25616 , \21977 , \21944 );
buf \U$13172 ( \21979 , \21978_nR25616 );
not \U$13173 ( \21980 , \21969 );
and \U$13174 ( \21981 , RIde4d6f8_4008, \21980 );
buf \U$13175 ( \21982 , RIb7c20c8_243);
and \U$13176 ( \21983 , \21982 , \21969 );
or \U$13177 ( \21984 , \21981 , \21983 );
and \U$13179 ( \21985 , \21984 , 1'b1 );
or \U$13181 ( \21986 , \21985 , 1'b0 );
buf \U$13182 ( \21987 , \21986 );
_DC r25618_GF_IsGateDCbyConstraint ( \21988_nR25618 , \21987 , \21944 );
buf \U$13183 ( \21989 , \21988_nR25618 );
not \U$13184 ( \21990 , \21969 );
and \U$13185 ( \21991 , RIde431f8_4020, \21990 );
buf \U$13186 ( \21992 , RIb7c5728_242);
and \U$13187 ( \21993 , \21992 , \21969 );
or \U$13188 ( \21994 , \21991 , \21993 );
and \U$13190 ( \21995 , \21994 , 1'b1 );
or \U$13192 ( \21996 , \21995 , 1'b0 );
buf \U$13193 ( \21997 , \21996 );
_DC r2561a_GF_IsGateDCbyConstraint ( \21998_nR2561a , \21997 , \21944 );
buf \U$13194 ( \21999 , \21998_nR2561a );
not \U$13195 ( \22000 , \21969 );
and \U$13196 ( \22001 , RIde43f90_4019, \22000 );
buf \U$13197 ( \22002 , RIb7c57a0_241);
and \U$13198 ( \22003 , \22002 , \21969 );
or \U$13199 ( \22004 , \22001 , \22003 );
and \U$13201 ( \22005 , \22004 , 1'b1 );
or \U$13203 ( \22006 , \22005 , 1'b0 );
buf \U$13204 ( \22007 , \22006 );
_DC r2561c_GF_IsGateDCbyConstraint ( \22008_nR2561c , \22007 , \21944 );
buf \U$13205 ( \22009 , \22008_nR2561c );
not \U$13206 ( \22010 , \21969 );
and \U$13207 ( \22011 , RIde44da0_4018, \22010 );
buf \U$13208 ( \22012 , RIb7c5818_240);
and \U$13209 ( \22013 , \22012 , \21969 );
or \U$13210 ( \22014 , \22011 , \22013 );
and \U$13212 ( \22015 , \22014 , 1'b1 );
or \U$13214 ( \22016 , \22015 , 1'b0 );
buf \U$13215 ( \22017 , \22016 );
_DC r2561e_GF_IsGateDCbyConstraint ( \22018_nR2561e , \22017 , \21944 );
buf \U$13216 ( \22019 , \22018_nR2561e );
not \U$13217 ( \22020 , \21969 );
and \U$13218 ( \22021 , RIde45ac0_4017, \22020 );
buf \U$13219 ( \22022 , RIb7c5890_239);
and \U$13220 ( \22023 , \22022 , \21969 );
or \U$13221 ( \22024 , \22021 , \22023 );
and \U$13223 ( \22025 , \22024 , 1'b1 );
or \U$13225 ( \22026 , \22025 , 1'b0 );
buf \U$13226 ( \22027 , \22026 );
_DC r25620_GF_IsGateDCbyConstraint ( \22028_nR25620 , \22027 , \21944 );
buf \U$13227 ( \22029 , \22028_nR25620 );
not \U$13228 ( \22030 , \21969 );
and \U$13229 ( \22031 , RIde468d0_4016, \22030 );
buf \U$13230 ( \22032 , RIb7c5908_238);
and \U$13231 ( \22033 , \22032 , \21969 );
or \U$13232 ( \22034 , \22031 , \22033 );
and \U$13234 ( \22035 , \22034 , 1'b1 );
or \U$13236 ( \22036 , \22035 , 1'b0 );
buf \U$13237 ( \22037 , \22036 );
_DC r25622_GF_IsGateDCbyConstraint ( \22038_nR25622 , \22037 , \21944 );
buf \U$13238 ( \22039 , \22038_nR25622 );
not \U$13239 ( \22040 , \21969 );
and \U$13240 ( \22041 , RIde4fb10_4005, \22040 );
buf \U$13241 ( \22042 , RIb7a09f0_266);
and \U$13242 ( \22043 , \22042 , \21969 );
or \U$13243 ( \22044 , \22041 , \22043 );
and \U$13245 ( \22045 , \22044 , 1'b1 );
or \U$13247 ( \22046 , \22045 , 1'b0 );
buf \U$13248 ( \22047 , \22046 );
_DC r25612_GF_IsGateDCbyConstraint ( \22048_nR25612 , \22047 , \21944 );
buf \U$13249 ( \22049 , \22048_nR25612 );
not \U$13250 ( \22050 , \21969 );
and \U$13251 ( \22051 , RIde49300_4013, \22050 );
buf \U$13252 ( \22052 , RIb7a0a68_265);
and \U$13253 ( \22053 , \22052 , \21969 );
or \U$13254 ( \22054 , \22051 , \22053 );
and \U$13256 ( \22055 , \22054 , 1'b1 );
or \U$13258 ( \22056 , \22055 , 1'b0 );
buf \U$13259 ( \22057 , \22056 );
_DC r25624_GF_IsGateDCbyConstraint ( \22058_nR25624 , \22057 , \21944 );
buf \U$13260 ( \22059 , \22058_nR25624 );
not \U$13261 ( \22060 , \21969 );
and \U$13262 ( \22061 , RIde4a020_4012, \22060 );
buf \U$13263 ( \22062 , RIb7a0ae0_264);
and \U$13264 ( \22063 , \22062 , \21969 );
or \U$13265 ( \22064 , \22061 , \22063 );
and \U$13267 ( \22065 , \22064 , 1'b1 );
or \U$13269 ( \22066 , \22065 , 1'b0 );
buf \U$13270 ( \22067 , \22066 );
_DC r25626_GF_IsGateDCbyConstraint ( \22068_nR25626 , \22067 , \21944 );
buf \U$13271 ( \22069 , \22068_nR25626 );
not \U$13272 ( \22070 , \21969 );
and \U$13273 ( \22071 , RIde4ae30_4011, \22070 );
buf \U$13274 ( \22072 , RIb7a0b58_263);
and \U$13275 ( \22073 , \22072 , \21969 );
or \U$13276 ( \22074 , \22071 , \22073 );
and \U$13278 ( \22075 , \22074 , 1'b1 );
or \U$13280 ( \22076 , \22075 , 1'b0 );
buf \U$13281 ( \22077 , \22076 );
_DC r25628_GF_IsGateDCbyConstraint ( \22078_nR25628 , \22077 , \21944 );
buf \U$13282 ( \22079 , \22078_nR25628 );
not \U$13283 ( \22080 , \21969 );
and \U$13284 ( \22081 , RIde4bb50_4010, \22080 );
buf \U$13285 ( \22082 , RIb7a0bd0_262);
and \U$13286 ( \22083 , \22082 , \21969 );
or \U$13287 ( \22084 , \22081 , \22083 );
and \U$13289 ( \22085 , \22084 , 1'b1 );
or \U$13291 ( \22086 , \22085 , 1'b0 );
buf \U$13292 ( \22087 , \22086 );
_DC r2562a_GF_IsGateDCbyConstraint ( \22088_nR2562a , \22087 , \21944 );
buf \U$13293 ( \22089 , \22088_nR2562a );
buf \U$13294 ( \22090 , \21816 );
not \U$13295 ( \22091 , RIb839b90_145);
and \U$13296 ( \22092 , RIb839848_152, \22091 );
and \U$13297 ( \22093 , RIb8396e0_155, RIb839b90_145);
or \U$13298 ( \22094 , \22092 , \22093 );
not \U$13299 ( \22095 , \22094 );
not \U$13300 ( \22096 , \22095 );
buf \U$13301 ( \22097 , \22096 );
buf \U$13302 ( \22098 , \22097 );
nand \U$13303 ( \22099 , \22090 , \22098 );
buf \U$13304 ( \22100 , \8826 );
buf \U$13305 ( \22101 , \21696 );
nand \U$13306 ( \22102 , \22100 , \22101 );
nand \U$13307 ( \22103 , \22099 , \22102 );
buf \U$13308 ( \22104 , \22103 );
buf \U$13309 ( \22105 , \22104 );
not \U$13310 ( \22106 , \22105 );
and \U$13311 ( \22107 , RIdbee210_3713, \22106 );
not \U$13312 ( \22108 , RIdbee210_3713);
buf \U$13313 ( \22109 , RIe667bb0_6885);
buf \U$13314 ( \22110 , \22109 );
buf \U$13315 ( \22111 , RIe667f70_6886);
not \U$13316 ( \22112 , \22111 );
not \U$13317 ( \22113 , \22112 );
or \U$13318 ( \22114 , \22110 , \22113 );
not \U$13319 ( \22115 , \22114 );
nand \U$13320 ( \22116 , \22102 , \22115 );
buf \U$13321 ( \22117 , RIea91768_6889);
not \U$13322 ( \22118 , \22117 );
not \U$13323 ( \22119 , RIeab7058_6894);
not \U$13324 ( \22120 , \22119 );
buf \U$13325 ( \22121 , \22120 );
not \U$13326 ( \22122 , \22121 );
not \U$13327 ( \22123 , \22102 );
and \U$13328 ( \22124 , \22118 , \22122 , \22123 );
not \U$13329 ( \22125 , \22124 );
buf \U$13330 ( \22126 , \22125 );
and \U$13331 ( \22127 , \22116 , \22126 );
not \U$13332 ( \22128 , \22127 );
or \U$13333 ( \22129 , \22108 , \22128 );
not \U$13334 ( \22130 , \22116 );
buf \U$13335 ( \22131 , RIb87eb00_69);
buf \U$13336 ( \22132 , \22131 );
and \U$13337 ( \22133 , \22130 , \22132 );
buf \U$13338 ( \22134 , RIb7c5980_237);
buf \U$13339 ( \22135 , \22134 );
not \U$13340 ( \22136 , \22126 );
and \U$13341 ( \22137 , \22135 , \22136 );
nor \U$13342 ( \22138 , \22133 , \22137 );
nand \U$13343 ( \22139 , \22129 , \22138 );
and \U$13344 ( \22140 , \22139 , \22105 );
or \U$13345 ( \22141 , \22107 , \22140 );
and \U$13347 ( \22142 , \22141 , 1'b1 );
or \U$13349 ( \22143 , \22142 , 1'b0 );
buf \U$13350 ( \22144 , \22143 );
_DC r253fc_GF_IsGateDCbyConstraint ( \22145_nR253fc , \22144 , \21944 );
buf \U$13351 ( \22146 , \22145_nR253fc );
not \U$13352 ( \22147 , \22105 );
and \U$13353 ( \22148 , RIdbecc08_3714, \22147 );
not \U$13354 ( \22149 , RIdbecc08_3714);
not \U$13355 ( \22150 , \22117 );
not \U$13356 ( \22151 , \22121 );
and \U$13357 ( \22152 , \22150 , \22151 , \22123 );
not \U$13358 ( \22153 , \22152 );
buf \U$13359 ( \22154 , \22153 );
and \U$13360 ( \22155 , \22116 , \22154 );
not \U$13361 ( \22156 , \22155 );
or \U$13362 ( \22157 , \22149 , \22156 );
buf \U$13363 ( \22158 , \22130 );
buf \U$13364 ( \22159 , RIb87eb78_68);
and \U$13365 ( \22160 , \22158 , \22159 );
buf \U$13366 ( \22161 , RIb7c59f8_236);
buf \U$13367 ( \22162 , \22161 );
buf \U$13368 ( \22163 , \22125 );
not \U$13369 ( \22164 , \22163 );
and \U$13370 ( \22165 , \22162 , \22164 );
nor \U$13371 ( \22166 , \22160 , \22165 );
nand \U$13372 ( \22167 , \22157 , \22166 );
and \U$13373 ( \22168 , \22167 , \22105 );
or \U$13374 ( \22169 , \22148 , \22168 );
and \U$13376 ( \22170 , \22169 , 1'b1 );
or \U$13378 ( \22171 , \22170 , 1'b0 );
buf \U$13379 ( \22172 , \22171 );
_DC r25412_GF_IsGateDCbyConstraint ( \22173_nR25412 , \22172 , \21944 );
buf \U$13380 ( \22174 , \22173_nR25412 );
not \U$13381 ( \22175 , \22105 );
and \U$13382 ( \22176 , RIdbebab0_3715, \22175 );
not \U$13383 ( \22177 , RIdbebab0_3715);
or \U$13384 ( \22178 , \22177 , \22128 );
buf \U$13385 ( \22179 , RIb87ebf0_67);
buf \U$13386 ( \22180 , \22179 );
and \U$13387 ( \22181 , \22158 , \22180 );
buf \U$13388 ( \22182 , RIb7c5a70_235);
buf \U$13389 ( \22183 , \22182 );
not \U$13390 ( \22184 , \22126 );
and \U$13391 ( \22185 , \22183 , \22184 );
nor \U$13392 ( \22186 , \22181 , \22185 );
nand \U$13393 ( \22187 , \22178 , \22186 );
and \U$13394 ( \22188 , \22187 , \22105 );
or \U$13395 ( \22189 , \22176 , \22188 );
and \U$13397 ( \22190 , \22189 , 1'b1 );
or \U$13399 ( \22191 , \22190 , 1'b0 );
buf \U$13400 ( \22192 , \22191 );
_DC r25428_GF_IsGateDCbyConstraint ( \22193_nR25428 , \22192 , \21944 );
buf \U$13401 ( \22194 , \22193_nR25428 );
buf \U$13402 ( \22195 , \22103 );
buf \U$13403 ( \22196 , \22195 );
not \U$13404 ( \22197 , \22196 );
and \U$13405 ( \22198 , RIdbea4a8_3716, \22197 );
not \U$13406 ( \22199 , RIdbea4a8_3716);
or \U$13407 ( \22200 , \22199 , \22156 );
buf \U$13408 ( \22201 , \22130 );
buf \U$13409 ( \22202 , RIb882ca0_66);
buf \U$13410 ( \22203 , \22202 );
and \U$13411 ( \22204 , \22201 , \22203 );
buf \U$13412 ( \22205 , RIb7cade0_234);
buf \U$13413 ( \22206 , \22205 );
not \U$13414 ( \22207 , \22154 );
and \U$13415 ( \22208 , \22206 , \22207 );
nor \U$13416 ( \22209 , \22204 , \22208 );
nand \U$13417 ( \22210 , \22200 , \22209 );
and \U$13418 ( \22211 , \22210 , \22196 );
or \U$13419 ( \22212 , \22198 , \22211 );
and \U$13421 ( \22213 , \22212 , 1'b1 );
or \U$13423 ( \22214 , \22213 , 1'b0 );
buf \U$13424 ( \22215 , \22214 );
_DC r2543e_GF_IsGateDCbyConstraint ( \22216_nR2543e , \22215 , \21944 );
buf \U$13425 ( \22217 , \22216_nR2543e );
not \U$13426 ( \22218 , \22196 );
and \U$13427 ( \22219 , RIdbe9350_3717, \22218 );
not \U$13428 ( \22220 , RIdbe9350_3717);
not \U$13429 ( \22221 , \22127 );
or \U$13430 ( \22222 , \22220 , \22221 );
buf \U$13431 ( \22223 , RIb885310_65);
buf \U$13432 ( \22224 , \22223 );
and \U$13433 ( \22225 , \22130 , \22224 );
buf \U$13434 ( \22226 , RIb7cae58_233);
buf \U$13435 ( \22227 , \22226 );
not \U$13436 ( \22228 , \22163 );
and \U$13437 ( \22229 , \22227 , \22228 );
nor \U$13438 ( \22230 , \22225 , \22229 );
nand \U$13439 ( \22231 , \22222 , \22230 );
and \U$13440 ( \22232 , \22231 , \22196 );
or \U$13441 ( \22233 , \22219 , \22232 );
and \U$13443 ( \22234 , \22233 , 1'b1 );
or \U$13445 ( \22235 , \22234 , 1'b0 );
buf \U$13446 ( \22236 , \22235 );
_DC r25454_GF_IsGateDCbyConstraint ( \22237_nR25454 , \22236 , \21944 );
buf \U$13447 ( \22238 , \22237_nR25454 );
not \U$13448 ( \22239 , \22105 );
and \U$13449 ( \22240 , RIdbe7d48_3718, \22239 );
not \U$13450 ( \22241 , RIdbe7d48_3718);
not \U$13451 ( \22242 , \22155 );
or \U$13452 ( \22243 , \22241 , \22242 );
buf \U$13453 ( \22244 , \22130 );
buf \U$13454 ( \22245 , RIb885388_64);
buf \U$13455 ( \22246 , \22245 );
and \U$13456 ( \22247 , \22244 , \22246 );
buf \U$13457 ( \22248 , RIb7caed0_232);
buf \U$13458 ( \22249 , \22248 );
not \U$13459 ( \22250 , \22117 );
not \U$13460 ( \22251 , \22121 );
and \U$13461 ( \22252 , \22250 , \22251 , \22123 );
not \U$13462 ( \22253 , \22252 );
buf \U$13463 ( \22254 , \22253 );
not \U$13464 ( \22255 , \22254 );
and \U$13465 ( \22256 , \22249 , \22255 );
nor \U$13466 ( \22257 , \22247 , \22256 );
nand \U$13467 ( \22258 , \22243 , \22257 );
and \U$13468 ( \22259 , \22258 , \22105 );
or \U$13469 ( \22260 , \22240 , \22259 );
and \U$13471 ( \22261 , \22260 , 1'b1 );
or \U$13473 ( \22262 , \22261 , 1'b0 );
buf \U$13474 ( \22263 , \22262 );
_DC r2546a_GF_IsGateDCbyConstraint ( \22264_nR2546a , \22263 , \21944 );
buf \U$13475 ( \22265 , \22264_nR2546a );
not \U$13476 ( \22266 , \22105 );
and \U$13477 ( \22267 , RIdbe6bf0_3719, \22266 );
not \U$13478 ( \22268 , RIdbe6bf0_3719);
not \U$13479 ( \22269 , \22127 );
or \U$13480 ( \22270 , \22268 , \22269 );
buf \U$13481 ( \22271 , RIb885400_63);
buf \U$13482 ( \22272 , \22271 );
and \U$13483 ( \22273 , \22130 , \22272 );
buf \U$13484 ( \22274 , RIb7caf48_231);
buf \U$13485 ( \22275 , \22274 );
not \U$13486 ( \22276 , \22154 );
and \U$13487 ( \22277 , \22275 , \22276 );
nor \U$13488 ( \22278 , \22273 , \22277 );
nand \U$13489 ( \22279 , \22270 , \22278 );
and \U$13490 ( \22280 , \22279 , \22105 );
or \U$13491 ( \22281 , \22267 , \22280 );
and \U$13493 ( \22282 , \22281 , 1'b1 );
or \U$13495 ( \22283 , \22282 , 1'b0 );
buf \U$13496 ( \22284 , \22283 );
_DC r25474_GF_IsGateDCbyConstraint ( \22285_nR25474 , \22284 , \21944 );
buf \U$13497 ( \22286 , \22285_nR25474 );
not \U$13498 ( \22287 , \22105 );
and \U$13499 ( \22288 , RIdbe5a98_3720, \22287 );
not \U$13500 ( \22289 , RIdbe5a98_3720);
or \U$13501 ( \22290 , \22289 , \22156 );
not \U$13502 ( \22291 , \22116 );
buf \U$13503 ( \22292 , RIb885478_62);
and \U$13504 ( \22293 , \22291 , \22292 );
buf \U$13505 ( \22294 , RIb7cafc0_230);
buf \U$13506 ( \22295 , \22294 );
buf \U$13507 ( \22296 , \22253 );
not \U$13508 ( \22297 , \22296 );
and \U$13509 ( \22298 , \22295 , \22297 );
nor \U$13510 ( \22299 , \22293 , \22298 );
nand \U$13511 ( \22300 , \22290 , \22299 );
and \U$13512 ( \22301 , \22300 , \22105 );
or \U$13513 ( \22302 , \22288 , \22301 );
and \U$13515 ( \22303 , \22302 , 1'b1 );
or \U$13517 ( \22304 , \22303 , 1'b0 );
buf \U$13518 ( \22305 , \22304 );
_DC r25476_GF_IsGateDCbyConstraint ( \22306_nR25476 , \22305 , \21944 );
buf \U$13519 ( \22307 , \22306_nR25476 );
buf \U$13520 ( \22308 , \22104 );
not \U$13521 ( \22309 , \22308 );
and \U$13522 ( \22310 , RIdbe4490_3721, \22309 );
not \U$13523 ( \22311 , RIdbe4490_3721);
or \U$13524 ( \22312 , \22311 , \22156 );
buf \U$13525 ( \22313 , RIb8854f0_61);
buf \U$13526 ( \22314 , \22313 );
and \U$13527 ( \22315 , \22244 , \22314 );
buf \U$13528 ( \22316 , RIb7cb038_229);
buf \U$13529 ( \22317 , \22316 );
buf \U$13530 ( \22318 , \22253 );
not \U$13531 ( \22319 , \22318 );
and \U$13532 ( \22320 , \22317 , \22319 );
nor \U$13533 ( \22321 , \22315 , \22320 );
nand \U$13534 ( \22322 , \22312 , \22321 );
and \U$13535 ( \22323 , \22322 , \22308 );
or \U$13536 ( \22324 , \22310 , \22323 );
and \U$13538 ( \22325 , \22324 , 1'b1 );
or \U$13540 ( \22326 , \22325 , 1'b0 );
buf \U$13541 ( \22327 , \22326 );
_DC r25478_GF_IsGateDCbyConstraint ( \22328_nR25478 , \22327 , \21944 );
buf \U$13542 ( \22329 , \22328_nR25478 );
not \U$13543 ( \22330 , \22196 );
and \U$13544 ( \22331 , RIdbe3338_3722, \22330 );
not \U$13545 ( \22332 , RIdbe3338_3722);
or \U$13546 ( \22333 , \22332 , \22156 );
buf \U$13547 ( \22334 , RIb885568_60);
buf \U$13548 ( \22335 , \22334 );
and \U$13549 ( \22336 , \22130 , \22335 );
buf \U$13550 ( \22337 , RIb7cb0b0_228);
buf \U$13551 ( \22338 , \22337 );
buf \U$13552 ( \22339 , \22153 );
not \U$13553 ( \22340 , \22339 );
and \U$13554 ( \22341 , \22338 , \22340 );
nor \U$13555 ( \22342 , \22336 , \22341 );
nand \U$13556 ( \22343 , \22333 , \22342 );
and \U$13557 ( \22344 , \22343 , \22196 );
or \U$13558 ( \22345 , \22331 , \22344 );
and \U$13560 ( \22346 , \22345 , 1'b1 );
or \U$13562 ( \22347 , \22346 , 1'b0 );
buf \U$13563 ( \22348 , \22347 );
_DC r2547a_GF_IsGateDCbyConstraint ( \22349_nR2547a , \22348 , \21944 );
buf \U$13564 ( \22350 , \22349_nR2547a );
not \U$13565 ( \22351 , \22105 );
and \U$13566 ( \22352 , RIdbe1d30_3723, \22351 );
not \U$13567 ( \22353 , RIdbe1d30_3723);
not \U$13568 ( \22354 , \22127 );
or \U$13569 ( \22355 , \22353 , \22354 );
buf \U$13570 ( \22356 , RIb8855e0_59);
buf \U$13571 ( \22357 , \22356 );
and \U$13572 ( \22358 , \22158 , \22357 );
buf \U$13573 ( \22359 , RIb7cb128_227);
buf \U$13574 ( \22360 , \22359 );
not \U$13575 ( \22361 , \22254 );
and \U$13576 ( \22362 , \22360 , \22361 );
nor \U$13577 ( \22363 , \22358 , \22362 );
nand \U$13578 ( \22364 , \22355 , \22363 );
and \U$13579 ( \22365 , \22364 , \22105 );
or \U$13580 ( \22366 , \22352 , \22365 );
and \U$13582 ( \22367 , \22366 , 1'b1 );
or \U$13584 ( \22368 , \22367 , 1'b0 );
buf \U$13585 ( \22369 , \22368 );
_DC r253fe_GF_IsGateDCbyConstraint ( \22370_nR253fe , \22369 , \21944 );
buf \U$13586 ( \22371 , \22370_nR253fe );
not \U$13587 ( \22372 , \22308 );
and \U$13588 ( \22373 , RIdbe0bd8_3724, \22372 );
not \U$13589 ( \22374 , RIdbe0bd8_3724);
or \U$13590 ( \22375 , \22374 , \22221 );
buf \U$13591 ( \22376 , RIb885658_58);
buf \U$13592 ( \22377 , \22376 );
and \U$13593 ( \22378 , \22158 , \22377 );
buf \U$13594 ( \22379 , RIb7d00d8_226);
buf \U$13595 ( \22380 , \22379 );
not \U$13596 ( \22381 , \22296 );
and \U$13597 ( \22382 , \22380 , \22381 );
nor \U$13598 ( \22383 , \22378 , \22382 );
nand \U$13599 ( \22384 , \22375 , \22383 );
and \U$13600 ( \22385 , \22384 , \22308 );
or \U$13601 ( \22386 , \22373 , \22385 );
and \U$13603 ( \22387 , \22386 , 1'b1 );
or \U$13605 ( \22388 , \22387 , 1'b0 );
buf \U$13606 ( \22389 , \22388 );
_DC r25400_GF_IsGateDCbyConstraint ( \22390_nR25400 , \22389 , \21944 );
buf \U$13607 ( \22391 , \22390_nR25400 );
not \U$13608 ( \22392 , \22105 );
and \U$13609 ( \22393 , RIdaab098_3725, \22392 );
not \U$13610 ( \22394 , RIdaab098_3725);
not \U$13611 ( \22395 , \22127 );
or \U$13612 ( \22396 , \22394 , \22395 );
buf \U$13613 ( \22397 , RIb8856d0_57);
buf \U$13614 ( \22398 , \22397 );
and \U$13615 ( \22399 , \22158 , \22398 );
buf \U$13616 ( \22400 , RIb8263d8_225);
buf \U$13617 ( \22401 , \22400 );
not \U$13618 ( \22402 , \22318 );
and \U$13619 ( \22403 , \22401 , \22402 );
nor \U$13620 ( \22404 , \22399 , \22403 );
nand \U$13621 ( \22405 , \22396 , \22404 );
and \U$13622 ( \22406 , \22405 , \22105 );
or \U$13623 ( \22407 , \22393 , \22406 );
and \U$13625 ( \22408 , \22407 , 1'b1 );
or \U$13627 ( \22409 , \22408 , 1'b0 );
buf \U$13628 ( \22410 , \22409 );
_DC r25402_GF_IsGateDCbyConstraint ( \22411_nR25402 , \22410 , \21944 );
buf \U$13629 ( \22412 , \22411_nR25402 );
not \U$13630 ( \22413 , \22105 );
and \U$13631 ( \22414 , RIdaaf0d0_3726, \22413 );
not \U$13632 ( \22415 , RIdaaf0d0_3726);
or \U$13633 ( \22416 , \22415 , \22242 );
buf \U$13634 ( \22417 , RIb885748_56);
buf \U$13635 ( \22418 , \22417 );
and \U$13636 ( \22419 , \22158 , \22418 );
buf \U$13637 ( \22420 , RIb826e28_224);
buf \U$13638 ( \22421 , \22420 );
buf \U$13639 ( \22422 , \22153 );
not \U$13640 ( \22423 , \22422 );
and \U$13641 ( \22424 , \22421 , \22423 );
nor \U$13642 ( \22425 , \22419 , \22424 );
nand \U$13643 ( \22426 , \22416 , \22425 );
and \U$13644 ( \22427 , \22426 , \22105 );
or \U$13645 ( \22428 , \22414 , \22427 );
and \U$13647 ( \22429 , \22428 , 1'b1 );
or \U$13649 ( \22430 , \22429 , 1'b0 );
buf \U$13650 ( \22431 , \22430 );
_DC r25404_GF_IsGateDCbyConstraint ( \22432_nR25404 , \22431 , \21944 );
buf \U$13651 ( \22433 , \22432_nR25404 );
not \U$13652 ( \22434 , \22308 );
and \U$13653 ( \22435 , RIdab2fa0_3727, \22434 );
not \U$13654 ( \22436 , RIdab2fa0_3727);
or \U$13655 ( \22437 , \22436 , \22242 );
buf \U$13656 ( \22438 , RIb8857c0_55);
and \U$13657 ( \22439 , \22158 , \22438 );
buf \U$13658 ( \22440 , RIb826ea0_223);
buf \U$13659 ( \22441 , \22440 );
not \U$13660 ( \22442 , \22339 );
and \U$13661 ( \22443 , \22441 , \22442 );
nor \U$13662 ( \22444 , \22439 , \22443 );
nand \U$13663 ( \22445 , \22437 , \22444 );
and \U$13664 ( \22446 , \22445 , \22308 );
or \U$13665 ( \22447 , \22435 , \22446 );
and \U$13667 ( \22448 , \22447 , 1'b1 );
or \U$13669 ( \22449 , \22448 , 1'b0 );
buf \U$13670 ( \22450 , \22449 );
_DC r25406_GF_IsGateDCbyConstraint ( \22451_nR25406 , \22450 , \21944 );
buf \U$13671 ( \22452 , \22451_nR25406 );
not \U$13672 ( \22453 , \22196 );
and \U$13673 ( \22454 , RIdab8e50_3728, \22453 );
not \U$13674 ( \22455 , RIdab8e50_3728);
or \U$13675 ( \22456 , \22455 , \22128 );
buf \U$13676 ( \22457 , RIb885838_54);
buf \U$13677 ( \22458 , \22457 );
and \U$13678 ( \22459 , \22201 , \22458 );
buf \U$13679 ( \22460 , RIb826f18_222);
buf \U$13680 ( \22461 , \22460 );
not \U$13681 ( \22462 , \22154 );
and \U$13682 ( \22463 , \22461 , \22462 );
nor \U$13683 ( \22464 , \22459 , \22463 );
nand \U$13684 ( \22465 , \22456 , \22464 );
and \U$13685 ( \22466 , \22465 , \22196 );
or \U$13686 ( \22467 , \22454 , \22466 );
and \U$13688 ( \22468 , \22467 , 1'b1 );
or \U$13690 ( \22469 , \22468 , 1'b0 );
buf \U$13691 ( \22470 , \22469 );
_DC r25408_GF_IsGateDCbyConstraint ( \22471_nR25408 , \22470 , \21944 );
buf \U$13692 ( \22472 , \22471_nR25408 );
not \U$13693 ( \22473 , \22196 );
and \U$13694 ( \22474 , RIdabcf00_3729, \22473 );
not \U$13695 ( \22475 , RIdabcf00_3729);
or \U$13696 ( \22476 , \22475 , \22354 );
buf \U$13697 ( \22477 , RIb8858b0_53);
buf \U$13698 ( \22478 , \22477 );
and \U$13699 ( \22479 , \22158 , \22478 );
buf \U$13700 ( \22480 , RIb826f90_221);
buf \U$13701 ( \22481 , \22480 );
not \U$13702 ( \22482 , \22163 );
and \U$13703 ( \22483 , \22481 , \22482 );
nor \U$13704 ( \22484 , \22479 , \22483 );
nand \U$13705 ( \22485 , \22476 , \22484 );
and \U$13706 ( \22486 , \22485 , \22196 );
or \U$13707 ( \22487 , \22474 , \22486 );
and \U$13709 ( \22488 , \22487 , 1'b1 );
or \U$13711 ( \22489 , \22488 , 1'b0 );
buf \U$13712 ( \22490 , \22489 );
_DC r2540a_GF_IsGateDCbyConstraint ( \22491_nR2540a , \22490 , \21944 );
buf \U$13713 ( \22492 , \22491_nR2540a );
not \U$13714 ( \22493 , \22308 );
and \U$13715 ( \22494 , RIdac3788_3730, \22493 );
not \U$13716 ( \22495 , RIdac3788_3730);
or \U$13717 ( \22496 , \22495 , \22221 );
buf \U$13718 ( \22497 , RIb885928_52);
buf \U$13719 ( \22498 , \22497 );
and \U$13720 ( \22499 , \22158 , \22498 );
buf \U$13721 ( \22500 , RIb8293a8_220);
buf \U$13722 ( \22501 , \22500 );
buf \U$13723 ( \22502 , \22125 );
not \U$13724 ( \22503 , \22502 );
and \U$13725 ( \22504 , \22501 , \22503 );
nor \U$13726 ( \22505 , \22499 , \22504 );
nand \U$13727 ( \22506 , \22496 , \22505 );
and \U$13728 ( \22507 , \22506 , \22308 );
or \U$13729 ( \22508 , \22494 , \22507 );
and \U$13731 ( \22509 , \22508 , 1'b1 );
or \U$13733 ( \22510 , \22509 , 1'b0 );
buf \U$13734 ( \22511 , \22510 );
_DC r2540c_GF_IsGateDCbyConstraint ( \22512_nR2540c , \22511 , \21944 );
buf \U$13735 ( \22513 , \22512_nR2540c );
not \U$13736 ( \22514 , \22196 );
and \U$13737 ( \22515 , RIdac8eb8_3731, \22514 );
not \U$13738 ( \22516 , RIdac8eb8_3731);
or \U$13739 ( \22517 , \22516 , \22395 );
buf \U$13740 ( \22518 , RIb8859a0_51);
buf \U$13741 ( \22519 , \22518 );
and \U$13742 ( \22520 , \22244 , \22519 );
buf \U$13743 ( \22521 , RIb829420_219);
buf \U$13744 ( \22522 , \22521 );
not \U$13745 ( \22523 , \22163 );
and \U$13746 ( \22524 , \22522 , \22523 );
nor \U$13747 ( \22525 , \22520 , \22524 );
nand \U$13748 ( \22526 , \22517 , \22525 );
and \U$13749 ( \22527 , \22526 , \22196 );
or \U$13750 ( \22528 , \22515 , \22527 );
and \U$13752 ( \22529 , \22528 , 1'b1 );
or \U$13754 ( \22530 , \22529 , 1'b0 );
buf \U$13755 ( \22531 , \22530 );
_DC r2540e_GF_IsGateDCbyConstraint ( \22532_nR2540e , \22531 , \21944 );
buf \U$13756 ( \22533 , \22532_nR2540e );
not \U$13757 ( \22534 , \22105 );
and \U$13758 ( \22535 , RIdacf650_3732, \22534 );
not \U$13759 ( \22536 , RIdacf650_3732);
or \U$13760 ( \22537 , \22536 , \22269 );
buf \U$13761 ( \22538 , RIb885a18_50);
buf \U$13762 ( \22539 , \22538 );
and \U$13763 ( \22540 , \22158 , \22539 );
buf \U$13764 ( \22541 , RIb829498_218);
buf \U$13765 ( \22542 , \22541 );
not \U$13766 ( \22543 , \22126 );
and \U$13767 ( \22544 , \22542 , \22543 );
nor \U$13768 ( \22545 , \22540 , \22544 );
nand \U$13769 ( \22546 , \22537 , \22545 );
and \U$13770 ( \22547 , \22546 , \22105 );
or \U$13771 ( \22548 , \22535 , \22547 );
and \U$13773 ( \22549 , \22548 , 1'b1 );
or \U$13775 ( \22550 , \22549 , 1'b0 );
buf \U$13776 ( \22551 , \22550 );
_DC r25410_GF_IsGateDCbyConstraint ( \22552_nR25410 , \22551 , \21944 );
buf \U$13777 ( \22553 , \22552_nR25410 );
not \U$13778 ( \22554 , \22308 );
and \U$13779 ( \22555 , RIdad4fd8_3733, \22554 );
not \U$13780 ( \22556 , RIdad4fd8_3733);
or \U$13781 ( \22557 , \22556 , \22156 );
buf \U$13782 ( \22558 , RIb885a90_49);
buf \U$13783 ( \22559 , \22558 );
and \U$13784 ( \22560 , \22201 , \22559 );
buf \U$13785 ( \22561 , RIb829510_217);
buf \U$13786 ( \22562 , \22561 );
not \U$13787 ( \22563 , \22502 );
and \U$13788 ( \22564 , \22562 , \22563 );
nor \U$13789 ( \22565 , \22560 , \22564 );
nand \U$13790 ( \22566 , \22557 , \22565 );
and \U$13791 ( \22567 , \22566 , \22308 );
or \U$13792 ( \22568 , \22555 , \22567 );
and \U$13794 ( \22569 , \22568 , 1'b1 );
or \U$13796 ( \22570 , \22569 , 1'b0 );
buf \U$13797 ( \22571 , \22570 );
_DC r25414_GF_IsGateDCbyConstraint ( \22572_nR25414 , \22571 , \21944 );
buf \U$13798 ( \22573 , \22572_nR25414 );
not \U$13799 ( \22574 , \22196 );
and \U$13800 ( \22575 , RIdadaf00_3734, \22574 );
not \U$13801 ( \22576 , RIdadaf00_3734);
or \U$13802 ( \22577 , \22576 , \22242 );
buf \U$13803 ( \22578 , RIb885b08_48);
buf \U$13804 ( \22579 , \22578 );
and \U$13805 ( \22580 , \22201 , \22579 );
buf \U$13806 ( \22581 , RIb829588_216);
buf \U$13807 ( \22582 , \22581 );
not \U$13808 ( \22583 , \22254 );
and \U$13809 ( \22584 , \22582 , \22583 );
nor \U$13810 ( \22585 , \22580 , \22584 );
nand \U$13811 ( \22586 , \22577 , \22585 );
and \U$13812 ( \22587 , \22586 , \22196 );
or \U$13813 ( \22588 , \22575 , \22587 );
and \U$13815 ( \22589 , \22588 , 1'b1 );
or \U$13817 ( \22590 , \22589 , 1'b0 );
buf \U$13818 ( \22591 , \22590 );
_DC r25416_GF_IsGateDCbyConstraint ( \22592_nR25416 , \22591 , \21944 );
buf \U$13819 ( \22593 , \22592_nR25416 );
not \U$13820 ( \22594 , \22196 );
and \U$13821 ( \22595 , RIdae2610_3735, \22594 );
not \U$13822 ( \22596 , RIdae2610_3735);
or \U$13823 ( \22597 , \22596 , \22269 );
buf \U$13824 ( \22598 , RIb885b80_47);
buf \U$13825 ( \22599 , \22598 );
and \U$13826 ( \22600 , \22244 , \22599 );
buf \U$13827 ( \22601 , RIb829600_215);
buf \U$13828 ( \22602 , \22601 );
not \U$13829 ( \22603 , \22296 );
and \U$13830 ( \22604 , \22602 , \22603 );
nor \U$13831 ( \22605 , \22600 , \22604 );
nand \U$13832 ( \22606 , \22597 , \22605 );
and \U$13833 ( \22607 , \22606 , \22196 );
or \U$13834 ( \22608 , \22595 , \22607 );
and \U$13836 ( \22609 , \22608 , 1'b1 );
or \U$13838 ( \22610 , \22609 , 1'b0 );
buf \U$13839 ( \22611 , \22610 );
_DC r25418_GF_IsGateDCbyConstraint ( \22612_nR25418 , \22611 , \21944 );
buf \U$13840 ( \22613 , \22612_nR25418 );
not \U$13841 ( \22614 , \22308 );
and \U$13842 ( \22615 , RIdae8268_3736, \22614 );
not \U$13843 ( \22616 , RIdae8268_3736);
or \U$13844 ( \22617 , \22616 , \22156 );
buf \U$13845 ( \22618 , RIb885bf8_46);
buf \U$13846 ( \22619 , \22618 );
and \U$13847 ( \22620 , \22201 , \22619 );
buf \U$13848 ( \22621 , RIb829678_214);
buf \U$13849 ( \22622 , \22621 );
not \U$13850 ( \22623 , \22318 );
and \U$13851 ( \22624 , \22622 , \22623 );
nor \U$13852 ( \22625 , \22620 , \22624 );
nand \U$13853 ( \22626 , \22617 , \22625 );
and \U$13854 ( \22627 , \22626 , \22308 );
or \U$13855 ( \22628 , \22615 , \22627 );
and \U$13857 ( \22629 , \22628 , 1'b1 );
or \U$13859 ( \22630 , \22629 , 1'b0 );
buf \U$13860 ( \22631 , \22630 );
_DC r2541a_GF_IsGateDCbyConstraint ( \22632_nR2541a , \22631 , \21944 );
buf \U$13861 ( \22633 , \22632_nR2541a );
not \U$13862 ( \22634 , \22105 );
and \U$13863 ( \22635 , RIdaef720_3737, \22634 );
not \U$13864 ( \22636 , RIdaef720_3737);
or \U$13865 ( \22637 , \22636 , \22156 );
not \U$13866 ( \22638 , \22116 );
buf \U$13867 ( \22639 , RIb885c70_45);
buf \U$13868 ( \22640 , \22639 );
and \U$13869 ( \22641 , \22638 , \22640 );
buf \U$13870 ( \22642 , RIb8296f0_213);
buf \U$13871 ( \22643 , \22642 );
not \U$13872 ( \22644 , \22254 );
and \U$13873 ( \22645 , \22643 , \22644 );
nor \U$13874 ( \22646 , \22641 , \22645 );
nand \U$13875 ( \22647 , \22637 , \22646 );
and \U$13876 ( \22648 , \22647 , \22105 );
or \U$13877 ( \22649 , \22635 , \22648 );
and \U$13879 ( \22650 , \22649 , 1'b1 );
or \U$13881 ( \22651 , \22650 , 1'b0 );
buf \U$13882 ( \22652 , \22651 );
_DC r2541c_GF_IsGateDCbyConstraint ( \22653_nR2541c , \22652 , \21944 );
buf \U$13883 ( \22654 , \22653_nR2541c );
not \U$13884 ( \22655 , \22105 );
and \U$13885 ( \22656 , RIdaf4e50_3738, \22655 );
not \U$13886 ( \22657 , RIdaf4e50_3738);
or \U$13887 ( \22658 , \22657 , \22242 );
buf \U$13888 ( \22659 , RIb885ce8_44);
buf \U$13889 ( \22660 , \22659 );
and \U$13890 ( \22661 , \22201 , \22660 );
buf \U$13891 ( \22662 , RIb82dae8_212);
buf \U$13892 ( \22663 , \22662 );
not \U$13893 ( \22664 , \22296 );
and \U$13894 ( \22665 , \22663 , \22664 );
nor \U$13895 ( \22666 , \22661 , \22665 );
nand \U$13896 ( \22667 , \22658 , \22666 );
and \U$13897 ( \22668 , \22667 , \22105 );
or \U$13898 ( \22669 , \22656 , \22668 );
and \U$13900 ( \22670 , \22669 , 1'b1 );
or \U$13902 ( \22671 , \22670 , 1'b0 );
buf \U$13903 ( \22672 , \22671 );
_DC r2541e_GF_IsGateDCbyConstraint ( \22673_nR2541e , \22672 , \21944 );
buf \U$13904 ( \22674 , \22673_nR2541e );
not \U$13905 ( \22675 , \22308 );
and \U$13906 ( \22676 , RIdafa508_3739, \22675 );
not \U$13907 ( \22677 , RIdafa508_3739);
or \U$13908 ( \22678 , \22677 , \22242 );
not \U$13909 ( \22679 , \22116 );
buf \U$13910 ( \22680 , RIb885d60_43);
buf \U$13911 ( \22681 , \22680 );
and \U$13912 ( \22682 , \22679 , \22681 );
buf \U$13913 ( \22683 , RIb82db60_211);
buf \U$13914 ( \22684 , \22683 );
not \U$13915 ( \22685 , \22502 );
and \U$13916 ( \22686 , \22684 , \22685 );
nor \U$13917 ( \22687 , \22682 , \22686 );
nand \U$13918 ( \22688 , \22678 , \22687 );
and \U$13919 ( \22689 , \22688 , \22308 );
or \U$13920 ( \22690 , \22676 , \22689 );
and \U$13922 ( \22691 , \22690 , 1'b1 );
or \U$13924 ( \22692 , \22691 , 1'b0 );
buf \U$13925 ( \22693 , \22692 );
_DC r25420_GF_IsGateDCbyConstraint ( \22694_nR25420 , \22693 , \21944 );
buf \U$13926 ( \22695 , \22694_nR25420 );
not \U$13927 ( \22696 , \22196 );
and \U$13928 ( \22697 , RIdafe630_3740, \22696 );
not \U$13929 ( \22698 , RIdafe630_3740);
or \U$13930 ( \22699 , \22698 , \22242 );
buf \U$13931 ( \22700 , RIb885dd8_42);
buf \U$13932 ( \22701 , \22700 );
and \U$13933 ( \22702 , \22244 , \22701 );
buf \U$13934 ( \22703 , RIb82dbd8_210);
buf \U$13935 ( \22704 , \22703 );
not \U$13936 ( \22705 , \22422 );
and \U$13937 ( \22706 , \22704 , \22705 );
nor \U$13938 ( \22707 , \22702 , \22706 );
nand \U$13939 ( \22708 , \22699 , \22707 );
and \U$13940 ( \22709 , \22708 , \22196 );
or \U$13941 ( \22710 , \22697 , \22709 );
and \U$13943 ( \22711 , \22710 , 1'b1 );
or \U$13945 ( \22712 , \22711 , 1'b0 );
buf \U$13946 ( \22713 , \22712 );
_DC r25422_GF_IsGateDCbyConstraint ( \22714_nR25422 , \22713 , \21944 );
buf \U$13947 ( \22715 , \22714_nR25422 );
buf \U$13948 ( \22716 , \22195 );
not \U$13949 ( \22717 , \22716 );
and \U$13950 ( \22718 , RIdb03b08_3741, \22717 );
not \U$13951 ( \22719 , RIdb03b08_3741);
or \U$13952 ( \22720 , \22719 , \22242 );
buf \U$13953 ( \22721 , RIb885e50_41);
and \U$13954 ( \22722 , \22158 , \22721 );
buf \U$13955 ( \22723 , RIb82dc50_209);
buf \U$13956 ( \22724 , \22723 );
not \U$13957 ( \22725 , \22339 );
and \U$13958 ( \22726 , \22724 , \22725 );
nor \U$13959 ( \22727 , \22722 , \22726 );
nand \U$13960 ( \22728 , \22720 , \22727 );
and \U$13961 ( \22729 , \22728 , \22716 );
or \U$13962 ( \22730 , \22718 , \22729 );
and \U$13964 ( \22731 , \22730 , 1'b1 );
or \U$13966 ( \22732 , \22731 , 1'b0 );
buf \U$13967 ( \22733 , \22732 );
_DC r25424_GF_IsGateDCbyConstraint ( \22734_nR25424 , \22733 , \21944 );
buf \U$13968 ( \22735 , \22734_nR25424 );
not \U$13969 ( \22736 , \22308 );
and \U$13970 ( \22737 , RIdb09d00_3742, \22736 );
not \U$13971 ( \22738 , RIdb09d00_3742);
or \U$13972 ( \22739 , \22738 , \22242 );
buf \U$13973 ( \22740 , RIb885ec8_40);
buf \U$13974 ( \22741 , \22740 );
and \U$13975 ( \22742 , \22158 , \22741 );
buf \U$13976 ( \22743 , RIb82dcc8_208);
buf \U$13977 ( \22744 , \22743 );
not \U$13978 ( \22745 , \22154 );
and \U$13979 ( \22746 , \22744 , \22745 );
nor \U$13980 ( \22747 , \22742 , \22746 );
nand \U$13981 ( \22748 , \22739 , \22747 );
and \U$13982 ( \22749 , \22748 , \22308 );
or \U$13983 ( \22750 , \22737 , \22749 );
and \U$13985 ( \22751 , \22750 , 1'b1 );
or \U$13987 ( \22752 , \22751 , 1'b0 );
buf \U$13988 ( \22753 , \22752 );
_DC r25426_GF_IsGateDCbyConstraint ( \22754_nR25426 , \22753 , \21944 );
buf \U$13989 ( \22755 , \22754_nR25426 );
buf \U$13990 ( \22756 , \22103 );
buf \U$13991 ( \22757 , \22756 );
not \U$13992 ( \22758 , \22757 );
and \U$13993 ( \22759 , RIdb0e440_3743, \22758 );
not \U$13994 ( \22760 , RIdb0e440_3743);
or \U$13995 ( \22761 , \22760 , \22354 );
buf \U$13996 ( \22762 , RIb885f40_39);
buf \U$13997 ( \22763 , \22762 );
and \U$13998 ( \22764 , \22201 , \22763 );
buf \U$13999 ( \22765 , RIb82dd40_207);
buf \U$14000 ( \22766 , \22765 );
not \U$14001 ( \22767 , \22163 );
and \U$14002 ( \22768 , \22766 , \22767 );
nor \U$14003 ( \22769 , \22764 , \22768 );
nand \U$14004 ( \22770 , \22761 , \22769 );
and \U$14005 ( \22771 , \22770 , \22757 );
or \U$14006 ( \22772 , \22759 , \22771 );
and \U$14008 ( \22773 , \22772 , 1'b1 );
or \U$14010 ( \22774 , \22773 , 1'b0 );
buf \U$14011 ( \22775 , \22774 );
_DC r2542a_GF_IsGateDCbyConstraint ( \22776_nR2542a , \22775 , \21944 );
buf \U$14012 ( \22777 , \22776_nR2542a );
not \U$14013 ( \22778 , \22757 );
and \U$14014 ( \22779 , RIdb13468_3744, \22778 );
not \U$14015 ( \22780 , RIdb13468_3744);
or \U$14016 ( \22781 , \22780 , \22128 );
buf \U$14017 ( \22782 , RIb885fb8_38);
buf \U$14018 ( \22783 , \22782 );
and \U$14019 ( \22784 , \22201 , \22783 );
buf \U$14020 ( \22785 , RIb82ddb8_206);
buf \U$14021 ( \22786 , \22785 );
not \U$14022 ( \22787 , \22502 );
and \U$14023 ( \22788 , \22786 , \22787 );
nor \U$14024 ( \22789 , \22784 , \22788 );
nand \U$14025 ( \22790 , \22781 , \22789 );
and \U$14026 ( \22791 , \22790 , \22757 );
or \U$14027 ( \22792 , \22779 , \22791 );
and \U$14029 ( \22793 , \22792 , 1'b1 );
or \U$14031 ( \22794 , \22793 , 1'b0 );
buf \U$14032 ( \22795 , \22794 );
_DC r2542c_GF_IsGateDCbyConstraint ( \22796_nR2542c , \22795 , \21944 );
buf \U$14033 ( \22797 , \22796_nR2542c );
not \U$14034 ( \22798 , \22308 );
and \U$14035 ( \22799 , RId9d7370_3745, \22798 );
not \U$14036 ( \22800 , RId9d7370_3745);
or \U$14037 ( \22801 , \22800 , \22354 );
buf \U$14038 ( \22802 , RIb886030_37);
buf \U$14039 ( \22803 , \22802 );
and \U$14040 ( \22804 , \22158 , \22803 );
buf \U$14041 ( \22805 , RIb82de30_205);
buf \U$14042 ( \22806 , \22805 );
not \U$14043 ( \22807 , \22318 );
and \U$14044 ( \22808 , \22806 , \22807 );
nor \U$14045 ( \22809 , \22804 , \22808 );
nand \U$14046 ( \22810 , \22801 , \22809 );
and \U$14047 ( \22811 , \22810 , \22308 );
or \U$14048 ( \22812 , \22799 , \22811 );
and \U$14050 ( \22813 , \22812 , 1'b1 );
or \U$14052 ( \22814 , \22813 , 1'b0 );
buf \U$14053 ( \22815 , \22814 );
_DC r2542e_GF_IsGateDCbyConstraint ( \22816_nR2542e , \22815 , \21944 );
buf \U$14054 ( \22817 , \22816_nR2542e );
not \U$14055 ( \22818 , \22716 );
and \U$14056 ( \22819 , RId9d25a0_3746, \22818 );
not \U$14057 ( \22820 , RId9d25a0_3746);
or \U$14058 ( \22821 , \22820 , \22221 );
buf \U$14059 ( \22822 , RIb8860a8_36);
buf \U$14060 ( \22823 , \22822 );
and \U$14061 ( \22824 , \22201 , \22823 );
buf \U$14062 ( \22825 , RIb832228_204);
buf \U$14063 ( \22826 , \22825 );
not \U$14064 ( \22827 , \22422 );
and \U$14065 ( \22828 , \22826 , \22827 );
nor \U$14066 ( \22829 , \22824 , \22828 );
nand \U$14067 ( \22830 , \22821 , \22829 );
and \U$14068 ( \22831 , \22830 , \22716 );
or \U$14069 ( \22832 , \22819 , \22831 );
and \U$14071 ( \22833 , \22832 , 1'b1 );
or \U$14073 ( \22834 , \22833 , 1'b0 );
buf \U$14074 ( \22835 , \22834 );
_DC r25430_GF_IsGateDCbyConstraint ( \22836_nR25430 , \22835 , \21944 );
buf \U$14075 ( \22837 , \22836_nR25430 );
not \U$14076 ( \22838 , \22757 );
and \U$14077 ( \22839 , RId9cd0c8_3747, \22838 );
not \U$14078 ( \22840 , RId9cd0c8_3747);
or \U$14079 ( \22841 , \22840 , \22395 );
buf \U$14080 ( \22842 , RIb886120_35);
buf \U$14081 ( \22843 , \22842 );
and \U$14082 ( \22844 , \22158 , \22843 );
buf \U$14083 ( \22845 , RIb8322a0_203);
buf \U$14084 ( \22846 , \22845 );
not \U$14085 ( \22847 , \22254 );
and \U$14086 ( \22848 , \22846 , \22847 );
nor \U$14087 ( \22849 , \22844 , \22848 );
nand \U$14088 ( \22850 , \22841 , \22849 );
and \U$14089 ( \22851 , \22850 , \22757 );
or \U$14090 ( \22852 , \22839 , \22851 );
and \U$14092 ( \22853 , \22852 , 1'b1 );
or \U$14094 ( \22854 , \22853 , 1'b0 );
buf \U$14095 ( \22855 , \22854 );
_DC r25432_GF_IsGateDCbyConstraint ( \22856_nR25432 , \22855 , \21944 );
buf \U$14096 ( \22857 , \22856_nR25432 );
not \U$14097 ( \22858 , \22308 );
and \U$14098 ( \22859 , RId9c86b8_3748, \22858 );
not \U$14099 ( \22860 , RId9c86b8_3748);
or \U$14100 ( \22861 , \22860 , \22269 );
buf \U$14101 ( \22862 , RIb886198_34);
buf \U$14102 ( \22863 , \22862 );
and \U$14103 ( \22864 , \22201 , \22863 );
buf \U$14104 ( \22865 , RIb832318_202);
buf \U$14105 ( \22866 , \22865 );
not \U$14106 ( \22867 , \22254 );
and \U$14107 ( \22868 , \22866 , \22867 );
nor \U$14108 ( \22869 , \22864 , \22868 );
nand \U$14109 ( \22870 , \22861 , \22869 );
and \U$14110 ( \22871 , \22870 , \22308 );
or \U$14111 ( \22872 , \22859 , \22871 );
and \U$14113 ( \22873 , \22872 , 1'b1 );
or \U$14115 ( \22874 , \22873 , 1'b0 );
buf \U$14116 ( \22875 , \22874 );
_DC r25434_GF_IsGateDCbyConstraint ( \22876_nR25434 , \22875 , \21944 );
buf \U$14117 ( \22877 , \22876_nR25434 );
not \U$14118 ( \22878 , \22757 );
and \U$14119 ( \22879 , RIda940a0_3749, \22878 );
not \U$14120 ( \22880 , RIda940a0_3749);
or \U$14121 ( \22881 , \22880 , \22156 );
buf \U$14122 ( \22882 , RIb886210_33);
buf \U$14123 ( \22883 , \22882 );
and \U$14124 ( \22884 , \22201 , \22883 );
buf \U$14125 ( \22885 , RIb832390_201);
buf \U$14126 ( \22886 , \22885 );
not \U$14127 ( \22887 , \22296 );
and \U$14128 ( \22888 , \22886 , \22887 );
nor \U$14129 ( \22889 , \22884 , \22888 );
nand \U$14130 ( \22890 , \22881 , \22889 );
and \U$14131 ( \22891 , \22890 , \22757 );
or \U$14132 ( \22892 , \22879 , \22891 );
and \U$14134 ( \22893 , \22892 , 1'b1 );
or \U$14136 ( \22894 , \22893 , 1'b0 );
buf \U$14137 ( \22895 , \22894 );
_DC r25436_GF_IsGateDCbyConstraint ( \22896_nR25436 , \22895 , \21944 );
buf \U$14138 ( \22897 , \22896_nR25436 );
not \U$14139 ( \22898 , \22757 );
and \U$14140 ( \22899 , RIda91850_3750, \22898 );
not \U$14141 ( \22900 , RIda91850_3750);
or \U$14142 ( \22901 , \22900 , \22221 );
not \U$14143 ( \22902 , \22201 );
not \U$14144 ( \22903 , \22902 );
buf \U$14145 ( \22904 , RIb886288_32);
buf \U$14146 ( \22905 , \22904 );
and \U$14147 ( \22906 , \22903 , \22905 );
buf \U$14148 ( \22907 , RIb832408_200);
buf \U$14149 ( \22908 , \22907 );
not \U$14150 ( \22909 , \22318 );
and \U$14151 ( \22910 , \22908 , \22909 );
nor \U$14152 ( \22911 , \22906 , \22910 );
nand \U$14153 ( \22912 , \22901 , \22911 );
and \U$14154 ( \22913 , \22912 , \22757 );
or \U$14155 ( \22914 , \22899 , \22913 );
and \U$14157 ( \22915 , \22914 , 1'b1 );
or \U$14159 ( \22916 , \22915 , 1'b0 );
buf \U$14160 ( \22917 , \22916 );
_DC r25438_GF_IsGateDCbyConstraint ( \22918_nR25438 , \22917 , \21944 );
buf \U$14161 ( \22919 , \22918_nR25438 );
not \U$14162 ( \22920 , \22308 );
and \U$14163 ( \22921 , RIda8dbd8_3751, \22920 );
not \U$14164 ( \22922 , RIda8dbd8_3751);
or \U$14165 ( \22923 , \22922 , \22395 );
buf \U$14166 ( \22924 , RIb886300_31);
buf \U$14167 ( \22925 , \22924 );
and \U$14168 ( \22926 , \22201 , \22925 );
buf \U$14169 ( \22927 , RIb832480_199);
buf \U$14170 ( \22928 , \22927 );
not \U$14171 ( \22929 , \22422 );
and \U$14172 ( \22930 , \22928 , \22929 );
nor \U$14173 ( \22931 , \22926 , \22930 );
nand \U$14174 ( \22932 , \22923 , \22931 );
and \U$14175 ( \22933 , \22932 , \22308 );
or \U$14176 ( \22934 , \22921 , \22933 );
and \U$14178 ( \22935 , \22934 , 1'b1 );
or \U$14180 ( \22936 , \22935 , 1'b0 );
buf \U$14181 ( \22937 , \22936 );
_DC r2543a_GF_IsGateDCbyConstraint ( \22938_nR2543a , \22937 , \21944 );
buf \U$14182 ( \22939 , \22938_nR2543a );
not \U$14183 ( \22940 , \22716 );
and \U$14184 ( \22941 , RIda8a7d0_3752, \22940 );
not \U$14185 ( \22942 , RIda8a7d0_3752);
or \U$14186 ( \22943 , \22942 , \22269 );
buf \U$14187 ( \22944 , RIb886378_30);
buf \U$14188 ( \22945 , \22944 );
and \U$14189 ( \22946 , \22201 , \22945 );
buf \U$14190 ( \22947 , RIb8324f8_198);
buf \U$14191 ( \22948 , \22947 );
not \U$14192 ( \22949 , \22339 );
and \U$14193 ( \22950 , \22948 , \22949 );
nor \U$14194 ( \22951 , \22946 , \22950 );
nand \U$14195 ( \22952 , \22943 , \22951 );
and \U$14196 ( \22953 , \22952 , \22716 );
or \U$14197 ( \22954 , \22941 , \22953 );
and \U$14199 ( \22955 , \22954 , 1'b1 );
or \U$14201 ( \22956 , \22955 , 1'b0 );
buf \U$14202 ( \22957 , \22956 );
_DC r2543c_GF_IsGateDCbyConstraint ( \22958_nR2543c , \22957 , \21944 );
buf \U$14203 ( \22959 , \22958_nR2543c );
not \U$14204 ( \22960 , \22716 );
and \U$14205 ( \22961 , RIda86978_3753, \22960 );
not \U$14206 ( \22962 , RIda86978_3753);
or \U$14207 ( \22963 , \22962 , \22156 );
buf \U$14208 ( \22964 , RIb8863f0_29);
buf \U$14209 ( \22965 , \22964 );
and \U$14210 ( \22966 , \22130 , \22965 );
buf \U$14211 ( \22967 , RIb832570_197);
buf \U$14212 ( \22968 , \22967 );
not \U$14213 ( \22969 , \22339 );
and \U$14214 ( \22970 , \22968 , \22969 );
nor \U$14215 ( \22971 , \22966 , \22970 );
nand \U$14216 ( \22972 , \22963 , \22971 );
and \U$14217 ( \22973 , \22972 , \22716 );
or \U$14218 ( \22974 , \22961 , \22973 );
and \U$14220 ( \22975 , \22974 , 1'b1 );
or \U$14222 ( \22976 , \22975 , 1'b0 );
buf \U$14223 ( \22977 , \22976 );
_DC r25440_GF_IsGateDCbyConstraint ( \22978_nR25440 , \22977 , \21944 );
buf \U$14224 ( \22979 , \22978_nR25440 );
not \U$14225 ( \22980 , \22308 );
and \U$14226 ( \22981 , RIda835e8_3754, \22980 );
not \U$14227 ( \22982 , RIda835e8_3754);
or \U$14228 ( \22983 , \22982 , \22156 );
buf \U$14229 ( \22984 , RIb886468_28);
and \U$14230 ( \22985 , \22244 , \22984 );
buf \U$14231 ( \22986 , RIb8383a8_196);
buf \U$14232 ( \22987 , \22986 );
not \U$14233 ( \22988 , \22154 );
and \U$14234 ( \22989 , \22987 , \22988 );
nor \U$14235 ( \22990 , \22985 , \22989 );
nand \U$14236 ( \22991 , \22983 , \22990 );
and \U$14237 ( \22992 , \22991 , \22308 );
or \U$14238 ( \22993 , \22981 , \22992 );
and \U$14240 ( \22994 , \22993 , 1'b1 );
or \U$14242 ( \22995 , \22994 , 1'b0 );
buf \U$14243 ( \22996 , \22995 );
_DC r25442_GF_IsGateDCbyConstraint ( \22997_nR25442 , \22996 , \21944 );
buf \U$14244 ( \22998 , \22997_nR25442 );
not \U$14245 ( \22999 , \22716 );
and \U$14246 ( \23000 , RIda80f00_3755, \22999 );
not \U$14247 ( \23001 , RIda80f00_3755);
or \U$14248 ( \23002 , \23001 , \22242 );
buf \U$14249 ( \23003 , RIb8864e0_27);
and \U$14250 ( \23004 , \22244 , \23003 );
buf \U$14251 ( \23005 , RIb838420_195);
buf \U$14252 ( \23006 , \23005 );
not \U$14253 ( \23007 , \22296 );
and \U$14254 ( \23008 , \23006 , \23007 );
nor \U$14255 ( \23009 , \23004 , \23008 );
nand \U$14256 ( \23010 , \23002 , \23009 );
and \U$14257 ( \23011 , \23010 , \22716 );
or \U$14258 ( \23012 , \23000 , \23011 );
and \U$14260 ( \23013 , \23012 , 1'b1 );
or \U$14262 ( \23014 , \23013 , 1'b0 );
buf \U$14263 ( \23015 , \23014 );
_DC r25444_GF_IsGateDCbyConstraint ( \23016_nR25444 , \23015 , \21944 );
buf \U$14264 ( \23017 , \23016_nR25444 );
not \U$14265 ( \23018 , \22757 );
and \U$14266 ( \23019 , RIda7daf8_3756, \23018 );
not \U$14267 ( \23020 , RIda7daf8_3756);
or \U$14268 ( \23021 , \23020 , \22242 );
buf \U$14269 ( \23022 , RIb886558_26);
buf \U$14270 ( \23023 , \23022 );
and \U$14271 ( \23024 , \22158 , \23023 );
buf \U$14272 ( \23025 , RIb838498_194);
buf \U$14273 ( \23026 , \23025 );
not \U$14274 ( \23027 , \22126 );
and \U$14275 ( \23028 , \23026 , \23027 );
nor \U$14276 ( \23029 , \23024 , \23028 );
nand \U$14277 ( \23030 , \23021 , \23029 );
and \U$14278 ( \23031 , \23030 , \22757 );
or \U$14279 ( \23032 , \23019 , \23031 );
and \U$14281 ( \23033 , \23032 , 1'b1 );
or \U$14283 ( \23034 , \23033 , 1'b0 );
buf \U$14284 ( \23035 , \23034 );
_DC r25446_GF_IsGateDCbyConstraint ( \23036_nR25446 , \23035 , \21944 );
buf \U$14285 ( \23037 , \23036_nR25446 );
buf \U$14286 ( \23038 , \22103 );
buf \U$14287 ( \23039 , \23038 );
not \U$14288 ( \23040 , \23039 );
and \U$14289 ( \23041 , RIda7a7e0_3757, \23040 );
not \U$14290 ( \23042 , RIda7a7e0_3757);
or \U$14291 ( \23043 , \23042 , \22128 );
buf \U$14292 ( \23044 , RIb8865d0_25);
buf \U$14293 ( \23045 , \23044 );
and \U$14294 ( \23046 , \22201 , \23045 );
buf \U$14295 ( \23047 , RIb838510_193);
buf \U$14296 ( \23048 , \23047 );
not \U$14297 ( \23049 , \22163 );
and \U$14298 ( \23050 , \23048 , \23049 );
nor \U$14299 ( \23051 , \23046 , \23050 );
nand \U$14300 ( \23052 , \23043 , \23051 );
and \U$14301 ( \23053 , \23052 , \23039 );
or \U$14302 ( \23054 , \23041 , \23053 );
and \U$14304 ( \23055 , \23054 , 1'b1 );
or \U$14306 ( \23056 , \23055 , 1'b0 );
buf \U$14307 ( \23057 , \23056 );
_DC r25448_GF_IsGateDCbyConstraint ( \23058_nR25448 , \23057 , \21944 );
buf \U$14308 ( \23059 , \23058_nR25448 );
not \U$14309 ( \23060 , \22716 );
and \U$14310 ( \23061 , RIda745e8_3758, \23060 );
not \U$14311 ( \23062 , RIda745e8_3758);
or \U$14312 ( \23063 , \23062 , \22354 );
buf \U$14313 ( \23064 , RIb886648_24);
buf \U$14314 ( \23065 , \23064 );
and \U$14315 ( \23066 , \22130 , \23065 );
buf \U$14316 ( \23067 , RIb838588_192);
buf \U$14317 ( \23068 , \23067 );
not \U$14318 ( \23069 , \22502 );
and \U$14319 ( \23070 , \23068 , \23069 );
nor \U$14320 ( \23071 , \23066 , \23070 );
nand \U$14321 ( \23072 , \23063 , \23071 );
and \U$14322 ( \23073 , \23072 , \22716 );
or \U$14323 ( \23074 , \23061 , \23073 );
and \U$14325 ( \23075 , \23074 , 1'b1 );
or \U$14327 ( \23076 , \23075 , 1'b0 );
buf \U$14328 ( \23077 , \23076 );
_DC r2544a_GF_IsGateDCbyConstraint ( \23078_nR2544a , \23077 , \21944 );
buf \U$14329 ( \23079 , \23078_nR2544a );
not \U$14330 ( \23080 , \22757 );
and \U$14331 ( \23081 , RIda6e018_3759, \23080 );
not \U$14332 ( \23082 , RIda6e018_3759);
or \U$14333 ( \23083 , \23082 , \22156 );
buf \U$14334 ( \23084 , RIb8866c0_23);
buf \U$14335 ( \23085 , \23084 );
and \U$14336 ( \23086 , \22244 , \23085 );
buf \U$14337 ( \23087 , RIb838600_191);
buf \U$14338 ( \23088 , \23087 );
not \U$14339 ( \23089 , \22254 );
and \U$14340 ( \23090 , \23088 , \23089 );
nor \U$14341 ( \23091 , \23086 , \23090 );
nand \U$14342 ( \23092 , \23083 , \23091 );
and \U$14343 ( \23093 , \23092 , \22757 );
or \U$14344 ( \23094 , \23081 , \23093 );
and \U$14346 ( \23095 , \23094 , 1'b1 );
or \U$14348 ( \23096 , \23095 , 1'b0 );
buf \U$14349 ( \23097 , \23096 );
_DC r2544c_GF_IsGateDCbyConstraint ( \23098_nR2544c , \23097 , \21944 );
buf \U$14350 ( \23099 , \23098_nR2544c );
not \U$14351 ( \23100 , \23039 );
and \U$14352 ( \23101 , RIda65e40_3760, \23100 );
not \U$14353 ( \23102 , RIda65e40_3760);
or \U$14354 ( \23103 , \23102 , \22156 );
buf \U$14355 ( \23104 , RIb886738_22);
buf \U$14356 ( \23105 , \23104 );
and \U$14357 ( \23106 , \22158 , \23105 );
buf \U$14358 ( \23107 , RIb838678_190);
buf \U$14359 ( \23108 , \23107 );
not \U$14360 ( \23109 , \22296 );
and \U$14361 ( \23110 , \23108 , \23109 );
nor \U$14362 ( \23111 , \23106 , \23110 );
nand \U$14363 ( \23112 , \23103 , \23111 );
and \U$14364 ( \23113 , \23112 , \23039 );
or \U$14365 ( \23114 , \23101 , \23113 );
and \U$14367 ( \23115 , \23114 , 1'b1 );
or \U$14369 ( \23116 , \23115 , 1'b0 );
buf \U$14370 ( \23117 , \23116 );
_DC r2544e_GF_IsGateDCbyConstraint ( \23118_nR2544e , \23117 , \21944 );
buf \U$14371 ( \23119 , \23118_nR2544e );
not \U$14372 ( \23120 , \22757 );
and \U$14373 ( \23121 , RIda5f888_3761, \23120 );
not \U$14374 ( \23122 , RIda5f888_3761);
or \U$14375 ( \23123 , \23122 , \22242 );
buf \U$14376 ( \23124 , RIb8867b0_21);
buf \U$14377 ( \23125 , \23124 );
and \U$14378 ( \23126 , \22244 , \23125 );
buf \U$14379 ( \23127 , RIb8386f0_189);
buf \U$14380 ( \23128 , \23127 );
not \U$14381 ( \23129 , \22318 );
and \U$14382 ( \23130 , \23128 , \23129 );
nor \U$14383 ( \23131 , \23126 , \23130 );
nand \U$14384 ( \23132 , \23123 , \23131 );
and \U$14385 ( \23133 , \23132 , \22757 );
or \U$14386 ( \23134 , \23121 , \23133 );
and \U$14388 ( \23135 , \23134 , 1'b1 );
or \U$14390 ( \23136 , \23135 , 1'b0 );
buf \U$14391 ( \23137 , \23136 );
_DC r25450_GF_IsGateDCbyConstraint ( \23138_nR25450 , \23137 , \21944 );
buf \U$14392 ( \23139 , \23138_nR25450 );
not \U$14393 ( \23140 , \22757 );
and \U$14394 ( \23141 , RIda59780_3762, \23140 );
not \U$14395 ( \23142 , RIda59780_3762);
or \U$14396 ( \23143 , \23142 , \22156 );
buf \U$14397 ( \23144 , RIb886828_20);
buf \U$14398 ( \23145 , \23144 );
and \U$14399 ( \23146 , \22201 , \23145 );
buf \U$14400 ( \23147 , RIb838768_188);
buf \U$14401 ( \23148 , \23147 );
not \U$14402 ( \23149 , \22126 );
and \U$14403 ( \23150 , \23148 , \23149 );
nor \U$14404 ( \23151 , \23146 , \23150 );
nand \U$14405 ( \23152 , \23143 , \23151 );
and \U$14406 ( \23153 , \23152 , \22757 );
or \U$14407 ( \23154 , \23141 , \23153 );
and \U$14409 ( \23155 , \23154 , 1'b1 );
or \U$14411 ( \23156 , \23155 , 1'b0 );
buf \U$14412 ( \23157 , \23156 );
_DC r25452_GF_IsGateDCbyConstraint ( \23158_nR25452 , \23157 , \21944 );
buf \U$14413 ( \23159 , \23158_nR25452 );
not \U$14414 ( \23160 , \23039 );
and \U$14415 ( \23161 , RIda510f8_3763, \23160 );
not \U$14416 ( \23162 , RIda510f8_3763);
or \U$14417 ( \23163 , \23162 , \22395 );
buf \U$14418 ( \23164 , RIb8868a0_19);
buf \U$14419 ( \23165 , \23164 );
and \U$14420 ( \23166 , \22244 , \23165 );
buf \U$14421 ( \23167 , RIb8387e0_187);
buf \U$14422 ( \23168 , \23167 );
not \U$14423 ( \23169 , \22318 );
and \U$14424 ( \23170 , \23168 , \23169 );
nor \U$14425 ( \23171 , \23166 , \23170 );
nand \U$14426 ( \23172 , \23163 , \23171 );
and \U$14427 ( \23173 , \23172 , \23039 );
or \U$14428 ( \23174 , \23161 , \23173 );
and \U$14430 ( \23175 , \23174 , 1'b1 );
or \U$14432 ( \23176 , \23175 , 1'b0 );
buf \U$14433 ( \23177 , \23176 );
_DC r25456_GF_IsGateDCbyConstraint ( \23178_nR25456 , \23177 , \21944 );
buf \U$14434 ( \23179 , \23178_nR25456 );
not \U$14435 ( \23180 , \22716 );
and \U$14436 ( \23181 , RIda4aff0_3764, \23180 );
not \U$14437 ( \23182 , RIda4aff0_3764);
or \U$14438 ( \23183 , \23182 , \22269 );
buf \U$14439 ( \23184 , RIb886918_18);
and \U$14440 ( \23185 , \22244 , \23184 );
buf \U$14441 ( \23186 , RIb838858_186);
buf \U$14442 ( \23187 , \23186 );
not \U$14443 ( \23188 , \22422 );
and \U$14444 ( \23189 , \23187 , \23188 );
nor \U$14445 ( \23190 , \23185 , \23189 );
nand \U$14446 ( \23191 , \23183 , \23190 );
and \U$14447 ( \23192 , \23191 , \22716 );
or \U$14448 ( \23193 , \23181 , \23192 );
and \U$14450 ( \23194 , \23193 , 1'b1 );
or \U$14452 ( \23195 , \23194 , 1'b0 );
buf \U$14453 ( \23196 , \23195 );
_DC r25458_GF_IsGateDCbyConstraint ( \23197_nR25458 , \23196 , \21944 );
buf \U$14454 ( \23198 , \23197_nR25458 );
not \U$14455 ( \23199 , \22716 );
and \U$14456 ( \23200 , RId927408_3765, \23199 );
not \U$14457 ( \23201 , RId927408_3765);
or \U$14458 ( \23202 , \23201 , \22156 );
buf \U$14459 ( \23203 , RIb886990_17);
buf \U$14460 ( \23204 , \23203 );
and \U$14461 ( \23205 , \22201 , \23204 );
buf \U$14462 ( \23206 , RIb8388d0_185);
buf \U$14463 ( \23207 , \23206 );
not \U$14464 ( \23208 , \22339 );
and \U$14465 ( \23209 , \23207 , \23208 );
nor \U$14466 ( \23210 , \23205 , \23209 );
nand \U$14467 ( \23211 , \23202 , \23210 );
and \U$14468 ( \23212 , \23211 , \22716 );
or \U$14469 ( \23213 , \23200 , \23212 );
and \U$14471 ( \23214 , \23213 , 1'b1 );
or \U$14473 ( \23215 , \23214 , 1'b0 );
buf \U$14474 ( \23216 , \23215 );
_DC r2545a_GF_IsGateDCbyConstraint ( \23217_nR2545a , \23216 , \21944 );
buf \U$14475 ( \23218 , \23217_nR2545a );
not \U$14476 ( \23219 , \23039 );
and \U$14477 ( \23220 , RId943680_3766, \23219 );
not \U$14478 ( \23221 , RId943680_3766);
or \U$14479 ( \23222 , \23221 , \22156 );
buf \U$14480 ( \23223 , RIb886a08_16);
buf \U$14481 ( \23224 , \23223 );
and \U$14482 ( \23225 , \22130 , \23224 );
buf \U$14483 ( \23226 , RIb838948_184);
buf \U$14484 ( \23227 , \23226 );
not \U$14485 ( \23228 , \22154 );
and \U$14486 ( \23229 , \23227 , \23228 );
nor \U$14487 ( \23230 , \23225 , \23229 );
nand \U$14488 ( \23231 , \23222 , \23230 );
and \U$14489 ( \23232 , \23231 , \23039 );
or \U$14490 ( \23233 , \23220 , \23232 );
and \U$14492 ( \23234 , \23233 , 1'b1 );
or \U$14494 ( \23235 , \23234 , 1'b0 );
buf \U$14495 ( \23236 , \23235 );
_DC r2545c_GF_IsGateDCbyConstraint ( \23237_nR2545c , \23236 , \21944 );
buf \U$14496 ( \23238 , \23237_nR2545c );
not \U$14497 ( \23239 , \22757 );
and \U$14498 ( \23240 , RId96ccd8_3767, \23239 );
not \U$14499 ( \23241 , RId96ccd8_3767);
or \U$14500 ( \23242 , \23241 , \22156 );
buf \U$14501 ( \23243 , RIb886a80_15);
buf \U$14502 ( \23244 , \23243 );
and \U$14503 ( \23245 , \22244 , \23244 );
buf \U$14504 ( \23246 , RIb8389c0_183);
buf \U$14505 ( \23247 , \23246 );
not \U$14506 ( \23248 , \22126 );
and \U$14507 ( \23249 , \23247 , \23248 );
nor \U$14508 ( \23250 , \23245 , \23249 );
nand \U$14509 ( \23251 , \23242 , \23250 );
and \U$14510 ( \23252 , \23251 , \22757 );
or \U$14511 ( \23253 , \23240 , \23252 );
and \U$14513 ( \23254 , \23253 , 1'b1 );
or \U$14515 ( \23255 , \23254 , 1'b0 );
buf \U$14516 ( \23256 , \23255 );
_DC r2545e_GF_IsGateDCbyConstraint ( \23257_nR2545e , \23256 , \21944 );
buf \U$14517 ( \23258 , \23257_nR2545e );
not \U$14518 ( \23259 , \22757 );
and \U$14519 ( \23260 , RId988b30_3768, \23259 );
not \U$14520 ( \23261 , RId988b30_3768);
or \U$14521 ( \23262 , \23261 , \22128 );
buf \U$14522 ( \23263 , RIb886af8_14);
buf \U$14523 ( \23264 , \23263 );
and \U$14524 ( \23265 , \22201 , \23264 );
buf \U$14525 ( \23266 , RIb838a38_182);
buf \U$14526 ( \23267 , \23266 );
not \U$14527 ( \23268 , \22163 );
and \U$14528 ( \23269 , \23267 , \23268 );
nor \U$14529 ( \23270 , \23265 , \23269 );
nand \U$14530 ( \23271 , \23262 , \23270 );
and \U$14531 ( \23272 , \23271 , \22757 );
or \U$14532 ( \23273 , \23260 , \23272 );
and \U$14534 ( \23274 , \23273 , 1'b1 );
or \U$14536 ( \23275 , \23274 , 1'b0 );
buf \U$14537 ( \23276 , \23275 );
_DC r25460_GF_IsGateDCbyConstraint ( \23277_nR25460 , \23276 , \21944 );
buf \U$14538 ( \23278 , \23277_nR25460 );
not \U$14539 ( \23279 , \23039 );
and \U$14540 ( \23280 , RId90bb68_3769, \23279 );
not \U$14541 ( \23281 , RId90bb68_3769);
or \U$14542 ( \23282 , \23281 , \22354 );
buf \U$14543 ( \23283 , RIb886b70_13);
buf \U$14544 ( \23284 , \23283 );
and \U$14545 ( \23285 , \22130 , \23284 );
buf \U$14546 ( \23286 , RIb838ab0_181);
buf \U$14547 ( \23287 , \23286 );
not \U$14548 ( \23288 , \22502 );
and \U$14549 ( \23289 , \23287 , \23288 );
nor \U$14550 ( \23290 , \23285 , \23289 );
nand \U$14551 ( \23291 , \23282 , \23290 );
and \U$14552 ( \23292 , \23291 , \23039 );
or \U$14553 ( \23293 , \23280 , \23292 );
and \U$14555 ( \23294 , \23293 , 1'b1 );
or \U$14557 ( \23295 , \23294 , 1'b0 );
buf \U$14558 ( \23296 , \23295 );
_DC r25462_GF_IsGateDCbyConstraint ( \23297_nR25462 , \23296 , \21944 );
buf \U$14559 ( \23298 , \23297_nR25462 );
not \U$14560 ( \23299 , \22716 );
and \U$14561 ( \23300 , RId8f7438_3770, \23299 );
not \U$14562 ( \23301 , RId8f7438_3770);
or \U$14563 ( \23302 , \23301 , \22221 );
buf \U$14564 ( \23303 , RIb886be8_12);
and \U$14565 ( \23304 , \22244 , \23303 );
buf \U$14566 ( \23305 , RIb838b28_180);
buf \U$14567 ( \23306 , \23305 );
not \U$14568 ( \23307 , \22502 );
and \U$14569 ( \23308 , \23306 , \23307 );
nor \U$14570 ( \23309 , \23304 , \23308 );
nand \U$14571 ( \23310 , \23302 , \23309 );
and \U$14572 ( \23311 , \23310 , \22716 );
or \U$14573 ( \23312 , \23300 , \23311 );
and \U$14575 ( \23313 , \23312 , 1'b1 );
or \U$14577 ( \23314 , \23313 , 1'b0 );
buf \U$14578 ( \23315 , \23314 );
_DC r25464_GF_IsGateDCbyConstraint ( \23316_nR25464 , \23315 , \21944 );
buf \U$14579 ( \23317 , \23316_nR25464 );
not \U$14580 ( \23318 , \22757 );
and \U$14581 ( \23319 , RId8d6dc8_3771, \23318 );
not \U$14582 ( \23320 , RId8d6dc8_3771);
or \U$14583 ( \23321 , \23320 , \22395 );
buf \U$14584 ( \23322 , RIb886c60_11);
buf \U$14585 ( \23323 , \23322 );
and \U$14586 ( \23324 , \22158 , \23323 );
buf \U$14587 ( \23325 , RIb838ba0_179);
buf \U$14588 ( \23326 , \23325 );
not \U$14589 ( \23327 , \22254 );
and \U$14590 ( \23328 , \23326 , \23327 );
nor \U$14591 ( \23329 , \23324 , \23328 );
nand \U$14592 ( \23330 , \23321 , \23329 );
and \U$14593 ( \23331 , \23330 , \22757 );
or \U$14594 ( \23332 , \23319 , \23331 );
and \U$14596 ( \23333 , \23332 , 1'b1 );
or \U$14598 ( \23334 , \23333 , 1'b0 );
buf \U$14599 ( \23335 , \23334 );
_DC r25466_GF_IsGateDCbyConstraint ( \23336_nR25466 , \23335 , \21944 );
buf \U$14600 ( \23337 , \23336_nR25466 );
not \U$14601 ( \23338 , \23039 );
and \U$14602 ( \23339 , RId6c4d70_3772, \23338 );
not \U$14603 ( \23340 , RId6c4d70_3772);
or \U$14604 ( \23341 , \23340 , \22242 );
buf \U$14605 ( \23342 , RIb886cd8_10);
buf \U$14606 ( \23343 , \23342 );
and \U$14607 ( \23344 , \22130 , \23343 );
buf \U$14608 ( \23345 , RIb838c18_178);
buf \U$14609 ( \23346 , \23345 );
not \U$14610 ( \23347 , \22422 );
and \U$14611 ( \23348 , \23346 , \23347 );
nor \U$14612 ( \23349 , \23344 , \23348 );
nand \U$14613 ( \23350 , \23341 , \23349 );
and \U$14614 ( \23351 , \23350 , \23039 );
or \U$14615 ( \23352 , \23339 , \23351 );
and \U$14617 ( \23353 , \23352 , 1'b1 );
or \U$14619 ( \23354 , \23353 , 1'b0 );
buf \U$14620 ( \23355 , \23354 );
_DC r25468_GF_IsGateDCbyConstraint ( \23356_nR25468 , \23355 , \21944 );
buf \U$14621 ( \23357 , \23356_nR25468 );
buf \U$14622 ( \23358 , \22756 );
not \U$14623 ( \23359 , \23358 );
and \U$14624 ( \23360 , RId6ae7c8_3773, \23359 );
not \U$14625 ( \23361 , RId6ae7c8_3773);
or \U$14626 ( \23362 , \23361 , \22128 );
buf \U$14627 ( \23363 , RIb886d50_9);
buf \U$14628 ( \23364 , \23363 );
and \U$14629 ( \23365 , \22244 , \23364 );
buf \U$14630 ( \23366 , RIb838c90_177);
buf \U$14631 ( \23367 , \23366 );
not \U$14632 ( \23368 , \22296 );
and \U$14633 ( \23369 , \23367 , \23368 );
nor \U$14634 ( \23370 , \23365 , \23369 );
nand \U$14635 ( \23371 , \23362 , \23370 );
and \U$14636 ( \23372 , \23371 , \23358 );
or \U$14637 ( \23373 , \23360 , \23372 );
and \U$14639 ( \23374 , \23373 , 1'b1 );
or \U$14641 ( \23375 , \23374 , 1'b0 );
buf \U$14642 ( \23376 , \23375 );
_DC r2546c_GF_IsGateDCbyConstraint ( \23377_nR2546c , \23376 , \21944 );
buf \U$14643 ( \23378 , \23377_nR2546c );
not \U$14644 ( \23379 , \23358 );
and \U$14645 ( \23380 , RId835578_3774, \23379 );
not \U$14646 ( \23381 , RId835578_3774);
or \U$14647 ( \23382 , \23381 , \22354 );
buf \U$14648 ( \23383 , RIb886dc8_8);
buf \U$14649 ( \23384 , \23383 );
and \U$14650 ( \23385 , \22130 , \23384 );
buf \U$14651 ( \23386 , RIb838d08_176);
buf \U$14652 ( \23387 , \23386 );
not \U$14653 ( \23388 , \22318 );
and \U$14654 ( \23389 , \23387 , \23388 );
nor \U$14655 ( \23390 , \23385 , \23389 );
nand \U$14656 ( \23391 , \23382 , \23390 );
and \U$14657 ( \23392 , \23391 , \23358 );
or \U$14658 ( \23393 , \23380 , \23392 );
and \U$14660 ( \23394 , \23393 , 1'b1 );
or \U$14662 ( \23395 , \23394 , 1'b0 );
buf \U$14663 ( \23396 , \23395 );
_DC r2546e_GF_IsGateDCbyConstraint ( \23397_nR2546e , \23396 , \21944 );
buf \U$14664 ( \23398 , \23397_nR2546e );
not \U$14665 ( \23399 , \23039 );
and \U$14666 ( \23400 , RId8a9d50_3775, \23399 );
not \U$14667 ( \23401 , RId8a9d50_3775);
or \U$14668 ( \23402 , \23401 , \22221 );
buf \U$14669 ( \23403 , RIb886e40_7);
buf \U$14670 ( \23404 , \23403 );
and \U$14671 ( \23405 , \22244 , \23404 );
buf \U$14672 ( \23406 , RIb838d80_175);
buf \U$14673 ( \23407 , \23406 );
not \U$14674 ( \23408 , \22422 );
and \U$14675 ( \23409 , \23407 , \23408 );
nor \U$14676 ( \23410 , \23405 , \23409 );
nand \U$14677 ( \23411 , \23402 , \23410 );
and \U$14678 ( \23412 , \23411 , \23039 );
or \U$14679 ( \23413 , \23400 , \23412 );
and \U$14681 ( \23414 , \23413 , 1'b1 );
or \U$14683 ( \23415 , \23414 , 1'b0 );
buf \U$14684 ( \23416 , \23415 );
_DC r25470_GF_IsGateDCbyConstraint ( \23417_nR25470 , \23416 , \21944 );
buf \U$14685 ( \23418 , \23417_nR25470 );
not \U$14686 ( \23419 , \22716 );
and \U$14687 ( \23420 , RId862aa0_3776, \23419 );
not \U$14688 ( \23421 , RId862aa0_3776);
or \U$14689 ( \23422 , \23421 , \22395 );
buf \U$14690 ( \23423 , RIb886eb8_6);
buf \U$14691 ( \23424 , \23423 );
and \U$14692 ( \23425 , \22130 , \23424 );
buf \U$14693 ( \23426 , RIb838df8_174);
buf \U$14694 ( \23427 , \23426 );
not \U$14695 ( \23428 , \22339 );
and \U$14696 ( \23429 , \23427 , \23428 );
nor \U$14697 ( \23430 , \23425 , \23429 );
nand \U$14698 ( \23431 , \23422 , \23430 );
and \U$14699 ( \23432 , \23431 , \22716 );
or \U$14700 ( \23433 , \23420 , \23432 );
and \U$14702 ( \23434 , \23433 , 1'b1 );
or \U$14704 ( \23435 , \23434 , 1'b0 );
buf \U$14705 ( \23436 , \23435 );
_DC r25472_GF_IsGateDCbyConstraint ( \23437_nR25472 , \23436 , \21944 );
buf \U$14706 ( \23438 , \23437_nR25472 );
not \U$14707 ( \23439 , \22716 );
and \U$14708 ( \23440 , RId99e778_3777, \23439 );
not \U$14709 ( \23441 , RId99e778_3777);
not \U$14710 ( \23442 , \22121 );
nor \U$14711 ( \23443 , \22117 , \23442 );
nand \U$14712 ( \23444 , \23443 , \22123 );
not \U$14713 ( \23445 , \23444 );
not \U$14714 ( \23446 , \22110 );
or \U$14715 ( \23447 , \22111 , \23446 );
not \U$14716 ( \23448 , \23447 );
nand \U$14717 ( \23449 , \22102 , \23448 );
not \U$14718 ( \23450 , \23449 );
or \U$14719 ( \23451 , \23445 , \23450 );
not \U$14720 ( \23452 , \23451 );
not \U$14721 ( \23453 , \23452 );
or \U$14722 ( \23454 , \23441 , \23453 );
not \U$14723 ( \23455 , \23444 );
not \U$14724 ( \23456 , \23455 );
not \U$14725 ( \23457 , \23456 );
and \U$14726 ( \23458 , \22135 , \23457 );
not \U$14727 ( \23459 , \23458 );
not \U$14728 ( \23460 , \22132 );
not \U$14729 ( \23461 , \23449 );
buf \U$14730 ( \23462 , \23461 );
not \U$14731 ( \23463 , \23462 );
or \U$14732 ( \23464 , \23460 , \23463 );
nand \U$14733 ( \23465 , \23454 , \23459 , \23464 );
and \U$14734 ( \23466 , \23465 , \22716 );
or \U$14735 ( \23467 , \23440 , \23466 );
and \U$14737 ( \23468 , \23467 , 1'b1 );
or \U$14739 ( \23469 , \23468 , 1'b0 );
buf \U$14740 ( \23470 , \23469 );
_DC r2547c_GF_IsGateDCbyConstraint ( \23471_nR2547c , \23470 , \21944 );
buf \U$14741 ( \23472 , \23471_nR2547c );
not \U$14742 ( \23473 , \23039 );
and \U$14743 ( \23474 , RId9ac620_3778, \23473 );
not \U$14744 ( \23475 , RId9ac620_3778);
not \U$14745 ( \23476 , \23452 );
or \U$14746 ( \23477 , \23475 , \23476 );
not \U$14747 ( \23478 , \23455 );
not \U$14748 ( \23479 , \23478 );
and \U$14749 ( \23480 , \22162 , \23479 );
not \U$14750 ( \23481 , \23480 );
not \U$14751 ( \23482 , \22159 );
not \U$14752 ( \23483 , \23461 );
or \U$14753 ( \23484 , \23482 , \23483 );
nand \U$14754 ( \23485 , \23477 , \23481 , \23484 );
and \U$14755 ( \23486 , \23485 , \23039 );
or \U$14756 ( \23487 , \23474 , \23486 );
and \U$14758 ( \23488 , \23487 , 1'b1 );
or \U$14760 ( \23489 , \23488 , 1'b0 );
buf \U$14761 ( \23490 , \23489 );
_DC r25492_GF_IsGateDCbyConstraint ( \23491_nR25492 , \23490 , \21944 );
buf \U$14762 ( \23492 , \23491_nR25492 );
not \U$14763 ( \23493 , \22716 );
and \U$14764 ( \23494 , RId9b8290_3779, \23493 );
not \U$14765 ( \23495 , RId9b8290_3779);
or \U$14766 ( \23496 , \23495 , \23476 );
not \U$14767 ( \23497 , \23456 );
and \U$14768 ( \23498 , \22183 , \23497 );
not \U$14769 ( \23499 , \23498 );
not \U$14770 ( \23500 , \22180 );
not \U$14771 ( \23501 , \23462 );
or \U$14772 ( \23502 , \23500 , \23501 );
nand \U$14773 ( \23503 , \23496 , \23499 , \23502 );
and \U$14774 ( \23504 , \23503 , \22716 );
or \U$14775 ( \23505 , \23494 , \23504 );
and \U$14777 ( \23506 , \23505 , 1'b1 );
or \U$14779 ( \23507 , \23506 , 1'b0 );
buf \U$14780 ( \23508 , \23507 );
_DC r254a8_GF_IsGateDCbyConstraint ( \23509_nR254a8 , \23508 , \21944 );
buf \U$14781 ( \23510 , \23509_nR254a8 );
not \U$14782 ( \23511 , \23358 );
and \U$14783 ( \23512 , RId9bdfd8_3780, \23511 );
not \U$14784 ( \23513 , RId9bdfd8_3780);
or \U$14785 ( \23514 , \23513 , \23476 );
not \U$14786 ( \23515 , \23478 );
and \U$14787 ( \23516 , \22206 , \23515 );
not \U$14788 ( \23517 , \23516 );
not \U$14789 ( \23518 , \22203 );
not \U$14790 ( \23519 , \23461 );
or \U$14791 ( \23520 , \23518 , \23519 );
nand \U$14792 ( \23521 , \23514 , \23517 , \23520 );
and \U$14793 ( \23522 , \23521 , \23358 );
or \U$14794 ( \23523 , \23512 , \23522 );
and \U$14796 ( \23524 , \23523 , 1'b1 );
or \U$14798 ( \23525 , \23524 , 1'b0 );
buf \U$14799 ( \23526 , \23525 );
_DC r254be_GF_IsGateDCbyConstraint ( \23527_nR254be , \23526 , \21944 );
buf \U$14800 ( \23528 , \23527_nR254be );
not \U$14801 ( \23529 , \23039 );
and \U$14802 ( \23530 , RId90fe70_3781, \23529 );
not \U$14803 ( \23531 , RId90fe70_3781);
not \U$14804 ( \23532 , \23452 );
or \U$14805 ( \23533 , \23531 , \23532 );
not \U$14806 ( \23534 , \23456 );
and \U$14807 ( \23535 , \22227 , \23534 );
not \U$14808 ( \23536 , \23535 );
not \U$14809 ( \23537 , \22224 );
buf \U$14810 ( \23538 , \23461 );
not \U$14811 ( \23539 , \23538 );
or \U$14812 ( \23540 , \23537 , \23539 );
nand \U$14813 ( \23541 , \23533 , \23536 , \23540 );
and \U$14814 ( \23542 , \23541 , \23039 );
or \U$14815 ( \23543 , \23530 , \23542 );
and \U$14817 ( \23544 , \23543 , 1'b1 );
or \U$14819 ( \23545 , \23544 , 1'b0 );
buf \U$14820 ( \23546 , \23545 );
_DC r254d4_GF_IsGateDCbyConstraint ( \23547_nR254d4 , \23546 , \21944 );
buf \U$14821 ( \23548 , \23547_nR254d4 );
buf \U$14822 ( \23549 , \22756 );
not \U$14823 ( \23550 , \23549 );
and \U$14824 ( \23551 , RId918b10_3782, \23550 );
not \U$14825 ( \23552 , RId918b10_3782);
not \U$14826 ( \23553 , \23452 );
or \U$14827 ( \23554 , \23552 , \23553 );
not \U$14828 ( \23555 , \23455 );
not \U$14829 ( \23556 , \23555 );
and \U$14830 ( \23557 , \22249 , \23556 );
not \U$14831 ( \23558 , \23557 );
not \U$14832 ( \23559 , \22246 );
not \U$14833 ( \23560 , \23462 );
or \U$14834 ( \23561 , \23559 , \23560 );
nand \U$14835 ( \23562 , \23554 , \23558 , \23561 );
and \U$14836 ( \23563 , \23562 , \23549 );
or \U$14837 ( \23564 , \23551 , \23563 );
and \U$14839 ( \23565 , \23564 , 1'b1 );
or \U$14841 ( \23566 , \23565 , 1'b0 );
buf \U$14842 ( \23567 , \23566 );
_DC r254ea_GF_IsGateDCbyConstraint ( \23568_nR254ea , \23567 , \21944 );
buf \U$14843 ( \23569 , \23568_nR254ea );
not \U$14844 ( \23570 , \23549 );
and \U$14845 ( \23571 , RIda42698_3783, \23570 );
not \U$14846 ( \23572 , RIda42698_3783);
or \U$14847 ( \23573 , \23572 , \23476 );
not \U$14848 ( \23574 , \23444 );
and \U$14849 ( \23575 , \22275 , \23574 );
not \U$14850 ( \23576 , \23575 );
not \U$14851 ( \23577 , \22272 );
not \U$14852 ( \23578 , \23538 );
or \U$14853 ( \23579 , \23577 , \23578 );
nand \U$14854 ( \23580 , \23573 , \23576 , \23579 );
and \U$14855 ( \23581 , \23580 , \23549 );
or \U$14856 ( \23582 , \23571 , \23581 );
and \U$14858 ( \23583 , \23582 , 1'b1 );
or \U$14860 ( \23584 , \23583 , 1'b0 );
buf \U$14861 ( \23585 , \23584 );
_DC r254f4_GF_IsGateDCbyConstraint ( \23586_nR254f4 , \23585 , \21944 );
buf \U$14862 ( \23587 , \23586_nR254f4 );
not \U$14863 ( \23588 , \23039 );
and \U$14864 ( \23589 , RIda33a58_3784, \23588 );
not \U$14865 ( \23590 , RIda33a58_3784);
or \U$14866 ( \23591 , \23590 , \23476 );
not \U$14867 ( \23592 , \23478 );
and \U$14868 ( \23593 , \22295 , \23592 );
not \U$14869 ( \23594 , \23593 );
not \U$14870 ( \23595 , \22292 );
buf \U$14871 ( \23596 , \23461 );
not \U$14872 ( \23597 , \23596 );
or \U$14873 ( \23598 , \23595 , \23597 );
nand \U$14874 ( \23599 , \23591 , \23594 , \23598 );
and \U$14875 ( \23600 , \23599 , \23039 );
or \U$14876 ( \23601 , \23589 , \23600 );
and \U$14878 ( \23602 , \23601 , 1'b1 );
or \U$14880 ( \23603 , \23602 , 1'b0 );
buf \U$14881 ( \23604 , \23603 );
_DC r254f6_GF_IsGateDCbyConstraint ( \23605_nR254f6 , \23604 , \21944 );
buf \U$14882 ( \23606 , \23605_nR254f6 );
not \U$14883 ( \23607 , \23358 );
and \U$14884 ( \23608 , RIda28b08_3785, \23607 );
not \U$14885 ( \23609 , RIda28b08_3785);
or \U$14886 ( \23610 , \23609 , \23453 );
not \U$14887 ( \23611 , \23555 );
and \U$14888 ( \23612 , \22317 , \23611 );
not \U$14889 ( \23613 , \23612 );
not \U$14890 ( \23614 , \22314 );
not \U$14891 ( \23615 , \23538 );
or \U$14892 ( \23616 , \23614 , \23615 );
nand \U$14893 ( \23617 , \23610 , \23613 , \23616 );
and \U$14894 ( \23618 , \23617 , \23358 );
or \U$14895 ( \23619 , \23608 , \23618 );
and \U$14897 ( \23620 , \23619 , 1'b1 );
or \U$14899 ( \23621 , \23620 , 1'b0 );
buf \U$14900 ( \23622 , \23621 );
_DC r254f8_GF_IsGateDCbyConstraint ( \23623_nR254f8 , \23622 , \21944 );
buf \U$14901 ( \23624 , \23623_nR254f8 );
not \U$14902 ( \23625 , \23358 );
and \U$14903 ( \23626 , RIda18aa0_3786, \23625 );
not \U$14904 ( \23627 , RIda18aa0_3786);
not \U$14905 ( \23628 , \23452 );
or \U$14906 ( \23629 , \23627 , \23628 );
not \U$14907 ( \23630 , \23455 );
not \U$14908 ( \23631 , \23630 );
and \U$14909 ( \23632 , \22338 , \23631 );
not \U$14910 ( \23633 , \23632 );
not \U$14911 ( \23634 , \22335 );
not \U$14912 ( \23635 , \23538 );
or \U$14913 ( \23636 , \23634 , \23635 );
nand \U$14914 ( \23637 , \23629 , \23633 , \23636 );
and \U$14915 ( \23638 , \23637 , \23358 );
or \U$14916 ( \23639 , \23626 , \23638 );
and \U$14918 ( \23640 , \23639 , 1'b1 );
or \U$14920 ( \23641 , \23640 , 1'b0 );
buf \U$14921 ( \23642 , \23641 );
_DC r254fa_GF_IsGateDCbyConstraint ( \23643_nR254fa , \23642 , \21944 );
buf \U$14922 ( \23644 , \23643_nR254fa );
not \U$14923 ( \23645 , \23039 );
and \U$14924 ( \23646 , RIda0b288_3787, \23645 );
not \U$14925 ( \23647 , RIda0b288_3787);
or \U$14926 ( \23648 , \23647 , \23532 );
not \U$14927 ( \23649 , \23455 );
not \U$14928 ( \23650 , \23649 );
and \U$14929 ( \23651 , \22360 , \23650 );
not \U$14930 ( \23652 , \23651 );
not \U$14931 ( \23653 , \22357 );
not \U$14932 ( \23654 , \23462 );
or \U$14933 ( \23655 , \23653 , \23654 );
nand \U$14934 ( \23656 , \23648 , \23652 , \23655 );
and \U$14935 ( \23657 , \23656 , \23039 );
or \U$14936 ( \23658 , \23646 , \23657 );
and \U$14938 ( \23659 , \23658 , 1'b1 );
or \U$14940 ( \23660 , \23659 , 1'b0 );
buf \U$14941 ( \23661 , \23660 );
_DC r2547e_GF_IsGateDCbyConstraint ( \23662_nR2547e , \23661 , \21944 );
buf \U$14942 ( \23663 , \23662_nR2547e );
not \U$14943 ( \23664 , \23549 );
and \U$14944 ( \23665 , RId9f8d18_3788, \23664 );
not \U$14945 ( \23666 , RId9f8d18_3788);
or \U$14946 ( \23667 , \23666 , \23553 );
not \U$14947 ( \23668 , \23649 );
and \U$14948 ( \23669 , \22380 , \23668 );
not \U$14949 ( \23670 , \23669 );
not \U$14950 ( \23671 , \22377 );
not \U$14951 ( \23672 , \23462 );
or \U$14952 ( \23673 , \23671 , \23672 );
nand \U$14953 ( \23674 , \23667 , \23670 , \23673 );
and \U$14954 ( \23675 , \23674 , \23549 );
or \U$14955 ( \23676 , \23665 , \23675 );
and \U$14957 ( \23677 , \23676 , 1'b1 );
or \U$14959 ( \23678 , \23677 , 1'b0 );
buf \U$14960 ( \23679 , \23678 );
_DC r25480_GF_IsGateDCbyConstraint ( \23680_nR25480 , \23679 , \21944 );
buf \U$14961 ( \23681 , \23680_nR25480 );
not \U$14962 ( \23682 , \23549 );
and \U$14963 ( \23683 , RId9ec9a0_3789, \23682 );
not \U$14964 ( \23684 , RId9ec9a0_3789);
or \U$14965 ( \23685 , \23684 , \23476 );
not \U$14966 ( \23686 , \23455 );
not \U$14967 ( \23687 , \23686 );
and \U$14968 ( \23688 , \22401 , \23687 );
not \U$14969 ( \23689 , \23688 );
not \U$14970 ( \23690 , \22398 );
not \U$14971 ( \23691 , \23461 );
or \U$14972 ( \23692 , \23690 , \23691 );
nand \U$14973 ( \23693 , \23685 , \23689 , \23692 );
and \U$14974 ( \23694 , \23693 , \23549 );
or \U$14975 ( \23695 , \23683 , \23694 );
and \U$14977 ( \23696 , \23695 , 1'b1 );
or \U$14979 ( \23697 , \23696 , 1'b0 );
buf \U$14980 ( \23698 , \23697 );
_DC r25482_GF_IsGateDCbyConstraint ( \23699_nR25482 , \23698 , \21944 );
buf \U$14981 ( \23700 , \23699_nR25482 );
not \U$14982 ( \23701 , \23039 );
and \U$14983 ( \23702 , RId9e3418_3790, \23701 );
not \U$14984 ( \23703 , RId9e3418_3790);
or \U$14985 ( \23704 , \23703 , \23628 );
not \U$14986 ( \23705 , \23456 );
and \U$14987 ( \23706 , \22421 , \23705 );
not \U$14988 ( \23707 , \23706 );
not \U$14989 ( \23708 , \22418 );
not \U$14990 ( \23709 , \23462 );
or \U$14991 ( \23710 , \23708 , \23709 );
nand \U$14992 ( \23711 , \23704 , \23707 , \23710 );
and \U$14993 ( \23712 , \23711 , \23039 );
or \U$14994 ( \23713 , \23702 , \23712 );
and \U$14996 ( \23714 , \23713 , 1'b1 );
or \U$14998 ( \23715 , \23714 , 1'b0 );
buf \U$14999 ( \23716 , \23715 );
_DC r25484_GF_IsGateDCbyConstraint ( \23717_nR25484 , \23716 , \21944 );
buf \U$15000 ( \23718 , \23717_nR25484 );
not \U$15001 ( \23719 , \23549 );
and \U$15002 ( \23720 , RIdb156a0_3791, \23719 );
not \U$15003 ( \23721 , RIdb156a0_3791);
or \U$15004 ( \23722 , \23721 , \23628 );
not \U$15005 ( \23723 , \23630 );
and \U$15006 ( \23724 , \22441 , \23723 );
not \U$15007 ( \23725 , \23724 );
not \U$15008 ( \23726 , \22438 );
not \U$15009 ( \23727 , \23461 );
or \U$15010 ( \23728 , \23726 , \23727 );
nand \U$15011 ( \23729 , \23722 , \23725 , \23728 );
and \U$15012 ( \23730 , \23729 , \23549 );
or \U$15013 ( \23731 , \23720 , \23730 );
and \U$15015 ( \23732 , \23731 , 1'b1 );
or \U$15017 ( \23733 , \23732 , 1'b0 );
buf \U$15018 ( \23734 , \23733 );
_DC r25486_GF_IsGateDCbyConstraint ( \23735_nR25486 , \23734 , \21944 );
buf \U$15019 ( \23736 , \23735_nR25486 );
not \U$15020 ( \23737 , \23358 );
and \U$15021 ( \23738 , RIdb17f68_3792, \23737 );
not \U$15022 ( \23739 , RIdb17f68_3792);
or \U$15023 ( \23740 , \23739 , \23628 );
not \U$15024 ( \23741 , \23649 );
and \U$15025 ( \23742 , \22461 , \23741 );
not \U$15026 ( \23743 , \23742 );
not \U$15027 ( \23744 , \22458 );
not \U$15028 ( \23745 , \23596 );
or \U$15029 ( \23746 , \23744 , \23745 );
nand \U$15030 ( \23747 , \23740 , \23743 , \23746 );
and \U$15031 ( \23748 , \23747 , \23358 );
or \U$15032 ( \23749 , \23738 , \23748 );
and \U$15034 ( \23750 , \23749 , 1'b1 );
or \U$15036 ( \23751 , \23750 , 1'b0 );
buf \U$15037 ( \23752 , \23751 );
_DC r25488_GF_IsGateDCbyConstraint ( \23753_nR25488 , \23752 , \21944 );
buf \U$15038 ( \23754 , \23753_nR25488 );
buf \U$15039 ( \23755 , \23038 );
not \U$15040 ( \23756 , \23755 );
and \U$15041 ( \23757 , RIdb1b640_3793, \23756 );
not \U$15042 ( \23758 , RIdb1b640_3793);
or \U$15043 ( \23759 , \23758 , \23453 );
not \U$15044 ( \23760 , \23555 );
and \U$15045 ( \23761 , \22481 , \23760 );
not \U$15046 ( \23762 , \23761 );
not \U$15047 ( \23763 , \22478 );
not \U$15048 ( \23764 , \23538 );
or \U$15049 ( \23765 , \23763 , \23764 );
nand \U$15050 ( \23766 , \23759 , \23762 , \23765 );
and \U$15051 ( \23767 , \23766 , \23755 );
or \U$15052 ( \23768 , \23757 , \23767 );
and \U$15054 ( \23769 , \23768 , 1'b1 );
or \U$15056 ( \23770 , \23769 , 1'b0 );
buf \U$15057 ( \23771 , \23770 );
_DC r2548a_GF_IsGateDCbyConstraint ( \23772_nR2548a , \23771 , \21944 );
buf \U$15058 ( \23773 , \23772_nR2548a );
not \U$15059 ( \23774 , \23549 );
and \U$15060 ( \23775 , RIdb1df08_3794, \23774 );
not \U$15061 ( \23776 , RIdb1df08_3794);
or \U$15062 ( \23777 , \23776 , \23476 );
not \U$15063 ( \23778 , \23444 );
and \U$15064 ( \23779 , \22501 , \23778 );
not \U$15065 ( \23780 , \23779 );
not \U$15066 ( \23781 , \22498 );
not \U$15067 ( \23782 , \23596 );
or \U$15068 ( \23783 , \23781 , \23782 );
nand \U$15069 ( \23784 , \23777 , \23780 , \23783 );
and \U$15070 ( \23785 , \23784 , \23549 );
or \U$15071 ( \23786 , \23775 , \23785 );
and \U$15073 ( \23787 , \23786 , 1'b1 );
or \U$15075 ( \23788 , \23787 , 1'b0 );
buf \U$15076 ( \23789 , \23788 );
_DC r2548c_GF_IsGateDCbyConstraint ( \23790_nR2548c , \23789 , \21944 );
buf \U$15077 ( \23791 , \23790_nR2548c );
not \U$15078 ( \23792 , \23358 );
and \U$15079 ( \23793 , RIdb215e0_3795, \23792 );
not \U$15080 ( \23794 , RIdb215e0_3795);
or \U$15081 ( \23795 , \23794 , \23453 );
not \U$15082 ( \23796 , \23686 );
and \U$15083 ( \23797 , \22522 , \23796 );
not \U$15084 ( \23798 , \23797 );
not \U$15085 ( \23799 , \22519 );
not \U$15086 ( \23800 , \23596 );
or \U$15087 ( \23801 , \23799 , \23800 );
nand \U$15088 ( \23802 , \23795 , \23798 , \23801 );
and \U$15089 ( \23803 , \23802 , \23358 );
or \U$15090 ( \23804 , \23793 , \23803 );
and \U$15092 ( \23805 , \23804 , 1'b1 );
or \U$15094 ( \23806 , \23805 , 1'b0 );
buf \U$15095 ( \23807 , \23806 );
_DC r2548e_GF_IsGateDCbyConstraint ( \23808_nR2548e , \23807 , \21944 );
buf \U$15096 ( \23809 , \23808_nR2548e );
not \U$15097 ( \23810 , \23755 );
and \U$15098 ( \23811 , RIdb23ea8_3796, \23810 );
not \U$15099 ( \23812 , RIdb23ea8_3796);
or \U$15100 ( \23813 , \23812 , \23553 );
not \U$15101 ( \23814 , \23444 );
and \U$15102 ( \23815 , \22542 , \23814 );
not \U$15103 ( \23816 , \23815 );
not \U$15104 ( \23817 , \22539 );
not \U$15105 ( \23818 , \23462 );
or \U$15106 ( \23819 , \23817 , \23818 );
nand \U$15107 ( \23820 , \23813 , \23816 , \23819 );
and \U$15108 ( \23821 , \23820 , \23755 );
or \U$15109 ( \23822 , \23811 , \23821 );
and \U$15111 ( \23823 , \23822 , 1'b1 );
or \U$15113 ( \23824 , \23823 , 1'b0 );
buf \U$15114 ( \23825 , \23824 );
_DC r25490_GF_IsGateDCbyConstraint ( \23826_nR25490 , \23825 , \21944 );
buf \U$15115 ( \23827 , \23826_nR25490 );
not \U$15116 ( \23828 , \23358 );
and \U$15117 ( \23829 , RIdb26c20_3797, \23828 );
not \U$15118 ( \23830 , RIdb26c20_3797);
or \U$15119 ( \23831 , \23830 , \23628 );
not \U$15120 ( \23832 , \23555 );
and \U$15121 ( \23833 , \22562 , \23832 );
not \U$15122 ( \23834 , \23833 );
not \U$15123 ( \23835 , \22559 );
not \U$15124 ( \23836 , \23596 );
or \U$15125 ( \23837 , \23835 , \23836 );
nand \U$15126 ( \23838 , \23831 , \23834 , \23837 );
and \U$15127 ( \23839 , \23838 , \23358 );
or \U$15128 ( \23840 , \23829 , \23839 );
and \U$15130 ( \23841 , \23840 , 1'b1 );
or \U$15132 ( \23842 , \23841 , 1'b0 );
buf \U$15133 ( \23843 , \23842 );
_DC r25494_GF_IsGateDCbyConstraint ( \23844_nR25494 , \23843 , \21944 );
buf \U$15134 ( \23845 , \23844_nR25494 );
not \U$15135 ( \23846 , \23358 );
and \U$15136 ( \23847 , RIdb29e48_3798, \23846 );
not \U$15137 ( \23848 , RIdb29e48_3798);
or \U$15138 ( \23849 , \23848 , \23553 );
not \U$15139 ( \23850 , \23630 );
and \U$15140 ( \23851 , \22582 , \23850 );
not \U$15141 ( \23852 , \23851 );
not \U$15142 ( \23853 , \22579 );
not \U$15143 ( \23854 , \23596 );
or \U$15144 ( \23855 , \23853 , \23854 );
nand \U$15145 ( \23856 , \23849 , \23852 , \23855 );
and \U$15146 ( \23857 , \23856 , \23358 );
or \U$15147 ( \23858 , \23847 , \23857 );
and \U$15149 ( \23859 , \23858 , 1'b1 );
or \U$15151 ( \23860 , \23859 , 1'b0 );
buf \U$15152 ( \23861 , \23860 );
_DC r25496_GF_IsGateDCbyConstraint ( \23862_nR25496 , \23861 , \21944 );
buf \U$15153 ( \23863 , \23862_nR25496 );
not \U$15154 ( \23864 , \23755 );
and \U$15155 ( \23865 , RIdb2cbc0_3799, \23864 );
not \U$15156 ( \23866 , RIdb2cbc0_3799);
or \U$15157 ( \23867 , \23866 , \23532 );
not \U$15158 ( \23868 , \23478 );
and \U$15159 ( \23869 , \22602 , \23868 );
not \U$15160 ( \23870 , \23869 );
not \U$15161 ( \23871 , \22599 );
not \U$15162 ( \23872 , \23462 );
or \U$15163 ( \23873 , \23871 , \23872 );
nand \U$15164 ( \23874 , \23867 , \23870 , \23873 );
and \U$15165 ( \23875 , \23874 , \23755 );
or \U$15166 ( \23876 , \23865 , \23875 );
and \U$15168 ( \23877 , \23876 , 1'b1 );
or \U$15170 ( \23878 , \23877 , 1'b0 );
buf \U$15171 ( \23879 , \23878 );
_DC r25498_GF_IsGateDCbyConstraint ( \23880_nR25498 , \23879 , \21944 );
buf \U$15172 ( \23881 , \23880_nR25498 );
not \U$15173 ( \23882 , \23549 );
and \U$15174 ( \23883 , RIdb2fde8_3800, \23882 );
not \U$15175 ( \23884 , RIdb2fde8_3800);
or \U$15176 ( \23885 , \23884 , \23532 );
not \U$15177 ( \23886 , \23555 );
and \U$15178 ( \23887 , \22622 , \23886 );
not \U$15179 ( \23888 , \23887 );
not \U$15180 ( \23889 , \22619 );
not \U$15181 ( \23890 , \23596 );
or \U$15182 ( \23891 , \23889 , \23890 );
nand \U$15183 ( \23892 , \23885 , \23888 , \23891 );
and \U$15184 ( \23893 , \23892 , \23549 );
or \U$15185 ( \23894 , \23883 , \23893 );
and \U$15187 ( \23895 , \23894 , 1'b1 );
or \U$15189 ( \23896 , \23895 , 1'b0 );
buf \U$15190 ( \23897 , \23896 );
_DC r2549a_GF_IsGateDCbyConstraint ( \23898_nR2549a , \23897 , \21944 );
buf \U$15191 ( \23899 , \23898_nR2549a );
not \U$15192 ( \23900 , \23549 );
and \U$15193 ( \23901 , RIdb32b60_3801, \23900 );
not \U$15194 ( \23902 , RIdb32b60_3801);
or \U$15195 ( \23903 , \23902 , \23453 );
not \U$15196 ( \23904 , \23630 );
and \U$15197 ( \23905 , \22643 , \23904 );
not \U$15198 ( \23906 , \23905 );
not \U$15199 ( \23907 , \22640 );
not \U$15200 ( \23908 , \23596 );
or \U$15201 ( \23909 , \23907 , \23908 );
nand \U$15202 ( \23910 , \23903 , \23906 , \23909 );
and \U$15203 ( \23911 , \23910 , \23549 );
or \U$15204 ( \23912 , \23901 , \23911 );
and \U$15206 ( \23913 , \23912 , 1'b1 );
or \U$15208 ( \23914 , \23913 , 1'b0 );
buf \U$15209 ( \23915 , \23914 );
_DC r2549c_GF_IsGateDCbyConstraint ( \23916_nR2549c , \23915 , \21944 );
buf \U$15210 ( \23917 , \23916_nR2549c );
not \U$15211 ( \23918 , \23755 );
and \U$15212 ( \23919 , RIdb35d88_3802, \23918 );
not \U$15213 ( \23920 , RIdb35d88_3802);
or \U$15214 ( \23921 , \23920 , \23532 );
not \U$15215 ( \23922 , \23686 );
and \U$15216 ( \23923 , \22663 , \23922 );
not \U$15217 ( \23924 , \23923 );
not \U$15218 ( \23925 , \22660 );
not \U$15219 ( \23926 , \23596 );
or \U$15220 ( \23927 , \23925 , \23926 );
nand \U$15221 ( \23928 , \23921 , \23924 , \23927 );
and \U$15222 ( \23929 , \23928 , \23755 );
or \U$15223 ( \23930 , \23919 , \23929 );
and \U$15225 ( \23931 , \23930 , 1'b1 );
or \U$15227 ( \23932 , \23931 , 1'b0 );
buf \U$15228 ( \23933 , \23932 );
_DC r2549e_GF_IsGateDCbyConstraint ( \23934_nR2549e , \23933 , \21944 );
buf \U$15229 ( \23935 , \23934_nR2549e );
not \U$15230 ( \23936 , \23549 );
and \U$15231 ( \23937 , RIdb38b00_3803, \23936 );
not \U$15232 ( \23938 , RIdb38b00_3803);
or \U$15233 ( \23939 , \23938 , \23453 );
not \U$15234 ( \23940 , \23455 );
not \U$15235 ( \23941 , \23940 );
and \U$15236 ( \23942 , \22684 , \23941 );
not \U$15237 ( \23943 , \23942 );
not \U$15238 ( \23944 , \22681 );
not \U$15239 ( \23945 , \23596 );
or \U$15240 ( \23946 , \23944 , \23945 );
nand \U$15241 ( \23947 , \23939 , \23943 , \23946 );
and \U$15242 ( \23948 , \23947 , \23549 );
or \U$15243 ( \23949 , \23937 , \23948 );
and \U$15245 ( \23950 , \23949 , 1'b1 );
or \U$15247 ( \23951 , \23950 , 1'b0 );
buf \U$15248 ( \23952 , \23951 );
_DC r254a0_GF_IsGateDCbyConstraint ( \23953_nR254a0 , \23952 , \21944 );
buf \U$15249 ( \23954 , \23953_nR254a0 );
not \U$15250 ( \23955 , \23358 );
and \U$15251 ( \23956 , RIdb3b3c8_3804, \23955 );
not \U$15252 ( \23957 , RIdb3b3c8_3804);
or \U$15253 ( \23958 , \23957 , \23553 );
not \U$15254 ( \23959 , \23940 );
and \U$15255 ( \23960 , \22704 , \23959 );
not \U$15256 ( \23961 , \23960 );
not \U$15257 ( \23962 , \22701 );
not \U$15258 ( \23963 , \23462 );
or \U$15259 ( \23964 , \23962 , \23963 );
nand \U$15260 ( \23965 , \23958 , \23961 , \23964 );
and \U$15261 ( \23966 , \23965 , \23358 );
or \U$15262 ( \23967 , \23956 , \23966 );
and \U$15264 ( \23968 , \23967 , 1'b1 );
or \U$15266 ( \23969 , \23968 , 1'b0 );
buf \U$15267 ( \23970 , \23969 );
_DC r254a2_GF_IsGateDCbyConstraint ( \23971_nR254a2 , \23970 , \21944 );
buf \U$15268 ( \23972 , \23971_nR254a2 );
not \U$15269 ( \23973 , \23755 );
and \U$15270 ( \23974 , RIdb3eaa0_3805, \23973 );
not \U$15271 ( \23975 , RIdb3eaa0_3805);
or \U$15272 ( \23976 , \23975 , \23628 );
not \U$15273 ( \23977 , \23686 );
and \U$15274 ( \23978 , \22724 , \23977 );
not \U$15275 ( \23979 , \23978 );
not \U$15276 ( \23980 , \22721 );
not \U$15277 ( \23981 , \23462 );
or \U$15278 ( \23982 , \23980 , \23981 );
nand \U$15279 ( \23983 , \23976 , \23979 , \23982 );
and \U$15280 ( \23984 , \23983 , \23755 );
or \U$15281 ( \23985 , \23974 , \23984 );
and \U$15283 ( \23986 , \23985 , 1'b1 );
or \U$15285 ( \23987 , \23986 , 1'b0 );
buf \U$15286 ( \23988 , \23987 );
_DC r254a4_GF_IsGateDCbyConstraint ( \23989_nR254a4 , \23988 , \21944 );
buf \U$15287 ( \23990 , \23989_nR254a4 );
not \U$15288 ( \23991 , \23549 );
and \U$15289 ( \23992 , RIdb404e0_3806, \23991 );
not \U$15290 ( \23993 , RIdb404e0_3806);
or \U$15291 ( \23994 , \23993 , \23453 );
not \U$15292 ( \23995 , \23940 );
and \U$15293 ( \23996 , \22744 , \23995 );
not \U$15294 ( \23997 , \23996 );
not \U$15295 ( \23998 , \22741 );
not \U$15296 ( \23999 , \23462 );
or \U$15297 ( \24000 , \23998 , \23999 );
nand \U$15298 ( \24001 , \23994 , \23997 , \24000 );
and \U$15299 ( \24002 , \24001 , \23549 );
or \U$15300 ( \24003 , \23992 , \24002 );
and \U$15302 ( \24004 , \24003 , 1'b1 );
or \U$15304 ( \24005 , \24004 , 1'b0 );
buf \U$15305 ( \24006 , \24005 );
_DC r254a6_GF_IsGateDCbyConstraint ( \24007_nR254a6 , \24006 , \21944 );
buf \U$15306 ( \24008 , \24007_nR254a6 );
not \U$15307 ( \24009 , \23549 );
and \U$15308 ( \24010 , RIdb422e0_3807, \24009 );
not \U$15309 ( \24011 , RIdb422e0_3807);
or \U$15310 ( \24012 , \24011 , \23628 );
not \U$15311 ( \24013 , \23555 );
and \U$15312 ( \24014 , \22766 , \24013 );
not \U$15313 ( \24015 , \24014 );
not \U$15314 ( \24016 , \22763 );
not \U$15315 ( \24017 , \23596 );
or \U$15316 ( \24018 , \24016 , \24017 );
nand \U$15317 ( \24019 , \24012 , \24015 , \24018 );
and \U$15318 ( \24020 , \24019 , \23549 );
or \U$15319 ( \24021 , \24010 , \24020 );
and \U$15321 ( \24022 , \24021 , 1'b1 );
or \U$15323 ( \24023 , \24022 , 1'b0 );
buf \U$15324 ( \24024 , \24023 );
_DC r254aa_GF_IsGateDCbyConstraint ( \24025_nR254aa , \24024 , \21944 );
buf \U$15325 ( \24026 , \24025_nR254aa );
not \U$15326 ( \24027 , \23755 );
and \U$15327 ( \24028 , RIdb43ac8_3808, \24027 );
not \U$15328 ( \24029 , RIdb43ac8_3808);
or \U$15329 ( \24030 , \24029 , \23453 );
not \U$15330 ( \24031 , \23456 );
and \U$15331 ( \24032 , \22786 , \24031 );
not \U$15332 ( \24033 , \24032 );
not \U$15333 ( \24034 , \22783 );
not \U$15334 ( \24035 , \23596 );
or \U$15335 ( \24036 , \24034 , \24035 );
nand \U$15336 ( \24037 , \24030 , \24033 , \24036 );
and \U$15337 ( \24038 , \24037 , \23755 );
or \U$15338 ( \24039 , \24028 , \24038 );
and \U$15340 ( \24040 , \24039 , 1'b1 );
or \U$15342 ( \24041 , \24040 , 1'b0 );
buf \U$15343 ( \24042 , \24041 );
_DC r254ac_GF_IsGateDCbyConstraint ( \24043_nR254ac , \24042 , \21944 );
buf \U$15344 ( \24044 , \24043_nR254ac );
not \U$15345 ( \24045 , \23358 );
and \U$15346 ( \24046 , RIdb45850_3809, \24045 );
not \U$15347 ( \24047 , RIdb45850_3809);
or \U$15348 ( \24048 , \24047 , \23532 );
not \U$15349 ( \24049 , \23649 );
and \U$15350 ( \24050 , \22806 , \24049 );
not \U$15351 ( \24051 , \24050 );
not \U$15352 ( \24052 , \22803 );
not \U$15353 ( \24053 , \23462 );
or \U$15354 ( \24054 , \24052 , \24053 );
nand \U$15355 ( \24055 , \24048 , \24051 , \24054 );
and \U$15356 ( \24056 , \24055 , \23358 );
or \U$15357 ( \24057 , \24046 , \24056 );
and \U$15359 ( \24058 , \24057 , 1'b1 );
or \U$15361 ( \24059 , \24058 , 1'b0 );
buf \U$15362 ( \24060 , \24059 );
_DC r254ae_GF_IsGateDCbyConstraint ( \24061_nR254ae , \24060 , \21944 );
buf \U$15363 ( \24062 , \24061_nR254ae );
not \U$15364 ( \24063 , \23358 );
and \U$15365 ( \24064 , RIdb47128_3810, \24063 );
not \U$15366 ( \24065 , RIdb47128_3810);
or \U$15367 ( \24066 , \24065 , \23553 );
not \U$15368 ( \24067 , \23649 );
and \U$15369 ( \24068 , \22826 , \24067 );
not \U$15370 ( \24069 , \24068 );
not \U$15371 ( \24070 , \22823 );
not \U$15372 ( \24071 , \23596 );
or \U$15373 ( \24072 , \24070 , \24071 );
nand \U$15374 ( \24073 , \24066 , \24069 , \24072 );
and \U$15375 ( \24074 , \24073 , \23358 );
or \U$15376 ( \24075 , \24064 , \24074 );
and \U$15378 ( \24076 , \24075 , 1'b1 );
or \U$15380 ( \24077 , \24076 , 1'b0 );
buf \U$15381 ( \24078 , \24077 );
_DC r254b0_GF_IsGateDCbyConstraint ( \24079_nR254b0 , \24078 , \21944 );
buf \U$15382 ( \24080 , \24079_nR254b0 );
not \U$15383 ( \24081 , \23755 );
and \U$15384 ( \24082 , RIdb483e8_3811, \24081 );
not \U$15385 ( \24083 , RIdb483e8_3811);
or \U$15386 ( \24084 , \24083 , \23553 );
not \U$15387 ( \24085 , \23940 );
and \U$15388 ( \24086 , \22846 , \24085 );
not \U$15389 ( \24087 , \24086 );
not \U$15390 ( \24088 , \22843 );
not \U$15391 ( \24089 , \23462 );
or \U$15392 ( \24090 , \24088 , \24089 );
nand \U$15393 ( \24091 , \24084 , \24087 , \24090 );
and \U$15394 ( \24092 , \24091 , \23755 );
or \U$15395 ( \24093 , \24082 , \24092 );
and \U$15397 ( \24094 , \24093 , 1'b1 );
or \U$15399 ( \24095 , \24094 , 1'b0 );
buf \U$15400 ( \24096 , \24095 );
_DC r254b2_GF_IsGateDCbyConstraint ( \24097_nR254b2 , \24096 , \21944 );
buf \U$15401 ( \24098 , \24097_nR254b2 );
not \U$15402 ( \24099 , \23549 );
and \U$15403 ( \24100 , RIdb49888_3812, \24099 );
not \U$15404 ( \24101 , RIdb49888_3812);
or \U$15405 ( \24102 , \24101 , \23476 );
not \U$15406 ( \24103 , \23444 );
and \U$15407 ( \24104 , \22866 , \24103 );
not \U$15408 ( \24105 , \24104 );
not \U$15409 ( \24106 , \22863 );
not \U$15410 ( \24107 , \23596 );
or \U$15411 ( \24108 , \24106 , \24107 );
nand \U$15412 ( \24109 , \24102 , \24105 , \24108 );
and \U$15413 ( \24110 , \24109 , \23549 );
or \U$15414 ( \24111 , \24100 , \24110 );
and \U$15416 ( \24112 , \24111 , 1'b1 );
or \U$15418 ( \24113 , \24112 , 1'b0 );
buf \U$15419 ( \24114 , \24113 );
_DC r254b4_GF_IsGateDCbyConstraint ( \24115_nR254b4 , \24114 , \21944 );
buf \U$15420 ( \24116 , \24115_nR254b4 );
buf \U$15421 ( \24117 , \22103 );
buf \U$15422 ( \24118 , \24117 );
not \U$15423 ( \24119 , \24118 );
and \U$15424 ( \24120 , RIdb4abc0_3813, \24119 );
not \U$15425 ( \24121 , RIdb4abc0_3813);
or \U$15426 ( \24122 , \24121 , \23476 );
not \U$15427 ( \24123 , \23456 );
and \U$15428 ( \24124 , \22886 , \24123 );
not \U$15429 ( \24125 , \24124 );
not \U$15430 ( \24126 , \22883 );
not \U$15431 ( \24127 , \23596 );
or \U$15432 ( \24128 , \24126 , \24127 );
nand \U$15433 ( \24129 , \24122 , \24125 , \24128 );
and \U$15434 ( \24130 , \24129 , \24118 );
or \U$15435 ( \24131 , \24120 , \24130 );
and \U$15437 ( \24132 , \24131 , 1'b1 );
or \U$15439 ( \24133 , \24132 , 1'b0 );
buf \U$15440 ( \24134 , \24133 );
_DC r254b6_GF_IsGateDCbyConstraint ( \24135_nR254b6 , \24134 , \21944 );
buf \U$15441 ( \24136 , \24135_nR254b6 );
not \U$15442 ( \24137 , \23755 );
and \U$15443 ( \24138 , RIdb4c330_3814, \24137 );
not \U$15444 ( \24139 , RIdb4c330_3814);
or \U$15445 ( \24140 , \24139 , \23553 );
not \U$15446 ( \24141 , \23649 );
and \U$15447 ( \24142 , \22908 , \24141 );
not \U$15448 ( \24143 , \24142 );
not \U$15449 ( \24144 , \22905 );
not \U$15450 ( \24145 , \23596 );
or \U$15451 ( \24146 , \24144 , \24145 );
nand \U$15452 ( \24147 , \24140 , \24143 , \24146 );
and \U$15453 ( \24148 , \24147 , \23755 );
or \U$15454 ( \24149 , \24138 , \24148 );
and \U$15456 ( \24150 , \24149 , 1'b1 );
or \U$15458 ( \24151 , \24150 , 1'b0 );
buf \U$15459 ( \24152 , \24151 );
_DC r254b8_GF_IsGateDCbyConstraint ( \24153_nR254b8 , \24152 , \21944 );
buf \U$15460 ( \24154 , \24153_nR254b8 );
buf \U$15461 ( \24155 , \22103 );
buf \U$15462 ( \24156 , \24155 );
not \U$15463 ( \24157 , \24156 );
and \U$15464 ( \24158 , RIdb4d410_3815, \24157 );
not \U$15465 ( \24159 , RIdb4d410_3815);
or \U$15466 ( \24160 , \24159 , \23532 );
not \U$15467 ( \24161 , \23630 );
and \U$15468 ( \24162 , \22928 , \24161 );
not \U$15469 ( \24163 , \24162 );
not \U$15470 ( \24164 , \22925 );
not \U$15471 ( \24165 , \23462 );
or \U$15472 ( \24166 , \24164 , \24165 );
nand \U$15473 ( \24167 , \24160 , \24163 , \24166 );
and \U$15474 ( \24168 , \24167 , \24156 );
or \U$15475 ( \24169 , \24158 , \24168 );
and \U$15477 ( \24170 , \24169 , 1'b1 );
or \U$15479 ( \24171 , \24170 , 1'b0 );
buf \U$15480 ( \24172 , \24171 );
_DC r254ba_GF_IsGateDCbyConstraint ( \24173_nR254ba , \24172 , \21944 );
buf \U$15481 ( \24174 , \24173_nR254ba );
not \U$15482 ( \24175 , \24156 );
and \U$15483 ( \24176 , RIdb4e5e0_3816, \24175 );
not \U$15484 ( \24177 , RIdb4e5e0_3816);
or \U$15485 ( \24178 , \24177 , \23628 );
not \U$15486 ( \24179 , \23444 );
and \U$15487 ( \24180 , \22948 , \24179 );
not \U$15488 ( \24181 , \24180 );
not \U$15489 ( \24182 , \22945 );
not \U$15490 ( \24183 , \23538 );
or \U$15491 ( \24184 , \24182 , \24183 );
nand \U$15492 ( \24185 , \24178 , \24181 , \24184 );
and \U$15493 ( \24186 , \24185 , \24156 );
or \U$15494 ( \24187 , \24176 , \24186 );
and \U$15496 ( \24188 , \24187 , 1'b1 );
or \U$15498 ( \24189 , \24188 , 1'b0 );
buf \U$15499 ( \24190 , \24189 );
_DC r254bc_GF_IsGateDCbyConstraint ( \24191_nR254bc , \24190 , \21944 );
buf \U$15500 ( \24192 , \24191_nR254bc );
not \U$15501 ( \24193 , \23755 );
and \U$15502 ( \24194 , RIdb4fa08_3817, \24193 );
not \U$15503 ( \24195 , RIdb4fa08_3817);
or \U$15504 ( \24196 , \24195 , \23628 );
not \U$15505 ( \24197 , \23478 );
and \U$15506 ( \24198 , \22968 , \24197 );
not \U$15507 ( \24199 , \24198 );
not \U$15508 ( \24200 , \22965 );
not \U$15509 ( \24201 , \23462 );
or \U$15510 ( \24202 , \24200 , \24201 );
nand \U$15511 ( \24203 , \24196 , \24199 , \24202 );
and \U$15512 ( \24204 , \24203 , \23755 );
or \U$15513 ( \24205 , \24194 , \24204 );
and \U$15515 ( \24206 , \24205 , 1'b1 );
or \U$15517 ( \24207 , \24206 , 1'b0 );
buf \U$15518 ( \24208 , \24207 );
_DC r254c0_GF_IsGateDCbyConstraint ( \24209_nR254c0 , \24208 , \21944 );
buf \U$15519 ( \24210 , \24209_nR254c0 );
not \U$15520 ( \24211 , \24118 );
and \U$15521 ( \24212 , RIdb51100_3818, \24211 );
not \U$15522 ( \24213 , RIdb51100_3818);
or \U$15523 ( \24214 , \24213 , \23532 );
not \U$15524 ( \24215 , \23555 );
and \U$15525 ( \24216 , \22987 , \24215 );
not \U$15526 ( \24217 , \24216 );
not \U$15527 ( \24218 , \22984 );
not \U$15528 ( \24219 , \23538 );
or \U$15529 ( \24220 , \24218 , \24219 );
nand \U$15530 ( \24221 , \24214 , \24217 , \24220 );
and \U$15531 ( \24222 , \24221 , \24118 );
or \U$15532 ( \24223 , \24212 , \24222 );
and \U$15534 ( \24224 , \24223 , 1'b1 );
or \U$15536 ( \24225 , \24224 , 1'b0 );
buf \U$15537 ( \24226 , \24225 );
_DC r254c2_GF_IsGateDCbyConstraint ( \24227_nR254c2 , \24226 , \21944 );
buf \U$15538 ( \24228 , \24227_nR254c2 );
not \U$15539 ( \24229 , \24156 );
and \U$15540 ( \24230 , RIdb52c30_3819, \24229 );
not \U$15541 ( \24231 , RIdb52c30_3819);
or \U$15542 ( \24232 , \24231 , \23476 );
not \U$15543 ( \24233 , \23630 );
and \U$15544 ( \24234 , \23006 , \24233 );
not \U$15545 ( \24235 , \24234 );
not \U$15546 ( \24236 , \23003 );
not \U$15547 ( \24237 , \23538 );
or \U$15548 ( \24238 , \24236 , \24237 );
nand \U$15549 ( \24239 , \24232 , \24235 , \24238 );
and \U$15550 ( \24240 , \24239 , \24156 );
or \U$15551 ( \24241 , \24230 , \24240 );
and \U$15553 ( \24242 , \24241 , 1'b1 );
or \U$15555 ( \24243 , \24242 , 1'b0 );
buf \U$15556 ( \24244 , \24243 );
_DC r254c4_GF_IsGateDCbyConstraint ( \24245_nR254c4 , \24244 , \21944 );
buf \U$15557 ( \24246 , \24245_nR254c4 );
not \U$15558 ( \24247 , \23755 );
and \U$15559 ( \24248 , RIdb541c0_3820, \24247 );
not \U$15560 ( \24249 , RIdb541c0_3820);
or \U$15561 ( \24250 , \24249 , \23628 );
not \U$15562 ( \24251 , \23686 );
and \U$15563 ( \24252 , \23026 , \24251 );
not \U$15564 ( \24253 , \24252 );
not \U$15565 ( \24254 , \23023 );
not \U$15566 ( \24255 , \23538 );
or \U$15567 ( \24256 , \24254 , \24255 );
nand \U$15568 ( \24257 , \24250 , \24253 , \24256 );
and \U$15569 ( \24258 , \24257 , \23755 );
or \U$15570 ( \24259 , \24248 , \24258 );
and \U$15572 ( \24260 , \24259 , 1'b1 );
or \U$15574 ( \24261 , \24260 , 1'b0 );
buf \U$15575 ( \24262 , \24261 );
_DC r254c6_GF_IsGateDCbyConstraint ( \24263_nR254c6 , \24262 , \21944 );
buf \U$15576 ( \24264 , \24263_nR254c6 );
not \U$15577 ( \24265 , \24156 );
and \U$15578 ( \24266 , RIdb559a8_3821, \24265 );
not \U$15579 ( \24267 , RIdb559a8_3821);
or \U$15580 ( \24268 , \24267 , \23532 );
not \U$15581 ( \24269 , \23940 );
and \U$15582 ( \24270 , \23048 , \24269 );
not \U$15583 ( \24271 , \24270 );
not \U$15584 ( \24272 , \23045 );
not \U$15585 ( \24273 , \23462 );
or \U$15586 ( \24274 , \24272 , \24273 );
nand \U$15587 ( \24275 , \24268 , \24271 , \24274 );
and \U$15588 ( \24276 , \24275 , \24156 );
or \U$15589 ( \24277 , \24266 , \24276 );
and \U$15591 ( \24278 , \24277 , 1'b1 );
or \U$15593 ( \24279 , \24278 , 1'b0 );
buf \U$15594 ( \24280 , \24279 );
_DC r254c8_GF_IsGateDCbyConstraint ( \24281_nR254c8 , \24280 , \21944 );
buf \U$15595 ( \24282 , \24281_nR254c8 );
not \U$15596 ( \24283 , \24156 );
and \U$15597 ( \24284 , RIdb56e48_3822, \24283 );
not \U$15598 ( \24285 , RIdb56e48_3822);
or \U$15599 ( \24286 , \24285 , \23453 );
not \U$15600 ( \24287 , \23686 );
and \U$15601 ( \24288 , \23068 , \24287 );
not \U$15602 ( \24289 , \24288 );
not \U$15603 ( \24290 , \23065 );
not \U$15604 ( \24291 , \23538 );
or \U$15605 ( \24292 , \24290 , \24291 );
nand \U$15606 ( \24293 , \24286 , \24289 , \24292 );
and \U$15607 ( \24294 , \24293 , \24156 );
or \U$15608 ( \24295 , \24284 , \24294 );
and \U$15610 ( \24296 , \24295 , 1'b1 );
or \U$15612 ( \24297 , \24296 , 1'b0 );
buf \U$15613 ( \24298 , \24297 );
_DC r254ca_GF_IsGateDCbyConstraint ( \24299_nR254ca , \24298 , \21944 );
buf \U$15614 ( \24300 , \24299_nR254ca );
not \U$15615 ( \24301 , \23755 );
and \U$15616 ( \24302 , RIdb58900_3823, \24301 );
not \U$15617 ( \24303 , RIdb58900_3823);
or \U$15618 ( \24304 , \24303 , \23532 );
not \U$15619 ( \24305 , \23555 );
and \U$15620 ( \24306 , \23088 , \24305 );
not \U$15621 ( \24307 , \24306 );
not \U$15622 ( \24308 , \23085 );
not \U$15623 ( \24309 , \23462 );
or \U$15624 ( \24310 , \24308 , \24309 );
nand \U$15625 ( \24311 , \24304 , \24307 , \24310 );
and \U$15626 ( \24312 , \24311 , \23755 );
or \U$15627 ( \24313 , \24302 , \24312 );
and \U$15629 ( \24314 , \24313 , 1'b1 );
or \U$15631 ( \24315 , \24314 , 1'b0 );
buf \U$15632 ( \24316 , \24315 );
_DC r254cc_GF_IsGateDCbyConstraint ( \24317_nR254cc , \24316 , \21944 );
buf \U$15633 ( \24318 , \24317_nR254cc );
not \U$15634 ( \24319 , \24118 );
and \U$15635 ( \24320 , RIdb5a070_3824, \24319 );
not \U$15636 ( \24321 , RIdb5a070_3824);
or \U$15637 ( \24322 , \24321 , \23553 );
not \U$15638 ( \24323 , \23630 );
and \U$15639 ( \24324 , \23108 , \24323 );
not \U$15640 ( \24325 , \24324 );
not \U$15641 ( \24326 , \23105 );
not \U$15642 ( \24327 , \23596 );
or \U$15643 ( \24328 , \24326 , \24327 );
nand \U$15644 ( \24329 , \24322 , \24325 , \24328 );
and \U$15645 ( \24330 , \24329 , \24118 );
or \U$15646 ( \24331 , \24320 , \24330 );
and \U$15648 ( \24332 , \24331 , 1'b1 );
or \U$15650 ( \24333 , \24332 , 1'b0 );
buf \U$15651 ( \24334 , \24333 );
_DC r254ce_GF_IsGateDCbyConstraint ( \24335_nR254ce , \24334 , \21944 );
buf \U$15652 ( \24336 , \24335_nR254ce );
not \U$15653 ( \24337 , \24118 );
and \U$15654 ( \24338 , RIdb5b588_3825, \24337 );
not \U$15655 ( \24339 , RIdb5b588_3825);
or \U$15656 ( \24340 , \24339 , \23453 );
not \U$15657 ( \24341 , \23686 );
and \U$15658 ( \24342 , \23128 , \24341 );
not \U$15659 ( \24343 , \24342 );
not \U$15660 ( \24344 , \23125 );
not \U$15661 ( \24345 , \23462 );
or \U$15662 ( \24346 , \24344 , \24345 );
nand \U$15663 ( \24347 , \24340 , \24343 , \24346 );
and \U$15664 ( \24348 , \24347 , \24118 );
or \U$15665 ( \24349 , \24338 , \24348 );
and \U$15667 ( \24350 , \24349 , 1'b1 );
or \U$15669 ( \24351 , \24350 , 1'b0 );
buf \U$15670 ( \24352 , \24351 );
_DC r254d0_GF_IsGateDCbyConstraint ( \24353_nR254d0 , \24352 , \21944 );
buf \U$15671 ( \24354 , \24353_nR254d0 );
not \U$15672 ( \24355 , \23755 );
and \U$15673 ( \24356 , RIdb5d0b8_3826, \24355 );
not \U$15674 ( \24357 , RIdb5d0b8_3826);
or \U$15675 ( \24358 , \24357 , \23453 );
not \U$15676 ( \24359 , \23940 );
and \U$15677 ( \24360 , \23148 , \24359 );
not \U$15678 ( \24361 , \24360 );
not \U$15679 ( \24362 , \23145 );
not \U$15680 ( \24363 , \23596 );
or \U$15681 ( \24364 , \24362 , \24363 );
nand \U$15682 ( \24365 , \24358 , \24361 , \24364 );
and \U$15683 ( \24366 , \24365 , \23755 );
or \U$15684 ( \24367 , \24356 , \24366 );
and \U$15686 ( \24368 , \24367 , 1'b1 );
or \U$15688 ( \24369 , \24368 , 1'b0 );
buf \U$15689 ( \24370 , \24369 );
_DC r254d2_GF_IsGateDCbyConstraint ( \24371_nR254d2 , \24370 , \21944 );
buf \U$15690 ( \24372 , \24371_nR254d2 );
not \U$15691 ( \24373 , \24118 );
and \U$15692 ( \24374 , RIdb5e3f0_3827, \24373 );
not \U$15693 ( \24375 , RIdb5e3f0_3827);
or \U$15694 ( \24376 , \24375 , \23553 );
not \U$15695 ( \24377 , \23555 );
and \U$15696 ( \24378 , \23168 , \24377 );
not \U$15697 ( \24379 , \24378 );
not \U$15698 ( \24380 , \23165 );
not \U$15699 ( \24381 , \23538 );
or \U$15700 ( \24382 , \24380 , \24381 );
nand \U$15701 ( \24383 , \24376 , \24379 , \24382 );
and \U$15702 ( \24384 , \24383 , \24118 );
or \U$15703 ( \24385 , \24374 , \24384 );
and \U$15705 ( \24386 , \24385 , 1'b1 );
or \U$15707 ( \24387 , \24386 , 1'b0 );
buf \U$15708 ( \24388 , \24387 );
_DC r254d6_GF_IsGateDCbyConstraint ( \24389_nR254d6 , \24388 , \21944 );
buf \U$15709 ( \24390 , \24389_nR254d6 );
not \U$15710 ( \24391 , \24156 );
and \U$15711 ( \24392 , RIda95720_3828, \24391 );
not \U$15712 ( \24393 , RIda95720_3828);
or \U$15713 ( \24394 , \24393 , \23532 );
not \U$15714 ( \24395 , \23649 );
and \U$15715 ( \24396 , \23187 , \24395 );
not \U$15716 ( \24397 , \24396 );
not \U$15717 ( \24398 , \23184 );
not \U$15718 ( \24399 , \23462 );
or \U$15719 ( \24400 , \24398 , \24399 );
nand \U$15720 ( \24401 , \24394 , \24397 , \24400 );
and \U$15721 ( \24402 , \24401 , \24156 );
or \U$15722 ( \24403 , \24392 , \24402 );
and \U$15724 ( \24404 , \24403 , 1'b1 );
or \U$15726 ( \24405 , \24404 , 1'b0 );
buf \U$15727 ( \24406 , \24405 );
_DC r254d8_GF_IsGateDCbyConstraint ( \24407_nR254d8 , \24406 , \21944 );
buf \U$15728 ( \24408 , \24407_nR254d8 );
buf \U$15729 ( \24409 , \24155 );
not \U$15730 ( \24410 , \24409 );
and \U$15731 ( \24411 , RIda97598_3829, \24410 );
not \U$15732 ( \24412 , RIda97598_3829);
or \U$15733 ( \24413 , \24412 , \23553 );
not \U$15734 ( \24414 , \23686 );
and \U$15735 ( \24415 , \23207 , \24414 );
not \U$15736 ( \24416 , \24415 );
not \U$15737 ( \24417 , \23204 );
not \U$15738 ( \24418 , \23461 );
or \U$15739 ( \24419 , \24417 , \24418 );
nand \U$15740 ( \24420 , \24413 , \24416 , \24419 );
and \U$15741 ( \24421 , \24420 , \24409 );
or \U$15742 ( \24422 , \24411 , \24421 );
and \U$15744 ( \24423 , \24422 , 1'b1 );
or \U$15746 ( \24424 , \24423 , 1'b0 );
buf \U$15747 ( \24425 , \24424 );
_DC r254da_GF_IsGateDCbyConstraint ( \24426_nR254da , \24425 , \21944 );
buf \U$15748 ( \24427 , \24426_nR254da );
not \U$15749 ( \24428 , \24118 );
and \U$15750 ( \24429 , RIda99a28_3830, \24428 );
not \U$15751 ( \24430 , RIda99a28_3830);
or \U$15752 ( \24431 , \24430 , \23453 );
not \U$15753 ( \24432 , \23444 );
and \U$15754 ( \24433 , \23227 , \24432 );
not \U$15755 ( \24434 , \24433 );
not \U$15756 ( \24435 , \23224 );
not \U$15757 ( \24436 , \23538 );
or \U$15758 ( \24437 , \24435 , \24436 );
nand \U$15759 ( \24438 , \24431 , \24434 , \24437 );
and \U$15760 ( \24439 , \24438 , \24118 );
or \U$15761 ( \24440 , \24429 , \24439 );
and \U$15763 ( \24441 , \24440 , 1'b1 );
or \U$15765 ( \24442 , \24441 , 1'b0 );
buf \U$15766 ( \24443 , \24442 );
_DC r254dc_GF_IsGateDCbyConstraint ( \24444_nR254dc , \24443 , \21944 );
buf \U$15767 ( \24445 , \24444_nR254dc );
not \U$15768 ( \24446 , \24118 );
and \U$15769 ( \24447 , RIda9bd50_3831, \24446 );
not \U$15770 ( \24448 , RIda9bd50_3831);
or \U$15771 ( \24449 , \24448 , \23476 );
not \U$15772 ( \24450 , \23649 );
and \U$15773 ( \24451 , \23247 , \24450 );
not \U$15774 ( \24452 , \24451 );
not \U$15775 ( \24453 , \23244 );
not \U$15776 ( \24454 , \23461 );
or \U$15777 ( \24455 , \24453 , \24454 );
nand \U$15778 ( \24456 , \24449 , \24452 , \24455 );
and \U$15779 ( \24457 , \24456 , \24118 );
or \U$15780 ( \24458 , \24447 , \24457 );
and \U$15782 ( \24459 , \24458 , 1'b1 );
or \U$15784 ( \24460 , \24459 , 1'b0 );
buf \U$15785 ( \24461 , \24460 );
_DC r254de_GF_IsGateDCbyConstraint ( \24462_nR254de , \24461 , \21944 );
buf \U$15786 ( \24463 , \24462_nR254de );
not \U$15787 ( \24464 , \24409 );
and \U$15788 ( \24465 , RIda9df10_3832, \24464 );
not \U$15789 ( \24466 , RIda9df10_3832);
or \U$15790 ( \24467 , \24466 , \23553 );
not \U$15791 ( \24468 , \23456 );
and \U$15792 ( \24469 , \23267 , \24468 );
not \U$15793 ( \24470 , \24469 );
not \U$15794 ( \24471 , \23264 );
not \U$15795 ( \24472 , \23538 );
or \U$15796 ( \24473 , \24471 , \24472 );
nand \U$15797 ( \24474 , \24467 , \24470 , \24473 );
and \U$15798 ( \24475 , \24474 , \24409 );
or \U$15799 ( \24476 , \24465 , \24475 );
and \U$15801 ( \24477 , \24476 , 1'b1 );
or \U$15803 ( \24478 , \24477 , 1'b0 );
buf \U$15804 ( \24479 , \24478 );
_DC r254e0_GF_IsGateDCbyConstraint ( \24480_nR254e0 , \24479 , \21944 );
buf \U$15805 ( \24481 , \24480_nR254e0 );
not \U$15806 ( \24482 , \24156 );
and \U$15807 ( \24483 , RIda9f4a0_3833, \24482 );
not \U$15808 ( \24484 , RIda9f4a0_3833);
or \U$15809 ( \24485 , \24484 , \23628 );
not \U$15810 ( \24486 , \23478 );
and \U$15811 ( \24487 , \23287 , \24486 );
not \U$15812 ( \24488 , \24487 );
not \U$15813 ( \24489 , \23284 );
not \U$15814 ( \24490 , \23538 );
or \U$15815 ( \24491 , \24489 , \24490 );
nand \U$15816 ( \24492 , \24485 , \24488 , \24491 );
and \U$15817 ( \24493 , \24492 , \24156 );
or \U$15818 ( \24494 , \24483 , \24493 );
and \U$15820 ( \24495 , \24494 , 1'b1 );
or \U$15822 ( \24496 , \24495 , 1'b0 );
buf \U$15823 ( \24497 , \24496 );
_DC r254e2_GF_IsGateDCbyConstraint ( \24498_nR254e2 , \24497 , \21944 );
buf \U$15824 ( \24499 , \24498_nR254e2 );
not \U$15825 ( \24500 , \24156 );
and \U$15826 ( \24501 , RIdaa1228_3834, \24500 );
not \U$15827 ( \24502 , RIdaa1228_3834);
or \U$15828 ( \24503 , \24502 , \23532 );
not \U$15829 ( \24504 , \23649 );
and \U$15830 ( \24505 , \23306 , \24504 );
not \U$15831 ( \24506 , \24505 );
not \U$15832 ( \24507 , \23303 );
not \U$15833 ( \24508 , \23462 );
or \U$15834 ( \24509 , \24507 , \24508 );
nand \U$15835 ( \24510 , \24503 , \24506 , \24509 );
and \U$15836 ( \24511 , \24510 , \24156 );
or \U$15837 ( \24512 , \24501 , \24511 );
and \U$15839 ( \24513 , \24512 , 1'b1 );
or \U$15841 ( \24514 , \24513 , 1'b0 );
buf \U$15842 ( \24515 , \24514 );
_DC r254e4_GF_IsGateDCbyConstraint ( \24516_nR254e4 , \24515 , \21944 );
buf \U$15843 ( \24517 , \24516_nR254e4 );
not \U$15844 ( \24518 , \24409 );
and \U$15845 ( \24519 , RIdaa2d58_3835, \24518 );
not \U$15846 ( \24520 , RIdaa2d58_3835);
or \U$15847 ( \24521 , \24520 , \23476 );
not \U$15848 ( \24522 , \23478 );
and \U$15849 ( \24523 , \23326 , \24522 );
not \U$15850 ( \24524 , \24523 );
not \U$15851 ( \24525 , \23323 );
not \U$15852 ( \24526 , \23538 );
or \U$15853 ( \24527 , \24525 , \24526 );
nand \U$15854 ( \24528 , \24521 , \24524 , \24527 );
and \U$15855 ( \24529 , \24528 , \24409 );
or \U$15856 ( \24530 , \24519 , \24529 );
and \U$15858 ( \24531 , \24530 , 1'b1 );
or \U$15860 ( \24532 , \24531 , 1'b0 );
buf \U$15861 ( \24533 , \24532 );
_DC r254e6_GF_IsGateDCbyConstraint ( \24534_nR254e6 , \24533 , \21944 );
buf \U$15862 ( \24535 , \24534_nR254e6 );
not \U$15863 ( \24536 , \24118 );
and \U$15864 ( \24537 , RIdaa4a68_3836, \24536 );
not \U$15865 ( \24538 , RIdaa4a68_3836);
or \U$15866 ( \24539 , \24538 , \23553 );
not \U$15867 ( \24540 , \23478 );
and \U$15868 ( \24541 , \23346 , \24540 );
not \U$15869 ( \24542 , \24541 );
not \U$15870 ( \24543 , \23343 );
not \U$15871 ( \24544 , \23538 );
or \U$15872 ( \24545 , \24543 , \24544 );
nand \U$15873 ( \24546 , \24539 , \24542 , \24545 );
and \U$15874 ( \24547 , \24546 , \24118 );
or \U$15875 ( \24548 , \24537 , \24547 );
and \U$15877 ( \24549 , \24548 , 1'b1 );
or \U$15879 ( \24550 , \24549 , 1'b0 );
buf \U$15880 ( \24551 , \24550 );
_DC r254e8_GF_IsGateDCbyConstraint ( \24552_nR254e8 , \24551 , \21944 );
buf \U$15881 ( \24553 , \24552_nR254e8 );
not \U$15882 ( \24554 , \24118 );
and \U$15883 ( \24555 , RIdaa6b38_3837, \24554 );
not \U$15884 ( \24556 , RIdaa6b38_3837);
or \U$15885 ( \24557 , \24556 , \23453 );
not \U$15886 ( \24558 , \23630 );
and \U$15887 ( \24559 , \23367 , \24558 );
not \U$15888 ( \24560 , \24559 );
not \U$15889 ( \24561 , \23364 );
not \U$15890 ( \24562 , \23538 );
or \U$15891 ( \24563 , \24561 , \24562 );
nand \U$15892 ( \24564 , \24557 , \24560 , \24563 );
and \U$15893 ( \24565 , \24564 , \24118 );
or \U$15894 ( \24566 , \24555 , \24565 );
and \U$15896 ( \24567 , \24566 , 1'b1 );
or \U$15898 ( \24568 , \24567 , 1'b0 );
buf \U$15899 ( \24569 , \24568 );
_DC r254ec_GF_IsGateDCbyConstraint ( \24570_nR254ec , \24569 , \21944 );
buf \U$15900 ( \24571 , \24570_nR254ec );
not \U$15901 ( \24572 , \24409 );
and \U$15902 ( \24573 , RIdaa89b0_3838, \24572 );
not \U$15903 ( \24574 , RIdaa89b0_3838);
or \U$15904 ( \24575 , \24574 , \23628 );
not \U$15905 ( \24576 , \23686 );
and \U$15906 ( \24577 , \23387 , \24576 );
not \U$15907 ( \24578 , \24577 );
not \U$15908 ( \24579 , \23384 );
not \U$15909 ( \24580 , \23538 );
or \U$15910 ( \24581 , \24579 , \24580 );
nand \U$15911 ( \24582 , \24575 , \24578 , \24581 );
and \U$15912 ( \24583 , \24582 , \24409 );
or \U$15913 ( \24584 , \24573 , \24583 );
and \U$15915 ( \24585 , \24584 , 1'b1 );
or \U$15917 ( \24586 , \24585 , 1'b0 );
buf \U$15918 ( \24587 , \24586 );
_DC r254ee_GF_IsGateDCbyConstraint ( \24588_nR254ee , \24587 , \21944 );
buf \U$15919 ( \24589 , \24588_nR254ee );
not \U$15920 ( \24590 , \24156 );
and \U$15921 ( \24591 , RIdbdf030_3839, \24590 );
not \U$15922 ( \24592 , RIdbdf030_3839);
or \U$15923 ( \24593 , \24592 , \23476 );
not \U$15924 ( \24594 , \23940 );
and \U$15925 ( \24595 , \23407 , \24594 );
not \U$15926 ( \24596 , \24595 );
not \U$15927 ( \24597 , \23404 );
not \U$15928 ( \24598 , \23538 );
or \U$15929 ( \24599 , \24597 , \24598 );
nand \U$15930 ( \24600 , \24593 , \24596 , \24599 );
and \U$15931 ( \24601 , \24600 , \24156 );
or \U$15932 ( \24602 , \24591 , \24601 );
and \U$15934 ( \24603 , \24602 , 1'b1 );
or \U$15936 ( \24604 , \24603 , 1'b0 );
buf \U$15937 ( \24605 , \24604 );
_DC r254f0_GF_IsGateDCbyConstraint ( \24606_nR254f0 , \24605 , \21944 );
buf \U$15938 ( \24607 , \24606_nR254f0 );
not \U$15939 ( \24608 , \24409 );
and \U$15940 ( \24609 , RIdbdcd80_3840, \24608 );
not \U$15941 ( \24610 , RIdbdcd80_3840);
or \U$15942 ( \24611 , \24610 , \23628 );
not \U$15943 ( \24612 , \23456 );
and \U$15944 ( \24613 , \23427 , \24612 );
not \U$15945 ( \24614 , \24613 );
not \U$15946 ( \24615 , \23424 );
not \U$15947 ( \24616 , \23538 );
or \U$15948 ( \24617 , \24615 , \24616 );
nand \U$15949 ( \24618 , \24611 , \24614 , \24617 );
and \U$15950 ( \24619 , \24618 , \24409 );
or \U$15951 ( \24620 , \24609 , \24619 );
and \U$15953 ( \24621 , \24620 , 1'b1 );
or \U$15955 ( \24622 , \24621 , 1'b0 );
buf \U$15956 ( \24623 , \24622 );
_DC r254f2_GF_IsGateDCbyConstraint ( \24624_nR254f2 , \24623 , \21944 );
buf \U$15957 ( \24625 , \24624_nR254f2 );
not \U$15958 ( \24626 , \24118 );
and \U$15959 ( \24627 , RIdbdaff8_3841, \24626 );
not \U$15960 ( \24628 , RIdbdaff8_3841);
not \U$15961 ( \24629 , \22117 );
nor \U$15962 ( \24630 , \22121 , \24629 );
nand \U$15963 ( \24631 , \24630 , \22123 );
not \U$15964 ( \24632 , \24631 );
not \U$15965 ( \24633 , \22111 );
or \U$15966 ( \24634 , \22110 , \24633 );
not \U$15967 ( \24635 , \24634 );
nand \U$15968 ( \24636 , \22102 , \24635 );
not \U$15969 ( \24637 , \24636 );
or \U$15970 ( \24638 , \24632 , \24637 );
not \U$15971 ( \24639 , \24638 );
not \U$15972 ( \24640 , \24639 );
or \U$15973 ( \24641 , \24628 , \24640 );
not \U$15974 ( \24642 , \24632 );
not \U$15975 ( \24643 , \24642 );
and \U$15976 ( \24644 , \22135 , \24643 );
not \U$15977 ( \24645 , \24644 );
not \U$15978 ( \24646 , \24636 );
buf \U$15979 ( \24647 , \24646 );
not \U$15980 ( \24648 , \24647 );
or \U$15981 ( \24649 , \23460 , \24648 );
nand \U$15982 ( \24650 , \24641 , \24645 , \24649 );
and \U$15983 ( \24651 , \24650 , \24118 );
or \U$15984 ( \24652 , \24627 , \24651 );
and \U$15986 ( \24653 , \24652 , 1'b1 );
or \U$15988 ( \24654 , \24653 , 1'b0 );
buf \U$15989 ( \24655 , \24654 );
_DC r254fc_GF_IsGateDCbyConstraint ( \24656_nR254fc , \24655 , \21944 );
buf \U$15990 ( \24657 , \24656_nR254fc );
not \U$15991 ( \24658 , \24409 );
and \U$15992 ( \24659 , RIdbd9540_3842, \24658 );
not \U$15993 ( \24660 , RIdbd9540_3842);
not \U$15994 ( \24661 , \24639 );
or \U$15995 ( \24662 , \24660 , \24661 );
not \U$15996 ( \24663 , \24642 );
and \U$15997 ( \24664 , \22162 , \24663 );
not \U$15998 ( \24665 , \24664 );
buf \U$15999 ( \24666 , \24646 );
not \U$16000 ( \24667 , \24666 );
or \U$16001 ( \24668 , \23482 , \24667 );
nand \U$16002 ( \24669 , \24662 , \24665 , \24668 );
and \U$16003 ( \24670 , \24669 , \24409 );
or \U$16004 ( \24671 , \24659 , \24670 );
and \U$16006 ( \24672 , \24671 , 1'b1 );
or \U$16008 ( \24673 , \24672 , 1'b0 );
buf \U$16009 ( \24674 , \24673 );
_DC r25512_GF_IsGateDCbyConstraint ( \24675_nR25512 , \24674 , \21944 );
buf \U$16010 ( \24676 , \24675_nR25512 );
not \U$16011 ( \24677 , \24156 );
and \U$16012 ( \24678 , RIdbd6e58_3843, \24677 );
not \U$16013 ( \24679 , RIdbd6e58_3843);
or \U$16014 ( \24680 , \24679 , \24661 );
not \U$16015 ( \24681 , \24642 );
and \U$16016 ( \24682 , \22183 , \24681 );
not \U$16017 ( \24683 , \24682 );
not \U$16018 ( \24684 , \24647 );
or \U$16019 ( \24685 , \23500 , \24684 );
nand \U$16020 ( \24686 , \24680 , \24683 , \24685 );
and \U$16021 ( \24687 , \24686 , \24156 );
or \U$16022 ( \24688 , \24678 , \24687 );
and \U$16024 ( \24689 , \24688 , 1'b1 );
or \U$16026 ( \24690 , \24689 , 1'b0 );
buf \U$16027 ( \24691 , \24690 );
_DC r25528_GF_IsGateDCbyConstraint ( \24692_nR25528 , \24691 , \21944 );
buf \U$16028 ( \24693 , \24692_nR25528 );
not \U$16029 ( \24694 , \24118 );
and \U$16030 ( \24695 , RIdbd4860_3844, \24694 );
not \U$16031 ( \24696 , RIdbd4860_3844);
or \U$16032 ( \24697 , \24696 , \24661 );
not \U$16033 ( \24698 , \24632 );
not \U$16034 ( \24699 , \24698 );
and \U$16035 ( \24700 , \22206 , \24699 );
not \U$16036 ( \24701 , \24700 );
not \U$16037 ( \24702 , \24666 );
or \U$16038 ( \24703 , \23518 , \24702 );
nand \U$16039 ( \24704 , \24697 , \24701 , \24703 );
and \U$16040 ( \24705 , \24704 , \24118 );
or \U$16041 ( \24706 , \24695 , \24705 );
and \U$16043 ( \24707 , \24706 , 1'b1 );
or \U$16045 ( \24708 , \24707 , 1'b0 );
buf \U$16046 ( \24709 , \24708 );
_DC r2553e_GF_IsGateDCbyConstraint ( \24710_nR2553e , \24709 , \21944 );
buf \U$16047 ( \24711 , \24710_nR2553e );
not \U$16048 ( \24712 , \24409 );
and \U$16049 ( \24713 , RIdbd25b0_3845, \24712 );
not \U$16050 ( \24714 , RIdbd25b0_3845);
not \U$16051 ( \24715 , \24639 );
or \U$16052 ( \24716 , \24714 , \24715 );
not \U$16053 ( \24717 , \24642 );
and \U$16054 ( \24718 , \22227 , \24717 );
not \U$16055 ( \24719 , \24718 );
buf \U$16056 ( \24720 , \24646 );
not \U$16057 ( \24721 , \24720 );
or \U$16058 ( \24722 , \23537 , \24721 );
nand \U$16059 ( \24723 , \24716 , \24719 , \24722 );
and \U$16060 ( \24724 , \24723 , \24409 );
or \U$16061 ( \24725 , \24713 , \24724 );
and \U$16063 ( \24726 , \24725 , 1'b1 );
or \U$16065 ( \24727 , \24726 , 1'b0 );
buf \U$16066 ( \24728 , \24727 );
_DC r25554_GF_IsGateDCbyConstraint ( \24729_nR25554 , \24728 , \21944 );
buf \U$16067 ( \24730 , \24729_nR25554 );
not \U$16068 ( \24731 , \24156 );
and \U$16069 ( \24732 , RIdbd0030_3846, \24731 );
not \U$16070 ( \24733 , RIdbd0030_3846);
not \U$16071 ( \24734 , \24639 );
or \U$16072 ( \24735 , \24733 , \24734 );
not \U$16073 ( \24736 , \24632 );
not \U$16074 ( \24737 , \24736 );
and \U$16075 ( \24738 , \22249 , \24737 );
not \U$16076 ( \24739 , \24738 );
nand \U$16077 ( \24740 , \22246 , \24666 );
nand \U$16078 ( \24741 , \24735 , \24739 , \24740 );
and \U$16079 ( \24742 , \24741 , \24156 );
or \U$16080 ( \24743 , \24732 , \24742 );
and \U$16082 ( \24744 , \24743 , 1'b1 );
or \U$16084 ( \24745 , \24744 , 1'b0 );
buf \U$16085 ( \24746 , \24745 );
_DC r2556a_GF_IsGateDCbyConstraint ( \24747_nR2556a , \24746 , \21944 );
buf \U$16086 ( \24748 , \24747_nR2556a );
not \U$16087 ( \24749 , \24118 );
and \U$16088 ( \24750 , RIdbcdc18_3847, \24749 );
not \U$16089 ( \24751 , RIdbcdc18_3847);
or \U$16090 ( \24752 , \24751 , \24661 );
not \U$16091 ( \24753 , \24632 );
not \U$16092 ( \24754 , \24753 );
and \U$16093 ( \24755 , \22275 , \24754 );
not \U$16094 ( \24756 , \24755 );
nand \U$16095 ( \24757 , \22272 , \24720 );
nand \U$16096 ( \24758 , \24752 , \24756 , \24757 );
and \U$16097 ( \24759 , \24758 , \24118 );
or \U$16098 ( \24760 , \24750 , \24759 );
and \U$16100 ( \24761 , \24760 , 1'b1 );
or \U$16102 ( \24762 , \24761 , 1'b0 );
buf \U$16103 ( \24763 , \24762 );
_DC r25574_GF_IsGateDCbyConstraint ( \24764_nR25574 , \24763 , \21944 );
buf \U$16104 ( \24765 , \24764_nR25574 );
not \U$16105 ( \24766 , \24409 );
and \U$16106 ( \24767 , RIdbcb800_3848, \24766 );
not \U$16107 ( \24768 , RIdbcb800_3848);
or \U$16108 ( \24769 , \24768 , \24661 );
not \U$16109 ( \24770 , \24698 );
and \U$16110 ( \24771 , \22295 , \24770 );
not \U$16111 ( \24772 , \24771 );
not \U$16112 ( \24773 , \24666 );
or \U$16113 ( \24774 , \23595 , \24773 );
nand \U$16114 ( \24775 , \24769 , \24772 , \24774 );
and \U$16115 ( \24776 , \24775 , \24409 );
or \U$16116 ( \24777 , \24767 , \24776 );
and \U$16118 ( \24778 , \24777 , 1'b1 );
or \U$16120 ( \24779 , \24778 , 1'b0 );
buf \U$16121 ( \24780 , \24779 );
_DC r25576_GF_IsGateDCbyConstraint ( \24781_nR25576 , \24780 , \21944 );
buf \U$16122 ( \24782 , \24781_nR25576 );
not \U$16123 ( \24783 , \24156 );
and \U$16124 ( \24784 , RIdbc9730_3849, \24783 );
not \U$16125 ( \24785 , RIdbc9730_3849);
or \U$16126 ( \24786 , \24785 , \24640 );
not \U$16127 ( \24787 , \24753 );
and \U$16128 ( \24788 , \22317 , \24787 );
not \U$16129 ( \24789 , \24788 );
not \U$16130 ( \24790 , \24720 );
or \U$16131 ( \24791 , \23614 , \24790 );
nand \U$16132 ( \24792 , \24786 , \24789 , \24791 );
and \U$16133 ( \24793 , \24792 , \24156 );
or \U$16134 ( \24794 , \24784 , \24793 );
and \U$16136 ( \24795 , \24794 , 1'b1 );
or \U$16138 ( \24796 , \24795 , 1'b0 );
buf \U$16139 ( \24797 , \24796 );
_DC r25578_GF_IsGateDCbyConstraint ( \24798_nR25578 , \24797 , \21944 );
buf \U$16140 ( \24799 , \24798_nR25578 );
not \U$16141 ( \24800 , \24117 );
and \U$16142 ( \24801 , RIdbc7a20_3850, \24800 );
not \U$16143 ( \24802 , RIdbc7a20_3850);
not \U$16144 ( \24803 , \24639 );
or \U$16145 ( \24804 , \24802 , \24803 );
not \U$16146 ( \24805 , \24753 );
and \U$16147 ( \24806 , \22338 , \24805 );
not \U$16148 ( \24807 , \24806 );
not \U$16149 ( \24808 , \24720 );
or \U$16150 ( \24809 , \23634 , \24808 );
nand \U$16151 ( \24810 , \24804 , \24807 , \24809 );
and \U$16152 ( \24811 , \24810 , \24117 );
or \U$16153 ( \24812 , \24801 , \24811 );
and \U$16155 ( \24813 , \24812 , 1'b1 );
or \U$16157 ( \24814 , \24813 , 1'b0 );
buf \U$16158 ( \24815 , \24814 );
_DC r2557a_GF_IsGateDCbyConstraint ( \24816_nR2557a , \24815 , \21944 );
buf \U$16159 ( \24817 , \24816_nR2557a );
not \U$16160 ( \24818 , \24409 );
and \U$16161 ( \24819 , RIdbc5e78_3851, \24818 );
not \U$16162 ( \24820 , RIdbc5e78_3851);
or \U$16163 ( \24821 , \24820 , \24715 );
not \U$16164 ( \24822 , \24632 );
not \U$16165 ( \24823 , \24822 );
and \U$16166 ( \24824 , \22360 , \24823 );
not \U$16167 ( \24825 , \24824 );
not \U$16168 ( \24826 , \24647 );
or \U$16169 ( \24827 , \23653 , \24826 );
nand \U$16170 ( \24828 , \24821 , \24825 , \24827 );
and \U$16171 ( \24829 , \24828 , \24409 );
or \U$16172 ( \24830 , \24819 , \24829 );
and \U$16174 ( \24831 , \24830 , 1'b1 );
or \U$16176 ( \24832 , \24831 , 1'b0 );
buf \U$16177 ( \24833 , \24832 );
_DC r254fe_GF_IsGateDCbyConstraint ( \24834_nR254fe , \24833 , \21944 );
buf \U$16178 ( \24835 , \24834_nR254fe );
not \U$16179 ( \24836 , \24156 );
and \U$16180 ( \24837 , RIdbc40f0_3852, \24836 );
not \U$16181 ( \24838 , RIdbc40f0_3852);
or \U$16182 ( \24839 , \24838 , \24734 );
not \U$16183 ( \24840 , \24822 );
and \U$16184 ( \24841 , \22380 , \24840 );
not \U$16185 ( \24842 , \24841 );
not \U$16186 ( \24843 , \24647 );
or \U$16187 ( \24844 , \23671 , \24843 );
nand \U$16188 ( \24845 , \24839 , \24842 , \24844 );
and \U$16189 ( \24846 , \24845 , \24156 );
or \U$16190 ( \24847 , \24837 , \24846 );
and \U$16192 ( \24848 , \24847 , 1'b1 );
or \U$16194 ( \24849 , \24848 , 1'b0 );
buf \U$16195 ( \24850 , \24849 );
_DC r25500_GF_IsGateDCbyConstraint ( \24851_nR25500 , \24850 , \21944 );
buf \U$16196 ( \24852 , \24851_nR25500 );
not \U$16197 ( \24853 , \24117 );
and \U$16198 ( \24854 , RIdbc1f30_3853, \24853 );
not \U$16199 ( \24855 , RIdbc1f30_3853);
or \U$16200 ( \24856 , \24855 , \24661 );
not \U$16201 ( \24857 , \24698 );
and \U$16202 ( \24858 , \22401 , \24857 );
not \U$16203 ( \24859 , \24858 );
not \U$16204 ( \24860 , \24666 );
or \U$16205 ( \24861 , \23690 , \24860 );
nand \U$16206 ( \24862 , \24856 , \24859 , \24861 );
and \U$16207 ( \24863 , \24862 , \24117 );
or \U$16208 ( \24864 , \24854 , \24863 );
and \U$16210 ( \24865 , \24864 , 1'b1 );
or \U$16212 ( \24866 , \24865 , 1'b0 );
buf \U$16213 ( \24867 , \24866 );
_DC r25502_GF_IsGateDCbyConstraint ( \24868_nR25502 , \24867 , \21944 );
buf \U$16214 ( \24869 , \24868_nR25502 );
not \U$16215 ( \24870 , \24409 );
and \U$16216 ( \24871 , RIdbbf938_3854, \24870 );
not \U$16217 ( \24872 , RIdbbf938_3854);
or \U$16218 ( \24873 , \24872 , \24803 );
not \U$16219 ( \24874 , \24642 );
and \U$16220 ( \24875 , \22421 , \24874 );
not \U$16221 ( \24876 , \24875 );
not \U$16222 ( \24877 , \24647 );
or \U$16223 ( \24878 , \23708 , \24877 );
nand \U$16224 ( \24879 , \24873 , \24876 , \24878 );
and \U$16225 ( \24880 , \24879 , \24409 );
or \U$16226 ( \24881 , \24871 , \24880 );
and \U$16228 ( \24882 , \24881 , 1'b1 );
or \U$16230 ( \24883 , \24882 , 1'b0 );
buf \U$16231 ( \24884 , \24883 );
_DC r25504_GF_IsGateDCbyConstraint ( \24885_nR25504 , \24884 , \21944 );
buf \U$16232 ( \24886 , \24885_nR25504 );
not \U$16233 ( \24887 , \24156 );
and \U$16234 ( \24888 , RIdbbd4a8_3855, \24887 );
not \U$16235 ( \24889 , RIdbbd4a8_3855);
or \U$16236 ( \24890 , \24889 , \24803 );
not \U$16237 ( \24891 , \24642 );
and \U$16238 ( \24892 , \22441 , \24891 );
not \U$16239 ( \24893 , \24892 );
not \U$16240 ( \24894 , \24666 );
or \U$16241 ( \24895 , \23726 , \24894 );
nand \U$16242 ( \24896 , \24890 , \24893 , \24895 );
and \U$16243 ( \24897 , \24896 , \24156 );
or \U$16244 ( \24898 , \24888 , \24897 );
and \U$16246 ( \24899 , \24898 , 1'b1 );
or \U$16248 ( \24900 , \24899 , 1'b0 );
buf \U$16249 ( \24901 , \24900 );
_DC r25506_GF_IsGateDCbyConstraint ( \24902_nR25506 , \24901 , \21944 );
buf \U$16250 ( \24903 , \24902_nR25506 );
not \U$16251 ( \24904 , \22756 );
and \U$16252 ( \24905 , RIdbba910_3856, \24904 );
not \U$16253 ( \24906 , RIdbba910_3856);
or \U$16254 ( \24907 , \24906 , \24803 );
not \U$16255 ( \24908 , \24822 );
and \U$16256 ( \24909 , \22461 , \24908 );
not \U$16257 ( \24910 , \24909 );
buf \U$16258 ( \24911 , \24646 );
not \U$16259 ( \24912 , \24911 );
or \U$16260 ( \24913 , \23744 , \24912 );
nand \U$16261 ( \24914 , \24907 , \24910 , \24913 );
and \U$16262 ( \24915 , \24914 , \22756 );
or \U$16263 ( \24916 , \24905 , \24915 );
and \U$16265 ( \24917 , \24916 , 1'b1 );
or \U$16267 ( \24918 , \24917 , 1'b0 );
buf \U$16268 ( \24919 , \24918 );
_DC r25508_GF_IsGateDCbyConstraint ( \24920_nR25508 , \24919 , \21944 );
buf \U$16269 ( \24921 , \24920_nR25508 );
not \U$16270 ( \24922 , \24409 );
and \U$16271 ( \24923 , RIdbb8480_3857, \24922 );
not \U$16272 ( \24924 , RIdbb8480_3857);
or \U$16273 ( \24925 , \24924 , \24640 );
not \U$16274 ( \24926 , \24698 );
and \U$16275 ( \24927 , \22481 , \24926 );
not \U$16276 ( \24928 , \24927 );
not \U$16277 ( \24929 , \24720 );
or \U$16278 ( \24930 , \23763 , \24929 );
nand \U$16279 ( \24931 , \24925 , \24928 , \24930 );
and \U$16280 ( \24932 , \24931 , \24409 );
or \U$16281 ( \24933 , \24923 , \24932 );
and \U$16283 ( \24934 , \24933 , 1'b1 );
or \U$16285 ( \24935 , \24934 , 1'b0 );
buf \U$16286 ( \24936 , \24935 );
_DC r2550a_GF_IsGateDCbyConstraint ( \24937_nR2550a , \24936 , \21944 );
buf \U$16287 ( \24938 , \24937_nR2550a );
not \U$16288 ( \24939 , \24155 );
and \U$16289 ( \24940 , RIdbb58e8_3858, \24939 );
not \U$16290 ( \24941 , RIdbb58e8_3858);
or \U$16291 ( \24942 , \24941 , \24661 );
not \U$16292 ( \24943 , \24753 );
and \U$16293 ( \24944 , \22501 , \24943 );
not \U$16294 ( \24945 , \24944 );
not \U$16295 ( \24946 , \24911 );
or \U$16296 ( \24947 , \23781 , \24946 );
nand \U$16297 ( \24948 , \24942 , \24945 , \24947 );
and \U$16298 ( \24949 , \24948 , \24155 );
or \U$16299 ( \24950 , \24940 , \24949 );
and \U$16301 ( \24951 , \24950 , 1'b1 );
or \U$16303 ( \24952 , \24951 , 1'b0 );
buf \U$16304 ( \24953 , \24952 );
_DC r2550c_GF_IsGateDCbyConstraint ( \24954_nR2550c , \24953 , \21944 );
buf \U$16305 ( \24955 , \24954_nR2550c );
not \U$16306 ( \24956 , \24117 );
and \U$16307 ( \24957 , RIdbb2648_3859, \24956 );
not \U$16308 ( \24958 , RIdbb2648_3859);
or \U$16309 ( \24959 , \24958 , \24640 );
not \U$16310 ( \24960 , \24698 );
and \U$16311 ( \24961 , \22522 , \24960 );
not \U$16312 ( \24962 , \24961 );
not \U$16313 ( \24963 , \24911 );
or \U$16314 ( \24964 , \23799 , \24963 );
nand \U$16315 ( \24965 , \24959 , \24962 , \24964 );
and \U$16316 ( \24966 , \24965 , \24117 );
or \U$16317 ( \24967 , \24957 , \24966 );
and \U$16319 ( \24968 , \24967 , 1'b1 );
or \U$16321 ( \24969 , \24968 , 1'b0 );
buf \U$16322 ( \24970 , \24969 );
_DC r2550e_GF_IsGateDCbyConstraint ( \24971_nR2550e , \24970 , \21944 );
buf \U$16323 ( \24972 , \24971_nR2550e );
not \U$16324 ( \24973 , \24409 );
and \U$16325 ( \24974 , RIdbb0758_3860, \24973 );
not \U$16326 ( \24975 , RIdbb0758_3860);
or \U$16327 ( \24976 , \24975 , \24734 );
not \U$16328 ( \24977 , \24642 );
and \U$16329 ( \24978 , \22542 , \24977 );
not \U$16330 ( \24979 , \24978 );
not \U$16331 ( \24980 , \24647 );
or \U$16332 ( \24981 , \23817 , \24980 );
nand \U$16333 ( \24982 , \24976 , \24979 , \24981 );
and \U$16334 ( \24983 , \24982 , \24409 );
or \U$16335 ( \24984 , \24974 , \24983 );
and \U$16337 ( \24985 , \24984 , 1'b1 );
or \U$16339 ( \24986 , \24985 , 1'b0 );
buf \U$16340 ( \24987 , \24986 );
_DC r25510_GF_IsGateDCbyConstraint ( \24988_nR25510 , \24987 , \21944 );
buf \U$16341 ( \24989 , \24988_nR25510 );
not \U$16342 ( \24990 , \24156 );
and \U$16343 ( \24991 , RIdbad788_3861, \24990 );
not \U$16344 ( \24992 , RIdbad788_3861);
or \U$16345 ( \24993 , \24992 , \24803 );
not \U$16346 ( \24994 , \24736 );
and \U$16347 ( \24995 , \22562 , \24994 );
not \U$16348 ( \24996 , \24995 );
not \U$16349 ( \24997 , \24911 );
or \U$16350 ( \24998 , \23835 , \24997 );
nand \U$16351 ( \24999 , \24993 , \24996 , \24998 );
and \U$16352 ( \25000 , \24999 , \24156 );
or \U$16353 ( \25001 , \24991 , \25000 );
and \U$16355 ( \25002 , \25001 , 1'b1 );
or \U$16357 ( \25003 , \25002 , 1'b0 );
buf \U$16358 ( \25004 , \25003 );
_DC r25514_GF_IsGateDCbyConstraint ( \25005_nR25514 , \25004 , \21944 );
buf \U$16359 ( \25006 , \25005_nR25514 );
not \U$16360 ( \25007 , \22756 );
and \U$16361 ( \25008 , RIdbaad58_3862, \25007 );
not \U$16362 ( \25009 , RIdbaad58_3862);
or \U$16363 ( \25010 , \25009 , \24734 );
not \U$16364 ( \25011 , \24753 );
and \U$16365 ( \25012 , \22582 , \25011 );
not \U$16366 ( \25013 , \25012 );
not \U$16367 ( \25014 , \24911 );
or \U$16368 ( \25015 , \23853 , \25014 );
nand \U$16369 ( \25016 , \25010 , \25013 , \25015 );
and \U$16370 ( \25017 , \25016 , \22756 );
or \U$16371 ( \25018 , \25008 , \25017 );
and \U$16373 ( \25019 , \25018 , 1'b1 );
or \U$16375 ( \25020 , \25019 , 1'b0 );
buf \U$16376 ( \25021 , \25020 );
_DC r25516_GF_IsGateDCbyConstraint ( \25022_nR25516 , \25021 , \21944 );
buf \U$16377 ( \25023 , \25022_nR25516 );
not \U$16378 ( \25024 , \22195 );
and \U$16379 ( \25025 , RIdba7d88_3863, \25024 );
not \U$16380 ( \25026 , RIdba7d88_3863);
or \U$16381 ( \25027 , \25026 , \24715 );
not \U$16382 ( \25028 , \24698 );
and \U$16383 ( \25029 , \22602 , \25028 );
not \U$16384 ( \25030 , \25029 );
not \U$16385 ( \25031 , \24647 );
or \U$16386 ( \25032 , \23871 , \25031 );
nand \U$16387 ( \25033 , \25027 , \25030 , \25032 );
and \U$16388 ( \25034 , \25033 , \22195 );
or \U$16389 ( \25035 , \25025 , \25034 );
and \U$16391 ( \25036 , \25035 , 1'b1 );
or \U$16393 ( \25037 , \25036 , 1'b0 );
buf \U$16394 ( \25038 , \25037 );
_DC r25518_GF_IsGateDCbyConstraint ( \25039_nR25518 , \25038 , \21944 );
buf \U$16395 ( \25040 , \25039_nR25518 );
not \U$16396 ( \25041 , \24156 );
and \U$16397 ( \25042 , RIdba55b0_3864, \25041 );
not \U$16398 ( \25043 , RIdba55b0_3864);
or \U$16399 ( \25044 , \25043 , \24715 );
not \U$16400 ( \25045 , \24753 );
and \U$16401 ( \25046 , \22622 , \25045 );
not \U$16402 ( \25047 , \25046 );
not \U$16403 ( \25048 , \24911 );
or \U$16404 ( \25049 , \23889 , \25048 );
nand \U$16405 ( \25050 , \25044 , \25047 , \25049 );
and \U$16406 ( \25051 , \25050 , \24156 );
or \U$16407 ( \25052 , \25042 , \25051 );
and \U$16409 ( \25053 , \25052 , 1'b1 );
or \U$16411 ( \25054 , \25053 , 1'b0 );
buf \U$16412 ( \25055 , \25054 );
_DC r2551a_GF_IsGateDCbyConstraint ( \25056_nR2551a , \25055 , \21944 );
buf \U$16413 ( \25057 , \25056_nR2551a );
not \U$16414 ( \25058 , \24117 );
and \U$16415 ( \25059 , RIdba2ce8_3865, \25058 );
not \U$16416 ( \25060 , RIdba2ce8_3865);
or \U$16417 ( \25061 , \25060 , \24640 );
not \U$16418 ( \25062 , \24753 );
and \U$16419 ( \25063 , \22643 , \25062 );
not \U$16420 ( \25064 , \25063 );
not \U$16421 ( \25065 , \24911 );
or \U$16422 ( \25066 , \23907 , \25065 );
nand \U$16423 ( \25067 , \25061 , \25064 , \25066 );
and \U$16424 ( \25068 , \25067 , \24117 );
or \U$16425 ( \25069 , \25059 , \25068 );
and \U$16427 ( \25070 , \25069 , 1'b1 );
or \U$16429 ( \25071 , \25070 , 1'b0 );
buf \U$16430 ( \25072 , \25071 );
_DC r2551c_GF_IsGateDCbyConstraint ( \25073_nR2551c , \25072 , \21944 );
buf \U$16431 ( \25074 , \25073_nR2551c );
not \U$16432 ( \25075 , \22195 );
and \U$16433 ( \25076 , RIdb9fe80_3866, \25075 );
not \U$16434 ( \25077 , RIdb9fe80_3866);
or \U$16435 ( \25078 , \25077 , \24715 );
not \U$16436 ( \25079 , \24698 );
and \U$16437 ( \25080 , \22663 , \25079 );
not \U$16438 ( \25081 , \25080 );
not \U$16439 ( \25082 , \24911 );
or \U$16440 ( \25083 , \23925 , \25082 );
nand \U$16441 ( \25084 , \25078 , \25081 , \25083 );
and \U$16442 ( \25085 , \25084 , \22195 );
or \U$16443 ( \25086 , \25076 , \25085 );
and \U$16445 ( \25087 , \25086 , 1'b1 );
or \U$16447 ( \25088 , \25087 , 1'b0 );
buf \U$16448 ( \25089 , \25088 );
_DC r2551e_GF_IsGateDCbyConstraint ( \25090_nR2551e , \25089 , \21944 );
buf \U$16449 ( \25091 , \25090_nR2551e );
not \U$16450 ( \25092 , \24156 );
and \U$16451 ( \25093 , RIdb9d4c8_3867, \25092 );
not \U$16452 ( \25094 , RIdb9d4c8_3867);
or \U$16453 ( \25095 , \25094 , \24640 );
not \U$16454 ( \25096 , \24736 );
and \U$16455 ( \25097 , \22684 , \25096 );
not \U$16456 ( \25098 , \25097 );
not \U$16457 ( \25099 , \24911 );
or \U$16458 ( \25100 , \23944 , \25099 );
nand \U$16459 ( \25101 , \25095 , \25098 , \25100 );
and \U$16460 ( \25102 , \25101 , \24156 );
or \U$16461 ( \25103 , \25093 , \25102 );
and \U$16463 ( \25104 , \25103 , 1'b1 );
or \U$16465 ( \25105 , \25104 , 1'b0 );
buf \U$16466 ( \25106 , \25105 );
_DC r25520_GF_IsGateDCbyConstraint ( \25107_nR25520 , \25106 , \21944 );
buf \U$16467 ( \25108 , \25107_nR25520 );
not \U$16468 ( \25109 , \24117 );
and \U$16469 ( \25110 , RIdb9acf0_3868, \25109 );
not \U$16470 ( \25111 , RIdb9acf0_3868);
or \U$16471 ( \25112 , \25111 , \24734 );
not \U$16472 ( \25113 , \24736 );
and \U$16473 ( \25114 , \22704 , \25113 );
not \U$16474 ( \25115 , \25114 );
not \U$16475 ( \25116 , \24647 );
or \U$16476 ( \25117 , \23962 , \25116 );
nand \U$16477 ( \25118 , \25112 , \25115 , \25117 );
and \U$16478 ( \25119 , \25118 , \24117 );
or \U$16479 ( \25120 , \25110 , \25119 );
and \U$16481 ( \25121 , \25120 , 1'b1 );
or \U$16483 ( \25122 , \25121 , 1'b0 );
buf \U$16484 ( \25123 , \25122 );
_DC r25522_GF_IsGateDCbyConstraint ( \25124_nR25522 , \25123 , \21944 );
buf \U$16485 ( \25125 , \25124_nR25522 );
not \U$16486 ( \25126 , \24117 );
and \U$16487 ( \25127 , RIdb98c20_3869, \25126 );
not \U$16488 ( \25128 , RIdb98c20_3869);
or \U$16489 ( \25129 , \25128 , \24803 );
not \U$16490 ( \25130 , \24698 );
and \U$16491 ( \25131 , \22724 , \25130 );
not \U$16492 ( \25132 , \25131 );
not \U$16493 ( \25133 , \24647 );
or \U$16494 ( \25134 , \23980 , \25133 );
nand \U$16495 ( \25135 , \25129 , \25132 , \25134 );
and \U$16496 ( \25136 , \25135 , \24117 );
or \U$16497 ( \25137 , \25127 , \25136 );
and \U$16499 ( \25138 , \25137 , 1'b1 );
or \U$16501 ( \25139 , \25138 , 1'b0 );
buf \U$16502 ( \25140 , \25139 );
_DC r25524_GF_IsGateDCbyConstraint ( \25141_nR25524 , \25140 , \21944 );
buf \U$16503 ( \25142 , \25141_nR25524 );
not \U$16504 ( \25143 , \24409 );
and \U$16505 ( \25144 , RIdb96178_3870, \25143 );
not \U$16506 ( \25145 , RIdb96178_3870);
or \U$16507 ( \25146 , \25145 , \24640 );
not \U$16508 ( \25147 , \24736 );
and \U$16509 ( \25148 , \22744 , \25147 );
not \U$16510 ( \25149 , \25148 );
not \U$16511 ( \25150 , \24647 );
or \U$16512 ( \25151 , \23998 , \25150 );
nand \U$16513 ( \25152 , \25146 , \25149 , \25151 );
and \U$16514 ( \25153 , \25152 , \24409 );
or \U$16515 ( \25154 , \25144 , \25153 );
and \U$16517 ( \25155 , \25154 , 1'b1 );
or \U$16519 ( \25156 , \25155 , 1'b0 );
buf \U$16520 ( \25157 , \25156 );
_DC r25526_GF_IsGateDCbyConstraint ( \25158_nR25526 , \25157 , \21944 );
buf \U$16521 ( \25159 , \25158_nR25526 );
not \U$16522 ( \25160 , \22756 );
and \U$16523 ( \25161 , RIdb93ce8_3871, \25160 );
not \U$16524 ( \25162 , RIdb93ce8_3871);
or \U$16525 ( \25163 , \25162 , \24803 );
not \U$16526 ( \25164 , \24753 );
and \U$16527 ( \25165 , \22766 , \25164 );
not \U$16528 ( \25166 , \25165 );
not \U$16529 ( \25167 , \24911 );
or \U$16530 ( \25168 , \24016 , \25167 );
nand \U$16531 ( \25169 , \25163 , \25166 , \25168 );
and \U$16532 ( \25170 , \25169 , \22756 );
or \U$16533 ( \25171 , \25161 , \25170 );
and \U$16535 ( \25172 , \25171 , 1'b1 );
or \U$16537 ( \25173 , \25172 , 1'b0 );
buf \U$16538 ( \25174 , \25173 );
_DC r2552a_GF_IsGateDCbyConstraint ( \25175_nR2552a , \25174 , \21944 );
buf \U$16539 ( \25176 , \25175_nR2552a );
not \U$16540 ( \25177 , \22756 );
and \U$16541 ( \25178 , RIdb916f0_3872, \25177 );
not \U$16542 ( \25179 , RIdb916f0_3872);
or \U$16543 ( \25180 , \25179 , \24640 );
not \U$16544 ( \25181 , \24642 );
and \U$16545 ( \25182 , \22786 , \25181 );
not \U$16546 ( \25183 , \25182 );
not \U$16547 ( \25184 , \24911 );
or \U$16548 ( \25185 , \24034 , \25184 );
nand \U$16549 ( \25186 , \25180 , \25183 , \25185 );
and \U$16550 ( \25187 , \25186 , \22756 );
or \U$16551 ( \25188 , \25178 , \25187 );
and \U$16553 ( \25189 , \25188 , 1'b1 );
or \U$16555 ( \25190 , \25189 , 1'b0 );
buf \U$16556 ( \25191 , \25190 );
_DC r2552c_GF_IsGateDCbyConstraint ( \25192_nR2552c , \25191 , \21944 );
buf \U$16557 ( \25193 , \25192_nR2552c );
not \U$16558 ( \25194 , \24409 );
and \U$16559 ( \25195 , RIdb8e2e8_3873, \25194 );
not \U$16560 ( \25196 , RIdb8e2e8_3873);
or \U$16561 ( \25197 , \25196 , \24715 );
not \U$16562 ( \25198 , \24642 );
and \U$16563 ( \25199 , \22806 , \25198 );
not \U$16564 ( \25200 , \25199 );
not \U$16565 ( \25201 , \24647 );
or \U$16566 ( \25202 , \24052 , \25201 );
nand \U$16567 ( \25203 , \25197 , \25200 , \25202 );
and \U$16568 ( \25204 , \25203 , \24409 );
or \U$16569 ( \25205 , \25195 , \25204 );
and \U$16571 ( \25206 , \25205 , 1'b1 );
or \U$16573 ( \25207 , \25206 , 1'b0 );
buf \U$16574 ( \25208 , \25207 );
_DC r2552e_GF_IsGateDCbyConstraint ( \25209_nR2552e , \25208 , \21944 );
buf \U$16575 ( \25210 , \25209_nR2552e );
not \U$16576 ( \25211 , \22756 );
and \U$16577 ( \25212 , RIdb8b840_3874, \25211 );
not \U$16578 ( \25213 , RIdb8b840_3874);
or \U$16579 ( \25214 , \25213 , \24734 );
not \U$16580 ( \25215 , \24822 );
and \U$16581 ( \25216 , \22826 , \25215 );
not \U$16582 ( \25217 , \25216 );
not \U$16583 ( \25218 , \24911 );
or \U$16584 ( \25219 , \24070 , \25218 );
nand \U$16585 ( \25220 , \25214 , \25217 , \25219 );
and \U$16586 ( \25221 , \25220 , \22756 );
or \U$16587 ( \25222 , \25212 , \25221 );
and \U$16589 ( \25223 , \25222 , 1'b1 );
or \U$16591 ( \25224 , \25223 , 1'b0 );
buf \U$16592 ( \25225 , \25224 );
_DC r25530_GF_IsGateDCbyConstraint ( \25226_nR25530 , \25225 , \21944 );
buf \U$16593 ( \25227 , \25226_nR25530 );
not \U$16594 ( \25228 , \24117 );
and \U$16595 ( \25229 , RIdb890e0_3875, \25228 );
not \U$16596 ( \25230 , RIdb890e0_3875);
or \U$16597 ( \25231 , \25230 , \24734 );
not \U$16598 ( \25232 , \24736 );
and \U$16599 ( \25233 , \22846 , \25232 );
not \U$16600 ( \25234 , \25233 );
not \U$16601 ( \25235 , \24647 );
or \U$16602 ( \25236 , \24088 , \25235 );
nand \U$16603 ( \25237 , \25231 , \25234 , \25236 );
and \U$16604 ( \25238 , \25237 , \24117 );
or \U$16605 ( \25239 , \25229 , \25238 );
and \U$16607 ( \25240 , \25239 , 1'b1 );
or \U$16609 ( \25241 , \25240 , 1'b0 );
buf \U$16610 ( \25242 , \25241 );
_DC r25532_GF_IsGateDCbyConstraint ( \25243_nR25532 , \25242 , \21944 );
buf \U$16611 ( \25244 , \25243_nR25532 );
not \U$16612 ( \25245 , \24409 );
and \U$16613 ( \25246 , RIdb86cc8_3876, \25245 );
not \U$16614 ( \25247 , RIdb86cc8_3876);
or \U$16615 ( \25248 , \25247 , \24661 );
not \U$16616 ( \25249 , \24753 );
and \U$16617 ( \25250 , \22866 , \25249 );
not \U$16618 ( \25251 , \25250 );
not \U$16619 ( \25252 , \24911 );
or \U$16620 ( \25253 , \24106 , \25252 );
nand \U$16621 ( \25254 , \25248 , \25251 , \25253 );
and \U$16622 ( \25255 , \25254 , \24409 );
or \U$16623 ( \25256 , \25246 , \25255 );
and \U$16625 ( \25257 , \25256 , 1'b1 );
or \U$16627 ( \25258 , \25257 , 1'b0 );
buf \U$16628 ( \25259 , \25258 );
_DC r25534_GF_IsGateDCbyConstraint ( \25260_nR25534 , \25259 , \21944 );
buf \U$16629 ( \25261 , \25260_nR25534 );
not \U$16630 ( \25262 , \22756 );
and \U$16631 ( \25263 , RIdb84ec8_3877, \25262 );
not \U$16632 ( \25264 , RIdb84ec8_3877);
or \U$16633 ( \25265 , \25264 , \24661 );
not \U$16634 ( \25266 , \24642 );
and \U$16635 ( \25267 , \22886 , \25266 );
not \U$16636 ( \25268 , \25267 );
not \U$16637 ( \25269 , \24911 );
or \U$16638 ( \25270 , \24126 , \25269 );
nand \U$16639 ( \25271 , \25265 , \25268 , \25270 );
and \U$16640 ( \25272 , \25271 , \22756 );
or \U$16641 ( \25273 , \25263 , \25272 );
and \U$16643 ( \25274 , \25273 , 1'b1 );
or \U$16645 ( \25275 , \25274 , 1'b0 );
buf \U$16646 ( \25276 , \25275 );
_DC r25536_GF_IsGateDCbyConstraint ( \25277_nR25536 , \25276 , \21944 );
buf \U$16647 ( \25278 , \25277_nR25536 );
not \U$16648 ( \25279 , \24117 );
and \U$16649 ( \25280 , RIdb83410_3878, \25279 );
not \U$16650 ( \25281 , RIdb83410_3878);
or \U$16651 ( \25282 , \25281 , \24734 );
not \U$16652 ( \25283 , \24822 );
and \U$16653 ( \25284 , \22908 , \25283 );
not \U$16654 ( \25285 , \25284 );
not \U$16655 ( \25286 , \24911 );
or \U$16656 ( \25287 , \24144 , \25286 );
nand \U$16657 ( \25288 , \25282 , \25285 , \25287 );
and \U$16658 ( \25289 , \25288 , \24117 );
or \U$16659 ( \25290 , \25280 , \25289 );
and \U$16661 ( \25291 , \25290 , 1'b1 );
or \U$16663 ( \25292 , \25291 , 1'b0 );
buf \U$16664 ( \25293 , \25292 );
_DC r25538_GF_IsGateDCbyConstraint ( \25294_nR25538 , \25293 , \21944 );
buf \U$16665 ( \25295 , \25294_nR25538 );
not \U$16666 ( \25296 , \24409 );
and \U$16667 ( \25297 , RIdb81700_3879, \25296 );
not \U$16668 ( \25298 , RIdb81700_3879);
or \U$16669 ( \25299 , \25298 , \24715 );
not \U$16670 ( \25300 , \24698 );
and \U$16671 ( \25301 , \22928 , \25300 );
not \U$16672 ( \25302 , \25301 );
not \U$16673 ( \25303 , \24666 );
or \U$16674 ( \25304 , \24164 , \25303 );
nand \U$16675 ( \25305 , \25299 , \25302 , \25304 );
and \U$16676 ( \25306 , \25305 , \24409 );
or \U$16677 ( \25307 , \25297 , \25306 );
and \U$16679 ( \25308 , \25307 , 1'b1 );
or \U$16681 ( \25309 , \25308 , 1'b0 );
buf \U$16682 ( \25310 , \25309 );
_DC r2553a_GF_IsGateDCbyConstraint ( \25311_nR2553a , \25310 , \21944 );
buf \U$16683 ( \25312 , \25311_nR2553a );
not \U$16684 ( \25313 , \24117 );
and \U$16685 ( \25314 , RIdb7fa68_3880, \25313 );
not \U$16686 ( \25315 , RIdb7fa68_3880);
or \U$16687 ( \25316 , \25315 , \24803 );
not \U$16688 ( \25317 , \24736 );
and \U$16689 ( \25318 , \22948 , \25317 );
not \U$16690 ( \25319 , \25318 );
not \U$16691 ( \25320 , \24720 );
or \U$16692 ( \25321 , \24182 , \25320 );
nand \U$16693 ( \25322 , \25316 , \25319 , \25321 );
and \U$16694 ( \25323 , \25322 , \24117 );
or \U$16695 ( \25324 , \25314 , \25323 );
and \U$16697 ( \25325 , \25324 , 1'b1 );
or \U$16699 ( \25326 , \25325 , 1'b0 );
buf \U$16700 ( \25327 , \25326 );
_DC r2553c_GF_IsGateDCbyConstraint ( \25328_nR2553c , \25327 , \21944 );
buf \U$16701 ( \25329 , \25328_nR2553c );
not \U$16702 ( \25330 , \24117 );
and \U$16703 ( \25331 , RIdb7db78_3881, \25330 );
not \U$16704 ( \25332 , RIdb7db78_3881);
or \U$16705 ( \25333 , \25332 , \24803 );
not \U$16706 ( \25334 , \24736 );
and \U$16707 ( \25335 , \22968 , \25334 );
not \U$16708 ( \25336 , \25335 );
not \U$16709 ( \25337 , \24647 );
or \U$16710 ( \25338 , \24200 , \25337 );
nand \U$16711 ( \25339 , \25333 , \25336 , \25338 );
and \U$16712 ( \25340 , \25339 , \24117 );
or \U$16713 ( \25341 , \25331 , \25340 );
and \U$16715 ( \25342 , \25341 , 1'b1 );
or \U$16717 ( \25343 , \25342 , 1'b0 );
buf \U$16718 ( \25344 , \25343 );
_DC r25540_GF_IsGateDCbyConstraint ( \25345_nR25540 , \25344 , \21944 );
buf \U$16719 ( \25346 , \25345_nR25540 );
not \U$16720 ( \25347 , \24409 );
and \U$16721 ( \25348 , RIdb7bb98_3882, \25347 );
not \U$16722 ( \25349 , RIdb7bb98_3882);
or \U$16723 ( \25350 , \25349 , \24715 );
not \U$16724 ( \25351 , \24698 );
and \U$16725 ( \25352 , \22987 , \25351 );
not \U$16726 ( \25353 , \25352 );
not \U$16727 ( \25354 , \24720 );
or \U$16728 ( \25355 , \24218 , \25354 );
nand \U$16729 ( \25356 , \25350 , \25353 , \25355 );
and \U$16730 ( \25357 , \25356 , \24409 );
or \U$16731 ( \25358 , \25348 , \25357 );
and \U$16733 ( \25359 , \25358 , 1'b1 );
or \U$16735 ( \25360 , \25359 , 1'b0 );
buf \U$16736 ( \25361 , \25360 );
_DC r25542_GF_IsGateDCbyConstraint ( \25362_nR25542 , \25361 , \21944 );
buf \U$16737 ( \25363 , \25362_nR25542 );
not \U$16738 ( \25364 , \24117 );
and \U$16739 ( \25365 , RIdb79e10_3883, \25364 );
not \U$16740 ( \25366 , RIdb79e10_3883);
or \U$16741 ( \25367 , \25366 , \24661 );
not \U$16742 ( \25368 , \24753 );
and \U$16743 ( \25369 , \23006 , \25368 );
not \U$16744 ( \25370 , \25369 );
not \U$16745 ( \25371 , \24666 );
or \U$16746 ( \25372 , \24236 , \25371 );
nand \U$16747 ( \25373 , \25367 , \25370 , \25372 );
and \U$16748 ( \25374 , \25373 , \24117 );
or \U$16749 ( \25375 , \25365 , \25374 );
and \U$16751 ( \25376 , \25375 , 1'b1 );
or \U$16753 ( \25377 , \25376 , 1'b0 );
buf \U$16754 ( \25378 , \25377 );
_DC r25544_GF_IsGateDCbyConstraint ( \25379_nR25544 , \25378 , \21944 );
buf \U$16755 ( \25380 , \25379_nR25544 );
not \U$16756 ( \25381 , \24155 );
and \U$16757 ( \25382 , RIdb78268_3884, \25381 );
not \U$16758 ( \25383 , RIdb78268_3884);
or \U$16759 ( \25384 , \25383 , \24803 );
not \U$16760 ( \25385 , \24698 );
and \U$16761 ( \25386 , \23026 , \25385 );
not \U$16762 ( \25387 , \25386 );
not \U$16763 ( \25388 , \24720 );
or \U$16764 ( \25389 , \24254 , \25388 );
nand \U$16765 ( \25390 , \25384 , \25387 , \25389 );
and \U$16766 ( \25391 , \25390 , \24155 );
or \U$16767 ( \25392 , \25382 , \25391 );
and \U$16769 ( \25393 , \25392 , 1'b1 );
or \U$16771 ( \25394 , \25393 , 1'b0 );
buf \U$16772 ( \25395 , \25394 );
_DC r25546_GF_IsGateDCbyConstraint ( \25396_nR25546 , \25395 , \21944 );
buf \U$16773 ( \25397 , \25396_nR25546 );
not \U$16774 ( \25398 , \24155 );
and \U$16775 ( \25399 , RIdb76828_3885, \25398 );
not \U$16776 ( \25400 , RIdb76828_3885);
or \U$16777 ( \25401 , \25400 , \24715 );
not \U$16778 ( \25402 , \24736 );
and \U$16779 ( \25403 , \23048 , \25402 );
not \U$16780 ( \25404 , \25403 );
not \U$16781 ( \25405 , \24647 );
or \U$16782 ( \25406 , \24272 , \25405 );
nand \U$16783 ( \25407 , \25401 , \25404 , \25406 );
and \U$16784 ( \25408 , \25407 , \24155 );
or \U$16785 ( \25409 , \25399 , \25408 );
and \U$16787 ( \25410 , \25409 , 1'b1 );
or \U$16789 ( \25411 , \25410 , 1'b0 );
buf \U$16790 ( \25412 , \25411 );
_DC r25548_GF_IsGateDCbyConstraint ( \25413_nR25548 , \25412 , \21944 );
buf \U$16791 ( \25414 , \25413_nR25548 );
not \U$16792 ( \25415 , \22756 );
and \U$16793 ( \25416 , RIdb746e0_3886, \25415 );
not \U$16794 ( \25417 , RIdb746e0_3886);
or \U$16795 ( \25418 , \25417 , \24640 );
not \U$16796 ( \25419 , \24753 );
and \U$16797 ( \25420 , \23068 , \25419 );
not \U$16798 ( \25421 , \25420 );
not \U$16799 ( \25422 , \24720 );
or \U$16800 ( \25423 , \24290 , \25422 );
nand \U$16801 ( \25424 , \25418 , \25421 , \25423 );
and \U$16802 ( \25425 , \25424 , \22756 );
or \U$16803 ( \25426 , \25416 , \25425 );
and \U$16805 ( \25427 , \25426 , 1'b1 );
or \U$16807 ( \25428 , \25427 , 1'b0 );
buf \U$16808 ( \25429 , \25428 );
_DC r2554a_GF_IsGateDCbyConstraint ( \25430_nR2554a , \25429 , \21944 );
buf \U$16809 ( \25431 , \25430_nR2554a );
not \U$16810 ( \25432 , \22195 );
and \U$16811 ( \25433 , RIdda9490_3887, \25432 );
not \U$16812 ( \25434 , RIdda9490_3887);
or \U$16813 ( \25435 , \25434 , \24715 );
not \U$16814 ( \25436 , \24736 );
and \U$16815 ( \25437 , \23088 , \25436 );
not \U$16816 ( \25438 , \25437 );
not \U$16817 ( \25439 , \24647 );
or \U$16818 ( \25440 , \24308 , \25439 );
nand \U$16819 ( \25441 , \25435 , \25438 , \25440 );
and \U$16820 ( \25442 , \25441 , \22195 );
or \U$16821 ( \25443 , \25433 , \25442 );
and \U$16823 ( \25444 , \25443 , 1'b1 );
or \U$16825 ( \25445 , \25444 , 1'b0 );
buf \U$16826 ( \25446 , \25445 );
_DC r2554c_GF_IsGateDCbyConstraint ( \25447_nR2554c , \25446 , \21944 );
buf \U$16827 ( \25448 , \25447_nR2554c );
buf \U$16828 ( \25449 , \23038 );
not \U$16829 ( \25450 , \25449 );
and \U$16830 ( \25451 , RIdda9c88_3888, \25450 );
not \U$16831 ( \25452 , RIdda9c88_3888);
or \U$16832 ( \25453 , \25452 , \24734 );
not \U$16833 ( \25454 , \24753 );
and \U$16834 ( \25455 , \23108 , \25454 );
not \U$16835 ( \25456 , \25455 );
not \U$16836 ( \25457 , \24911 );
or \U$16837 ( \25458 , \24326 , \25457 );
nand \U$16838 ( \25459 , \25453 , \25456 , \25458 );
and \U$16839 ( \25460 , \25459 , \25449 );
or \U$16840 ( \25461 , \25451 , \25460 );
and \U$16842 ( \25462 , \25461 , 1'b1 );
or \U$16844 ( \25463 , \25462 , 1'b0 );
buf \U$16845 ( \25464 , \25463 );
_DC r2554e_GF_IsGateDCbyConstraint ( \25465_nR2554e , \25464 , \21944 );
buf \U$16846 ( \25466 , \25465_nR2554e );
not \U$16847 ( \25467 , \23038 );
and \U$16848 ( \25468 , RIddaa480_3889, \25467 );
not \U$16849 ( \25469 , RIddaa480_3889);
or \U$16850 ( \25470 , \25469 , \24640 );
not \U$16851 ( \25471 , \24698 );
and \U$16852 ( \25472 , \23128 , \25471 );
not \U$16853 ( \25473 , \25472 );
not \U$16854 ( \25474 , \24647 );
or \U$16855 ( \25475 , \24344 , \25474 );
nand \U$16856 ( \25476 , \25470 , \25473 , \25475 );
and \U$16857 ( \25477 , \25476 , \23038 );
or \U$16858 ( \25478 , \25468 , \25477 );
and \U$16860 ( \25479 , \25478 , 1'b1 );
or \U$16862 ( \25480 , \25479 , 1'b0 );
buf \U$16863 ( \25481 , \25480 );
_DC r25550_GF_IsGateDCbyConstraint ( \25482_nR25550 , \25481 , \21944 );
buf \U$16864 ( \25483 , \25482_nR25550 );
not \U$16865 ( \25484 , \22756 );
and \U$16866 ( \25485 , RIddaac78_3890, \25484 );
not \U$16867 ( \25486 , RIddaac78_3890);
or \U$16868 ( \25487 , \25486 , \24640 );
not \U$16869 ( \25488 , \24736 );
and \U$16870 ( \25489 , \23148 , \25488 );
not \U$16871 ( \25490 , \25489 );
not \U$16872 ( \25491 , \24666 );
or \U$16873 ( \25492 , \24362 , \25491 );
nand \U$16874 ( \25493 , \25487 , \25490 , \25492 );
and \U$16875 ( \25494 , \25493 , \22756 );
or \U$16876 ( \25495 , \25485 , \25494 );
and \U$16878 ( \25496 , \25495 , 1'b1 );
or \U$16880 ( \25497 , \25496 , 1'b0 );
buf \U$16881 ( \25498 , \25497 );
_DC r25552_GF_IsGateDCbyConstraint ( \25499_nR25552 , \25498 , \21944 );
buf \U$16882 ( \25500 , \25499_nR25552 );
not \U$16883 ( \25501 , \25449 );
and \U$16884 ( \25502 , RIddab470_3891, \25501 );
not \U$16885 ( \25503 , RIddab470_3891);
or \U$16886 ( \25504 , \25503 , \24734 );
not \U$16887 ( \25505 , \24642 );
and \U$16888 ( \25506 , \23168 , \25505 );
not \U$16889 ( \25507 , \25506 );
not \U$16890 ( \25508 , \24720 );
or \U$16891 ( \25509 , \24380 , \25508 );
nand \U$16892 ( \25510 , \25504 , \25507 , \25509 );
and \U$16893 ( \25511 , \25510 , \25449 );
or \U$16894 ( \25512 , \25502 , \25511 );
and \U$16896 ( \25513 , \25512 , 1'b1 );
or \U$16898 ( \25514 , \25513 , 1'b0 );
buf \U$16899 ( \25515 , \25514 );
_DC r25556_GF_IsGateDCbyConstraint ( \25516_nR25556 , \25515 , \21944 );
buf \U$16900 ( \25517 , \25516_nR25556 );
not \U$16901 ( \25518 , \22104 );
and \U$16902 ( \25519 , RIddabc68_3892, \25518 );
not \U$16903 ( \25520 , RIddabc68_3892);
or \U$16904 ( \25521 , \25520 , \24715 );
not \U$16905 ( \25522 , \24822 );
and \U$16906 ( \25523 , \23187 , \25522 );
not \U$16907 ( \25524 , \25523 );
not \U$16908 ( \25525 , \24666 );
or \U$16909 ( \25526 , \24398 , \25525 );
nand \U$16910 ( \25527 , \25521 , \25524 , \25526 );
and \U$16911 ( \25528 , \25527 , \22104 );
or \U$16912 ( \25529 , \25519 , \25528 );
and \U$16914 ( \25530 , \25529 , 1'b1 );
or \U$16916 ( \25531 , \25530 , 1'b0 );
buf \U$16917 ( \25532 , \25531 );
_DC r25558_GF_IsGateDCbyConstraint ( \25533_nR25558 , \25532 , \21944 );
buf \U$16918 ( \25534 , \25533_nR25558 );
not \U$16919 ( \25535 , \22756 );
and \U$16920 ( \25536 , RIddac460_3893, \25535 );
not \U$16921 ( \25537 , RIddac460_3893);
or \U$16922 ( \25538 , \25537 , \24734 );
not \U$16923 ( \25539 , \24736 );
and \U$16924 ( \25540 , \23207 , \25539 );
not \U$16925 ( \25541 , \25540 );
not \U$16926 ( \25542 , \24666 );
or \U$16927 ( \25543 , \24417 , \25542 );
nand \U$16928 ( \25544 , \25538 , \25541 , \25543 );
and \U$16929 ( \25545 , \25544 , \22756 );
or \U$16930 ( \25546 , \25536 , \25545 );
and \U$16932 ( \25547 , \25546 , 1'b1 );
or \U$16934 ( \25548 , \25547 , 1'b0 );
buf \U$16935 ( \25549 , \25548 );
_DC r2555a_GF_IsGateDCbyConstraint ( \25550_nR2555a , \25549 , \21944 );
buf \U$16936 ( \25551 , \25550_nR2555a );
not \U$16937 ( \25552 , \25449 );
and \U$16938 ( \25553 , RIddacc58_3894, \25552 );
not \U$16939 ( \25554 , RIddacc58_3894);
or \U$16940 ( \25555 , \25554 , \24640 );
not \U$16941 ( \25556 , \24642 );
and \U$16942 ( \25557 , \23227 , \25556 );
not \U$16943 ( \25558 , \25557 );
not \U$16944 ( \25559 , \24720 );
or \U$16945 ( \25560 , \24435 , \25559 );
nand \U$16946 ( \25561 , \25555 , \25558 , \25560 );
and \U$16947 ( \25562 , \25561 , \25449 );
or \U$16948 ( \25563 , \25553 , \25562 );
and \U$16950 ( \25564 , \25563 , 1'b1 );
or \U$16952 ( \25565 , \25564 , 1'b0 );
buf \U$16953 ( \25566 , \25565 );
_DC r2555c_GF_IsGateDCbyConstraint ( \25567_nR2555c , \25566 , \21944 );
buf \U$16954 ( \25568 , \25567_nR2555c );
not \U$16955 ( \25569 , \22195 );
and \U$16956 ( \25570 , RIddad450_3895, \25569 );
not \U$16957 ( \25571 , RIddad450_3895);
or \U$16958 ( \25572 , \25571 , \24661 );
not \U$16959 ( \25573 , \24822 );
and \U$16960 ( \25574 , \23247 , \25573 );
not \U$16961 ( \25575 , \25574 );
not \U$16962 ( \25576 , \24666 );
or \U$16963 ( \25577 , \24453 , \25576 );
nand \U$16964 ( \25578 , \25572 , \25575 , \25577 );
and \U$16965 ( \25579 , \25578 , \22195 );
or \U$16966 ( \25580 , \25570 , \25579 );
and \U$16968 ( \25581 , \25580 , 1'b1 );
or \U$16970 ( \25582 , \25581 , 1'b0 );
buf \U$16971 ( \25583 , \25582 );
_DC r2555e_GF_IsGateDCbyConstraint ( \25584_nR2555e , \25583 , \21944 );
buf \U$16972 ( \25585 , \25584_nR2555e );
not \U$16973 ( \25586 , \23038 );
and \U$16974 ( \25587 , RIddadc48_3896, \25586 );
not \U$16975 ( \25588 , RIddadc48_3896);
or \U$16976 ( \25589 , \25588 , \24734 );
not \U$16977 ( \25590 , \24642 );
and \U$16978 ( \25591 , \23267 , \25590 );
not \U$16979 ( \25592 , \25591 );
not \U$16980 ( \25593 , \24720 );
or \U$16981 ( \25594 , \24471 , \25593 );
nand \U$16982 ( \25595 , \25589 , \25592 , \25594 );
and \U$16983 ( \25596 , \25595 , \23038 );
or \U$16984 ( \25597 , \25587 , \25596 );
and \U$16986 ( \25598 , \25597 , 1'b1 );
or \U$16988 ( \25599 , \25598 , 1'b0 );
buf \U$16989 ( \25600 , \25599 );
_DC r25560_GF_IsGateDCbyConstraint ( \25601_nR25560 , \25600 , \21944 );
buf \U$16990 ( \25602 , \25601_nR25560 );
not \U$16991 ( \25603 , \25449 );
and \U$16992 ( \25604 , RIddae440_3897, \25603 );
not \U$16993 ( \25605 , RIddae440_3897);
or \U$16994 ( \25606 , \25605 , \24803 );
not \U$16995 ( \25607 , \24753 );
and \U$16996 ( \25608 , \23287 , \25607 );
not \U$16997 ( \25609 , \25608 );
not \U$16998 ( \25610 , \24720 );
or \U$16999 ( \25611 , \24489 , \25610 );
nand \U$17000 ( \25612 , \25606 , \25609 , \25611 );
and \U$17001 ( \25613 , \25612 , \25449 );
or \U$17002 ( \25614 , \25604 , \25613 );
and \U$17004 ( \25615 , \25614 , 1'b1 );
or \U$17006 ( \25616 , \25615 , 1'b0 );
buf \U$17007 ( \25617 , \25616 );
_DC r25562_GF_IsGateDCbyConstraint ( \25618_nR25562 , \25617 , \21944 );
buf \U$17008 ( \25619 , \25618_nR25562 );
not \U$17009 ( \25620 , \24155 );
and \U$17010 ( \25621 , RIddaec38_3898, \25620 );
not \U$17011 ( \25622 , RIddaec38_3898);
or \U$17012 ( \25623 , \25622 , \24715 );
not \U$17013 ( \25624 , \24822 );
and \U$17014 ( \25625 , \23306 , \25624 );
not \U$17015 ( \25626 , \25625 );
not \U$17016 ( \25627 , \24666 );
or \U$17017 ( \25628 , \24507 , \25627 );
nand \U$17018 ( \25629 , \25623 , \25626 , \25628 );
and \U$17019 ( \25630 , \25629 , \24155 );
or \U$17020 ( \25631 , \25621 , \25630 );
and \U$17022 ( \25632 , \25631 , 1'b1 );
or \U$17024 ( \25633 , \25632 , 1'b0 );
buf \U$17025 ( \25634 , \25633 );
_DC r25564_GF_IsGateDCbyConstraint ( \25635_nR25564 , \25634 , \21944 );
buf \U$17026 ( \25636 , \25635_nR25564 );
buf \U$17027 ( \25637 , \24117 );
not \U$17028 ( \25638 , \25637 );
and \U$17029 ( \25639 , RIddaf430_3899, \25638 );
not \U$17030 ( \25640 , RIddaf430_3899);
or \U$17031 ( \25641 , \25640 , \24661 );
not \U$17032 ( \25642 , \24698 );
and \U$17033 ( \25643 , \23326 , \25642 );
not \U$17034 ( \25644 , \25643 );
not \U$17035 ( \25645 , \24666 );
or \U$17036 ( \25646 , \24525 , \25645 );
nand \U$17037 ( \25647 , \25641 , \25644 , \25646 );
and \U$17038 ( \25648 , \25647 , \25637 );
or \U$17039 ( \25649 , \25639 , \25648 );
and \U$17041 ( \25650 , \25649 , 1'b1 );
or \U$17043 ( \25651 , \25650 , 1'b0 );
buf \U$17044 ( \25652 , \25651 );
_DC r25566_GF_IsGateDCbyConstraint ( \25653_nR25566 , \25652 , \21944 );
buf \U$17045 ( \25654 , \25653_nR25566 );
not \U$17046 ( \25655 , \25449 );
and \U$17047 ( \25656 , RIddafc28_3900, \25655 );
not \U$17048 ( \25657 , RIddafc28_3900);
or \U$17049 ( \25658 , \25657 , \24734 );
not \U$17050 ( \25659 , \24631 );
and \U$17051 ( \25660 , \23346 , \25659 );
not \U$17052 ( \25661 , \25660 );
not \U$17053 ( \25662 , \24720 );
or \U$17054 ( \25663 , \24543 , \25662 );
nand \U$17055 ( \25664 , \25658 , \25661 , \25663 );
and \U$17056 ( \25665 , \25664 , \25449 );
or \U$17057 ( \25666 , \25656 , \25665 );
and \U$17059 ( \25667 , \25666 , 1'b1 );
or \U$17061 ( \25668 , \25667 , 1'b0 );
buf \U$17062 ( \25669 , \25668 );
_DC r25568_GF_IsGateDCbyConstraint ( \25670_nR25568 , \25669 , \21944 );
buf \U$17063 ( \25671 , \25670_nR25568 );
not \U$17064 ( \25672 , \22756 );
and \U$17065 ( \25673 , RIddb0420_3901, \25672 );
not \U$17066 ( \25674 , RIddb0420_3901);
or \U$17067 ( \25675 , \25674 , \24640 );
not \U$17068 ( \25676 , \24753 );
and \U$17069 ( \25677 , \23367 , \25676 );
not \U$17070 ( \25678 , \25677 );
not \U$17071 ( \25679 , \24720 );
or \U$17072 ( \25680 , \24561 , \25679 );
nand \U$17073 ( \25681 , \25675 , \25678 , \25680 );
and \U$17074 ( \25682 , \25681 , \22756 );
or \U$17075 ( \25683 , \25673 , \25682 );
and \U$17077 ( \25684 , \25683 , 1'b1 );
or \U$17079 ( \25685 , \25684 , 1'b0 );
buf \U$17080 ( \25686 , \25685 );
_DC r2556c_GF_IsGateDCbyConstraint ( \25687_nR2556c , \25686 , \21944 );
buf \U$17081 ( \25688 , \25687_nR2556c );
not \U$17082 ( \25689 , \25637 );
and \U$17083 ( \25690 , RIddb0c18_3902, \25689 );
not \U$17084 ( \25691 , RIddb0c18_3902);
or \U$17085 ( \25692 , \25691 , \24803 );
not \U$17086 ( \25693 , \24698 );
and \U$17087 ( \25694 , \23387 , \25693 );
not \U$17088 ( \25695 , \25694 );
not \U$17089 ( \25696 , \24720 );
or \U$17090 ( \25697 , \24579 , \25696 );
nand \U$17091 ( \25698 , \25692 , \25695 , \25697 );
and \U$17092 ( \25699 , \25698 , \25637 );
or \U$17093 ( \25700 , \25690 , \25699 );
and \U$17095 ( \25701 , \25700 , 1'b1 );
or \U$17097 ( \25702 , \25701 , 1'b0 );
buf \U$17098 ( \25703 , \25702 );
_DC r2556e_GF_IsGateDCbyConstraint ( \25704_nR2556e , \25703 , \21944 );
buf \U$17099 ( \25705 , \25704_nR2556e );
not \U$17100 ( \25706 , \25449 );
and \U$17101 ( \25707 , RIddb1410_3903, \25706 );
not \U$17102 ( \25708 , RIddb1410_3903);
or \U$17103 ( \25709 , \25708 , \24661 );
not \U$17104 ( \25710 , \24736 );
and \U$17105 ( \25711 , \23407 , \25710 );
not \U$17106 ( \25712 , \25711 );
not \U$17107 ( \25713 , \24666 );
or \U$17108 ( \25714 , \24597 , \25713 );
nand \U$17109 ( \25715 , \25709 , \25712 , \25714 );
and \U$17110 ( \25716 , \25715 , \25449 );
or \U$17111 ( \25717 , \25707 , \25716 );
and \U$17113 ( \25718 , \25717 , 1'b1 );
or \U$17115 ( \25719 , \25718 , 1'b0 );
buf \U$17116 ( \25720 , \25719 );
_DC r25570_GF_IsGateDCbyConstraint ( \25721_nR25570 , \25720 , \21944 );
buf \U$17117 ( \25722 , \25721_nR25570 );
not \U$17118 ( \25723 , \22195 );
and \U$17119 ( \25724 , RIddb1c08_3904, \25723 );
not \U$17120 ( \25725 , RIddb1c08_3904);
or \U$17121 ( \25726 , \25725 , \24803 );
not \U$17122 ( \25727 , \24736 );
and \U$17123 ( \25728 , \23427 , \25727 );
not \U$17124 ( \25729 , \25728 );
not \U$17125 ( \25730 , \24666 );
or \U$17126 ( \25731 , \24615 , \25730 );
nand \U$17127 ( \25732 , \25726 , \25729 , \25731 );
and \U$17128 ( \25733 , \25732 , \22195 );
or \U$17129 ( \25734 , \25724 , \25733 );
and \U$17131 ( \25735 , \25734 , 1'b1 );
or \U$17133 ( \25736 , \25735 , 1'b0 );
buf \U$17134 ( \25737 , \25736 );
_DC r25572_GF_IsGateDCbyConstraint ( \25738_nR25572 , \25737 , \21944 );
buf \U$17135 ( \25739 , \25738_nR25572 );
not \U$17136 ( \25740 , \25637 );
and \U$17137 ( \25741 , RIddb2400_3905, \25740 );
not \U$17138 ( \25742 , RIddb2400_3905);
nand \U$17139 ( \25743 , \22121 , \22117 );
not \U$17140 ( \25744 , \22123 );
or \U$17141 ( \25745 , \25743 , \25744 );
not \U$17142 ( \25746 , \25745 );
nand \U$17143 ( \25747 , \22111 , \22110 );
not \U$17144 ( \25748 , \25747 );
nand \U$17145 ( \25749 , \22102 , \25748 );
not \U$17146 ( \25750 , \25749 );
or \U$17147 ( \25751 , \25746 , \25750 );
buf \U$17148 ( \25752 , \25751 );
or \U$17149 ( \25753 , \25742 , \25752 );
not \U$17150 ( \25754 , \25749 );
buf \U$17151 ( \25755 , \25754 );
nand \U$17152 ( \25756 , \22132 , \25755 );
buf \U$17153 ( \25757 , \25746 );
nand \U$17154 ( \25758 , \22135 , \25757 );
nand \U$17155 ( \25759 , \25753 , \25756 , \25758 );
and \U$17156 ( \25760 , \25759 , \25637 );
or \U$17157 ( \25761 , \25741 , \25760 );
and \U$17159 ( \25762 , \25761 , 1'b1 );
or \U$17161 ( \25763 , \25762 , 1'b0 );
buf \U$17162 ( \25764 , \25763 );
_DC r2557c_GF_IsGateDCbyConstraint ( \25765_nR2557c , \25764 , \21944 );
buf \U$17163 ( \25766 , \25765_nR2557c );
not \U$17164 ( \25767 , \25449 );
and \U$17165 ( \25768 , RIddb2bf8_3906, \25767 );
not \U$17166 ( \25769 , RIddb2bf8_3906);
buf \U$17167 ( \25770 , \25751 );
or \U$17168 ( \25771 , \25769 , \25770 );
buf \U$17169 ( \25772 , \25754 );
nand \U$17170 ( \25773 , \22159 , \25772 );
nand \U$17171 ( \25774 , \22162 , \25757 );
nand \U$17172 ( \25775 , \25771 , \25773 , \25774 );
and \U$17173 ( \25776 , \25775 , \25449 );
or \U$17174 ( \25777 , \25768 , \25776 );
and \U$17176 ( \25778 , \25777 , 1'b1 );
or \U$17178 ( \25779 , \25778 , 1'b0 );
buf \U$17179 ( \25780 , \25779 );
_DC r25592_GF_IsGateDCbyConstraint ( \25781_nR25592 , \25780 , \21944 );
buf \U$17180 ( \25782 , \25781_nR25592 );
not \U$17181 ( \25783 , \22104 );
and \U$17182 ( \25784 , RIddb33f0_3907, \25783 );
not \U$17183 ( \25785 , RIddb33f0_3907);
buf \U$17184 ( \25786 , \25751 );
or \U$17185 ( \25787 , \25785 , \25786 );
buf \U$17186 ( \25788 , \25754 );
nand \U$17187 ( \25789 , \22180 , \25788 );
buf \U$17188 ( \25790 , \25746 );
nand \U$17189 ( \25791 , \22183 , \25790 );
nand \U$17190 ( \25792 , \25787 , \25789 , \25791 );
and \U$17191 ( \25793 , \25792 , \22104 );
or \U$17192 ( \25794 , \25784 , \25793 );
and \U$17194 ( \25795 , \25794 , 1'b1 );
or \U$17196 ( \25796 , \25795 , 1'b0 );
buf \U$17197 ( \25797 , \25796 );
_DC r255a8_GF_IsGateDCbyConstraint ( \25798_nR255a8 , \25797 , \21944 );
buf \U$17198 ( \25799 , \25798_nR255a8 );
not \U$17199 ( \25800 , \25637 );
and \U$17200 ( \25801 , RIddb3be8_3908, \25800 );
not \U$17201 ( \25802 , RIddb3be8_3908);
buf \U$17202 ( \25803 , \25751 );
or \U$17203 ( \25804 , \25802 , \25803 );
nand \U$17204 ( \25805 , \22203 , \25755 );
buf \U$17205 ( \25806 , \25746 );
nand \U$17206 ( \25807 , \22206 , \25806 );
nand \U$17207 ( \25808 , \25804 , \25805 , \25807 );
and \U$17208 ( \25809 , \25808 , \25637 );
or \U$17209 ( \25810 , \25801 , \25809 );
and \U$17211 ( \25811 , \25810 , 1'b1 );
or \U$17213 ( \25812 , \25811 , 1'b0 );
buf \U$17214 ( \25813 , \25812 );
_DC r255be_GF_IsGateDCbyConstraint ( \25814_nR255be , \25813 , \21944 );
buf \U$17215 ( \25815 , \25814_nR255be );
not \U$17216 ( \25816 , \25449 );
and \U$17217 ( \25817 , RIddb43e0_3909, \25816 );
not \U$17218 ( \25818 , RIddb43e0_3909);
or \U$17219 ( \25819 , \25818 , \25752 );
nand \U$17220 ( \25820 , \22224 , \25788 );
nand \U$17221 ( \25821 , \22227 , \25790 );
nand \U$17222 ( \25822 , \25819 , \25820 , \25821 );
and \U$17223 ( \25823 , \25822 , \25449 );
or \U$17224 ( \25824 , \25817 , \25823 );
and \U$17226 ( \25825 , \25824 , 1'b1 );
or \U$17228 ( \25826 , \25825 , 1'b0 );
buf \U$17229 ( \25827 , \25826 );
_DC r255d4_GF_IsGateDCbyConstraint ( \25828_nR255d4 , \25827 , \21944 );
buf \U$17230 ( \25829 , \25828_nR255d4 );
not \U$17231 ( \25830 , \24117 );
and \U$17232 ( \25831 , RIddb4bd8_3910, \25830 );
not \U$17233 ( \25832 , RIddb4bd8_3910);
or \U$17234 ( \25833 , \25832 , \25770 );
nand \U$17235 ( \25834 , \22246 , \25788 );
buf \U$17236 ( \25835 , \25746 );
nand \U$17237 ( \25836 , \22249 , \25835 );
nand \U$17238 ( \25837 , \25833 , \25834 , \25836 );
and \U$17239 ( \25838 , \25837 , \24117 );
or \U$17240 ( \25839 , \25831 , \25838 );
and \U$17242 ( \25840 , \25839 , 1'b1 );
or \U$17244 ( \25841 , \25840 , 1'b0 );
buf \U$17245 ( \25842 , \25841 );
_DC r255ea_GF_IsGateDCbyConstraint ( \25843_nR255ea , \25842 , \21944 );
buf \U$17246 ( \25844 , \25843_nR255ea );
not \U$17247 ( \25845 , \25637 );
and \U$17248 ( \25846 , RIddb53d0_3911, \25845 );
not \U$17249 ( \25847 , RIddb53d0_3911);
or \U$17250 ( \25848 , \25847 , \25786 );
nand \U$17251 ( \25849 , \22272 , \25772 );
nand \U$17252 ( \25850 , \22275 , \25757 );
nand \U$17253 ( \25851 , \25848 , \25849 , \25850 );
and \U$17254 ( \25852 , \25851 , \25637 );
or \U$17255 ( \25853 , \25846 , \25852 );
and \U$17257 ( \25854 , \25853 , 1'b1 );
or \U$17259 ( \25855 , \25854 , 1'b0 );
buf \U$17260 ( \25856 , \25855 );
_DC r255f4_GF_IsGateDCbyConstraint ( \25857_nR255f4 , \25856 , \21944 );
buf \U$17261 ( \25858 , \25857_nR255f4 );
not \U$17262 ( \25859 , \25449 );
and \U$17263 ( \25860 , RIddb5bc8_3912, \25859 );
not \U$17264 ( \25861 , RIddb5bc8_3912);
or \U$17265 ( \25862 , \25861 , \25770 );
nand \U$17266 ( \25863 , \22292 , \25755 );
nand \U$17267 ( \25864 , \22295 , \25757 );
nand \U$17268 ( \25865 , \25862 , \25863 , \25864 );
and \U$17269 ( \25866 , \25865 , \25449 );
or \U$17270 ( \25867 , \25860 , \25866 );
and \U$17272 ( \25868 , \25867 , 1'b1 );
or \U$17274 ( \25869 , \25868 , 1'b0 );
buf \U$17275 ( \25870 , \25869 );
_DC r255f6_GF_IsGateDCbyConstraint ( \25871_nR255f6 , \25870 , \21944 );
buf \U$17276 ( \25872 , \25871_nR255f6 );
not \U$17277 ( \25873 , \23038 );
and \U$17278 ( \25874 , RIddb63c0_3913, \25873 );
not \U$17279 ( \25875 , RIddb63c0_3913);
or \U$17280 ( \25876 , \25875 , \25752 );
nand \U$17281 ( \25877 , \22314 , \25754 );
nand \U$17282 ( \25878 , \22317 , \25806 );
nand \U$17283 ( \25879 , \25876 , \25877 , \25878 );
and \U$17284 ( \25880 , \25879 , \23038 );
or \U$17285 ( \25881 , \25874 , \25880 );
and \U$17287 ( \25882 , \25881 , 1'b1 );
or \U$17289 ( \25883 , \25882 , 1'b0 );
buf \U$17290 ( \25884 , \25883 );
_DC r255f8_GF_IsGateDCbyConstraint ( \25885_nR255f8 , \25884 , \21944 );
buf \U$17291 ( \25886 , \25885_nR255f8 );
not \U$17292 ( \25887 , \25637 );
and \U$17293 ( \25888 , RIddb6bb8_3914, \25887 );
not \U$17294 ( \25889 , RIddb6bb8_3914);
buf \U$17295 ( \25890 , \25751 );
or \U$17296 ( \25891 , \25889 , \25890 );
nand \U$17297 ( \25892 , \22335 , \25788 );
nand \U$17298 ( \25893 , \22338 , \25790 );
nand \U$17299 ( \25894 , \25891 , \25892 , \25893 );
and \U$17300 ( \25895 , \25894 , \25637 );
or \U$17301 ( \25896 , \25888 , \25895 );
and \U$17303 ( \25897 , \25896 , 1'b1 );
or \U$17305 ( \25898 , \25897 , 1'b0 );
buf \U$17306 ( \25899 , \25898 );
_DC r255fa_GF_IsGateDCbyConstraint ( \25900_nR255fa , \25899 , \21944 );
buf \U$17307 ( \25901 , \25900_nR255fa );
not \U$17308 ( \25902 , \25449 );
and \U$17309 ( \25903 , RIddb73b0_3915, \25902 );
not \U$17310 ( \25904 , RIddb73b0_3915);
or \U$17311 ( \25905 , \25904 , \25890 );
nand \U$17312 ( \25906 , \22357 , \25788 );
nand \U$17313 ( \25907 , \22360 , \25835 );
nand \U$17314 ( \25908 , \25905 , \25906 , \25907 );
and \U$17315 ( \25909 , \25908 , \25449 );
or \U$17316 ( \25910 , \25903 , \25909 );
and \U$17318 ( \25911 , \25910 , 1'b1 );
or \U$17320 ( \25912 , \25911 , 1'b0 );
buf \U$17321 ( \25913 , \25912 );
_DC r2557e_GF_IsGateDCbyConstraint ( \25914_nR2557e , \25913 , \21944 );
buf \U$17322 ( \25915 , \25914_nR2557e );
not \U$17323 ( \25916 , \24117 );
and \U$17324 ( \25917 , RIddb7ba8_3916, \25916 );
not \U$17325 ( \25918 , RIddb7ba8_3916);
or \U$17326 ( \25919 , \25918 , \25803 );
nand \U$17327 ( \25920 , \22377 , \25788 );
nand \U$17328 ( \25921 , \22380 , \25790 );
nand \U$17329 ( \25922 , \25919 , \25920 , \25921 );
and \U$17330 ( \25923 , \25922 , \24117 );
or \U$17331 ( \25924 , \25917 , \25923 );
and \U$17333 ( \25925 , \25924 , 1'b1 );
or \U$17335 ( \25926 , \25925 , 1'b0 );
buf \U$17336 ( \25927 , \25926 );
_DC r25580_GF_IsGateDCbyConstraint ( \25928_nR25580 , \25927 , \21944 );
buf \U$17337 ( \25929 , \25928_nR25580 );
not \U$17338 ( \25930 , \25637 );
and \U$17339 ( \25931 , RIddb83a0_3917, \25930 );
not \U$17340 ( \25932 , RIddb83a0_3917);
or \U$17341 ( \25933 , \25932 , \25786 );
nand \U$17342 ( \25934 , \22398 , \25772 );
nand \U$17343 ( \25935 , \22401 , \25835 );
nand \U$17344 ( \25936 , \25933 , \25934 , \25935 );
and \U$17345 ( \25937 , \25936 , \25637 );
or \U$17346 ( \25938 , \25931 , \25937 );
and \U$17348 ( \25939 , \25938 , 1'b1 );
or \U$17350 ( \25940 , \25939 , 1'b0 );
buf \U$17351 ( \25941 , \25940 );
_DC r25582_GF_IsGateDCbyConstraint ( \25942_nR25582 , \25941 , \21944 );
buf \U$17352 ( \25943 , \25942_nR25582 );
not \U$17353 ( \25944 , \25449 );
and \U$17354 ( \25945 , RIddb8b98_3918, \25944 );
not \U$17355 ( \25946 , RIddb8b98_3918);
or \U$17356 ( \25947 , \25946 , \25803 );
nand \U$17357 ( \25948 , \22418 , \25788 );
nand \U$17358 ( \25949 , \22421 , \25806 );
nand \U$17359 ( \25950 , \25947 , \25948 , \25949 );
and \U$17360 ( \25951 , \25950 , \25449 );
or \U$17361 ( \25952 , \25945 , \25951 );
and \U$17363 ( \25953 , \25952 , 1'b1 );
or \U$17365 ( \25954 , \25953 , 1'b0 );
buf \U$17366 ( \25955 , \25954 );
_DC r25584_GF_IsGateDCbyConstraint ( \25956_nR25584 , \25955 , \21944 );
buf \U$17367 ( \25957 , \25956_nR25584 );
not \U$17368 ( \25958 , \24155 );
and \U$17369 ( \25959 , RIddb9390_3919, \25958 );
not \U$17370 ( \25960 , RIddb9390_3919);
or \U$17371 ( \25961 , \25960 , \25770 );
nand \U$17372 ( \25962 , \22438 , \25755 );
nand \U$17373 ( \25963 , \22441 , \25790 );
nand \U$17374 ( \25964 , \25961 , \25962 , \25963 );
and \U$17375 ( \25965 , \25964 , \24155 );
or \U$17376 ( \25966 , \25959 , \25965 );
and \U$17378 ( \25967 , \25966 , 1'b1 );
or \U$17380 ( \25968 , \25967 , 1'b0 );
buf \U$17381 ( \25969 , \25968 );
_DC r25586_GF_IsGateDCbyConstraint ( \25970_nR25586 , \25969 , \21944 );
buf \U$17382 ( \25971 , \25970_nR25586 );
not \U$17383 ( \25972 , \25637 );
and \U$17384 ( \25973 , RIddb9b88_3920, \25972 );
not \U$17385 ( \25974 , RIddb9b88_3920);
or \U$17386 ( \25975 , \25974 , \25752 );
nand \U$17387 ( \25976 , \22458 , \25788 );
nand \U$17388 ( \25977 , \22461 , \25835 );
nand \U$17389 ( \25978 , \25975 , \25976 , \25977 );
and \U$17390 ( \25979 , \25978 , \25637 );
or \U$17391 ( \25980 , \25973 , \25979 );
and \U$17393 ( \25981 , \25980 , 1'b1 );
or \U$17395 ( \25982 , \25981 , 1'b0 );
buf \U$17396 ( \25983 , \25982 );
_DC r25588_GF_IsGateDCbyConstraint ( \25984_nR25588 , \25983 , \21944 );
buf \U$17397 ( \25985 , \25984_nR25588 );
not \U$17398 ( \25986 , \25449 );
and \U$17399 ( \25987 , RIddba380_3921, \25986 );
not \U$17400 ( \25988 , RIddba380_3921);
or \U$17401 ( \25989 , \25988 , \25890 );
nand \U$17402 ( \25990 , \22478 , \25788 );
nand \U$17403 ( \25991 , \22481 , \25757 );
nand \U$17404 ( \25992 , \25989 , \25990 , \25991 );
and \U$17405 ( \25993 , \25992 , \25449 );
or \U$17406 ( \25994 , \25987 , \25993 );
and \U$17408 ( \25995 , \25994 , 1'b1 );
or \U$17410 ( \25996 , \25995 , 1'b0 );
buf \U$17411 ( \25997 , \25996 );
_DC r2558a_GF_IsGateDCbyConstraint ( \25998_nR2558a , \25997 , \21944 );
buf \U$17412 ( \25999 , \25998_nR2558a );
not \U$17413 ( \26000 , \22756 );
and \U$17414 ( \26001 , RIddbab78_3922, \26000 );
not \U$17415 ( \26002 , RIddbab78_3922);
or \U$17416 ( \26003 , \26002 , \25803 );
nand \U$17417 ( \26004 , \22498 , \25772 );
nand \U$17418 ( \26005 , \22501 , \25806 );
nand \U$17419 ( \26006 , \26003 , \26004 , \26005 );
and \U$17420 ( \26007 , \26006 , \22756 );
or \U$17421 ( \26008 , \26001 , \26007 );
and \U$17423 ( \26009 , \26008 , 1'b1 );
or \U$17425 ( \26010 , \26009 , 1'b0 );
buf \U$17426 ( \26011 , \26010 );
_DC r2558c_GF_IsGateDCbyConstraint ( \26012_nR2558c , \26011 , \21944 );
buf \U$17427 ( \26013 , \26012_nR2558c );
not \U$17428 ( \26014 , \25637 );
and \U$17429 ( \26015 , RIddbb370_3923, \26014 );
not \U$17430 ( \26016 , RIddbb370_3923);
or \U$17431 ( \26017 , \26016 , \25786 );
nand \U$17432 ( \26018 , \22519 , \25755 );
nand \U$17433 ( \26019 , \22522 , \25806 );
nand \U$17434 ( \26020 , \26017 , \26018 , \26019 );
and \U$17435 ( \26021 , \26020 , \25637 );
or \U$17436 ( \26022 , \26015 , \26021 );
and \U$17438 ( \26023 , \26022 , 1'b1 );
or \U$17440 ( \26024 , \26023 , 1'b0 );
buf \U$17441 ( \26025 , \26024 );
_DC r2558e_GF_IsGateDCbyConstraint ( \26026_nR2558e , \26025 , \21944 );
buf \U$17442 ( \26027 , \26026_nR2558e );
buf \U$17443 ( \26028 , \22104 );
not \U$17444 ( \26029 , \26028 );
and \U$17445 ( \26030 , RIddbbb68_3924, \26029 );
not \U$17446 ( \26031 , RIddbbb68_3924);
or \U$17447 ( \26032 , \26031 , \25786 );
nand \U$17448 ( \26033 , \22539 , \25755 );
nand \U$17449 ( \26034 , \22542 , \25790 );
nand \U$17450 ( \26035 , \26032 , \26033 , \26034 );
and \U$17451 ( \26036 , \26035 , \26028 );
or \U$17452 ( \26037 , \26030 , \26036 );
and \U$17454 ( \26038 , \26037 , 1'b1 );
or \U$17456 ( \26039 , \26038 , 1'b0 );
buf \U$17457 ( \26040 , \26039 );
_DC r25590_GF_IsGateDCbyConstraint ( \26041_nR25590 , \26040 , \21944 );
buf \U$17458 ( \26042 , \26041_nR25590 );
not \U$17459 ( \26043 , \22756 );
and \U$17460 ( \26044 , RIddbc360_3925, \26043 );
not \U$17461 ( \26045 , RIddbc360_3925);
or \U$17462 ( \26046 , \26045 , \25752 );
nand \U$17463 ( \26047 , \22559 , \25788 );
nand \U$17464 ( \26048 , \22562 , \25790 );
nand \U$17465 ( \26049 , \26046 , \26047 , \26048 );
and \U$17466 ( \26050 , \26049 , \22756 );
or \U$17467 ( \26051 , \26044 , \26050 );
and \U$17469 ( \26052 , \26051 , 1'b1 );
or \U$17471 ( \26053 , \26052 , 1'b0 );
buf \U$17472 ( \26054 , \26053 );
_DC r25594_GF_IsGateDCbyConstraint ( \26055_nR25594 , \26054 , \21944 );
buf \U$17473 ( \26056 , \26055_nR25594 );
not \U$17474 ( \26057 , \25637 );
and \U$17475 ( \26058 , RIddbcb58_3926, \26057 );
not \U$17476 ( \26059 , RIddbcb58_3926);
or \U$17477 ( \26060 , \26059 , \25890 );
nand \U$17478 ( \26061 , \22579 , \25755 );
nand \U$17479 ( \26062 , \22582 , \25835 );
nand \U$17480 ( \26063 , \26060 , \26061 , \26062 );
and \U$17481 ( \26064 , \26063 , \25637 );
or \U$17482 ( \26065 , \26058 , \26064 );
and \U$17484 ( \26066 , \26065 , 1'b1 );
or \U$17486 ( \26067 , \26066 , 1'b0 );
buf \U$17487 ( \26068 , \26067 );
_DC r25596_GF_IsGateDCbyConstraint ( \26069_nR25596 , \26068 , \21944 );
buf \U$17488 ( \26070 , \26069_nR25596 );
not \U$17489 ( \26071 , \26028 );
and \U$17490 ( \26072 , RIddbd350_3927, \26071 );
not \U$17491 ( \26073 , RIddbd350_3927);
or \U$17492 ( \26074 , \26073 , \25770 );
nand \U$17493 ( \26075 , \22599 , \25788 );
nand \U$17494 ( \26076 , \22602 , \25757 );
nand \U$17495 ( \26077 , \26074 , \26075 , \26076 );
and \U$17496 ( \26078 , \26077 , \26028 );
or \U$17497 ( \26079 , \26072 , \26078 );
and \U$17499 ( \26080 , \26079 , 1'b1 );
or \U$17501 ( \26081 , \26080 , 1'b0 );
buf \U$17502 ( \26082 , \26081 );
_DC r25598_GF_IsGateDCbyConstraint ( \26083_nR25598 , \26082 , \21944 );
buf \U$17503 ( \26084 , \26083_nR25598 );
not \U$17504 ( \26085 , \22104 );
and \U$17505 ( \26086 , RIddbdb48_3928, \26085 );
not \U$17506 ( \26087 , RIddbdb48_3928);
or \U$17507 ( \26088 , \26087 , \25803 );
nand \U$17508 ( \26089 , \22619 , \25772 );
nand \U$17509 ( \26090 , \22622 , \25790 );
nand \U$17510 ( \26091 , \26088 , \26089 , \26090 );
and \U$17511 ( \26092 , \26091 , \22104 );
or \U$17512 ( \26093 , \26086 , \26092 );
and \U$17514 ( \26094 , \26093 , 1'b1 );
or \U$17516 ( \26095 , \26094 , 1'b0 );
buf \U$17517 ( \26096 , \26095 );
_DC r2559a_GF_IsGateDCbyConstraint ( \26097_nR2559a , \26096 , \21944 );
buf \U$17518 ( \26098 , \26097_nR2559a );
not \U$17519 ( \26099 , \25637 );
and \U$17520 ( \26100 , RIddbe340_3929, \26099 );
not \U$17521 ( \26101 , RIddbe340_3929);
or \U$17522 ( \26102 , \26101 , \25786 );
nand \U$17523 ( \26103 , \22640 , \25755 );
nand \U$17524 ( \26104 , \22643 , \25806 );
nand \U$17525 ( \26105 , \26102 , \26103 , \26104 );
and \U$17526 ( \26106 , \26105 , \25637 );
or \U$17527 ( \26107 , \26100 , \26106 );
and \U$17529 ( \26108 , \26107 , 1'b1 );
or \U$17531 ( \26109 , \26108 , 1'b0 );
buf \U$17532 ( \26110 , \26109 );
_DC r2559c_GF_IsGateDCbyConstraint ( \26111_nR2559c , \26110 , \21944 );
buf \U$17533 ( \26112 , \26111_nR2559c );
not \U$17534 ( \26113 , \26028 );
and \U$17535 ( \26114 , RIddbeb38_3930, \26113 );
not \U$17536 ( \26115 , RIddbeb38_3930);
or \U$17537 ( \26116 , \26115 , \25770 );
nand \U$17538 ( \26117 , \22660 , \25755 );
nand \U$17539 ( \26118 , \22663 , \25835 );
nand \U$17540 ( \26119 , \26116 , \26117 , \26118 );
and \U$17541 ( \26120 , \26119 , \26028 );
or \U$17542 ( \26121 , \26114 , \26120 );
and \U$17544 ( \26122 , \26121 , 1'b1 );
or \U$17546 ( \26123 , \26122 , 1'b0 );
buf \U$17547 ( \26124 , \26123 );
_DC r2559e_GF_IsGateDCbyConstraint ( \26125_nR2559e , \26124 , \21944 );
buf \U$17548 ( \26126 , \26125_nR2559e );
not \U$17549 ( \26127 , \23038 );
and \U$17550 ( \26128 , RIddbf330_3931, \26127 );
not \U$17551 ( \26129 , RIddbf330_3931);
or \U$17552 ( \26130 , \26129 , \25752 );
nand \U$17553 ( \26131 , \22681 , \25772 );
nand \U$17554 ( \26132 , \22684 , \25835 );
nand \U$17555 ( \26133 , \26130 , \26131 , \26132 );
and \U$17556 ( \26134 , \26133 , \23038 );
or \U$17557 ( \26135 , \26128 , \26134 );
and \U$17559 ( \26136 , \26135 , 1'b1 );
or \U$17561 ( \26137 , \26136 , 1'b0 );
buf \U$17562 ( \26138 , \26137 );
_DC r255a0_GF_IsGateDCbyConstraint ( \26139_nR255a0 , \26138 , \21944 );
buf \U$17563 ( \26140 , \26139_nR255a0 );
not \U$17564 ( \26141 , \25637 );
and \U$17565 ( \26142 , RIddbfb28_3932, \26141 );
not \U$17566 ( \26143 , RIddbfb28_3932);
or \U$17567 ( \26144 , \26143 , \25752 );
nand \U$17568 ( \26145 , \22701 , \25755 );
nand \U$17569 ( \26146 , \22704 , \25757 );
nand \U$17570 ( \26147 , \26144 , \26145 , \26146 );
and \U$17571 ( \26148 , \26147 , \25637 );
or \U$17572 ( \26149 , \26142 , \26148 );
and \U$17574 ( \26150 , \26149 , 1'b1 );
or \U$17576 ( \26151 , \26150 , 1'b0 );
buf \U$17577 ( \26152 , \26151 );
_DC r255a2_GF_IsGateDCbyConstraint ( \26153_nR255a2 , \26152 , \21944 );
buf \U$17578 ( \26154 , \26153_nR255a2 );
not \U$17579 ( \26155 , \26028 );
and \U$17580 ( \26156 , RIddc0320_3933, \26155 );
not \U$17581 ( \26157 , RIddc0320_3933);
or \U$17582 ( \26158 , \26157 , \25890 );
nand \U$17583 ( \26159 , \22721 , \25788 );
nand \U$17584 ( \26160 , \22724 , \25806 );
nand \U$17585 ( \26161 , \26158 , \26159 , \26160 );
and \U$17586 ( \26162 , \26161 , \26028 );
or \U$17587 ( \26163 , \26156 , \26162 );
and \U$17589 ( \26164 , \26163 , 1'b1 );
or \U$17591 ( \26165 , \26164 , 1'b0 );
buf \U$17592 ( \26166 , \26165 );
_DC r255a4_GF_IsGateDCbyConstraint ( \26167_nR255a4 , \26166 , \21944 );
buf \U$17593 ( \26168 , \26167_nR255a4 );
not \U$17594 ( \26169 , \22104 );
and \U$17595 ( \26170 , RIddc0b18_3934, \26169 );
not \U$17596 ( \26171 , RIddc0b18_3934);
or \U$17597 ( \26172 , \26171 , \25803 );
nand \U$17598 ( \26173 , \22741 , \25755 );
nand \U$17599 ( \26174 , \22744 , \25757 );
nand \U$17600 ( \26175 , \26172 , \26173 , \26174 );
and \U$17601 ( \26176 , \26175 , \22104 );
or \U$17602 ( \26177 , \26170 , \26176 );
and \U$17604 ( \26178 , \26177 , 1'b1 );
or \U$17606 ( \26179 , \26178 , 1'b0 );
buf \U$17607 ( \26180 , \26179 );
_DC r255a6_GF_IsGateDCbyConstraint ( \26181_nR255a6 , \26180 , \21944 );
buf \U$17608 ( \26182 , \26181_nR255a6 );
buf \U$17609 ( \26183 , \24117 );
not \U$17610 ( \26184 , \26183 );
and \U$17611 ( \26185 , RIddc1310_3935, \26184 );
not \U$17612 ( \26186 , RIddc1310_3935);
or \U$17613 ( \26187 , \26186 , \25770 );
nand \U$17614 ( \26188 , \22763 , \25772 );
nand \U$17615 ( \26189 , \22766 , \25806 );
nand \U$17616 ( \26190 , \26187 , \26188 , \26189 );
and \U$17617 ( \26191 , \26190 , \26183 );
or \U$17618 ( \26192 , \26185 , \26191 );
and \U$17620 ( \26193 , \26192 , 1'b1 );
or \U$17622 ( \26194 , \26193 , 1'b0 );
buf \U$17623 ( \26195 , \26194 );
_DC r255aa_GF_IsGateDCbyConstraint ( \26196_nR255aa , \26195 , \21944 );
buf \U$17624 ( \26197 , \26196_nR255aa );
not \U$17625 ( \26198 , \26028 );
and \U$17626 ( \26199 , RIddc1b08_3936, \26198 );
not \U$17627 ( \26200 , RIddc1b08_3936);
or \U$17628 ( \26201 , \26200 , \25890 );
nand \U$17629 ( \26202 , \22783 , \25755 );
nand \U$17630 ( \26203 , \22786 , \25757 );
nand \U$17631 ( \26204 , \26201 , \26202 , \26203 );
and \U$17632 ( \26205 , \26204 , \26028 );
or \U$17633 ( \26206 , \26199 , \26205 );
and \U$17635 ( \26207 , \26206 , 1'b1 );
or \U$17637 ( \26208 , \26207 , 1'b0 );
buf \U$17638 ( \26209 , \26208 );
_DC r255ac_GF_IsGateDCbyConstraint ( \26210_nR255ac , \26209 , \21944 );
buf \U$17639 ( \26211 , \26210_nR255ac );
not \U$17640 ( \26212 , \22756 );
and \U$17641 ( \26213 , RIddc2300_3937, \26212 );
not \U$17642 ( \26214 , RIddc2300_3937);
or \U$17643 ( \26215 , \26214 , \25752 );
nand \U$17644 ( \26216 , \22803 , \25772 );
nand \U$17645 ( \26217 , \22806 , \25835 );
nand \U$17646 ( \26218 , \26215 , \26216 , \26217 );
and \U$17647 ( \26219 , \26218 , \22756 );
or \U$17648 ( \26220 , \26213 , \26219 );
and \U$17650 ( \26221 , \26220 , 1'b1 );
or \U$17652 ( \26222 , \26221 , 1'b0 );
buf \U$17653 ( \26223 , \26222 );
_DC r255ae_GF_IsGateDCbyConstraint ( \26224_nR255ae , \26223 , \21944 );
buf \U$17654 ( \26225 , \26224_nR255ae );
not \U$17655 ( \26226 , \26183 );
and \U$17656 ( \26227 , RIddc2af8_3938, \26226 );
not \U$17657 ( \26228 , RIddc2af8_3938);
or \U$17658 ( \26229 , \26228 , \25890 );
nand \U$17659 ( \26230 , \22823 , \25788 );
nand \U$17660 ( \26231 , \22826 , \25790 );
nand \U$17661 ( \26232 , \26229 , \26230 , \26231 );
and \U$17662 ( \26233 , \26232 , \26183 );
or \U$17663 ( \26234 , \26227 , \26233 );
and \U$17665 ( \26235 , \26234 , 1'b1 );
or \U$17667 ( \26236 , \26235 , 1'b0 );
buf \U$17668 ( \26237 , \26236 );
_DC r255b0_GF_IsGateDCbyConstraint ( \26238_nR255b0 , \26237 , \21944 );
buf \U$17669 ( \26239 , \26238_nR255b0 );
not \U$17670 ( \26240 , \26028 );
and \U$17671 ( \26241 , RIddc32f0_3939, \26240 );
not \U$17672 ( \26242 , RIddc32f0_3939);
or \U$17673 ( \26243 , \26242 , \25803 );
nand \U$17674 ( \26244 , \22843 , \25788 );
nand \U$17675 ( \26245 , \22846 , \25835 );
nand \U$17676 ( \26246 , \26243 , \26244 , \26245 );
and \U$17677 ( \26247 , \26246 , \26028 );
or \U$17678 ( \26248 , \26241 , \26247 );
and \U$17680 ( \26249 , \26248 , 1'b1 );
or \U$17682 ( \26250 , \26249 , 1'b0 );
buf \U$17683 ( \26251 , \26250 );
_DC r255b2_GF_IsGateDCbyConstraint ( \26252_nR255b2 , \26251 , \21944 );
buf \U$17684 ( \26253 , \26252_nR255b2 );
not \U$17685 ( \26254 , \22195 );
and \U$17686 ( \26255 , RIddc3ae8_3940, \26254 );
not \U$17687 ( \26256 , RIddc3ae8_3940);
or \U$17688 ( \26257 , \26256 , \25786 );
nand \U$17689 ( \26258 , \22863 , \25772 );
nand \U$17690 ( \26259 , \22866 , \25806 );
nand \U$17691 ( \26260 , \26257 , \26258 , \26259 );
and \U$17692 ( \26261 , \26260 , \22195 );
or \U$17693 ( \26262 , \26255 , \26261 );
and \U$17695 ( \26263 , \26262 , 1'b1 );
or \U$17697 ( \26264 , \26263 , 1'b0 );
buf \U$17698 ( \26265 , \26264 );
_DC r255b4_GF_IsGateDCbyConstraint ( \26266_nR255b4 , \26265 , \21944 );
buf \U$17699 ( \26267 , \26266_nR255b4 );
not \U$17700 ( \26268 , \26183 );
and \U$17701 ( \26269 , RIddc42e0_3941, \26268 );
not \U$17702 ( \26270 , RIddc42e0_3941);
or \U$17703 ( \26271 , \26270 , \25803 );
nand \U$17704 ( \26272 , \22883 , \25788 );
nand \U$17705 ( \26273 , \22886 , \25790 );
nand \U$17706 ( \26274 , \26271 , \26272 , \26273 );
and \U$17707 ( \26275 , \26274 , \26183 );
or \U$17708 ( \26276 , \26269 , \26275 );
and \U$17710 ( \26277 , \26276 , 1'b1 );
or \U$17712 ( \26278 , \26277 , 1'b0 );
buf \U$17713 ( \26279 , \26278 );
_DC r255b6_GF_IsGateDCbyConstraint ( \26280_nR255b6 , \26279 , \21944 );
buf \U$17714 ( \26281 , \26280_nR255b6 );
not \U$17715 ( \26282 , \26028 );
and \U$17716 ( \26283 , RIddc4ad8_3942, \26282 );
not \U$17717 ( \26284 , RIddc4ad8_3942);
or \U$17718 ( \26285 , \26284 , \25770 );
nand \U$17719 ( \26286 , \22905 , \25755 );
nand \U$17720 ( \26287 , \22908 , \25835 );
nand \U$17721 ( \26288 , \26285 , \26286 , \26287 );
and \U$17722 ( \26289 , \26288 , \26028 );
or \U$17723 ( \26290 , \26283 , \26289 );
and \U$17725 ( \26291 , \26290 , 1'b1 );
or \U$17727 ( \26292 , \26291 , 1'b0 );
buf \U$17728 ( \26293 , \26292 );
_DC r255b8_GF_IsGateDCbyConstraint ( \26294_nR255b8 , \26293 , \21944 );
buf \U$17729 ( \26295 , \26294_nR255b8 );
not \U$17730 ( \26296 , \22104 );
and \U$17731 ( \26297 , RIddc52d0_3943, \26296 );
not \U$17732 ( \26298 , RIddc52d0_3943);
or \U$17733 ( \26299 , \26298 , \25752 );
nand \U$17734 ( \26300 , \22925 , \25755 );
nand \U$17735 ( \26301 , \22928 , \25757 );
nand \U$17736 ( \26302 , \26299 , \26300 , \26301 );
and \U$17737 ( \26303 , \26302 , \22104 );
or \U$17738 ( \26304 , \26297 , \26303 );
and \U$17740 ( \26305 , \26304 , 1'b1 );
or \U$17742 ( \26306 , \26305 , 1'b0 );
buf \U$17743 ( \26307 , \26306 );
_DC r255ba_GF_IsGateDCbyConstraint ( \26308_nR255ba , \26307 , \21944 );
buf \U$17744 ( \26309 , \26308_nR255ba );
not \U$17745 ( \26310 , \26183 );
and \U$17746 ( \26311 , RIddc5ac8_3944, \26310 );
not \U$17747 ( \26312 , RIddc5ac8_3944);
or \U$17748 ( \26313 , \26312 , \25890 );
nand \U$17749 ( \26314 , \22945 , \25755 );
nand \U$17750 ( \26315 , \22948 , \25790 );
nand \U$17751 ( \26316 , \26313 , \26314 , \26315 );
and \U$17752 ( \26317 , \26316 , \26183 );
or \U$17753 ( \26318 , \26311 , \26317 );
and \U$17755 ( \26319 , \26318 , 1'b1 );
or \U$17757 ( \26320 , \26319 , 1'b0 );
buf \U$17758 ( \26321 , \26320 );
_DC r255bc_GF_IsGateDCbyConstraint ( \26322_nR255bc , \26321 , \21944 );
buf \U$17759 ( \26323 , \26322_nR255bc );
not \U$17760 ( \26324 , \26028 );
and \U$17761 ( \26325 , RIddc62c0_3945, \26324 );
not \U$17762 ( \26326 , RIddc62c0_3945);
or \U$17763 ( \26327 , \26326 , \25786 );
nand \U$17764 ( \26328 , \22965 , \25755 );
nand \U$17765 ( \26329 , \22968 , \25806 );
nand \U$17766 ( \26330 , \26327 , \26328 , \26329 );
and \U$17767 ( \26331 , \26330 , \26028 );
or \U$17768 ( \26332 , \26325 , \26331 );
and \U$17770 ( \26333 , \26332 , 1'b1 );
or \U$17772 ( \26334 , \26333 , 1'b0 );
buf \U$17773 ( \26335 , \26334 );
_DC r255c0_GF_IsGateDCbyConstraint ( \26336_nR255c0 , \26335 , \21944 );
buf \U$17774 ( \26337 , \26336_nR255c0 );
not \U$17775 ( \26338 , \24117 );
and \U$17776 ( \26339 , RIddc6ab8_3946, \26338 );
not \U$17777 ( \26340 , RIddc6ab8_3946);
or \U$17778 ( \26341 , \26340 , \25786 );
nand \U$17779 ( \26342 , \22984 , \25772 );
nand \U$17780 ( \26343 , \22987 , \25835 );
nand \U$17781 ( \26344 , \26341 , \26342 , \26343 );
and \U$17782 ( \26345 , \26344 , \24117 );
or \U$17783 ( \26346 , \26339 , \26345 );
and \U$17785 ( \26347 , \26346 , 1'b1 );
or \U$17787 ( \26348 , \26347 , 1'b0 );
buf \U$17788 ( \26349 , \26348 );
_DC r255c2_GF_IsGateDCbyConstraint ( \26350_nR255c2 , \26349 , \21944 );
buf \U$17789 ( \26351 , \26350_nR255c2 );
not \U$17790 ( \26352 , \26183 );
and \U$17791 ( \26353 , RIddc72b0_3947, \26352 );
not \U$17792 ( \26354 , RIddc72b0_3947);
or \U$17793 ( \26355 , \26354 , \25770 );
nand \U$17794 ( \26356 , \23003 , \25772 );
nand \U$17795 ( \26357 , \23006 , \25757 );
nand \U$17796 ( \26358 , \26355 , \26356 , \26357 );
and \U$17797 ( \26359 , \26358 , \26183 );
or \U$17798 ( \26360 , \26353 , \26359 );
and \U$17800 ( \26361 , \26360 , 1'b1 );
or \U$17802 ( \26362 , \26361 , 1'b0 );
buf \U$17803 ( \26363 , \26362 );
_DC r255c4_GF_IsGateDCbyConstraint ( \26364_nR255c4 , \26363 , \21944 );
buf \U$17804 ( \26365 , \26364_nR255c4 );
not \U$17805 ( \26366 , \26028 );
and \U$17806 ( \26367 , RIddc7aa8_3948, \26366 );
not \U$17807 ( \26368 , RIddc7aa8_3948);
or \U$17808 ( \26369 , \26368 , \25752 );
nand \U$17809 ( \26370 , \23023 , \25772 );
nand \U$17810 ( \26371 , \23026 , \25757 );
nand \U$17811 ( \26372 , \26369 , \26370 , \26371 );
and \U$17812 ( \26373 , \26372 , \26028 );
or \U$17813 ( \26374 , \26367 , \26373 );
and \U$17815 ( \26375 , \26374 , 1'b1 );
or \U$17817 ( \26376 , \26375 , 1'b0 );
buf \U$17818 ( \26377 , \26376 );
_DC r255c6_GF_IsGateDCbyConstraint ( \26378_nR255c6 , \26377 , \21944 );
buf \U$17819 ( \26379 , \26378_nR255c6 );
not \U$17820 ( \26380 , \22195 );
and \U$17821 ( \26381 , RIddc82a0_3949, \26380 );
not \U$17822 ( \26382 , RIddc82a0_3949);
or \U$17823 ( \26383 , \26382 , \25890 );
nand \U$17824 ( \26384 , \23045 , \25772 );
nand \U$17825 ( \26385 , \23048 , \25806 );
nand \U$17826 ( \26386 , \26383 , \26384 , \26385 );
and \U$17827 ( \26387 , \26386 , \22195 );
or \U$17828 ( \26388 , \26381 , \26387 );
and \U$17830 ( \26389 , \26388 , 1'b1 );
or \U$17832 ( \26390 , \26389 , 1'b0 );
buf \U$17833 ( \26391 , \26390 );
_DC r255c8_GF_IsGateDCbyConstraint ( \26392_nR255c8 , \26391 , \21944 );
buf \U$17834 ( \26393 , \26392_nR255c8 );
not \U$17835 ( \26394 , \26183 );
and \U$17836 ( \26395 , RIddc8a98_3950, \26394 );
not \U$17837 ( \26396 , RIddc8a98_3950);
or \U$17838 ( \26397 , \26396 , \25770 );
nand \U$17839 ( \26398 , \23065 , \25788 );
nand \U$17840 ( \26399 , \23068 , \25790 );
nand \U$17841 ( \26400 , \26397 , \26398 , \26399 );
and \U$17842 ( \26401 , \26400 , \26183 );
or \U$17843 ( \26402 , \26395 , \26401 );
and \U$17845 ( \26403 , \26402 , 1'b1 );
or \U$17847 ( \26404 , \26403 , 1'b0 );
buf \U$17848 ( \26405 , \26404 );
_DC r255ca_GF_IsGateDCbyConstraint ( \26406_nR255ca , \26405 , \21944 );
buf \U$17849 ( \26407 , \26406_nR255ca );
not \U$17850 ( \26408 , \26028 );
and \U$17851 ( \26409 , RIddc9290_3951, \26408 );
not \U$17852 ( \26410 , RIddc9290_3951);
or \U$17853 ( \26411 , \26410 , \25803 );
nand \U$17854 ( \26412 , \23085 , \25772 );
nand \U$17855 ( \26413 , \23088 , \25790 );
nand \U$17856 ( \26414 , \26411 , \26412 , \26413 );
and \U$17857 ( \26415 , \26414 , \26028 );
or \U$17858 ( \26416 , \26409 , \26415 );
and \U$17860 ( \26417 , \26416 , 1'b1 );
or \U$17862 ( \26418 , \26417 , 1'b0 );
buf \U$17863 ( \26419 , \26418 );
_DC r255cc_GF_IsGateDCbyConstraint ( \26420_nR255cc , \26419 , \21944 );
buf \U$17864 ( \26421 , \26420_nR255cc );
not \U$17865 ( \26422 , \23038 );
and \U$17866 ( \26423 , RIddc9a88_3952, \26422 );
not \U$17867 ( \26424 , RIddc9a88_3952);
or \U$17868 ( \26425 , \26424 , \25786 );
nand \U$17869 ( \26426 , \23105 , \25772 );
nand \U$17870 ( \26427 , \23108 , \25757 );
nand \U$17871 ( \26428 , \26425 , \26426 , \26427 );
and \U$17872 ( \26429 , \26428 , \23038 );
or \U$17873 ( \26430 , \26423 , \26429 );
and \U$17875 ( \26431 , \26430 , 1'b1 );
or \U$17877 ( \26432 , \26431 , 1'b0 );
buf \U$17878 ( \26433 , \26432 );
_DC r255ce_GF_IsGateDCbyConstraint ( \26434_nR255ce , \26433 , \21944 );
buf \U$17879 ( \26435 , \26434_nR255ce );
not \U$17880 ( \26436 , \26183 );
and \U$17881 ( \26437 , RIddca280_3953, \26436 );
not \U$17882 ( \26438 , RIddca280_3953);
or \U$17883 ( \26439 , \26438 , \25770 );
nand \U$17884 ( \26440 , \23125 , \25788 );
nand \U$17885 ( \26441 , \23128 , \25835 );
nand \U$17886 ( \26442 , \26439 , \26440 , \26441 );
and \U$17887 ( \26443 , \26442 , \26183 );
or \U$17888 ( \26444 , \26437 , \26443 );
and \U$17890 ( \26445 , \26444 , 1'b1 );
or \U$17892 ( \26446 , \26445 , 1'b0 );
buf \U$17893 ( \26447 , \26446 );
_DC r255d0_GF_IsGateDCbyConstraint ( \26448_nR255d0 , \26447 , \21944 );
buf \U$17894 ( \26449 , \26448_nR255d0 );
not \U$17895 ( \26450 , \26028 );
and \U$17896 ( \26451 , RIddcaa78_3954, \26450 );
not \U$17897 ( \26452 , RIddcaa78_3954);
or \U$17898 ( \26453 , \26452 , \25752 );
nand \U$17899 ( \26454 , \23145 , \25788 );
nand \U$17900 ( \26455 , \23148 , \25835 );
nand \U$17901 ( \26456 , \26453 , \26454 , \26455 );
and \U$17902 ( \26457 , \26456 , \26028 );
or \U$17903 ( \26458 , \26451 , \26457 );
and \U$17905 ( \26459 , \26458 , 1'b1 );
or \U$17907 ( \26460 , \26459 , 1'b0 );
buf \U$17908 ( \26461 , \26460 );
_DC r255d2_GF_IsGateDCbyConstraint ( \26462_nR255d2 , \26461 , \21944 );
buf \U$17909 ( \26463 , \26462_nR255d2 );
not \U$17910 ( \26464 , \22756 );
and \U$17911 ( \26465 , RIddcb270_3955, \26464 );
not \U$17912 ( \26466 , RIddcb270_3955);
or \U$17913 ( \26467 , \26466 , \25890 );
nand \U$17914 ( \26468 , \23165 , \25755 );
nand \U$17915 ( \26469 , \23168 , \25806 );
nand \U$17916 ( \26470 , \26467 , \26468 , \26469 );
and \U$17917 ( \26471 , \26470 , \22756 );
or \U$17918 ( \26472 , \26465 , \26471 );
and \U$17920 ( \26473 , \26472 , 1'b1 );
or \U$17922 ( \26474 , \26473 , 1'b0 );
buf \U$17923 ( \26475 , \26474 );
_DC r255d6_GF_IsGateDCbyConstraint ( \26476_nR255d6 , \26475 , \21944 );
buf \U$17924 ( \26477 , \26476_nR255d6 );
not \U$17925 ( \26478 , \26183 );
and \U$17926 ( \26479 , RIddcba68_3956, \26478 );
not \U$17927 ( \26480 , RIddcba68_3956);
or \U$17928 ( \26481 , \26480 , \25803 );
nand \U$17929 ( \26482 , \23184 , \25788 );
nand \U$17930 ( \26483 , \23187 , \25806 );
nand \U$17931 ( \26484 , \26481 , \26482 , \26483 );
and \U$17932 ( \26485 , \26484 , \26183 );
or \U$17933 ( \26486 , \26479 , \26485 );
and \U$17935 ( \26487 , \26486 , 1'b1 );
or \U$17937 ( \26488 , \26487 , 1'b0 );
buf \U$17938 ( \26489 , \26488 );
_DC r255d8_GF_IsGateDCbyConstraint ( \26490_nR255d8 , \26489 , \21944 );
buf \U$17939 ( \26491 , \26490_nR255d8 );
not \U$17940 ( \26492 , \26028 );
and \U$17941 ( \26493 , RIddcc260_3957, \26492 );
not \U$17942 ( \26494 , RIddcc260_3957);
or \U$17943 ( \26495 , \26494 , \25786 );
nand \U$17944 ( \26496 , \23204 , \25772 );
nand \U$17945 ( \26497 , \23207 , \25835 );
nand \U$17946 ( \26498 , \26495 , \26496 , \26497 );
and \U$17947 ( \26499 , \26498 , \26028 );
or \U$17948 ( \26500 , \26493 , \26499 );
and \U$17950 ( \26501 , \26500 , 1'b1 );
or \U$17952 ( \26502 , \26501 , 1'b0 );
buf \U$17953 ( \26503 , \26502 );
_DC r255da_GF_IsGateDCbyConstraint ( \26504_nR255da , \26503 , \21944 );
buf \U$17954 ( \26505 , \26504_nR255da );
not \U$17955 ( \26506 , \24155 );
and \U$17956 ( \26507 , RIddcca58_3958, \26506 );
not \U$17957 ( \26508 , RIddcca58_3958);
or \U$17958 ( \26509 , \26508 , \25770 );
nand \U$17959 ( \26510 , \23224 , \25772 );
nand \U$17960 ( \26511 , \23227 , \25757 );
nand \U$17961 ( \26512 , \26509 , \26510 , \26511 );
and \U$17962 ( \26513 , \26512 , \24155 );
or \U$17963 ( \26514 , \26507 , \26513 );
and \U$17965 ( \26515 , \26514 , 1'b1 );
or \U$17967 ( \26516 , \26515 , 1'b0 );
buf \U$17968 ( \26517 , \26516 );
_DC r255dc_GF_IsGateDCbyConstraint ( \26518_nR255dc , \26517 , \21944 );
buf \U$17969 ( \26519 , \26518_nR255dc );
not \U$17970 ( \26520 , \26183 );
and \U$17971 ( \26521 , RIddcd250_3959, \26520 );
not \U$17972 ( \26522 , RIddcd250_3959);
or \U$17973 ( \26523 , \26522 , \25890 );
nand \U$17974 ( \26524 , \23244 , \25772 );
nand \U$17975 ( \26525 , \23247 , \25757 );
nand \U$17976 ( \26526 , \26523 , \26524 , \26525 );
and \U$17977 ( \26527 , \26526 , \26183 );
or \U$17978 ( \26528 , \26521 , \26527 );
and \U$17980 ( \26529 , \26528 , 1'b1 );
or \U$17982 ( \26530 , \26529 , 1'b0 );
buf \U$17983 ( \26531 , \26530 );
_DC r255de_GF_IsGateDCbyConstraint ( \26532_nR255de , \26531 , \21944 );
buf \U$17984 ( \26533 , \26532_nR255de );
not \U$17985 ( \26534 , \22196 );
and \U$17986 ( \26535 , RIddcda48_3960, \26534 );
not \U$17987 ( \26536 , RIddcda48_3960);
or \U$17988 ( \26537 , \26536 , \25752 );
nand \U$17989 ( \26538 , \23264 , \25755 );
nand \U$17990 ( \26539 , \23267 , \25806 );
nand \U$17991 ( \26540 , \26537 , \26538 , \26539 );
and \U$17992 ( \26541 , \26540 , \22196 );
or \U$17993 ( \26542 , \26535 , \26541 );
and \U$17995 ( \26543 , \26542 , 1'b1 );
or \U$17997 ( \26544 , \26543 , 1'b0 );
buf \U$17998 ( \26545 , \26544 );
_DC r255e0_GF_IsGateDCbyConstraint ( \26546_nR255e0 , \26545 , \21944 );
buf \U$17999 ( \26547 , \26546_nR255e0 );
not \U$18000 ( \26548 , \22756 );
and \U$18001 ( \26549 , RIddce240_3961, \26548 );
not \U$18002 ( \26550 , RIddce240_3961);
or \U$18003 ( \26551 , \26550 , \25890 );
nand \U$18004 ( \26552 , \23284 , \25755 );
nand \U$18005 ( \26553 , \23287 , \25790 );
nand \U$18006 ( \26554 , \26551 , \26552 , \26553 );
and \U$18007 ( \26555 , \26554 , \22756 );
or \U$18008 ( \26556 , \26549 , \26555 );
and \U$18010 ( \26557 , \26556 , 1'b1 );
or \U$18012 ( \26558 , \26557 , 1'b0 );
buf \U$18013 ( \26559 , \26558 );
_DC r255e2_GF_IsGateDCbyConstraint ( \26560_nR255e2 , \26559 , \21944 );
buf \U$18014 ( \26561 , \26560_nR255e2 );
not \U$18015 ( \26562 , \26183 );
and \U$18016 ( \26563 , RIddcea38_3962, \26562 );
not \U$18017 ( \26564 , RIddcea38_3962);
or \U$18018 ( \26565 , \26564 , \25803 );
nand \U$18019 ( \26566 , \23303 , \25788 );
nand \U$18020 ( \26567 , \23306 , \25790 );
nand \U$18021 ( \26568 , \26565 , \26566 , \26567 );
and \U$18022 ( \26569 , \26568 , \26183 );
or \U$18023 ( \26570 , \26563 , \26569 );
and \U$18025 ( \26571 , \26570 , 1'b1 );
or \U$18027 ( \26572 , \26571 , 1'b0 );
buf \U$18028 ( \26573 , \26572 );
_DC r255e4_GF_IsGateDCbyConstraint ( \26574_nR255e4 , \26573 , \21944 );
buf \U$18029 ( \26575 , \26574_nR255e4 );
not \U$18030 ( \26576 , \22196 );
and \U$18031 ( \26577 , RIddcf230_3963, \26576 );
not \U$18032 ( \26578 , RIddcf230_3963);
or \U$18033 ( \26579 , \26578 , \25786 );
nand \U$18034 ( \26580 , \23323 , \25772 );
nand \U$18035 ( \26581 , \23326 , \25757 );
nand \U$18036 ( \26582 , \26579 , \26580 , \26581 );
and \U$18037 ( \26583 , \26582 , \22196 );
or \U$18038 ( \26584 , \26577 , \26583 );
and \U$18040 ( \26585 , \26584 , 1'b1 );
or \U$18042 ( \26586 , \26585 , 1'b0 );
buf \U$18043 ( \26587 , \26586 );
_DC r255e6_GF_IsGateDCbyConstraint ( \26588_nR255e6 , \26587 , \21944 );
buf \U$18044 ( \26589 , \26588_nR255e6 );
not \U$18045 ( \26590 , \22756 );
and \U$18046 ( \26591 , RIddcfa28_3964, \26590 );
not \U$18047 ( \26592 , RIddcfa28_3964);
or \U$18048 ( \26593 , \26592 , \25803 );
nand \U$18049 ( \26594 , \23343 , \25754 );
nand \U$18050 ( \26595 , \23346 , \25835 );
nand \U$18051 ( \26596 , \26593 , \26594 , \26595 );
and \U$18052 ( \26597 , \26596 , \22756 );
or \U$18053 ( \26598 , \26591 , \26597 );
and \U$18055 ( \26599 , \26598 , 1'b1 );
or \U$18057 ( \26600 , \26599 , 1'b0 );
buf \U$18058 ( \26601 , \26600 );
_DC r255e8_GF_IsGateDCbyConstraint ( \26602_nR255e8 , \26601 , \21944 );
buf \U$18059 ( \26603 , \26602_nR255e8 );
not \U$18060 ( \26604 , \26183 );
and \U$18061 ( \26605 , RIddd0220_3965, \26604 );
not \U$18062 ( \26606 , RIddd0220_3965);
or \U$18063 ( \26607 , \26606 , \25752 );
nand \U$18064 ( \26608 , \23364 , \25772 );
nand \U$18065 ( \26609 , \23367 , \25790 );
nand \U$18066 ( \26610 , \26607 , \26608 , \26609 );
and \U$18067 ( \26611 , \26610 , \26183 );
or \U$18068 ( \26612 , \26605 , \26611 );
and \U$18070 ( \26613 , \26612 , 1'b1 );
or \U$18072 ( \26614 , \26613 , 1'b0 );
buf \U$18073 ( \26615 , \26614 );
_DC r255ec_GF_IsGateDCbyConstraint ( \26616_nR255ec , \26615 , \21944 );
buf \U$18074 ( \26617 , \26616_nR255ec );
not \U$18075 ( \26618 , \22196 );
and \U$18076 ( \26619 , RIddd0a18_3966, \26618 );
not \U$18077 ( \26620 , RIddd0a18_3966);
or \U$18078 ( \26621 , \26620 , \25890 );
nand \U$18079 ( \26622 , \23384 , \25754 );
nand \U$18080 ( \26623 , \23387 , \25806 );
nand \U$18081 ( \26624 , \26621 , \26622 , \26623 );
and \U$18082 ( \26625 , \26624 , \22196 );
or \U$18083 ( \26626 , \26619 , \26625 );
and \U$18085 ( \26627 , \26626 , 1'b1 );
or \U$18087 ( \26628 , \26627 , 1'b0 );
buf \U$18088 ( \26629 , \26628 );
_DC r255ee_GF_IsGateDCbyConstraint ( \26630_nR255ee , \26629 , \21944 );
buf \U$18089 ( \26631 , \26630_nR255ee );
not \U$18090 ( \26632 , \24117 );
and \U$18091 ( \26633 , RIddd1210_3967, \26632 );
not \U$18092 ( \26634 , RIddd1210_3967);
or \U$18093 ( \26635 , \26634 , \25803 );
nand \U$18094 ( \26636 , \23404 , \25754 );
nand \U$18095 ( \26637 , \23407 , \25806 );
nand \U$18096 ( \26638 , \26635 , \26636 , \26637 );
and \U$18097 ( \26639 , \26638 , \24117 );
or \U$18098 ( \26640 , \26633 , \26639 );
and \U$18100 ( \26641 , \26640 , 1'b1 );
or \U$18102 ( \26642 , \26641 , 1'b0 );
buf \U$18103 ( \26643 , \26642 );
_DC r255f0_GF_IsGateDCbyConstraint ( \26644_nR255f0 , \26643 , \21944 );
buf \U$18104 ( \26645 , \26644_nR255f0 );
not \U$18105 ( \26646 , \26183 );
and \U$18106 ( \26647 , RIddd1a08_3968, \26646 );
not \U$18107 ( \26648 , RIddd1a08_3968);
or \U$18108 ( \26649 , \26648 , \25786 );
nand \U$18109 ( \26650 , \23424 , \25755 );
nand \U$18110 ( \26651 , \23427 , \25835 );
nand \U$18111 ( \26652 , \26649 , \26650 , \26651 );
and \U$18112 ( \26653 , \26652 , \26183 );
or \U$18113 ( \26654 , \26647 , \26653 );
and \U$18115 ( \26655 , \26654 , 1'b1 );
or \U$18117 ( \26656 , \26655 , 1'b0 );
buf \U$18118 ( \26657 , \26656 );
_DC r255f2_GF_IsGateDCbyConstraint ( \26658_nR255f2 , \26657 , \21944 );
buf \U$18119 ( \26659 , \26658_nR255f2 );
nor \U$18120 ( \26660 , \22123 , \22099 );
buf \U$18121 ( \26661 , \26660 );
not \U$18122 ( \26662 , \26661 );
and \U$18123 ( \26663 , RIdc0fbb8_3681, \26662 );
not \U$18124 ( \26664 , RIdc0fbb8_3681);
not \U$18125 ( \26665 , \26664 );
not \U$18126 ( \26666 , \22115 );
and \U$18127 ( \26667 , \26665 , \26666 );
buf \U$18128 ( \26668 , RIb86fc68_77);
buf \U$18129 ( \26669 , \26668 );
and \U$18130 ( \26670 , \26669 , \22115 );
or \U$18131 ( \26671 , \26667 , \26670 );
and \U$18132 ( \26672 , \26671 , \26661 );
or \U$18133 ( \26673 , \26663 , \26672 );
and \U$18135 ( \26674 , \26673 , 1'b1 );
or \U$18137 ( \26675 , \26674 , 1'b0 );
buf \U$18138 ( \26676 , \26675 );
_DC r253bc_GF_IsGateDCbyConstraint ( \26677_nR253bc , \26676 , \21944 );
buf \U$18139 ( \26678 , \26677_nR253bc );
buf \U$18140 ( \26679 , \26660 );
not \U$18141 ( \26680 , \26679 );
and \U$18142 ( \26681 , RIdc0f0f0_3682, \26680 );
not \U$18143 ( \26682 , RIdc0f0f0_3682);
not \U$18144 ( \26683 , \26682 );
not \U$18145 ( \26684 , \22115 );
and \U$18146 ( \26685 , \26683 , \26684 );
buf \U$18147 ( \26686 , RIb86fce0_76);
buf \U$18148 ( \26687 , \26686 );
and \U$18149 ( \26688 , \26687 , \22115 );
or \U$18150 ( \26689 , \26685 , \26688 );
and \U$18151 ( \26690 , \26689 , \26679 );
or \U$18152 ( \26691 , \26681 , \26690 );
and \U$18154 ( \26692 , \26691 , 1'b1 );
or \U$18156 ( \26693 , \26692 , 1'b0 );
buf \U$18157 ( \26694 , \26693 );
_DC r253be_GF_IsGateDCbyConstraint ( \26695_nR253be , \26694 , \21944 );
buf \U$18158 ( \26696 , \26695_nR253be );
not \U$18159 ( \26697 , \26661 );
and \U$18160 ( \26698 , RIdc0e5b0_3683, \26697 );
not \U$18161 ( \26699 , RIdc0e5b0_3683);
not \U$18162 ( \26700 , \26699 );
not \U$18163 ( \26701 , \22115 );
and \U$18164 ( \26702 , \26700 , \26701 );
buf \U$18165 ( \26703 , RIb86fd58_75);
buf \U$18166 ( \26704 , \26703 );
and \U$18167 ( \26705 , \26704 , \22115 );
or \U$18168 ( \26706 , \26702 , \26705 );
and \U$18169 ( \26707 , \26706 , \26661 );
or \U$18170 ( \26708 , \26698 , \26707 );
and \U$18172 ( \26709 , \26708 , 1'b1 );
or \U$18174 ( \26710 , \26709 , 1'b0 );
buf \U$18175 ( \26711 , \26710 );
_DC r253c0_GF_IsGateDCbyConstraint ( \26712_nR253c0 , \26711 , \21944 );
buf \U$18176 ( \26713 , \26712_nR253c0 );
not \U$18177 ( \26714 , \26679 );
and \U$18178 ( \26715 , RIdc0dae8_3684, \26714 );
not \U$18179 ( \26716 , RIdc0dae8_3684);
not \U$18180 ( \26717 , \26716 );
not \U$18181 ( \26718 , \22115 );
and \U$18182 ( \26719 , \26717 , \26718 );
buf \U$18183 ( \26720 , RIb87e8a8_74);
buf \U$18184 ( \26721 , \26720 );
and \U$18185 ( \26722 , \26721 , \22115 );
or \U$18186 ( \26723 , \26719 , \26722 );
and \U$18187 ( \26724 , \26723 , \26679 );
or \U$18188 ( \26725 , \26715 , \26724 );
and \U$18190 ( \26726 , \26725 , 1'b1 );
or \U$18192 ( \26727 , \26726 , 1'b0 );
buf \U$18193 ( \26728 , \26727 );
_DC r253c2_GF_IsGateDCbyConstraint ( \26729_nR253c2 , \26728 , \21944 );
buf \U$18194 ( \26730 , \26729_nR253c2 );
not \U$18195 ( \26731 , \26661 );
and \U$18196 ( \26732 , RIdc0cfa8_3685, \26731 );
not \U$18197 ( \26733 , RIdc0cfa8_3685);
not \U$18198 ( \26734 , \26733 );
not \U$18199 ( \26735 , \22115 );
and \U$18200 ( \26736 , \26734 , \26735 );
buf \U$18201 ( \26737 , RIb87e920_73);
buf \U$18202 ( \26738 , \26737 );
and \U$18203 ( \26739 , \26738 , \22115 );
or \U$18204 ( \26740 , \26736 , \26739 );
and \U$18205 ( \26741 , \26740 , \26661 );
or \U$18206 ( \26742 , \26732 , \26741 );
and \U$18208 ( \26743 , \26742 , 1'b1 );
or \U$18210 ( \26744 , \26743 , 1'b0 );
buf \U$18211 ( \26745 , \26744 );
_DC r253c4_GF_IsGateDCbyConstraint ( \26746_nR253c4 , \26745 , \21944 );
buf \U$18212 ( \26747 , \26746_nR253c4 );
not \U$18213 ( \26748 , \26679 );
and \U$18214 ( \26749 , RIdc0c3f0_3686, \26748 );
not \U$18215 ( \26750 , RIdc0c3f0_3686);
not \U$18216 ( \26751 , \26750 );
not \U$18217 ( \26752 , \22115 );
and \U$18218 ( \26753 , \26751 , \26752 );
buf \U$18219 ( \26754 , RIb87e998_72);
buf \U$18220 ( \26755 , \26754 );
and \U$18221 ( \26756 , \26755 , \22115 );
or \U$18222 ( \26757 , \26753 , \26756 );
and \U$18223 ( \26758 , \26757 , \26679 );
or \U$18224 ( \26759 , \26749 , \26758 );
and \U$18226 ( \26760 , \26759 , 1'b1 );
or \U$18228 ( \26761 , \26760 , 1'b0 );
buf \U$18229 ( \26762 , \26761 );
_DC r253c6_GF_IsGateDCbyConstraint ( \26763_nR253c6 , \26762 , \21944 );
buf \U$18230 ( \26764 , \26763_nR253c6 );
not \U$18231 ( \26765 , \26661 );
and \U$18232 ( \26766 , RIdc0b7c0_3687, \26765 );
not \U$18233 ( \26767 , RIdc0b7c0_3687);
not \U$18234 ( \26768 , \26767 );
not \U$18235 ( \26769 , \22115 );
and \U$18236 ( \26770 , \26768 , \26769 );
buf \U$18237 ( \26771 , RIb87ea10_71);
buf \U$18238 ( \26772 , \26771 );
and \U$18239 ( \26773 , \26772 , \22115 );
or \U$18240 ( \26774 , \26770 , \26773 );
and \U$18241 ( \26775 , \26774 , \26661 );
or \U$18242 ( \26776 , \26766 , \26775 );
and \U$18244 ( \26777 , \26776 , 1'b1 );
or \U$18246 ( \26778 , \26777 , 1'b0 );
buf \U$18247 ( \26779 , \26778 );
_DC r253c8_GF_IsGateDCbyConstraint ( \26780_nR253c8 , \26779 , \21944 );
buf \U$18248 ( \26781 , \26780_nR253c8 );
not \U$18249 ( \26782 , \26679 );
and \U$18250 ( \26783 , RIdc0ac08_3688, \26782 );
not \U$18251 ( \26784 , RIdc0ac08_3688);
not \U$18252 ( \26785 , \26784 );
not \U$18253 ( \26786 , \22115 );
and \U$18254 ( \26787 , \26785 , \26786 );
buf \U$18255 ( \26788 , RIb87ea88_70);
buf \U$18256 ( \26789 , \26788 );
and \U$18257 ( \26790 , \26789 , \22115 );
or \U$18258 ( \26791 , \26787 , \26790 );
and \U$18259 ( \26792 , \26791 , \26679 );
or \U$18260 ( \26793 , \26783 , \26792 );
and \U$18262 ( \26794 , \26793 , 1'b1 );
or \U$18264 ( \26795 , \26794 , 1'b0 );
buf \U$18265 ( \26796 , \26795 );
_DC r253ca_GF_IsGateDCbyConstraint ( \26797_nR253ca , \26796 , \21944 );
buf \U$18266 ( \26798 , \26797_nR253ca );
not \U$18267 ( \26799 , \26661 );
and \U$18268 ( \26800 , RIdc09f60_3689, \26799 );
not \U$18269 ( \26801 , RIdc09f60_3689);
not \U$18270 ( \26802 , \26801 );
not \U$18271 ( \26803 , \23448 );
and \U$18272 ( \26804 , \26802 , \26803 );
and \U$18273 ( \26805 , \26669 , \23448 );
or \U$18274 ( \26806 , \26804 , \26805 );
and \U$18275 ( \26807 , \26806 , \26661 );
or \U$18276 ( \26808 , \26800 , \26807 );
and \U$18278 ( \26809 , \26808 , 1'b1 );
or \U$18280 ( \26810 , \26809 , 1'b0 );
buf \U$18281 ( \26811 , \26810 );
_DC r253cc_GF_IsGateDCbyConstraint ( \26812_nR253cc , \26811 , \21944 );
buf \U$18282 ( \26813 , \26812_nR253cc );
not \U$18283 ( \26814 , \26679 );
and \U$18284 ( \26815 , RIdc093a8_3690, \26814 );
not \U$18285 ( \26816 , RIdc093a8_3690);
not \U$18286 ( \26817 , \26816 );
not \U$18287 ( \26818 , \23448 );
and \U$18288 ( \26819 , \26817 , \26818 );
and \U$18289 ( \26820 , \26687 , \23448 );
or \U$18290 ( \26821 , \26819 , \26820 );
and \U$18291 ( \26822 , \26821 , \26679 );
or \U$18292 ( \26823 , \26815 , \26822 );
and \U$18294 ( \26824 , \26823 , 1'b1 );
or \U$18296 ( \26825 , \26824 , 1'b0 );
buf \U$18297 ( \26826 , \26825 );
_DC r253ce_GF_IsGateDCbyConstraint ( \26827_nR253ce , \26826 , \21944 );
buf \U$18298 ( \26828 , \26827_nR253ce );
not \U$18299 ( \26829 , \26661 );
and \U$18300 ( \26830 , RIdc08700_3691, \26829 );
not \U$18301 ( \26831 , RIdc08700_3691);
not \U$18302 ( \26832 , \26831 );
not \U$18303 ( \26833 , \23448 );
and \U$18304 ( \26834 , \26832 , \26833 );
and \U$18305 ( \26835 , \26704 , \23448 );
or \U$18306 ( \26836 , \26834 , \26835 );
and \U$18307 ( \26837 , \26836 , \26661 );
or \U$18308 ( \26838 , \26830 , \26837 );
and \U$18310 ( \26839 , \26838 , 1'b1 );
or \U$18312 ( \26840 , \26839 , 1'b0 );
buf \U$18313 ( \26841 , \26840 );
_DC r253d0_GF_IsGateDCbyConstraint ( \26842_nR253d0 , \26841 , \21944 );
buf \U$18314 ( \26843 , \26842_nR253d0 );
not \U$18315 ( \26844 , \26679 );
and \U$18316 ( \26845 , RIdc07878_3692, \26844 );
not \U$18317 ( \26846 , RIdc07878_3692);
not \U$18318 ( \26847 , \26846 );
not \U$18319 ( \26848 , \23448 );
and \U$18320 ( \26849 , \26847 , \26848 );
and \U$18321 ( \26850 , \26721 , \23448 );
or \U$18322 ( \26851 , \26849 , \26850 );
and \U$18323 ( \26852 , \26851 , \26679 );
or \U$18324 ( \26853 , \26845 , \26852 );
and \U$18326 ( \26854 , \26853 , 1'b1 );
or \U$18328 ( \26855 , \26854 , 1'b0 );
buf \U$18329 ( \26856 , \26855 );
_DC r253d2_GF_IsGateDCbyConstraint ( \26857_nR253d2 , \26856 , \21944 );
buf \U$18330 ( \26858 , \26857_nR253d2 );
not \U$18331 ( \26859 , \26661 );
and \U$18332 ( \26860 , RIdc06270_3693, \26859 );
not \U$18333 ( \26861 , RIdc06270_3693);
not \U$18334 ( \26862 , \26861 );
not \U$18335 ( \26863 , \23448 );
and \U$18336 ( \26864 , \26862 , \26863 );
and \U$18337 ( \26865 , \26738 , \23448 );
or \U$18338 ( \26866 , \26864 , \26865 );
and \U$18339 ( \26867 , \26866 , \26661 );
or \U$18340 ( \26868 , \26860 , \26867 );
and \U$18342 ( \26869 , \26868 , 1'b1 );
or \U$18344 ( \26870 , \26869 , 1'b0 );
buf \U$18345 ( \26871 , \26870 );
_DC r253d4_GF_IsGateDCbyConstraint ( \26872_nR253d4 , \26871 , \21944 );
buf \U$18346 ( \26873 , \26872_nR253d4 );
not \U$18347 ( \26874 , \26679 );
and \U$18348 ( \26875 , RIdc05118_3694, \26874 );
not \U$18349 ( \26876 , RIdc05118_3694);
not \U$18350 ( \26877 , \26876 );
not \U$18351 ( \26878 , \23448 );
and \U$18352 ( \26879 , \26877 , \26878 );
and \U$18353 ( \26880 , \26755 , \23448 );
or \U$18354 ( \26881 , \26879 , \26880 );
and \U$18355 ( \26882 , \26881 , \26679 );
or \U$18356 ( \26883 , \26875 , \26882 );
and \U$18358 ( \26884 , \26883 , 1'b1 );
or \U$18360 ( \26885 , \26884 , 1'b0 );
buf \U$18361 ( \26886 , \26885 );
_DC r253d6_GF_IsGateDCbyConstraint ( \26887_nR253d6 , \26886 , \21944 );
buf \U$18362 ( \26888 , \26887_nR253d6 );
not \U$18363 ( \26889 , \26661 );
and \U$18364 ( \26890 , RIdc03b10_3695, \26889 );
not \U$18365 ( \26891 , RIdc03b10_3695);
not \U$18366 ( \26892 , \26891 );
not \U$18367 ( \26893 , \23448 );
and \U$18368 ( \26894 , \26892 , \26893 );
and \U$18369 ( \26895 , \26772 , \23448 );
or \U$18370 ( \26896 , \26894 , \26895 );
and \U$18371 ( \26897 , \26896 , \26661 );
or \U$18372 ( \26898 , \26890 , \26897 );
and \U$18374 ( \26899 , \26898 , 1'b1 );
or \U$18376 ( \26900 , \26899 , 1'b0 );
buf \U$18377 ( \26901 , \26900 );
_DC r253d8_GF_IsGateDCbyConstraint ( \26902_nR253d8 , \26901 , \21944 );
buf \U$18378 ( \26903 , \26902_nR253d8 );
not \U$18379 ( \26904 , \26679 );
and \U$18380 ( \26905 , RIdc029b8_3696, \26904 );
not \U$18381 ( \26906 , RIdc029b8_3696);
not \U$18382 ( \26907 , \26906 );
not \U$18383 ( \26908 , \23448 );
and \U$18384 ( \26909 , \26907 , \26908 );
and \U$18385 ( \26910 , \26789 , \23448 );
or \U$18386 ( \26911 , \26909 , \26910 );
and \U$18387 ( \26912 , \26911 , \26679 );
or \U$18388 ( \26913 , \26905 , \26912 );
and \U$18390 ( \26914 , \26913 , 1'b1 );
or \U$18392 ( \26915 , \26914 , 1'b0 );
buf \U$18393 ( \26916 , \26915 );
_DC r253da_GF_IsGateDCbyConstraint ( \26917_nR253da , \26916 , \21944 );
buf \U$18394 ( \26918 , \26917_nR253da );
not \U$18395 ( \26919 , \26661 );
and \U$18396 ( \26920 , RIdc013b0_3697, \26919 );
not \U$18397 ( \26921 , RIdc013b0_3697);
not \U$18398 ( \26922 , \26921 );
not \U$18399 ( \26923 , \24635 );
and \U$18400 ( \26924 , \26922 , \26923 );
and \U$18401 ( \26925 , \26669 , \24635 );
or \U$18402 ( \26926 , \26924 , \26925 );
and \U$18403 ( \26927 , \26926 , \26661 );
or \U$18404 ( \26928 , \26920 , \26927 );
and \U$18406 ( \26929 , \26928 , 1'b1 );
or \U$18408 ( \26930 , \26929 , 1'b0 );
buf \U$18409 ( \26931 , \26930 );
_DC r253dc_GF_IsGateDCbyConstraint ( \26932_nR253dc , \26931 , \21944 );
buf \U$18410 ( \26933 , \26932_nR253dc );
not \U$18411 ( \26934 , \26661 );
and \U$18412 ( \26935 , RIdc00258_3698, \26934 );
not \U$18413 ( \26936 , RIdc00258_3698);
not \U$18414 ( \26937 , \26936 );
not \U$18415 ( \26938 , \24635 );
and \U$18416 ( \26939 , \26937 , \26938 );
and \U$18417 ( \26940 , \26687 , \24635 );
or \U$18418 ( \26941 , \26939 , \26940 );
and \U$18419 ( \26942 , \26941 , \26661 );
or \U$18420 ( \26943 , \26935 , \26942 );
and \U$18422 ( \26944 , \26943 , 1'b1 );
or \U$18424 ( \26945 , \26944 , 1'b0 );
buf \U$18425 ( \26946 , \26945 );
_DC r253de_GF_IsGateDCbyConstraint ( \26947_nR253de , \26946 , \21944 );
buf \U$18426 ( \26948 , \26947_nR253de );
not \U$18427 ( \26949 , \26661 );
and \U$18428 ( \26950 , RIdbff100_3699, \26949 );
not \U$18429 ( \26951 , RIdbff100_3699);
not \U$18430 ( \26952 , \26951 );
not \U$18431 ( \26953 , \24635 );
and \U$18432 ( \26954 , \26952 , \26953 );
and \U$18433 ( \26955 , \26704 , \24635 );
or \U$18434 ( \26956 , \26954 , \26955 );
and \U$18435 ( \26957 , \26956 , \26661 );
or \U$18436 ( \26958 , \26950 , \26957 );
and \U$18438 ( \26959 , \26958 , 1'b1 );
or \U$18440 ( \26960 , \26959 , 1'b0 );
buf \U$18441 ( \26961 , \26960 );
_DC r253e0_GF_IsGateDCbyConstraint ( \26962_nR253e0 , \26961 , \21944 );
buf \U$18442 ( \26963 , \26962_nR253e0 );
not \U$18443 ( \26964 , \26661 );
and \U$18444 ( \26965 , RIdbfdaf8_3700, \26964 );
not \U$18445 ( \26966 , RIdbfdaf8_3700);
not \U$18446 ( \26967 , \26966 );
not \U$18447 ( \26968 , \24635 );
and \U$18448 ( \26969 , \26967 , \26968 );
and \U$18449 ( \26970 , \26721 , \24635 );
or \U$18450 ( \26971 , \26969 , \26970 );
and \U$18451 ( \26972 , \26971 , \26661 );
or \U$18452 ( \26973 , \26965 , \26972 );
and \U$18454 ( \26974 , \26973 , 1'b1 );
or \U$18456 ( \26975 , \26974 , 1'b0 );
buf \U$18457 ( \26976 , \26975 );
_DC r253e2_GF_IsGateDCbyConstraint ( \26977_nR253e2 , \26976 , \21944 );
buf \U$18458 ( \26978 , \26977_nR253e2 );
not \U$18459 ( \26979 , \26661 );
and \U$18460 ( \26980 , RIdbfc9a0_3701, \26979 );
not \U$18461 ( \26981 , RIdbfc9a0_3701);
not \U$18462 ( \26982 , \26981 );
not \U$18463 ( \26983 , \24635 );
and \U$18464 ( \26984 , \26982 , \26983 );
and \U$18465 ( \26985 , \26738 , \24635 );
or \U$18466 ( \26986 , \26984 , \26985 );
and \U$18467 ( \26987 , \26986 , \26661 );
or \U$18468 ( \26988 , \26980 , \26987 );
and \U$18470 ( \26989 , \26988 , 1'b1 );
or \U$18472 ( \26990 , \26989 , 1'b0 );
buf \U$18473 ( \26991 , \26990 );
_DC r253e4_GF_IsGateDCbyConstraint ( \26992_nR253e4 , \26991 , \21944 );
buf \U$18474 ( \26993 , \26992_nR253e4 );
not \U$18475 ( \26994 , \26661 );
and \U$18476 ( \26995 , RIdbfb398_3702, \26994 );
not \U$18477 ( \26996 , RIdbfb398_3702);
not \U$18478 ( \26997 , \26996 );
not \U$18479 ( \26998 , \24635 );
and \U$18480 ( \26999 , \26997 , \26998 );
and \U$18481 ( \27000 , \26755 , \24635 );
or \U$18482 ( \27001 , \26999 , \27000 );
and \U$18483 ( \27002 , \27001 , \26661 );
or \U$18484 ( \27003 , \26995 , \27002 );
and \U$18486 ( \27004 , \27003 , 1'b1 );
or \U$18488 ( \27005 , \27004 , 1'b0 );
buf \U$18489 ( \27006 , \27005 );
_DC r253e6_GF_IsGateDCbyConstraint ( \27007_nR253e6 , \27006 , \21944 );
buf \U$18490 ( \27008 , \27007_nR253e6 );
not \U$18491 ( \27009 , \26661 );
and \U$18492 ( \27010 , RIdbfa240_3703, \27009 );
not \U$18493 ( \27011 , RIdbfa240_3703);
not \U$18494 ( \27012 , \27011 );
not \U$18495 ( \27013 , \24635 );
and \U$18496 ( \27014 , \27012 , \27013 );
and \U$18497 ( \27015 , \26772 , \24635 );
or \U$18498 ( \27016 , \27014 , \27015 );
and \U$18499 ( \27017 , \27016 , \26661 );
or \U$18500 ( \27018 , \27010 , \27017 );
and \U$18502 ( \27019 , \27018 , 1'b1 );
or \U$18504 ( \27020 , \27019 , 1'b0 );
buf \U$18505 ( \27021 , \27020 );
_DC r253e8_GF_IsGateDCbyConstraint ( \27022_nR253e8 , \27021 , \21944 );
buf \U$18506 ( \27023 , \27022_nR253e8 );
not \U$18507 ( \27024 , \26661 );
and \U$18508 ( \27025 , RIdbf8c38_3704, \27024 );
not \U$18509 ( \27026 , RIdbf8c38_3704);
not \U$18510 ( \27027 , \27026 );
not \U$18511 ( \27028 , \24635 );
and \U$18512 ( \27029 , \27027 , \27028 );
and \U$18513 ( \27030 , \26789 , \24635 );
or \U$18514 ( \27031 , \27029 , \27030 );
and \U$18515 ( \27032 , \27031 , \26661 );
or \U$18516 ( \27033 , \27025 , \27032 );
and \U$18518 ( \27034 , \27033 , 1'b1 );
or \U$18520 ( \27035 , \27034 , 1'b0 );
buf \U$18521 ( \27036 , \27035 );
_DC r253ea_GF_IsGateDCbyConstraint ( \27037_nR253ea , \27036 , \21944 );
buf \U$18522 ( \27038 , \27037_nR253ea );
not \U$18523 ( \27039 , \26679 );
and \U$18524 ( \27040 , RIdbf7ae0_3705, \27039 );
not \U$18525 ( \27041 , RIdbf7ae0_3705);
not \U$18526 ( \27042 , \27041 );
not \U$18527 ( \27043 , \25748 );
and \U$18528 ( \27044 , \27042 , \27043 );
and \U$18529 ( \27045 , \26669 , \25748 );
or \U$18530 ( \27046 , \27044 , \27045 );
and \U$18531 ( \27047 , \27046 , \26679 );
or \U$18532 ( \27048 , \27040 , \27047 );
and \U$18534 ( \27049 , \27048 , 1'b1 );
or \U$18536 ( \27050 , \27049 , 1'b0 );
buf \U$18537 ( \27051 , \27050 );
_DC r253ec_GF_IsGateDCbyConstraint ( \27052_nR253ec , \27051 , \21944 );
buf \U$18538 ( \27053 , \27052_nR253ec );
not \U$18539 ( \27054 , \26679 );
and \U$18540 ( \27055 , RIdbf6988_3706, \27054 );
not \U$18541 ( \27056 , RIdbf6988_3706);
not \U$18542 ( \27057 , \27056 );
not \U$18543 ( \27058 , \25748 );
and \U$18544 ( \27059 , \27057 , \27058 );
and \U$18545 ( \27060 , \26687 , \25748 );
or \U$18546 ( \27061 , \27059 , \27060 );
and \U$18547 ( \27062 , \27061 , \26679 );
or \U$18548 ( \27063 , \27055 , \27062 );
and \U$18550 ( \27064 , \27063 , 1'b1 );
or \U$18552 ( \27065 , \27064 , 1'b0 );
buf \U$18553 ( \27066 , \27065 );
_DC r253ee_GF_IsGateDCbyConstraint ( \27067_nR253ee , \27066 , \21944 );
buf \U$18554 ( \27068 , \27067_nR253ee );
not \U$18555 ( \27069 , \26679 );
and \U$18556 ( \27070 , RIdbf5380_3707, \27069 );
not \U$18557 ( \27071 , RIdbf5380_3707);
not \U$18558 ( \27072 , \27071 );
not \U$18559 ( \27073 , \25748 );
and \U$18560 ( \27074 , \27072 , \27073 );
and \U$18561 ( \27075 , \26704 , \25748 );
or \U$18562 ( \27076 , \27074 , \27075 );
and \U$18563 ( \27077 , \27076 , \26679 );
or \U$18564 ( \27078 , \27070 , \27077 );
and \U$18566 ( \27079 , \27078 , 1'b1 );
or \U$18568 ( \27080 , \27079 , 1'b0 );
buf \U$18569 ( \27081 , \27080 );
_DC r253f0_GF_IsGateDCbyConstraint ( \27082_nR253f0 , \27081 , \21944 );
buf \U$18570 ( \27083 , \27082_nR253f0 );
not \U$18571 ( \27084 , \26679 );
and \U$18572 ( \27085 , RIdbf4228_3708, \27084 );
not \U$18573 ( \27086 , RIdbf4228_3708);
not \U$18574 ( \27087 , \27086 );
not \U$18575 ( \27088 , \25748 );
and \U$18576 ( \27089 , \27087 , \27088 );
and \U$18577 ( \27090 , \26721 , \25748 );
or \U$18578 ( \27091 , \27089 , \27090 );
and \U$18579 ( \27092 , \27091 , \26679 );
or \U$18580 ( \27093 , \27085 , \27092 );
and \U$18582 ( \27094 , \27093 , 1'b1 );
or \U$18584 ( \27095 , \27094 , 1'b0 );
buf \U$18585 ( \27096 , \27095 );
_DC r253f2_GF_IsGateDCbyConstraint ( \27097_nR253f2 , \27096 , \21944 );
buf \U$18586 ( \27098 , \27097_nR253f2 );
not \U$18587 ( \27099 , \26679 );
and \U$18588 ( \27100 , RIdbf2c20_3709, \27099 );
not \U$18589 ( \27101 , RIdbf2c20_3709);
not \U$18590 ( \27102 , \27101 );
not \U$18591 ( \27103 , \25748 );
and \U$18592 ( \27104 , \27102 , \27103 );
and \U$18593 ( \27105 , \26738 , \25748 );
or \U$18594 ( \27106 , \27104 , \27105 );
and \U$18595 ( \27107 , \27106 , \26679 );
or \U$18596 ( \27108 , \27100 , \27107 );
and \U$18598 ( \27109 , \27108 , 1'b1 );
or \U$18600 ( \27110 , \27109 , 1'b0 );
buf \U$18601 ( \27111 , \27110 );
_DC r253f4_GF_IsGateDCbyConstraint ( \27112_nR253f4 , \27111 , \21944 );
buf \U$18602 ( \27113 , \27112_nR253f4 );
not \U$18603 ( \27114 , \26679 );
and \U$18604 ( \27115 , RIdbf1ac8_3710, \27114 );
not \U$18605 ( \27116 , RIdbf1ac8_3710);
not \U$18606 ( \27117 , \27116 );
not \U$18607 ( \27118 , \25748 );
and \U$18608 ( \27119 , \27117 , \27118 );
and \U$18609 ( \27120 , \26755 , \25748 );
or \U$18610 ( \27121 , \27119 , \27120 );
and \U$18611 ( \27122 , \27121 , \26679 );
or \U$18612 ( \27123 , \27115 , \27122 );
and \U$18614 ( \27124 , \27123 , 1'b1 );
or \U$18616 ( \27125 , \27124 , 1'b0 );
buf \U$18617 ( \27126 , \27125 );
_DC r253f6_GF_IsGateDCbyConstraint ( \27127_nR253f6 , \27126 , \21944 );
buf \U$18618 ( \27128 , \27127_nR253f6 );
not \U$18619 ( \27129 , \26679 );
and \U$18620 ( \27130 , RIdbf04c0_3711, \27129 );
not \U$18621 ( \27131 , RIdbf04c0_3711);
not \U$18622 ( \27132 , \27131 );
not \U$18623 ( \27133 , \25748 );
and \U$18624 ( \27134 , \27132 , \27133 );
and \U$18625 ( \27135 , \26772 , \25748 );
or \U$18626 ( \27136 , \27134 , \27135 );
and \U$18627 ( \27137 , \27136 , \26679 );
or \U$18628 ( \27138 , \27130 , \27137 );
and \U$18630 ( \27139 , \27138 , 1'b1 );
or \U$18632 ( \27140 , \27139 , 1'b0 );
buf \U$18633 ( \27141 , \27140 );
_DC r253f8_GF_IsGateDCbyConstraint ( \27142_nR253f8 , \27141 , \21944 );
buf \U$18634 ( \27143 , \27142_nR253f8 );
not \U$18635 ( \27144 , \26679 );
and \U$18636 ( \27145 , RIdbef368_3712, \27144 );
not \U$18637 ( \27146 , RIdbef368_3712);
not \U$18638 ( \27147 , \27146 );
not \U$18639 ( \27148 , \25748 );
and \U$18640 ( \27149 , \27147 , \27148 );
and \U$18641 ( \27150 , \26789 , \25748 );
or \U$18642 ( \27151 , \27149 , \27150 );
and \U$18643 ( \27152 , \27151 , \26679 );
or \U$18644 ( \27153 , \27145 , \27152 );
and \U$18646 ( \27154 , \27153 , 1'b1 );
or \U$18648 ( \27155 , \27154 , 1'b0 );
buf \U$18649 ( \27156 , \27155 );
_DC r253fa_GF_IsGateDCbyConstraint ( \27157_nR253fa , \27156 , \21944 );
buf \U$18650 ( \27158 , \27157_nR253fa );
nand \U$18651 ( \27159 , RIb79b428_272, \21694 );
or \U$18652 ( \27160 , \21458 , \27159 );
not \U$18653 ( \27161 , \10986 );
and \U$18654 ( \27162 , \27160 , \27161 );
not \U$18655 ( \27163 , \21814 );
buf \U$18656 ( \27164 , RIb8396e0_155);
not \U$18657 ( \27165 , \27164 );
not \U$18658 ( \27166 , \21809 );
not \U$18659 ( \27167 , \27166 );
or \U$18660 ( \27168 , \27165 , \27167 );
not \U$18661 ( \27169 , \27168 );
and \U$18662 ( \27170 , \27163 , \27169 );
nor \U$18663 ( \27171 , \27162 , \27170 );
and \U$18665 ( \27172 , \27171 , 1'b1 );
or \U$18667 ( \27173 , \27172 , 1'b0 );
_DC r25666_GF_IsGateDCbyConstraint ( \27174_nR25666 , \27173 , \21944 );
buf \U$18668 ( \27175 , \27174_nR25666 );
buf \U$18669 ( \27176 , RIdda31a8_3581);
not \U$18670 ( \27177 , \27176 );
nand \U$18671 ( \27178 , \21455 , \21360 );
not \U$18672 ( \27179 , \27178 );
not \U$18673 ( \27180 , \27179 );
or \U$18674 ( \27181 , \21275 , \27180 );
or \U$18675 ( \27182 , \27177 , \27181 );
buf \U$18676 ( \27183 , RIdbd9c48_3186);
not \U$18677 ( \27184 , \27183 );
not \U$18678 ( \27185 , \21273 );
not \U$18679 ( \27186 , \27185 );
or \U$18680 ( \27187 , \21172 , \27186 );
not \U$18681 ( \27188 , \21455 );
nand \U$18682 ( \27189 , \21361 , \27188 );
not \U$18683 ( \27190 , \27189 );
not \U$18684 ( \27191 , \27190 );
or \U$18685 ( \27192 , \27187 , \27191 );
or \U$18686 ( \27193 , \27184 , \27192 );
nand \U$18687 ( \27194 , \27182 , \27193 );
buf \U$18688 ( \27195 , RIe036f80_4371);
not \U$18689 ( \27196 , \27195 );
nand \U$18690 ( \27197 , \27188 , \21360 );
not \U$18691 ( \27198 , \27197 );
not \U$18692 ( \27199 , \27198 );
or \U$18693 ( \27200 , \21275 , \27199 );
or \U$18694 ( \27201 , \27196 , \27200 );
buf \U$18695 ( \27202 , RIe100460_4766);
not \U$18696 ( \27203 , \27202 );
not \U$18697 ( \27204 , \27190 );
or \U$18698 ( \27205 , \21275 , \27204 );
or \U$18699 ( \27206 , \27203 , \27205 );
nand \U$18700 ( \27207 , \27201 , \27206 );
nor \U$18701 ( \27208 , \27194 , \27207 );
buf \U$18702 ( \27209 , RIda3bc30_2396);
not \U$18703 ( \27210 , \27209 );
not \U$18704 ( \27211 , \21456 );
or \U$18705 ( \27212 , \27187 , \27211 );
or \U$18706 ( \27213 , \27210 , \27212 );
buf \U$18707 ( \27214 , RIde6b9c8_3976);
not \U$18708 ( \27215 , \27214 );
or \U$18709 ( \27216 , \27215 , \21458 );
nand \U$18710 ( \27217 , \27213 , \27216 );
buf \U$18711 ( \27218 , RIdb0e968_2791);
not \U$18712 ( \27219 , \27218 );
or \U$18713 ( \27220 , \27187 , \27197 );
or \U$18714 ( \27221 , \27219 , \27220 );
buf \U$18715 ( \27222 , RId987e10_2001);
not \U$18716 ( \27223 , \27222 );
not \U$18717 ( \27224 , \27179 );
or \U$18718 ( \27225 , \27187 , \27224 );
or \U$18719 ( \27226 , \27223 , \27225 );
nand \U$18720 ( \27227 , \27221 , \27226 );
nor \U$18721 ( \27228 , \27217 , \27227 );
not \U$18722 ( \27229 , \27185 );
or \U$18723 ( \27230 , \21173 , \27229 );
or \U$18724 ( \27231 , \27230 , \27189 );
not \U$18725 ( \27232 , \27231 );
buf \U$18726 ( \27233 , RIe527288_6346);
and \U$18727 ( \27234 , \27232 , \27233 );
buf \U$18728 ( \27235 , RIe45e528_5951);
not \U$18729 ( \27236 , \27198 );
or \U$18730 ( \27237 , \27230 , \27236 );
not \U$18731 ( \27238 , \27237 );
and \U$18732 ( \27239 , \27235 , \27238 );
nor \U$18733 ( \27240 , \27234 , \27239 );
not \U$18734 ( \27241 , \21456 );
or \U$18735 ( \27242 , \27230 , \27241 );
not \U$18736 ( \27243 , \27242 );
buf \U$18737 ( \27244 , RIe395df8_5556);
and \U$18738 ( \27245 , \27243 , \27244 );
buf \U$18739 ( \27246 , RIe1ca840_5161);
or \U$18740 ( \27247 , \27230 , \27178 );
not \U$18741 ( \27248 , \27247 );
and \U$18742 ( \27249 , \27246 , \27248 );
nor \U$18743 ( \27250 , \27245 , \27249 );
nand \U$18744 ( \27251 , \27240 , \27250 );
not \U$18745 ( \27252 , \27251 );
not \U$18746 ( \27253 , \21273 );
or \U$18747 ( \27254 , \21172 , \27253 );
not \U$18748 ( \27255 , \21456 );
or \U$18749 ( \27256 , \27254 , \27255 );
not \U$18750 ( \27257 , \27256 );
buf \U$18751 ( \27258 , RId72b4a8_816);
and \U$18752 ( \27259 , \27257 , \27258 );
buf \U$18753 ( \27260 , RIe5efc28_6741);
not \U$18754 ( \27261 , \27179 );
or \U$18755 ( \27262 , \27254 , \27261 );
not \U$18756 ( \27263 , \27262 );
and \U$18757 ( \27264 , \27260 , \27263 );
nor \U$18758 ( \27265 , \27259 , \27264 );
not \U$18759 ( \27266 , \27190 );
or \U$18760 ( \27267 , \27254 , \27266 );
not \U$18761 ( \27268 , \27267 );
buf \U$18762 ( \27269 , RId8bc950_1606);
and \U$18763 ( \27270 , \27268 , \27269 );
buf \U$18764 ( \27271 , RId7f4028_1211);
not \U$18765 ( \27272 , \27198 );
or \U$18766 ( \27273 , \27254 , \27272 );
not \U$18767 ( \27274 , \27273 );
and \U$18768 ( \27275 , \27271 , \27274 );
nor \U$18769 ( \27276 , \27270 , \27275 );
and \U$18770 ( \27277 , \27252 , \27265 , \27276 );
nand \U$18771 ( \27278 , \27208 , \27228 , \27277 );
_DC r22c68_GF_IsGateDCbyConstraint ( \27279_nR22c68 , \27278 , \21944 );
buf \U$18772 ( \27280 , \27279_nR22c68 );
buf \U$18773 ( \27281 , RId710748_846);
not \U$18774 ( \27282 , \27281 );
or \U$18775 ( \27283 , \27256 , \27282 );
buf \U$18776 ( \27284 , RId96d278_2032);
not \U$18777 ( \27285 , \27284 );
or \U$18778 ( \27286 , \27225 , \27285 );
nand \U$18779 ( \27287 , \27283 , \27286 );
buf \U$18780 ( \27288 , RId8aa728_1632);
not \U$18781 ( \27289 , \27288 );
or \U$18782 ( \27290 , \27267 , \27289 );
buf \U$18783 ( \27291 , RId7dcb80_1235);
not \U$18784 ( \27292 , \27291 );
or \U$18785 ( \27293 , \27273 , \27292 );
nand \U$18786 ( \27294 , \27290 , \27293 );
nor \U$18787 ( \27295 , \27287 , \27294 );
buf \U$18788 ( \27296 , RIdbc4870_3212);
not \U$18789 ( \27297 , \27296 );
or \U$18790 ( \27298 , \27192 , \27297 );
buf \U$18791 ( \27299 , RIdd8ba30_3609);
not \U$18792 ( \27300 , \27299 );
or \U$18793 ( \27301 , \27181 , \27300 );
nand \U$18794 ( \27302 , \27298 , \27301 );
buf \U$18795 ( \27303 , RIda25c28_2423);
not \U$18796 ( \27304 , \27303 );
or \U$18797 ( \27305 , \27212 , \27304 );
buf \U$18798 ( \27306 , RIdaf5f30_2820);
not \U$18799 ( \27307 , \27306 );
or \U$18800 ( \27308 , \27220 , \27307 );
nand \U$18801 ( \27309 , \27305 , \27308 );
nor \U$18802 ( \27310 , \27302 , \27309 );
nand \U$18803 ( \27311 , \27295 , \27310 );
not \U$18804 ( \27312 , \27311 );
buf \U$18805 ( \27313 , RIe022a30_4393);
not \U$18806 ( \27314 , \27313 );
or \U$18807 ( \27315 , \27200 , \27314 );
buf \U$18808 ( \27316 , RIe0e8ec8_4791);
not \U$18809 ( \27317 , \27316 );
or \U$18810 ( \27318 , \27205 , \27317 );
nand \U$18811 ( \27319 , \27315 , \27318 );
buf \U$18812 ( \27320 , RIe1ac2a0_5191);
not \U$18813 ( \27321 , \27320 );
or \U$18814 ( \27322 , \27247 , \27321 );
buf \U$18815 ( \27323 , RIde4ec88_4006);
not \U$18816 ( \27324 , \27323 );
or \U$18817 ( \27325 , \21458 , \27324 );
nand \U$18818 ( \27326 , \27322 , \27325 );
nor \U$18819 ( \27327 , \27319 , \27326 );
buf \U$18820 ( \27328 , RIe444fb0_5975);
not \U$18821 ( \27329 , \27328 );
or \U$18822 ( \27330 , \27237 , \27329 );
buf \U$18823 ( \27331 , RIe37f9b8_5584);
not \U$18824 ( \27332 , \27331 );
or \U$18825 ( \27333 , \27242 , \27332 );
nand \U$18826 ( \27334 , \27330 , \27333 );
buf \U$18827 ( \27335 , RIe5d6d40_6768);
not \U$18828 ( \27336 , \27335 );
or \U$18829 ( \27337 , \27262 , \27336 );
buf \U$18830 ( \27338 , RIe5117a8_6369);
not \U$18831 ( \27339 , \27338 );
or \U$18832 ( \27340 , \27231 , \27339 );
nand \U$18833 ( \27341 , \27337 , \27340 );
nor \U$18834 ( \27342 , \27334 , \27341 );
and \U$18835 ( \27343 , \27312 , \27327 , \27342 );
_DC r22c59_GF_IsGateDCbyConstraint ( \27344_nR22c59 , \27343 , \21944 );
buf \U$18836 ( \27345 , \27344_nR22c59 );
nor \U$18837 ( \27346 , \21812 , \21810 );
nand \U$18838 ( \27347 , RIe546098_6850, \27346 );
nor \U$18839 ( \27348 , \21809 , \27347 );
buf \U$18840 ( \27349 , \27348 );
buf \U$18841 ( \27350 , \27349 );
not \U$18842 ( \27351 , \22095 );
buf \U$18843 ( \27352 , \27351 );
buf \U$18844 ( \27353 , \27352 );
nand \U$18845 ( \27354 , \27350 , \27353 );
buf \U$18846 ( \27355 , RIb79b518_270);
buf \U$18847 ( \27356 , \27355 );
buf \U$18848 ( \27357 , \27356 );
not \U$18849 ( \27358 , \27231 );
and \U$18850 ( \27359 , \27358 , \21694 );
buf \U$18851 ( \27360 , \27359 );
buf \U$18852 ( \27361 , \27360 );
nand \U$18853 ( \27362 , \27357 , \27361 );
nand \U$18854 ( \27363 , \27354 , \27362 );
buf \U$18855 ( \27364 , \27363 );
buf \U$18856 ( \27365 , \27364 );
not \U$18857 ( \27366 , \27365 );
and \U$18858 ( \27367 , RIe3ac2b0_6083, \27366 );
not \U$18859 ( \27368 , RIe3ac2b0_6083);
buf \U$18860 ( \27369 , RIe667bb0_6885);
buf \U$18861 ( \27370 , \27369 );
buf \U$18862 ( \27371 , RIe667f70_6886);
buf \U$18863 ( \27372 , \27371 );
not \U$18864 ( \27373 , \27372 );
not \U$18865 ( \27374 , \27373 );
or \U$18866 ( \27375 , \27370 , \27374 );
not \U$18867 ( \27376 , \27375 );
nand \U$18868 ( \27377 , \27362 , \27376 );
not \U$18869 ( \27378 , RIea91768_6889);
not \U$18870 ( \27379 , \27378 );
buf \U$18871 ( \27380 , \27379 );
not \U$18872 ( \27381 , \27380 );
not \U$18873 ( \27382 , \22119 );
buf \U$18874 ( \27383 , \27382 );
not \U$18875 ( \27384 , \27383 );
not \U$18876 ( \27385 , \27362 );
and \U$18877 ( \27386 , \27381 , \27384 , \27385 );
not \U$18878 ( \27387 , \27386 );
and \U$18879 ( \27388 , \27377 , \27387 );
not \U$18880 ( \27389 , \27388 );
or \U$18881 ( \27390 , \27368 , \27389 );
not \U$18882 ( \27391 , \27377 );
buf \U$18883 ( \27392 , \27391 );
buf \U$18884 ( \27393 , \22131 );
and \U$18885 ( \27394 , \27392 , \27393 );
buf \U$18886 ( \27395 , RIb7c5980_237);
not \U$18887 ( \27396 , \27380 );
not \U$18888 ( \27397 , \27383 );
and \U$18889 ( \27398 , \27396 , \27397 , \27385 );
not \U$18890 ( \27399 , \27398 );
buf \U$18891 ( \27400 , \27399 );
not \U$18892 ( \27401 , \27400 );
and \U$18893 ( \27402 , \27395 , \27401 );
nor \U$18894 ( \27403 , \27394 , \27402 );
nand \U$18895 ( \27404 , \27390 , \27403 );
and \U$18896 ( \27405 , \27404 , \27365 );
or \U$18897 ( \27406 , \27367 , \27405 );
and \U$18899 ( \27407 , \27406 , 1'b1 );
or \U$18901 ( \27408 , \27407 , 1'b0 );
buf \U$18902 ( \27409 , \27408 );
_DC r23ca4_GF_IsGateDCbyConstraint ( \27410_nR23ca4 , \27409 , \21944 );
buf \U$18903 ( \27411 , \27410_nR23ca4 );
not \U$18904 ( \27412 , \27365 );
and \U$18905 ( \27413 , RIe3aaca8_6084, \27412 );
not \U$18906 ( \27414 , RIe3aaca8_6084);
not \U$18907 ( \27415 , \27380 );
not \U$18908 ( \27416 , \27383 );
and \U$18909 ( \27417 , \27415 , \27416 , \27385 );
not \U$18910 ( \27418 , \27417 );
buf \U$18911 ( \27419 , \27418 );
and \U$18912 ( \27420 , \27377 , \27419 );
not \U$18913 ( \27421 , \27420 );
or \U$18914 ( \27422 , \27414 , \27421 );
buf \U$18915 ( \27423 , \27391 );
buf \U$18916 ( \27424 , RIb87eb78_68);
and \U$18917 ( \27425 , \27423 , \27424 );
buf \U$18918 ( \27426 , RIb7c59f8_236);
buf \U$18919 ( \27427 , \27426 );
buf \U$18920 ( \27428 , \27399 );
not \U$18921 ( \27429 , \27428 );
and \U$18922 ( \27430 , \27427 , \27429 );
nor \U$18923 ( \27431 , \27425 , \27430 );
nand \U$18924 ( \27432 , \27422 , \27431 );
and \U$18925 ( \27433 , \27432 , \27365 );
or \U$18926 ( \27434 , \27413 , \27433 );
and \U$18928 ( \27435 , \27434 , 1'b1 );
or \U$18930 ( \27436 , \27435 , 1'b0 );
buf \U$18931 ( \27437 , \27436 );
_DC r23cba_GF_IsGateDCbyConstraint ( \27438_nR23cba , \27437 , \21944 );
buf \U$18932 ( \27439 , \27438_nR23cba );
not \U$18933 ( \27440 , \27365 );
and \U$18934 ( \27441 , RIe3a9b50_6085, \27440 );
not \U$18935 ( \27442 , RIe3a9b50_6085);
or \U$18936 ( \27443 , \27442 , \27389 );
buf \U$18937 ( \27444 , \22179 );
and \U$18938 ( \27445 , \27423 , \27444 );
buf \U$18939 ( \27446 , RIb7c5a70_235);
not \U$18940 ( \27447 , \27400 );
and \U$18941 ( \27448 , \27446 , \27447 );
nor \U$18942 ( \27449 , \27445 , \27448 );
nand \U$18943 ( \27450 , \27443 , \27449 );
and \U$18944 ( \27451 , \27450 , \27365 );
or \U$18945 ( \27452 , \27441 , \27451 );
and \U$18947 ( \27453 , \27452 , 1'b1 );
or \U$18949 ( \27454 , \27453 , 1'b0 );
buf \U$18950 ( \27455 , \27454 );
_DC r23cd0_GF_IsGateDCbyConstraint ( \27456_nR23cd0 , \27455 , \21944 );
buf \U$18951 ( \27457 , \27456_nR23cd0 );
buf \U$18952 ( \27458 , \27363 );
buf \U$18953 ( \27459 , \27458 );
not \U$18954 ( \27460 , \27459 );
and \U$18955 ( \27461 , RIe3a8548_6086, \27460 );
not \U$18956 ( \27462 , RIe3a8548_6086);
or \U$18957 ( \27463 , \27462 , \27421 );
buf \U$18958 ( \27464 , \27391 );
buf \U$18959 ( \27465 , \22202 );
and \U$18960 ( \27466 , \27464 , \27465 );
buf \U$18961 ( \27467 , \22205 );
not \U$18962 ( \27468 , \27419 );
and \U$18963 ( \27469 , \27467 , \27468 );
nor \U$18964 ( \27470 , \27466 , \27469 );
nand \U$18965 ( \27471 , \27463 , \27470 );
and \U$18966 ( \27472 , \27471 , \27459 );
or \U$18967 ( \27473 , \27461 , \27472 );
and \U$18969 ( \27474 , \27473 , 1'b1 );
or \U$18971 ( \27475 , \27474 , 1'b0 );
buf \U$18972 ( \27476 , \27475 );
_DC r23ce6_GF_IsGateDCbyConstraint ( \27477_nR23ce6 , \27476 , \21944 );
buf \U$18973 ( \27478 , \27477_nR23ce6 );
not \U$18974 ( \27479 , \27459 );
and \U$18975 ( \27480 , RIe3a73f0_6087, \27479 );
not \U$18976 ( \27481 , RIe3a73f0_6087);
not \U$18977 ( \27482 , \27388 );
or \U$18978 ( \27483 , \27481 , \27482 );
buf \U$18979 ( \27484 , \22223 );
and \U$18980 ( \27485 , \27392 , \27484 );
buf \U$18981 ( \27486 , RIb7cae58_233);
buf \U$18982 ( \27487 , \27418 );
not \U$18983 ( \27488 , \27487 );
and \U$18984 ( \27489 , \27486 , \27488 );
nor \U$18985 ( \27490 , \27485 , \27489 );
nand \U$18986 ( \27491 , \27483 , \27490 );
and \U$18987 ( \27492 , \27491 , \27459 );
or \U$18988 ( \27493 , \27480 , \27492 );
and \U$18990 ( \27494 , \27493 , 1'b1 );
or \U$18992 ( \27495 , \27494 , 1'b0 );
buf \U$18993 ( \27496 , \27495 );
_DC r23cfc_GF_IsGateDCbyConstraint ( \27497_nR23cfc , \27496 , \21944 );
buf \U$18994 ( \27498 , \27497_nR23cfc );
not \U$18995 ( \27499 , \27365 );
and \U$18996 ( \27500 , RIe3a6298_6088, \27499 );
not \U$18997 ( \27501 , RIe3a6298_6088);
not \U$18998 ( \27502 , \27420 );
or \U$18999 ( \27503 , \27501 , \27502 );
buf \U$19000 ( \27504 , \22245 );
and \U$19001 ( \27505 , \27464 , \27504 );
buf \U$19002 ( \27506 , RIb7caed0_232);
buf \U$19003 ( \27507 , \27506 );
buf \U$19004 ( \27508 , \27399 );
not \U$19005 ( \27509 , \27508 );
and \U$19006 ( \27510 , \27507 , \27509 );
nor \U$19007 ( \27511 , \27505 , \27510 );
nand \U$19008 ( \27512 , \27503 , \27511 );
and \U$19009 ( \27513 , \27512 , \27365 );
or \U$19010 ( \27514 , \27500 , \27513 );
and \U$19012 ( \27515 , \27514 , 1'b1 );
or \U$19014 ( \27516 , \27515 , 1'b0 );
buf \U$19015 ( \27517 , \27516 );
_DC r23d12_GF_IsGateDCbyConstraint ( \27518_nR23d12 , \27517 , \21944 );
buf \U$19016 ( \27519 , \27518_nR23d12 );
not \U$19017 ( \27520 , \27365 );
and \U$19018 ( \27521 , RIe3a4c90_6089, \27520 );
not \U$19019 ( \27522 , RIe3a4c90_6089);
not \U$19020 ( \27523 , \27388 );
or \U$19021 ( \27524 , \27522 , \27523 );
buf \U$19022 ( \27525 , \22271 );
and \U$19023 ( \27526 , \27392 , \27525 );
buf \U$19024 ( \27527 , RIb7caf48_231);
not \U$19025 ( \27528 , \27419 );
and \U$19026 ( \27529 , \27527 , \27528 );
nor \U$19027 ( \27530 , \27526 , \27529 );
nand \U$19028 ( \27531 , \27524 , \27530 );
and \U$19029 ( \27532 , \27531 , \27365 );
or \U$19030 ( \27533 , \27521 , \27532 );
and \U$19032 ( \27534 , \27533 , 1'b1 );
or \U$19034 ( \27535 , \27534 , 1'b0 );
buf \U$19035 ( \27536 , \27535 );
_DC r23d1c_GF_IsGateDCbyConstraint ( \27537_nR23d1c , \27536 , \21944 );
buf \U$19036 ( \27538 , \27537_nR23d1c );
not \U$19037 ( \27539 , \27365 );
and \U$19038 ( \27540 , RIe3a3b38_6090, \27539 );
not \U$19039 ( \27541 , RIe3a3b38_6090);
or \U$19040 ( \27542 , \27541 , \27421 );
buf \U$19041 ( \27543 , RIb885478_62);
and \U$19042 ( \27544 , \27464 , \27543 );
buf \U$19043 ( \27545 , RIb7cafc0_230);
buf \U$19044 ( \27546 , \27545 );
not \U$19045 ( \27547 , \27428 );
and \U$19046 ( \27548 , \27546 , \27547 );
nor \U$19047 ( \27549 , \27544 , \27548 );
nand \U$19048 ( \27550 , \27542 , \27549 );
and \U$19049 ( \27551 , \27550 , \27365 );
or \U$19050 ( \27552 , \27540 , \27551 );
and \U$19052 ( \27553 , \27552 , 1'b1 );
or \U$19054 ( \27554 , \27553 , 1'b0 );
buf \U$19055 ( \27555 , \27554 );
_DC r23d1e_GF_IsGateDCbyConstraint ( \27556_nR23d1e , \27555 , \21944 );
buf \U$19056 ( \27557 , \27556_nR23d1e );
buf \U$19057 ( \27558 , \27364 );
not \U$19058 ( \27559 , \27558 );
and \U$19059 ( \27560 , RIe3a2530_6091, \27559 );
not \U$19060 ( \27561 , RIe3a2530_6091);
not \U$19061 ( \27562 , \27420 );
or \U$19062 ( \27563 , \27561 , \27562 );
buf \U$19063 ( \27564 , RIb8854f0_61);
buf \U$19064 ( \27565 , \27564 );
and \U$19065 ( \27566 , \27464 , \27565 );
buf \U$19066 ( \27567 , RIb7cb038_229);
buf \U$19067 ( \27568 , \27567 );
not \U$19068 ( \27569 , \27400 );
and \U$19069 ( \27570 , \27568 , \27569 );
nor \U$19070 ( \27571 , \27566 , \27570 );
nand \U$19071 ( \27572 , \27563 , \27571 );
and \U$19072 ( \27573 , \27572 , \27558 );
or \U$19073 ( \27574 , \27560 , \27573 );
and \U$19075 ( \27575 , \27574 , 1'b1 );
or \U$19077 ( \27576 , \27575 , 1'b0 );
buf \U$19078 ( \27577 , \27576 );
_DC r23d20_GF_IsGateDCbyConstraint ( \27578_nR23d20 , \27577 , \21944 );
buf \U$19079 ( \27579 , \27578_nR23d20 );
not \U$19080 ( \27580 , \27459 );
and \U$19081 ( \27581 , RIe3a13d8_6092, \27580 );
not \U$19082 ( \27582 , RIe3a13d8_6092);
not \U$19083 ( \27583 , \27420 );
or \U$19084 ( \27584 , \27582 , \27583 );
buf \U$19085 ( \27585 , \22334 );
and \U$19086 ( \27586 , \27392 , \27585 );
buf \U$19087 ( \27587 , RIb7cb0b0_228);
buf \U$19088 ( \27588 , \27587 );
buf \U$19089 ( \27589 , \27418 );
not \U$19090 ( \27590 , \27589 );
and \U$19091 ( \27591 , \27588 , \27590 );
nor \U$19092 ( \27592 , \27586 , \27591 );
nand \U$19093 ( \27593 , \27584 , \27592 );
and \U$19094 ( \27594 , \27593 , \27459 );
or \U$19095 ( \27595 , \27581 , \27594 );
and \U$19097 ( \27596 , \27595 , 1'b1 );
or \U$19099 ( \27597 , \27596 , 1'b0 );
buf \U$19100 ( \27598 , \27597 );
_DC r23d22_GF_IsGateDCbyConstraint ( \27599_nR23d22 , \27598 , \21944 );
buf \U$19101 ( \27600 , \27599_nR23d22 );
not \U$19102 ( \27601 , \27365 );
and \U$19103 ( \27602 , RIe39fdd0_6093, \27601 );
not \U$19104 ( \27603 , RIe39fdd0_6093);
not \U$19105 ( \27604 , \27388 );
or \U$19106 ( \27605 , \27603 , \27604 );
buf \U$19107 ( \27606 , RIb8855e0_59);
and \U$19108 ( \27607 , \27464 , \27606 );
buf \U$19109 ( \27608 , RIb7cb128_227);
buf \U$19110 ( \27609 , \27608 );
not \U$19111 ( \27610 , \27508 );
and \U$19112 ( \27611 , \27609 , \27610 );
nor \U$19113 ( \27612 , \27607 , \27611 );
nand \U$19114 ( \27613 , \27605 , \27612 );
and \U$19115 ( \27614 , \27613 , \27365 );
or \U$19116 ( \27615 , \27602 , \27614 );
and \U$19118 ( \27616 , \27615 , 1'b1 );
or \U$19120 ( \27617 , \27616 , 1'b0 );
buf \U$19121 ( \27618 , \27617 );
_DC r23ca6_GF_IsGateDCbyConstraint ( \27619_nR23ca6 , \27618 , \21944 );
buf \U$19122 ( \27620 , \27619_nR23ca6 );
not \U$19123 ( \27621 , \27558 );
and \U$19124 ( \27622 , RIe39ec78_6094, \27621 );
not \U$19125 ( \27623 , RIe39ec78_6094);
or \U$19126 ( \27624 , \27623 , \27482 );
buf \U$19127 ( \27625 , \22376 );
and \U$19128 ( \27626 , \27423 , \27625 );
buf \U$19129 ( \27627 , RIb7d00d8_226);
buf \U$19130 ( \27628 , \27627 );
not \U$19131 ( \27629 , \27428 );
and \U$19132 ( \27630 , \27628 , \27629 );
nor \U$19133 ( \27631 , \27626 , \27630 );
nand \U$19134 ( \27632 , \27624 , \27631 );
and \U$19135 ( \27633 , \27632 , \27558 );
or \U$19136 ( \27634 , \27622 , \27633 );
and \U$19138 ( \27635 , \27634 , 1'b1 );
or \U$19140 ( \27636 , \27635 , 1'b0 );
buf \U$19141 ( \27637 , \27636 );
_DC r23ca8_GF_IsGateDCbyConstraint ( \27638_nR23ca8 , \27637 , \21944 );
buf \U$19142 ( \27639 , \27638_nR23ca8 );
not \U$19143 ( \27640 , \27365 );
and \U$19144 ( \27641 , RIe39db20_6095, \27640 );
not \U$19145 ( \27642 , RIe39db20_6095);
not \U$19146 ( \27643 , \27388 );
or \U$19147 ( \27644 , \27642 , \27643 );
buf \U$19148 ( \27645 , RIb8856d0_57);
and \U$19149 ( \27646 , \27423 , \27645 );
buf \U$19150 ( \27647 , RIb8263d8_225);
buf \U$19151 ( \27648 , \27647 );
not \U$19152 ( \27649 , \27400 );
and \U$19153 ( \27650 , \27648 , \27649 );
nor \U$19154 ( \27651 , \27646 , \27650 );
nand \U$19155 ( \27652 , \27644 , \27651 );
and \U$19156 ( \27653 , \27652 , \27365 );
or \U$19157 ( \27654 , \27641 , \27653 );
and \U$19159 ( \27655 , \27654 , 1'b1 );
or \U$19161 ( \27656 , \27655 , 1'b0 );
buf \U$19162 ( \27657 , \27656 );
_DC r23caa_GF_IsGateDCbyConstraint ( \27658_nR23caa , \27657 , \21944 );
buf \U$19163 ( \27659 , \27658_nR23caa );
not \U$19164 ( \27660 , \27365 );
and \U$19165 ( \27661 , RIe39c518_6096, \27660 );
not \U$19166 ( \27662 , RIe39c518_6096);
not \U$19167 ( \27663 , \27420 );
or \U$19168 ( \27664 , \27662 , \27663 );
buf \U$19169 ( \27665 , \22417 );
and \U$19170 ( \27666 , \27423 , \27665 );
buf \U$19171 ( \27667 , RIb826e28_224);
buf \U$19172 ( \27668 , \27667 );
not \U$19173 ( \27669 , \27487 );
and \U$19174 ( \27670 , \27668 , \27669 );
nor \U$19175 ( \27671 , \27666 , \27670 );
nand \U$19176 ( \27672 , \27664 , \27671 );
and \U$19177 ( \27673 , \27672 , \27365 );
or \U$19178 ( \27674 , \27661 , \27673 );
and \U$19180 ( \27675 , \27674 , 1'b1 );
or \U$19182 ( \27676 , \27675 , 1'b0 );
buf \U$19183 ( \27677 , \27676 );
_DC r23cac_GF_IsGateDCbyConstraint ( \27678_nR23cac , \27677 , \21944 );
buf \U$19184 ( \27679 , \27678_nR23cac );
not \U$19185 ( \27680 , \27558 );
and \U$19186 ( \27681 , RIe1694d8_6097, \27680 );
not \U$19187 ( \27682 , RIe1694d8_6097);
or \U$19188 ( \27683 , \27682 , \27502 );
buf \U$19189 ( \27684 , RIb8857c0_55);
and \U$19190 ( \27685 , \27464 , \27684 );
buf \U$19191 ( \27686 , RIb826ea0_223);
not \U$19192 ( \27687 , \27589 );
and \U$19193 ( \27688 , \27686 , \27687 );
nor \U$19194 ( \27689 , \27685 , \27688 );
nand \U$19195 ( \27690 , \27683 , \27689 );
and \U$19196 ( \27691 , \27690 , \27558 );
or \U$19197 ( \27692 , \27681 , \27691 );
and \U$19199 ( \27693 , \27692 , 1'b1 );
or \U$19201 ( \27694 , \27693 , 1'b0 );
buf \U$19202 ( \27695 , \27694 );
_DC r23cae_GF_IsGateDCbyConstraint ( \27696_nR23cae , \27695 , \21944 );
buf \U$19203 ( \27697 , \27696_nR23cae );
not \U$19204 ( \27698 , \27459 );
and \U$19205 ( \27699 , RIe16e398_6098, \27698 );
not \U$19206 ( \27700 , RIe16e398_6098);
or \U$19207 ( \27701 , \27700 , \27389 );
buf \U$19208 ( \27702 , \22457 );
and \U$19209 ( \27703 , \27391 , \27702 );
buf \U$19210 ( \27704 , \22460 );
not \U$19211 ( \27705 , \27419 );
and \U$19212 ( \27706 , \27704 , \27705 );
nor \U$19213 ( \27707 , \27703 , \27706 );
nand \U$19214 ( \27708 , \27701 , \27707 );
and \U$19215 ( \27709 , \27708 , \27459 );
or \U$19216 ( \27710 , \27699 , \27709 );
and \U$19218 ( \27711 , \27710 , 1'b1 );
or \U$19220 ( \27712 , \27711 , 1'b0 );
buf \U$19221 ( \27713 , \27712 );
_DC r23cb0_GF_IsGateDCbyConstraint ( \27714_nR23cb0 , \27713 , \21944 );
buf \U$19222 ( \27715 , \27714_nR23cb0 );
not \U$19223 ( \27716 , \27459 );
and \U$19224 ( \27717 , RIe173270_6099, \27716 );
not \U$19225 ( \27718 , RIe173270_6099);
or \U$19226 ( \27719 , \27718 , \27604 );
buf \U$19227 ( \27720 , \22477 );
and \U$19228 ( \27721 , \27392 , \27720 );
buf \U$19229 ( \27722 , \22480 );
not \U$19230 ( \27723 , \27589 );
and \U$19231 ( \27724 , \27722 , \27723 );
nor \U$19232 ( \27725 , \27721 , \27724 );
nand \U$19233 ( \27726 , \27719 , \27725 );
and \U$19234 ( \27727 , \27726 , \27459 );
or \U$19235 ( \27728 , \27717 , \27727 );
and \U$19237 ( \27729 , \27728 , 1'b1 );
or \U$19239 ( \27730 , \27729 , 1'b0 );
buf \U$19240 ( \27731 , \27730 );
_DC r23cb2_GF_IsGateDCbyConstraint ( \27732_nR23cb2 , \27731 , \21944 );
buf \U$19241 ( \27733 , \27732_nR23cb2 );
not \U$19242 ( \27734 , \27558 );
and \U$19243 ( \27735 , RIe178388_6100, \27734 );
not \U$19244 ( \27736 , RIe178388_6100);
or \U$19245 ( \27737 , \27736 , \27482 );
buf \U$19246 ( \27738 , RIb885928_52);
and \U$19247 ( \27739 , \27423 , \27738 );
buf \U$19248 ( \27740 , RIb8293a8_220);
buf \U$19249 ( \27741 , \27740 );
not \U$19250 ( \27742 , \27589 );
and \U$19251 ( \27743 , \27741 , \27742 );
nor \U$19252 ( \27744 , \27739 , \27743 );
nand \U$19253 ( \27745 , \27737 , \27744 );
and \U$19254 ( \27746 , \27745 , \27558 );
or \U$19255 ( \27747 , \27735 , \27746 );
and \U$19257 ( \27748 , \27747 , 1'b1 );
or \U$19259 ( \27749 , \27748 , 1'b0 );
buf \U$19260 ( \27750 , \27749 );
_DC r23cb4_GF_IsGateDCbyConstraint ( \27751_nR23cb4 , \27750 , \21944 );
buf \U$19261 ( \27752 , \27751_nR23cb4 );
not \U$19262 ( \27753 , \27459 );
and \U$19263 ( \27754 , RIe17c780_6101, \27753 );
not \U$19264 ( \27755 , RIe17c780_6101);
or \U$19265 ( \27756 , \27755 , \27643 );
buf \U$19266 ( \27757 , RIb8859a0_51);
and \U$19267 ( \27758 , \27423 , \27757 );
buf \U$19268 ( \27759 , RIb829420_219);
buf \U$19269 ( \27760 , \27759 );
not \U$19270 ( \27761 , \27508 );
and \U$19271 ( \27762 , \27760 , \27761 );
nor \U$19272 ( \27763 , \27758 , \27762 );
nand \U$19273 ( \27764 , \27756 , \27763 );
and \U$19274 ( \27765 , \27764 , \27459 );
or \U$19275 ( \27766 , \27754 , \27765 );
and \U$19277 ( \27767 , \27766 , 1'b1 );
or \U$19279 ( \27768 , \27767 , 1'b0 );
buf \U$19280 ( \27769 , \27768 );
_DC r23cb6_GF_IsGateDCbyConstraint ( \27770_nR23cb6 , \27769 , \21944 );
buf \U$19281 ( \27771 , \27770_nR23cb6 );
not \U$19282 ( \27772 , \27365 );
and \U$19283 ( \27773 , RIe1805d8_6102, \27772 );
not \U$19284 ( \27774 , RIe1805d8_6102);
or \U$19285 ( \27775 , \27774 , \27523 );
buf \U$19286 ( \27776 , \22538 );
and \U$19287 ( \27777 , \27423 , \27776 );
buf \U$19288 ( \27778 , RIb829498_218);
buf \U$19289 ( \27779 , \27778 );
not \U$19290 ( \27780 , \27400 );
and \U$19291 ( \27781 , \27779 , \27780 );
nor \U$19292 ( \27782 , \27777 , \27781 );
nand \U$19293 ( \27783 , \27775 , \27782 );
and \U$19294 ( \27784 , \27783 , \27365 );
or \U$19295 ( \27785 , \27773 , \27784 );
and \U$19297 ( \27786 , \27785 , 1'b1 );
or \U$19299 ( \27787 , \27786 , 1'b0 );
buf \U$19300 ( \27788 , \27787 );
_DC r23cb8_GF_IsGateDCbyConstraint ( \27789_nR23cb8 , \27788 , \21944 );
buf \U$19301 ( \27790 , \27789_nR23cb8 );
not \U$19302 ( \27791 , \27558 );
and \U$19303 ( \27792 , RIe1877c0_6103, \27791 );
not \U$19304 ( \27793 , RIe1877c0_6103);
or \U$19305 ( \27794 , \27793 , \27562 );
buf \U$19306 ( \27795 , RIb885a90_49);
buf \U$19307 ( \27796 , \27795 );
and \U$19308 ( \27797 , \27391 , \27796 );
buf \U$19309 ( \27798 , RIb829510_217);
buf \U$19310 ( \27799 , \27798 );
not \U$19311 ( \27800 , \27589 );
and \U$19312 ( \27801 , \27799 , \27800 );
nor \U$19313 ( \27802 , \27797 , \27801 );
nand \U$19314 ( \27803 , \27794 , \27802 );
and \U$19315 ( \27804 , \27803 , \27558 );
or \U$19316 ( \27805 , \27792 , \27804 );
and \U$19318 ( \27806 , \27805 , 1'b1 );
or \U$19320 ( \27807 , \27806 , 1'b0 );
buf \U$19321 ( \27808 , \27807 );
_DC r23cbc_GF_IsGateDCbyConstraint ( \27809_nR23cbc , \27808 , \21944 );
buf \U$19322 ( \27810 , \27809_nR23cbc );
not \U$19323 ( \27811 , \27459 );
and \U$19324 ( \27812 , RIe18c9c8_6104, \27811 );
not \U$19325 ( \27813 , RIe18c9c8_6104);
or \U$19326 ( \27814 , \27813 , \27583 );
buf \U$19327 ( \27815 , \22578 );
and \U$19328 ( \27816 , \27391 , \27815 );
buf \U$19329 ( \27817 , \22581 );
not \U$19330 ( \27818 , \27508 );
and \U$19331 ( \27819 , \27817 , \27818 );
nor \U$19332 ( \27820 , \27816 , \27819 );
nand \U$19333 ( \27821 , \27814 , \27820 );
and \U$19334 ( \27822 , \27821 , \27459 );
or \U$19335 ( \27823 , \27812 , \27822 );
and \U$19337 ( \27824 , \27823 , 1'b1 );
or \U$19339 ( \27825 , \27824 , 1'b0 );
buf \U$19340 ( \27826 , \27825 );
_DC r23cbe_GF_IsGateDCbyConstraint ( \27827_nR23cbe , \27826 , \21944 );
buf \U$19341 ( \27828 , \27827_nR23cbe );
not \U$19342 ( \27829 , \27459 );
and \U$19343 ( \27830 , RIe192ff8_6105, \27829 );
not \U$19344 ( \27831 , RIe192ff8_6105);
or \U$19345 ( \27832 , \27831 , \27523 );
buf \U$19346 ( \27833 , \22598 );
and \U$19347 ( \27834 , \27464 , \27833 );
buf \U$19348 ( \27835 , \22601 );
not \U$19349 ( \27836 , \27428 );
and \U$19350 ( \27837 , \27835 , \27836 );
nor \U$19351 ( \27838 , \27834 , \27837 );
nand \U$19352 ( \27839 , \27832 , \27838 );
and \U$19353 ( \27840 , \27839 , \27459 );
or \U$19354 ( \27841 , \27830 , \27840 );
and \U$19356 ( \27842 , \27841 , 1'b1 );
or \U$19358 ( \27843 , \27842 , 1'b0 );
buf \U$19359 ( \27844 , \27843 );
_DC r23cc0_GF_IsGateDCbyConstraint ( \27845_nR23cc0 , \27844 , \21944 );
buf \U$19360 ( \27846 , \27845_nR23cc0 );
not \U$19361 ( \27847 , \27558 );
and \U$19362 ( \27848 , RIe198cc8_6106, \27847 );
not \U$19363 ( \27849 , RIe198cc8_6106);
or \U$19364 ( \27850 , \27849 , \27421 );
buf \U$19365 ( \27851 , RIb885bf8_46);
and \U$19366 ( \27852 , \27392 , \27851 );
buf \U$19367 ( \27853 , RIb829678_214);
buf \U$19368 ( \27854 , \27853 );
not \U$19369 ( \27855 , \27400 );
and \U$19370 ( \27856 , \27854 , \27855 );
nor \U$19371 ( \27857 , \27852 , \27856 );
nand \U$19372 ( \27858 , \27850 , \27857 );
and \U$19373 ( \27859 , \27858 , \27558 );
or \U$19374 ( \27860 , \27848 , \27859 );
and \U$19376 ( \27861 , \27860 , 1'b1 );
or \U$19378 ( \27862 , \27861 , 1'b0 );
buf \U$19379 ( \27863 , \27862 );
_DC r23cc2_GF_IsGateDCbyConstraint ( \27864_nR23cc2 , \27863 , \21944 );
buf \U$19380 ( \27865 , \27864_nR23cc2 );
not \U$19381 ( \27866 , \27365 );
and \U$19382 ( \27867 , RIe1a05b8_6107, \27866 );
not \U$19383 ( \27868 , RIe1a05b8_6107);
or \U$19384 ( \27869 , \27868 , \27562 );
buf \U$19385 ( \27870 , RIb885c70_45);
and \U$19386 ( \27871 , \27391 , \27870 );
buf \U$19387 ( \27872 , RIb8296f0_213);
buf \U$19388 ( \27873 , \27872 );
not \U$19389 ( \27874 , \27508 );
and \U$19390 ( \27875 , \27873 , \27874 );
nor \U$19391 ( \27876 , \27871 , \27875 );
nand \U$19392 ( \27877 , \27869 , \27876 );
and \U$19393 ( \27878 , \27877 , \27365 );
or \U$19394 ( \27879 , \27867 , \27878 );
and \U$19396 ( \27880 , \27879 , 1'b1 );
or \U$19398 ( \27881 , \27880 , 1'b0 );
buf \U$19399 ( \27882 , \27881 );
_DC r23cc4_GF_IsGateDCbyConstraint ( \27883_nR23cc4 , \27882 , \21944 );
buf \U$19400 ( \27884 , \27883_nR23cc4 );
not \U$19401 ( \27885 , \27365 );
and \U$19402 ( \27886 , RIe1a6300_6108, \27885 );
not \U$19403 ( \27887 , RIe1a6300_6108);
or \U$19404 ( \27888 , \27887 , \27583 );
buf \U$19405 ( \27889 , \22659 );
and \U$19406 ( \27890 , \27423 , \27889 );
buf \U$19407 ( \27891 , RIb82dae8_212);
buf \U$19408 ( \27892 , \27891 );
not \U$19409 ( \27893 , \27428 );
and \U$19410 ( \27894 , \27892 , \27893 );
nor \U$19411 ( \27895 , \27890 , \27894 );
nand \U$19412 ( \27896 , \27888 , \27895 );
and \U$19413 ( \27897 , \27896 , \27365 );
or \U$19414 ( \27898 , \27886 , \27897 );
and \U$19416 ( \27899 , \27898 , 1'b1 );
or \U$19418 ( \27900 , \27899 , 1'b0 );
buf \U$19419 ( \27901 , \27900 );
_DC r23cc6_GF_IsGateDCbyConstraint ( \27902_nR23cc6 , \27901 , \21944 );
buf \U$19420 ( \27903 , \27902_nR23cc6 );
not \U$19421 ( \27904 , \27558 );
and \U$19422 ( \27905 , RIe1ac318_6109, \27904 );
not \U$19423 ( \27906 , RIe1ac318_6109);
or \U$19424 ( \27907 , \27906 , \27663 );
buf \U$19425 ( \27908 , \22680 );
and \U$19426 ( \27909 , \27391 , \27908 );
buf \U$19427 ( \27910 , RIb82db60_211);
buf \U$19428 ( \27911 , \27910 );
not \U$19429 ( \27912 , \27589 );
and \U$19430 ( \27913 , \27911 , \27912 );
nor \U$19431 ( \27914 , \27909 , \27913 );
nand \U$19432 ( \27915 , \27907 , \27914 );
and \U$19433 ( \27916 , \27915 , \27558 );
or \U$19434 ( \27917 , \27905 , \27916 );
and \U$19436 ( \27918 , \27917 , 1'b1 );
or \U$19438 ( \27919 , \27918 , 1'b0 );
buf \U$19439 ( \27920 , \27919 );
_DC r23cc8_GF_IsGateDCbyConstraint ( \27921_nR23cc8 , \27920 , \21944 );
buf \U$19440 ( \27922 , \27921_nR23cc8 );
not \U$19441 ( \27923 , \27459 );
and \U$19442 ( \27924 , RIe1b2420_6110, \27923 );
not \U$19443 ( \27925 , RIe1b2420_6110);
or \U$19444 ( \27926 , \27925 , \27502 );
buf \U$19445 ( \27927 , \22700 );
and \U$19446 ( \27928 , \27392 , \27927 );
buf \U$19447 ( \27929 , RIb82dbd8_210);
buf \U$19448 ( \27930 , \27929 );
not \U$19449 ( \27931 , \27487 );
and \U$19450 ( \27932 , \27930 , \27931 );
nor \U$19451 ( \27933 , \27928 , \27932 );
nand \U$19452 ( \27934 , \27926 , \27933 );
and \U$19453 ( \27935 , \27934 , \27459 );
or \U$19454 ( \27936 , \27924 , \27935 );
and \U$19456 ( \27937 , \27936 , 1'b1 );
or \U$19458 ( \27938 , \27937 , 1'b0 );
buf \U$19459 ( \27939 , \27938 );
_DC r23cca_GF_IsGateDCbyConstraint ( \27940_nR23cca , \27939 , \21944 );
buf \U$19460 ( \27941 , \27940_nR23cca );
buf \U$19461 ( \27942 , \27458 );
not \U$19462 ( \27943 , \27942 );
and \U$19463 ( \27944 , RIe1b7970_6111, \27943 );
not \U$19464 ( \27945 , RIe1b7970_6111);
or \U$19465 ( \27946 , \27945 , \27663 );
buf \U$19466 ( \27947 , RIb885e50_41);
and \U$19467 ( \27948 , \27423 , \27947 );
buf \U$19468 ( \27949 , \22723 );
not \U$19469 ( \27950 , \27589 );
and \U$19470 ( \27951 , \27949 , \27950 );
nor \U$19471 ( \27952 , \27948 , \27951 );
nand \U$19472 ( \27953 , \27946 , \27952 );
and \U$19473 ( \27954 , \27953 , \27942 );
or \U$19474 ( \27955 , \27944 , \27954 );
and \U$19476 ( \27956 , \27955 , 1'b1 );
or \U$19478 ( \27957 , \27956 , 1'b0 );
buf \U$19479 ( \27958 , \27957 );
_DC r23ccc_GF_IsGateDCbyConstraint ( \27959_nR23ccc , \27958 , \21944 );
buf \U$19480 ( \27960 , \27959_nR23ccc );
not \U$19481 ( \27961 , \27558 );
and \U$19482 ( \27962 , RIe1bce48_6112, \27961 );
not \U$19483 ( \27963 , RIe1bce48_6112);
or \U$19484 ( \27964 , \27963 , \27502 );
buf \U$19485 ( \27965 , RIb885ec8_40);
buf \U$19486 ( \27966 , \27965 );
and \U$19487 ( \27967 , \27423 , \27966 );
buf \U$19488 ( \27968 , \22743 );
not \U$19489 ( \27969 , \27419 );
and \U$19490 ( \27970 , \27968 , \27969 );
nor \U$19491 ( \27971 , \27967 , \27970 );
nand \U$19492 ( \27972 , \27964 , \27971 );
and \U$19493 ( \27973 , \27972 , \27558 );
or \U$19494 ( \27974 , \27962 , \27973 );
and \U$19496 ( \27975 , \27974 , 1'b1 );
or \U$19498 ( \27976 , \27975 , 1'b0 );
buf \U$19499 ( \27977 , \27976 );
_DC r23cce_GF_IsGateDCbyConstraint ( \27978_nR23cce , \27977 , \21944 );
buf \U$19500 ( \27979 , \27978_nR23cce );
buf \U$19501 ( \27980 , \27364 );
not \U$19502 ( \27981 , \27980 );
and \U$19503 ( \27982 , RIe1c12b8_6113, \27981 );
not \U$19504 ( \27983 , RIe1c12b8_6113);
or \U$19505 ( \27984 , \27983 , \27604 );
buf \U$19506 ( \27985 , \22762 );
and \U$19507 ( \27986 , \27391 , \27985 );
buf \U$19508 ( \27987 , RIb82dd40_207);
buf \U$19509 ( \27988 , \27987 );
not \U$19510 ( \27989 , \27487 );
and \U$19511 ( \27990 , \27988 , \27989 );
nor \U$19512 ( \27991 , \27986 , \27990 );
nand \U$19513 ( \27992 , \27984 , \27991 );
and \U$19514 ( \27993 , \27992 , \27980 );
or \U$19515 ( \27994 , \27982 , \27993 );
and \U$19517 ( \27995 , \27994 , 1'b1 );
or \U$19519 ( \27996 , \27995 , 1'b0 );
buf \U$19520 ( \27997 , \27996 );
_DC r23cd2_GF_IsGateDCbyConstraint ( \27998_nR23cd2 , \27997 , \21944 );
buf \U$19521 ( \27999 , \27998_nR23cd2 );
not \U$19522 ( \28000 , \27980 );
and \U$19523 ( \28001 , RIe1c7960_6114, \28000 );
not \U$19524 ( \28002 , RIe1c7960_6114);
or \U$19525 ( \28003 , \28002 , \27389 );
not \U$19526 ( \28004 , \27391 );
not \U$19527 ( \28005 , \28004 );
buf \U$19528 ( \28006 , RIb885fb8_38);
and \U$19529 ( \28007 , \28005 , \28006 );
buf \U$19530 ( \28008 , RIb82ddb8_206);
buf \U$19531 ( \28009 , \28008 );
not \U$19532 ( \28010 , \27589 );
and \U$19533 ( \28011 , \28009 , \28010 );
nor \U$19534 ( \28012 , \28007 , \28011 );
nand \U$19535 ( \28013 , \28003 , \28012 );
and \U$19536 ( \28014 , \28013 , \27980 );
or \U$19537 ( \28015 , \28001 , \28014 );
and \U$19539 ( \28016 , \28015 , 1'b1 );
or \U$19541 ( \28017 , \28016 , 1'b0 );
buf \U$19542 ( \28018 , \28017 );
_DC r23cd4_GF_IsGateDCbyConstraint ( \28019_nR23cd4 , \28018 , \21944 );
buf \U$19543 ( \28020 , \28019_nR23cd4 );
not \U$19544 ( \28021 , \27558 );
and \U$19545 ( \28022 , RIe1cc820_6115, \28021 );
not \U$19546 ( \28023 , RIe1cc820_6115);
or \U$19547 ( \28024 , \28023 , \27604 );
not \U$19548 ( \28025 , \28004 );
buf \U$19549 ( \28026 , \22802 );
and \U$19550 ( \28027 , \28025 , \28026 );
buf \U$19551 ( \28028 , RIb82de30_205);
buf \U$19552 ( \28029 , \28028 );
not \U$19553 ( \28030 , \27400 );
and \U$19554 ( \28031 , \28029 , \28030 );
nor \U$19555 ( \28032 , \28027 , \28031 );
nand \U$19556 ( \28033 , \28024 , \28032 );
and \U$19557 ( \28034 , \28033 , \27558 );
or \U$19558 ( \28035 , \28022 , \28034 );
and \U$19560 ( \28036 , \28035 , 1'b1 );
or \U$19562 ( \28037 , \28036 , 1'b0 );
buf \U$19563 ( \28038 , \28037 );
_DC r23cd6_GF_IsGateDCbyConstraint ( \28039_nR23cd6 , \28038 , \21944 );
buf \U$19564 ( \28040 , \28039_nR23cd6 );
not \U$19565 ( \28041 , \27942 );
and \U$19566 ( \28042 , RIe1d0fd8_6116, \28041 );
not \U$19567 ( \28043 , RIe1d0fd8_6116);
or \U$19568 ( \28044 , \28043 , \27482 );
buf \U$19569 ( \28045 , RIb8860a8_36);
and \U$19570 ( \28046 , \27391 , \28045 );
buf \U$19571 ( \28047 , RIb832228_204);
buf \U$19572 ( \28048 , \28047 );
not \U$19573 ( \28049 , \27487 );
and \U$19574 ( \28050 , \28048 , \28049 );
nor \U$19575 ( \28051 , \28046 , \28050 );
nand \U$19576 ( \28052 , \28044 , \28051 );
and \U$19577 ( \28053 , \28052 , \27942 );
or \U$19578 ( \28054 , \28042 , \28053 );
and \U$19580 ( \28055 , \28054 , 1'b1 );
or \U$19582 ( \28056 , \28055 , 1'b0 );
buf \U$19583 ( \28057 , \28056 );
_DC r23cd8_GF_IsGateDCbyConstraint ( \28058_nR23cd8 , \28057 , \21944 );
buf \U$19584 ( \28059 , \28058_nR23cd8 );
not \U$19585 ( \28060 , \27980 );
and \U$19586 ( \28061 , RIe094940_6117, \28060 );
not \U$19587 ( \28062 , RIe094940_6117);
or \U$19588 ( \28063 , \28062 , \27643 );
buf \U$19589 ( \28064 , \22842 );
and \U$19590 ( \28065 , \27423 , \28064 );
buf \U$19591 ( \28066 , \22845 );
not \U$19592 ( \28067 , \27508 );
and \U$19593 ( \28068 , \28066 , \28067 );
nor \U$19594 ( \28069 , \28065 , \28068 );
nand \U$19595 ( \28070 , \28063 , \28069 );
and \U$19596 ( \28071 , \28070 , \27980 );
or \U$19597 ( \28072 , \28061 , \28071 );
and \U$19599 ( \28073 , \28072 , 1'b1 );
or \U$19601 ( \28074 , \28073 , 1'b0 );
buf \U$19602 ( \28075 , \28074 );
_DC r23cda_GF_IsGateDCbyConstraint ( \28076_nR23cda , \28075 , \21944 );
buf \U$19603 ( \28077 , \28076_nR23cda );
not \U$19604 ( \28078 , \27558 );
and \U$19605 ( \28079 , RIe090368_6118, \28078 );
not \U$19606 ( \28080 , RIe090368_6118);
or \U$19607 ( \28081 , \28080 , \27523 );
buf \U$19608 ( \28082 , RIb886198_34);
and \U$19609 ( \28083 , \27391 , \28082 );
buf \U$19610 ( \28084 , RIb832318_202);
buf \U$19611 ( \28085 , \28084 );
not \U$19612 ( \28086 , \27508 );
and \U$19613 ( \28087 , \28085 , \28086 );
nor \U$19614 ( \28088 , \28083 , \28087 );
nand \U$19615 ( \28089 , \28081 , \28088 );
and \U$19616 ( \28090 , \28089 , \27558 );
or \U$19617 ( \28091 , \28079 , \28090 );
and \U$19619 ( \28092 , \28091 , 1'b1 );
or \U$19621 ( \28093 , \28092 , 1'b0 );
buf \U$19622 ( \28094 , \28093 );
_DC r23cdc_GF_IsGateDCbyConstraint ( \28095_nR23cdc , \28094 , \21944 );
buf \U$19623 ( \28096 , \28095_nR23cdc );
not \U$19624 ( \28097 , \27980 );
and \U$19625 ( \28098 , RIe08b700_6119, \28097 );
not \U$19626 ( \28099 , RIe08b700_6119);
or \U$19627 ( \28100 , \28099 , \27421 );
buf \U$19628 ( \28101 , RIb886210_33);
and \U$19629 ( \28102 , \27391 , \28101 );
buf \U$19630 ( \28103 , RIb832390_201);
buf \U$19631 ( \28104 , \28103 );
not \U$19632 ( \28105 , \27428 );
and \U$19633 ( \28106 , \28104 , \28105 );
nor \U$19634 ( \28107 , \28102 , \28106 );
nand \U$19635 ( \28108 , \28100 , \28107 );
and \U$19636 ( \28109 , \28108 , \27980 );
or \U$19637 ( \28110 , \28098 , \28109 );
and \U$19639 ( \28111 , \28110 , 1'b1 );
or \U$19641 ( \28112 , \28111 , 1'b0 );
buf \U$19642 ( \28113 , \28112 );
_DC r23cde_GF_IsGateDCbyConstraint ( \28114_nR23cde , \28113 , \21944 );
buf \U$19643 ( \28115 , \28114_nR23cde );
not \U$19644 ( \28116 , \27980 );
and \U$19645 ( \28117 , RIe087a10_6120, \28116 );
not \U$19646 ( \28118 , RIe087a10_6120);
or \U$19647 ( \28119 , \28118 , \27482 );
buf \U$19648 ( \28120 , RIb886288_32);
and \U$19649 ( \28121 , \27391 , \28120 );
buf \U$19650 ( \28122 , RIb832408_200);
buf \U$19651 ( \28123 , \28122 );
not \U$19652 ( \28124 , \27400 );
and \U$19653 ( \28125 , \28123 , \28124 );
nor \U$19654 ( \28126 , \28121 , \28125 );
nand \U$19655 ( \28127 , \28119 , \28126 );
and \U$19656 ( \28128 , \28127 , \27980 );
or \U$19657 ( \28129 , \28117 , \28128 );
and \U$19659 ( \28130 , \28129 , 1'b1 );
or \U$19661 ( \28131 , \28130 , 1'b0 );
buf \U$19662 ( \28132 , \28131 );
_DC r23ce0_GF_IsGateDCbyConstraint ( \28133_nR23ce0 , \28132 , \21944 );
buf \U$19663 ( \28134 , \28133_nR23ce0 );
not \U$19664 ( \28135 , \27558 );
and \U$19665 ( \28136 , RIe14c9f0_6121, \28135 );
not \U$19666 ( \28137 , RIe14c9f0_6121);
or \U$19667 ( \28138 , \28137 , \27643 );
buf \U$19668 ( \28139 , RIb886300_31);
and \U$19669 ( \28140 , \27392 , \28139 );
buf \U$19670 ( \28141 , RIb832480_199);
buf \U$19671 ( \28142 , \28141 );
not \U$19672 ( \28143 , \27487 );
and \U$19673 ( \28144 , \28142 , \28143 );
nor \U$19674 ( \28145 , \28140 , \28144 );
nand \U$19675 ( \28146 , \28138 , \28145 );
and \U$19676 ( \28147 , \28146 , \27558 );
or \U$19677 ( \28148 , \28136 , \28147 );
and \U$19679 ( \28149 , \28148 , 1'b1 );
or \U$19681 ( \28150 , \28149 , 1'b0 );
buf \U$19682 ( \28151 , \28150 );
_DC r23ce2_GF_IsGateDCbyConstraint ( \28152_nR23ce2 , \28151 , \21944 );
buf \U$19683 ( \28153 , \28152_nR23ce2 );
not \U$19684 ( \28154 , \27942 );
and \U$19685 ( \28155 , RIe1495e8_6122, \28154 );
not \U$19686 ( \28156 , RIe1495e8_6122);
or \U$19687 ( \28157 , \28156 , \27523 );
buf \U$19688 ( \28158 , RIb886378_30);
and \U$19689 ( \28159 , \27423 , \28158 );
buf \U$19690 ( \28160 , RIb8324f8_198);
buf \U$19691 ( \28161 , \28160 );
not \U$19692 ( \28162 , \27589 );
and \U$19693 ( \28163 , \28161 , \28162 );
nor \U$19694 ( \28164 , \28159 , \28163 );
nand \U$19695 ( \28165 , \28157 , \28164 );
and \U$19696 ( \28166 , \28165 , \27942 );
or \U$19697 ( \28167 , \28155 , \28166 );
and \U$19699 ( \28168 , \28167 , 1'b1 );
or \U$19701 ( \28169 , \28168 , 1'b0 );
buf \U$19702 ( \28170 , \28169 );
_DC r23ce4_GF_IsGateDCbyConstraint ( \28171_nR23ce4 , \28170 , \21944 );
buf \U$19703 ( \28172 , \28171_nR23ce4 );
not \U$19704 ( \28173 , \27942 );
and \U$19705 ( \28174 , RIe146348_6123, \28173 );
not \U$19706 ( \28175 , RIe146348_6123);
or \U$19707 ( \28176 , \28175 , \27562 );
buf \U$19708 ( \28177 , \22964 );
and \U$19709 ( \28178 , \27423 , \28177 );
buf \U$19710 ( \28179 , RIb832570_197);
buf \U$19711 ( \28180 , \28179 );
not \U$19712 ( \28181 , \27589 );
and \U$19713 ( \28182 , \28180 , \28181 );
nor \U$19714 ( \28183 , \28178 , \28182 );
nand \U$19715 ( \28184 , \28176 , \28183 );
and \U$19716 ( \28185 , \28184 , \27942 );
or \U$19717 ( \28186 , \28174 , \28185 );
and \U$19719 ( \28187 , \28186 , 1'b1 );
or \U$19721 ( \28188 , \28187 , 1'b0 );
buf \U$19722 ( \28189 , \28188 );
_DC r23ce8_GF_IsGateDCbyConstraint ( \28190_nR23ce8 , \28189 , \21944 );
buf \U$19723 ( \28191 , \28190_nR23ce8 );
not \U$19724 ( \28192 , \27558 );
and \U$19725 ( \28193 , RIe143210_6124, \28192 );
not \U$19726 ( \28194 , RIe143210_6124);
or \U$19727 ( \28195 , \28194 , \27583 );
buf \U$19728 ( \28196 , RIb886468_28);
and \U$19729 ( \28197 , \27464 , \28196 );
buf \U$19730 ( \28198 , RIb8383a8_196);
buf \U$19731 ( \28199 , \28198 );
not \U$19732 ( \28200 , \27419 );
and \U$19733 ( \28201 , \28199 , \28200 );
nor \U$19734 ( \28202 , \28197 , \28201 );
nand \U$19735 ( \28203 , \28195 , \28202 );
and \U$19736 ( \28204 , \28203 , \27558 );
or \U$19737 ( \28205 , \28193 , \28204 );
and \U$19739 ( \28206 , \28205 , 1'b1 );
or \U$19741 ( \28207 , \28206 , 1'b0 );
buf \U$19742 ( \28208 , \28207 );
_DC r23cea_GF_IsGateDCbyConstraint ( \28209_nR23cea , \28208 , \21944 );
buf \U$19743 ( \28210 , \28209_nR23cea );
not \U$19744 ( \28211 , \27942 );
and \U$19745 ( \28212 , RIe140a38_6125, \28211 );
not \U$19746 ( \28213 , RIe140a38_6125);
or \U$19747 ( \28214 , \28213 , \27663 );
buf \U$19748 ( \28215 , RIb8864e0_27);
and \U$19749 ( \28216 , \27464 , \28215 );
buf \U$19750 ( \28217 , RIb838420_195);
buf \U$19751 ( \28218 , \28217 );
not \U$19752 ( \28219 , \27428 );
and \U$19753 ( \28220 , \28218 , \28219 );
nor \U$19754 ( \28221 , \28216 , \28220 );
nand \U$19755 ( \28222 , \28214 , \28221 );
and \U$19756 ( \28223 , \28222 , \27942 );
or \U$19757 ( \28224 , \28212 , \28223 );
and \U$19759 ( \28225 , \28224 , 1'b1 );
or \U$19761 ( \28226 , \28225 , 1'b0 );
buf \U$19762 ( \28227 , \28226 );
_DC r23cec_GF_IsGateDCbyConstraint ( \28228_nR23cec , \28227 , \21944 );
buf \U$19763 ( \28229 , \28228_nR23cec );
not \U$19764 ( \28230 , \27980 );
and \U$19765 ( \28231 , RIe13d4c8_6126, \28230 );
not \U$19766 ( \28232 , RIe13d4c8_6126);
or \U$19767 ( \28233 , \28232 , \27502 );
not \U$19768 ( \28234 , \27377 );
buf \U$19769 ( \28235 , \23022 );
and \U$19770 ( \28236 , \28234 , \28235 );
buf \U$19771 ( \28237 , \23025 );
not \U$19772 ( \28238 , \27387 );
and \U$19773 ( \28239 , \28237 , \28238 );
nor \U$19774 ( \28240 , \28236 , \28239 );
nand \U$19775 ( \28241 , \28233 , \28240 );
and \U$19776 ( \28242 , \28241 , \27980 );
or \U$19777 ( \28243 , \28231 , \28242 );
and \U$19779 ( \28244 , \28243 , 1'b1 );
or \U$19781 ( \28245 , \28244 , 1'b0 );
buf \U$19782 ( \28246 , \28245 );
_DC r23cee_GF_IsGateDCbyConstraint ( \28247_nR23cee , \28246 , \21944 );
buf \U$19783 ( \28248 , \28247_nR23cee );
buf \U$19784 ( \28249 , \27363 );
not \U$19785 ( \28250 , \28249 );
and \U$19786 ( \28251 , RIe13a660_6127, \28250 );
not \U$19787 ( \28252 , RIe13a660_6127);
or \U$19788 ( \28253 , \28252 , \27389 );
buf \U$19789 ( \28254 , \23044 );
and \U$19790 ( \28255 , \27423 , \28254 );
buf \U$19791 ( \28256 , RIb838510_193);
buf \U$19792 ( \28257 , \28256 );
not \U$19793 ( \28258 , \27487 );
and \U$19794 ( \28259 , \28257 , \28258 );
nor \U$19795 ( \28260 , \28255 , \28259 );
nand \U$19796 ( \28261 , \28253 , \28260 );
and \U$19797 ( \28262 , \28261 , \28249 );
or \U$19798 ( \28263 , \28251 , \28262 );
and \U$19800 ( \28264 , \28263 , 1'b1 );
or \U$19802 ( \28265 , \28264 , 1'b0 );
buf \U$19803 ( \28266 , \28265 );
_DC r23cf0_GF_IsGateDCbyConstraint ( \28267_nR23cf0 , \28266 , \21944 );
buf \U$19804 ( \28268 , \28267_nR23cf0 );
not \U$19805 ( \28269 , \27942 );
and \U$19806 ( \28270 , RIe137168_6128, \28269 );
not \U$19807 ( \28271 , RIe137168_6128);
or \U$19808 ( \28272 , \28271 , \27604 );
buf \U$19809 ( \28273 , \23064 );
and \U$19810 ( \28274 , \27464 , \28273 );
buf \U$19811 ( \28275 , RIb838588_192);
buf \U$19812 ( \28276 , \28275 );
not \U$19813 ( \28277 , \27589 );
and \U$19814 ( \28278 , \28276 , \28277 );
nor \U$19815 ( \28279 , \28274 , \28278 );
nand \U$19816 ( \28280 , \28272 , \28279 );
and \U$19817 ( \28281 , \28280 , \27942 );
or \U$19818 ( \28282 , \28270 , \28281 );
and \U$19820 ( \28283 , \28282 , 1'b1 );
or \U$19822 ( \28284 , \28283 , 1'b0 );
buf \U$19823 ( \28285 , \28284 );
_DC r23cf2_GF_IsGateDCbyConstraint ( \28286_nR23cf2 , \28285 , \21944 );
buf \U$19824 ( \28287 , \28286_nR23cf2 );
not \U$19825 ( \28288 , \27980 );
and \U$19826 ( \28289 , RIe133a18_6129, \28288 );
not \U$19827 ( \28290 , RIe133a18_6129);
or \U$19828 ( \28291 , \28290 , \27562 );
buf \U$19829 ( \28292 , \23084 );
and \U$19830 ( \28293 , \27392 , \28292 );
buf \U$19831 ( \28294 , RIb838600_191);
buf \U$19832 ( \28295 , \28294 );
not \U$19833 ( \28296 , \27508 );
and \U$19834 ( \28297 , \28295 , \28296 );
nor \U$19835 ( \28298 , \28293 , \28297 );
nand \U$19836 ( \28299 , \28291 , \28298 );
and \U$19837 ( \28300 , \28299 , \27980 );
or \U$19838 ( \28301 , \28289 , \28300 );
and \U$19840 ( \28302 , \28301 , 1'b1 );
or \U$19842 ( \28303 , \28302 , 1'b0 );
buf \U$19843 ( \28304 , \28303 );
_DC r23cf4_GF_IsGateDCbyConstraint ( \28305_nR23cf4 , \28304 , \21944 );
buf \U$19844 ( \28306 , \28305_nR23cf4 );
buf \U$19845 ( \28307 , \27363 );
not \U$19846 ( \28308 , \28307 );
and \U$19847 ( \28309 , RIe12fda0_6130, \28308 );
not \U$19848 ( \28310 , RIe12fda0_6130);
or \U$19849 ( \28311 , \28310 , \27583 );
buf \U$19850 ( \28312 , \23104 );
and \U$19851 ( \28313 , \27423 , \28312 );
buf \U$19852 ( \28314 , \23107 );
not \U$19853 ( \28315 , \27428 );
and \U$19854 ( \28316 , \28314 , \28315 );
nor \U$19855 ( \28317 , \28313 , \28316 );
nand \U$19856 ( \28318 , \28311 , \28317 );
and \U$19857 ( \28319 , \28318 , \28307 );
or \U$19858 ( \28320 , \28309 , \28319 );
and \U$19860 ( \28321 , \28320 , 1'b1 );
or \U$19862 ( \28322 , \28321 , 1'b0 );
buf \U$19863 ( \28323 , \28322 );
_DC r23cf6_GF_IsGateDCbyConstraint ( \28324_nR23cf6 , \28323 , \21944 );
buf \U$19864 ( \28325 , \28324_nR23cf6 );
not \U$19865 ( \28326 , \27980 );
and \U$19866 ( \28327 , RIe1280f0_6131, \28326 );
not \U$19867 ( \28328 , RIe1280f0_6131);
or \U$19868 ( \28329 , \28328 , \27663 );
buf \U$19869 ( \28330 , RIb8867b0_21);
and \U$19870 ( \28331 , \27464 , \28330 );
buf \U$19871 ( \28332 , RIb8386f0_189);
buf \U$19872 ( \28333 , \28332 );
not \U$19873 ( \28334 , \27400 );
and \U$19874 ( \28335 , \28333 , \28334 );
nor \U$19875 ( \28336 , \28331 , \28335 );
nand \U$19876 ( \28337 , \28329 , \28336 );
and \U$19877 ( \28338 , \28337 , \27980 );
or \U$19878 ( \28339 , \28327 , \28338 );
and \U$19880 ( \28340 , \28339 , 1'b1 );
or \U$19882 ( \28341 , \28340 , 1'b0 );
buf \U$19883 ( \28342 , \28341 );
_DC r23cf8_GF_IsGateDCbyConstraint ( \28343_nR23cf8 , \28342 , \21944 );
buf \U$19884 ( \28344 , \28343_nR23cf8 );
not \U$19885 ( \28345 , \27980 );
and \U$19886 ( \28346 , RIe121b38_6132, \28345 );
not \U$19887 ( \28347 , RIe121b38_6132);
or \U$19888 ( \28348 , \28347 , \27502 );
buf \U$19889 ( \28349 , \23144 );
and \U$19890 ( \28350 , \27392 , \28349 );
buf \U$19891 ( \28351 , RIb838768_188);
buf \U$19892 ( \28352 , \28351 );
not \U$19893 ( \28353 , \27400 );
and \U$19894 ( \28354 , \28352 , \28353 );
nor \U$19895 ( \28355 , \28350 , \28354 );
nand \U$19896 ( \28356 , \28348 , \28355 );
and \U$19897 ( \28357 , \28356 , \27980 );
or \U$19898 ( \28358 , \28346 , \28357 );
and \U$19900 ( \28359 , \28358 , 1'b1 );
or \U$19902 ( \28360 , \28359 , 1'b0 );
buf \U$19903 ( \28361 , \28360 );
_DC r23cfa_GF_IsGateDCbyConstraint ( \28362_nR23cfa , \28361 , \21944 );
buf \U$19904 ( \28363 , \28362_nR23cfa );
not \U$19905 ( \28364 , \27458 );
and \U$19906 ( \28365 , RIe1194b0_6133, \28364 );
not \U$19907 ( \28366 , RIe1194b0_6133);
or \U$19908 ( \28367 , \28366 , \27643 );
not \U$19909 ( \28368 , \27377 );
buf \U$19910 ( \28369 , \23164 );
and \U$19911 ( \28370 , \28368 , \28369 );
buf \U$19912 ( \28371 , RIb8387e0_187);
buf \U$19913 ( \28372 , \28371 );
not \U$19914 ( \28373 , \27400 );
and \U$19915 ( \28374 , \28372 , \28373 );
nor \U$19916 ( \28375 , \28370 , \28374 );
nand \U$19917 ( \28376 , \28367 , \28375 );
and \U$19918 ( \28377 , \28376 , \27458 );
or \U$19919 ( \28378 , \28365 , \28377 );
and \U$19921 ( \28379 , \28378 , 1'b1 );
or \U$19923 ( \28380 , \28379 , 1'b0 );
buf \U$19924 ( \28381 , \28380 );
_DC r23cfe_GF_IsGateDCbyConstraint ( \28382_nR23cfe , \28381 , \21944 );
buf \U$19925 ( \28383 , \28382_nR23cfe );
not \U$19926 ( \28384 , \27942 );
and \U$19927 ( \28385 , RIe1133a8_6134, \28384 );
not \U$19928 ( \28386 , RIe1133a8_6134);
or \U$19929 ( \28387 , \28386 , \27523 );
not \U$19930 ( \28388 , \27377 );
buf \U$19931 ( \28389 , RIb886918_18);
and \U$19932 ( \28390 , \28388 , \28389 );
buf \U$19933 ( \28391 , RIb838858_186);
buf \U$19934 ( \28392 , \28391 );
not \U$19935 ( \28393 , \27487 );
and \U$19936 ( \28394 , \28392 , \28393 );
nor \U$19937 ( \28395 , \28390 , \28394 );
nand \U$19938 ( \28396 , \28387 , \28395 );
and \U$19939 ( \28397 , \28396 , \27942 );
or \U$19940 ( \28398 , \28385 , \28397 );
and \U$19942 ( \28399 , \28398 , 1'b1 );
or \U$19944 ( \28400 , \28399 , 1'b0 );
buf \U$19945 ( \28401 , \28400 );
_DC r23d00_GF_IsGateDCbyConstraint ( \28402_nR23d00 , \28401 , \21944 );
buf \U$19946 ( \28403 , \28402_nR23d00 );
not \U$19947 ( \28404 , \27942 );
and \U$19948 ( \28405 , RIe10ad20_6135, \28404 );
not \U$19949 ( \28406 , RIe10ad20_6135);
or \U$19950 ( \28407 , \28406 , \27421 );
buf \U$19951 ( \28408 , RIb886990_17);
buf \U$19952 ( \28409 , \28408 );
and \U$19953 ( \28410 , \27392 , \28409 );
buf \U$19954 ( \28411 , RIb8388d0_185);
buf \U$19955 ( \28412 , \28411 );
not \U$19956 ( \28413 , \27589 );
and \U$19957 ( \28414 , \28412 , \28413 );
nor \U$19958 ( \28415 , \28410 , \28414 );
nand \U$19959 ( \28416 , \28407 , \28415 );
and \U$19960 ( \28417 , \28416 , \27942 );
or \U$19961 ( \28418 , \28405 , \28417 );
and \U$19963 ( \28419 , \28418 , 1'b1 );
or \U$19965 ( \28420 , \28419 , 1'b0 );
buf \U$19966 ( \28421 , \28420 );
_DC r23d02_GF_IsGateDCbyConstraint ( \28422_nR23d02 , \28421 , \21944 );
buf \U$19967 ( \28423 , \28422_nR23d02 );
not \U$19968 ( \28424 , \27458 );
and \U$19969 ( \28425 , RIdfd70d0_6136, \28424 );
not \U$19970 ( \28426 , RIdfd70d0_6136);
or \U$19971 ( \28427 , \28426 , \27562 );
not \U$19972 ( \28428 , \27377 );
buf \U$19973 ( \28429 , \23223 );
and \U$19974 ( \28430 , \28428 , \28429 );
buf \U$19975 ( \28431 , RIb838948_184);
buf \U$19976 ( \28432 , \28431 );
not \U$19977 ( \28433 , \27419 );
and \U$19978 ( \28434 , \28432 , \28433 );
nor \U$19979 ( \28435 , \28430 , \28434 );
nand \U$19980 ( \28436 , \28427 , \28435 );
and \U$19981 ( \28437 , \28436 , \27458 );
or \U$19982 ( \28438 , \28425 , \28437 );
and \U$19984 ( \28439 , \28438 , 1'b1 );
or \U$19986 ( \28440 , \28439 , 1'b0 );
buf \U$19987 ( \28441 , \28440 );
_DC r23d04_GF_IsGateDCbyConstraint ( \28442_nR23d04 , \28441 , \21944 );
buf \U$19988 ( \28443 , \28442_nR23d04 );
not \U$19989 ( \28444 , \27980 );
and \U$19990 ( \28445 , RIdff52b0_6137, \28444 );
not \U$19991 ( \28446 , RIdff52b0_6137);
or \U$19992 ( \28447 , \28446 , \27583 );
not \U$19993 ( \28448 , \27377 );
buf \U$19994 ( \28449 , RIb886a80_15);
and \U$19995 ( \28450 , \28448 , \28449 );
buf \U$19996 ( \28451 , RIb8389c0_183);
buf \U$19997 ( \28452 , \28451 );
not \U$19998 ( \28453 , \27400 );
and \U$19999 ( \28454 , \28452 , \28453 );
nor \U$20000 ( \28455 , \28450 , \28454 );
nand \U$20001 ( \28456 , \28447 , \28455 );
and \U$20002 ( \28457 , \28456 , \27980 );
or \U$20003 ( \28458 , \28445 , \28457 );
and \U$20005 ( \28459 , \28458 , 1'b1 );
or \U$20007 ( \28460 , \28459 , 1'b0 );
buf \U$20008 ( \28461 , \28460 );
_DC r23d06_GF_IsGateDCbyConstraint ( \28462_nR23d06 , \28461 , \21944 );
buf \U$20009 ( \28463 , \28462_nR23d06 );
not \U$20010 ( \28464 , \27980 );
and \U$20011 ( \28465 , RIe01ea70_6138, \28464 );
not \U$20012 ( \28466 , RIe01ea70_6138);
or \U$20013 ( \28467 , \28466 , \27389 );
buf \U$20014 ( \28468 , \23263 );
and \U$20015 ( \28469 , \27391 , \28468 );
buf \U$20016 ( \28470 , RIb838a38_182);
buf \U$20017 ( \28471 , \28470 );
not \U$20018 ( \28472 , \27487 );
and \U$20019 ( \28473 , \28471 , \28472 );
nor \U$20020 ( \28474 , \28469 , \28473 );
nand \U$20021 ( \28475 , \28467 , \28474 );
and \U$20022 ( \28476 , \28475 , \27980 );
or \U$20023 ( \28477 , \28465 , \28476 );
and \U$20025 ( \28478 , \28477 , 1'b1 );
or \U$20027 ( \28479 , \28478 , 1'b0 );
buf \U$20028 ( \28480 , \28479 );
_DC r23d08_GF_IsGateDCbyConstraint ( \28481_nR23d08 , \28480 , \21944 );
buf \U$20029 ( \28482 , \28481_nR23d08 );
buf \U$20030 ( \28483 , \27363 );
not \U$20031 ( \28484 , \28483 );
and \U$20032 ( \28485 , RIe03a5e0_6139, \28484 );
not \U$20033 ( \28486 , RIe03a5e0_6139);
or \U$20034 ( \28487 , \28486 , \27604 );
buf \U$20035 ( \28488 , \23283 );
and \U$20036 ( \28489 , \27392 , \28488 );
buf \U$20037 ( \28490 , \23286 );
not \U$20038 ( \28491 , \27589 );
and \U$20039 ( \28492 , \28490 , \28491 );
nor \U$20040 ( \28493 , \28489 , \28492 );
nand \U$20041 ( \28494 , \28487 , \28493 );
and \U$20042 ( \28495 , \28494 , \28483 );
or \U$20043 ( \28496 , \28485 , \28495 );
and \U$20045 ( \28497 , \28496 , 1'b1 );
or \U$20047 ( \28498 , \28497 , 1'b0 );
buf \U$20048 ( \28499 , \28498 );
_DC r23d0a_GF_IsGateDCbyConstraint ( \28500_nR23d0a , \28499 , \21944 );
buf \U$20049 ( \28501 , \28500_nR23d0a );
not \U$20050 ( \28502 , \27942 );
and \U$20051 ( \28503 , RIdfb6cb8_6140, \28502 );
not \U$20052 ( \28504 , RIdfb6cb8_6140);
or \U$20053 ( \28505 , \28504 , \27482 );
buf \U$20054 ( \28506 , RIb886be8_12);
buf \U$20055 ( \28507 , \28506 );
and \U$20056 ( \28508 , \27464 , \28507 );
buf \U$20057 ( \28509 , RIb838b28_180);
buf \U$20058 ( \28510 , \28509 );
not \U$20059 ( \28511 , \27589 );
and \U$20060 ( \28512 , \28510 , \28511 );
nor \U$20061 ( \28513 , \28508 , \28512 );
nand \U$20062 ( \28514 , \28505 , \28513 );
and \U$20063 ( \28515 , \28514 , \27942 );
or \U$20064 ( \28516 , \28503 , \28515 );
and \U$20066 ( \28517 , \28516 , 1'b1 );
or \U$20068 ( \28518 , \28517 , 1'b0 );
buf \U$20069 ( \28519 , \28518 );
_DC r23d0c_GF_IsGateDCbyConstraint ( \28520_nR23d0c , \28519 , \21944 );
buf \U$20070 ( \28521 , \28520_nR23d0c );
not \U$20071 ( \28522 , \27980 );
and \U$20072 ( \28523 , RIdfa46d0_6141, \28522 );
not \U$20073 ( \28524 , RIdfa46d0_6141);
or \U$20074 ( \28525 , \28524 , \27643 );
buf \U$20075 ( \28526 , RIb886c60_11);
and \U$20076 ( \28527 , \27423 , \28526 );
buf \U$20077 ( \28528 , RIb838ba0_179);
buf \U$20078 ( \28529 , \28528 );
not \U$20079 ( \28530 , \27508 );
and \U$20080 ( \28531 , \28529 , \28530 );
nor \U$20081 ( \28532 , \28527 , \28531 );
nand \U$20082 ( \28533 , \28525 , \28532 );
and \U$20083 ( \28534 , \28533 , \27980 );
or \U$20084 ( \28535 , \28523 , \28534 );
and \U$20086 ( \28536 , \28535 , 1'b1 );
or \U$20088 ( \28537 , \28536 , 1'b0 );
buf \U$20089 ( \28538 , \28537 );
_DC r23d0e_GF_IsGateDCbyConstraint ( \28539_nR23d0e , \28538 , \21944 );
buf \U$20090 ( \28540 , \28539_nR23d0e );
buf \U$20091 ( \28541 , \27363 );
not \U$20092 ( \28542 , \28541 );
and \U$20093 ( \28543 , RIdf7c7e8_6142, \28542 );
not \U$20094 ( \28544 , RIdf7c7e8_6142);
or \U$20095 ( \28545 , \28544 , \27663 );
not \U$20096 ( \28546 , \27377 );
buf \U$20097 ( \28547 , RIb886cd8_10);
buf \U$20098 ( \28548 , \28547 );
and \U$20099 ( \28549 , \28546 , \28548 );
buf \U$20100 ( \28550 , RIb838c18_178);
buf \U$20101 ( \28551 , \28550 );
not \U$20102 ( \28552 , \27487 );
and \U$20103 ( \28553 , \28551 , \28552 );
nor \U$20104 ( \28554 , \28549 , \28553 );
nand \U$20105 ( \28555 , \28545 , \28554 );
and \U$20106 ( \28556 , \28555 , \28541 );
or \U$20107 ( \28557 , \28543 , \28556 );
and \U$20109 ( \28558 , \28557 , 1'b1 );
or \U$20111 ( \28559 , \28558 , 1'b0 );
buf \U$20112 ( \28560 , \28559 );
_DC r23d10_GF_IsGateDCbyConstraint ( \28561_nR23d10 , \28560 , \21944 );
buf \U$20113 ( \28562 , \28561_nR23d10 );
buf \U$20114 ( \28563 , \28541 );
not \U$20115 ( \28564 , \28563 );
and \U$20116 ( \28565 , RIdc22218_6143, \28564 );
not \U$20117 ( \28566 , RIdc22218_6143);
or \U$20118 ( \28567 , \28566 , \27389 );
buf \U$20119 ( \28568 , RIb886d50_9);
buf \U$20120 ( \28569 , \28568 );
and \U$20121 ( \28570 , \27464 , \28569 );
buf \U$20122 ( \28571 , RIb838c90_177);
not \U$20123 ( \28572 , \27428 );
and \U$20124 ( \28573 , \28571 , \28572 );
nor \U$20125 ( \28574 , \28570 , \28573 );
nand \U$20126 ( \28575 , \28567 , \28574 );
and \U$20127 ( \28576 , \28575 , \28563 );
or \U$20128 ( \28577 , \28565 , \28576 );
and \U$20130 ( \28578 , \28577 , 1'b1 );
or \U$20132 ( \28579 , \28578 , 1'b0 );
buf \U$20133 ( \28580 , \28579 );
_DC r23d14_GF_IsGateDCbyConstraint ( \28581_nR23d14 , \28580 , \21944 );
buf \U$20134 ( \28582 , \28581_nR23d14 );
not \U$20135 ( \28583 , \28563 );
and \U$20136 ( \28584 , RIda953d8_6144, \28583 );
not \U$20137 ( \28585 , RIda953d8_6144);
or \U$20138 ( \28586 , \28585 , \27604 );
buf \U$20139 ( \28587 , RIb886dc8_8);
and \U$20140 ( \28588 , \27392 , \28587 );
buf \U$20141 ( \28589 , \23386 );
not \U$20142 ( \28590 , \27400 );
and \U$20143 ( \28591 , \28589 , \28590 );
nor \U$20144 ( \28592 , \28588 , \28591 );
nand \U$20145 ( \28593 , \28586 , \28592 );
and \U$20146 ( \28594 , \28593 , \28563 );
or \U$20147 ( \28595 , \28584 , \28594 );
and \U$20149 ( \28596 , \28595 , 1'b1 );
or \U$20151 ( \28597 , \28596 , 1'b0 );
buf \U$20152 ( \28598 , \28597 );
_DC r23d16_GF_IsGateDCbyConstraint ( \28599_nR23d16 , \28598 , \21944 );
buf \U$20153 ( \28600 , \28599_nR23d16 );
not \U$20154 ( \28601 , \28541 );
and \U$20155 ( \28602 , RIddeaf80_6145, \28601 );
not \U$20156 ( \28603 , RIddeaf80_6145);
or \U$20157 ( \28604 , \28603 , \27482 );
buf \U$20158 ( \28605 , RIb886e40_7);
buf \U$20159 ( \28606 , \28605 );
and \U$20160 ( \28607 , \27464 , \28606 );
buf \U$20161 ( \28608 , \23406 );
not \U$20162 ( \28609 , \27487 );
and \U$20163 ( \28610 , \28608 , \28609 );
nor \U$20164 ( \28611 , \28607 , \28610 );
nand \U$20165 ( \28612 , \28604 , \28611 );
and \U$20166 ( \28613 , \28612 , \28541 );
or \U$20167 ( \28614 , \28602 , \28613 );
and \U$20169 ( \28615 , \28614 , 1'b1 );
or \U$20171 ( \28616 , \28615 , 1'b0 );
buf \U$20172 ( \28617 , \28616 );
_DC r23d18_GF_IsGateDCbyConstraint ( \28618_nR23d18 , \28617 , \21944 );
buf \U$20173 ( \28619 , \28618_nR23d18 );
not \U$20174 ( \28620 , \27942 );
and \U$20175 ( \28621 , RIde58a80_6146, \28620 );
not \U$20176 ( \28622 , RIde58a80_6146);
or \U$20177 ( \28623 , \28622 , \27643 );
buf \U$20178 ( \28624 , \23423 );
and \U$20179 ( \28625 , \27392 , \28624 );
buf \U$20180 ( \28626 , RIb838df8_174);
not \U$20181 ( \28627 , \27589 );
and \U$20182 ( \28628 , \28626 , \28627 );
nor \U$20183 ( \28629 , \28625 , \28628 );
nand \U$20184 ( \28630 , \28623 , \28629 );
and \U$20185 ( \28631 , \28630 , \27942 );
or \U$20186 ( \28632 , \28621 , \28631 );
and \U$20188 ( \28633 , \28632 , 1'b1 );
or \U$20190 ( \28634 , \28633 , 1'b0 );
buf \U$20191 ( \28635 , \28634 );
_DC r23d1a_GF_IsGateDCbyConstraint ( \28636_nR23d1a , \28635 , \21944 );
buf \U$20192 ( \28637 , \28636_nR23d1a );
not \U$20193 ( \28638 , \27942 );
and \U$20194 ( \28639 , RIe03fa40_6147, \28638 );
not \U$20195 ( \28640 , RIe03fa40_6147);
not \U$20196 ( \28641 , \27383 );
nor \U$20197 ( \28642 , \27380 , \28641 );
and \U$20198 ( \28643 , \28642 , \27385 );
not \U$20199 ( \28644 , \27370 );
or \U$20200 ( \28645 , \27372 , \28644 );
not \U$20201 ( \28646 , \28645 );
nand \U$20202 ( \28647 , \27362 , \28646 );
not \U$20203 ( \28648 , \28647 );
or \U$20204 ( \28649 , \28643 , \28648 );
not \U$20205 ( \28650 , \28649 );
not \U$20206 ( \28651 , \28650 );
or \U$20207 ( \28652 , \28640 , \28651 );
not \U$20208 ( \28653 , \28643 );
not \U$20209 ( \28654 , \28653 );
and \U$20210 ( \28655 , \27395 , \28654 );
not \U$20211 ( \28656 , \28655 );
not \U$20212 ( \28657 , \27393 );
not \U$20213 ( \28658 , \28647 );
buf \U$20214 ( \28659 , \28658 );
not \U$20215 ( \28660 , \28659 );
or \U$20216 ( \28661 , \28657 , \28660 );
nand \U$20217 ( \28662 , \28652 , \28656 , \28661 );
and \U$20218 ( \28663 , \28662 , \27942 );
or \U$20219 ( \28664 , \28639 , \28663 );
and \U$20221 ( \28665 , \28664 , 1'b1 );
or \U$20223 ( \28666 , \28665 , 1'b0 );
buf \U$20224 ( \28667 , \28666 );
_DC r23d24_GF_IsGateDCbyConstraint ( \28668_nR23d24 , \28667 , \21944 );
buf \U$20225 ( \28669 , \28668_nR23d24 );
not \U$20226 ( \28670 , \28541 );
and \U$20227 ( \28671 , RIe04e338_6148, \28670 );
not \U$20228 ( \28672 , RIe04e338_6148);
not \U$20229 ( \28673 , \28650 );
or \U$20230 ( \28674 , \28672 , \28673 );
not \U$20231 ( \28675 , \28643 );
not \U$20232 ( \28676 , \28675 );
and \U$20233 ( \28677 , \27427 , \28676 );
not \U$20234 ( \28678 , \28677 );
not \U$20235 ( \28679 , \27424 );
buf \U$20236 ( \28680 , \28658 );
not \U$20237 ( \28681 , \28680 );
or \U$20238 ( \28682 , \28679 , \28681 );
nand \U$20239 ( \28683 , \28674 , \28678 , \28682 );
and \U$20240 ( \28684 , \28683 , \28541 );
or \U$20241 ( \28685 , \28671 , \28684 );
and \U$20243 ( \28686 , \28685 , 1'b1 );
or \U$20245 ( \28687 , \28686 , 1'b0 );
buf \U$20246 ( \28688 , \28687 );
_DC r23d3a_GF_IsGateDCbyConstraint ( \28689_nR23d3a , \28688 , \21944 );
buf \U$20247 ( \28690 , \28689_nR23d3a );
not \U$20248 ( \28691 , \27942 );
and \U$20249 ( \28692 , RIe0629f0_6149, \28691 );
not \U$20250 ( \28693 , RIe0629f0_6149);
not \U$20251 ( \28694 , \28650 );
or \U$20252 ( \28695 , \28693 , \28694 );
not \U$20253 ( \28696 , \28675 );
and \U$20254 ( \28697 , \27446 , \28696 );
not \U$20255 ( \28698 , \28697 );
not \U$20256 ( \28699 , \27444 );
not \U$20257 ( \28700 , \28659 );
or \U$20258 ( \28701 , \28699 , \28700 );
nand \U$20259 ( \28702 , \28695 , \28698 , \28701 );
and \U$20260 ( \28703 , \28702 , \27942 );
or \U$20261 ( \28704 , \28692 , \28703 );
and \U$20263 ( \28705 , \28704 , 1'b1 );
or \U$20265 ( \28706 , \28705 , 1'b0 );
buf \U$20266 ( \28707 , \28706 );
_DC r23d50_GF_IsGateDCbyConstraint ( \28708_nR23d50 , \28707 , \21944 );
buf \U$20267 ( \28709 , \28708_nR23d50 );
not \U$20268 ( \28710 , \28563 );
and \U$20269 ( \28711 , RIe06c608_6150, \28710 );
not \U$20270 ( \28712 , RIe06c608_6150);
not \U$20271 ( \28713 , \28650 );
or \U$20272 ( \28714 , \28712 , \28713 );
not \U$20273 ( \28715 , \28643 );
not \U$20274 ( \28716 , \28715 );
and \U$20275 ( \28717 , \27467 , \28716 );
not \U$20276 ( \28718 , \28717 );
not \U$20277 ( \28719 , \27465 );
not \U$20278 ( \28720 , \28659 );
or \U$20279 ( \28721 , \28719 , \28720 );
nand \U$20280 ( \28722 , \28714 , \28718 , \28721 );
and \U$20281 ( \28723 , \28722 , \28563 );
or \U$20282 ( \28724 , \28711 , \28723 );
and \U$20284 ( \28725 , \28724 , 1'b1 );
or \U$20286 ( \28726 , \28725 , 1'b0 );
buf \U$20287 ( \28727 , \28726 );
_DC r23d66_GF_IsGateDCbyConstraint ( \28728_nR23d66 , \28727 , \21944 );
buf \U$20288 ( \28729 , \28728_nR23d66 );
not \U$20289 ( \28730 , \28249 );
and \U$20290 ( \28731 , RIe0732e0_6151, \28730 );
not \U$20291 ( \28732 , RIe0732e0_6151);
or \U$20292 ( \28733 , \28732 , \28713 );
not \U$20293 ( \28734 , \28653 );
and \U$20294 ( \28735 , \27486 , \28734 );
not \U$20295 ( \28736 , \28735 );
not \U$20296 ( \28737 , \27484 );
buf \U$20297 ( \28738 , \28658 );
not \U$20298 ( \28739 , \28738 );
or \U$20299 ( \28740 , \28737 , \28739 );
nand \U$20300 ( \28741 , \28733 , \28736 , \28740 );
and \U$20301 ( \28742 , \28741 , \28249 );
or \U$20302 ( \28743 , \28731 , \28742 );
and \U$20304 ( \28744 , \28743 , 1'b1 );
or \U$20306 ( \28745 , \28744 , 1'b0 );
buf \U$20307 ( \28746 , \28745 );
_DC r23d7c_GF_IsGateDCbyConstraint ( \28747_nR23d7c , \28746 , \21944 );
buf \U$20308 ( \28748 , \28747_nR23d7c );
buf \U$20309 ( \28749 , \28307 );
not \U$20310 ( \28750 , \28749 );
and \U$20311 ( \28751 , RIe07d0d8_6152, \28750 );
not \U$20312 ( \28752 , RIe07d0d8_6152);
or \U$20313 ( \28753 , \28752 , \28713 );
not \U$20314 ( \28754 , \28643 );
not \U$20315 ( \28755 , \28754 );
and \U$20316 ( \28756 , \27507 , \28755 );
not \U$20317 ( \28757 , \28756 );
not \U$20318 ( \28758 , \27504 );
not \U$20319 ( \28759 , \28738 );
or \U$20320 ( \28760 , \28758 , \28759 );
nand \U$20321 ( \28761 , \28753 , \28757 , \28760 );
and \U$20322 ( \28762 , \28761 , \28749 );
or \U$20323 ( \28763 , \28751 , \28762 );
and \U$20325 ( \28764 , \28763 , 1'b1 );
or \U$20327 ( \28765 , \28764 , 1'b0 );
buf \U$20328 ( \28766 , \28765 );
_DC r23d92_GF_IsGateDCbyConstraint ( \28767_nR23d92 , \28766 , \21944 );
buf \U$20329 ( \28768 , \28767_nR23d92 );
not \U$20330 ( \28769 , \28749 );
and \U$20331 ( \28770 , RIe084158_6153, \28769 );
not \U$20332 ( \28771 , RIe084158_6153);
or \U$20333 ( \28772 , \28771 , \28673 );
not \U$20334 ( \28773 , \28643 );
not \U$20335 ( \28774 , \28773 );
and \U$20336 ( \28775 , \27527 , \28774 );
not \U$20337 ( \28776 , \28775 );
not \U$20338 ( \28777 , \27525 );
not \U$20339 ( \28778 , \28680 );
or \U$20340 ( \28779 , \28777 , \28778 );
nand \U$20341 ( \28780 , \28772 , \28776 , \28779 );
and \U$20342 ( \28781 , \28780 , \28749 );
or \U$20343 ( \28782 , \28770 , \28781 );
and \U$20345 ( \28783 , \28782 , 1'b1 );
or \U$20347 ( \28784 , \28783 , 1'b0 );
buf \U$20348 ( \28785 , \28784 );
_DC r23d9c_GF_IsGateDCbyConstraint ( \28786_nR23d9c , \28785 , \21944 );
buf \U$20349 ( \28787 , \28786_nR23d9c );
not \U$20350 ( \28788 , \28483 );
and \U$20351 ( \28789 , RIdfc61e0_6154, \28788 );
not \U$20352 ( \28790 , RIdfc61e0_6154);
or \U$20353 ( \28791 , \28790 , \28713 );
not \U$20354 ( \28792 , \28715 );
and \U$20355 ( \28793 , \27546 , \28792 );
not \U$20356 ( \28794 , \28793 );
not \U$20357 ( \28795 , \27543 );
not \U$20358 ( \28796 , \28738 );
or \U$20359 ( \28797 , \28795 , \28796 );
nand \U$20360 ( \28798 , \28791 , \28794 , \28797 );
and \U$20361 ( \28799 , \28798 , \28483 );
or \U$20362 ( \28800 , \28789 , \28799 );
and \U$20364 ( \28801 , \28800 , 1'b1 );
or \U$20366 ( \28802 , \28801 , 1'b0 );
buf \U$20367 ( \28803 , \28802 );
_DC r23d9e_GF_IsGateDCbyConstraint ( \28804_nR23d9e , \28803 , \21944 );
buf \U$20368 ( \28805 , \28804_nR23d9e );
not \U$20369 ( \28806 , \28563 );
and \U$20370 ( \28807 , RIe106838_6155, \28806 );
not \U$20371 ( \28808 , RIe106838_6155);
or \U$20372 ( \28809 , \28808 , \28651 );
not \U$20373 ( \28810 , \28754 );
and \U$20374 ( \28811 , \27568 , \28810 );
not \U$20375 ( \28812 , \28811 );
not \U$20376 ( \28813 , \27565 );
not \U$20377 ( \28814 , \28738 );
or \U$20378 ( \28815 , \28813 , \28814 );
nand \U$20379 ( \28816 , \28809 , \28812 , \28815 );
and \U$20380 ( \28817 , \28816 , \28563 );
or \U$20381 ( \28818 , \28807 , \28817 );
and \U$20383 ( \28819 , \28818 , 1'b1 );
or \U$20385 ( \28820 , \28819 , 1'b0 );
buf \U$20386 ( \28821 , \28820 );
_DC r23da0_GF_IsGateDCbyConstraint ( \28822_nR23da0 , \28821 , \21944 );
buf \U$20387 ( \28823 , \28822_nR23da0 );
not \U$20388 ( \28824 , \28563 );
and \U$20389 ( \28825 , RIe0f8198_6156, \28824 );
not \U$20390 ( \28826 , RIe0f8198_6156);
or \U$20391 ( \28827 , \28826 , \28651 );
not \U$20392 ( \28828 , \28675 );
and \U$20393 ( \28829 , \27588 , \28828 );
not \U$20394 ( \28830 , \28829 );
nand \U$20395 ( \28831 , \27585 , \28680 );
nand \U$20396 ( \28832 , \28827 , \28830 , \28831 );
and \U$20397 ( \28833 , \28832 , \28563 );
or \U$20398 ( \28834 , \28825 , \28833 );
and \U$20400 ( \28835 , \28834 , 1'b1 );
or \U$20402 ( \28836 , \28835 , 1'b0 );
buf \U$20403 ( \28837 , \28836 );
_DC r23da2_GF_IsGateDCbyConstraint ( \28838_nR23da2 , \28837 , \21944 );
buf \U$20404 ( \28839 , \28838_nR23da2 );
not \U$20405 ( \28840 , \28307 );
and \U$20406 ( \28841 , RIe0eed00_6157, \28840 );
not \U$20407 ( \28842 , RIe0eed00_6157);
not \U$20408 ( \28843 , \28650 );
or \U$20409 ( \28844 , \28842 , \28843 );
not \U$20410 ( \28845 , \28754 );
and \U$20411 ( \28846 , \27609 , \28845 );
not \U$20412 ( \28847 , \28846 );
nand \U$20413 ( \28848 , \27606 , \28738 );
nand \U$20414 ( \28849 , \28844 , \28847 , \28848 );
and \U$20415 ( \28850 , \28849 , \28307 );
or \U$20416 ( \28851 , \28841 , \28850 );
and \U$20418 ( \28852 , \28851 , 1'b1 );
or \U$20420 ( \28853 , \28852 , 1'b0 );
buf \U$20421 ( \28854 , \28853 );
_DC r23d26_GF_IsGateDCbyConstraint ( \28855_nR23d26 , \28854 , \21944 );
buf \U$20422 ( \28856 , \28855_nR23d26 );
not \U$20423 ( \28857 , \28749 );
and \U$20424 ( \28858 , RIe0e2b68_6158, \28857 );
not \U$20425 ( \28859 , RIe0e2b68_6158);
or \U$20426 ( \28860 , \28859 , \28673 );
not \U$20427 ( \28861 , \28653 );
and \U$20428 ( \28862 , \27628 , \28861 );
not \U$20429 ( \28863 , \28862 );
nand \U$20430 ( \28864 , \27625 , \28659 );
nand \U$20431 ( \28865 , \28860 , \28863 , \28864 );
and \U$20432 ( \28866 , \28865 , \28749 );
or \U$20433 ( \28867 , \28858 , \28866 );
and \U$20435 ( \28868 , \28867 , 1'b1 );
or \U$20437 ( \28869 , \28868 , 1'b0 );
buf \U$20438 ( \28870 , \28869 );
_DC r23d28_GF_IsGateDCbyConstraint ( \28871_nR23d28 , \28870 , \21944 );
buf \U$20439 ( \28872 , \28871_nR23d28 );
not \U$20440 ( \28873 , \28749 );
and \U$20441 ( \28874 , RIe0d0b98_6159, \28873 );
not \U$20442 ( \28875 , RIe0d0b98_6159);
or \U$20443 ( \28876 , \28875 , \28673 );
not \U$20444 ( \28877 , \28773 );
and \U$20445 ( \28878 , \27648 , \28877 );
not \U$20446 ( \28879 , \28878 );
nand \U$20447 ( \28880 , \27645 , \28738 );
nand \U$20448 ( \28881 , \28876 , \28879 , \28880 );
and \U$20449 ( \28882 , \28881 , \28749 );
or \U$20450 ( \28883 , \28874 , \28882 );
and \U$20452 ( \28884 , \28883 , 1'b1 );
or \U$20454 ( \28885 , \28884 , 1'b0 );
buf \U$20455 ( \28886 , \28885 );
_DC r23d2a_GF_IsGateDCbyConstraint ( \28887_nR23d2a , \28886 , \21944 );
buf \U$20456 ( \28888 , \28887_nR23d2a );
buf \U$20457 ( \28889 , \27363 );
not \U$20458 ( \28890 , \28889 );
and \U$20459 ( \28891 , RIe0c3998_6160, \28890 );
not \U$20460 ( \28892 , RIe0c3998_6160);
or \U$20461 ( \28893 , \28892 , \28673 );
not \U$20462 ( \28894 , \28773 );
and \U$20463 ( \28895 , \27668 , \28894 );
not \U$20464 ( \28896 , \28895 );
nand \U$20465 ( \28897 , \27665 , \28659 );
nand \U$20466 ( \28898 , \28893 , \28896 , \28897 );
and \U$20467 ( \28899 , \28898 , \28889 );
or \U$20468 ( \28900 , \28891 , \28899 );
and \U$20470 ( \28901 , \28900 , 1'b1 );
or \U$20472 ( \28902 , \28901 , 1'b0 );
buf \U$20473 ( \28903 , \28902 );
_DC r23d2c_GF_IsGateDCbyConstraint ( \28904_nR23d2c , \28903 , \21944 );
buf \U$20474 ( \28905 , \28904_nR23d2c );
not \U$20475 ( \28906 , \28749 );
and \U$20476 ( \28907 , RIe0b0960_6161, \28906 );
not \U$20477 ( \28908 , RIe0b0960_6161);
or \U$20478 ( \28909 , \28908 , \28651 );
not \U$20479 ( \28910 , \28754 );
and \U$20480 ( \28911 , \27686 , \28910 );
not \U$20481 ( \28912 , \28911 );
nand \U$20482 ( \28913 , \27684 , \28680 );
nand \U$20483 ( \28914 , \28909 , \28912 , \28913 );
and \U$20484 ( \28915 , \28914 , \28749 );
or \U$20485 ( \28916 , \28907 , \28915 );
and \U$20487 ( \28917 , \28916 , 1'b1 );
or \U$20489 ( \28918 , \28917 , 1'b0 );
buf \U$20490 ( \28919 , \28918 );
_DC r23d2e_GF_IsGateDCbyConstraint ( \28920_nR23d2e , \28919 , \21944 );
buf \U$20491 ( \28921 , \28920_nR23d2e );
not \U$20492 ( \28922 , \28563 );
and \U$20493 ( \28923 , RIe0a6988_6162, \28922 );
not \U$20494 ( \28924 , RIe0a6988_6162);
or \U$20495 ( \28925 , \28924 , \28651 );
not \U$20496 ( \28926 , \28653 );
and \U$20497 ( \28927 , \27704 , \28926 );
not \U$20498 ( \28928 , \28927 );
buf \U$20499 ( \28929 , \28658 );
nand \U$20500 ( \28930 , \27702 , \28929 );
nand \U$20501 ( \28931 , \28925 , \28928 , \28930 );
and \U$20502 ( \28932 , \28931 , \28563 );
or \U$20503 ( \28933 , \28923 , \28932 );
and \U$20505 ( \28934 , \28933 , 1'b1 );
or \U$20507 ( \28935 , \28934 , 1'b0 );
buf \U$20508 ( \28936 , \28935 );
_DC r23d30_GF_IsGateDCbyConstraint ( \28937_nR23d30 , \28936 , \21944 );
buf \U$20509 ( \28938 , \28937_nR23d30 );
buf \U$20510 ( \28939 , \28541 );
not \U$20511 ( \28940 , \28939 );
and \U$20512 ( \28941 , RIe099440_6163, \28940 );
not \U$20513 ( \28942 , RIe099440_6163);
or \U$20514 ( \28943 , \28942 , \28843 );
not \U$20515 ( \28944 , \28653 );
and \U$20516 ( \28945 , \27722 , \28944 );
not \U$20517 ( \28946 , \28945 );
nand \U$20518 ( \28947 , \27720 , \28929 );
nand \U$20519 ( \28948 , \28943 , \28946 , \28947 );
and \U$20520 ( \28949 , \28948 , \28939 );
or \U$20521 ( \28950 , \28941 , \28949 );
and \U$20523 ( \28951 , \28950 , 1'b1 );
or \U$20525 ( \28952 , \28951 , 1'b0 );
buf \U$20526 ( \28953 , \28952 );
_DC r23d32_GF_IsGateDCbyConstraint ( \28954_nR23d32 , \28953 , \21944 );
buf \U$20527 ( \28955 , \28954_nR23d32 );
not \U$20528 ( \28956 , \28749 );
and \U$20529 ( \28957 , RIe1d3c60_6164, \28956 );
not \U$20530 ( \28958 , RIe1d3c60_6164);
or \U$20531 ( \28959 , \28958 , \28673 );
not \U$20532 ( \28960 , \28773 );
and \U$20533 ( \28961 , \27741 , \28960 );
not \U$20534 ( \28962 , \28961 );
nand \U$20535 ( \28963 , \27738 , \28659 );
nand \U$20536 ( \28964 , \28959 , \28962 , \28963 );
and \U$20537 ( \28965 , \28964 , \28749 );
or \U$20538 ( \28966 , \28957 , \28965 );
and \U$20540 ( \28967 , \28966 , 1'b1 );
or \U$20542 ( \28968 , \28967 , 1'b0 );
buf \U$20543 ( \28969 , \28968 );
_DC r23d34_GF_IsGateDCbyConstraint ( \28970_nR23d34 , \28969 , \21944 );
buf \U$20544 ( \28971 , \28970_nR23d34 );
not \U$20545 ( \28972 , \28563 );
and \U$20546 ( \28973 , RIe1d69d8_6165, \28972 );
not \U$20547 ( \28974 , RIe1d69d8_6165);
or \U$20548 ( \28975 , \28974 , \28694 );
not \U$20549 ( \28976 , \28715 );
and \U$20550 ( \28977 , \27760 , \28976 );
not \U$20551 ( \28978 , \28977 );
nand \U$20552 ( \28979 , \27757 , \28929 );
nand \U$20553 ( \28980 , \28975 , \28978 , \28979 );
and \U$20554 ( \28981 , \28980 , \28563 );
or \U$20555 ( \28982 , \28973 , \28981 );
and \U$20557 ( \28983 , \28982 , 1'b1 );
or \U$20559 ( \28984 , \28983 , 1'b0 );
buf \U$20560 ( \28985 , \28984 );
_DC r23d36_GF_IsGateDCbyConstraint ( \28986_nR23d36 , \28985 , \21944 );
buf \U$20561 ( \28987 , \28986_nR23d36 );
not \U$20562 ( \28988 , \28939 );
and \U$20563 ( \28989 , RIe1d9c00_6166, \28988 );
not \U$20564 ( \28990 , RIe1d9c00_6166);
or \U$20565 ( \28991 , \28990 , \28713 );
not \U$20566 ( \28992 , \28773 );
and \U$20567 ( \28993 , \27779 , \28992 );
not \U$20568 ( \28994 , \28993 );
not \U$20569 ( \28995 , \27776 );
not \U$20570 ( \28996 , \28929 );
or \U$20571 ( \28997 , \28995 , \28996 );
nand \U$20572 ( \28998 , \28991 , \28994 , \28997 );
and \U$20573 ( \28999 , \28998 , \28939 );
or \U$20574 ( \29000 , \28989 , \28999 );
and \U$20576 ( \29001 , \29000 , 1'b1 );
or \U$20578 ( \29002 , \29001 , 1'b0 );
buf \U$20579 ( \29003 , \29002 );
_DC r23d38_GF_IsGateDCbyConstraint ( \29004_nR23d38 , \29003 , \21944 );
buf \U$20580 ( \29005 , \29004_nR23d38 );
not \U$20581 ( \29006 , \28563 );
and \U$20582 ( \29007 , RIe1dc978_6167, \29006 );
not \U$20583 ( \29008 , RIe1dc978_6167);
or \U$20584 ( \29009 , \29008 , \28651 );
not \U$20585 ( \29010 , \28754 );
and \U$20586 ( \29011 , \27799 , \29010 );
not \U$20587 ( \29012 , \29011 );
not \U$20588 ( \29013 , \27796 );
not \U$20589 ( \29014 , \28659 );
or \U$20590 ( \29015 , \29013 , \29014 );
nand \U$20591 ( \29016 , \29009 , \29012 , \29015 );
and \U$20592 ( \29017 , \29016 , \28563 );
or \U$20593 ( \29018 , \29007 , \29017 );
and \U$20595 ( \29019 , \29018 , 1'b1 );
or \U$20597 ( \29020 , \29019 , 1'b0 );
buf \U$20598 ( \29021 , \29020 );
_DC r23d3c_GF_IsGateDCbyConstraint ( \29022_nR23d3c , \29021 , \21944 );
buf \U$20599 ( \29023 , \29022_nR23d3c );
not \U$20600 ( \29024 , \28563 );
and \U$20601 ( \29025 , RIe1dfba0_6168, \29024 );
not \U$20602 ( \29026 , RIe1dfba0_6168);
or \U$20603 ( \29027 , \29026 , \28694 );
not \U$20604 ( \29028 , \28675 );
and \U$20605 ( \29029 , \27817 , \29028 );
not \U$20606 ( \29030 , \29029 );
not \U$20607 ( \29031 , \27815 );
not \U$20608 ( \29032 , \28659 );
or \U$20609 ( \29033 , \29031 , \29032 );
nand \U$20610 ( \29034 , \29027 , \29030 , \29033 );
and \U$20611 ( \29035 , \29034 , \28563 );
or \U$20612 ( \29036 , \29025 , \29035 );
and \U$20614 ( \29037 , \29036 , 1'b1 );
or \U$20616 ( \29038 , \29037 , 1'b0 );
buf \U$20617 ( \29039 , \29038 );
_DC r23d3e_GF_IsGateDCbyConstraint ( \29040_nR23d3e , \29039 , \21944 );
buf \U$20618 ( \29041 , \29040_nR23d3e );
not \U$20619 ( \29042 , \28939 );
and \U$20620 ( \29043 , RIe1e2918_6169, \29042 );
not \U$20621 ( \29044 , RIe1e2918_6169);
or \U$20622 ( \29045 , \29044 , \28843 );
not \U$20623 ( \29046 , \28715 );
and \U$20624 ( \29047 , \27835 , \29046 );
not \U$20625 ( \29048 , \29047 );
not \U$20626 ( \29049 , \27833 );
not \U$20627 ( \29050 , \28659 );
or \U$20628 ( \29051 , \29049 , \29050 );
nand \U$20629 ( \29052 , \29045 , \29048 , \29051 );
and \U$20630 ( \29053 , \29052 , \28939 );
or \U$20631 ( \29054 , \29043 , \29053 );
and \U$20633 ( \29055 , \29054 , 1'b1 );
or \U$20635 ( \29056 , \29055 , 1'b0 );
buf \U$20636 ( \29057 , \29056 );
_DC r23d40_GF_IsGateDCbyConstraint ( \29058_nR23d40 , \29057 , \21944 );
buf \U$20637 ( \29059 , \29058_nR23d40 );
not \U$20638 ( \29060 , \28749 );
and \U$20639 ( \29061 , RIe1e5b40_6170, \29060 );
not \U$20640 ( \29062 , RIe1e5b40_6170);
or \U$20641 ( \29063 , \29062 , \28843 );
not \U$20642 ( \29064 , \28754 );
and \U$20643 ( \29065 , \27854 , \29064 );
not \U$20644 ( \29066 , \29065 );
not \U$20645 ( \29067 , \27851 );
not \U$20646 ( \29068 , \28659 );
or \U$20647 ( \29069 , \29067 , \29068 );
nand \U$20648 ( \29070 , \29063 , \29066 , \29069 );
and \U$20649 ( \29071 , \29070 , \28749 );
or \U$20650 ( \29072 , \29061 , \29071 );
and \U$20652 ( \29073 , \29072 , 1'b1 );
or \U$20654 ( \29074 , \29073 , 1'b0 );
buf \U$20655 ( \29075 , \29074 );
_DC r23d42_GF_IsGateDCbyConstraint ( \29076_nR23d42 , \29075 , \21944 );
buf \U$20656 ( \29077 , \29076_nR23d42 );
not \U$20657 ( \29078 , \28749 );
and \U$20658 ( \29079 , RIe1e88b8_6171, \29078 );
not \U$20659 ( \29080 , RIe1e88b8_6171);
or \U$20660 ( \29081 , \29080 , \28713 );
not \U$20661 ( \29082 , \28675 );
and \U$20662 ( \29083 , \27873 , \29082 );
not \U$20663 ( \29084 , \29083 );
not \U$20664 ( \29085 , \27870 );
not \U$20665 ( \29086 , \28929 );
or \U$20666 ( \29087 , \29085 , \29086 );
nand \U$20667 ( \29088 , \29081 , \29084 , \29087 );
and \U$20668 ( \29089 , \29088 , \28749 );
or \U$20669 ( \29090 , \29079 , \29089 );
and \U$20671 ( \29091 , \29090 , 1'b1 );
or \U$20673 ( \29092 , \29091 , 1'b0 );
buf \U$20674 ( \29093 , \29092 );
_DC r23d44_GF_IsGateDCbyConstraint ( \29094_nR23d44 , \29093 , \21944 );
buf \U$20675 ( \29095 , \29094_nR23d44 );
not \U$20676 ( \29096 , \28939 );
and \U$20677 ( \29097 , RIe1eb180_6172, \29096 );
not \U$20678 ( \29098 , RIe1eb180_6172);
or \U$20679 ( \29099 , \29098 , \28843 );
not \U$20680 ( \29100 , \28715 );
and \U$20681 ( \29101 , \27892 , \29100 );
not \U$20682 ( \29102 , \29101 );
not \U$20683 ( \29103 , \27889 );
not \U$20684 ( \29104 , \28659 );
or \U$20685 ( \29105 , \29103 , \29104 );
nand \U$20686 ( \29106 , \29099 , \29102 , \29105 );
and \U$20687 ( \29107 , \29106 , \28939 );
or \U$20688 ( \29108 , \29097 , \29107 );
and \U$20690 ( \29109 , \29108 , 1'b1 );
or \U$20692 ( \29110 , \29109 , 1'b0 );
buf \U$20693 ( \29111 , \29110 );
_DC r23d46_GF_IsGateDCbyConstraint ( \29112_nR23d46 , \29111 , \21944 );
buf \U$20694 ( \29113 , \29112_nR23d46 );
not \U$20695 ( \29114 , \28749 );
and \U$20696 ( \29115 , RIe1ee858_6173, \29114 );
not \U$20697 ( \29116 , RIe1ee858_6173);
or \U$20698 ( \29117 , \29116 , \28694 );
not \U$20699 ( \29118 , \28715 );
and \U$20700 ( \29119 , \27911 , \29118 );
not \U$20701 ( \29120 , \29119 );
not \U$20702 ( \29121 , \27908 );
not \U$20703 ( \29122 , \28929 );
or \U$20704 ( \29123 , \29121 , \29122 );
nand \U$20705 ( \29124 , \29117 , \29120 , \29123 );
and \U$20706 ( \29125 , \29124 , \28749 );
or \U$20707 ( \29126 , \29115 , \29125 );
and \U$20709 ( \29127 , \29126 , 1'b1 );
or \U$20711 ( \29128 , \29127 , 1'b0 );
buf \U$20712 ( \29129 , \29128 );
_DC r23d48_GF_IsGateDCbyConstraint ( \29130_nR23d48 , \29129 , \21944 );
buf \U$20713 ( \29131 , \29130_nR23d48 );
not \U$20714 ( \29132 , \28563 );
and \U$20715 ( \29133 , RIe1f1120_6174, \29132 );
not \U$20716 ( \29134 , RIe1f1120_6174);
or \U$20717 ( \29135 , \29134 , \28713 );
not \U$20718 ( \29136 , \28773 );
and \U$20719 ( \29137 , \27930 , \29136 );
not \U$20720 ( \29138 , \29137 );
not \U$20721 ( \29139 , \27927 );
not \U$20722 ( \29140 , \28738 );
or \U$20723 ( \29141 , \29139 , \29140 );
nand \U$20724 ( \29142 , \29135 , \29138 , \29141 );
and \U$20725 ( \29143 , \29142 , \28563 );
or \U$20726 ( \29144 , \29133 , \29143 );
and \U$20728 ( \29145 , \29144 , 1'b1 );
or \U$20730 ( \29146 , \29145 , 1'b0 );
buf \U$20731 ( \29147 , \29146 );
_DC r23d4a_GF_IsGateDCbyConstraint ( \29148_nR23d4a , \29147 , \21944 );
buf \U$20732 ( \29149 , \29148_nR23d4a );
not \U$20733 ( \29150 , \28939 );
and \U$20734 ( \29151 , RIe1f47f8_6175, \29150 );
not \U$20735 ( \29152 , RIe1f47f8_6175);
or \U$20736 ( \29153 , \29152 , \28694 );
not \U$20737 ( \29154 , \28715 );
and \U$20738 ( \29155 , \27949 , \29154 );
not \U$20739 ( \29156 , \29155 );
not \U$20740 ( \29157 , \27947 );
not \U$20741 ( \29158 , \28929 );
or \U$20742 ( \29159 , \29157 , \29158 );
nand \U$20743 ( \29160 , \29153 , \29156 , \29159 );
and \U$20744 ( \29161 , \29160 , \28939 );
or \U$20745 ( \29162 , \29151 , \29161 );
and \U$20747 ( \29163 , \29162 , 1'b1 );
or \U$20749 ( \29164 , \29163 , 1'b0 );
buf \U$20750 ( \29165 , \29164 );
_DC r23d4c_GF_IsGateDCbyConstraint ( \29166_nR23d4c , \29165 , \21944 );
buf \U$20751 ( \29167 , \29166_nR23d4c );
not \U$20752 ( \29168 , \28749 );
and \U$20753 ( \29169 , RIe1f70c0_6176, \29168 );
not \U$20754 ( \29170 , RIe1f70c0_6176);
or \U$20755 ( \29171 , \29170 , \28713 );
not \U$20756 ( \29172 , \28675 );
and \U$20757 ( \29173 , \27968 , \29172 );
not \U$20758 ( \29174 , \29173 );
not \U$20759 ( \29175 , \27966 );
not \U$20760 ( \29176 , \28659 );
or \U$20761 ( \29177 , \29175 , \29176 );
nand \U$20762 ( \29178 , \29171 , \29174 , \29177 );
and \U$20763 ( \29179 , \29178 , \28749 );
or \U$20764 ( \29180 , \29169 , \29179 );
and \U$20766 ( \29181 , \29180 , 1'b1 );
or \U$20768 ( \29182 , \29181 , 1'b0 );
buf \U$20769 ( \29183 , \29182 );
_DC r23d4e_GF_IsGateDCbyConstraint ( \29184_nR23d4e , \29183 , \21944 );
buf \U$20770 ( \29185 , \29184_nR23d4e );
not \U$20771 ( \29186 , \28749 );
and \U$20772 ( \29187 , RIe1fa180_6177, \29186 );
not \U$20773 ( \29188 , RIe1fa180_6177);
or \U$20774 ( \29189 , \29188 , \28843 );
not \U$20775 ( \29190 , \28754 );
and \U$20776 ( \29191 , \27988 , \29190 );
not \U$20777 ( \29192 , \29191 );
not \U$20778 ( \29193 , \27985 );
not \U$20779 ( \29194 , \28929 );
or \U$20780 ( \29195 , \29193 , \29194 );
nand \U$20781 ( \29196 , \29189 , \29192 , \29195 );
and \U$20782 ( \29197 , \29196 , \28749 );
or \U$20783 ( \29198 , \29187 , \29197 );
and \U$20785 ( \29199 , \29198 , 1'b1 );
or \U$20787 ( \29200 , \29199 , 1'b0 );
buf \U$20788 ( \29201 , \29200 );
_DC r23d52_GF_IsGateDCbyConstraint ( \29202_nR23d52 , \29201 , \21944 );
buf \U$20789 ( \29203 , \29202_nR23d52 );
not \U$20790 ( \29204 , \28939 );
and \U$20791 ( \29205 , RIe1fbad0_6178, \29204 );
not \U$20792 ( \29206 , RIe1fbad0_6178);
or \U$20793 ( \29207 , \29206 , \28673 );
not \U$20794 ( \29208 , \28653 );
and \U$20795 ( \29209 , \28009 , \29208 );
not \U$20796 ( \29210 , \29209 );
not \U$20797 ( \29211 , \28006 );
not \U$20798 ( \29212 , \28659 );
or \U$20799 ( \29213 , \29211 , \29212 );
nand \U$20800 ( \29214 , \29207 , \29210 , \29213 );
and \U$20801 ( \29215 , \29214 , \28939 );
or \U$20802 ( \29216 , \29205 , \29215 );
and \U$20804 ( \29217 , \29216 , 1'b1 );
or \U$20806 ( \29218 , \29217 , 1'b0 );
buf \U$20807 ( \29219 , \29218 );
_DC r23d54_GF_IsGateDCbyConstraint ( \29220_nR23d54 , \29219 , \21944 );
buf \U$20808 ( \29221 , \29220_nR23d54 );
not \U$20809 ( \29222 , \28563 );
and \U$20810 ( \29223 , RIe1fd330_6179, \29222 );
not \U$20811 ( \29224 , RIe1fd330_6179);
or \U$20812 ( \29225 , \29224 , \28673 );
not \U$20813 ( \29226 , \28754 );
and \U$20814 ( \29227 , \28029 , \29226 );
not \U$20815 ( \29228 , \29227 );
not \U$20816 ( \29229 , \28026 );
not \U$20817 ( \29230 , \28929 );
or \U$20818 ( \29231 , \29229 , \29230 );
nand \U$20819 ( \29232 , \29225 , \29228 , \29231 );
and \U$20820 ( \29233 , \29232 , \28563 );
or \U$20821 ( \29234 , \29223 , \29233 );
and \U$20823 ( \29235 , \29234 , 1'b1 );
or \U$20825 ( \29236 , \29235 , 1'b0 );
buf \U$20826 ( \29237 , \29236 );
_DC r23d56_GF_IsGateDCbyConstraint ( \29238_nR23d56 , \29237 , \21944 );
buf \U$20827 ( \29239 , \29238_nR23d56 );
not \U$20828 ( \29240 , \28563 );
and \U$20829 ( \29241 , RIe1ff568_6180, \29240 );
not \U$20830 ( \29242 , RIe1ff568_6180);
or \U$20831 ( \29243 , \29242 , \28694 );
not \U$20832 ( \29244 , \28653 );
and \U$20833 ( \29245 , \28048 , \29244 );
not \U$20834 ( \29246 , \29245 );
not \U$20835 ( \29247 , \28045 );
not \U$20836 ( \29248 , \28659 );
or \U$20837 ( \29249 , \29247 , \29248 );
nand \U$20838 ( \29250 , \29243 , \29246 , \29249 );
and \U$20839 ( \29251 , \29250 , \28563 );
or \U$20840 ( \29252 , \29241 , \29251 );
and \U$20842 ( \29253 , \29252 , 1'b1 );
or \U$20844 ( \29254 , \29253 , 1'b0 );
buf \U$20845 ( \29255 , \29254 );
_DC r23d58_GF_IsGateDCbyConstraint ( \29256_nR23d58 , \29255 , \21944 );
buf \U$20846 ( \29257 , \29256_nR23d58 );
not \U$20847 ( \29258 , \28939 );
and \U$20848 ( \29259 , RIe2012f0_6181, \29258 );
not \U$20849 ( \29260 , RIe2012f0_6181);
or \U$20850 ( \29261 , \29260 , \28651 );
not \U$20851 ( \29262 , \28653 );
and \U$20852 ( \29263 , \28066 , \29262 );
not \U$20853 ( \29264 , \29263 );
not \U$20854 ( \29265 , \28064 );
not \U$20855 ( \29266 , \28659 );
or \U$20856 ( \29267 , \29265 , \29266 );
nand \U$20857 ( \29268 , \29261 , \29264 , \29267 );
and \U$20858 ( \29269 , \29268 , \28939 );
or \U$20859 ( \29270 , \29259 , \29269 );
and \U$20861 ( \29271 , \29270 , 1'b1 );
or \U$20863 ( \29272 , \29271 , 1'b0 );
buf \U$20864 ( \29273 , \29272 );
_DC r23d5a_GF_IsGateDCbyConstraint ( \29274_nR23d5a , \29273 , \21944 );
buf \U$20865 ( \29275 , \29274_nR23d5a );
not \U$20866 ( \29276 , \28749 );
and \U$20867 ( \29277 , RIe203000_6182, \29276 );
not \U$20868 ( \29278 , RIe203000_6182);
or \U$20869 ( \29279 , \29278 , \28694 );
not \U$20870 ( \29280 , \28773 );
and \U$20871 ( \29281 , \28085 , \29280 );
not \U$20872 ( \29282 , \29281 );
not \U$20873 ( \29283 , \28082 );
not \U$20874 ( \29284 , \28929 );
or \U$20875 ( \29285 , \29283 , \29284 );
nand \U$20876 ( \29286 , \29279 , \29282 , \29285 );
and \U$20877 ( \29287 , \29286 , \28749 );
or \U$20878 ( \29288 , \29277 , \29287 );
and \U$20880 ( \29289 , \29288 , 1'b1 );
or \U$20882 ( \29290 , \29289 , 1'b0 );
buf \U$20883 ( \29291 , \29290 );
_DC r23d5c_GF_IsGateDCbyConstraint ( \29292_nR23d5c , \29291 , \21944 );
buf \U$20884 ( \29293 , \29292_nR23d5c );
buf \U$20885 ( \29294 , \28307 );
not \U$20886 ( \29295 , \29294 );
and \U$20887 ( \29296 , RIe203f00_6183, \29295 );
not \U$20888 ( \29297 , RIe203f00_6183);
or \U$20889 ( \29298 , \29297 , \28713 );
not \U$20890 ( \29299 , \28675 );
and \U$20891 ( \29300 , \28104 , \29299 );
not \U$20892 ( \29301 , \29300 );
not \U$20893 ( \29302 , \28101 );
not \U$20894 ( \29303 , \28929 );
or \U$20895 ( \29304 , \29302 , \29303 );
nand \U$20896 ( \29305 , \29298 , \29301 , \29304 );
and \U$20897 ( \29306 , \29305 , \29294 );
or \U$20898 ( \29307 , \29296 , \29306 );
and \U$20900 ( \29308 , \29307 , 1'b1 );
or \U$20902 ( \29309 , \29308 , 1'b0 );
buf \U$20903 ( \29310 , \29309 );
_DC r23d5e_GF_IsGateDCbyConstraint ( \29311_nR23d5e , \29310 , \21944 );
buf \U$20904 ( \29312 , \29311_nR23d5e );
not \U$20905 ( \29313 , \28939 );
and \U$20906 ( \29314 , RIe2053a0_6184, \29313 );
not \U$20907 ( \29315 , RIe2053a0_6184);
or \U$20908 ( \29316 , \29315 , \28694 );
not \U$20909 ( \29317 , \28653 );
and \U$20910 ( \29318 , \28123 , \29317 );
not \U$20911 ( \29319 , \29318 );
nand \U$20912 ( \29320 , \28120 , \28929 );
nand \U$20913 ( \29321 , \29316 , \29319 , \29320 );
and \U$20914 ( \29322 , \29321 , \28939 );
or \U$20915 ( \29323 , \29314 , \29322 );
and \U$20917 ( \29324 , \29323 , 1'b1 );
or \U$20919 ( \29325 , \29324 , 1'b0 );
buf \U$20920 ( \29326 , \29325 );
_DC r23d60_GF_IsGateDCbyConstraint ( \29327_nR23d60 , \29326 , \21944 );
buf \U$20921 ( \29328 , \29327_nR23d60 );
buf \U$20922 ( \29329 , \27363 );
buf \U$20923 ( \29330 , \29329 );
not \U$20924 ( \29331 , \29330 );
and \U$20925 ( \29332 , RIe2066d8_6185, \29331 );
not \U$20926 ( \29333 , RIe2066d8_6185);
or \U$20927 ( \29334 , \29333 , \28673 );
not \U$20928 ( \29335 , \28653 );
and \U$20929 ( \29336 , \28142 , \29335 );
not \U$20930 ( \29337 , \29336 );
nand \U$20931 ( \29338 , \28139 , \28680 );
nand \U$20932 ( \29339 , \29334 , \29337 , \29338 );
and \U$20933 ( \29340 , \29339 , \29330 );
or \U$20934 ( \29341 , \29332 , \29340 );
and \U$20936 ( \29342 , \29341 , 1'b1 );
or \U$20938 ( \29343 , \29342 , 1'b0 );
buf \U$20939 ( \29344 , \29343 );
_DC r23d62_GF_IsGateDCbyConstraint ( \29345_nR23d62 , \29344 , \21944 );
buf \U$20940 ( \29346 , \29345_nR23d62 );
not \U$20941 ( \29347 , \29330 );
and \U$20942 ( \29348 , RIe207920_6186, \29347 );
not \U$20943 ( \29349 , RIe207920_6186);
or \U$20944 ( \29350 , \29349 , \28843 );
not \U$20945 ( \29351 , \28773 );
and \U$20946 ( \29352 , \28161 , \29351 );
not \U$20947 ( \29353 , \29352 );
nand \U$20948 ( \29354 , \28158 , \28659 );
nand \U$20949 ( \29355 , \29350 , \29353 , \29354 );
and \U$20950 ( \29356 , \29355 , \29330 );
or \U$20951 ( \29357 , \29348 , \29356 );
and \U$20953 ( \29358 , \29357 , 1'b1 );
or \U$20955 ( \29359 , \29358 , 1'b0 );
buf \U$20956 ( \29360 , \29359 );
_DC r23d64_GF_IsGateDCbyConstraint ( \29361_nR23d64 , \29360 , \21944 );
buf \U$20957 ( \29362 , \29361_nR23d64 );
not \U$20958 ( \29363 , \28939 );
and \U$20959 ( \29364 , RIe208be0_6187, \29363 );
not \U$20960 ( \29365 , RIe208be0_6187);
or \U$20961 ( \29366 , \29365 , \28843 );
not \U$20962 ( \29367 , \28715 );
and \U$20963 ( \29368 , \28180 , \29367 );
not \U$20964 ( \29369 , \29368 );
nand \U$20965 ( \29370 , \28177 , \28929 );
nand \U$20966 ( \29371 , \29366 , \29369 , \29370 );
and \U$20967 ( \29372 , \29371 , \28939 );
or \U$20968 ( \29373 , \29364 , \29372 );
and \U$20970 ( \29374 , \29373 , 1'b1 );
or \U$20972 ( \29375 , \29374 , 1'b0 );
buf \U$20973 ( \29376 , \29375 );
_DC r23d68_GF_IsGateDCbyConstraint ( \29377_nR23d68 , \29376 , \21944 );
buf \U$20974 ( \29378 , \29377_nR23d68 );
not \U$20975 ( \29379 , \29294 );
and \U$20976 ( \29380 , RIe209d38_6188, \29379 );
not \U$20977 ( \29381 , RIe209d38_6188);
or \U$20978 ( \29382 , \29381 , \28651 );
not \U$20979 ( \29383 , \28754 );
and \U$20980 ( \29384 , \28199 , \29383 );
not \U$20981 ( \29385 , \29384 );
nand \U$20982 ( \29386 , \28196 , \28929 );
nand \U$20983 ( \29387 , \29382 , \29385 , \29386 );
and \U$20984 ( \29388 , \29387 , \29294 );
or \U$20985 ( \29389 , \29380 , \29388 );
and \U$20987 ( \29390 , \29389 , 1'b1 );
or \U$20989 ( \29391 , \29390 , 1'b0 );
buf \U$20990 ( \29392 , \29391 );
_DC r23d6a_GF_IsGateDCbyConstraint ( \29393_nR23d6a , \29392 , \21944 );
buf \U$20991 ( \29394 , \29393_nR23d6a );
not \U$20992 ( \29395 , \29330 );
and \U$20993 ( \29396 , RIe20b958_6189, \29395 );
not \U$20994 ( \29397 , RIe20b958_6189);
or \U$20995 ( \29398 , \29397 , \28673 );
not \U$20996 ( \29399 , \28675 );
and \U$20997 ( \29400 , \28218 , \29399 );
not \U$20998 ( \29401 , \29400 );
nand \U$20999 ( \29402 , \28215 , \28680 );
nand \U$21000 ( \29403 , \29398 , \29401 , \29402 );
and \U$21001 ( \29404 , \29403 , \29330 );
or \U$21002 ( \29405 , \29396 , \29404 );
and \U$21004 ( \29406 , \29405 , 1'b1 );
or \U$21006 ( \29407 , \29406 , 1'b0 );
buf \U$21007 ( \29408 , \29407 );
_DC r23d6c_GF_IsGateDCbyConstraint ( \29409_nR23d6c , \29408 , \21944 );
buf \U$21008 ( \29410 , \29409_nR23d6c );
not \U$21009 ( \29411 , \28939 );
and \U$21010 ( \29412 , RIe20cf60_6190, \29411 );
not \U$21011 ( \29413 , RIe20cf60_6190);
or \U$21012 ( \29414 , \29413 , \28673 );
not \U$21013 ( \29415 , \28715 );
and \U$21014 ( \29416 , \28237 , \29415 );
not \U$21015 ( \29417 , \29416 );
nand \U$21016 ( \29418 , \28235 , \28680 );
nand \U$21017 ( \29419 , \29414 , \29417 , \29418 );
and \U$21018 ( \29420 , \29419 , \28939 );
or \U$21019 ( \29421 , \29412 , \29420 );
and \U$21021 ( \29422 , \29421 , 1'b1 );
or \U$21023 ( \29423 , \29422 , 1'b0 );
buf \U$21024 ( \29424 , \29423 );
_DC r23d6e_GF_IsGateDCbyConstraint ( \29425_nR23d6e , \29424 , \21944 );
buf \U$21025 ( \29426 , \29425_nR23d6e );
not \U$21026 ( \29427 , \29330 );
and \U$21027 ( \29428 , RIe20e4f0_6191, \29427 );
not \U$21028 ( \29429 , RIe20e4f0_6191);
or \U$21029 ( \29430 , \29429 , \28713 );
not \U$21030 ( \29431 , \28675 );
and \U$21031 ( \29432 , \28257 , \29431 );
not \U$21032 ( \29433 , \29432 );
not \U$21033 ( \29434 , \28254 );
not \U$21034 ( \29435 , \28738 );
or \U$21035 ( \29436 , \29434 , \29435 );
nand \U$21036 ( \29437 , \29430 , \29433 , \29436 );
and \U$21037 ( \29438 , \29437 , \29330 );
or \U$21038 ( \29439 , \29428 , \29438 );
and \U$21040 ( \29440 , \29439 , 1'b1 );
or \U$21042 ( \29441 , \29440 , 1'b0 );
buf \U$21043 ( \29442 , \29441 );
_DC r23d70_GF_IsGateDCbyConstraint ( \29443_nR23d70 , \29442 , \21944 );
buf \U$21044 ( \29444 , \29443_nR23d70 );
not \U$21045 ( \29445 , \29330 );
and \U$21046 ( \29446 , RIe20f5d0_6192, \29445 );
not \U$21047 ( \29447 , RIe20f5d0_6192);
or \U$21048 ( \29448 , \29447 , \28651 );
not \U$21049 ( \29449 , \28754 );
and \U$21050 ( \29450 , \28276 , \29449 );
not \U$21051 ( \29451 , \29450 );
not \U$21052 ( \29452 , \28273 );
not \U$21053 ( \29453 , \28929 );
or \U$21054 ( \29454 , \29452 , \29453 );
nand \U$21055 ( \29455 , \29448 , \29451 , \29454 );
and \U$21056 ( \29456 , \29455 , \29330 );
or \U$21057 ( \29457 , \29446 , \29456 );
and \U$21059 ( \29458 , \29457 , 1'b1 );
or \U$21061 ( \29459 , \29458 , 1'b0 );
buf \U$21062 ( \29460 , \29459 );
_DC r23d72_GF_IsGateDCbyConstraint ( \29461_nR23d72 , \29460 , \21944 );
buf \U$21063 ( \29462 , \29461_nR23d72 );
not \U$21064 ( \29463 , \28939 );
and \U$21065 ( \29464 , RIe211178_6193, \29463 );
not \U$21066 ( \29465 , RIe211178_6193);
or \U$21067 ( \29466 , \29465 , \28843 );
not \U$21068 ( \29467 , \28754 );
and \U$21069 ( \29468 , \28295 , \29467 );
not \U$21070 ( \29469 , \29468 );
not \U$21071 ( \29470 , \28292 );
not \U$21072 ( \29471 , \28738 );
or \U$21073 ( \29472 , \29470 , \29471 );
nand \U$21074 ( \29473 , \29466 , \29469 , \29472 );
and \U$21075 ( \29474 , \29473 , \28939 );
or \U$21076 ( \29475 , \29464 , \29474 );
and \U$21078 ( \29476 , \29475 , 1'b1 );
or \U$21080 ( \29477 , \29476 , 1'b0 );
buf \U$21081 ( \29478 , \29477 );
_DC r23d74_GF_IsGateDCbyConstraint ( \29479_nR23d74 , \29478 , \21944 );
buf \U$21082 ( \29480 , \29479_nR23d74 );
not \U$21083 ( \29481 , \29294 );
and \U$21084 ( \29482 , RIe212c30_6194, \29481 );
not \U$21085 ( \29483 , RIe212c30_6194);
or \U$21086 ( \29484 , \29483 , \28694 );
not \U$21087 ( \29485 , \28675 );
and \U$21088 ( \29486 , \28314 , \29485 );
not \U$21089 ( \29487 , \29486 );
not \U$21090 ( \29488 , \28312 );
not \U$21091 ( \29489 , \28929 );
or \U$21092 ( \29490 , \29488 , \29489 );
nand \U$21093 ( \29491 , \29484 , \29487 , \29490 );
and \U$21094 ( \29492 , \29491 , \29294 );
or \U$21095 ( \29493 , \29482 , \29492 );
and \U$21097 ( \29494 , \29493 , 1'b1 );
or \U$21099 ( \29495 , \29494 , 1'b0 );
buf \U$21100 ( \29496 , \29495 );
_DC r23d76_GF_IsGateDCbyConstraint ( \29497_nR23d76 , \29496 , \21944 );
buf \U$21101 ( \29498 , \29497_nR23d76 );
not \U$21102 ( \29499 , \29294 );
and \U$21103 ( \29500 , RIe214148_6195, \29499 );
not \U$21104 ( \29501 , RIe214148_6195);
or \U$21105 ( \29502 , \29501 , \28651 );
not \U$21106 ( \29503 , \28715 );
and \U$21107 ( \29504 , \28333 , \29503 );
not \U$21108 ( \29505 , \29504 );
not \U$21109 ( \29506 , \28330 );
not \U$21110 ( \29507 , \28680 );
or \U$21111 ( \29508 , \29506 , \29507 );
nand \U$21112 ( \29509 , \29502 , \29505 , \29508 );
and \U$21113 ( \29510 , \29509 , \29294 );
or \U$21114 ( \29511 , \29500 , \29510 );
and \U$21116 ( \29512 , \29511 , 1'b1 );
or \U$21118 ( \29513 , \29512 , 1'b0 );
buf \U$21119 ( \29514 , \29513 );
_DC r23d78_GF_IsGateDCbyConstraint ( \29515_nR23d78 , \29514 , \21944 );
buf \U$21120 ( \29516 , \29515_nR23d78 );
not \U$21121 ( \29517 , \28939 );
and \U$21122 ( \29518 , RIe215c00_6196, \29517 );
not \U$21123 ( \29519 , RIe215c00_6196);
or \U$21124 ( \29520 , \29519 , \28673 );
not \U$21125 ( \29521 , \28675 );
and \U$21126 ( \29522 , \28352 , \29521 );
not \U$21127 ( \29523 , \29522 );
not \U$21128 ( \29524 , \28349 );
not \U$21129 ( \29525 , \28738 );
or \U$21130 ( \29526 , \29524 , \29525 );
nand \U$21131 ( \29527 , \29520 , \29523 , \29526 );
and \U$21132 ( \29528 , \29527 , \28939 );
or \U$21133 ( \29529 , \29518 , \29528 );
and \U$21135 ( \29530 , \29529 , 1'b1 );
or \U$21137 ( \29531 , \29530 , 1'b0 );
buf \U$21138 ( \29532 , \29531 );
_DC r23d7a_GF_IsGateDCbyConstraint ( \29533_nR23d7a , \29532 , \21944 );
buf \U$21139 ( \29534 , \29533_nR23d7a );
not \U$21140 ( \29535 , \29294 );
and \U$21141 ( \29536 , RIe217460_6197, \29535 );
not \U$21142 ( \29537 , RIe217460_6197);
or \U$21143 ( \29538 , \29537 , \28694 );
not \U$21144 ( \29539 , \28754 );
and \U$21145 ( \29540 , \28372 , \29539 );
not \U$21146 ( \29541 , \29540 );
not \U$21147 ( \29542 , \28369 );
not \U$21148 ( \29543 , \28680 );
or \U$21149 ( \29544 , \29542 , \29543 );
nand \U$21150 ( \29545 , \29538 , \29541 , \29544 );
and \U$21151 ( \29546 , \29545 , \29294 );
or \U$21152 ( \29547 , \29536 , \29546 );
and \U$21154 ( \29548 , \29547 , 1'b1 );
or \U$21156 ( \29549 , \29548 , 1'b0 );
buf \U$21157 ( \29550 , \29549 );
_DC r23d7e_GF_IsGateDCbyConstraint ( \29551_nR23d7e , \29550 , \21944 );
buf \U$21158 ( \29552 , \29551_nR23d7e );
not \U$21159 ( \29553 , \29330 );
and \U$21160 ( \29554 , RIe218798_6198, \29553 );
not \U$21161 ( \29555 , RIe218798_6198);
or \U$21162 ( \29556 , \29555 , \28713 );
not \U$21163 ( \29557 , \28653 );
and \U$21164 ( \29558 , \28392 , \29557 );
not \U$21165 ( \29559 , \29558 );
not \U$21166 ( \29560 , \28389 );
not \U$21167 ( \29561 , \28738 );
or \U$21168 ( \29562 , \29560 , \29561 );
nand \U$21169 ( \29563 , \29556 , \29559 , \29562 );
and \U$21170 ( \29564 , \29563 , \29330 );
or \U$21171 ( \29565 , \29554 , \29564 );
and \U$21173 ( \29566 , \29565 , 1'b1 );
or \U$21175 ( \29567 , \29566 , 1'b0 );
buf \U$21176 ( \29568 , \29567 );
_DC r23d80_GF_IsGateDCbyConstraint ( \29569_nR23d80 , \29568 , \21944 );
buf \U$21177 ( \29570 , \29569_nR23d80 );
buf \U$21178 ( \29571 , \27363 );
not \U$21179 ( \29572 , \29571 );
and \U$21180 ( \29573 , RIe2199e0_6199, \29572 );
not \U$21181 ( \29574 , RIe2199e0_6199);
or \U$21182 ( \29575 , \29574 , \28651 );
not \U$21183 ( \29576 , \28653 );
and \U$21184 ( \29577 , \28412 , \29576 );
not \U$21185 ( \29578 , \29577 );
not \U$21186 ( \29579 , \28409 );
not \U$21187 ( \29580 , \28680 );
or \U$21188 ( \29581 , \29579 , \29580 );
nand \U$21189 ( \29582 , \29575 , \29578 , \29581 );
and \U$21190 ( \29583 , \29582 , \29571 );
or \U$21191 ( \29584 , \29573 , \29583 );
and \U$21193 ( \29585 , \29584 , 1'b1 );
or \U$21195 ( \29586 , \29585 , 1'b0 );
buf \U$21196 ( \29587 , \29586 );
_DC r23d82_GF_IsGateDCbyConstraint ( \29588_nR23d82 , \29587 , \21944 );
buf \U$21197 ( \29589 , \29588_nR23d82 );
not \U$21198 ( \29590 , \29294 );
and \U$21199 ( \29591 , RIe14e868_6200, \29590 );
not \U$21200 ( \29592 , RIe14e868_6200);
or \U$21201 ( \29593 , \29592 , \28651 );
not \U$21202 ( \29594 , \28773 );
and \U$21203 ( \29595 , \28432 , \29594 );
not \U$21204 ( \29596 , \29595 );
not \U$21205 ( \29597 , \28429 );
not \U$21206 ( \29598 , \28680 );
or \U$21207 ( \29599 , \29597 , \29598 );
nand \U$21208 ( \29600 , \29593 , \29596 , \29599 );
and \U$21209 ( \29601 , \29600 , \29294 );
or \U$21210 ( \29602 , \29591 , \29601 );
and \U$21212 ( \29603 , \29602 , 1'b1 );
or \U$21214 ( \29604 , \29603 , 1'b0 );
buf \U$21215 ( \29605 , \29604 );
_DC r23d84_GF_IsGateDCbyConstraint ( \29606_nR23d84 , \29605 , \21944 );
buf \U$21216 ( \29607 , \29606_nR23d84 );
not \U$21217 ( \29608 , \29294 );
and \U$21218 ( \29609 , RIe151130_6201, \29608 );
not \U$21219 ( \29610 , RIe151130_6201);
or \U$21220 ( \29611 , \29610 , \28843 );
not \U$21221 ( \29612 , \28653 );
and \U$21222 ( \29613 , \28452 , \29612 );
not \U$21223 ( \29614 , \29613 );
not \U$21224 ( \29615 , \28449 );
not \U$21225 ( \29616 , \28738 );
or \U$21226 ( \29617 , \29615 , \29616 );
nand \U$21227 ( \29618 , \29611 , \29614 , \29617 );
and \U$21228 ( \29619 , \29618 , \29294 );
or \U$21229 ( \29620 , \29609 , \29619 );
and \U$21231 ( \29621 , \29620 , 1'b1 );
or \U$21233 ( \29622 , \29621 , 1'b0 );
buf \U$21234 ( \29623 , \29622 );
_DC r23d86_GF_IsGateDCbyConstraint ( \29624_nR23d86 , \29623 , \21944 );
buf \U$21235 ( \29625 , \29624_nR23d86 );
not \U$21236 ( \29626 , \29571 );
and \U$21237 ( \29627 , RIe153020_6202, \29626 );
not \U$21238 ( \29628 , RIe153020_6202);
or \U$21239 ( \29629 , \29628 , \28843 );
not \U$21240 ( \29630 , \28675 );
and \U$21241 ( \29631 , \28471 , \29630 );
not \U$21242 ( \29632 , \29631 );
not \U$21243 ( \29633 , \28468 );
not \U$21244 ( \29634 , \28738 );
or \U$21245 ( \29635 , \29633 , \29634 );
nand \U$21246 ( \29636 , \29629 , \29632 , \29635 );
and \U$21247 ( \29637 , \29636 , \29571 );
or \U$21248 ( \29638 , \29627 , \29637 );
and \U$21250 ( \29639 , \29638 , 1'b1 );
or \U$21252 ( \29640 , \29639 , 1'b0 );
buf \U$21253 ( \29641 , \29640 );
_DC r23d88_GF_IsGateDCbyConstraint ( \29642_nR23d88 , \29641 , \21944 );
buf \U$21254 ( \29643 , \29642_nR23d88 );
not \U$21255 ( \29644 , \29330 );
and \U$21256 ( \29645 , RIe154ad8_6203, \29644 );
not \U$21257 ( \29646 , RIe154ad8_6203);
or \U$21258 ( \29647 , \29646 , \28694 );
not \U$21259 ( \29648 , \28754 );
and \U$21260 ( \29649 , \28490 , \29648 );
not \U$21261 ( \29650 , \29649 );
not \U$21262 ( \29651 , \28488 );
not \U$21263 ( \29652 , \28680 );
or \U$21264 ( \29653 , \29651 , \29652 );
nand \U$21265 ( \29654 , \29647 , \29650 , \29653 );
and \U$21266 ( \29655 , \29654 , \29330 );
or \U$21267 ( \29656 , \29645 , \29655 );
and \U$21269 ( \29657 , \29656 , 1'b1 );
or \U$21271 ( \29658 , \29657 , 1'b0 );
buf \U$21272 ( \29659 , \29658 );
_DC r23d8a_GF_IsGateDCbyConstraint ( \29660_nR23d8a , \29659 , \21944 );
buf \U$21273 ( \29661 , \29660_nR23d8a );
not \U$21274 ( \29662 , \29330 );
and \U$21275 ( \29663 , RIe156518_6204, \29662 );
not \U$21276 ( \29664 , RIe156518_6204);
or \U$21277 ( \29665 , \29664 , \28713 );
not \U$21278 ( \29666 , \28653 );
and \U$21279 ( \29667 , \28510 , \29666 );
not \U$21280 ( \29668 , \29667 );
not \U$21281 ( \29669 , \28507 );
not \U$21282 ( \29670 , \28738 );
or \U$21283 ( \29671 , \29669 , \29670 );
nand \U$21284 ( \29672 , \29665 , \29668 , \29671 );
and \U$21285 ( \29673 , \29672 , \29330 );
or \U$21286 ( \29674 , \29663 , \29673 );
and \U$21288 ( \29675 , \29674 , 1'b1 );
or \U$21290 ( \29676 , \29675 , 1'b0 );
buf \U$21291 ( \29677 , \29676 );
_DC r23d8c_GF_IsGateDCbyConstraint ( \29678_nR23d8c , \29677 , \21944 );
buf \U$21292 ( \29679 , \29678_nR23d8c );
not \U$21293 ( \29680 , \29571 );
and \U$21294 ( \29681 , RIe158228_6205, \29680 );
not \U$21295 ( \29682 , RIe158228_6205);
or \U$21296 ( \29683 , \29682 , \28713 );
not \U$21297 ( \29684 , \28653 );
and \U$21298 ( \29685 , \28529 , \29684 );
not \U$21299 ( \29686 , \29685 );
not \U$21300 ( \29687 , \28526 );
not \U$21301 ( \29688 , \28680 );
or \U$21302 ( \29689 , \29687 , \29688 );
nand \U$21303 ( \29690 , \29683 , \29686 , \29689 );
and \U$21304 ( \29691 , \29690 , \29571 );
or \U$21305 ( \29692 , \29681 , \29691 );
and \U$21307 ( \29693 , \29692 , 1'b1 );
or \U$21309 ( \29694 , \29693 , 1'b0 );
buf \U$21310 ( \29695 , \29694 );
_DC r23d8e_GF_IsGateDCbyConstraint ( \29696_nR23d8e , \29695 , \21944 );
buf \U$21311 ( \29697 , \29696_nR23d8e );
not \U$21312 ( \29698 , \29294 );
and \U$21313 ( \29699 , RIe15a280_6206, \29698 );
not \U$21314 ( \29700 , RIe15a280_6206);
or \U$21315 ( \29701 , \29700 , \28843 );
not \U$21316 ( \29702 , \28715 );
and \U$21317 ( \29703 , \28551 , \29702 );
not \U$21318 ( \29704 , \29703 );
not \U$21319 ( \29705 , \28548 );
not \U$21320 ( \29706 , \28680 );
or \U$21321 ( \29707 , \29705 , \29706 );
nand \U$21322 ( \29708 , \29701 , \29704 , \29707 );
and \U$21323 ( \29709 , \29708 , \29294 );
or \U$21324 ( \29710 , \29699 , \29709 );
and \U$21326 ( \29711 , \29710 , 1'b1 );
or \U$21328 ( \29712 , \29711 , 1'b0 );
buf \U$21329 ( \29713 , \29712 );
_DC r23d90_GF_IsGateDCbyConstraint ( \29714_nR23d90 , \29713 , \21944 );
buf \U$21330 ( \29715 , \29714_nR23d90 );
not \U$21331 ( \29716 , \29294 );
and \U$21332 ( \29717 , RIe15c3c8_6207, \29716 );
not \U$21333 ( \29718 , RIe15c3c8_6207);
or \U$21334 ( \29719 , \29718 , \28694 );
not \U$21335 ( \29720 , \28675 );
and \U$21336 ( \29721 , \28571 , \29720 );
not \U$21337 ( \29722 , \29721 );
not \U$21338 ( \29723 , \28569 );
not \U$21339 ( \29724 , \28738 );
or \U$21340 ( \29725 , \29723 , \29724 );
nand \U$21341 ( \29726 , \29719 , \29722 , \29725 );
and \U$21342 ( \29727 , \29726 , \29294 );
or \U$21343 ( \29728 , \29717 , \29727 );
and \U$21345 ( \29729 , \29728 , 1'b1 );
or \U$21347 ( \29730 , \29729 , 1'b0 );
buf \U$21348 ( \29731 , \29730 );
_DC r23d94_GF_IsGateDCbyConstraint ( \29732_nR23d94 , \29731 , \21944 );
buf \U$21349 ( \29733 , \29732_nR23d94 );
not \U$21350 ( \29734 , \29571 );
and \U$21351 ( \29735 , RIe15ef60_6208, \29734 );
not \U$21352 ( \29736 , RIe15ef60_6208);
or \U$21353 ( \29737 , \29736 , \28673 );
not \U$21354 ( \29738 , \28715 );
and \U$21355 ( \29739 , \28589 , \29738 );
not \U$21356 ( \29740 , \29739 );
not \U$21357 ( \29741 , \28587 );
not \U$21358 ( \29742 , \28680 );
or \U$21359 ( \29743 , \29741 , \29742 );
nand \U$21360 ( \29744 , \29737 , \29740 , \29743 );
and \U$21361 ( \29745 , \29744 , \29571 );
or \U$21362 ( \29746 , \29735 , \29745 );
and \U$21364 ( \29747 , \29746 , 1'b1 );
or \U$21366 ( \29748 , \29747 , 1'b0 );
buf \U$21367 ( \29749 , \29748 );
_DC r23d96_GF_IsGateDCbyConstraint ( \29750_nR23d96 , \29749 , \21944 );
buf \U$21368 ( \29751 , \29750_nR23d96 );
not \U$21369 ( \29752 , \29330 );
and \U$21370 ( \29753 , RIe1616c0_6209, \29752 );
not \U$21371 ( \29754 , RIe1616c0_6209);
or \U$21372 ( \29755 , \29754 , \28843 );
not \U$21373 ( \29756 , \28675 );
and \U$21374 ( \29757 , \28608 , \29756 );
not \U$21375 ( \29758 , \29757 );
not \U$21376 ( \29759 , \28606 );
not \U$21377 ( \29760 , \28738 );
or \U$21378 ( \29761 , \29759 , \29760 );
nand \U$21379 ( \29762 , \29755 , \29758 , \29761 );
and \U$21380 ( \29763 , \29762 , \29330 );
or \U$21381 ( \29764 , \29753 , \29763 );
and \U$21383 ( \29765 , \29764 , 1'b1 );
or \U$21385 ( \29766 , \29765 , 1'b0 );
buf \U$21386 ( \29767 , \29766 );
_DC r23d98_GF_IsGateDCbyConstraint ( \29768_nR23d98 , \29767 , \21944 );
buf \U$21387 ( \29769 , \29768_nR23d98 );
not \U$21388 ( \29770 , \29571 );
and \U$21389 ( \29771 , RIe164168_6210, \29770 );
not \U$21390 ( \29772 , RIe164168_6210);
or \U$21391 ( \29773 , \29772 , \28694 );
not \U$21392 ( \29774 , \28715 );
and \U$21393 ( \29775 , \28626 , \29774 );
not \U$21394 ( \29776 , \29775 );
not \U$21395 ( \29777 , \28624 );
not \U$21396 ( \29778 , \28680 );
or \U$21397 ( \29779 , \29777 , \29778 );
nand \U$21398 ( \29780 , \29773 , \29776 , \29779 );
and \U$21399 ( \29781 , \29780 , \29571 );
or \U$21400 ( \29782 , \29771 , \29781 );
and \U$21402 ( \29783 , \29782 , 1'b1 );
or \U$21404 ( \29784 , \29783 , 1'b0 );
buf \U$21405 ( \29785 , \29784 );
_DC r23d9a_GF_IsGateDCbyConstraint ( \29786_nR23d9a , \29785 , \21944 );
buf \U$21406 ( \29787 , \29786_nR23d9a );
not \U$21407 ( \29788 , \29294 );
and \U$21408 ( \29789 , RIe166c10_6211, \29788 );
not \U$21409 ( \29790 , RIe166c10_6211);
not \U$21410 ( \29791 , \27380 );
nor \U$21411 ( \29792 , \27383 , \29791 );
and \U$21412 ( \29793 , \29792 , \27385 );
not \U$21413 ( \29794 , \27372 );
or \U$21414 ( \29795 , \27370 , \29794 );
not \U$21415 ( \29796 , \29795 );
nand \U$21416 ( \29797 , \27362 , \29796 );
not \U$21417 ( \29798 , \29797 );
or \U$21418 ( \29799 , \29793 , \29798 );
not \U$21419 ( \29800 , \29799 );
not \U$21420 ( \29801 , \29800 );
or \U$21421 ( \29802 , \29790 , \29801 );
not \U$21422 ( \29803 , \29793 );
not \U$21423 ( \29804 , \29803 );
and \U$21424 ( \29805 , \27395 , \29804 );
not \U$21425 ( \29806 , \29805 );
not \U$21426 ( \29807 , \29797 );
buf \U$21427 ( \29808 , \29807 );
not \U$21428 ( \29809 , \29808 );
or \U$21429 ( \29810 , \28657 , \29809 );
nand \U$21430 ( \29811 , \29802 , \29806 , \29810 );
and \U$21431 ( \29812 , \29811 , \29294 );
or \U$21432 ( \29813 , \29789 , \29812 );
and \U$21434 ( \29814 , \29813 , 1'b1 );
or \U$21436 ( \29815 , \29814 , 1'b0 );
buf \U$21437 ( \29816 , \29815 );
_DC r23da4_GF_IsGateDCbyConstraint ( \29817_nR23da4 , \29816 , \21944 );
buf \U$21438 ( \29818 , \29817_nR23da4 );
not \U$21439 ( \29819 , \29571 );
and \U$21440 ( \29820 , RIe39a100_6212, \29819 );
not \U$21441 ( \29821 , RIe39a100_6212);
not \U$21442 ( \29822 , \29800 );
or \U$21443 ( \29823 , \29821 , \29822 );
not \U$21444 ( \29824 , \29793 );
not \U$21445 ( \29825 , \29824 );
and \U$21446 ( \29826 , \27427 , \29825 );
not \U$21447 ( \29827 , \29826 );
buf \U$21448 ( \29828 , \29807 );
not \U$21449 ( \29829 , \29828 );
or \U$21450 ( \29830 , \28679 , \29829 );
nand \U$21451 ( \29831 , \29823 , \29827 , \29830 );
and \U$21452 ( \29832 , \29831 , \29571 );
or \U$21453 ( \29833 , \29820 , \29832 );
and \U$21455 ( \29834 , \29833 , 1'b1 );
or \U$21457 ( \29835 , \29834 , 1'b0 );
buf \U$21458 ( \29836 , \29835 );
_DC r23dba_GF_IsGateDCbyConstraint ( \29837_nR23dba , \29836 , \21944 );
buf \U$21459 ( \29838 , \29837_nR23dba );
not \U$21460 ( \29839 , \29330 );
and \U$21461 ( \29840 , RIe3984e0_6213, \29839 );
not \U$21462 ( \29841 , RIe3984e0_6213);
not \U$21463 ( \29842 , \29800 );
or \U$21464 ( \29843 , \29841 , \29842 );
not \U$21465 ( \29844 , \29824 );
and \U$21466 ( \29845 , \27446 , \29844 );
not \U$21467 ( \29846 , \29845 );
not \U$21468 ( \29847 , \29808 );
or \U$21469 ( \29848 , \28699 , \29847 );
nand \U$21470 ( \29849 , \29843 , \29846 , \29848 );
and \U$21471 ( \29850 , \29849 , \29330 );
or \U$21472 ( \29851 , \29840 , \29850 );
and \U$21474 ( \29852 , \29851 , 1'b1 );
or \U$21476 ( \29853 , \29852 , 1'b0 );
buf \U$21477 ( \29854 , \29853 );
_DC r23dd0_GF_IsGateDCbyConstraint ( \29855_nR23dd0 , \29854 , \21944 );
buf \U$21478 ( \29856 , \29855_nR23dd0 );
not \U$21479 ( \29857 , \29294 );
and \U$21480 ( \29858 , RIe3967d0_6214, \29857 );
not \U$21481 ( \29859 , RIe3967d0_6214);
not \U$21482 ( \29860 , \29800 );
or \U$21483 ( \29861 , \29859 , \29860 );
not \U$21484 ( \29862 , \29824 );
and \U$21485 ( \29863 , \27467 , \29862 );
not \U$21486 ( \29864 , \29863 );
not \U$21487 ( \29865 , \29808 );
or \U$21488 ( \29866 , \28719 , \29865 );
nand \U$21489 ( \29867 , \29861 , \29864 , \29866 );
and \U$21490 ( \29868 , \29867 , \29294 );
or \U$21491 ( \29869 , \29858 , \29868 );
and \U$21493 ( \29870 , \29869 , 1'b1 );
or \U$21495 ( \29871 , \29870 , 1'b0 );
buf \U$21496 ( \29872 , \29871 );
_DC r23de6_GF_IsGateDCbyConstraint ( \29873_nR23de6 , \29872 , \21944 );
buf \U$21497 ( \29874 , \29873_nR23de6 );
not \U$21498 ( \29875 , \29571 );
and \U$21499 ( \29876 , RIe3941d8_6215, \29875 );
not \U$21500 ( \29877 , RIe3941d8_6215);
or \U$21501 ( \29878 , \29877 , \29860 );
not \U$21502 ( \29879 , \29824 );
and \U$21503 ( \29880 , \27486 , \29879 );
not \U$21504 ( \29881 , \29880 );
buf \U$21505 ( \29882 , \29807 );
not \U$21506 ( \29883 , \29882 );
or \U$21507 ( \29884 , \28737 , \29883 );
nand \U$21508 ( \29885 , \29878 , \29881 , \29884 );
and \U$21509 ( \29886 , \29885 , \29571 );
or \U$21510 ( \29887 , \29876 , \29886 );
and \U$21512 ( \29888 , \29887 , 1'b1 );
or \U$21514 ( \29889 , \29888 , 1'b0 );
buf \U$21515 ( \29890 , \29889 );
_DC r23dfc_GF_IsGateDCbyConstraint ( \29891_nR23dfc , \29890 , \21944 );
buf \U$21516 ( \29892 , \29891_nR23dfc );
not \U$21517 ( \29893 , \29330 );
and \U$21518 ( \29894 , RIe391c58_6216, \29893 );
not \U$21519 ( \29895 , RIe391c58_6216);
or \U$21520 ( \29896 , \29895 , \29860 );
not \U$21521 ( \29897 , \29793 );
not \U$21522 ( \29898 , \29897 );
and \U$21523 ( \29899 , \27507 , \29898 );
not \U$21524 ( \29900 , \29899 );
buf \U$21525 ( \29901 , \29807 );
not \U$21526 ( \29902 , \29901 );
or \U$21527 ( \29903 , \28758 , \29902 );
nand \U$21528 ( \29904 , \29896 , \29900 , \29903 );
and \U$21529 ( \29905 , \29904 , \29330 );
or \U$21530 ( \29906 , \29894 , \29905 );
and \U$21532 ( \29907 , \29906 , 1'b1 );
or \U$21534 ( \29908 , \29907 , 1'b0 );
buf \U$21535 ( \29909 , \29908 );
_DC r23e12_GF_IsGateDCbyConstraint ( \29910_nR23e12 , \29909 , \21944 );
buf \U$21536 ( \29911 , \29910_nR23e12 );
not \U$21537 ( \29912 , \29294 );
and \U$21538 ( \29913 , RIe38f5e8_6217, \29912 );
not \U$21539 ( \29914 , RIe38f5e8_6217);
or \U$21540 ( \29915 , \29914 , \29822 );
not \U$21541 ( \29916 , \29793 );
not \U$21542 ( \29917 , \29916 );
and \U$21543 ( \29918 , \27527 , \29917 );
not \U$21544 ( \29919 , \29918 );
not \U$21545 ( \29920 , \29882 );
or \U$21546 ( \29921 , \28777 , \29920 );
nand \U$21547 ( \29922 , \29915 , \29919 , \29921 );
and \U$21548 ( \29923 , \29922 , \29294 );
or \U$21549 ( \29924 , \29913 , \29923 );
and \U$21551 ( \29925 , \29924 , 1'b1 );
or \U$21553 ( \29926 , \29925 , 1'b0 );
buf \U$21554 ( \29927 , \29926 );
_DC r23e1c_GF_IsGateDCbyConstraint ( \29928_nR23e1c , \29927 , \21944 );
buf \U$21555 ( \29929 , \29928_nR23e1c );
not \U$21556 ( \29930 , \29571 );
and \U$21557 ( \29931 , RIe38d428_6218, \29930 );
not \U$21558 ( \29932 , RIe38d428_6218);
or \U$21559 ( \29933 , \29932 , \29860 );
not \U$21560 ( \29934 , \29824 );
and \U$21561 ( \29935 , \27546 , \29934 );
not \U$21562 ( \29936 , \29935 );
not \U$21563 ( \29937 , \29901 );
or \U$21564 ( \29938 , \28795 , \29937 );
nand \U$21565 ( \29939 , \29933 , \29936 , \29938 );
and \U$21566 ( \29940 , \29939 , \29571 );
or \U$21567 ( \29941 , \29931 , \29940 );
and \U$21569 ( \29942 , \29941 , 1'b1 );
or \U$21571 ( \29943 , \29942 , 1'b0 );
buf \U$21572 ( \29944 , \29943 );
_DC r23e1e_GF_IsGateDCbyConstraint ( \29945_nR23e1e , \29944 , \21944 );
buf \U$21573 ( \29946 , \29945_nR23e1e );
not \U$21574 ( \29947 , \29330 );
and \U$21575 ( \29948 , RIe38ae30_6219, \29947 );
not \U$21576 ( \29949 , RIe38ae30_6219);
or \U$21577 ( \29950 , \29949 , \29801 );
not \U$21578 ( \29951 , \29897 );
and \U$21579 ( \29952 , \27568 , \29951 );
not \U$21580 ( \29953 , \29952 );
not \U$21581 ( \29954 , \29882 );
or \U$21582 ( \29955 , \28813 , \29954 );
nand \U$21583 ( \29956 , \29950 , \29953 , \29955 );
and \U$21584 ( \29957 , \29956 , \29330 );
or \U$21585 ( \29958 , \29948 , \29957 );
and \U$21587 ( \29959 , \29958 , 1'b1 );
or \U$21589 ( \29960 , \29959 , 1'b0 );
buf \U$21590 ( \29961 , \29960 );
_DC r23e20_GF_IsGateDCbyConstraint ( \29962_nR23e20 , \29961 , \21944 );
buf \U$21591 ( \29963 , \29962_nR23e20 );
buf \U$21592 ( \29964 , \28249 );
not \U$21593 ( \29965 , \29964 );
and \U$21594 ( \29966 , RIe389030_6220, \29965 );
not \U$21595 ( \29967 , RIe389030_6220);
or \U$21596 ( \29968 , \29967 , \29801 );
not \U$21597 ( \29969 , \29803 );
and \U$21598 ( \29970 , \27588 , \29969 );
not \U$21599 ( \29971 , \29970 );
not \U$21600 ( \29972 , \27585 );
not \U$21601 ( \29973 , \29882 );
or \U$21602 ( \29974 , \29972 , \29973 );
nand \U$21603 ( \29975 , \29968 , \29971 , \29974 );
and \U$21604 ( \29976 , \29975 , \29964 );
or \U$21605 ( \29977 , \29966 , \29976 );
and \U$21607 ( \29978 , \29977 , 1'b1 );
or \U$21609 ( \29979 , \29978 , 1'b0 );
buf \U$21610 ( \29980 , \29979 );
_DC r23e22_GF_IsGateDCbyConstraint ( \29981_nR23e22 , \29980 , \21944 );
buf \U$21611 ( \29982 , \29981_nR23e22 );
not \U$21612 ( \29983 , \29571 );
and \U$21613 ( \29984 , RIe386fd8_6221, \29983 );
not \U$21614 ( \29985 , RIe386fd8_6221);
not \U$21615 ( \29986 , \29800 );
or \U$21616 ( \29987 , \29985 , \29986 );
not \U$21617 ( \29988 , \29916 );
and \U$21618 ( \29989 , \27609 , \29988 );
not \U$21619 ( \29990 , \29989 );
nand \U$21620 ( \29991 , \27606 , \29882 );
nand \U$21621 ( \29992 , \29987 , \29990 , \29991 );
and \U$21622 ( \29993 , \29992 , \29571 );
or \U$21623 ( \29994 , \29984 , \29993 );
and \U$21625 ( \29995 , \29994 , 1'b1 );
or \U$21627 ( \29996 , \29995 , 1'b0 );
buf \U$21628 ( \29997 , \29996 );
_DC r23da6_GF_IsGateDCbyConstraint ( \29998_nR23da6 , \29997 , \21944 );
buf \U$21629 ( \29999 , \29998_nR23da6 );
buf \U$21630 ( \30000 , \29329 );
not \U$21631 ( \30001 , \30000 );
and \U$21632 ( \30002 , RIe384ff8_6222, \30001 );
not \U$21633 ( \30003 , RIe384ff8_6222);
or \U$21634 ( \30004 , \30003 , \29822 );
not \U$21635 ( \30005 , \29824 );
and \U$21636 ( \30006 , \27628 , \30005 );
not \U$21637 ( \30007 , \30006 );
nand \U$21638 ( \30008 , \27625 , \29808 );
nand \U$21639 ( \30009 , \30004 , \30007 , \30008 );
and \U$21640 ( \30010 , \30009 , \30000 );
or \U$21641 ( \30011 , \30002 , \30010 );
and \U$21643 ( \30012 , \30011 , 1'b1 );
or \U$21645 ( \30013 , \30012 , 1'b0 );
buf \U$21646 ( \30014 , \30013 );
_DC r23da8_GF_IsGateDCbyConstraint ( \30015_nR23da8 , \30014 , \21944 );
buf \U$21647 ( \30016 , \30015_nR23da8 );
not \U$21648 ( \30017 , \29964 );
and \U$21649 ( \30018 , RIe3832e8_6223, \30017 );
not \U$21650 ( \30019 , RIe3832e8_6223);
or \U$21651 ( \30020 , \30019 , \29822 );
not \U$21652 ( \30021 , \29803 );
and \U$21653 ( \30022 , \27648 , \30021 );
not \U$21654 ( \30023 , \30022 );
nand \U$21655 ( \30024 , \27645 , \29901 );
nand \U$21656 ( \30025 , \30020 , \30023 , \30024 );
and \U$21657 ( \30026 , \30025 , \29964 );
or \U$21658 ( \30027 , \30018 , \30026 );
and \U$21660 ( \30028 , \30027 , 1'b1 );
or \U$21662 ( \30029 , \30028 , 1'b0 );
buf \U$21663 ( \30030 , \30029 );
_DC r23daa_GF_IsGateDCbyConstraint ( \30031_nR23daa , \30030 , \21944 );
buf \U$21664 ( \30032 , \30031_nR23daa );
not \U$21665 ( \30033 , \29571 );
and \U$21666 ( \30034 , RIe381218_6224, \30033 );
not \U$21667 ( \30035 , RIe381218_6224);
or \U$21668 ( \30036 , \30035 , \29822 );
not \U$21669 ( \30037 , \29916 );
and \U$21670 ( \30038 , \27668 , \30037 );
not \U$21671 ( \30039 , \30038 );
nand \U$21672 ( \30040 , \27665 , \29808 );
nand \U$21673 ( \30041 , \30036 , \30039 , \30040 );
and \U$21674 ( \30042 , \30041 , \29571 );
or \U$21675 ( \30043 , \30034 , \30042 );
and \U$21677 ( \30044 , \30043 , 1'b1 );
or \U$21679 ( \30045 , \30044 , 1'b0 );
buf \U$21680 ( \30046 , \30045 );
_DC r23dac_GF_IsGateDCbyConstraint ( \30047_nR23dac , \30046 , \21944 );
buf \U$21681 ( \30048 , \30047_nR23dac );
not \U$21682 ( \30049 , \30000 );
and \U$21683 ( \30050 , RIe37f148_6225, \30049 );
not \U$21684 ( \30051 , RIe37f148_6225);
or \U$21685 ( \30052 , \30051 , \29801 );
not \U$21686 ( \30053 , \29916 );
and \U$21687 ( \30054 , \27686 , \30053 );
not \U$21688 ( \30055 , \30054 );
nand \U$21689 ( \30056 , \27684 , \29808 );
nand \U$21690 ( \30057 , \30052 , \30055 , \30056 );
and \U$21691 ( \30058 , \30057 , \30000 );
or \U$21692 ( \30059 , \30050 , \30058 );
and \U$21694 ( \30060 , \30059 , 1'b1 );
or \U$21696 ( \30061 , \30060 , 1'b0 );
buf \U$21697 ( \30062 , \30061 );
_DC r23dae_GF_IsGateDCbyConstraint ( \30063_nR23dae , \30062 , \21944 );
buf \U$21698 ( \30064 , \30063_nR23dae );
not \U$21699 ( \30065 , \29964 );
and \U$21700 ( \30066 , RIe37ce20_6226, \30065 );
not \U$21701 ( \30067 , RIe37ce20_6226);
or \U$21702 ( \30068 , \30067 , \29801 );
not \U$21703 ( \30069 , \29897 );
and \U$21704 ( \30070 , \27704 , \30069 );
not \U$21705 ( \30071 , \30070 );
nand \U$21706 ( \30072 , \27702 , \29828 );
nand \U$21707 ( \30073 , \30068 , \30071 , \30072 );
and \U$21708 ( \30074 , \30073 , \29964 );
or \U$21709 ( \30075 , \30066 , \30074 );
and \U$21711 ( \30076 , \30075 , 1'b1 );
or \U$21713 ( \30077 , \30076 , 1'b0 );
buf \U$21714 ( \30078 , \30077 );
_DC r23db0_GF_IsGateDCbyConstraint ( \30079_nR23db0 , \30078 , \21944 );
buf \U$21715 ( \30080 , \30079_nR23db0 );
not \U$21716 ( \30081 , \29571 );
and \U$21717 ( \30082 , RIe37aeb8_6227, \30081 );
not \U$21718 ( \30083 , RIe37aeb8_6227);
or \U$21719 ( \30084 , \30083 , \29986 );
not \U$21720 ( \30085 , \29916 );
and \U$21721 ( \30086 , \27722 , \30085 );
not \U$21722 ( \30087 , \30086 );
nand \U$21723 ( \30088 , \27720 , \29828 );
nand \U$21724 ( \30089 , \30084 , \30087 , \30088 );
and \U$21725 ( \30090 , \30089 , \29571 );
or \U$21726 ( \30091 , \30082 , \30090 );
and \U$21728 ( \30092 , \30091 , 1'b1 );
or \U$21730 ( \30093 , \30092 , 1'b0 );
buf \U$21731 ( \30094 , \30093 );
_DC r23db2_GF_IsGateDCbyConstraint ( \30095_nR23db2 , \30094 , \21944 );
buf \U$21732 ( \30096 , \30095_nR23db2 );
not \U$21733 ( \30097 , \30000 );
and \U$21734 ( \30098 , RIe378668_6228, \30097 );
not \U$21735 ( \30099 , RIe378668_6228);
or \U$21736 ( \30100 , \30099 , \29822 );
not \U$21737 ( \30101 , \29916 );
and \U$21738 ( \30102 , \27741 , \30101 );
not \U$21739 ( \30103 , \30102 );
nand \U$21740 ( \30104 , \27738 , \29828 );
nand \U$21741 ( \30105 , \30100 , \30103 , \30104 );
and \U$21742 ( \30106 , \30105 , \30000 );
or \U$21743 ( \30107 , \30098 , \30106 );
and \U$21745 ( \30108 , \30107 , 1'b1 );
or \U$21747 ( \30109 , \30108 , 1'b0 );
buf \U$21748 ( \30110 , \30109 );
_DC r23db4_GF_IsGateDCbyConstraint ( \30111_nR23db4 , \30110 , \21944 );
buf \U$21749 ( \30112 , \30111_nR23db4 );
not \U$21750 ( \30113 , \29964 );
and \U$21751 ( \30114 , RIe3755a8_6229, \30113 );
not \U$21752 ( \30115 , RIe3755a8_6229);
or \U$21753 ( \30116 , \30115 , \29842 );
not \U$21754 ( \30117 , \29793 );
not \U$21755 ( \30118 , \30117 );
and \U$21756 ( \30119 , \27760 , \30118 );
not \U$21757 ( \30120 , \30119 );
nand \U$21758 ( \30121 , \27757 , \29901 );
nand \U$21759 ( \30122 , \30116 , \30120 , \30121 );
and \U$21760 ( \30123 , \30122 , \29964 );
or \U$21761 ( \30124 , \30114 , \30123 );
and \U$21763 ( \30125 , \30124 , 1'b1 );
or \U$21765 ( \30126 , \30125 , 1'b0 );
buf \U$21766 ( \30127 , \30126 );
_DC r23db6_GF_IsGateDCbyConstraint ( \30128_nR23db6 , \30127 , \21944 );
buf \U$21767 ( \30129 , \30128_nR23db6 );
not \U$21768 ( \30130 , \29571 );
and \U$21769 ( \30131 , RIe372c68_6230, \30130 );
not \U$21770 ( \30132 , RIe372c68_6230);
or \U$21771 ( \30133 , \30132 , \29860 );
not \U$21772 ( \30134 , \29916 );
and \U$21773 ( \30135 , \27779 , \30134 );
not \U$21774 ( \30136 , \30135 );
nand \U$21775 ( \30137 , \27776 , \29808 );
nand \U$21776 ( \30138 , \30133 , \30136 , \30137 );
and \U$21777 ( \30139 , \30138 , \29571 );
or \U$21778 ( \30140 , \30131 , \30139 );
and \U$21780 ( \30141 , \30140 , 1'b1 );
or \U$21782 ( \30142 , \30141 , 1'b0 );
buf \U$21783 ( \30143 , \30142 );
_DC r23db8_GF_IsGateDCbyConstraint ( \30144_nR23db8 , \30143 , \21944 );
buf \U$21784 ( \30145 , \30144_nR23db8 );
not \U$21785 ( \30146 , \30000 );
and \U$21786 ( \30147 , RIe2703f8_6231, \30146 );
not \U$21787 ( \30148 , RIe2703f8_6231);
or \U$21788 ( \30149 , \30148 , \29801 );
not \U$21789 ( \30150 , \29897 );
and \U$21790 ( \30151 , \27799 , \30150 );
not \U$21791 ( \30152 , \30151 );
not \U$21792 ( \30153 , \29828 );
or \U$21793 ( \30154 , \29013 , \30153 );
nand \U$21794 ( \30155 , \30149 , \30152 , \30154 );
and \U$21795 ( \30156 , \30155 , \30000 );
or \U$21796 ( \30157 , \30147 , \30156 );
and \U$21798 ( \30158 , \30157 , 1'b1 );
or \U$21800 ( \30159 , \30158 , 1'b0 );
buf \U$21801 ( \30160 , \30159 );
_DC r23dbc_GF_IsGateDCbyConstraint ( \30161_nR23dbc , \30160 , \21944 );
buf \U$21802 ( \30162 , \30161_nR23dbc );
not \U$21803 ( \30163 , \29964 );
and \U$21804 ( \30164 , RIe26d4a0_6232, \30163 );
not \U$21805 ( \30165 , RIe26d4a0_6232);
or \U$21806 ( \30166 , \30165 , \29842 );
not \U$21807 ( \30167 , \29803 );
and \U$21808 ( \30168 , \27817 , \30167 );
not \U$21809 ( \30169 , \30168 );
not \U$21810 ( \30170 , \29828 );
or \U$21811 ( \30171 , \29031 , \30170 );
nand \U$21812 ( \30172 , \30166 , \30169 , \30171 );
and \U$21813 ( \30173 , \30172 , \29964 );
or \U$21814 ( \30174 , \30164 , \30173 );
and \U$21816 ( \30175 , \30174 , 1'b1 );
or \U$21818 ( \30176 , \30175 , 1'b0 );
buf \U$21819 ( \30177 , \30176 );
_DC r23dbe_GF_IsGateDCbyConstraint ( \30178_nR23dbe , \30177 , \21944 );
buf \U$21820 ( \30179 , \30178_nR23dbe );
not \U$21821 ( \30180 , \27458 );
and \U$21822 ( \30181 , RIe26aae8_6233, \30180 );
not \U$21823 ( \30182 , RIe26aae8_6233);
or \U$21824 ( \30183 , \30182 , \29986 );
not \U$21825 ( \30184 , \29824 );
and \U$21826 ( \30185 , \27835 , \30184 );
not \U$21827 ( \30186 , \30185 );
not \U$21828 ( \30187 , \29808 );
or \U$21829 ( \30188 , \29049 , \30187 );
nand \U$21830 ( \30189 , \30183 , \30186 , \30188 );
and \U$21831 ( \30190 , \30189 , \27458 );
or \U$21832 ( \30191 , \30181 , \30190 );
and \U$21834 ( \30192 , \30191 , 1'b1 );
or \U$21836 ( \30193 , \30192 , 1'b0 );
buf \U$21837 ( \30194 , \30193 );
_DC r23dc0_GF_IsGateDCbyConstraint ( \30195_nR23dc0 , \30194 , \21944 );
buf \U$21838 ( \30196 , \30195_nR23dc0 );
not \U$21839 ( \30197 , \30000 );
and \U$21840 ( \30198 , RIe2686d0_6234, \30197 );
not \U$21841 ( \30199 , RIe2686d0_6234);
or \U$21842 ( \30200 , \30199 , \29986 );
not \U$21843 ( \30201 , \29897 );
and \U$21844 ( \30202 , \27854 , \30201 );
not \U$21845 ( \30203 , \30202 );
not \U$21846 ( \30204 , \29882 );
or \U$21847 ( \30205 , \29067 , \30204 );
nand \U$21848 ( \30206 , \30200 , \30203 , \30205 );
and \U$21849 ( \30207 , \30206 , \30000 );
or \U$21850 ( \30208 , \30198 , \30207 );
and \U$21852 ( \30209 , \30208 , 1'b1 );
or \U$21854 ( \30210 , \30209 , 1'b0 );
buf \U$21855 ( \30211 , \30210 );
_DC r23dc2_GF_IsGateDCbyConstraint ( \30212_nR23dc2 , \30211 , \21944 );
buf \U$21856 ( \30213 , \30212_nR23dc2 );
not \U$21857 ( \30214 , \29964 );
and \U$21858 ( \30215 , RIe265ca0_6235, \30214 );
not \U$21859 ( \30216 , RIe265ca0_6235);
or \U$21860 ( \30217 , \30216 , \29860 );
not \U$21861 ( \30218 , \29803 );
and \U$21862 ( \30219 , \27873 , \30218 );
not \U$21863 ( \30220 , \30219 );
not \U$21864 ( \30221 , \29828 );
or \U$21865 ( \30222 , \29085 , \30221 );
nand \U$21866 ( \30223 , \30217 , \30220 , \30222 );
and \U$21867 ( \30224 , \30223 , \29964 );
or \U$21868 ( \30225 , \30215 , \30224 );
and \U$21870 ( \30226 , \30225 , 1'b1 );
or \U$21872 ( \30227 , \30226 , 1'b0 );
buf \U$21873 ( \30228 , \30227 );
_DC r23dc4_GF_IsGateDCbyConstraint ( \30229_nR23dc4 , \30228 , \21944 );
buf \U$21874 ( \30230 , \30229_nR23dc4 );
not \U$21875 ( \30231 , \27458 );
and \U$21876 ( \30232 , RIe264170_6236, \30231 );
not \U$21877 ( \30233 , RIe264170_6236);
or \U$21878 ( \30234 , \30233 , \29986 );
not \U$21879 ( \30235 , \30117 );
and \U$21880 ( \30236 , \27892 , \30235 );
not \U$21881 ( \30237 , \30236 );
not \U$21882 ( \30238 , \29882 );
or \U$21883 ( \30239 , \29103 , \30238 );
nand \U$21884 ( \30240 , \30234 , \30237 , \30239 );
and \U$21885 ( \30241 , \30240 , \27458 );
or \U$21886 ( \30242 , \30232 , \30241 );
and \U$21888 ( \30243 , \30242 , 1'b1 );
or \U$21890 ( \30244 , \30243 , 1'b0 );
buf \U$21891 ( \30245 , \30244 );
_DC r23dc6_GF_IsGateDCbyConstraint ( \30246_nR23dc6 , \30245 , \21944 );
buf \U$21892 ( \30247 , \30246_nR23dc6 );
not \U$21893 ( \30248 , \30000 );
and \U$21894 ( \30249 , RIe2616c8_6237, \30248 );
not \U$21895 ( \30250 , RIe2616c8_6237);
or \U$21896 ( \30251 , \30250 , \29842 );
not \U$21897 ( \30252 , \29803 );
and \U$21898 ( \30253 , \27911 , \30252 );
not \U$21899 ( \30254 , \30253 );
not \U$21900 ( \30255 , \29828 );
or \U$21901 ( \30256 , \29121 , \30255 );
nand \U$21902 ( \30257 , \30251 , \30254 , \30256 );
and \U$21903 ( \30258 , \30257 , \30000 );
or \U$21904 ( \30259 , \30249 , \30258 );
and \U$21906 ( \30260 , \30259 , 1'b1 );
or \U$21908 ( \30261 , \30260 , 1'b0 );
buf \U$21909 ( \30262 , \30261 );
_DC r23dc8_GF_IsGateDCbyConstraint ( \30263_nR23dc8 , \30262 , \21944 );
buf \U$21910 ( \30264 , \30263_nR23dc8 );
not \U$21911 ( \30265 , \29964 );
and \U$21912 ( \30266 , RIe25f238_6238, \30265 );
not \U$21913 ( \30267 , RIe25f238_6238);
or \U$21914 ( \30268 , \30267 , \29860 );
not \U$21915 ( \30269 , \29824 );
and \U$21916 ( \30270 , \27930 , \30269 );
not \U$21917 ( \30271 , \30270 );
not \U$21918 ( \30272 , \29828 );
or \U$21919 ( \30273 , \29139 , \30272 );
nand \U$21920 ( \30274 , \30268 , \30271 , \30273 );
and \U$21921 ( \30275 , \30274 , \29964 );
or \U$21922 ( \30276 , \30266 , \30275 );
and \U$21924 ( \30277 , \30276 , 1'b1 );
or \U$21926 ( \30278 , \30277 , 1'b0 );
buf \U$21927 ( \30279 , \30278 );
_DC r23dca_GF_IsGateDCbyConstraint ( \30280_nR23dca , \30279 , \21944 );
buf \U$21928 ( \30281 , \30280_nR23dca );
not \U$21929 ( \30282 , \27363 );
and \U$21930 ( \30283 , RIe25c6a0_6239, \30282 );
not \U$21931 ( \30284 , RIe25c6a0_6239);
or \U$21932 ( \30285 , \30284 , \29842 );
not \U$21933 ( \30286 , \30117 );
and \U$21934 ( \30287 , \27949 , \30286 );
not \U$21935 ( \30288 , \30287 );
not \U$21936 ( \30289 , \29808 );
or \U$21937 ( \30290 , \29157 , \30289 );
nand \U$21938 ( \30291 , \30285 , \30288 , \30290 );
and \U$21939 ( \30292 , \30291 , \27363 );
or \U$21940 ( \30293 , \30283 , \30292 );
and \U$21942 ( \30294 , \30293 , 1'b1 );
or \U$21944 ( \30295 , \30294 , 1'b0 );
buf \U$21945 ( \30296 , \30295 );
_DC r23dcc_GF_IsGateDCbyConstraint ( \30297_nR23dcc , \30296 , \21944 );
buf \U$21946 ( \30298 , \30297_nR23dcc );
not \U$21947 ( \30299 , \30000 );
and \U$21948 ( \30300 , RIe259ec8_6240, \30299 );
not \U$21949 ( \30301 , RIe259ec8_6240);
or \U$21950 ( \30302 , \30301 , \29860 );
not \U$21951 ( \30303 , \29897 );
and \U$21952 ( \30304 , \27968 , \30303 );
not \U$21953 ( \30305 , \30304 );
not \U$21954 ( \30306 , \29808 );
or \U$21955 ( \30307 , \29175 , \30306 );
nand \U$21956 ( \30308 , \30302 , \30305 , \30307 );
and \U$21957 ( \30309 , \30308 , \30000 );
or \U$21958 ( \30310 , \30300 , \30309 );
and \U$21960 ( \30311 , \30310 , 1'b1 );
or \U$21962 ( \30312 , \30311 , 1'b0 );
buf \U$21963 ( \30313 , \30312 );
_DC r23dce_GF_IsGateDCbyConstraint ( \30314_nR23dce , \30313 , \21944 );
buf \U$21964 ( \30315 , \30314_nR23dce );
not \U$21965 ( \30316 , \29964 );
and \U$21966 ( \30317 , RIe257240_6241, \30316 );
not \U$21967 ( \30318 , RIe257240_6241);
or \U$21968 ( \30319 , \30318 , \29986 );
not \U$21969 ( \30320 , \29803 );
and \U$21970 ( \30321 , \27988 , \30320 );
not \U$21971 ( \30322 , \30321 );
not \U$21972 ( \30323 , \29828 );
or \U$21973 ( \30324 , \29193 , \30323 );
nand \U$21974 ( \30325 , \30319 , \30322 , \30324 );
and \U$21975 ( \30326 , \30325 , \29964 );
or \U$21976 ( \30327 , \30317 , \30326 );
and \U$21978 ( \30328 , \30327 , 1'b1 );
or \U$21980 ( \30329 , \30328 , 1'b0 );
buf \U$21981 ( \30330 , \30329 );
_DC r23dd2_GF_IsGateDCbyConstraint ( \30331_nR23dd2 , \30330 , \21944 );
buf \U$21982 ( \30332 , \30331_nR23dd2 );
not \U$21983 ( \30333 , \27363 );
and \U$21984 ( \30334 , RIe254018_6242, \30333 );
not \U$21985 ( \30335 , RIe254018_6242);
or \U$21986 ( \30336 , \30335 , \29822 );
not \U$21987 ( \30337 , \29897 );
and \U$21988 ( \30338 , \28009 , \30337 );
not \U$21989 ( \30339 , \30338 );
not \U$21990 ( \30340 , \29828 );
or \U$21991 ( \30341 , \29211 , \30340 );
nand \U$21992 ( \30342 , \30336 , \30339 , \30341 );
and \U$21993 ( \30343 , \30342 , \27363 );
or \U$21994 ( \30344 , \30334 , \30343 );
and \U$21996 ( \30345 , \30344 , 1'b1 );
or \U$21998 ( \30346 , \30345 , 1'b0 );
buf \U$21999 ( \30347 , \30346 );
_DC r23dd4_GF_IsGateDCbyConstraint ( \30348_nR23dd4 , \30347 , \21944 );
buf \U$22000 ( \30349 , \30348_nR23dd4 );
not \U$22001 ( \30350 , \30000 );
and \U$22002 ( \30351 , RIe251408_6243, \30350 );
not \U$22003 ( \30352 , RIe251408_6243);
or \U$22004 ( \30353 , \30352 , \29822 );
not \U$22005 ( \30354 , \29897 );
and \U$22006 ( \30355 , \28029 , \30354 );
not \U$22007 ( \30356 , \30355 );
not \U$22008 ( \30357 , \29808 );
or \U$22009 ( \30358 , \29229 , \30357 );
nand \U$22010 ( \30359 , \30353 , \30356 , \30358 );
and \U$22011 ( \30360 , \30359 , \30000 );
or \U$22012 ( \30361 , \30351 , \30360 );
and \U$22014 ( \30362 , \30361 , 1'b1 );
or \U$22016 ( \30363 , \30362 , 1'b0 );
buf \U$22017 ( \30364 , \30363 );
_DC r23dd6_GF_IsGateDCbyConstraint ( \30365_nR23dd6 , \30364 , \21944 );
buf \U$22018 ( \30366 , \30365_nR23dd6 );
not \U$22019 ( \30367 , \29964 );
and \U$22020 ( \30368 , RIe24e8e8_6244, \30367 );
not \U$22021 ( \30369 , RIe24e8e8_6244);
or \U$22022 ( \30370 , \30369 , \29842 );
not \U$22023 ( \30371 , \29916 );
and \U$22024 ( \30372 , \28048 , \30371 );
not \U$22025 ( \30373 , \30372 );
not \U$22026 ( \30374 , \29828 );
or \U$22027 ( \30375 , \29247 , \30374 );
nand \U$22028 ( \30376 , \30370 , \30373 , \30375 );
and \U$22029 ( \30377 , \30376 , \29964 );
or \U$22030 ( \30378 , \30368 , \30377 );
and \U$22032 ( \30379 , \30378 , 1'b1 );
or \U$22034 ( \30380 , \30379 , 1'b0 );
buf \U$22035 ( \30381 , \30380 );
_DC r23dd8_GF_IsGateDCbyConstraint ( \30382_nR23dd8 , \30381 , \21944 );
buf \U$22036 ( \30383 , \30382_nR23dd8 );
not \U$22037 ( \30384 , \27363 );
and \U$22038 ( \30385 , RIe24c110_6245, \30384 );
not \U$22039 ( \30386 , RIe24c110_6245);
or \U$22040 ( \30387 , \30386 , \29801 );
not \U$22041 ( \30388 , \29916 );
and \U$22042 ( \30389 , \28066 , \30388 );
not \U$22043 ( \30390 , \30389 );
not \U$22044 ( \30391 , \29808 );
or \U$22045 ( \30392 , \29265 , \30391 );
nand \U$22046 ( \30393 , \30387 , \30390 , \30392 );
and \U$22047 ( \30394 , \30393 , \27363 );
or \U$22048 ( \30395 , \30385 , \30394 );
and \U$22050 ( \30396 , \30395 , 1'b1 );
or \U$22052 ( \30397 , \30396 , 1'b0 );
buf \U$22053 ( \30398 , \30397 );
_DC r23dda_GF_IsGateDCbyConstraint ( \30399_nR23dda , \30398 , \21944 );
buf \U$22054 ( \30400 , \30399_nR23dda );
not \U$22055 ( \30401 , \30000 );
and \U$22056 ( \30402 , RIe248d08_6246, \30401 );
not \U$22057 ( \30403 , RIe248d08_6246);
or \U$22058 ( \30404 , \30403 , \29842 );
not \U$22059 ( \30405 , \29916 );
and \U$22060 ( \30406 , \28085 , \30405 );
not \U$22061 ( \30407 , \30406 );
nand \U$22062 ( \30408 , \28082 , \29828 );
nand \U$22063 ( \30409 , \30404 , \30407 , \30408 );
and \U$22064 ( \30410 , \30409 , \30000 );
or \U$22065 ( \30411 , \30402 , \30410 );
and \U$22067 ( \30412 , \30411 , 1'b1 );
or \U$22069 ( \30413 , \30412 , 1'b0 );
buf \U$22070 ( \30414 , \30413 );
_DC r23ddc_GF_IsGateDCbyConstraint ( \30415_nR23ddc , \30414 , \21944 );
buf \U$22071 ( \30416 , \30415_nR23ddc );
not \U$22072 ( \30417 , \29964 );
and \U$22073 ( \30418 , RIe246170_6247, \30417 );
not \U$22074 ( \30419 , RIe246170_6247);
or \U$22075 ( \30420 , \30419 , \29860 );
not \U$22076 ( \30421 , \29916 );
and \U$22077 ( \30422 , \28104 , \30421 );
not \U$22078 ( \30423 , \30422 );
nand \U$22079 ( \30424 , \28101 , \29828 );
nand \U$22080 ( \30425 , \30420 , \30423 , \30424 );
and \U$22081 ( \30426 , \30425 , \29964 );
or \U$22082 ( \30427 , \30418 , \30426 );
and \U$22084 ( \30428 , \30427 , 1'b1 );
or \U$22086 ( \30429 , \30428 , 1'b0 );
buf \U$22087 ( \30430 , \30429 );
_DC r23dde_GF_IsGateDCbyConstraint ( \30431_nR23dde , \30430 , \21944 );
buf \U$22088 ( \30432 , \30431_nR23dde );
not \U$22089 ( \30433 , \27363 );
and \U$22090 ( \30434 , RIe2435d8_6248, \30433 );
not \U$22091 ( \30435 , RIe2435d8_6248);
or \U$22092 ( \30436 , \30435 , \29842 );
not \U$22093 ( \30437 , \29897 );
and \U$22094 ( \30438 , \28123 , \30437 );
not \U$22095 ( \30439 , \30438 );
nand \U$22096 ( \30440 , \28120 , \29828 );
nand \U$22097 ( \30441 , \30436 , \30439 , \30440 );
and \U$22098 ( \30442 , \30441 , \27363 );
or \U$22099 ( \30443 , \30434 , \30442 );
and \U$22101 ( \30444 , \30443 , 1'b1 );
or \U$22103 ( \30445 , \30444 , 1'b0 );
buf \U$22104 ( \30446 , \30445 );
_DC r23de0_GF_IsGateDCbyConstraint ( \30447_nR23de0 , \30446 , \21944 );
buf \U$22105 ( \30448 , \30447_nR23de0 );
not \U$22106 ( \30449 , \30000 );
and \U$22107 ( \30450 , RIe2418c8_6249, \30449 );
not \U$22108 ( \30451 , RIe2418c8_6249);
or \U$22109 ( \30452 , \30451 , \29822 );
not \U$22110 ( \30453 , \29824 );
and \U$22111 ( \30454 , \28142 , \30453 );
not \U$22112 ( \30455 , \30454 );
nand \U$22113 ( \30456 , \28139 , \29901 );
nand \U$22114 ( \30457 , \30452 , \30455 , \30456 );
and \U$22115 ( \30458 , \30457 , \30000 );
or \U$22116 ( \30459 , \30450 , \30458 );
and \U$22118 ( \30460 , \30459 , 1'b1 );
or \U$22120 ( \30461 , \30460 , 1'b0 );
buf \U$22121 ( \30462 , \30461 );
_DC r23de2_GF_IsGateDCbyConstraint ( \30463_nR23de2 , \30462 , \21944 );
buf \U$22122 ( \30464 , \30463_nR23de2 );
not \U$22123 ( \30465 , \29964 );
and \U$22124 ( \30466 , RIe23fb40_6250, \30465 );
not \U$22125 ( \30467 , RIe23fb40_6250);
or \U$22126 ( \30468 , \30467 , \29986 );
not \U$22127 ( \30469 , \29916 );
and \U$22128 ( \30470 , \28161 , \30469 );
not \U$22129 ( \30471 , \30470 );
nand \U$22130 ( \30472 , \28158 , \29882 );
nand \U$22131 ( \30473 , \30468 , \30471 , \30472 );
and \U$22132 ( \30474 , \30473 , \29964 );
or \U$22133 ( \30475 , \30466 , \30474 );
and \U$22135 ( \30476 , \30475 , 1'b1 );
or \U$22137 ( \30477 , \30476 , 1'b0 );
buf \U$22138 ( \30478 , \30477 );
_DC r23de4_GF_IsGateDCbyConstraint ( \30479_nR23de4 , \30478 , \21944 );
buf \U$22139 ( \30480 , \30479_nR23de4 );
not \U$22140 ( \30481 , \27363 );
and \U$22141 ( \30482 , RIe23dcc8_6251, \30481 );
not \U$22142 ( \30483 , RIe23dcc8_6251);
or \U$22143 ( \30484 , \30483 , \29986 );
not \U$22144 ( \30485 , \29824 );
and \U$22145 ( \30486 , \28180 , \30485 );
not \U$22146 ( \30487 , \30486 );
nand \U$22147 ( \30488 , \28177 , \29808 );
nand \U$22148 ( \30489 , \30484 , \30487 , \30488 );
and \U$22149 ( \30490 , \30489 , \27363 );
or \U$22150 ( \30491 , \30482 , \30490 );
and \U$22152 ( \30492 , \30491 , 1'b1 );
or \U$22154 ( \30493 , \30492 , 1'b0 );
buf \U$22155 ( \30494 , \30493 );
_DC r23de8_GF_IsGateDCbyConstraint ( \30495_nR23de8 , \30494 , \21944 );
buf \U$22156 ( \30496 , \30495_nR23de8 );
not \U$22157 ( \30497 , \30000 );
and \U$22158 ( \30498 , RIe23ba18_6252, \30497 );
not \U$22159 ( \30499 , RIe23ba18_6252);
or \U$22160 ( \30500 , \30499 , \29801 );
not \U$22161 ( \30501 , \29897 );
and \U$22162 ( \30502 , \28199 , \30501 );
not \U$22163 ( \30503 , \30502 );
nand \U$22164 ( \30504 , \28196 , \29808 );
nand \U$22165 ( \30505 , \30500 , \30503 , \30504 );
and \U$22166 ( \30506 , \30505 , \30000 );
or \U$22167 ( \30507 , \30498 , \30506 );
and \U$22169 ( \30508 , \30507 , 1'b1 );
or \U$22171 ( \30509 , \30508 , 1'b0 );
buf \U$22172 ( \30510 , \30509 );
_DC r23dea_GF_IsGateDCbyConstraint ( \30511_nR23dea , \30510 , \21944 );
buf \U$22173 ( \30512 , \30511_nR23dea );
not \U$22174 ( \30513 , \29964 );
and \U$22175 ( \30514 , RIe239948_6253, \30513 );
not \U$22176 ( \30515 , RIe239948_6253);
or \U$22177 ( \30516 , \30515 , \29822 );
not \U$22178 ( \30517 , \29803 );
and \U$22179 ( \30518 , \28218 , \30517 );
not \U$22180 ( \30519 , \30518 );
not \U$22181 ( \30520 , \28215 );
not \U$22182 ( \30521 , \29901 );
or \U$22183 ( \30522 , \30520 , \30521 );
nand \U$22184 ( \30523 , \30516 , \30519 , \30522 );
and \U$22185 ( \30524 , \30523 , \29964 );
or \U$22186 ( \30525 , \30514 , \30524 );
and \U$22188 ( \30526 , \30525 , 1'b1 );
or \U$22190 ( \30527 , \30526 , 1'b0 );
buf \U$22191 ( \30528 , \30527 );
_DC r23dec_GF_IsGateDCbyConstraint ( \30529_nR23dec , \30528 , \21944 );
buf \U$22192 ( \30530 , \30529_nR23dec );
not \U$22193 ( \30531 , \27363 );
and \U$22194 ( \30532 , RIe2381d8_6254, \30531 );
not \U$22195 ( \30533 , RIe2381d8_6254);
or \U$22196 ( \30534 , \30533 , \29822 );
not \U$22197 ( \30535 , \30117 );
and \U$22198 ( \30536 , \28237 , \30535 );
not \U$22199 ( \30537 , \30536 );
not \U$22200 ( \30538 , \28235 );
not \U$22201 ( \30539 , \29808 );
or \U$22202 ( \30540 , \30538 , \30539 );
nand \U$22203 ( \30541 , \30534 , \30537 , \30540 );
and \U$22204 ( \30542 , \30541 , \27363 );
or \U$22205 ( \30543 , \30532 , \30542 );
and \U$22207 ( \30544 , \30543 , 1'b1 );
or \U$22209 ( \30545 , \30544 , 1'b0 );
buf \U$22210 ( \30546 , \30545 );
_DC r23dee_GF_IsGateDCbyConstraint ( \30547_nR23dee , \30546 , \21944 );
buf \U$22211 ( \30548 , \30547_nR23dee );
not \U$22212 ( \30549 , \30000 );
and \U$22213 ( \30550 , RIe236720_6255, \30549 );
not \U$22214 ( \30551 , RIe236720_6255);
or \U$22215 ( \30552 , \30551 , \29860 );
not \U$22216 ( \30553 , \29803 );
and \U$22217 ( \30554 , \28257 , \30553 );
not \U$22218 ( \30555 , \30554 );
not \U$22219 ( \30556 , \29828 );
or \U$22220 ( \30557 , \29434 , \30556 );
nand \U$22221 ( \30558 , \30552 , \30555 , \30557 );
and \U$22222 ( \30559 , \30558 , \30000 );
or \U$22223 ( \30560 , \30550 , \30559 );
and \U$22225 ( \30561 , \30560 , 1'b1 );
or \U$22227 ( \30562 , \30561 , 1'b0 );
buf \U$22228 ( \30563 , \30562 );
_DC r23df0_GF_IsGateDCbyConstraint ( \30564_nR23df0 , \30563 , \21944 );
buf \U$22229 ( \30565 , \30564_nR23df0 );
buf \U$22230 ( \30566 , \28249 );
not \U$22231 ( \30567 , \30566 );
and \U$22232 ( \30568 , RIe2346c8_6256, \30567 );
not \U$22233 ( \30569 , RIe2346c8_6256);
or \U$22234 ( \30570 , \30569 , \29801 );
not \U$22235 ( \30571 , \29916 );
and \U$22236 ( \30572 , \28276 , \30571 );
not \U$22237 ( \30573 , \30572 );
not \U$22238 ( \30574 , \29882 );
or \U$22239 ( \30575 , \29452 , \30574 );
nand \U$22240 ( \30576 , \30570 , \30573 , \30575 );
and \U$22241 ( \30577 , \30576 , \30566 );
or \U$22242 ( \30578 , \30568 , \30577 );
and \U$22244 ( \30579 , \30578 , 1'b1 );
or \U$22246 ( \30580 , \30579 , 1'b0 );
buf \U$22247 ( \30581 , \30580 );
_DC r23df2_GF_IsGateDCbyConstraint ( \30582_nR23df2 , \30581 , \21944 );
buf \U$22248 ( \30583 , \30582_nR23df2 );
not \U$22249 ( \30584 , \27363 );
and \U$22250 ( \30585 , RIe232a30_6257, \30584 );
not \U$22251 ( \30586 , RIe232a30_6257);
or \U$22252 ( \30587 , \30586 , \29986 );
not \U$22253 ( \30588 , \29897 );
and \U$22254 ( \30589 , \28295 , \30588 );
not \U$22255 ( \30590 , \30589 );
not \U$22256 ( \30591 , \29901 );
or \U$22257 ( \30592 , \29470 , \30591 );
nand \U$22258 ( \30593 , \30587 , \30590 , \30592 );
and \U$22259 ( \30594 , \30593 , \27363 );
or \U$22260 ( \30595 , \30585 , \30594 );
and \U$22262 ( \30596 , \30595 , 1'b1 );
or \U$22264 ( \30597 , \30596 , 1'b0 );
buf \U$22265 ( \30598 , \30597 );
_DC r23df4_GF_IsGateDCbyConstraint ( \30599_nR23df4 , \30598 , \21944 );
buf \U$22266 ( \30600 , \30599_nR23df4 );
buf \U$22267 ( \30601 , \28889 );
not \U$22268 ( \30602 , \30601 );
and \U$22269 ( \30603 , RIe230bb8_6258, \30602 );
not \U$22270 ( \30604 , RIe230bb8_6258);
or \U$22271 ( \30605 , \30604 , \29842 );
not \U$22272 ( \30606 , \29803 );
and \U$22273 ( \30607 , \28314 , \30606 );
not \U$22274 ( \30608 , \30607 );
not \U$22275 ( \30609 , \29901 );
or \U$22276 ( \30610 , \29488 , \30609 );
nand \U$22277 ( \30611 , \30605 , \30608 , \30610 );
and \U$22278 ( \30612 , \30611 , \30601 );
or \U$22279 ( \30613 , \30603 , \30612 );
and \U$22281 ( \30614 , \30613 , 1'b1 );
or \U$22283 ( \30615 , \30614 , 1'b0 );
buf \U$22284 ( \30616 , \30615 );
_DC r23df6_GF_IsGateDCbyConstraint ( \30617_nR23df6 , \30616 , \21944 );
buf \U$22285 ( \30618 , \30617_nR23df6 );
not \U$22286 ( \30619 , \30566 );
and \U$22287 ( \30620 , RIe465cb0_6259, \30619 );
not \U$22288 ( \30621 , RIe465cb0_6259);
or \U$22289 ( \30622 , \30621 , \29801 );
not \U$22290 ( \30623 , \30117 );
and \U$22291 ( \30624 , \28333 , \30623 );
not \U$22292 ( \30625 , \30624 );
not \U$22293 ( \30626 , \29808 );
or \U$22294 ( \30627 , \29506 , \30626 );
nand \U$22295 ( \30628 , \30622 , \30625 , \30627 );
and \U$22296 ( \30629 , \30628 , \30566 );
or \U$22297 ( \30630 , \30620 , \30629 );
and \U$22299 ( \30631 , \30630 , 1'b1 );
or \U$22301 ( \30632 , \30631 , 1'b0 );
buf \U$22302 ( \30633 , \30632 );
_DC r23df8_GF_IsGateDCbyConstraint ( \30634_nR23df8 , \30633 , \21944 );
buf \U$22303 ( \30635 , \30634_nR23df8 );
not \U$22304 ( \30636 , \27458 );
and \U$22305 ( \30637 , RIe4664a8_6260, \30636 );
not \U$22306 ( \30638 , RIe4664a8_6260);
or \U$22307 ( \30639 , \30638 , \29822 );
not \U$22308 ( \30640 , \29897 );
and \U$22309 ( \30641 , \28352 , \30640 );
not \U$22310 ( \30642 , \30641 );
not \U$22311 ( \30643 , \29901 );
or \U$22312 ( \30644 , \29524 , \30643 );
nand \U$22313 ( \30645 , \30639 , \30642 , \30644 );
and \U$22314 ( \30646 , \30645 , \27458 );
or \U$22315 ( \30647 , \30637 , \30646 );
and \U$22317 ( \30648 , \30647 , 1'b1 );
or \U$22319 ( \30649 , \30648 , 1'b0 );
buf \U$22320 ( \30650 , \30649 );
_DC r23dfa_GF_IsGateDCbyConstraint ( \30651_nR23dfa , \30650 , \21944 );
buf \U$22321 ( \30652 , \30651_nR23dfa );
not \U$22322 ( \30653 , \30601 );
and \U$22323 ( \30654 , RIe466ca0_6261, \30653 );
not \U$22324 ( \30655 , RIe466ca0_6261);
or \U$22325 ( \30656 , \30655 , \29842 );
not \U$22326 ( \30657 , \29897 );
and \U$22327 ( \30658 , \28372 , \30657 );
not \U$22328 ( \30659 , \30658 );
not \U$22329 ( \30660 , \29882 );
or \U$22330 ( \30661 , \29542 , \30660 );
nand \U$22331 ( \30662 , \30656 , \30659 , \30661 );
and \U$22332 ( \30663 , \30662 , \30601 );
or \U$22333 ( \30664 , \30654 , \30663 );
and \U$22335 ( \30665 , \30664 , 1'b1 );
or \U$22337 ( \30666 , \30665 , 1'b0 );
buf \U$22338 ( \30667 , \30666 );
_DC r23dfe_GF_IsGateDCbyConstraint ( \30668_nR23dfe , \30667 , \21944 );
buf \U$22339 ( \30669 , \30668_nR23dfe );
not \U$22340 ( \30670 , \30566 );
and \U$22341 ( \30671 , RIe467498_6262, \30670 );
not \U$22342 ( \30672 , RIe467498_6262);
or \U$22343 ( \30673 , \30672 , \29860 );
not \U$22344 ( \30674 , \29897 );
and \U$22345 ( \30675 , \28392 , \30674 );
not \U$22346 ( \30676 , \30675 );
not \U$22347 ( \30677 , \29901 );
or \U$22348 ( \30678 , \29560 , \30677 );
nand \U$22349 ( \30679 , \30673 , \30676 , \30678 );
and \U$22350 ( \30680 , \30679 , \30566 );
or \U$22351 ( \30681 , \30671 , \30680 );
and \U$22353 ( \30682 , \30681 , 1'b1 );
or \U$22355 ( \30683 , \30682 , 1'b0 );
buf \U$22356 ( \30684 , \30683 );
_DC r23e00_GF_IsGateDCbyConstraint ( \30685_nR23e00 , \30684 , \21944 );
buf \U$22357 ( \30686 , \30685_nR23e00 );
not \U$22358 ( \30687 , \27363 );
and \U$22359 ( \30688 , RIe467c90_6263, \30687 );
not \U$22360 ( \30689 , RIe467c90_6263);
or \U$22361 ( \30690 , \30689 , \29801 );
not \U$22362 ( \30691 , \29803 );
and \U$22363 ( \30692 , \28412 , \30691 );
not \U$22364 ( \30693 , \30692 );
not \U$22365 ( \30694 , \29901 );
or \U$22366 ( \30695 , \29579 , \30694 );
nand \U$22367 ( \30696 , \30690 , \30693 , \30695 );
and \U$22368 ( \30697 , \30696 , \27363 );
or \U$22369 ( \30698 , \30688 , \30697 );
and \U$22371 ( \30699 , \30698 , 1'b1 );
or \U$22373 ( \30700 , \30699 , 1'b0 );
buf \U$22374 ( \30701 , \30700 );
_DC r23e02_GF_IsGateDCbyConstraint ( \30702_nR23e02 , \30701 , \21944 );
buf \U$22375 ( \30703 , \30702_nR23e02 );
not \U$22376 ( \30704 , \30601 );
and \U$22377 ( \30705 , RIe468488_6264, \30704 );
not \U$22378 ( \30706 , RIe468488_6264);
or \U$22379 ( \30707 , \30706 , \29801 );
not \U$22380 ( \30708 , \29916 );
and \U$22381 ( \30709 , \28432 , \30708 );
not \U$22382 ( \30710 , \30709 );
not \U$22383 ( \30711 , \29882 );
or \U$22384 ( \30712 , \29597 , \30711 );
nand \U$22385 ( \30713 , \30707 , \30710 , \30712 );
and \U$22386 ( \30714 , \30713 , \30601 );
or \U$22387 ( \30715 , \30705 , \30714 );
and \U$22389 ( \30716 , \30715 , 1'b1 );
or \U$22391 ( \30717 , \30716 , 1'b0 );
buf \U$22392 ( \30718 , \30717 );
_DC r23e04_GF_IsGateDCbyConstraint ( \30719_nR23e04 , \30718 , \21944 );
buf \U$22393 ( \30720 , \30719_nR23e04 );
not \U$22394 ( \30721 , \30566 );
and \U$22395 ( \30722 , RIe468c80_6265, \30721 );
not \U$22396 ( \30723 , RIe468c80_6265);
or \U$22397 ( \30724 , \30723 , \29986 );
not \U$22398 ( \30725 , \29897 );
and \U$22399 ( \30726 , \28452 , \30725 );
not \U$22400 ( \30727 , \30726 );
not \U$22401 ( \30728 , \29901 );
or \U$22402 ( \30729 , \29615 , \30728 );
nand \U$22403 ( \30730 , \30724 , \30727 , \30729 );
and \U$22404 ( \30731 , \30730 , \30566 );
or \U$22405 ( \30732 , \30722 , \30731 );
and \U$22407 ( \30733 , \30732 , 1'b1 );
or \U$22409 ( \30734 , \30733 , 1'b0 );
buf \U$22410 ( \30735 , \30734 );
_DC r23e06_GF_IsGateDCbyConstraint ( \30736_nR23e06 , \30735 , \21944 );
buf \U$22411 ( \30737 , \30736_nR23e06 );
not \U$22412 ( \30738 , \27363 );
and \U$22413 ( \30739 , RIe469478_6266, \30738 );
not \U$22414 ( \30740 , RIe469478_6266);
or \U$22415 ( \30741 , \30740 , \29986 );
not \U$22416 ( \30742 , \29824 );
and \U$22417 ( \30743 , \28471 , \30742 );
not \U$22418 ( \30744 , \30743 );
not \U$22419 ( \30745 , \29882 );
or \U$22420 ( \30746 , \29633 , \30745 );
nand \U$22421 ( \30747 , \30741 , \30744 , \30746 );
and \U$22422 ( \30748 , \30747 , \27363 );
or \U$22423 ( \30749 , \30739 , \30748 );
and \U$22425 ( \30750 , \30749 , 1'b1 );
or \U$22427 ( \30751 , \30750 , 1'b0 );
buf \U$22428 ( \30752 , \30751 );
_DC r23e08_GF_IsGateDCbyConstraint ( \30753_nR23e08 , \30752 , \21944 );
buf \U$22429 ( \30754 , \30753_nR23e08 );
not \U$22430 ( \30755 , \30601 );
and \U$22431 ( \30756 , RIe469c70_6267, \30755 );
not \U$22432 ( \30757 , RIe469c70_6267);
or \U$22433 ( \30758 , \30757 , \29842 );
not \U$22434 ( \30759 , \29897 );
and \U$22435 ( \30760 , \28490 , \30759 );
not \U$22436 ( \30761 , \30760 );
not \U$22437 ( \30762 , \29882 );
or \U$22438 ( \30763 , \29651 , \30762 );
nand \U$22439 ( \30764 , \30758 , \30761 , \30763 );
and \U$22440 ( \30765 , \30764 , \30601 );
or \U$22441 ( \30766 , \30756 , \30765 );
and \U$22443 ( \30767 , \30766 , 1'b1 );
or \U$22445 ( \30768 , \30767 , 1'b0 );
buf \U$22446 ( \30769 , \30768 );
_DC r23e0a_GF_IsGateDCbyConstraint ( \30770_nR23e0a , \30769 , \21944 );
buf \U$22447 ( \30771 , \30770_nR23e0a );
not \U$22448 ( \30772 , \30566 );
and \U$22449 ( \30773 , RIe46a468_6268, \30772 );
not \U$22450 ( \30774 , RIe46a468_6268);
or \U$22451 ( \30775 , \30774 , \29860 );
not \U$22452 ( \30776 , \29897 );
and \U$22453 ( \30777 , \28510 , \30776 );
not \U$22454 ( \30778 , \30777 );
not \U$22455 ( \30779 , \29901 );
or \U$22456 ( \30780 , \29669 , \30779 );
nand \U$22457 ( \30781 , \30775 , \30778 , \30780 );
and \U$22458 ( \30782 , \30781 , \30566 );
or \U$22459 ( \30783 , \30773 , \30782 );
and \U$22461 ( \30784 , \30783 , 1'b1 );
or \U$22463 ( \30785 , \30784 , 1'b0 );
buf \U$22464 ( \30786 , \30785 );
_DC r23e0c_GF_IsGateDCbyConstraint ( \30787_nR23e0c , \30786 , \21944 );
buf \U$22465 ( \30788 , \30787_nR23e0c );
buf \U$22466 ( \30789 , \28483 );
not \U$22467 ( \30790 , \30789 );
and \U$22468 ( \30791 , RIe46ac60_6269, \30790 );
not \U$22469 ( \30792 , RIe46ac60_6269);
or \U$22470 ( \30793 , \30792 , \29860 );
not \U$22471 ( \30794 , \29824 );
and \U$22472 ( \30795 , \28529 , \30794 );
not \U$22473 ( \30796 , \30795 );
not \U$22474 ( \30797 , \29901 );
or \U$22475 ( \30798 , \29687 , \30797 );
nand \U$22476 ( \30799 , \30793 , \30796 , \30798 );
and \U$22477 ( \30800 , \30799 , \30789 );
or \U$22478 ( \30801 , \30791 , \30800 );
and \U$22480 ( \30802 , \30801 , 1'b1 );
or \U$22482 ( \30803 , \30802 , 1'b0 );
buf \U$22483 ( \30804 , \30803 );
_DC r23e0e_GF_IsGateDCbyConstraint ( \30805_nR23e0e , \30804 , \21944 );
buf \U$22484 ( \30806 , \30805_nR23e0e );
not \U$22485 ( \30807 , \30601 );
and \U$22486 ( \30808 , RIe46b458_6270, \30807 );
not \U$22487 ( \30809 , RIe46b458_6270);
or \U$22488 ( \30810 , \30809 , \29986 );
not \U$22489 ( \30811 , \29824 );
and \U$22490 ( \30812 , \28551 , \30811 );
not \U$22491 ( \30813 , \30812 );
not \U$22492 ( \30814 , \29882 );
or \U$22493 ( \30815 , \29705 , \30814 );
nand \U$22494 ( \30816 , \30810 , \30813 , \30815 );
and \U$22495 ( \30817 , \30816 , \30601 );
or \U$22496 ( \30818 , \30808 , \30817 );
and \U$22498 ( \30819 , \30818 , 1'b1 );
or \U$22500 ( \30820 , \30819 , 1'b0 );
buf \U$22501 ( \30821 , \30820 );
_DC r23e10_GF_IsGateDCbyConstraint ( \30822_nR23e10 , \30821 , \21944 );
buf \U$22502 ( \30823 , \30822_nR23e10 );
not \U$22503 ( \30824 , \30566 );
and \U$22504 ( \30825 , RIe46bc50_6271, \30824 );
not \U$22505 ( \30826 , RIe46bc50_6271);
or \U$22506 ( \30827 , \30826 , \29842 );
not \U$22507 ( \30828 , \29803 );
and \U$22508 ( \30829 , \28571 , \30828 );
not \U$22509 ( \30830 , \30829 );
not \U$22510 ( \30831 , \29882 );
or \U$22511 ( \30832 , \29723 , \30831 );
nand \U$22512 ( \30833 , \30827 , \30830 , \30832 );
and \U$22513 ( \30834 , \30833 , \30566 );
or \U$22514 ( \30835 , \30825 , \30834 );
and \U$22516 ( \30836 , \30835 , 1'b1 );
or \U$22518 ( \30837 , \30836 , 1'b0 );
buf \U$22519 ( \30838 , \30837 );
_DC r23e14_GF_IsGateDCbyConstraint ( \30839_nR23e14 , \30838 , \21944 );
buf \U$22520 ( \30840 , \30839_nR23e14 );
not \U$22521 ( \30841 , \30789 );
and \U$22522 ( \30842 , RIe46c448_6272, \30841 );
not \U$22523 ( \30843 , RIe46c448_6272);
or \U$22524 ( \30844 , \30843 , \29822 );
not \U$22525 ( \30845 , \30117 );
and \U$22526 ( \30846 , \28589 , \30845 );
not \U$22527 ( \30847 , \30846 );
not \U$22528 ( \30848 , \29882 );
or \U$22529 ( \30849 , \29741 , \30848 );
nand \U$22530 ( \30850 , \30844 , \30847 , \30849 );
and \U$22531 ( \30851 , \30850 , \30789 );
or \U$22532 ( \30852 , \30842 , \30851 );
and \U$22534 ( \30853 , \30852 , 1'b1 );
or \U$22536 ( \30854 , \30853 , 1'b0 );
buf \U$22537 ( \30855 , \30854 );
_DC r23e16_GF_IsGateDCbyConstraint ( \30856_nR23e16 , \30855 , \21944 );
buf \U$22538 ( \30857 , \30856_nR23e16 );
not \U$22539 ( \30858 , \30601 );
and \U$22540 ( \30859 , RIe46cc40_6273, \30858 );
not \U$22541 ( \30860 , RIe46cc40_6273);
or \U$22542 ( \30861 , \30860 , \29986 );
not \U$22543 ( \30862 , \30117 );
and \U$22544 ( \30863 , \28608 , \30862 );
not \U$22545 ( \30864 , \30863 );
not \U$22546 ( \30865 , \29901 );
or \U$22547 ( \30866 , \29759 , \30865 );
nand \U$22548 ( \30867 , \30861 , \30864 , \30866 );
and \U$22549 ( \30868 , \30867 , \30601 );
or \U$22550 ( \30869 , \30859 , \30868 );
and \U$22552 ( \30870 , \30869 , 1'b1 );
or \U$22554 ( \30871 , \30870 , 1'b0 );
buf \U$22555 ( \30872 , \30871 );
_DC r23e18_GF_IsGateDCbyConstraint ( \30873_nR23e18 , \30872 , \21944 );
buf \U$22556 ( \30874 , \30873_nR23e18 );
not \U$22557 ( \30875 , \30566 );
and \U$22558 ( \30876 , RIe46d438_6274, \30875 );
not \U$22559 ( \30877 , RIe46d438_6274);
or \U$22560 ( \30878 , \30877 , \29842 );
not \U$22561 ( \30879 , \29916 );
and \U$22562 ( \30880 , \28626 , \30879 );
not \U$22563 ( \30881 , \30880 );
not \U$22564 ( \30882 , \29901 );
or \U$22565 ( \30883 , \29777 , \30882 );
nand \U$22566 ( \30884 , \30878 , \30881 , \30883 );
and \U$22567 ( \30885 , \30884 , \30566 );
or \U$22568 ( \30886 , \30876 , \30885 );
and \U$22570 ( \30887 , \30886 , 1'b1 );
or \U$22572 ( \30888 , \30887 , 1'b0 );
buf \U$22573 ( \30889 , \30888 );
_DC r23e1a_GF_IsGateDCbyConstraint ( \30890_nR23e1a , \30889 , \21944 );
buf \U$22574 ( \30891 , \30890_nR23e1a );
not \U$22575 ( \30892 , \30789 );
and \U$22576 ( \30893 , RIe46dc30_6275, \30892 );
not \U$22577 ( \30894 , RIe46dc30_6275);
nand \U$22578 ( \30895 , \27383 , \27380 );
not \U$22579 ( \30896 , \27385 );
or \U$22580 ( \30897 , \30895 , \30896 );
nand \U$22581 ( \30898 , \27372 , \27370 );
not \U$22582 ( \30899 , \30898 );
nand \U$22583 ( \30900 , \27362 , \30899 );
nand \U$22584 ( \30901 , \30897 , \30900 );
buf \U$22585 ( \30902 , \30901 );
or \U$22586 ( \30903 , \30894 , \30902 );
not \U$22587 ( \30904 , \30900 );
buf \U$22588 ( \30905 , \30904 );
nand \U$22589 ( \30906 , \27393 , \30905 );
not \U$22590 ( \30907 , \30897 );
buf \U$22591 ( \30908 , \30907 );
nand \U$22592 ( \30909 , \27395 , \30908 );
nand \U$22593 ( \30910 , \30903 , \30906 , \30909 );
and \U$22594 ( \30911 , \30910 , \30789 );
or \U$22595 ( \30912 , \30893 , \30911 );
and \U$22597 ( \30913 , \30912 , 1'b1 );
or \U$22599 ( \30914 , \30913 , 1'b0 );
buf \U$22600 ( \30915 , \30914 );
_DC r23e24_GF_IsGateDCbyConstraint ( \30916_nR23e24 , \30915 , \21944 );
buf \U$22601 ( \30917 , \30916_nR23e24 );
not \U$22602 ( \30918 , \30601 );
and \U$22603 ( \30919 , RIe46e428_6276, \30918 );
not \U$22604 ( \30920 , RIe46e428_6276);
buf \U$22605 ( \30921 , \30901 );
or \U$22606 ( \30922 , \30920 , \30921 );
buf \U$22607 ( \30923 , \30904 );
nand \U$22608 ( \30924 , \27424 , \30923 );
nand \U$22609 ( \30925 , \27427 , \30908 );
nand \U$22610 ( \30926 , \30922 , \30924 , \30925 );
and \U$22611 ( \30927 , \30926 , \30601 );
or \U$22612 ( \30928 , \30919 , \30927 );
and \U$22614 ( \30929 , \30928 , 1'b1 );
or \U$22616 ( \30930 , \30929 , 1'b0 );
buf \U$22617 ( \30931 , \30930 );
_DC r23e3a_GF_IsGateDCbyConstraint ( \30932_nR23e3a , \30931 , \21944 );
buf \U$22618 ( \30933 , \30932_nR23e3a );
not \U$22619 ( \30934 , \30566 );
and \U$22620 ( \30935 , RIe46ec20_6277, \30934 );
not \U$22621 ( \30936 , RIe46ec20_6277);
buf \U$22622 ( \30937 , \30901 );
or \U$22623 ( \30938 , \30936 , \30937 );
nand \U$22624 ( \30939 , \27444 , \30904 );
buf \U$22625 ( \30940 , \30907 );
nand \U$22626 ( \30941 , \27446 , \30940 );
nand \U$22627 ( \30942 , \30938 , \30939 , \30941 );
and \U$22628 ( \30943 , \30942 , \30566 );
or \U$22629 ( \30944 , \30935 , \30943 );
and \U$22631 ( \30945 , \30944 , 1'b1 );
or \U$22633 ( \30946 , \30945 , 1'b0 );
buf \U$22634 ( \30947 , \30946 );
_DC r23e50_GF_IsGateDCbyConstraint ( \30948_nR23e50 , \30947 , \21944 );
buf \U$22635 ( \30949 , \30948_nR23e50 );
not \U$22636 ( \30950 , \30789 );
and \U$22637 ( \30951 , RIe46f418_6278, \30950 );
not \U$22638 ( \30952 , RIe46f418_6278);
buf \U$22639 ( \30953 , \30901 );
or \U$22640 ( \30954 , \30952 , \30953 );
buf \U$22641 ( \30955 , \30904 );
nand \U$22642 ( \30956 , \27465 , \30955 );
buf \U$22643 ( \30957 , \30907 );
nand \U$22644 ( \30958 , \27467 , \30957 );
nand \U$22645 ( \30959 , \30954 , \30956 , \30958 );
and \U$22646 ( \30960 , \30959 , \30789 );
or \U$22647 ( \30961 , \30951 , \30960 );
and \U$22649 ( \30962 , \30961 , 1'b1 );
or \U$22651 ( \30963 , \30962 , 1'b0 );
buf \U$22652 ( \30964 , \30963 );
_DC r23e66_GF_IsGateDCbyConstraint ( \30965_nR23e66 , \30964 , \21944 );
buf \U$22653 ( \30966 , \30965_nR23e66 );
not \U$22654 ( \30967 , \30601 );
and \U$22655 ( \30968 , RIe46fc10_6279, \30967 );
not \U$22656 ( \30969 , RIe46fc10_6279);
or \U$22657 ( \30970 , \30969 , \30902 );
buf \U$22658 ( \30971 , \30904 );
nand \U$22659 ( \30972 , \27484 , \30971 );
nand \U$22660 ( \30973 , \27486 , \30940 );
nand \U$22661 ( \30974 , \30970 , \30972 , \30973 );
and \U$22662 ( \30975 , \30974 , \30601 );
or \U$22663 ( \30976 , \30968 , \30975 );
and \U$22665 ( \30977 , \30976 , 1'b1 );
or \U$22667 ( \30978 , \30977 , 1'b0 );
buf \U$22668 ( \30979 , \30978 );
_DC r23e7c_GF_IsGateDCbyConstraint ( \30980_nR23e7c , \30979 , \21944 );
buf \U$22669 ( \30981 , \30980_nR23e7c );
not \U$22670 ( \30982 , \30566 );
and \U$22671 ( \30983 , RIe470408_6280, \30982 );
not \U$22672 ( \30984 , RIe470408_6280);
or \U$22673 ( \30985 , \30984 , \30921 );
nand \U$22674 ( \30986 , \27504 , \30923 );
buf \U$22675 ( \30987 , \30907 );
nand \U$22676 ( \30988 , \27507 , \30987 );
nand \U$22677 ( \30989 , \30985 , \30986 , \30988 );
and \U$22678 ( \30990 , \30989 , \30566 );
or \U$22679 ( \30991 , \30983 , \30990 );
and \U$22681 ( \30992 , \30991 , 1'b1 );
or \U$22683 ( \30993 , \30992 , 1'b0 );
buf \U$22684 ( \30994 , \30993 );
_DC r23e92_GF_IsGateDCbyConstraint ( \30995_nR23e92 , \30994 , \21944 );
buf \U$22685 ( \30996 , \30995_nR23e92 );
not \U$22686 ( \30997 , \30789 );
and \U$22687 ( \30998 , RIe470c00_6281, \30997 );
not \U$22688 ( \30999 , RIe470c00_6281);
or \U$22689 ( \31000 , \30999 , \30937 );
nand \U$22690 ( \31001 , \27525 , \30955 );
nand \U$22691 ( \31002 , \27527 , \30908 );
nand \U$22692 ( \31003 , \31000 , \31001 , \31002 );
and \U$22693 ( \31004 , \31003 , \30789 );
or \U$22694 ( \31005 , \30998 , \31004 );
and \U$22696 ( \31006 , \31005 , 1'b1 );
or \U$22698 ( \31007 , \31006 , 1'b0 );
buf \U$22699 ( \31008 , \31007 );
_DC r23e9c_GF_IsGateDCbyConstraint ( \31009_nR23e9c , \31008 , \21944 );
buf \U$22700 ( \31010 , \31009_nR23e9c );
not \U$22701 ( \31011 , \30601 );
and \U$22702 ( \31012 , RIe4713f8_6282, \31011 );
not \U$22703 ( \31013 , RIe4713f8_6282);
or \U$22704 ( \31014 , \31013 , \30921 );
nand \U$22705 ( \31015 , \27543 , \30923 );
nand \U$22706 ( \31016 , \27546 , \30908 );
nand \U$22707 ( \31017 , \31014 , \31015 , \31016 );
and \U$22708 ( \31018 , \31017 , \30601 );
or \U$22709 ( \31019 , \31012 , \31018 );
and \U$22711 ( \31020 , \31019 , 1'b1 );
or \U$22713 ( \31021 , \31020 , 1'b0 );
buf \U$22714 ( \31022 , \31021 );
_DC r23e9e_GF_IsGateDCbyConstraint ( \31023_nR23e9e , \31022 , \21944 );
buf \U$22715 ( \31024 , \31023_nR23e9e );
not \U$22716 ( \31025 , \30566 );
and \U$22717 ( \31026 , RIe471bf0_6283, \31025 );
not \U$22718 ( \31027 , RIe471bf0_6283);
or \U$22719 ( \31028 , \31027 , \30902 );
nand \U$22720 ( \31029 , \27565 , \30971 );
nand \U$22721 ( \31030 , \27568 , \30957 );
nand \U$22722 ( \31031 , \31028 , \31029 , \31030 );
and \U$22723 ( \31032 , \31031 , \30566 );
or \U$22724 ( \31033 , \31026 , \31032 );
and \U$22726 ( \31034 , \31033 , 1'b1 );
or \U$22728 ( \31035 , \31034 , 1'b0 );
buf \U$22729 ( \31036 , \31035 );
_DC r23ea0_GF_IsGateDCbyConstraint ( \31037_nR23ea0 , \31036 , \21944 );
buf \U$22730 ( \31038 , \31037_nR23ea0 );
not \U$22731 ( \31039 , \30789 );
and \U$22732 ( \31040 , RIe4723e8_6284, \31039 );
not \U$22733 ( \31041 , RIe4723e8_6284);
buf \U$22734 ( \31042 , \30901 );
or \U$22735 ( \31043 , \31041 , \31042 );
nand \U$22736 ( \31044 , \27585 , \30905 );
nand \U$22737 ( \31045 , \27588 , \30940 );
nand \U$22738 ( \31046 , \31043 , \31044 , \31045 );
and \U$22739 ( \31047 , \31046 , \30789 );
or \U$22740 ( \31048 , \31040 , \31047 );
and \U$22742 ( \31049 , \31048 , 1'b1 );
or \U$22744 ( \31050 , \31049 , 1'b0 );
buf \U$22745 ( \31051 , \31050 );
_DC r23ea2_GF_IsGateDCbyConstraint ( \31052_nR23ea2 , \31051 , \21944 );
buf \U$22746 ( \31053 , \31052_nR23ea2 );
not \U$22747 ( \31054 , \30601 );
and \U$22748 ( \31055 , RIe472bf8_6285, \31054 );
not \U$22749 ( \31056 , RIe472bf8_6285);
or \U$22750 ( \31057 , \31056 , \31042 );
nand \U$22751 ( \31058 , \27606 , \30905 );
nand \U$22752 ( \31059 , \27609 , \30987 );
nand \U$22753 ( \31060 , \31057 , \31058 , \31059 );
and \U$22754 ( \31061 , \31060 , \30601 );
or \U$22755 ( \31062 , \31055 , \31061 );
and \U$22757 ( \31063 , \31062 , 1'b1 );
or \U$22759 ( \31064 , \31063 , 1'b0 );
buf \U$22760 ( \31065 , \31064 );
_DC r23e26_GF_IsGateDCbyConstraint ( \31066_nR23e26 , \31065 , \21944 );
buf \U$22761 ( \31067 , \31066_nR23e26 );
not \U$22762 ( \31068 , \30566 );
and \U$22763 ( \31069 , RIe4733f0_6286, \31068 );
not \U$22764 ( \31070 , RIe4733f0_6286);
or \U$22765 ( \31071 , \31070 , \30953 );
nand \U$22766 ( \31072 , \27625 , \30904 );
nand \U$22767 ( \31073 , \27628 , \30940 );
nand \U$22768 ( \31074 , \31071 , \31072 , \31073 );
and \U$22769 ( \31075 , \31074 , \30566 );
or \U$22770 ( \31076 , \31069 , \31075 );
and \U$22772 ( \31077 , \31076 , 1'b1 );
or \U$22774 ( \31078 , \31077 , 1'b0 );
buf \U$22775 ( \31079 , \31078 );
_DC r23e28_GF_IsGateDCbyConstraint ( \31080_nR23e28 , \31079 , \21944 );
buf \U$22776 ( \31081 , \31080_nR23e28 );
not \U$22777 ( \31082 , \30789 );
and \U$22778 ( \31083 , RIe473be8_6287, \31082 );
not \U$22779 ( \31084 , RIe473be8_6287);
or \U$22780 ( \31085 , \31084 , \30937 );
nand \U$22781 ( \31086 , \27645 , \30923 );
nand \U$22782 ( \31087 , \27648 , \30987 );
nand \U$22783 ( \31088 , \31085 , \31086 , \31087 );
and \U$22784 ( \31089 , \31088 , \30789 );
or \U$22785 ( \31090 , \31083 , \31089 );
and \U$22787 ( \31091 , \31090 , 1'b1 );
or \U$22789 ( \31092 , \31091 , 1'b0 );
buf \U$22790 ( \31093 , \31092 );
_DC r23e2a_GF_IsGateDCbyConstraint ( \31094_nR23e2a , \31093 , \21944 );
buf \U$22791 ( \31095 , \31094_nR23e2a );
not \U$22792 ( \31096 , \30601 );
and \U$22793 ( \31097 , RIe4743e0_6288, \31096 );
not \U$22794 ( \31098 , RIe4743e0_6288);
or \U$22795 ( \31099 , \31098 , \30953 );
nand \U$22796 ( \31100 , \27665 , \30971 );
nand \U$22797 ( \31101 , \27668 , \30957 );
nand \U$22798 ( \31102 , \31099 , \31100 , \31101 );
and \U$22799 ( \31103 , \31102 , \30601 );
or \U$22800 ( \31104 , \31097 , \31103 );
and \U$22802 ( \31105 , \31104 , 1'b1 );
or \U$22804 ( \31106 , \31105 , 1'b0 );
buf \U$22805 ( \31107 , \31106 );
_DC r23e2c_GF_IsGateDCbyConstraint ( \31108_nR23e2c , \31107 , \21944 );
buf \U$22806 ( \31109 , \31108_nR23e2c );
not \U$22807 ( \31110 , \30566 );
and \U$22808 ( \31111 , RIe474bd8_6289, \31110 );
not \U$22809 ( \31112 , RIe474bd8_6289);
or \U$22810 ( \31113 , \31112 , \30921 );
nand \U$22811 ( \31114 , \27684 , \30923 );
nand \U$22812 ( \31115 , \27686 , \30940 );
nand \U$22813 ( \31116 , \31113 , \31114 , \31115 );
and \U$22814 ( \31117 , \31116 , \30566 );
or \U$22815 ( \31118 , \31111 , \31117 );
and \U$22817 ( \31119 , \31118 , 1'b1 );
or \U$22819 ( \31120 , \31119 , 1'b0 );
buf \U$22820 ( \31121 , \31120 );
_DC r23e2e_GF_IsGateDCbyConstraint ( \31122_nR23e2e , \31121 , \21944 );
buf \U$22821 ( \31123 , \31122_nR23e2e );
not \U$22822 ( \31124 , \30789 );
and \U$22823 ( \31125 , RIe4753d0_6290, \31124 );
not \U$22824 ( \31126 , RIe4753d0_6290);
or \U$22825 ( \31127 , \31126 , \30902 );
nand \U$22826 ( \31128 , \27702 , \30955 );
nand \U$22827 ( \31129 , \27704 , \30987 );
nand \U$22828 ( \31130 , \31127 , \31128 , \31129 );
and \U$22829 ( \31131 , \31130 , \30789 );
or \U$22830 ( \31132 , \31125 , \31131 );
and \U$22832 ( \31133 , \31132 , 1'b1 );
or \U$22834 ( \31134 , \31133 , 1'b0 );
buf \U$22835 ( \31135 , \31134 );
_DC r23e30_GF_IsGateDCbyConstraint ( \31136_nR23e30 , \31135 , \21944 );
buf \U$22836 ( \31137 , \31136_nR23e30 );
not \U$22837 ( \31138 , \30601 );
and \U$22838 ( \31139 , RIe475bc8_6291, \31138 );
not \U$22839 ( \31140 , RIe475bc8_6291);
or \U$22840 ( \31141 , \31140 , \31042 );
nand \U$22841 ( \31142 , \27720 , \30923 );
nand \U$22842 ( \31143 , \27722 , \30908 );
nand \U$22843 ( \31144 , \31141 , \31142 , \31143 );
and \U$22844 ( \31145 , \31144 , \30601 );
or \U$22845 ( \31146 , \31139 , \31145 );
and \U$22847 ( \31147 , \31146 , 1'b1 );
or \U$22849 ( \31148 , \31147 , 1'b0 );
buf \U$22850 ( \31149 , \31148 );
_DC r23e32_GF_IsGateDCbyConstraint ( \31150_nR23e32 , \31149 , \21944 );
buf \U$22851 ( \31151 , \31150_nR23e32 );
not \U$22852 ( \31152 , \29571 );
and \U$22853 ( \31153 , RIe4763c0_6292, \31152 );
not \U$22854 ( \31154 , RIe4763c0_6292);
or \U$22855 ( \31155 , \31154 , \30953 );
nand \U$22856 ( \31156 , \27738 , \30971 );
nand \U$22857 ( \31157 , \27741 , \30957 );
nand \U$22858 ( \31158 , \31155 , \31156 , \31157 );
and \U$22859 ( \31159 , \31158 , \29571 );
or \U$22860 ( \31160 , \31153 , \31159 );
and \U$22862 ( \31161 , \31160 , 1'b1 );
or \U$22864 ( \31162 , \31161 , 1'b0 );
buf \U$22865 ( \31163 , \31162 );
_DC r23e34_GF_IsGateDCbyConstraint ( \31164_nR23e34 , \31163 , \21944 );
buf \U$22866 ( \31165 , \31164_nR23e34 );
not \U$22867 ( \31166 , \30789 );
and \U$22868 ( \31167 , RIe476bb8_6293, \31166 );
not \U$22869 ( \31168 , RIe476bb8_6293);
or \U$22870 ( \31169 , \31168 , \30937 );
nand \U$22871 ( \31170 , \27757 , \30923 );
nand \U$22872 ( \31171 , \27760 , \30957 );
nand \U$22873 ( \31172 , \31169 , \31170 , \31171 );
and \U$22874 ( \31173 , \31172 , \30789 );
or \U$22875 ( \31174 , \31167 , \31173 );
and \U$22877 ( \31175 , \31174 , 1'b1 );
or \U$22879 ( \31176 , \31175 , 1'b0 );
buf \U$22880 ( \31177 , \31176 );
_DC r23e36_GF_IsGateDCbyConstraint ( \31178_nR23e36 , \31177 , \21944 );
buf \U$22881 ( \31179 , \31178_nR23e36 );
buf \U$22882 ( \31180 , \28889 );
not \U$22883 ( \31181 , \31180 );
and \U$22884 ( \31182 , RIe4773b0_6294, \31181 );
not \U$22885 ( \31183 , RIe4773b0_6294);
or \U$22886 ( \31184 , \31183 , \30937 );
nand \U$22887 ( \31185 , \27776 , \30923 );
nand \U$22888 ( \31186 , \27779 , \30940 );
nand \U$22889 ( \31187 , \31184 , \31185 , \31186 );
and \U$22890 ( \31188 , \31187 , \31180 );
or \U$22891 ( \31189 , \31182 , \31188 );
and \U$22893 ( \31190 , \31189 , 1'b1 );
or \U$22895 ( \31191 , \31190 , 1'b0 );
buf \U$22896 ( \31192 , \31191 );
_DC r23e38_GF_IsGateDCbyConstraint ( \31193_nR23e38 , \31192 , \21944 );
buf \U$22897 ( \31194 , \31193_nR23e38 );
not \U$22898 ( \31195 , \29571 );
and \U$22899 ( \31196 , RIe477ba8_6295, \31195 );
not \U$22900 ( \31197 , RIe477ba8_6295);
or \U$22901 ( \31198 , \31197 , \30902 );
nand \U$22902 ( \31199 , \27796 , \30955 );
nand \U$22903 ( \31200 , \27799 , \30940 );
nand \U$22904 ( \31201 , \31198 , \31199 , \31200 );
and \U$22905 ( \31202 , \31201 , \29571 );
or \U$22906 ( \31203 , \31196 , \31202 );
and \U$22908 ( \31204 , \31203 , 1'b1 );
or \U$22910 ( \31205 , \31204 , 1'b0 );
buf \U$22911 ( \31206 , \31205 );
_DC r23e3c_GF_IsGateDCbyConstraint ( \31207_nR23e3c , \31206 , \21944 );
buf \U$22912 ( \31208 , \31207_nR23e3c );
not \U$22913 ( \31209 , \30789 );
and \U$22914 ( \31210 , RIe4783a0_6296, \31209 );
not \U$22915 ( \31211 , RIe4783a0_6296);
or \U$22916 ( \31212 , \31211 , \31042 );
nand \U$22917 ( \31213 , \27815 , \30955 );
nand \U$22918 ( \31214 , \27817 , \30987 );
nand \U$22919 ( \31215 , \31212 , \31213 , \31214 );
and \U$22920 ( \31216 , \31215 , \30789 );
or \U$22921 ( \31217 , \31210 , \31216 );
and \U$22923 ( \31218 , \31217 , 1'b1 );
or \U$22925 ( \31219 , \31218 , 1'b0 );
buf \U$22926 ( \31220 , \31219 );
_DC r23e3e_GF_IsGateDCbyConstraint ( \31221_nR23e3e , \31220 , \21944 );
buf \U$22927 ( \31222 , \31221_nR23e3e );
not \U$22928 ( \31223 , \31180 );
and \U$22929 ( \31224 , RIe478b98_6297, \31223 );
not \U$22930 ( \31225 , RIe478b98_6297);
or \U$22931 ( \31226 , \31225 , \30921 );
nand \U$22932 ( \31227 , \27833 , \30955 );
nand \U$22933 ( \31228 , \27835 , \30908 );
nand \U$22934 ( \31229 , \31226 , \31227 , \31228 );
and \U$22935 ( \31230 , \31229 , \31180 );
or \U$22936 ( \31231 , \31224 , \31230 );
and \U$22938 ( \31232 , \31231 , 1'b1 );
or \U$22940 ( \31233 , \31232 , 1'b0 );
buf \U$22941 ( \31234 , \31233 );
_DC r23e40_GF_IsGateDCbyConstraint ( \31235_nR23e40 , \31234 , \21944 );
buf \U$22942 ( \31236 , \31235_nR23e40 );
not \U$22943 ( \31237 , \27458 );
and \U$22944 ( \31238 , RIe479390_6298, \31237 );
not \U$22945 ( \31239 , RIe479390_6298);
or \U$22946 ( \31240 , \31239 , \30953 );
nand \U$22947 ( \31241 , \27851 , \30971 );
nand \U$22948 ( \31242 , \27854 , \30940 );
nand \U$22949 ( \31243 , \31240 , \31241 , \31242 );
and \U$22950 ( \31244 , \31243 , \27458 );
or \U$22951 ( \31245 , \31238 , \31244 );
and \U$22953 ( \31246 , \31245 , 1'b1 );
or \U$22955 ( \31247 , \31246 , 1'b0 );
buf \U$22956 ( \31248 , \31247 );
_DC r23e42_GF_IsGateDCbyConstraint ( \31249_nR23e42 , \31248 , \21944 );
buf \U$22957 ( \31250 , \31249_nR23e42 );
not \U$22958 ( \31251 , \30789 );
and \U$22959 ( \31252 , RIe479b88_6299, \31251 );
not \U$22960 ( \31253 , RIe479b88_6299);
or \U$22961 ( \31254 , \31253 , \30937 );
nand \U$22962 ( \31255 , \27870 , \30905 );
nand \U$22963 ( \31256 , \27873 , \30957 );
nand \U$22964 ( \31257 , \31254 , \31255 , \31256 );
and \U$22965 ( \31258 , \31257 , \30789 );
or \U$22966 ( \31259 , \31252 , \31258 );
and \U$22968 ( \31260 , \31259 , 1'b1 );
or \U$22970 ( \31261 , \31260 , 1'b0 );
buf \U$22971 ( \31262 , \31261 );
_DC r23e44_GF_IsGateDCbyConstraint ( \31263_nR23e44 , \31262 , \21944 );
buf \U$22972 ( \31264 , \31263_nR23e44 );
not \U$22973 ( \31265 , \31180 );
and \U$22974 ( \31266 , RIe47a380_6300, \31265 );
not \U$22975 ( \31267 , RIe47a380_6300);
or \U$22976 ( \31268 , \31267 , \30921 );
nand \U$22977 ( \31269 , \27889 , \30971 );
nand \U$22978 ( \31270 , \27892 , \30987 );
nand \U$22979 ( \31271 , \31268 , \31269 , \31270 );
and \U$22980 ( \31272 , \31271 , \31180 );
or \U$22981 ( \31273 , \31266 , \31272 );
and \U$22983 ( \31274 , \31273 , 1'b1 );
or \U$22985 ( \31275 , \31274 , 1'b0 );
buf \U$22986 ( \31276 , \31275 );
_DC r23e46_GF_IsGateDCbyConstraint ( \31277_nR23e46 , \31276 , \21944 );
buf \U$22987 ( \31278 , \31277_nR23e46 );
not \U$22988 ( \31279 , \29571 );
and \U$22989 ( \31280 , RIe47ab78_6301, \31279 );
not \U$22990 ( \31281 , RIe47ab78_6301);
or \U$22991 ( \31282 , \31281 , \30902 );
nand \U$22992 ( \31283 , \27908 , \30971 );
nand \U$22993 ( \31284 , \27911 , \30987 );
nand \U$22994 ( \31285 , \31282 , \31283 , \31284 );
and \U$22995 ( \31286 , \31285 , \29571 );
or \U$22996 ( \31287 , \31280 , \31286 );
and \U$22998 ( \31288 , \31287 , 1'b1 );
or \U$23000 ( \31289 , \31288 , 1'b0 );
buf \U$23001 ( \31290 , \31289 );
_DC r23e48_GF_IsGateDCbyConstraint ( \31291_nR23e48 , \31290 , \21944 );
buf \U$23002 ( \31292 , \31291_nR23e48 );
not \U$23003 ( \31293 , \30789 );
and \U$23004 ( \31294 , RIe47b370_6302, \31293 );
not \U$23005 ( \31295 , RIe47b370_6302);
or \U$23006 ( \31296 , \31295 , \30902 );
nand \U$23007 ( \31297 , \27927 , \30905 );
nand \U$23008 ( \31298 , \27930 , \30908 );
nand \U$23009 ( \31299 , \31296 , \31297 , \31298 );
and \U$23010 ( \31300 , \31299 , \30789 );
or \U$23011 ( \31301 , \31294 , \31300 );
and \U$23013 ( \31302 , \31301 , 1'b1 );
or \U$23015 ( \31303 , \31302 , 1'b0 );
buf \U$23016 ( \31304 , \31303 );
_DC r23e4a_GF_IsGateDCbyConstraint ( \31305_nR23e4a , \31304 , \21944 );
buf \U$23017 ( \31306 , \31305_nR23e4a );
not \U$23018 ( \31307 , \31180 );
and \U$23019 ( \31308 , RIe47bb68_6303, \31307 );
not \U$23020 ( \31309 , RIe47bb68_6303);
or \U$23021 ( \31310 , \31309 , \31042 );
nand \U$23022 ( \31311 , \27947 , \30971 );
nand \U$23023 ( \31312 , \27949 , \30957 );
nand \U$23024 ( \31313 , \31310 , \31311 , \31312 );
and \U$23025 ( \31314 , \31313 , \31180 );
or \U$23026 ( \31315 , \31308 , \31314 );
and \U$23028 ( \31316 , \31315 , 1'b1 );
or \U$23030 ( \31317 , \31316 , 1'b0 );
buf \U$23031 ( \31318 , \31317 );
_DC r23e4c_GF_IsGateDCbyConstraint ( \31319_nR23e4c , \31318 , \21944 );
buf \U$23032 ( \31320 , \31319_nR23e4c );
not \U$23033 ( \31321 , \27458 );
and \U$23034 ( \31322 , RIe47c360_6304, \31321 );
not \U$23035 ( \31323 , RIe47c360_6304);
or \U$23036 ( \31324 , \31323 , \30953 );
nand \U$23037 ( \31325 , \27966 , \30905 );
nand \U$23038 ( \31326 , \27968 , \30908 );
nand \U$23039 ( \31327 , \31324 , \31325 , \31326 );
and \U$23040 ( \31328 , \31327 , \27458 );
or \U$23041 ( \31329 , \31322 , \31328 );
and \U$23043 ( \31330 , \31329 , 1'b1 );
or \U$23045 ( \31331 , \31330 , 1'b0 );
buf \U$23046 ( \31332 , \31331 );
_DC r23e4e_GF_IsGateDCbyConstraint ( \31333_nR23e4e , \31332 , \21944 );
buf \U$23047 ( \31334 , \31333_nR23e4e );
buf \U$23048 ( \31335 , \28483 );
not \U$23049 ( \31336 , \31335 );
and \U$23050 ( \31337 , RIe47cb58_6305, \31336 );
not \U$23051 ( \31338 , RIe47cb58_6305);
or \U$23052 ( \31339 , \31338 , \30921 );
nand \U$23053 ( \31340 , \27985 , \30923 );
nand \U$23054 ( \31341 , \27988 , \30957 );
nand \U$23055 ( \31342 , \31339 , \31340 , \31341 );
and \U$23056 ( \31343 , \31342 , \31335 );
or \U$23057 ( \31344 , \31337 , \31343 );
and \U$23059 ( \31345 , \31344 , 1'b1 );
or \U$23061 ( \31346 , \31345 , 1'b0 );
buf \U$23062 ( \31347 , \31346 );
_DC r23e52_GF_IsGateDCbyConstraint ( \31348_nR23e52 , \31347 , \21944 );
buf \U$23063 ( \31349 , \31348_nR23e52 );
not \U$23064 ( \31350 , \31180 );
and \U$23065 ( \31351 , RIe47d350_6306, \31350 );
not \U$23066 ( \31352 , RIe47d350_6306);
or \U$23067 ( \31353 , \31352 , \31042 );
nand \U$23068 ( \31354 , \28006 , \30905 );
nand \U$23069 ( \31355 , \28009 , \30908 );
nand \U$23070 ( \31356 , \31353 , \31354 , \31355 );
and \U$23071 ( \31357 , \31356 , \31180 );
or \U$23072 ( \31358 , \31351 , \31357 );
and \U$23074 ( \31359 , \31358 , 1'b1 );
or \U$23076 ( \31360 , \31359 , 1'b0 );
buf \U$23077 ( \31361 , \31360 );
_DC r23e54_GF_IsGateDCbyConstraint ( \31362_nR23e54 , \31361 , \21944 );
buf \U$23078 ( \31363 , \31362_nR23e54 );
not \U$23079 ( \31364 , \27458 );
and \U$23080 ( \31365 , RIe47db48_6307, \31364 );
not \U$23081 ( \31366 , RIe47db48_6307);
or \U$23082 ( \31367 , \31366 , \30902 );
nand \U$23083 ( \31368 , \28026 , \30923 );
nand \U$23084 ( \31369 , \28029 , \30987 );
nand \U$23085 ( \31370 , \31367 , \31368 , \31369 );
and \U$23086 ( \31371 , \31370 , \27458 );
or \U$23087 ( \31372 , \31365 , \31371 );
and \U$23089 ( \31373 , \31372 , 1'b1 );
or \U$23091 ( \31374 , \31373 , 1'b0 );
buf \U$23092 ( \31375 , \31374 );
_DC r23e56_GF_IsGateDCbyConstraint ( \31376_nR23e56 , \31375 , \21944 );
buf \U$23093 ( \31377 , \31376_nR23e56 );
not \U$23094 ( \31378 , \31335 );
and \U$23095 ( \31379 , RIe47e340_6308, \31378 );
not \U$23096 ( \31380 , RIe47e340_6308);
or \U$23097 ( \31381 , \31380 , \31042 );
nand \U$23098 ( \31382 , \28045 , \30971 );
nand \U$23099 ( \31383 , \28048 , \30940 );
nand \U$23100 ( \31384 , \31381 , \31382 , \31383 );
and \U$23101 ( \31385 , \31384 , \31335 );
or \U$23102 ( \31386 , \31379 , \31385 );
and \U$23104 ( \31387 , \31386 , 1'b1 );
or \U$23106 ( \31388 , \31387 , 1'b0 );
buf \U$23107 ( \31389 , \31388 );
_DC r23e58_GF_IsGateDCbyConstraint ( \31390_nR23e58 , \31389 , \21944 );
buf \U$23108 ( \31391 , \31390_nR23e58 );
not \U$23109 ( \31392 , \31180 );
and \U$23110 ( \31393 , RIe47eb38_6309, \31392 );
not \U$23111 ( \31394 , RIe47eb38_6309);
or \U$23112 ( \31395 , \31394 , \30953 );
nand \U$23113 ( \31396 , \28064 , \30971 );
nand \U$23114 ( \31397 , \28066 , \30987 );
nand \U$23115 ( \31398 , \31395 , \31396 , \31397 );
and \U$23116 ( \31399 , \31398 , \31180 );
or \U$23117 ( \31400 , \31393 , \31399 );
and \U$23119 ( \31401 , \31400 , 1'b1 );
or \U$23121 ( \31402 , \31401 , 1'b0 );
buf \U$23122 ( \31403 , \31402 );
_DC r23e5a_GF_IsGateDCbyConstraint ( \31404_nR23e5a , \31403 , \21944 );
buf \U$23123 ( \31405 , \31404_nR23e5a );
not \U$23124 ( \31406 , \29571 );
and \U$23125 ( \31407 , RIe47f330_6310, \31406 );
not \U$23126 ( \31408 , RIe47f330_6310);
or \U$23127 ( \31409 , \31408 , \30937 );
nand \U$23128 ( \31410 , \28082 , \30923 );
nand \U$23129 ( \31411 , \28085 , \30957 );
nand \U$23130 ( \31412 , \31409 , \31410 , \31411 );
and \U$23131 ( \31413 , \31412 , \29571 );
or \U$23132 ( \31414 , \31407 , \31413 );
and \U$23134 ( \31415 , \31414 , 1'b1 );
or \U$23136 ( \31416 , \31415 , 1'b0 );
buf \U$23137 ( \31417 , \31416 );
_DC r23e5c_GF_IsGateDCbyConstraint ( \31418_nR23e5c , \31417 , \21944 );
buf \U$23138 ( \31419 , \31418_nR23e5c );
not \U$23139 ( \31420 , \31335 );
and \U$23140 ( \31421 , RIe47fb28_6311, \31420 );
not \U$23141 ( \31422 , RIe47fb28_6311);
or \U$23142 ( \31423 , \31422 , \30953 );
nand \U$23143 ( \31424 , \28101 , \30955 );
nand \U$23144 ( \31425 , \28104 , \30940 );
nand \U$23145 ( \31426 , \31423 , \31424 , \31425 );
and \U$23146 ( \31427 , \31426 , \31335 );
or \U$23147 ( \31428 , \31421 , \31427 );
and \U$23149 ( \31429 , \31428 , 1'b1 );
or \U$23151 ( \31430 , \31429 , 1'b0 );
buf \U$23152 ( \31431 , \31430 );
_DC r23e5e_GF_IsGateDCbyConstraint ( \31432_nR23e5e , \31431 , \21944 );
buf \U$23153 ( \31433 , \31432_nR23e5e );
not \U$23154 ( \31434 , \31180 );
and \U$23155 ( \31435 , RIe480320_6312, \31434 );
not \U$23156 ( \31436 , RIe480320_6312);
or \U$23157 ( \31437 , \31436 , \30921 );
nand \U$23158 ( \31438 , \28120 , \30971 );
nand \U$23159 ( \31439 , \28123 , \30987 );
nand \U$23160 ( \31440 , \31437 , \31438 , \31439 );
and \U$23161 ( \31441 , \31440 , \31180 );
or \U$23162 ( \31442 , \31435 , \31441 );
and \U$23164 ( \31443 , \31442 , 1'b1 );
or \U$23166 ( \31444 , \31443 , 1'b0 );
buf \U$23167 ( \31445 , \31444 );
_DC r23e60_GF_IsGateDCbyConstraint ( \31446_nR23e60 , \31445 , \21944 );
buf \U$23168 ( \31447 , \31446_nR23e60 );
not \U$23169 ( \31448 , \29571 );
and \U$23170 ( \31449 , RIe480b18_6313, \31448 );
not \U$23171 ( \31450 , RIe480b18_6313);
or \U$23172 ( \31451 , \31450 , \30902 );
nand \U$23173 ( \31452 , \28139 , \30955 );
nand \U$23174 ( \31453 , \28142 , \30908 );
nand \U$23175 ( \31454 , \31451 , \31452 , \31453 );
and \U$23176 ( \31455 , \31454 , \29571 );
or \U$23177 ( \31456 , \31449 , \31455 );
and \U$23179 ( \31457 , \31456 , 1'b1 );
or \U$23181 ( \31458 , \31457 , 1'b0 );
buf \U$23182 ( \31459 , \31458 );
_DC r23e62_GF_IsGateDCbyConstraint ( \31460_nR23e62 , \31459 , \21944 );
buf \U$23183 ( \31461 , \31460_nR23e62 );
not \U$23184 ( \31462 , \31335 );
and \U$23185 ( \31463 , RIe481310_6314, \31462 );
not \U$23186 ( \31464 , RIe481310_6314);
or \U$23187 ( \31465 , \31464 , \31042 );
nand \U$23188 ( \31466 , \28158 , \30905 );
nand \U$23189 ( \31467 , \28161 , \30940 );
nand \U$23190 ( \31468 , \31465 , \31466 , \31467 );
and \U$23191 ( \31469 , \31468 , \31335 );
or \U$23192 ( \31470 , \31463 , \31469 );
and \U$23194 ( \31471 , \31470 , 1'b1 );
or \U$23196 ( \31472 , \31471 , 1'b0 );
buf \U$23197 ( \31473 , \31472 );
_DC r23e64_GF_IsGateDCbyConstraint ( \31474_nR23e64 , \31473 , \21944 );
buf \U$23198 ( \31475 , \31474_nR23e64 );
not \U$23199 ( \31476 , \31180 );
and \U$23200 ( \31477 , RIe481b08_6315, \31476 );
not \U$23201 ( \31478 , RIe481b08_6315);
or \U$23202 ( \31479 , \31478 , \30937 );
nand \U$23203 ( \31480 , \28177 , \30971 );
nand \U$23204 ( \31481 , \28180 , \30957 );
nand \U$23205 ( \31482 , \31479 , \31480 , \31481 );
and \U$23206 ( \31483 , \31482 , \31180 );
or \U$23207 ( \31484 , \31477 , \31483 );
and \U$23209 ( \31485 , \31484 , 1'b1 );
or \U$23211 ( \31486 , \31485 , 1'b0 );
buf \U$23212 ( \31487 , \31486 );
_DC r23e68_GF_IsGateDCbyConstraint ( \31488_nR23e68 , \31487 , \21944 );
buf \U$23213 ( \31489 , \31488_nR23e68 );
not \U$23214 ( \31490 , \29571 );
and \U$23215 ( \31491 , RIe482300_6316, \31490 );
not \U$23216 ( \31492 , RIe482300_6316);
or \U$23217 ( \31493 , \31492 , \30937 );
nand \U$23218 ( \31494 , \28196 , \30905 );
nand \U$23219 ( \31495 , \28199 , \30987 );
nand \U$23220 ( \31496 , \31493 , \31494 , \31495 );
and \U$23221 ( \31497 , \31496 , \29571 );
or \U$23222 ( \31498 , \31491 , \31497 );
and \U$23224 ( \31499 , \31498 , 1'b1 );
or \U$23226 ( \31500 , \31499 , 1'b0 );
buf \U$23227 ( \31501 , \31500 );
_DC r23e6a_GF_IsGateDCbyConstraint ( \31502_nR23e6a , \31501 , \21944 );
buf \U$23228 ( \31503 , \31502_nR23e6a );
not \U$23229 ( \31504 , \31335 );
and \U$23230 ( \31505 , RIe482af8_6317, \31504 );
not \U$23231 ( \31506 , RIe482af8_6317);
or \U$23232 ( \31507 , \31506 , \30921 );
nand \U$23233 ( \31508 , \28215 , \30971 );
nand \U$23234 ( \31509 , \28218 , \30908 );
nand \U$23235 ( \31510 , \31507 , \31508 , \31509 );
and \U$23236 ( \31511 , \31510 , \31335 );
or \U$23237 ( \31512 , \31505 , \31511 );
and \U$23239 ( \31513 , \31512 , 1'b1 );
or \U$23241 ( \31514 , \31513 , 1'b0 );
buf \U$23242 ( \31515 , \31514 );
_DC r23e6c_GF_IsGateDCbyConstraint ( \31516_nR23e6c , \31515 , \21944 );
buf \U$23243 ( \31517 , \31516_nR23e6c );
not \U$23244 ( \31518 , \31180 );
and \U$23245 ( \31519 , RIe4832f0_6318, \31518 );
not \U$23246 ( \31520 , RIe4832f0_6318);
or \U$23247 ( \31521 , \31520 , \30902 );
nand \U$23248 ( \31522 , \28235 , \30923 );
nand \U$23249 ( \31523 , \28237 , \30908 );
nand \U$23250 ( \31524 , \31521 , \31522 , \31523 );
and \U$23251 ( \31525 , \31524 , \31180 );
or \U$23252 ( \31526 , \31519 , \31525 );
and \U$23254 ( \31527 , \31526 , 1'b1 );
or \U$23256 ( \31528 , \31527 , 1'b0 );
buf \U$23257 ( \31529 , \31528 );
_DC r23e6e_GF_IsGateDCbyConstraint ( \31530_nR23e6e , \31529 , \21944 );
buf \U$23258 ( \31531 , \31530_nR23e6e );
not \U$23259 ( \31532 , \29571 );
and \U$23260 ( \31533 , RIe483ae8_6319, \31532 );
not \U$23261 ( \31534 , RIe483ae8_6319);
or \U$23262 ( \31535 , \31534 , \31042 );
nand \U$23263 ( \31536 , \28254 , \30905 );
nand \U$23264 ( \31537 , \28257 , \30957 );
nand \U$23265 ( \31538 , \31535 , \31536 , \31537 );
and \U$23266 ( \31539 , \31538 , \29571 );
or \U$23267 ( \31540 , \31533 , \31539 );
and \U$23269 ( \31541 , \31540 , 1'b1 );
or \U$23271 ( \31542 , \31541 , 1'b0 );
buf \U$23272 ( \31543 , \31542 );
_DC r23e70_GF_IsGateDCbyConstraint ( \31544_nR23e70 , \31543 , \21944 );
buf \U$23273 ( \31545 , \31544_nR23e70 );
not \U$23274 ( \31546 , \31335 );
and \U$23275 ( \31547 , RIe4842e0_6320, \31546 );
not \U$23276 ( \31548 , RIe4842e0_6320);
or \U$23277 ( \31549 , \31548 , \30921 );
nand \U$23278 ( \31550 , \28273 , \30955 );
nand \U$23279 ( \31551 , \28276 , \30940 );
nand \U$23280 ( \31552 , \31549 , \31550 , \31551 );
and \U$23281 ( \31553 , \31552 , \31335 );
or \U$23282 ( \31554 , \31547 , \31553 );
and \U$23284 ( \31555 , \31554 , 1'b1 );
or \U$23286 ( \31556 , \31555 , 1'b0 );
buf \U$23287 ( \31557 , \31556 );
_DC r23e72_GF_IsGateDCbyConstraint ( \31558_nR23e72 , \31557 , \21944 );
buf \U$23288 ( \31559 , \31558_nR23e72 );
not \U$23289 ( \31560 , \31180 );
and \U$23290 ( \31561 , RIe484ad8_6321, \31560 );
not \U$23291 ( \31562 , RIe484ad8_6321);
or \U$23292 ( \31563 , \31562 , \30953 );
nand \U$23293 ( \31564 , \28292 , \30955 );
nand \U$23294 ( \31565 , \28295 , \30940 );
nand \U$23295 ( \31566 , \31563 , \31564 , \31565 );
and \U$23296 ( \31567 , \31566 , \31180 );
or \U$23297 ( \31568 , \31561 , \31567 );
and \U$23299 ( \31569 , \31568 , 1'b1 );
or \U$23301 ( \31570 , \31569 , 1'b0 );
buf \U$23302 ( \31571 , \31570 );
_DC r23e74_GF_IsGateDCbyConstraint ( \31572_nR23e74 , \31571 , \21944 );
buf \U$23303 ( \31573 , \31572_nR23e74 );
not \U$23304 ( \31574 , \29571 );
and \U$23305 ( \31575 , RIe4852d0_6322, \31574 );
not \U$23306 ( \31576 , RIe4852d0_6322);
or \U$23307 ( \31577 , \31576 , \30937 );
nand \U$23308 ( \31578 , \28312 , \30955 );
nand \U$23309 ( \31579 , \28314 , \30908 );
nand \U$23310 ( \31580 , \31577 , \31578 , \31579 );
and \U$23311 ( \31581 , \31580 , \29571 );
or \U$23312 ( \31582 , \31575 , \31581 );
and \U$23314 ( \31583 , \31582 , 1'b1 );
or \U$23316 ( \31584 , \31583 , 1'b0 );
buf \U$23317 ( \31585 , \31584 );
_DC r23e76_GF_IsGateDCbyConstraint ( \31586_nR23e76 , \31585 , \21944 );
buf \U$23318 ( \31587 , \31586_nR23e76 );
not \U$23319 ( \31588 , \31335 );
and \U$23320 ( \31589 , RIe485ac8_6323, \31588 );
not \U$23321 ( \31590 , RIe485ac8_6323);
or \U$23322 ( \31591 , \31590 , \30921 );
nand \U$23323 ( \31592 , \28330 , \30971 );
nand \U$23324 ( \31593 , \28333 , \30987 );
nand \U$23325 ( \31594 , \31591 , \31592 , \31593 );
and \U$23326 ( \31595 , \31594 , \31335 );
or \U$23327 ( \31596 , \31589 , \31595 );
and \U$23329 ( \31597 , \31596 , 1'b1 );
or \U$23331 ( \31598 , \31597 , 1'b0 );
buf \U$23332 ( \31599 , \31598 );
_DC r23e78_GF_IsGateDCbyConstraint ( \31600_nR23e78 , \31599 , \21944 );
buf \U$23333 ( \31601 , \31600_nR23e78 );
not \U$23334 ( \31602 , \31180 );
and \U$23335 ( \31603 , RIe4862c0_6324, \31602 );
not \U$23336 ( \31604 , RIe4862c0_6324);
or \U$23337 ( \31605 , \31604 , \30902 );
nand \U$23338 ( \31606 , \28349 , \30971 );
nand \U$23339 ( \31607 , \28352 , \30987 );
nand \U$23340 ( \31608 , \31605 , \31606 , \31607 );
and \U$23341 ( \31609 , \31608 , \31180 );
or \U$23342 ( \31610 , \31603 , \31609 );
and \U$23344 ( \31611 , \31610 , 1'b1 );
or \U$23346 ( \31612 , \31611 , 1'b0 );
buf \U$23347 ( \31613 , \31612 );
_DC r23e7a_GF_IsGateDCbyConstraint ( \31614_nR23e7a , \31613 , \21944 );
buf \U$23348 ( \31615 , \31614_nR23e7a );
not \U$23349 ( \31616 , \27458 );
and \U$23350 ( \31617 , RIe486ab8_6325, \31616 );
not \U$23351 ( \31618 , RIe486ab8_6325);
or \U$23352 ( \31619 , \31618 , \31042 );
nand \U$23353 ( \31620 , \28369 , \30971 );
nand \U$23354 ( \31621 , \28372 , \30957 );
nand \U$23355 ( \31622 , \31619 , \31620 , \31621 );
and \U$23356 ( \31623 , \31622 , \27458 );
or \U$23357 ( \31624 , \31617 , \31623 );
and \U$23359 ( \31625 , \31624 , 1'b1 );
or \U$23361 ( \31626 , \31625 , 1'b0 );
buf \U$23362 ( \31627 , \31626 );
_DC r23e7e_GF_IsGateDCbyConstraint ( \31628_nR23e7e , \31627 , \21944 );
buf \U$23363 ( \31629 , \31628_nR23e7e );
not \U$23364 ( \31630 , \31335 );
and \U$23365 ( \31631 , RIe4872b0_6326, \31630 );
not \U$23366 ( \31632 , RIe4872b0_6326);
or \U$23367 ( \31633 , \31632 , \30953 );
nand \U$23368 ( \31634 , \28389 , \30955 );
nand \U$23369 ( \31635 , \28392 , \30957 );
nand \U$23370 ( \31636 , \31633 , \31634 , \31635 );
and \U$23371 ( \31637 , \31636 , \31335 );
or \U$23372 ( \31638 , \31631 , \31637 );
and \U$23374 ( \31639 , \31638 , 1'b1 );
or \U$23376 ( \31640 , \31639 , 1'b0 );
buf \U$23377 ( \31641 , \31640 );
_DC r23e80_GF_IsGateDCbyConstraint ( \31642_nR23e80 , \31641 , \21944 );
buf \U$23378 ( \31643 , \31642_nR23e80 );
not \U$23379 ( \31644 , \31180 );
and \U$23380 ( \31645 , RIe487aa8_6327, \31644 );
not \U$23381 ( \31646 , RIe487aa8_6327);
or \U$23382 ( \31647 , \31646 , \30937 );
nand \U$23383 ( \31648 , \28409 , \30905 );
nand \U$23384 ( \31649 , \28412 , \30987 );
nand \U$23385 ( \31650 , \31647 , \31648 , \31649 );
and \U$23386 ( \31651 , \31650 , \31180 );
or \U$23387 ( \31652 , \31645 , \31651 );
and \U$23389 ( \31653 , \31652 , 1'b1 );
or \U$23391 ( \31654 , \31653 , 1'b0 );
buf \U$23392 ( \31655 , \31654 );
_DC r23e82_GF_IsGateDCbyConstraint ( \31656_nR23e82 , \31655 , \21944 );
buf \U$23393 ( \31657 , \31656_nR23e82 );
not \U$23394 ( \31658 , \27364 );
and \U$23395 ( \31659 , RIe4882a0_6328, \31658 );
not \U$23396 ( \31660 , RIe4882a0_6328);
or \U$23397 ( \31661 , \31660 , \30921 );
nand \U$23398 ( \31662 , \28429 , \30971 );
nand \U$23399 ( \31663 , \28432 , \30908 );
nand \U$23400 ( \31664 , \31661 , \31662 , \31663 );
and \U$23401 ( \31665 , \31664 , \27364 );
or \U$23402 ( \31666 , \31659 , \31665 );
and \U$23404 ( \31667 , \31666 , 1'b1 );
or \U$23406 ( \31668 , \31667 , 1'b0 );
buf \U$23407 ( \31669 , \31668 );
_DC r23e84_GF_IsGateDCbyConstraint ( \31670_nR23e84 , \31669 , \21944 );
buf \U$23408 ( \31671 , \31670_nR23e84 );
not \U$23409 ( \31672 , \31335 );
and \U$23410 ( \31673 , RIe488a98_6329, \31672 );
not \U$23411 ( \31674 , RIe488a98_6329);
or \U$23412 ( \31675 , \31674 , \31042 );
nand \U$23413 ( \31676 , \28449 , \30955 );
nand \U$23414 ( \31677 , \28452 , \30908 );
nand \U$23415 ( \31678 , \31675 , \31676 , \31677 );
and \U$23416 ( \31679 , \31678 , \31335 );
or \U$23417 ( \31680 , \31673 , \31679 );
and \U$23419 ( \31681 , \31680 , 1'b1 );
or \U$23421 ( \31682 , \31681 , 1'b0 );
buf \U$23422 ( \31683 , \31682 );
_DC r23e86_GF_IsGateDCbyConstraint ( \31684_nR23e86 , \31683 , \21944 );
buf \U$23423 ( \31685 , \31684_nR23e86 );
not \U$23424 ( \31686 , \27459 );
and \U$23425 ( \31687 , RIe489290_6330, \31686 );
not \U$23426 ( \31688 , RIe489290_6330);
or \U$23427 ( \31689 , \31688 , \30902 );
nand \U$23428 ( \31690 , \28468 , \30905 );
nand \U$23429 ( \31691 , \28471 , \30957 );
nand \U$23430 ( \31692 , \31689 , \31690 , \31691 );
and \U$23431 ( \31693 , \31692 , \27459 );
or \U$23432 ( \31694 , \31687 , \31693 );
and \U$23434 ( \31695 , \31694 , 1'b1 );
or \U$23436 ( \31696 , \31695 , 1'b0 );
buf \U$23437 ( \31697 , \31696 );
_DC r23e88_GF_IsGateDCbyConstraint ( \31698_nR23e88 , \31697 , \21944 );
buf \U$23438 ( \31699 , \31698_nR23e88 );
not \U$23439 ( \31700 , \29329 );
and \U$23440 ( \31701 , RIe489a88_6331, \31700 );
not \U$23441 ( \31702 , RIe489a88_6331);
or \U$23442 ( \31703 , \31702 , \31042 );
nand \U$23443 ( \31704 , \28488 , \30955 );
nand \U$23444 ( \31705 , \28490 , \30940 );
nand \U$23445 ( \31706 , \31703 , \31704 , \31705 );
and \U$23446 ( \31707 , \31706 , \29329 );
or \U$23447 ( \31708 , \31701 , \31707 );
and \U$23449 ( \31709 , \31708 , 1'b1 );
or \U$23451 ( \31710 , \31709 , 1'b0 );
buf \U$23452 ( \31711 , \31710 );
_DC r23e8a_GF_IsGateDCbyConstraint ( \31712_nR23e8a , \31711 , \21944 );
buf \U$23453 ( \31713 , \31712_nR23e8a );
not \U$23454 ( \31714 , \31335 );
and \U$23455 ( \31715 , RIe48a280_6332, \31714 );
not \U$23456 ( \31716 , RIe48a280_6332);
or \U$23457 ( \31717 , \31716 , \30953 );
nand \U$23458 ( \31718 , \28507 , \30923 );
nand \U$23459 ( \31719 , \28510 , \30940 );
nand \U$23460 ( \31720 , \31717 , \31718 , \31719 );
and \U$23461 ( \31721 , \31720 , \31335 );
or \U$23462 ( \31722 , \31715 , \31721 );
and \U$23464 ( \31723 , \31722 , 1'b1 );
or \U$23466 ( \31724 , \31723 , 1'b0 );
buf \U$23467 ( \31725 , \31724 );
_DC r23e8c_GF_IsGateDCbyConstraint ( \31726_nR23e8c , \31725 , \21944 );
buf \U$23468 ( \31727 , \31726_nR23e8c );
not \U$23469 ( \31728 , \27459 );
and \U$23470 ( \31729 , RIe48aa78_6333, \31728 );
not \U$23471 ( \31730 , RIe48aa78_6333);
or \U$23472 ( \31731 , \31730 , \30937 );
nand \U$23473 ( \31732 , \28526 , \30905 );
nand \U$23474 ( \31733 , \28529 , \30908 );
nand \U$23475 ( \31734 , \31731 , \31732 , \31733 );
and \U$23476 ( \31735 , \31734 , \27459 );
or \U$23477 ( \31736 , \31729 , \31735 );
and \U$23479 ( \31737 , \31736 , 1'b1 );
or \U$23481 ( \31738 , \31737 , 1'b0 );
buf \U$23482 ( \31739 , \31738 );
_DC r23e8e_GF_IsGateDCbyConstraint ( \31740_nR23e8e , \31739 , \21944 );
buf \U$23483 ( \31741 , \31740_nR23e8e );
not \U$23484 ( \31742 , \27364 );
and \U$23485 ( \31743 , RIe48b270_6334, \31742 );
not \U$23486 ( \31744 , RIe48b270_6334);
or \U$23487 ( \31745 , \31744 , \30953 );
nand \U$23488 ( \31746 , \28548 , \30971 );
nand \U$23489 ( \31747 , \28551 , \30987 );
nand \U$23490 ( \31748 , \31745 , \31746 , \31747 );
and \U$23491 ( \31749 , \31748 , \27364 );
or \U$23492 ( \31750 , \31743 , \31749 );
and \U$23494 ( \31751 , \31750 , 1'b1 );
or \U$23496 ( \31752 , \31751 , 1'b0 );
buf \U$23497 ( \31753 , \31752 );
_DC r23e90_GF_IsGateDCbyConstraint ( \31754_nR23e90 , \31753 , \21944 );
buf \U$23498 ( \31755 , \31754_nR23e90 );
not \U$23499 ( \31756 , \31335 );
and \U$23500 ( \31757 , RIe48ba68_6335, \31756 );
not \U$23501 ( \31758 , RIe48ba68_6335);
or \U$23502 ( \31759 , \31758 , \30902 );
nand \U$23503 ( \31760 , \28569 , \30971 );
nand \U$23504 ( \31761 , \28571 , \30940 );
nand \U$23505 ( \31762 , \31759 , \31760 , \31761 );
and \U$23506 ( \31763 , \31762 , \31335 );
or \U$23507 ( \31764 , \31757 , \31763 );
and \U$23509 ( \31765 , \31764 , 1'b1 );
or \U$23511 ( \31766 , \31765 , 1'b0 );
buf \U$23512 ( \31767 , \31766 );
_DC r23e94_GF_IsGateDCbyConstraint ( \31768_nR23e94 , \31767 , \21944 );
buf \U$23513 ( \31769 , \31768_nR23e94 );
not \U$23514 ( \31770 , \27459 );
and \U$23515 ( \31771 , RIe48c260_6336, \31770 );
not \U$23516 ( \31772 , RIe48c260_6336);
or \U$23517 ( \31773 , \31772 , \31042 );
nand \U$23518 ( \31774 , \28587 , \30905 );
nand \U$23519 ( \31775 , \28589 , \30957 );
nand \U$23520 ( \31776 , \31773 , \31774 , \31775 );
and \U$23521 ( \31777 , \31776 , \27459 );
or \U$23522 ( \31778 , \31771 , \31777 );
and \U$23524 ( \31779 , \31778 , 1'b1 );
or \U$23526 ( \31780 , \31779 , 1'b0 );
buf \U$23527 ( \31781 , \31780 );
_DC r23e96_GF_IsGateDCbyConstraint ( \31782_nR23e96 , \31781 , \21944 );
buf \U$23528 ( \31783 , \31782_nR23e96 );
not \U$23529 ( \31784 , \29329 );
and \U$23530 ( \31785 , RIe48ca58_6337, \31784 );
not \U$23531 ( \31786 , RIe48ca58_6337);
or \U$23532 ( \31787 , \31786 , \30953 );
nand \U$23533 ( \31788 , \28606 , \30923 );
nand \U$23534 ( \31789 , \28608 , \30957 );
nand \U$23535 ( \31790 , \31787 , \31788 , \31789 );
and \U$23536 ( \31791 , \31790 , \29329 );
or \U$23537 ( \31792 , \31785 , \31791 );
and \U$23539 ( \31793 , \31792 , 1'b1 );
or \U$23541 ( \31794 , \31793 , 1'b0 );
buf \U$23542 ( \31795 , \31794 );
_DC r23e98_GF_IsGateDCbyConstraint ( \31796_nR23e98 , \31795 , \21944 );
buf \U$23543 ( \31797 , \31796_nR23e98 );
not \U$23544 ( \31798 , \31335 );
and \U$23545 ( \31799 , RIe48d250_6338, \31798 );
not \U$23546 ( \31800 , RIe48d250_6338);
or \U$23547 ( \31801 , \31800 , \30937 );
nand \U$23548 ( \31802 , \28624 , \30905 );
nand \U$23549 ( \31803 , \28626 , \30987 );
nand \U$23550 ( \31804 , \31801 , \31802 , \31803 );
and \U$23551 ( \31805 , \31804 , \31335 );
or \U$23552 ( \31806 , \31799 , \31805 );
and \U$23554 ( \31807 , \31806 , 1'b1 );
or \U$23556 ( \31808 , \31807 , 1'b0 );
buf \U$23557 ( \31809 , \31808 );
_DC r23e9a_GF_IsGateDCbyConstraint ( \31810_nR23e9a , \31809 , \21944 );
buf \U$23558 ( \31811 , \31810_nR23e9a );
nor \U$23559 ( \31812 , \27354 , \27385 );
not \U$23560 ( \31813 , \31812 );
not \U$23561 ( \31814 , \31813 );
not \U$23562 ( \31815 , \31814 );
and \U$23563 ( \31816 , RIe3cd190_6051, \31815 );
not \U$23564 ( \31817 , RIe3cd190_6051);
not \U$23565 ( \31818 , \31817 );
not \U$23566 ( \31819 , \27376 );
and \U$23567 ( \31820 , \31818 , \31819 );
buf \U$23568 ( \31821 , \26668 );
and \U$23569 ( \31822 , \31821 , \27376 );
or \U$23570 ( \31823 , \31820 , \31822 );
and \U$23571 ( \31824 , \31823 , \31814 );
or \U$23572 ( \31825 , \31816 , \31824 );
and \U$23574 ( \31826 , \31825 , 1'b1 );
or \U$23576 ( \31827 , \31826 , 1'b0 );
buf \U$23577 ( \31828 , \31827 );
_DC r23c64_GF_IsGateDCbyConstraint ( \31829_nR23c64 , \31828 , \21944 );
buf \U$23578 ( \31830 , \31829_nR23c64 );
not \U$23579 ( \31831 , \31813 );
not \U$23580 ( \31832 , \31831 );
and \U$23581 ( \31833 , RIe3cc3f8_6052, \31832 );
not \U$23582 ( \31834 , RIe3cc3f8_6052);
not \U$23583 ( \31835 , \31834 );
not \U$23584 ( \31836 , \27376 );
and \U$23585 ( \31837 , \31835 , \31836 );
buf \U$23586 ( \31838 , \26686 );
and \U$23587 ( \31839 , \31838 , \27376 );
or \U$23588 ( \31840 , \31837 , \31839 );
and \U$23589 ( \31841 , \31840 , \31831 );
or \U$23590 ( \31842 , \31833 , \31841 );
and \U$23592 ( \31843 , \31842 , 1'b1 );
or \U$23594 ( \31844 , \31843 , 1'b0 );
buf \U$23595 ( \31845 , \31844 );
_DC r23c66_GF_IsGateDCbyConstraint ( \31846_nR23c66 , \31845 , \21944 );
buf \U$23596 ( \31847 , \31846_nR23c66 );
not \U$23597 ( \31848 , \31814 );
and \U$23598 ( \31849 , RIe3cb750_6053, \31848 );
not \U$23599 ( \31850 , RIe3cb750_6053);
not \U$23600 ( \31851 , \31850 );
not \U$23601 ( \31852 , \27376 );
and \U$23602 ( \31853 , \31851 , \31852 );
buf \U$23603 ( \31854 , RIb86fd58_75);
and \U$23604 ( \31855 , \31854 , \27376 );
or \U$23605 ( \31856 , \31853 , \31855 );
and \U$23606 ( \31857 , \31856 , \31814 );
or \U$23607 ( \31858 , \31849 , \31857 );
and \U$23609 ( \31859 , \31858 , 1'b1 );
or \U$23611 ( \31860 , \31859 , 1'b0 );
buf \U$23612 ( \31861 , \31860 );
_DC r23c68_GF_IsGateDCbyConstraint ( \31862_nR23c68 , \31861 , \21944 );
buf \U$23613 ( \31863 , \31862_nR23c68 );
not \U$23614 ( \31864 , \31814 );
and \U$23615 ( \31865 , RIe3ca9b8_6054, \31864 );
not \U$23616 ( \31866 , RIe3ca9b8_6054);
not \U$23617 ( \31867 , \31866 );
not \U$23618 ( \31868 , \27376 );
and \U$23619 ( \31869 , \31867 , \31868 );
buf \U$23620 ( \31870 , \26720 );
and \U$23621 ( \31871 , \31870 , \27376 );
or \U$23622 ( \31872 , \31869 , \31871 );
and \U$23623 ( \31873 , \31872 , \31814 );
or \U$23624 ( \31874 , \31865 , \31873 );
and \U$23626 ( \31875 , \31874 , 1'b1 );
or \U$23628 ( \31876 , \31875 , 1'b0 );
buf \U$23629 ( \31877 , \31876 );
_DC r23c6a_GF_IsGateDCbyConstraint ( \31878_nR23c6a , \31877 , \21944 );
buf \U$23630 ( \31879 , \31878_nR23c6a );
not \U$23631 ( \31880 , \31814 );
and \U$23632 ( \31881 , RIe3c9e00_6055, \31880 );
not \U$23633 ( \31882 , RIe3c9e00_6055);
not \U$23634 ( \31883 , \31882 );
not \U$23635 ( \31884 , \27376 );
and \U$23636 ( \31885 , \31883 , \31884 );
buf \U$23637 ( \31886 , \26737 );
and \U$23638 ( \31887 , \31886 , \27376 );
or \U$23639 ( \31888 , \31885 , \31887 );
and \U$23640 ( \31889 , \31888 , \31814 );
or \U$23641 ( \31890 , \31881 , \31889 );
and \U$23643 ( \31891 , \31890 , 1'b1 );
or \U$23645 ( \31892 , \31891 , 1'b0 );
buf \U$23646 ( \31893 , \31892 );
_DC r23c6c_GF_IsGateDCbyConstraint ( \31894_nR23c6c , \31893 , \21944 );
buf \U$23647 ( \31895 , \31894_nR23c6c );
not \U$23648 ( \31896 , \31831 );
and \U$23649 ( \31897 , RIe3c9248_6056, \31896 );
not \U$23650 ( \31898 , RIe3c9248_6056);
not \U$23651 ( \31899 , \31898 );
not \U$23652 ( \31900 , \27376 );
and \U$23653 ( \31901 , \31899 , \31900 );
buf \U$23654 ( \31902 , \26754 );
and \U$23655 ( \31903 , \31902 , \27376 );
or \U$23656 ( \31904 , \31901 , \31903 );
and \U$23657 ( \31905 , \31904 , \31831 );
or \U$23658 ( \31906 , \31897 , \31905 );
and \U$23660 ( \31907 , \31906 , 1'b1 );
or \U$23662 ( \31908 , \31907 , 1'b0 );
buf \U$23663 ( \31909 , \31908 );
_DC r23c6e_GF_IsGateDCbyConstraint ( \31910_nR23c6e , \31909 , \21944 );
buf \U$23664 ( \31911 , \31910_nR23c6e );
not \U$23665 ( \31912 , \31814 );
and \U$23666 ( \31913 , RIe3c8708_6057, \31912 );
not \U$23667 ( \31914 , RIe3c8708_6057);
not \U$23668 ( \31915 , \31914 );
not \U$23669 ( \31916 , \27376 );
and \U$23670 ( \31917 , \31915 , \31916 );
buf \U$23671 ( \31918 , \26771 );
and \U$23672 ( \31919 , \31918 , \27376 );
or \U$23673 ( \31920 , \31917 , \31919 );
and \U$23674 ( \31921 , \31920 , \31814 );
or \U$23675 ( \31922 , \31913 , \31921 );
and \U$23677 ( \31923 , \31922 , 1'b1 );
or \U$23679 ( \31924 , \31923 , 1'b0 );
buf \U$23680 ( \31925 , \31924 );
_DC r23c70_GF_IsGateDCbyConstraint ( \31926_nR23c70 , \31925 , \21944 );
buf \U$23681 ( \31927 , \31926_nR23c70 );
not \U$23682 ( \31928 , \31831 );
and \U$23683 ( \31929 , RIe3c7bc8_6058, \31928 );
not \U$23684 ( \31930 , RIe3c7bc8_6058);
not \U$23685 ( \31931 , \31930 );
not \U$23686 ( \31932 , \27376 );
and \U$23687 ( \31933 , \31931 , \31932 );
buf \U$23688 ( \31934 , \26788 );
and \U$23689 ( \31935 , \31934 , \27376 );
or \U$23690 ( \31936 , \31933 , \31935 );
and \U$23691 ( \31937 , \31936 , \31831 );
or \U$23692 ( \31938 , \31929 , \31937 );
and \U$23694 ( \31939 , \31938 , 1'b1 );
or \U$23696 ( \31940 , \31939 , 1'b0 );
buf \U$23697 ( \31941 , \31940 );
_DC r23c72_GF_IsGateDCbyConstraint ( \31942_nR23c72 , \31941 , \21944 );
buf \U$23698 ( \31943 , \31942_nR23c72 );
not \U$23699 ( \31944 , \31814 );
and \U$23700 ( \31945 , RIe3c7100_6059, \31944 );
not \U$23701 ( \31946 , RIe3c7100_6059);
not \U$23702 ( \31947 , \31946 );
not \U$23703 ( \31948 , \28646 );
and \U$23704 ( \31949 , \31947 , \31948 );
and \U$23705 ( \31950 , \31821 , \28646 );
or \U$23706 ( \31951 , \31949 , \31950 );
and \U$23707 ( \31952 , \31951 , \31814 );
or \U$23708 ( \31953 , \31945 , \31952 );
and \U$23710 ( \31954 , \31953 , 1'b1 );
or \U$23712 ( \31955 , \31954 , 1'b0 );
buf \U$23713 ( \31956 , \31955 );
_DC r23c74_GF_IsGateDCbyConstraint ( \31957_nR23c74 , \31956 , \21944 );
buf \U$23714 ( \31958 , \31957_nR23c74 );
not \U$23715 ( \31959 , \31831 );
and \U$23716 ( \31960 , RIe3c6638_6060, \31959 );
not \U$23717 ( \31961 , RIe3c6638_6060);
not \U$23718 ( \31962 , \31961 );
not \U$23719 ( \31963 , \28646 );
and \U$23720 ( \31964 , \31962 , \31963 );
and \U$23721 ( \31965 , \31838 , \28646 );
or \U$23722 ( \31966 , \31964 , \31965 );
and \U$23723 ( \31967 , \31966 , \31831 );
or \U$23724 ( \31968 , \31960 , \31967 );
and \U$23726 ( \31969 , \31968 , 1'b1 );
or \U$23728 ( \31970 , \31969 , 1'b0 );
buf \U$23729 ( \31971 , \31970 );
_DC r23c76_GF_IsGateDCbyConstraint ( \31972_nR23c76 , \31971 , \21944 );
buf \U$23730 ( \31973 , \31972_nR23c76 );
not \U$23731 ( \31974 , \31814 );
and \U$23732 ( \31975 , RIe3c5af8_6061, \31974 );
not \U$23733 ( \31976 , RIe3c5af8_6061);
not \U$23734 ( \31977 , \31976 );
not \U$23735 ( \31978 , \28646 );
and \U$23736 ( \31979 , \31977 , \31978 );
and \U$23737 ( \31980 , \31854 , \28646 );
or \U$23738 ( \31981 , \31979 , \31980 );
and \U$23739 ( \31982 , \31981 , \31814 );
or \U$23740 ( \31983 , \31975 , \31982 );
and \U$23742 ( \31984 , \31983 , 1'b1 );
or \U$23744 ( \31985 , \31984 , 1'b0 );
buf \U$23745 ( \31986 , \31985 );
_DC r23c78_GF_IsGateDCbyConstraint ( \31987_nR23c78 , \31986 , \21944 );
buf \U$23746 ( \31988 , \31987_nR23c78 );
not \U$23747 ( \31989 , \31831 );
and \U$23748 ( \31990 , RIe3c4ec8_6062, \31989 );
not \U$23749 ( \31991 , RIe3c4ec8_6062);
not \U$23750 ( \31992 , \31991 );
not \U$23751 ( \31993 , \28646 );
and \U$23752 ( \31994 , \31992 , \31993 );
and \U$23753 ( \31995 , \31870 , \28646 );
or \U$23754 ( \31996 , \31994 , \31995 );
and \U$23755 ( \31997 , \31996 , \31831 );
or \U$23756 ( \31998 , \31990 , \31997 );
and \U$23758 ( \31999 , \31998 , 1'b1 );
or \U$23760 ( \32000 , \31999 , 1'b0 );
buf \U$23761 ( \32001 , \32000 );
_DC r23c7a_GF_IsGateDCbyConstraint ( \32002_nR23c7a , \32001 , \21944 );
buf \U$23762 ( \32003 , \32002_nR23c7a );
not \U$23763 ( \32004 , \31814 );
and \U$23764 ( \32005 , RIe3c4130_6063, \32004 );
not \U$23765 ( \32006 , RIe3c4130_6063);
not \U$23766 ( \32007 , \32006 );
not \U$23767 ( \32008 , \28646 );
and \U$23768 ( \32009 , \32007 , \32008 );
and \U$23769 ( \32010 , \31886 , \28646 );
or \U$23770 ( \32011 , \32009 , \32010 );
and \U$23771 ( \32012 , \32011 , \31814 );
or \U$23772 ( \32013 , \32005 , \32012 );
and \U$23774 ( \32014 , \32013 , 1'b1 );
or \U$23776 ( \32015 , \32014 , 1'b0 );
buf \U$23777 ( \32016 , \32015 );
_DC r23c7c_GF_IsGateDCbyConstraint ( \32017_nR23c7c , \32016 , \21944 );
buf \U$23778 ( \32018 , \32017_nR23c7c );
not \U$23779 ( \32019 , \31831 );
and \U$23780 ( \32020 , RIe3c31b8_6064, \32019 );
not \U$23781 ( \32021 , RIe3c31b8_6064);
not \U$23782 ( \32022 , \32021 );
not \U$23783 ( \32023 , \28646 );
and \U$23784 ( \32024 , \32022 , \32023 );
and \U$23785 ( \32025 , \31902 , \28646 );
or \U$23786 ( \32026 , \32024 , \32025 );
and \U$23787 ( \32027 , \32026 , \31831 );
or \U$23788 ( \32028 , \32020 , \32027 );
and \U$23790 ( \32029 , \32028 , 1'b1 );
or \U$23792 ( \32030 , \32029 , 1'b0 );
buf \U$23793 ( \32031 , \32030 );
_DC r23c7e_GF_IsGateDCbyConstraint ( \32032_nR23c7e , \32031 , \21944 );
buf \U$23794 ( \32033 , \32032_nR23c7e );
not \U$23795 ( \32034 , \31814 );
and \U$23796 ( \32035 , RIe3c1bb0_6065, \32034 );
not \U$23797 ( \32036 , RIe3c1bb0_6065);
not \U$23798 ( \32037 , \32036 );
not \U$23799 ( \32038 , \28646 );
and \U$23800 ( \32039 , \32037 , \32038 );
and \U$23801 ( \32040 , \31918 , \28646 );
or \U$23802 ( \32041 , \32039 , \32040 );
and \U$23803 ( \32042 , \32041 , \31814 );
or \U$23804 ( \32043 , \32035 , \32042 );
and \U$23806 ( \32044 , \32043 , 1'b1 );
or \U$23808 ( \32045 , \32044 , 1'b0 );
buf \U$23809 ( \32046 , \32045 );
_DC r23c80_GF_IsGateDCbyConstraint ( \32047_nR23c80 , \32046 , \21944 );
buf \U$23810 ( \32048 , \32047_nR23c80 );
not \U$23811 ( \32049 , \31831 );
and \U$23812 ( \32050 , RIe3c0a58_6066, \32049 );
not \U$23813 ( \32051 , RIe3c0a58_6066);
not \U$23814 ( \32052 , \32051 );
not \U$23815 ( \32053 , \28646 );
and \U$23816 ( \32054 , \32052 , \32053 );
and \U$23817 ( \32055 , \31934 , \28646 );
or \U$23818 ( \32056 , \32054 , \32055 );
and \U$23819 ( \32057 , \32056 , \31831 );
or \U$23820 ( \32058 , \32050 , \32057 );
and \U$23822 ( \32059 , \32058 , 1'b1 );
or \U$23824 ( \32060 , \32059 , 1'b0 );
buf \U$23825 ( \32061 , \32060 );
_DC r23c82_GF_IsGateDCbyConstraint ( \32062_nR23c82 , \32061 , \21944 );
buf \U$23826 ( \32063 , \32062_nR23c82 );
not \U$23827 ( \32064 , \31814 );
and \U$23828 ( \32065 , RIe3bf900_6067, \32064 );
not \U$23829 ( \32066 , RIe3bf900_6067);
not \U$23830 ( \32067 , \32066 );
not \U$23831 ( \32068 , \29796 );
and \U$23832 ( \32069 , \32067 , \32068 );
and \U$23833 ( \32070 , \31821 , \29796 );
or \U$23834 ( \32071 , \32069 , \32070 );
and \U$23835 ( \32072 , \32071 , \31814 );
or \U$23836 ( \32073 , \32065 , \32072 );
and \U$23838 ( \32074 , \32073 , 1'b1 );
or \U$23840 ( \32075 , \32074 , 1'b0 );
buf \U$23841 ( \32076 , \32075 );
_DC r23c84_GF_IsGateDCbyConstraint ( \32077_nR23c84 , \32076 , \21944 );
buf \U$23842 ( \32078 , \32077_nR23c84 );
not \U$23843 ( \32079 , \31814 );
and \U$23844 ( \32080 , RIe3be2f8_6068, \32079 );
not \U$23845 ( \32081 , RIe3be2f8_6068);
not \U$23846 ( \32082 , \32081 );
not \U$23847 ( \32083 , \29796 );
and \U$23848 ( \32084 , \32082 , \32083 );
and \U$23849 ( \32085 , \31838 , \29796 );
or \U$23850 ( \32086 , \32084 , \32085 );
and \U$23851 ( \32087 , \32086 , \31814 );
or \U$23852 ( \32088 , \32080 , \32087 );
and \U$23854 ( \32089 , \32088 , 1'b1 );
or \U$23856 ( \32090 , \32089 , 1'b0 );
buf \U$23857 ( \32091 , \32090 );
_DC r23c86_GF_IsGateDCbyConstraint ( \32092_nR23c86 , \32091 , \21944 );
buf \U$23858 ( \32093 , \32092_nR23c86 );
not \U$23859 ( \32094 , \31814 );
and \U$23860 ( \32095 , RIe3bd1a0_6069, \32094 );
not \U$23861 ( \32096 , RIe3bd1a0_6069);
not \U$23862 ( \32097 , \32096 );
not \U$23863 ( \32098 , \29796 );
and \U$23864 ( \32099 , \32097 , \32098 );
and \U$23865 ( \32100 , \31854 , \29796 );
or \U$23866 ( \32101 , \32099 , \32100 );
and \U$23867 ( \32102 , \32101 , \31814 );
or \U$23868 ( \32103 , \32095 , \32102 );
and \U$23870 ( \32104 , \32103 , 1'b1 );
or \U$23872 ( \32105 , \32104 , 1'b0 );
buf \U$23873 ( \32106 , \32105 );
_DC r23c88_GF_IsGateDCbyConstraint ( \32107_nR23c88 , \32106 , \21944 );
buf \U$23874 ( \32108 , \32107_nR23c88 );
not \U$23875 ( \32109 , \31814 );
and \U$23876 ( \32110 , RIe3bbb98_6070, \32109 );
not \U$23877 ( \32111 , RIe3bbb98_6070);
not \U$23878 ( \32112 , \32111 );
not \U$23879 ( \32113 , \29796 );
and \U$23880 ( \32114 , \32112 , \32113 );
and \U$23881 ( \32115 , \31870 , \29796 );
or \U$23882 ( \32116 , \32114 , \32115 );
and \U$23883 ( \32117 , \32116 , \31814 );
or \U$23884 ( \32118 , \32110 , \32117 );
and \U$23886 ( \32119 , \32118 , 1'b1 );
or \U$23888 ( \32120 , \32119 , 1'b0 );
buf \U$23889 ( \32121 , \32120 );
_DC r23c8a_GF_IsGateDCbyConstraint ( \32122_nR23c8a , \32121 , \21944 );
buf \U$23890 ( \32123 , \32122_nR23c8a );
not \U$23891 ( \32124 , \31814 );
and \U$23892 ( \32125 , RIe3baa40_6071, \32124 );
not \U$23893 ( \32126 , RIe3baa40_6071);
not \U$23894 ( \32127 , \32126 );
not \U$23895 ( \32128 , \29796 );
and \U$23896 ( \32129 , \32127 , \32128 );
and \U$23897 ( \32130 , \31886 , \29796 );
or \U$23898 ( \32131 , \32129 , \32130 );
and \U$23899 ( \32132 , \32131 , \31814 );
or \U$23900 ( \32133 , \32125 , \32132 );
and \U$23902 ( \32134 , \32133 , 1'b1 );
or \U$23904 ( \32135 , \32134 , 1'b0 );
buf \U$23905 ( \32136 , \32135 );
_DC r23c8c_GF_IsGateDCbyConstraint ( \32137_nR23c8c , \32136 , \21944 );
buf \U$23906 ( \32138 , \32137_nR23c8c );
not \U$23907 ( \32139 , \31814 );
and \U$23908 ( \32140 , RIe3b9438_6072, \32139 );
not \U$23909 ( \32141 , RIe3b9438_6072);
not \U$23910 ( \32142 , \32141 );
not \U$23911 ( \32143 , \29796 );
and \U$23912 ( \32144 , \32142 , \32143 );
and \U$23913 ( \32145 , \31902 , \29796 );
or \U$23914 ( \32146 , \32144 , \32145 );
and \U$23915 ( \32147 , \32146 , \31814 );
or \U$23916 ( \32148 , \32140 , \32147 );
and \U$23918 ( \32149 , \32148 , 1'b1 );
or \U$23920 ( \32150 , \32149 , 1'b0 );
buf \U$23921 ( \32151 , \32150 );
_DC r23c8e_GF_IsGateDCbyConstraint ( \32152_nR23c8e , \32151 , \21944 );
buf \U$23922 ( \32153 , \32152_nR23c8e );
not \U$23923 ( \32154 , \31814 );
and \U$23924 ( \32155 , RIe3b82e0_6073, \32154 );
not \U$23925 ( \32156 , RIe3b82e0_6073);
not \U$23926 ( \32157 , \32156 );
not \U$23927 ( \32158 , \29796 );
and \U$23928 ( \32159 , \32157 , \32158 );
and \U$23929 ( \32160 , \31918 , \29796 );
or \U$23930 ( \32161 , \32159 , \32160 );
and \U$23931 ( \32162 , \32161 , \31814 );
or \U$23932 ( \32163 , \32155 , \32162 );
and \U$23934 ( \32164 , \32163 , 1'b1 );
or \U$23936 ( \32165 , \32164 , 1'b0 );
buf \U$23937 ( \32166 , \32165 );
_DC r23c90_GF_IsGateDCbyConstraint ( \32167_nR23c90 , \32166 , \21944 );
buf \U$23938 ( \32168 , \32167_nR23c90 );
not \U$23939 ( \32169 , \31814 );
and \U$23940 ( \32170 , RIe3b7188_6074, \32169 );
not \U$23941 ( \32171 , RIe3b7188_6074);
not \U$23942 ( \32172 , \32171 );
not \U$23943 ( \32173 , \29796 );
and \U$23944 ( \32174 , \32172 , \32173 );
and \U$23945 ( \32175 , \31934 , \29796 );
or \U$23946 ( \32176 , \32174 , \32175 );
and \U$23947 ( \32177 , \32176 , \31814 );
or \U$23948 ( \32178 , \32170 , \32177 );
and \U$23950 ( \32179 , \32178 , 1'b1 );
or \U$23952 ( \32180 , \32179 , 1'b0 );
buf \U$23953 ( \32181 , \32180 );
_DC r23c92_GF_IsGateDCbyConstraint ( \32182_nR23c92 , \32181 , \21944 );
buf \U$23954 ( \32183 , \32182_nR23c92 );
not \U$23955 ( \32184 , \31814 );
and \U$23956 ( \32185 , RIe3b5b80_6075, \32184 );
not \U$23957 ( \32186 , RIe3b5b80_6075);
not \U$23958 ( \32187 , \32186 );
not \U$23959 ( \32188 , \30899 );
and \U$23960 ( \32189 , \32187 , \32188 );
and \U$23961 ( \32190 , \31821 , \30899 );
or \U$23962 ( \32191 , \32189 , \32190 );
and \U$23963 ( \32192 , \32191 , \31814 );
or \U$23964 ( \32193 , \32185 , \32192 );
and \U$23966 ( \32194 , \32193 , 1'b1 );
or \U$23968 ( \32195 , \32194 , 1'b0 );
buf \U$23969 ( \32196 , \32195 );
_DC r23c94_GF_IsGateDCbyConstraint ( \32197_nR23c94 , \32196 , \21944 );
buf \U$23970 ( \32198 , \32197_nR23c94 );
not \U$23971 ( \32199 , \31831 );
and \U$23972 ( \32200 , RIe3b4a28_6076, \32199 );
not \U$23973 ( \32201 , RIe3b4a28_6076);
not \U$23974 ( \32202 , \32201 );
not \U$23975 ( \32203 , \30899 );
and \U$23976 ( \32204 , \32202 , \32203 );
and \U$23977 ( \32205 , \31838 , \30899 );
or \U$23978 ( \32206 , \32204 , \32205 );
and \U$23979 ( \32207 , \32206 , \31831 );
or \U$23980 ( \32208 , \32200 , \32207 );
and \U$23982 ( \32209 , \32208 , 1'b1 );
or \U$23984 ( \32210 , \32209 , 1'b0 );
buf \U$23985 ( \32211 , \32210 );
_DC r23c96_GF_IsGateDCbyConstraint ( \32212_nR23c96 , \32211 , \21944 );
buf \U$23986 ( \32213 , \32212_nR23c96 );
not \U$23987 ( \32214 , \31831 );
and \U$23988 ( \32215 , RIe3b3420_6077, \32214 );
not \U$23989 ( \32216 , RIe3b3420_6077);
not \U$23990 ( \32217 , \32216 );
not \U$23991 ( \32218 , \30899 );
and \U$23992 ( \32219 , \32217 , \32218 );
and \U$23993 ( \32220 , \31854 , \30899 );
or \U$23994 ( \32221 , \32219 , \32220 );
and \U$23995 ( \32222 , \32221 , \31831 );
or \U$23996 ( \32223 , \32215 , \32222 );
and \U$23998 ( \32224 , \32223 , 1'b1 );
or \U$24000 ( \32225 , \32224 , 1'b0 );
buf \U$24001 ( \32226 , \32225 );
_DC r23c98_GF_IsGateDCbyConstraint ( \32227_nR23c98 , \32226 , \21944 );
buf \U$24002 ( \32228 , \32227_nR23c98 );
not \U$24003 ( \32229 , \31831 );
and \U$24004 ( \32230 , RIe3b22c8_6078, \32229 );
not \U$24005 ( \32231 , RIe3b22c8_6078);
not \U$24006 ( \32232 , \32231 );
not \U$24007 ( \32233 , \30899 );
and \U$24008 ( \32234 , \32232 , \32233 );
and \U$24009 ( \32235 , \31870 , \30899 );
or \U$24010 ( \32236 , \32234 , \32235 );
and \U$24011 ( \32237 , \32236 , \31831 );
or \U$24012 ( \32238 , \32230 , \32237 );
and \U$24014 ( \32239 , \32238 , 1'b1 );
or \U$24016 ( \32240 , \32239 , 1'b0 );
buf \U$24017 ( \32241 , \32240 );
_DC r23c9a_GF_IsGateDCbyConstraint ( \32242_nR23c9a , \32241 , \21944 );
buf \U$24018 ( \32243 , \32242_nR23c9a );
not \U$24019 ( \32244 , \31831 );
and \U$24020 ( \32245 , RIe3b0cc0_6079, \32244 );
not \U$24021 ( \32246 , RIe3b0cc0_6079);
not \U$24022 ( \32247 , \32246 );
not \U$24023 ( \32248 , \30899 );
and \U$24024 ( \32249 , \32247 , \32248 );
and \U$24025 ( \32250 , \31886 , \30899 );
or \U$24026 ( \32251 , \32249 , \32250 );
and \U$24027 ( \32252 , \32251 , \31831 );
or \U$24028 ( \32253 , \32245 , \32252 );
and \U$24030 ( \32254 , \32253 , 1'b1 );
or \U$24032 ( \32255 , \32254 , 1'b0 );
buf \U$24033 ( \32256 , \32255 );
_DC r23c9c_GF_IsGateDCbyConstraint ( \32257_nR23c9c , \32256 , \21944 );
buf \U$24034 ( \32258 , \32257_nR23c9c );
not \U$24035 ( \32259 , \31831 );
and \U$24036 ( \32260 , RIe3afb68_6080, \32259 );
not \U$24037 ( \32261 , RIe3afb68_6080);
not \U$24038 ( \32262 , \32261 );
not \U$24039 ( \32263 , \30899 );
and \U$24040 ( \32264 , \32262 , \32263 );
and \U$24041 ( \32265 , \31902 , \30899 );
or \U$24042 ( \32266 , \32264 , \32265 );
and \U$24043 ( \32267 , \32266 , \31831 );
or \U$24044 ( \32268 , \32260 , \32267 );
and \U$24046 ( \32269 , \32268 , 1'b1 );
or \U$24048 ( \32270 , \32269 , 1'b0 );
buf \U$24049 ( \32271 , \32270 );
_DC r23c9e_GF_IsGateDCbyConstraint ( \32272_nR23c9e , \32271 , \21944 );
buf \U$24050 ( \32273 , \32272_nR23c9e );
not \U$24051 ( \32274 , \31831 );
and \U$24052 ( \32275 , RIe3aea10_6081, \32274 );
not \U$24053 ( \32276 , RIe3aea10_6081);
not \U$24054 ( \32277 , \32276 );
not \U$24055 ( \32278 , \30899 );
and \U$24056 ( \32279 , \32277 , \32278 );
and \U$24057 ( \32280 , \31918 , \30899 );
or \U$24058 ( \32281 , \32279 , \32280 );
and \U$24059 ( \32282 , \32281 , \31831 );
or \U$24060 ( \32283 , \32275 , \32282 );
and \U$24062 ( \32284 , \32283 , 1'b1 );
or \U$24064 ( \32285 , \32284 , 1'b0 );
buf \U$24065 ( \32286 , \32285 );
_DC r23ca0_GF_IsGateDCbyConstraint ( \32287_nR23ca0 , \32286 , \21944 );
buf \U$24066 ( \32288 , \32287_nR23ca0 );
not \U$24067 ( \32289 , \31814 );
and \U$24068 ( \32290 , RIe3ad408_6082, \32289 );
not \U$24069 ( \32291 , RIe3ad408_6082);
not \U$24070 ( \32292 , \32291 );
not \U$24071 ( \32293 , \30899 );
and \U$24072 ( \32294 , \32292 , \32293 );
and \U$24073 ( \32295 , \31934 , \30899 );
or \U$24074 ( \32296 , \32294 , \32295 );
and \U$24075 ( \32297 , \32296 , \31814 );
or \U$24076 ( \32298 , \32290 , \32297 );
and \U$24078 ( \32299 , \32298 , 1'b1 );
or \U$24080 ( \32300 , \32299 , 1'b0 );
buf \U$24081 ( \32301 , \32300 );
_DC r23ca2_GF_IsGateDCbyConstraint ( \32302_nR23ca2 , \32301 , \21944 );
buf \U$24082 ( \32303 , \32302_nR23ca2 );
buf \U$24083 ( \32304 , RIb7b9680_245);
buf \U$24084 ( \32305 , RIb79b3b0_273);
nand \U$24085 ( \32306 , \32305 , \27360 );
not \U$24086 ( \32307 , \32306 );
and \U$24087 ( \32308 , \32304 , \32307 );
and \U$24088 ( \32309 , RIe51b690_6365, \32306 );
or \U$24089 ( \32310 , \32308 , \32309 );
and \U$24091 ( \32311 , \32310 , 1'b1 );
or \U$24093 ( \32312 , \32311 , 1'b0 );
buf \U$24094 ( \32313 , \32312 );
_DC r23ebc_GF_IsGateDCbyConstraint ( \32314_nR23ebc , \32313 , \21944 );
buf \U$24095 ( \32315 , \32314_nR23ebc );
not \U$24096 ( \32316 , \32306 );
not \U$24097 ( \32317 , \32316 );
and \U$24098 ( \32318 , RIe500d68_6388, \32317 );
buf \U$24099 ( \32319 , RIb7b96f8_244);
and \U$24100 ( \32320 , \32319 , \32316 );
or \U$24101 ( \32321 , \32318 , \32320 );
and \U$24103 ( \32322 , \32321 , 1'b1 );
or \U$24105 ( \32323 , \32322 , 1'b0 );
buf \U$24106 ( \32324 , \32323 );
_DC r23ebe_GF_IsGateDCbyConstraint ( \32325_nR23ebe , \32324 , \21944 );
buf \U$24107 ( \32326 , \32325_nR23ebe );
not \U$24108 ( \32327 , \32316 );
and \U$24109 ( \32328 , RIe501998_6387, \32327 );
buf \U$24110 ( \32329 , RIb7c20c8_243);
and \U$24111 ( \32330 , \32329 , \32316 );
or \U$24112 ( \32331 , \32328 , \32330 );
and \U$24114 ( \32332 , \32331 , 1'b1 );
or \U$24116 ( \32333 , \32332 , 1'b0 );
buf \U$24117 ( \32334 , \32333 );
_DC r23ec0_GF_IsGateDCbyConstraint ( \32335_nR23ec0 , \32334 , \21944 );
buf \U$24118 ( \32336 , \32335_nR23ec0 );
not \U$24119 ( \32337 , \32316 );
and \U$24120 ( \32338 , RIe5026b8_6386, \32337 );
buf \U$24121 ( \32339 , RIb7c5728_242);
and \U$24122 ( \32340 , \32339 , \32316 );
or \U$24123 ( \32341 , \32338 , \32340 );
and \U$24125 ( \32342 , \32341 , 1'b1 );
or \U$24127 ( \32343 , \32342 , 1'b0 );
buf \U$24128 ( \32344 , \32343 );
_DC r23ec2_GF_IsGateDCbyConstraint ( \32345_nR23ec2 , \32344 , \21944 );
buf \U$24129 ( \32346 , \32345_nR23ec2 );
not \U$24130 ( \32347 , \32316 );
and \U$24131 ( \32348 , RIe5032e8_6385, \32347 );
buf \U$24132 ( \32349 , RIb7c57a0_241);
and \U$24133 ( \32350 , \32349 , \32316 );
or \U$24134 ( \32351 , \32348 , \32350 );
and \U$24136 ( \32352 , \32351 , 1'b1 );
or \U$24138 ( \32353 , \32352 , 1'b0 );
buf \U$24139 ( \32354 , \32353 );
_DC r23ec4_GF_IsGateDCbyConstraint ( \32355_nR23ec4 , \32354 , \21944 );
buf \U$24140 ( \32356 , \32355_nR23ec4 );
not \U$24141 ( \32357 , \32316 );
and \U$24142 ( \32358 , RIe503f90_6384, \32357 );
buf \U$24143 ( \32359 , RIb7c5818_240);
and \U$24144 ( \32360 , \32359 , \32316 );
or \U$24145 ( \32361 , \32358 , \32360 );
and \U$24147 ( \32362 , \32361 , 1'b1 );
or \U$24149 ( \32363 , \32362 , 1'b0 );
buf \U$24150 ( \32364 , \32363 );
_DC r23ec6_GF_IsGateDCbyConstraint ( \32365_nR23ec6 , \32364 , \21944 );
buf \U$24151 ( \32366 , \32365_nR23ec6 );
not \U$24152 ( \32367 , \32316 );
and \U$24153 ( \32368 , RIe504d28_6383, \32367 );
buf \U$24154 ( \32369 , RIb7c5890_239);
and \U$24155 ( \32370 , \32369 , \32316 );
or \U$24156 ( \32371 , \32368 , \32370 );
and \U$24158 ( \32372 , \32371 , 1'b1 );
or \U$24160 ( \32373 , \32372 , 1'b0 );
buf \U$24161 ( \32374 , \32373 );
_DC r23ec8_GF_IsGateDCbyConstraint ( \32375_nR23ec8 , \32374 , \21944 );
buf \U$24162 ( \32376 , \32375_nR23ec8 );
not \U$24163 ( \32377 , \32316 );
and \U$24164 ( \32378 , RIe505958_6382, \32377 );
buf \U$24165 ( \32379 , RIb7c5908_238);
and \U$24166 ( \32380 , \32379 , \32316 );
or \U$24167 ( \32381 , \32378 , \32380 );
and \U$24169 ( \32382 , \32381 , 1'b1 );
or \U$24171 ( \32383 , \32382 , 1'b0 );
buf \U$24172 ( \32384 , \32383 );
_DC r23eca_GF_IsGateDCbyConstraint ( \32385_nR23eca , \32384 , \21944 );
buf \U$24173 ( \32386 , \32385_nR23eca );
not \U$24174 ( \32387 , \32316 );
and \U$24175 ( \32388 , RIe50ef58_6371, \32387 );
buf \U$24176 ( \32389 , RIb7a09f0_266);
and \U$24177 ( \32390 , \32389 , \32316 );
or \U$24178 ( \32391 , \32388 , \32390 );
and \U$24180 ( \32392 , \32391 , 1'b1 );
or \U$24182 ( \32393 , \32392 , 1'b0 );
buf \U$24183 ( \32394 , \32393 );
_DC r23eba_GF_IsGateDCbyConstraint ( \32395_nR23eba , \32394 , \21944 );
buf \U$24184 ( \32396 , \32395_nR23eba );
not \U$24185 ( \32397 , \32316 );
and \U$24186 ( \32398 , RIe50ac50_6376, \32397 );
buf \U$24187 ( \32399 , RIb7a0a68_265);
and \U$24188 ( \32400 , \32399 , \32316 );
or \U$24189 ( \32401 , \32398 , \32400 );
and \U$24191 ( \32402 , \32401 , 1'b1 );
or \U$24193 ( \32403 , \32402 , 1'b0 );
buf \U$24194 ( \32404 , \32403 );
_DC r23ecc_GF_IsGateDCbyConstraint ( \32405_nR23ecc , \32404 , \21944 );
buf \U$24195 ( \32406 , \32405_nR23ecc );
not \U$24196 ( \32407 , \32316 );
and \U$24197 ( \32408 , RIe50b880_6375, \32407 );
buf \U$24198 ( \32409 , RIb7a0ae0_264);
and \U$24199 ( \32410 , \32409 , \32316 );
or \U$24200 ( \32411 , \32408 , \32410 );
and \U$24202 ( \32412 , \32411 , 1'b1 );
or \U$24204 ( \32413 , \32412 , 1'b0 );
buf \U$24205 ( \32414 , \32413 );
_DC r23ece_GF_IsGateDCbyConstraint ( \32415_nR23ece , \32414 , \21944 );
buf \U$24206 ( \32416 , \32415_nR23ece );
not \U$24207 ( \32417 , \32316 );
and \U$24208 ( \32418 , RIe50c690_6374, \32417 );
buf \U$24209 ( \32419 , RIb7a0b58_263);
and \U$24210 ( \32420 , \32419 , \32316 );
or \U$24211 ( \32421 , \32418 , \32420 );
and \U$24213 ( \32422 , \32421 , 1'b1 );
or \U$24215 ( \32423 , \32422 , 1'b0 );
buf \U$24216 ( \32424 , \32423 );
_DC r23ed0_GF_IsGateDCbyConstraint ( \32425_nR23ed0 , \32424 , \21944 );
buf \U$24217 ( \32426 , \32425_nR23ed0 );
not \U$24218 ( \32427 , \32316 );
and \U$24219 ( \32428 , RIe50d428_6373, \32427 );
buf \U$24220 ( \32429 , RIb7a0bd0_262);
and \U$24221 ( \32430 , \32429 , \32316 );
or \U$24222 ( \32431 , \32428 , \32430 );
and \U$24224 ( \32432 , \32431 , 1'b1 );
or \U$24226 ( \32433 , \32432 , 1'b0 );
buf \U$24227 ( \32434 , \32433 );
_DC r23ed2_GF_IsGateDCbyConstraint ( \32435_nR23ed2 , \32434 , \21944 );
buf \U$24228 ( \32436 , \32435_nR23ed2 );
not \U$24229 ( \32437 , RIe523688_6352);
not \U$24230 ( \32438 , \32437 );
or \U$24231 ( \32439 , RIe524060_6351, \32438 );
not \U$24232 ( \32440 , \32439 );
and \U$24233 ( \32441 , \32440 , RIe524948_6350);
nand \U$24234 ( \32442 , \27356 , \27360 );
not \U$24235 ( \32443 , \32442 );
not \U$24236 ( \32444 , RIe5117a8_6369);
or \U$24237 ( \32445 , \32304 , \32444 );
nand \U$24238 ( \32446 , \32445 , \27356 , \27360 );
buf \U$24239 ( \32447 , RIb79b4a0_271);
nor \U$24240 ( \32448 , RIea91330_6888, \9126 );
buf \U$24241 ( \32449 , \32448 );
nand \U$24242 ( \32450 , \32447 , \32449 );
not \U$24243 ( \32451 , \32450 );
buf \U$24244 ( \32452 , \21709 );
nand \U$24245 ( \32453 , \32449 , \32452 );
not \U$24246 ( \32454 , \32453 );
nor \U$24247 ( \32455 , \32451 , \32454 );
nand \U$24248 ( \32456 , \32443 , \32446 , \32455 );
or \U$24249 ( \32457 , \32441 , \32456 );
nand \U$24250 ( \32458 , \27356 , \27360 );
not \U$24251 ( \32459 , \32458 );
not \U$24252 ( \32460 , \32459 );
and \U$24253 ( \32461 , \32453 , \32451 );
not \U$24254 ( \32462 , \32439 );
not \U$24255 ( \32463 , \32462 );
or \U$24256 ( \32464 , RIe524948_6350, \32463 );
nand \U$24257 ( \32465 , \32460 , \32461 , \32464 );
nand \U$24258 ( \32466 , \32457 , \32465 );
not \U$24259 ( \32467 , \32466 );
or \U$24260 ( \32468 , \32459 , \32462 );
not \U$24261 ( \32469 , \32437 );
nand \U$24262 ( \32470 , RIe524060_6351, \32469 );
nand \U$24263 ( \32471 , \32468 , \32470 );
xnor \U$24264 ( \32472 , \32471 , \32458 );
nor \U$24265 ( \32473 , \32467 , \32472 );
not \U$24266 ( \32474 , \32473 );
not \U$24267 ( \32475 , RIe524948_6350);
and \U$24268 ( \32476 , \32474 , \32475 );
not \U$24269 ( \32477 , \32454 );
not \U$24270 ( \32478 , \32446 );
not \U$24271 ( \32479 , \32478 );
xnor \U$24272 ( \32480 , \32451 , \32459 );
and \U$24273 ( \32481 , \32477 , \32479 , \32480 );
not \U$24274 ( \32482 , \32481 );
not \U$24275 ( \32483 , \32482 );
not \U$24276 ( \32484 , \32483 );
not \U$24277 ( \32485 , \32472 );
and \U$24278 ( \32486 , \32484 , \32485 );
nand \U$24279 ( \32487 , \32456 , \32465 );
nor \U$24280 ( \32488 , \32483 , \32487 );
nor \U$24281 ( \32489 , \32486 , \32488 );
not \U$24282 ( \32490 , \32489 );
and \U$24283 ( \32491 , \32490 , RIe524948_6350);
or \U$24284 ( \32492 , \32476 , \32491 );
not \U$24285 ( \32493 , RIe51d5f8_6362);
nand \U$24286 ( \32494 , \32478 , \32453 );
not \U$24287 ( \32495 , \32494 );
not \U$24288 ( \32496 , \32495 );
or \U$24289 ( \32497 , \32493 , \32496 );
not \U$24290 ( \32498 , \32494 );
and \U$24291 ( \32499 , RIe51c158_6364, \32498 );
not \U$24292 ( \32500 , \32483 );
not \U$24293 ( \32501 , \32437 );
and \U$24294 ( \32502 , \32500 , \32501 );
not \U$24295 ( \32503 , \32466 );
and \U$24296 ( \32504 , \32503 , \32437 );
or \U$24297 ( \32505 , \32502 , \32504 );
not \U$24298 ( \32506 , \32505 );
or \U$24299 ( \32507 , \32499 , \32506 );
nand \U$24300 ( \32508 , \32462 , \32458 );
not \U$24301 ( \32509 , \32459 );
or \U$24302 ( \32510 , \32437 , \32509 );
not \U$24303 ( \32511 , \32510 );
not \U$24304 ( \32512 , RIe524060_6351);
and \U$24305 ( \32513 , \32511 , \32512 );
xnor \U$24306 ( \32514 , \32459 , \32469 );
not \U$24307 ( \32515 , \32514 );
and \U$24308 ( \32516 , \32515 , RIe524060_6351);
or \U$24309 ( \32517 , \32513 , \32516 );
not \U$24310 ( \32518 , \32517 );
and \U$24311 ( \32519 , \32508 , \32518 );
or \U$24312 ( \32520 , \32467 , \32519 );
and \U$24313 ( \32521 , \32483 , RIe524060_6351);
not \U$24314 ( \32522 , \32494 );
and \U$24315 ( \32523 , RIe51cc20_6363, \32522 );
nor \U$24316 ( \32524 , \32521 , \32523 );
nand \U$24317 ( \32525 , \32520 , \32524 );
nor \U$24318 ( \32526 , \32507 , \32525 );
and \U$24319 ( \32527 , \32492 , \32497 , \32526 );
buf \U$24320 ( \32528 , RIb839668_156);
buf \U$24321 ( \32529 , \32528 );
not \U$24322 ( \32530 , \32529 );
not \U$24323 ( \32531 , \32530 );
buf \U$24324 ( \32532 , RIb839848_152);
and \U$24325 ( \32533 , \32532 , \27349 );
buf \U$24326 ( \32534 , RIb8396e0_155);
nand \U$24327 ( \32535 , \32534 , \27349 );
not \U$24328 ( \32536 , \32535 );
buf \U$24329 ( \32537 , \32536 );
or \U$24330 ( \32538 , \32531 , \32533 , \32537 );
nand \U$24331 ( \32539 , \32538 , \27349 );
not \U$24332 ( \32540 , \32539 );
not \U$24333 ( \32541 , RIe51f290_6359);
or \U$24334 ( \32542 , \32540 , \32541 );
nand \U$24335 ( \32543 , \32535 , \32530 );
not \U$24336 ( \32544 , RIe51e840_6360);
not \U$24337 ( \32545 , \32544 );
or \U$24338 ( \32546 , \32541 , \32545 );
not \U$24339 ( \32547 , \32546 );
nand \U$24340 ( \32548 , RIe51dee0_6361, \32547 );
or \U$24341 ( \32549 , \32543 , \32548 );
xor \U$24342 ( \32550 , \32541 , \32544 );
nor \U$24343 ( \32551 , \32550 , \32547 );
nand \U$24344 ( \32552 , \27349 , \32535 , \32529 );
or \U$24345 ( \32553 , \32551 , \32552 );
not \U$24346 ( \32554 , \32543 );
nand \U$24347 ( \32555 , \32533 , \32548 , \32554 );
not \U$24348 ( \32556 , RIe51dee0_6361);
nor \U$24349 ( \32557 , \32544 , \32556 );
xor \U$24350 ( \32558 , \32541 , \32557 );
or \U$24351 ( \32559 , \32555 , \32558 );
nand \U$24352 ( \32560 , \32542 , \32549 , \32553 , \32559 );
not \U$24353 ( \32561 , RIe525410_6349);
not \U$24354 ( \32562 , RIe525d70_6348);
not \U$24355 ( \32563 , RIe5267c0_6347);
not \U$24356 ( \32564 , \32563 );
nand \U$24357 ( \32565 , \32561 , \32562 , \32564 );
not \U$24358 ( \32566 , \32565 );
not \U$24359 ( \32567 , \32566 );
not \U$24360 ( \32568 , \32451 );
and \U$24361 ( \32569 , \32564 , \32568 );
nor \U$24362 ( \32570 , \32562 , \32561 );
xnor \U$24363 ( \32571 , \32563 , \32570 );
and \U$24364 ( \32572 , \32571 , \32451 );
or \U$24365 ( \32573 , \32569 , \32572 );
not \U$24366 ( \32574 , \32573 );
and \U$24367 ( \32575 , \32567 , \32574 );
nor \U$24368 ( \32576 , \32575 , \32454 );
not \U$24369 ( \32577 , \32576 );
or \U$24370 ( \32578 , \32560 , \32577 );
or \U$24371 ( \32579 , \32540 , \32556 );
or \U$24372 ( \32580 , \32543 , \32548 );
or \U$24373 ( \32581 , \32555 , RIe51dee0_6361);
nand \U$24374 ( \32582 , \32529 , \27349 );
not \U$24375 ( \32583 , \32582 );
nand \U$24376 ( \32584 , \32583 , \32534 );
not \U$24377 ( \32585 , \32584 );
nand \U$24378 ( \32586 , RIe51dee0_6361, \32546 );
and \U$24379 ( \32587 , \32548 , \32586 );
or \U$24380 ( \32588 , \32587 , \32582 );
and \U$24381 ( \32589 , \32588 , \32535 );
or \U$24382 ( \32590 , \32585 , \32589 );
nand \U$24383 ( \32591 , \32579 , \32580 , \32581 , \32590 );
not \U$24384 ( \32592 , \32591 );
xor \U$24385 ( \32593 , \32544 , \32556 );
not \U$24386 ( \32594 , \32555 );
and \U$24387 ( \32595 , \32593 , \32594 );
not \U$24388 ( \32596 , \32544 );
not \U$24389 ( \32597 , \32596 );
not \U$24390 ( \32598 , \32539 );
or \U$24391 ( \32599 , \32597 , \32598 );
not \U$24392 ( \32600 , \32552 );
nand \U$24393 ( \32601 , \32544 , \32546 , \32600 );
nand \U$24394 ( \32602 , \32599 , \32601 , \32584 );
or \U$24395 ( \32603 , \32595 , \32602 );
xor \U$24396 ( \32604 , \32562 , \32561 );
and \U$24397 ( \32605 , \32604 , \32565 , \32461 );
not \U$24398 ( \32606 , \32562 );
and \U$24399 ( \32607 , \32450 , \32606 , \32453 );
or \U$24400 ( \32608 , \32605 , \32607 );
not \U$24401 ( \32609 , \32608 );
or \U$24402 ( \32610 , \32603 , \32609 );
and \U$24403 ( \32611 , \32561 , \32565 , \32461 );
not \U$24404 ( \32612 , \32561 );
and \U$24405 ( \32613 , \32450 , \32612 , \32453 );
nor \U$24406 ( \32614 , \32611 , \32613 );
nand \U$24407 ( \32615 , \32610 , \32614 );
or \U$24408 ( \32616 , \32592 , \32615 );
nand \U$24409 ( \32617 , \32603 , \32609 );
nand \U$24410 ( \32618 , \32616 , \32617 );
nand \U$24411 ( \32619 , \32578 , \32618 );
and \U$24412 ( \32620 , \32560 , \32577 );
not \U$24413 ( \32621 , RIe5117a8_6369);
not \U$24414 ( \32622 , \32310 );
nor \U$24415 ( \32623 , \32620 , \32621 , \32622 );
and \U$24416 ( \32624 , \32619 , \32623 );
nor \U$24417 ( \32625 , \32527 , \32624 );
and \U$24419 ( \32626 , \32625 , 1'b1 );
or \U$24421 ( \32627 , \32626 , 1'b0 );
buf \U$24422 ( \32628 , \32627 );
_DC r23eb8_GF_IsGateDCbyConstraint ( \32629_nR23eb8 , \32628 , \21944 );
buf \U$24423 ( \32630 , \32629_nR23eb8 );
and \U$24425 ( \32631 , \32507 , 1'b1 );
or \U$24427 ( \32632 , \32631 , 1'b0 );
buf \U$24428 ( \32633 , \32632 );
_DC r23eea_GF_IsGateDCbyConstraint ( \32634_nR23eea , \32633 , \21944 );
buf \U$24429 ( \32635 , \32634_nR23eea );
and \U$24431 ( \32636 , \32525 , 1'b1 );
or \U$24433 ( \32637 , \32636 , 1'b0 );
buf \U$24434 ( \32638 , \32637 );
_DC r23eec_GF_IsGateDCbyConstraint ( \32639_nR23eec , \32638 , \21944 );
buf \U$24435 ( \32640 , \32639_nR23eec );
not \U$24436 ( \32641 , \32497 );
not \U$24437 ( \32642 , \32492 );
or \U$24438 ( \32643 , \32641 , \32642 );
and \U$24440 ( \32644 , \32643 , 1'b1 );
or \U$24442 ( \32645 , \32644 , 1'b0 );
buf \U$24443 ( \32646 , \32645 );
_DC r23eee_GF_IsGateDCbyConstraint ( \32647_nR23eee , \32646 , \21944 );
buf \U$24444 ( \32648 , \32647_nR23eee );
not \U$24445 ( \32649 , \21812 );
nand \U$24446 ( \32650 , \32649 , \21810 , RIe546098_6850);
nor \U$24447 ( \32651 , \21809 , \32650 );
buf \U$24448 ( \32652 , \32651 );
buf \U$24449 ( \32653 , \32652 );
not \U$24450 ( \32654 , \22095 );
buf \U$24451 ( \32655 , \32654 );
buf \U$24452 ( \32656 , \32655 );
nand \U$24453 ( \32657 , \32653 , \32656 );
buf \U$24454 ( \32658 , \8825 );
buf \U$24455 ( \32659 , \32658 );
not \U$24456 ( \32660 , \27237 );
and \U$24457 ( \32661 , \32660 , \21694 );
buf \U$24458 ( \32662 , \32661 );
buf \U$24459 ( \32663 , \32662 );
nand \U$24460 ( \32664 , \32659 , \32663 );
nand \U$24461 ( \32665 , \32657 , \32664 );
buf \U$24462 ( \32666 , \32665 );
not \U$24463 ( \32667 , \32666 );
and \U$24464 ( \32668 , RIe1e2210_5688, \32667 );
not \U$24465 ( \32669 , RIe1e2210_5688);
buf \U$24466 ( \32670 , \27369 );
buf \U$24467 ( \32671 , RIe667f70_6886);
buf \U$24468 ( \32672 , \32671 );
not \U$24469 ( \32673 , \32672 );
not \U$24470 ( \32674 , \32673 );
or \U$24471 ( \32675 , \32670 , \32674 );
not \U$24472 ( \32676 , \32675 );
nand \U$24473 ( \32677 , \32664 , \32676 );
buf \U$24474 ( \32678 , \27379 );
not \U$24475 ( \32679 , \32678 );
buf \U$24476 ( \32680 , \22120 );
not \U$24477 ( \32681 , \32680 );
not \U$24478 ( \32682 , \32664 );
and \U$24479 ( \32683 , \32679 , \32681 , \32682 );
not \U$24480 ( \32684 , \32683 );
buf \U$24481 ( \32685 , \32684 );
nand \U$24482 ( \32686 , \32677 , \32685 );
not \U$24483 ( \32687 , \32686 );
not \U$24484 ( \32688 , \32687 );
or \U$24485 ( \32689 , \32669 , \32688 );
not \U$24486 ( \32690 , \32677 );
buf \U$24487 ( \32691 , RIb87eb00_69);
and \U$24488 ( \32692 , \32690 , \32691 );
buf \U$24489 ( \32693 , RIb7c5980_237);
buf \U$24490 ( \32694 , \32693 );
not \U$24491 ( \32695 , \32685 );
and \U$24492 ( \32696 , \32694 , \32695 );
nor \U$24493 ( \32697 , \32692 , \32696 );
nand \U$24494 ( \32698 , \32689 , \32697 );
and \U$24495 ( \32699 , \32698 , \32666 );
or \U$24496 ( \32700 , \32668 , \32699 );
and \U$24498 ( \32701 , \32700 , 1'b1 );
or \U$24500 ( \32702 , \32701 , 1'b0 );
buf \U$24501 ( \32703 , \32702 );
_DC r23a0c_GF_IsGateDCbyConstraint ( \32704_nR23a0c , \32703 , \21944 );
buf \U$24502 ( \32705 , \32704_nR23a0c );
not \U$24503 ( \32706 , \32666 );
and \U$24504 ( \32707 , RIe1e10b8_5689, \32706 );
not \U$24505 ( \32708 , RIe1e10b8_5689);
not \U$24506 ( \32709 , \32678 );
not \U$24507 ( \32710 , \32680 );
and \U$24508 ( \32711 , \32709 , \32710 , \32682 );
not \U$24509 ( \32712 , \32711 );
buf \U$24510 ( \32713 , \32712 );
and \U$24511 ( \32714 , \32677 , \32713 );
not \U$24512 ( \32715 , \32714 );
or \U$24513 ( \32716 , \32708 , \32715 );
buf \U$24514 ( \32717 , \32690 );
buf \U$24515 ( \32718 , RIb87eb78_68);
buf \U$24516 ( \32719 , \32718 );
and \U$24517 ( \32720 , \32717 , \32719 );
buf \U$24518 ( \32721 , RIb7c59f8_236);
buf \U$24519 ( \32722 , \32721 );
buf \U$24520 ( \32723 , \32684 );
not \U$24521 ( \32724 , \32723 );
and \U$24522 ( \32725 , \32722 , \32724 );
nor \U$24523 ( \32726 , \32720 , \32725 );
nand \U$24524 ( \32727 , \32716 , \32726 );
and \U$24525 ( \32728 , \32727 , \32666 );
or \U$24526 ( \32729 , \32707 , \32728 );
and \U$24528 ( \32730 , \32729 , 1'b1 );
or \U$24530 ( \32731 , \32730 , 1'b0 );
buf \U$24531 ( \32732 , \32731 );
_DC r23a22_GF_IsGateDCbyConstraint ( \32733_nR23a22 , \32732 , \21944 );
buf \U$24532 ( \32734 , \32733_nR23a22 );
not \U$24533 ( \32735 , \32666 );
and \U$24534 ( \32736 , RIe1dfab0_5690, \32735 );
not \U$24535 ( \32737 , RIe1dfab0_5690);
or \U$24536 ( \32738 , \32737 , \32688 );
buf \U$24537 ( \32739 , \32690 );
buf \U$24538 ( \32740 , RIb87ebf0_67);
and \U$24539 ( \32741 , \32739 , \32740 );
buf \U$24540 ( \32742 , RIb7c5a70_235);
buf \U$24541 ( \32743 , \32742 );
not \U$24542 ( \32744 , \32685 );
and \U$24543 ( \32745 , \32743 , \32744 );
nor \U$24544 ( \32746 , \32741 , \32745 );
nand \U$24545 ( \32747 , \32738 , \32746 );
and \U$24546 ( \32748 , \32747 , \32666 );
or \U$24547 ( \32749 , \32736 , \32748 );
and \U$24549 ( \32750 , \32749 , 1'b1 );
or \U$24551 ( \32751 , \32750 , 1'b0 );
buf \U$24552 ( \32752 , \32751 );
_DC r23a38_GF_IsGateDCbyConstraint ( \32753_nR23a38 , \32752 , \21944 );
buf \U$24553 ( \32754 , \32753_nR23a38 );
buf \U$24554 ( \32755 , \32665 );
buf \U$24555 ( \32756 , \32755 );
not \U$24556 ( \32757 , \32756 );
and \U$24557 ( \32758 , RIe1de958_5691, \32757 );
not \U$24558 ( \32759 , RIe1de958_5691);
or \U$24559 ( \32760 , \32759 , \32715 );
buf \U$24560 ( \32761 , RIb882ca0_66);
and \U$24561 ( \32762 , \32690 , \32761 );
buf \U$24562 ( \32763 , RIb7cade0_234);
buf \U$24563 ( \32764 , \32763 );
not \U$24564 ( \32765 , \32713 );
and \U$24565 ( \32766 , \32764 , \32765 );
nor \U$24566 ( \32767 , \32762 , \32766 );
nand \U$24567 ( \32768 , \32760 , \32767 );
and \U$24568 ( \32769 , \32768 , \32756 );
or \U$24569 ( \32770 , \32758 , \32769 );
and \U$24571 ( \32771 , \32770 , 1'b1 );
or \U$24573 ( \32772 , \32771 , 1'b0 );
buf \U$24574 ( \32773 , \32772 );
_DC r23a4e_GF_IsGateDCbyConstraint ( \32774_nR23a4e , \32773 , \21944 );
buf \U$24575 ( \32775 , \32774_nR23a4e );
not \U$24576 ( \32776 , \32756 );
and \U$24577 ( \32777 , RIe1dd350_5692, \32776 );
not \U$24578 ( \32778 , RIe1dd350_5692);
not \U$24579 ( \32779 , \32687 );
or \U$24580 ( \32780 , \32778 , \32779 );
buf \U$24581 ( \32781 , \32690 );
buf \U$24582 ( \32782 , RIb885310_65);
buf \U$24583 ( \32783 , \32782 );
and \U$24584 ( \32784 , \32781 , \32783 );
buf \U$24585 ( \32785 , RIb7cae58_233);
buf \U$24586 ( \32786 , \32785 );
not \U$24587 ( \32787 , \32723 );
and \U$24588 ( \32788 , \32786 , \32787 );
nor \U$24589 ( \32789 , \32784 , \32788 );
nand \U$24590 ( \32790 , \32780 , \32789 );
and \U$24591 ( \32791 , \32790 , \32756 );
or \U$24592 ( \32792 , \32777 , \32791 );
and \U$24594 ( \32793 , \32792 , 1'b1 );
or \U$24596 ( \32794 , \32793 , 1'b0 );
buf \U$24597 ( \32795 , \32794 );
_DC r23a64_GF_IsGateDCbyConstraint ( \32796_nR23a64 , \32795 , \21944 );
buf \U$24598 ( \32797 , \32796_nR23a64 );
not \U$24599 ( \32798 , \32666 );
and \U$24600 ( \32799 , RIe1dc1f8_5693, \32798 );
not \U$24601 ( \32800 , RIe1dc1f8_5693);
not \U$24602 ( \32801 , \32714 );
or \U$24603 ( \32802 , \32800 , \32801 );
buf \U$24604 ( \32803 , RIb885388_64);
buf \U$24605 ( \32804 , \32803 );
and \U$24606 ( \32805 , \32781 , \32804 );
buf \U$24607 ( \32806 , \22248 );
not \U$24608 ( \32807 , \32678 );
not \U$24609 ( \32808 , \32680 );
and \U$24610 ( \32809 , \32807 , \32808 , \32682 );
not \U$24611 ( \32810 , \32809 );
buf \U$24612 ( \32811 , \32810 );
not \U$24613 ( \32812 , \32811 );
and \U$24614 ( \32813 , \32806 , \32812 );
nor \U$24615 ( \32814 , \32805 , \32813 );
nand \U$24616 ( \32815 , \32802 , \32814 );
and \U$24617 ( \32816 , \32815 , \32666 );
or \U$24618 ( \32817 , \32799 , \32816 );
and \U$24620 ( \32818 , \32817 , 1'b1 );
or \U$24622 ( \32819 , \32818 , 1'b0 );
buf \U$24623 ( \32820 , \32819 );
_DC r23a7a_GF_IsGateDCbyConstraint ( \32821_nR23a7a , \32820 , \21944 );
buf \U$24624 ( \32822 , \32821_nR23a7a );
not \U$24625 ( \32823 , \32666 );
and \U$24626 ( \32824 , RIe1dabf0_5694, \32823 );
not \U$24627 ( \32825 , RIe1dabf0_5694);
or \U$24628 ( \32826 , \32825 , \32686 );
buf \U$24629 ( \32827 , RIb885400_63);
and \U$24630 ( \32828 , \32739 , \32827 );
buf \U$24631 ( \32829 , \22274 );
not \U$24632 ( \32830 , \32713 );
and \U$24633 ( \32831 , \32829 , \32830 );
nor \U$24634 ( \32832 , \32828 , \32831 );
nand \U$24635 ( \32833 , \32826 , \32832 );
and \U$24636 ( \32834 , \32833 , \32666 );
or \U$24637 ( \32835 , \32824 , \32834 );
and \U$24639 ( \32836 , \32835 , 1'b1 );
or \U$24641 ( \32837 , \32836 , 1'b0 );
buf \U$24642 ( \32838 , \32837 );
_DC r23a84_GF_IsGateDCbyConstraint ( \32839_nR23a84 , \32838 , \21944 );
buf \U$24643 ( \32840 , \32839_nR23a84 );
buf \U$24644 ( \32841 , \32665 );
buf \U$24645 ( \32842 , \32841 );
not \U$24646 ( \32843 , \32842 );
and \U$24647 ( \32844 , RIe1d9a98_5695, \32843 );
not \U$24648 ( \32845 , RIe1d9a98_5695);
or \U$24649 ( \32846 , \32845 , \32715 );
buf \U$24650 ( \32847 , RIb885478_62);
buf \U$24651 ( \32848 , \32847 );
and \U$24652 ( \32849 , \32781 , \32848 );
buf \U$24653 ( \32850 , RIb7cafc0_230);
buf \U$24654 ( \32851 , \32850 );
buf \U$24655 ( \32852 , \32810 );
not \U$24656 ( \32853 , \32852 );
and \U$24657 ( \32854 , \32851 , \32853 );
nor \U$24658 ( \32855 , \32849 , \32854 );
nand \U$24659 ( \32856 , \32846 , \32855 );
and \U$24660 ( \32857 , \32856 , \32842 );
or \U$24661 ( \32858 , \32844 , \32857 );
and \U$24663 ( \32859 , \32858 , 1'b1 );
or \U$24665 ( \32860 , \32859 , 1'b0 );
buf \U$24666 ( \32861 , \32860 );
_DC r23a86_GF_IsGateDCbyConstraint ( \32862_nR23a86 , \32861 , \21944 );
buf \U$24667 ( \32863 , \32862_nR23a86 );
buf \U$24668 ( \32864 , \32841 );
not \U$24669 ( \32865 , \32864 );
and \U$24670 ( \32866 , RIe1d8940_5696, \32865 );
not \U$24671 ( \32867 , RIe1d8940_5696);
not \U$24672 ( \32868 , \32714 );
or \U$24673 ( \32869 , \32867 , \32868 );
buf \U$24674 ( \32870 , \27564 );
and \U$24675 ( \32871 , \32690 , \32870 );
buf \U$24676 ( \32872 , RIb7cb038_229);
buf \U$24677 ( \32873 , \32872 );
buf \U$24678 ( \32874 , \32810 );
not \U$24679 ( \32875 , \32874 );
and \U$24680 ( \32876 , \32873 , \32875 );
nor \U$24681 ( \32877 , \32871 , \32876 );
nand \U$24682 ( \32878 , \32869 , \32877 );
and \U$24683 ( \32879 , \32878 , \32864 );
or \U$24684 ( \32880 , \32866 , \32879 );
and \U$24686 ( \32881 , \32880 , 1'b1 );
or \U$24688 ( \32882 , \32881 , 1'b0 );
buf \U$24689 ( \32883 , \32882 );
_DC r23a88_GF_IsGateDCbyConstraint ( \32884_nR23a88 , \32883 , \21944 );
buf \U$24690 ( \32885 , \32884_nR23a88 );
not \U$24691 ( \32886 , \32756 );
and \U$24692 ( \32887 , RIe1d7338_5697, \32886 );
not \U$24693 ( \32888 , RIe1d7338_5697);
not \U$24694 ( \32889 , \32714 );
or \U$24695 ( \32890 , \32888 , \32889 );
buf \U$24696 ( \32891 , \22334 );
and \U$24697 ( \32892 , \32781 , \32891 );
buf \U$24698 ( \32893 , RIb7cb0b0_228);
buf \U$24699 ( \32894 , \32893 );
buf \U$24700 ( \32895 , \32712 );
not \U$24701 ( \32896 , \32895 );
and \U$24702 ( \32897 , \32894 , \32896 );
nor \U$24703 ( \32898 , \32892 , \32897 );
nand \U$24704 ( \32899 , \32890 , \32898 );
and \U$24705 ( \32900 , \32899 , \32756 );
or \U$24706 ( \32901 , \32887 , \32900 );
and \U$24708 ( \32902 , \32901 , 1'b1 );
or \U$24710 ( \32903 , \32902 , 1'b0 );
buf \U$24711 ( \32904 , \32903 );
_DC r23a8a_GF_IsGateDCbyConstraint ( \32905_nR23a8a , \32904 , \21944 );
buf \U$24712 ( \32906 , \32905_nR23a8a );
not \U$24713 ( \32907 , \32666 );
and \U$24714 ( \32908 , RIe1d61e0_5698, \32907 );
not \U$24715 ( \32909 , RIe1d61e0_5698);
not \U$24716 ( \32910 , \32687 );
or \U$24717 ( \32911 , \32909 , \32910 );
buf \U$24718 ( \32912 , \22356 );
and \U$24719 ( \32913 , \32717 , \32912 );
buf \U$24720 ( \32914 , \22359 );
not \U$24721 ( \32915 , \32811 );
and \U$24722 ( \32916 , \32914 , \32915 );
nor \U$24723 ( \32917 , \32913 , \32916 );
nand \U$24724 ( \32918 , \32911 , \32917 );
and \U$24725 ( \32919 , \32918 , \32666 );
or \U$24726 ( \32920 , \32908 , \32919 );
and \U$24728 ( \32921 , \32920 , 1'b1 );
or \U$24730 ( \32922 , \32921 , 1'b0 );
buf \U$24731 ( \32923 , \32922 );
_DC r23a0e_GF_IsGateDCbyConstraint ( \32924_nR23a0e , \32923 , \21944 );
buf \U$24732 ( \32925 , \32924_nR23a0e );
not \U$24733 ( \32926 , \32842 );
and \U$24734 ( \32927 , RIe1d4bd8_5699, \32926 );
not \U$24735 ( \32928 , RIe1d4bd8_5699);
or \U$24736 ( \32929 , \32928 , \32779 );
buf \U$24737 ( \32930 , RIb885658_58);
buf \U$24738 ( \32931 , \32930 );
and \U$24739 ( \32932 , \32739 , \32931 );
buf \U$24740 ( \32933 , RIb7d00d8_226);
buf \U$24741 ( \32934 , \32933 );
not \U$24742 ( \32935 , \32852 );
and \U$24743 ( \32936 , \32934 , \32935 );
nor \U$24744 ( \32937 , \32932 , \32936 );
nand \U$24745 ( \32938 , \32929 , \32937 );
and \U$24746 ( \32939 , \32938 , \32842 );
or \U$24747 ( \32940 , \32927 , \32939 );
and \U$24749 ( \32941 , \32940 , 1'b1 );
or \U$24751 ( \32942 , \32941 , 1'b0 );
buf \U$24752 ( \32943 , \32942 );
_DC r23a10_GF_IsGateDCbyConstraint ( \32944_nR23a10 , \32943 , \21944 );
buf \U$24753 ( \32945 , \32944_nR23a10 );
not \U$24754 ( \32946 , \32666 );
and \U$24755 ( \32947 , RIe1d3a80_5700, \32946 );
not \U$24756 ( \32948 , RIe1d3a80_5700);
not \U$24757 ( \32949 , \32687 );
or \U$24758 ( \32950 , \32948 , \32949 );
buf \U$24759 ( \32951 , \22397 );
and \U$24760 ( \32952 , \32717 , \32951 );
buf \U$24761 ( \32953 , \22400 );
not \U$24762 ( \32954 , \32874 );
and \U$24763 ( \32955 , \32953 , \32954 );
nor \U$24764 ( \32956 , \32952 , \32955 );
nand \U$24765 ( \32957 , \32950 , \32956 );
and \U$24766 ( \32958 , \32957 , \32666 );
or \U$24767 ( \32959 , \32947 , \32958 );
and \U$24769 ( \32960 , \32959 , 1'b1 );
or \U$24771 ( \32961 , \32960 , 1'b0 );
buf \U$24772 ( \32962 , \32961 );
_DC r23a12_GF_IsGateDCbyConstraint ( \32963_nR23a12 , \32962 , \21944 );
buf \U$24773 ( \32964 , \32963_nR23a12 );
not \U$24774 ( \32965 , \32666 );
and \U$24775 ( \32966 , RIe1d2478_5701, \32965 );
not \U$24776 ( \32967 , RIe1d2478_5701);
not \U$24777 ( \32968 , \32714 );
or \U$24778 ( \32969 , \32967 , \32968 );
buf \U$24779 ( \32970 , \22417 );
and \U$24780 ( \32971 , \32717 , \32970 );
buf \U$24781 ( \32972 , RIb826e28_224);
buf \U$24782 ( \32973 , \32972 );
buf \U$24783 ( \32974 , \32712 );
not \U$24784 ( \32975 , \32974 );
and \U$24785 ( \32976 , \32973 , \32975 );
nor \U$24786 ( \32977 , \32971 , \32976 );
nand \U$24787 ( \32978 , \32969 , \32977 );
and \U$24788 ( \32979 , \32978 , \32666 );
or \U$24789 ( \32980 , \32966 , \32979 );
and \U$24791 ( \32981 , \32980 , 1'b1 );
or \U$24793 ( \32982 , \32981 , 1'b0 );
buf \U$24794 ( \32983 , \32982 );
_DC r23a14_GF_IsGateDCbyConstraint ( \32984_nR23a14 , \32983 , \21944 );
buf \U$24795 ( \32985 , \32984_nR23a14 );
not \U$24796 ( \32986 , \32666 );
and \U$24797 ( \32987 , RIe099530_5702, \32986 );
not \U$24798 ( \32988 , RIe099530_5702);
or \U$24799 ( \32989 , \32988 , \32801 );
buf \U$24800 ( \32990 , RIb8857c0_55);
buf \U$24801 ( \32991 , \32990 );
and \U$24802 ( \32992 , \32781 , \32991 );
buf \U$24803 ( \32993 , RIb826ea0_223);
buf \U$24804 ( \32994 , \32993 );
not \U$24805 ( \32995 , \32895 );
and \U$24806 ( \32996 , \32994 , \32995 );
nor \U$24807 ( \32997 , \32992 , \32996 );
nand \U$24808 ( \32998 , \32989 , \32997 );
and \U$24809 ( \32999 , \32998 , \32666 );
or \U$24810 ( \33000 , \32987 , \32999 );
and \U$24812 ( \33001 , \33000 , 1'b1 );
or \U$24814 ( \33002 , \33001 , 1'b0 );
buf \U$24815 ( \33003 , \33002 );
_DC r23a16_GF_IsGateDCbyConstraint ( \33004_nR23a16 , \33003 , \21944 );
buf \U$24816 ( \33005 , \33004_nR23a16 );
not \U$24817 ( \33006 , \32756 );
and \U$24818 ( \33007 , RIe09d298_5703, \33006 );
not \U$24819 ( \33008 , RIe09d298_5703);
or \U$24820 ( \33009 , \33008 , \32688 );
buf \U$24821 ( \33010 , RIb885838_54);
buf \U$24822 ( \33011 , \33010 );
and \U$24823 ( \33012 , \32717 , \33011 );
buf \U$24824 ( \33013 , RIb826f18_222);
buf \U$24825 ( \33014 , \33013 );
not \U$24826 ( \33015 , \32713 );
and \U$24827 ( \33016 , \33014 , \33015 );
nor \U$24828 ( \33017 , \33012 , \33016 );
nand \U$24829 ( \33018 , \33009 , \33017 );
and \U$24830 ( \33019 , \33018 , \32756 );
or \U$24831 ( \33020 , \33007 , \33019 );
and \U$24833 ( \33021 , \33020 , 1'b1 );
or \U$24835 ( \33022 , \33021 , 1'b0 );
buf \U$24836 ( \33023 , \33022 );
_DC r23a18_GF_IsGateDCbyConstraint ( \33024_nR23a18 , \33023 , \21944 );
buf \U$24837 ( \33025 , \33024_nR23a18 );
not \U$24838 ( \33026 , \32756 );
and \U$24839 ( \33027 , RIe0a2338_5704, \33026 );
not \U$24840 ( \33028 , RIe0a2338_5704);
or \U$24841 ( \33029 , \33028 , \32910 );
buf \U$24842 ( \33030 , RIb8858b0_53);
and \U$24843 ( \33031 , \32717 , \33030 );
buf \U$24844 ( \33032 , RIb826f90_221);
buf \U$24845 ( \33033 , \33032 );
not \U$24846 ( \33034 , \32723 );
and \U$24847 ( \33035 , \33033 , \33034 );
nor \U$24848 ( \33036 , \33031 , \33035 );
nand \U$24849 ( \33037 , \33029 , \33036 );
and \U$24850 ( \33038 , \33037 , \32756 );
or \U$24851 ( \33039 , \33027 , \33038 );
and \U$24853 ( \33040 , \33039 , 1'b1 );
or \U$24855 ( \33041 , \33040 , 1'b0 );
buf \U$24856 ( \33042 , \33041 );
_DC r23a1a_GF_IsGateDCbyConstraint ( \33043_nR23a1a , \33042 , \21944 );
buf \U$24857 ( \33044 , \33043_nR23a1a );
not \U$24858 ( \33045 , \32666 );
and \U$24859 ( \33046 , RIe0a6fa0_5705, \33045 );
not \U$24860 ( \33047 , RIe0a6fa0_5705);
or \U$24861 ( \33048 , \33047 , \32779 );
buf \U$24862 ( \33049 , RIb885928_52);
buf \U$24863 ( \33050 , \33049 );
and \U$24864 ( \33051 , \32781 , \33050 );
buf \U$24865 ( \33052 , \22500 );
buf \U$24866 ( \33053 , \32684 );
not \U$24867 ( \33054 , \33053 );
and \U$24868 ( \33055 , \33052 , \33054 );
nor \U$24869 ( \33056 , \33051 , \33055 );
nand \U$24870 ( \33057 , \33048 , \33056 );
and \U$24871 ( \33058 , \33057 , \32666 );
or \U$24872 ( \33059 , \33046 , \33058 );
and \U$24874 ( \33060 , \33059 , 1'b1 );
or \U$24876 ( \33061 , \33060 , 1'b0 );
buf \U$24877 ( \33062 , \33061 );
_DC r23a1c_GF_IsGateDCbyConstraint ( \33063_nR23a1c , \33062 , \21944 );
buf \U$24878 ( \33064 , \33063_nR23a1c );
not \U$24879 ( \33065 , \32756 );
and \U$24880 ( \33066 , RIe0ac310_5706, \33065 );
not \U$24881 ( \33067 , RIe0ac310_5706);
or \U$24882 ( \33068 , \33067 , \32949 );
buf \U$24883 ( \33069 , \22518 );
and \U$24884 ( \33070 , \32739 , \33069 );
buf \U$24885 ( \33071 , \22521 );
not \U$24886 ( \33072 , \32723 );
and \U$24887 ( \33073 , \33071 , \33072 );
nor \U$24888 ( \33074 , \33070 , \33073 );
nand \U$24889 ( \33075 , \33068 , \33074 );
and \U$24890 ( \33076 , \33075 , \32756 );
or \U$24891 ( \33077 , \33066 , \33076 );
and \U$24893 ( \33078 , \33077 , 1'b1 );
or \U$24895 ( \33079 , \33078 , 1'b0 );
buf \U$24896 ( \33080 , \33079 );
_DC r23a1e_GF_IsGateDCbyConstraint ( \33081_nR23a1e , \33080 , \21944 );
buf \U$24897 ( \33082 , \33081_nR23a1e );
not \U$24898 ( \33083 , \32666 );
and \U$24899 ( \33084 , RIe0b16f8_5707, \33083 );
not \U$24900 ( \33085 , RIe0b16f8_5707);
or \U$24901 ( \33086 , \33085 , \32686 );
buf \U$24902 ( \33087 , RIb885a18_50);
buf \U$24903 ( \33088 , \33087 );
and \U$24904 ( \33089 , \32717 , \33088 );
buf \U$24905 ( \33090 , RIb829498_218);
buf \U$24906 ( \33091 , \33090 );
not \U$24907 ( \33092 , \32685 );
and \U$24908 ( \33093 , \33091 , \33092 );
nor \U$24909 ( \33094 , \33089 , \33093 );
nand \U$24910 ( \33095 , \33086 , \33094 );
and \U$24911 ( \33096 , \33095 , \32666 );
or \U$24912 ( \33097 , \33084 , \33096 );
and \U$24914 ( \33098 , \33097 , 1'b1 );
or \U$24916 ( \33099 , \33098 , 1'b0 );
buf \U$24917 ( \33100 , \33099 );
_DC r23a20_GF_IsGateDCbyConstraint ( \33101_nR23a20 , \33100 , \21944 );
buf \U$24918 ( \33102 , \33101_nR23a20 );
not \U$24919 ( \33103 , \32666 );
and \U$24920 ( \33104 , RIe0b9240_5708, \33103 );
not \U$24921 ( \33105 , RIe0b9240_5708);
or \U$24922 ( \33106 , \33105 , \32868 );
buf \U$24923 ( \33107 , \27795 );
and \U$24924 ( \33108 , \32739 , \33107 );
buf \U$24925 ( \33109 , RIb829510_217);
buf \U$24926 ( \33110 , \33109 );
not \U$24927 ( \33111 , \33053 );
and \U$24928 ( \33112 , \33110 , \33111 );
nor \U$24929 ( \33113 , \33108 , \33112 );
nand \U$24930 ( \33114 , \33106 , \33113 );
and \U$24931 ( \33115 , \33114 , \32666 );
or \U$24932 ( \33116 , \33104 , \33115 );
and \U$24934 ( \33117 , \33116 , 1'b1 );
or \U$24936 ( \33118 , \33117 , 1'b0 );
buf \U$24937 ( \33119 , \33118 );
_DC r23a24_GF_IsGateDCbyConstraint ( \33120_nR23a24 , \33119 , \21944 );
buf \U$24938 ( \33121 , \33120_nR23a24 );
not \U$24939 ( \33122 , \32756 );
and \U$24940 ( \33123 , RIe0bf438_5709, \33122 );
not \U$24941 ( \33124 , RIe0bf438_5709);
or \U$24942 ( \33125 , \33124 , \32889 );
buf \U$24943 ( \33126 , RIb885b08_48);
and \U$24944 ( \33127 , \32739 , \33126 );
buf \U$24945 ( \33128 , RIb829588_216);
buf \U$24946 ( \33129 , \33128 );
not \U$24947 ( \33130 , \32811 );
and \U$24948 ( \33131 , \33129 , \33130 );
nor \U$24949 ( \33132 , \33127 , \33131 );
nand \U$24950 ( \33133 , \33125 , \33132 );
and \U$24951 ( \33134 , \33133 , \32756 );
or \U$24952 ( \33135 , \33123 , \33134 );
and \U$24954 ( \33136 , \33135 , 1'b1 );
or \U$24956 ( \33137 , \33136 , 1'b0 );
buf \U$24957 ( \33138 , \33137 );
_DC r23a26_GF_IsGateDCbyConstraint ( \33139_nR23a26 , \33138 , \21944 );
buf \U$24958 ( \33140 , \33139_nR23a26 );
not \U$24959 ( \33141 , \32756 );
and \U$24960 ( \33142 , RIe0c4730_5710, \33141 );
not \U$24961 ( \33143 , RIe0c4730_5710);
or \U$24962 ( \33144 , \33143 , \32686 );
buf \U$24963 ( \33145 , RIb885b80_47);
buf \U$24964 ( \33146 , \33145 );
and \U$24965 ( \33147 , \32739 , \33146 );
buf \U$24966 ( \33148 , RIb829600_215);
buf \U$24967 ( \33149 , \33148 );
not \U$24968 ( \33150 , \32852 );
and \U$24969 ( \33151 , \33149 , \33150 );
nor \U$24970 ( \33152 , \33147 , \33151 );
nand \U$24971 ( \33153 , \33144 , \33152 );
and \U$24972 ( \33154 , \33153 , \32756 );
or \U$24973 ( \33155 , \33142 , \33154 );
and \U$24975 ( \33156 , \33155 , 1'b1 );
or \U$24977 ( \33157 , \33156 , 1'b0 );
buf \U$24978 ( \33158 , \33157 );
_DC r23a28_GF_IsGateDCbyConstraint ( \33159_nR23a28 , \33158 , \21944 );
buf \U$24979 ( \33160 , \33159_nR23a28 );
not \U$24980 ( \33161 , \32666 );
and \U$24981 ( \33162 , RIe0cb0a8_5711, \33161 );
not \U$24982 ( \33163 , RIe0cb0a8_5711);
or \U$24983 ( \33164 , \33163 , \32715 );
buf \U$24984 ( \33165 , \22618 );
and \U$24985 ( \33166 , \32717 , \33165 );
buf \U$24986 ( \33167 , \22621 );
not \U$24987 ( \33168 , \32874 );
and \U$24988 ( \33169 , \33167 , \33168 );
nor \U$24989 ( \33170 , \33166 , \33169 );
nand \U$24990 ( \33171 , \33164 , \33170 );
and \U$24991 ( \33172 , \33171 , \32666 );
or \U$24992 ( \33173 , \33162 , \33172 );
and \U$24994 ( \33174 , \33173 , 1'b1 );
or \U$24996 ( \33175 , \33174 , 1'b0 );
buf \U$24997 ( \33176 , \33175 );
_DC r23a2a_GF_IsGateDCbyConstraint ( \33177_nR23a2a , \33176 , \21944 );
buf \U$24998 ( \33178 , \33177_nR23a2a );
not \U$24999 ( \33179 , \32666 );
and \U$25000 ( \33180 , RIe0d0df0_5712, \33179 );
not \U$25001 ( \33181 , RIe0d0df0_5712);
or \U$25002 ( \33182 , \33181 , \32868 );
buf \U$25003 ( \33183 , RIb885c70_45);
buf \U$25004 ( \33184 , \33183 );
and \U$25005 ( \33185 , \32739 , \33184 );
buf \U$25006 ( \33186 , RIb8296f0_213);
buf \U$25007 ( \33187 , \33186 );
not \U$25008 ( \33188 , \32811 );
and \U$25009 ( \33189 , \33187 , \33188 );
nor \U$25010 ( \33190 , \33185 , \33189 );
nand \U$25011 ( \33191 , \33182 , \33190 );
and \U$25012 ( \33192 , \33191 , \32666 );
or \U$25013 ( \33193 , \33180 , \33192 );
and \U$25015 ( \33194 , \33193 , 1'b1 );
or \U$25017 ( \33195 , \33194 , 1'b0 );
buf \U$25018 ( \33196 , \33195 );
_DC r23a2c_GF_IsGateDCbyConstraint ( \33197_nR23a2c , \33196 , \21944 );
buf \U$25019 ( \33198 , \33197_nR23a2c );
not \U$25020 ( \33199 , \32666 );
and \U$25021 ( \33200 , RIe0d8aa0_5713, \33199 );
not \U$25022 ( \33201 , RIe0d8aa0_5713);
or \U$25023 ( \33202 , \33201 , \32889 );
buf \U$25024 ( \33203 , \22659 );
and \U$25025 ( \33204 , \32739 , \33203 );
buf \U$25026 ( \33205 , \22662 );
not \U$25027 ( \33206 , \32852 );
and \U$25028 ( \33207 , \33205 , \33206 );
nor \U$25029 ( \33208 , \33204 , \33207 );
nand \U$25030 ( \33209 , \33202 , \33208 );
and \U$25031 ( \33210 , \33209 , \32666 );
or \U$25032 ( \33211 , \33200 , \33210 );
and \U$25034 ( \33212 , \33211 , 1'b1 );
or \U$25036 ( \33213 , \33212 , 1'b0 );
buf \U$25037 ( \33214 , \33213 );
_DC r23a2e_GF_IsGateDCbyConstraint ( \33215_nR23a2e , \33214 , \21944 );
buf \U$25038 ( \33216 , \33215_nR23a2e );
buf \U$25039 ( \33217 , \32665 );
buf \U$25040 ( \33218 , \33217 );
not \U$25041 ( \33219 , \33218 );
and \U$25042 ( \33220 , RIe0de608_5714, \33219 );
not \U$25043 ( \33221 , RIe0de608_5714);
or \U$25044 ( \33222 , \33221 , \32968 );
buf \U$25045 ( \33223 , \22680 );
and \U$25046 ( \33224 , \32739 , \33223 );
buf \U$25047 ( \33225 , RIb82db60_211);
buf \U$25048 ( \33226 , \33225 );
not \U$25049 ( \33227 , \33053 );
and \U$25050 ( \33228 , \33226 , \33227 );
nor \U$25051 ( \33229 , \33224 , \33228 );
nand \U$25052 ( \33230 , \33222 , \33229 );
and \U$25053 ( \33231 , \33230 , \33218 );
or \U$25054 ( \33232 , \33220 , \33231 );
and \U$25056 ( \33233 , \33232 , 1'b1 );
or \U$25058 ( \33234 , \33233 , 1'b0 );
buf \U$25059 ( \33235 , \33234 );
_DC r23a30_GF_IsGateDCbyConstraint ( \33236_nR23a30 , \33235 , \21944 );
buf \U$25060 ( \33237 , \33236_nR23a30 );
not \U$25061 ( \33238 , \32756 );
and \U$25062 ( \33239 , RIe0e5ca0_5715, \33238 );
not \U$25063 ( \33240 , RIe0e5ca0_5715);
or \U$25064 ( \33241 , \33240 , \32801 );
buf \U$25065 ( \33242 , \22700 );
and \U$25066 ( \33243 , \32739 , \33242 );
buf \U$25067 ( \33244 , RIb82dbd8_210);
buf \U$25068 ( \33245 , \33244 );
not \U$25069 ( \33246 , \32974 );
and \U$25070 ( \33247 , \33245 , \33246 );
nor \U$25071 ( \33248 , \33243 , \33247 );
nand \U$25072 ( \33249 , \33241 , \33248 );
and \U$25073 ( \33250 , \33249 , \32756 );
or \U$25074 ( \33251 , \33239 , \33250 );
and \U$25076 ( \33252 , \33251 , 1'b1 );
or \U$25078 ( \33253 , \33252 , 1'b0 );
buf \U$25079 ( \33254 , \33253 );
_DC r23a32_GF_IsGateDCbyConstraint ( \33255_nR23a32 , \33254 , \21944 );
buf \U$25080 ( \33256 , \33255_nR23a32 );
buf \U$25081 ( \33257 , \32755 );
not \U$25082 ( \33258 , \33257 );
and \U$25083 ( \33259 , RIe0eb358_5716, \33258 );
not \U$25084 ( \33260 , RIe0eb358_5716);
or \U$25085 ( \33261 , \33260 , \32968 );
buf \U$25086 ( \33262 , RIb885e50_41);
and \U$25087 ( \33263 , \32690 , \33262 );
buf \U$25088 ( \33264 , RIb82dc50_209);
buf \U$25089 ( \33265 , \33264 );
not \U$25090 ( \33266 , \32895 );
and \U$25091 ( \33267 , \33265 , \33266 );
nor \U$25092 ( \33268 , \33263 , \33267 );
nand \U$25093 ( \33269 , \33261 , \33268 );
and \U$25094 ( \33270 , \33269 , \33257 );
or \U$25095 ( \33271 , \33259 , \33270 );
and \U$25097 ( \33272 , \33271 , 1'b1 );
or \U$25099 ( \33273 , \33272 , 1'b0 );
buf \U$25100 ( \33274 , \33273 );
_DC r23a34_GF_IsGateDCbyConstraint ( \33275_nR23a34 , \33274 , \21944 );
buf \U$25101 ( \33276 , \33275_nR23a34 );
not \U$25102 ( \33277 , \32666 );
and \U$25103 ( \33278 , RIe0ef138_5717, \33277 );
not \U$25104 ( \33279 , RIe0ef138_5717);
or \U$25105 ( \33280 , \33279 , \32801 );
buf \U$25106 ( \33281 , RIb885ec8_40);
and \U$25107 ( \33282 , \32717 , \33281 );
buf \U$25108 ( \33283 , RIb82dcc8_208);
buf \U$25109 ( \33284 , \33283 );
not \U$25110 ( \33285 , \32713 );
and \U$25111 ( \33286 , \33284 , \33285 );
nor \U$25112 ( \33287 , \33282 , \33286 );
nand \U$25113 ( \33288 , \33280 , \33287 );
and \U$25114 ( \33289 , \33288 , \32666 );
or \U$25115 ( \33290 , \33278 , \33289 );
and \U$25117 ( \33291 , \33290 , 1'b1 );
or \U$25119 ( \33292 , \33291 , 1'b0 );
buf \U$25120 ( \33293 , \33292 );
_DC r23a36_GF_IsGateDCbyConstraint ( \33294_nR23a36 , \33293 , \21944 );
buf \U$25121 ( \33295 , \33294_nR23a36 );
buf \U$25122 ( \33296 , \32665 );
buf \U$25123 ( \33297 , \33296 );
not \U$25124 ( \33298 , \33297 );
and \U$25125 ( \33299 , RIe0f3bc0_5718, \33298 );
not \U$25126 ( \33300 , RIe0f3bc0_5718);
or \U$25127 ( \33301 , \33300 , \32910 );
buf \U$25128 ( \33302 , RIb885f40_39);
buf \U$25129 ( \33303 , \33302 );
and \U$25130 ( \33304 , \32717 , \33303 );
buf \U$25131 ( \33305 , \22765 );
not \U$25132 ( \33306 , \32723 );
and \U$25133 ( \33307 , \33305 , \33306 );
nor \U$25134 ( \33308 , \33304 , \33307 );
nand \U$25135 ( \33309 , \33301 , \33308 );
and \U$25136 ( \33310 , \33309 , \33297 );
or \U$25137 ( \33311 , \33299 , \33310 );
and \U$25139 ( \33312 , \33311 , 1'b1 );
or \U$25141 ( \33313 , \33312 , 1'b0 );
buf \U$25142 ( \33314 , \33313 );
_DC r23a3a_GF_IsGateDCbyConstraint ( \33315_nR23a3a , \33314 , \21944 );
buf \U$25143 ( \33316 , \33315_nR23a3a );
not \U$25144 ( \33317 , \33297 );
and \U$25145 ( \33318 , RIe0f8300_5719, \33317 );
not \U$25146 ( \33319 , RIe0f8300_5719);
or \U$25147 ( \33320 , \33319 , \32688 );
buf \U$25148 ( \33321 , RIb885fb8_38);
and \U$25149 ( \33322 , \32717 , \33321 );
buf \U$25150 ( \33323 , RIb82ddb8_206);
buf \U$25151 ( \33324 , \33323 );
not \U$25152 ( \33325 , \33053 );
and \U$25153 ( \33326 , \33324 , \33325 );
nor \U$25154 ( \33327 , \33322 , \33326 );
nand \U$25155 ( \33328 , \33320 , \33327 );
and \U$25156 ( \33329 , \33328 , \33297 );
or \U$25157 ( \33330 , \33318 , \33329 );
and \U$25159 ( \33331 , \33330 , 1'b1 );
or \U$25161 ( \33332 , \33331 , 1'b0 );
buf \U$25162 ( \33333 , \33332 );
_DC r23a3c_GF_IsGateDCbyConstraint ( \33334_nR23a3c , \33333 , \21944 );
buf \U$25163 ( \33335 , \33334_nR23a3c );
buf \U$25164 ( \33336 , \33217 );
not \U$25165 ( \33337 , \33336 );
and \U$25166 ( \33338 , RIe0ff380_5720, \33337 );
not \U$25167 ( \33339 , RIe0ff380_5720);
or \U$25168 ( \33340 , \33339 , \32910 );
buf \U$25169 ( \33341 , \22802 );
and \U$25170 ( \33342 , \32739 , \33341 );
buf \U$25171 ( \33343 , RIb82de30_205);
buf \U$25172 ( \33344 , \33343 );
not \U$25173 ( \33345 , \32874 );
and \U$25174 ( \33346 , \33344 , \33345 );
nor \U$25175 ( \33347 , \33342 , \33346 );
nand \U$25176 ( \33348 , \33340 , \33347 );
and \U$25177 ( \33349 , \33348 , \33336 );
or \U$25178 ( \33350 , \33338 , \33349 );
and \U$25180 ( \33351 , \33350 , 1'b1 );
or \U$25182 ( \33352 , \33351 , 1'b0 );
buf \U$25183 ( \33353 , \33352 );
_DC r23a3e_GF_IsGateDCbyConstraint ( \33354_nR23a3e , \33353 , \21944 );
buf \U$25184 ( \33355 , \33354_nR23a3e );
not \U$25185 ( \33356 , \33257 );
and \U$25186 ( \33357 , RIe103430_5721, \33356 );
not \U$25187 ( \33358 , RIe103430_5721);
or \U$25188 ( \33359 , \33358 , \32779 );
buf \U$25189 ( \33360 , RIb8860a8_36);
and \U$25190 ( \33361 , \32717 , \33360 );
buf \U$25191 ( \33362 , RIb832228_204);
buf \U$25192 ( \33363 , \33362 );
not \U$25193 ( \33364 , \32974 );
and \U$25194 ( \33365 , \33363 , \33364 );
nor \U$25195 ( \33366 , \33361 , \33365 );
nand \U$25196 ( \33367 , \33359 , \33366 );
and \U$25197 ( \33368 , \33367 , \33257 );
or \U$25198 ( \33369 , \33357 , \33368 );
and \U$25200 ( \33370 , \33369 , 1'b1 );
or \U$25202 ( \33371 , \33370 , 1'b0 );
buf \U$25203 ( \33372 , \33371 );
_DC r23a40_GF_IsGateDCbyConstraint ( \33373_nR23a40 , \33372 , \21944 );
buf \U$25204 ( \33374 , \33373_nR23a40 );
not \U$25205 ( \33375 , \33297 );
and \U$25206 ( \33376 , RIdfce868_5722, \33375 );
not \U$25207 ( \33377 , RIdfce868_5722);
or \U$25208 ( \33378 , \33377 , \32949 );
buf \U$25209 ( \33379 , RIb886120_35);
and \U$25210 ( \33380 , \32717 , \33379 );
buf \U$25211 ( \33381 , RIb8322a0_203);
buf \U$25212 ( \33382 , \33381 );
not \U$25213 ( \33383 , \32811 );
and \U$25214 ( \33384 , \33382 , \33383 );
nor \U$25215 ( \33385 , \33380 , \33384 );
nand \U$25216 ( \33386 , \33378 , \33385 );
and \U$25217 ( \33387 , \33386 , \33297 );
or \U$25218 ( \33388 , \33376 , \33387 );
and \U$25220 ( \33389 , \33388 , 1'b1 );
or \U$25222 ( \33390 , \33389 , 1'b0 );
buf \U$25223 ( \33391 , \33390 );
_DC r23a42_GF_IsGateDCbyConstraint ( \33392_nR23a42 , \33391 , \21944 );
buf \U$25224 ( \33393 , \33392_nR23a42 );
not \U$25225 ( \33394 , \32666 );
and \U$25226 ( \33395 , RIdfc9fc0_5723, \33394 );
not \U$25227 ( \33396 , RIdfc9fc0_5723);
or \U$25228 ( \33397 , \33396 , \32686 );
buf \U$25229 ( \33398 , RIb886198_34);
buf \U$25230 ( \33399 , \33398 );
and \U$25231 ( \33400 , \32739 , \33399 );
buf \U$25232 ( \33401 , RIb832318_202);
buf \U$25233 ( \33402 , \33401 );
not \U$25234 ( \33403 , \32811 );
and \U$25235 ( \33404 , \33402 , \33403 );
nor \U$25236 ( \33405 , \33400 , \33404 );
nand \U$25237 ( \33406 , \33397 , \33405 );
and \U$25238 ( \33407 , \33406 , \32666 );
or \U$25239 ( \33408 , \33395 , \33407 );
and \U$25241 ( \33409 , \33408 , 1'b1 );
or \U$25243 ( \33410 , \33409 , 1'b0 );
buf \U$25244 ( \33411 , \33410 );
_DC r23a44_GF_IsGateDCbyConstraint ( \33412_nR23a44 , \33411 , \21944 );
buf \U$25245 ( \33413 , \33412_nR23a44 );
not \U$25246 ( \33414 , \33297 );
and \U$25247 ( \33415 , RIdfc6000_5724, \33414 );
not \U$25248 ( \33416 , RIdfc6000_5724);
or \U$25249 ( \33417 , \33416 , \32715 );
buf \U$25250 ( \33418 , RIb886210_33);
buf \U$25251 ( \33419 , \33418 );
and \U$25252 ( \33420 , \32717 , \33419 );
buf \U$25253 ( \33421 , RIb832390_201);
buf \U$25254 ( \33422 , \33421 );
not \U$25255 ( \33423 , \32852 );
and \U$25256 ( \33424 , \33422 , \33423 );
nor \U$25257 ( \33425 , \33420 , \33424 );
nand \U$25258 ( \33426 , \33417 , \33425 );
and \U$25259 ( \33427 , \33426 , \33297 );
or \U$25260 ( \33428 , \33415 , \33427 );
and \U$25262 ( \33429 , \33428 , 1'b1 );
or \U$25264 ( \33430 , \33429 , 1'b0 );
buf \U$25265 ( \33431 , \33430 );
_DC r23a46_GF_IsGateDCbyConstraint ( \33432_nR23a46 , \33431 , \21944 );
buf \U$25266 ( \33433 , \33432_nR23a46 );
not \U$25267 ( \33434 , \33297 );
and \U$25268 ( \33435 , RIdfc1410_5725, \33434 );
not \U$25269 ( \33436 , RIdfc1410_5725);
or \U$25270 ( \33437 , \33436 , \32779 );
buf \U$25271 ( \33438 , \22904 );
and \U$25272 ( \33439 , \32739 , \33438 );
buf \U$25273 ( \33440 , \22907 );
not \U$25274 ( \33441 , \32874 );
and \U$25275 ( \33442 , \33440 , \33441 );
nor \U$25276 ( \33443 , \33439 , \33442 );
nand \U$25277 ( \33444 , \33437 , \33443 );
and \U$25278 ( \33445 , \33444 , \33297 );
or \U$25279 ( \33446 , \33435 , \33445 );
and \U$25281 ( \33447 , \33446 , 1'b1 );
or \U$25283 ( \33448 , \33447 , 1'b0 );
buf \U$25284 ( \33449 , \33448 );
_DC r23a48_GF_IsGateDCbyConstraint ( \33450_nR23a48 , \33449 , \21944 );
buf \U$25285 ( \33451 , \33450_nR23a48 );
not \U$25286 ( \33452 , \32666 );
and \U$25287 ( \33453 , RIdfbcc58_5726, \33452 );
not \U$25288 ( \33454 , RIdfbcc58_5726);
or \U$25289 ( \33455 , \33454 , \32949 );
buf \U$25290 ( \33456 , \22924 );
and \U$25291 ( \33457 , \32781 , \33456 );
buf \U$25292 ( \33458 , RIb832480_199);
buf \U$25293 ( \33459 , \33458 );
not \U$25294 ( \33460 , \32974 );
and \U$25295 ( \33461 , \33459 , \33460 );
nor \U$25296 ( \33462 , \33457 , \33461 );
nand \U$25297 ( \33463 , \33455 , \33462 );
and \U$25298 ( \33464 , \33463 , \32666 );
or \U$25299 ( \33465 , \33453 , \33464 );
and \U$25301 ( \33466 , \33465 , 1'b1 );
or \U$25303 ( \33467 , \33466 , 1'b0 );
buf \U$25304 ( \33468 , \33467 );
_DC r23a4a_GF_IsGateDCbyConstraint ( \33469_nR23a4a , \33468 , \21944 );
buf \U$25305 ( \33470 , \33469_nR23a4a );
not \U$25306 ( \33471 , \33257 );
and \U$25307 ( \33472 , RIe082f10_5727, \33471 );
not \U$25308 ( \33473 , RIe082f10_5727);
or \U$25309 ( \33474 , \33473 , \32686 );
buf \U$25310 ( \33475 , \22944 );
and \U$25311 ( \33476 , \32690 , \33475 );
buf \U$25312 ( \33477 , RIb8324f8_198);
buf \U$25313 ( \33478 , \33477 );
not \U$25314 ( \33479 , \32895 );
and \U$25315 ( \33480 , \33478 , \33479 );
nor \U$25316 ( \33481 , \33476 , \33480 );
nand \U$25317 ( \33482 , \33474 , \33481 );
and \U$25318 ( \33483 , \33482 , \33257 );
or \U$25319 ( \33484 , \33472 , \33483 );
and \U$25321 ( \33485 , \33484 , 1'b1 );
or \U$25323 ( \33486 , \33485 , 1'b0 );
buf \U$25324 ( \33487 , \33486 );
_DC r23a4c_GF_IsGateDCbyConstraint ( \33488_nR23a4c , \33487 , \21944 );
buf \U$25325 ( \33489 , \33488_nR23a4c );
not \U$25326 ( \33490 , \33257 );
and \U$25327 ( \33491 , RIe0800a8_5728, \33490 );
not \U$25328 ( \33492 , RIe0800a8_5728);
or \U$25329 ( \33493 , \33492 , \32868 );
buf \U$25330 ( \33494 , RIb8863f0_29);
and \U$25331 ( \33495 , \32781 , \33494 );
buf \U$25332 ( \33496 , RIb832570_197);
buf \U$25333 ( \33497 , \33496 );
not \U$25334 ( \33498 , \32895 );
and \U$25335 ( \33499 , \33497 , \33498 );
nor \U$25336 ( \33500 , \33495 , \33499 );
nand \U$25337 ( \33501 , \33493 , \33500 );
and \U$25338 ( \33502 , \33501 , \33257 );
or \U$25339 ( \33503 , \33491 , \33502 );
and \U$25341 ( \33504 , \33503 , 1'b1 );
or \U$25343 ( \33505 , \33504 , 1'b0 );
buf \U$25344 ( \33506 , \33505 );
_DC r23a50_GF_IsGateDCbyConstraint ( \33507_nR23a50 , \33506 , \21944 );
buf \U$25345 ( \33508 , \33507_nR23a50 );
not \U$25346 ( \33509 , \32666 );
and \U$25347 ( \33510 , RIe07bd28_5729, \33509 );
not \U$25348 ( \33511 , RIe07bd28_5729);
or \U$25349 ( \33512 , \33511 , \32889 );
buf \U$25350 ( \33513 , RIb886468_28);
buf \U$25351 ( \33514 , \33513 );
and \U$25352 ( \33515 , \32690 , \33514 );
buf \U$25353 ( \33516 , RIb8383a8_196);
buf \U$25354 ( \33517 , \33516 );
not \U$25355 ( \33518 , \32713 );
and \U$25356 ( \33519 , \33517 , \33518 );
nor \U$25357 ( \33520 , \33515 , \33519 );
nand \U$25358 ( \33521 , \33512 , \33520 );
and \U$25359 ( \33522 , \33521 , \32666 );
or \U$25360 ( \33523 , \33510 , \33522 );
and \U$25362 ( \33524 , \33523 , 1'b1 );
or \U$25364 ( \33525 , \33524 , 1'b0 );
buf \U$25365 ( \33526 , \33525 );
_DC r23a52_GF_IsGateDCbyConstraint ( \33527_nR23a52 , \33526 , \21944 );
buf \U$25366 ( \33528 , \33527_nR23a52 );
not \U$25367 ( \33529 , \33257 );
and \U$25368 ( \33530 , RIe078ec0_5730, \33529 );
not \U$25369 ( \33531 , RIe078ec0_5730);
or \U$25370 ( \33532 , \33531 , \32968 );
buf \U$25371 ( \33533 , RIb8864e0_27);
buf \U$25372 ( \33534 , \33533 );
and \U$25373 ( \33535 , \32781 , \33534 );
buf \U$25374 ( \33536 , RIb838420_195);
buf \U$25375 ( \33537 , \33536 );
not \U$25376 ( \33538 , \32852 );
and \U$25377 ( \33539 , \33537 , \33538 );
nor \U$25378 ( \33540 , \33535 , \33539 );
nand \U$25379 ( \33541 , \33532 , \33540 );
and \U$25380 ( \33542 , \33541 , \33257 );
or \U$25381 ( \33543 , \33530 , \33542 );
and \U$25383 ( \33544 , \33543 , 1'b1 );
or \U$25385 ( \33545 , \33544 , 1'b0 );
buf \U$25386 ( \33546 , \33545 );
_DC r23a54_GF_IsGateDCbyConstraint ( \33547_nR23a54 , \33546 , \21944 );
buf \U$25387 ( \33548 , \33547_nR23a54 );
not \U$25388 ( \33549 , \33297 );
and \U$25389 ( \33550 , RIe075ab8_5731, \33549 );
not \U$25390 ( \33551 , RIe075ab8_5731);
or \U$25391 ( \33552 , \33551 , \32801 );
buf \U$25392 ( \33553 , RIb886558_26);
and \U$25393 ( \33554 , \32739 , \33553 );
buf \U$25394 ( \33555 , RIb838498_194);
buf \U$25395 ( \33556 , \33555 );
not \U$25396 ( \33557 , \32685 );
and \U$25397 ( \33558 , \33556 , \33557 );
nor \U$25398 ( \33559 , \33554 , \33558 );
nand \U$25399 ( \33560 , \33552 , \33559 );
and \U$25400 ( \33561 , \33560 , \33297 );
or \U$25401 ( \33562 , \33550 , \33561 );
and \U$25403 ( \33563 , \33562 , 1'b1 );
or \U$25405 ( \33564 , \33563 , 1'b0 );
buf \U$25406 ( \33565 , \33564 );
_DC r23a56_GF_IsGateDCbyConstraint ( \33566_nR23a56 , \33565 , \21944 );
buf \U$25407 ( \33567 , \33566_nR23a56 );
buf \U$25408 ( \33568 , \32665 );
buf \U$25409 ( \33569 , \33568 );
not \U$25410 ( \33570 , \33569 );
and \U$25411 ( \33571 , RIe071f18_5732, \33570 );
not \U$25412 ( \33572 , RIe071f18_5732);
or \U$25413 ( \33573 , \33572 , \32688 );
buf \U$25414 ( \33574 , \23044 );
and \U$25415 ( \33575 , \32781 , \33574 );
buf \U$25416 ( \33576 , \23047 );
not \U$25417 ( \33577 , \32723 );
and \U$25418 ( \33578 , \33576 , \33577 );
nor \U$25419 ( \33579 , \33575 , \33578 );
nand \U$25420 ( \33580 , \33573 , \33579 );
and \U$25421 ( \33581 , \33580 , \33569 );
or \U$25422 ( \33582 , \33571 , \33581 );
and \U$25424 ( \33583 , \33582 , 1'b1 );
or \U$25426 ( \33584 , \33583 , 1'b0 );
buf \U$25427 ( \33585 , \33584 );
_DC r23a58_GF_IsGateDCbyConstraint ( \33586_nR23a58 , \33585 , \21944 );
buf \U$25428 ( \33587 , \33586_nR23a58 );
not \U$25429 ( \33588 , \33257 );
and \U$25430 ( \33589 , RIe06f308_5733, \33588 );
not \U$25431 ( \33590 , RIe06f308_5733);
or \U$25432 ( \33591 , \33590 , \32910 );
buf \U$25433 ( \33592 , \23064 );
and \U$25434 ( \33593 , \32739 , \33592 );
buf \U$25435 ( \33594 , \23067 );
not \U$25436 ( \33595 , \33053 );
and \U$25437 ( \33596 , \33594 , \33595 );
nor \U$25438 ( \33597 , \33593 , \33596 );
nand \U$25439 ( \33598 , \33591 , \33597 );
and \U$25440 ( \33599 , \33598 , \33257 );
or \U$25441 ( \33600 , \33589 , \33599 );
and \U$25443 ( \33601 , \33600 , 1'b1 );
or \U$25445 ( \33602 , \33601 , 1'b0 );
buf \U$25446 ( \33603 , \33602 );
_DC r23a5a_GF_IsGateDCbyConstraint ( \33604_nR23a5a , \33603 , \21944 );
buf \U$25447 ( \33605 , \33604_nR23a5a );
not \U$25448 ( \33606 , \33297 );
and \U$25449 ( \33607 , RIe06b0f0_5734, \33606 );
not \U$25450 ( \33608 , RIe06b0f0_5734);
or \U$25451 ( \33609 , \33608 , \32868 );
buf \U$25452 ( \33610 , \23084 );
and \U$25453 ( \33611 , \32739 , \33610 );
buf \U$25454 ( \33612 , \23087 );
not \U$25455 ( \33613 , \32811 );
and \U$25456 ( \33614 , \33612 , \33613 );
nor \U$25457 ( \33615 , \33611 , \33614 );
nand \U$25458 ( \33616 , \33609 , \33615 );
and \U$25459 ( \33617 , \33616 , \33297 );
or \U$25460 ( \33618 , \33607 , \33617 );
and \U$25462 ( \33619 , \33618 , 1'b1 );
or \U$25464 ( \33620 , \33619 , 1'b0 );
buf \U$25465 ( \33621 , \33620 );
_DC r23a5c_GF_IsGateDCbyConstraint ( \33622_nR23a5c , \33621 , \21944 );
buf \U$25466 ( \33623 , \33622_nR23a5c );
not \U$25467 ( \33624 , \33569 );
and \U$25468 ( \33625 , RIe067928_5735, \33624 );
not \U$25469 ( \33626 , RIe067928_5735);
or \U$25470 ( \33627 , \33626 , \32889 );
buf \U$25471 ( \33628 , RIb886738_22);
buf \U$25472 ( \33629 , \33628 );
and \U$25473 ( \33630 , \32717 , \33629 );
buf \U$25474 ( \33631 , RIb838678_190);
buf \U$25475 ( \33632 , \33631 );
not \U$25476 ( \33633 , \32852 );
and \U$25477 ( \33634 , \33632 , \33633 );
nor \U$25478 ( \33635 , \33630 , \33634 );
nand \U$25479 ( \33636 , \33627 , \33635 );
and \U$25480 ( \33637 , \33636 , \33569 );
or \U$25481 ( \33638 , \33625 , \33637 );
and \U$25483 ( \33639 , \33638 , 1'b1 );
or \U$25485 ( \33640 , \33639 , 1'b0 );
buf \U$25486 ( \33641 , \33640 );
_DC r23a5e_GF_IsGateDCbyConstraint ( \33642_nR23a5e , \33641 , \21944 );
buf \U$25487 ( \33643 , \33642_nR23a5e );
not \U$25488 ( \33644 , \33297 );
and \U$25489 ( \33645 , RIe0608a8_5736, \33644 );
not \U$25490 ( \33646 , RIe0608a8_5736);
or \U$25491 ( \33647 , \33646 , \32968 );
buf \U$25492 ( \33648 , \23124 );
and \U$25493 ( \33649 , \32781 , \33648 );
buf \U$25494 ( \33650 , RIb8386f0_189);
buf \U$25495 ( \33651 , \33650 );
not \U$25496 ( \33652 , \32874 );
and \U$25497 ( \33653 , \33651 , \33652 );
nor \U$25498 ( \33654 , \33649 , \33653 );
nand \U$25499 ( \33655 , \33647 , \33654 );
and \U$25500 ( \33656 , \33655 , \33297 );
or \U$25501 ( \33657 , \33645 , \33656 );
and \U$25503 ( \33658 , \33657 , 1'b1 );
or \U$25505 ( \33659 , \33658 , 1'b0 );
buf \U$25506 ( \33660 , \33659 );
_DC r23a60_GF_IsGateDCbyConstraint ( \33661_nR23a60 , \33660 , \21944 );
buf \U$25507 ( \33662 , \33661_nR23a60 );
not \U$25508 ( \33663 , \33297 );
and \U$25509 ( \33664 , RIe05a2f0_5737, \33663 );
not \U$25510 ( \33665 , RIe05a2f0_5737);
or \U$25511 ( \33666 , \33665 , \32801 );
buf \U$25512 ( \33667 , RIb886828_20);
buf \U$25513 ( \33668 , \33667 );
and \U$25514 ( \33669 , \32739 , \33668 );
buf \U$25515 ( \33670 , RIb838768_188);
buf \U$25516 ( \33671 , \33670 );
not \U$25517 ( \33672 , \32685 );
and \U$25518 ( \33673 , \33671 , \33672 );
nor \U$25519 ( \33674 , \33669 , \33673 );
nand \U$25520 ( \33675 , \33666 , \33674 );
and \U$25521 ( \33676 , \33675 , \33297 );
or \U$25522 ( \33677 , \33664 , \33676 );
and \U$25524 ( \33678 , \33677 , 1'b1 );
or \U$25526 ( \33679 , \33678 , 1'b0 );
buf \U$25527 ( \33680 , \33679 );
_DC r23a62_GF_IsGateDCbyConstraint ( \33681_nR23a62 , \33680 , \21944 );
buf \U$25528 ( \33682 , \33681_nR23a62 );
not \U$25529 ( \33683 , \33569 );
and \U$25530 ( \33684 , RIe0541e8_5738, \33683 );
not \U$25531 ( \33685 , RIe0541e8_5738);
or \U$25532 ( \33686 , \33685 , \32949 );
buf \U$25533 ( \33687 , RIb8868a0_19);
buf \U$25534 ( \33688 , \33687 );
and \U$25535 ( \33689 , \32690 , \33688 );
buf \U$25536 ( \33690 , RIb8387e0_187);
buf \U$25537 ( \33691 , \33690 );
not \U$25538 ( \33692 , \32874 );
and \U$25539 ( \33693 , \33691 , \33692 );
nor \U$25540 ( \33694 , \33689 , \33693 );
nand \U$25541 ( \33695 , \33686 , \33694 );
and \U$25542 ( \33696 , \33695 , \33569 );
or \U$25543 ( \33697 , \33684 , \33696 );
and \U$25545 ( \33698 , \33697 , 1'b1 );
or \U$25547 ( \33699 , \33698 , 1'b0 );
buf \U$25548 ( \33700 , \33699 );
_DC r23a66_GF_IsGateDCbyConstraint ( \33701_nR23a66 , \33700 , \21944 );
buf \U$25549 ( \33702 , \33701_nR23a66 );
not \U$25550 ( \33703 , \33257 );
and \U$25551 ( \33704 , RIe04bb60_5739, \33703 );
not \U$25552 ( \33705 , RIe04bb60_5739);
or \U$25553 ( \33706 , \33705 , \32686 );
buf \U$25554 ( \33707 , RIb886918_18);
and \U$25555 ( \33708 , \32781 , \33707 );
buf \U$25556 ( \33709 , \23186 );
not \U$25557 ( \33710 , \32974 );
and \U$25558 ( \33711 , \33709 , \33710 );
nor \U$25559 ( \33712 , \33708 , \33711 );
nand \U$25560 ( \33713 , \33706 , \33712 );
and \U$25561 ( \33714 , \33713 , \33257 );
or \U$25562 ( \33715 , \33704 , \33714 );
and \U$25564 ( \33716 , \33715 , 1'b1 );
or \U$25566 ( \33717 , \33716 , 1'b0 );
buf \U$25567 ( \33718 , \33717 );
_DC r23a68_GF_IsGateDCbyConstraint ( \33719_nR23a68 , \33718 , \21944 );
buf \U$25568 ( \33720 , \33719_nR23a68 );
not \U$25569 ( \33721 , \33257 );
and \U$25570 ( \33722 , RIe045a58_5740, \33721 );
not \U$25571 ( \33723 , RIe045a58_5740);
or \U$25572 ( \33724 , \33723 , \32715 );
buf \U$25573 ( \33725 , RIb886990_17);
and \U$25574 ( \33726 , \32690 , \33725 );
buf \U$25575 ( \33727 , RIb8388d0_185);
buf \U$25576 ( \33728 , \33727 );
not \U$25577 ( \33729 , \32895 );
and \U$25578 ( \33730 , \33728 , \33729 );
nor \U$25579 ( \33731 , \33726 , \33730 );
nand \U$25580 ( \33732 , \33724 , \33731 );
and \U$25581 ( \33733 , \33732 , \33257 );
or \U$25582 ( \33734 , \33722 , \33733 );
and \U$25584 ( \33735 , \33734 , 1'b1 );
or \U$25586 ( \33736 , \33735 , 1'b0 );
buf \U$25587 ( \33737 , \33736 );
_DC r23a6a_GF_IsGateDCbyConstraint ( \33738_nR23a6a , \33737 , \21944 );
buf \U$25588 ( \33739 , \33738_nR23a6a );
not \U$25589 ( \33740 , \33569 );
and \U$25590 ( \33741 , RIe03d3d0_5741, \33740 );
not \U$25591 ( \33742 , RIe03d3d0_5741);
or \U$25592 ( \33743 , \33742 , \32868 );
buf \U$25593 ( \33744 , \23223 );
and \U$25594 ( \33745 , \32717 , \33744 );
buf \U$25595 ( \33746 , \23226 );
not \U$25596 ( \33747 , \32713 );
and \U$25597 ( \33748 , \33746 , \33747 );
nor \U$25598 ( \33749 , \33745 , \33748 );
nand \U$25599 ( \33750 , \33743 , \33749 );
and \U$25600 ( \33751 , \33750 , \33569 );
or \U$25601 ( \33752 , \33741 , \33751 );
and \U$25603 ( \33753 , \33752 , 1'b1 );
or \U$25605 ( \33754 , \33753 , 1'b0 );
buf \U$25606 ( \33755 , \33754 );
_DC r23a6c_GF_IsGateDCbyConstraint ( \33756_nR23a6c , \33755 , \21944 );
buf \U$25607 ( \33757 , \33756_nR23a6c );
not \U$25608 ( \33758 , \33297 );
and \U$25609 ( \33759 , RIde1d908_5742, \33758 );
not \U$25610 ( \33760 , RIde1d908_5742);
or \U$25611 ( \33761 , \33760 , \32889 );
buf \U$25612 ( \33762 , RIb886a80_15);
buf \U$25613 ( \33763 , \33762 );
and \U$25614 ( \33764 , \32781 , \33763 );
buf \U$25615 ( \33765 , RIb8389c0_183);
buf \U$25616 ( \33766 , \33765 );
not \U$25617 ( \33767 , \32685 );
and \U$25618 ( \33768 , \33766 , \33767 );
nor \U$25619 ( \33769 , \33764 , \33768 );
nand \U$25620 ( \33770 , \33761 , \33769 );
and \U$25621 ( \33771 , \33770 , \33297 );
or \U$25622 ( \33772 , \33759 , \33771 );
and \U$25624 ( \33773 , \33772 , 1'b1 );
or \U$25626 ( \33774 , \33773 , 1'b0 );
buf \U$25627 ( \33775 , \33774 );
_DC r23a6e_GF_IsGateDCbyConstraint ( \33776_nR23a6e , \33775 , \21944 );
buf \U$25628 ( \33777 , \33776_nR23a6e );
not \U$25629 ( \33778 , \33297 );
and \U$25630 ( \33779 , RIde4a200_5743, \33778 );
not \U$25631 ( \33780 , RIde4a200_5743);
or \U$25632 ( \33781 , \33780 , \32688 );
buf \U$25633 ( \33782 , RIb886af8_14);
buf \U$25634 ( \33783 , \33782 );
and \U$25635 ( \33784 , \32690 , \33783 );
buf \U$25636 ( \33785 , RIb838a38_182);
buf \U$25637 ( \33786 , \33785 );
not \U$25638 ( \33787 , \32723 );
and \U$25639 ( \33788 , \33786 , \33787 );
nor \U$25640 ( \33789 , \33784 , \33788 );
nand \U$25641 ( \33790 , \33781 , \33789 );
and \U$25642 ( \33791 , \33790 , \33297 );
or \U$25643 ( \33792 , \33779 , \33791 );
and \U$25645 ( \33793 , \33792 , 1'b1 );
or \U$25647 ( \33794 , \33793 , 1'b0 );
buf \U$25648 ( \33795 , \33794 );
_DC r23a70_GF_IsGateDCbyConstraint ( \33796_nR23a70 , \33795 , \21944 );
buf \U$25649 ( \33797 , \33796_nR23a70 );
not \U$25650 ( \33798 , \33569 );
and \U$25651 ( \33799 , RIde62e18_5744, \33798 );
not \U$25652 ( \33800 , RIde62e18_5744);
or \U$25653 ( \33801 , \33800 , \32910 );
buf \U$25654 ( \33802 , \23283 );
and \U$25655 ( \33803 , \32739 , \33802 );
buf \U$25656 ( \33804 , RIb838ab0_181);
buf \U$25657 ( \33805 , \33804 );
not \U$25658 ( \33806 , \33053 );
and \U$25659 ( \33807 , \33805 , \33806 );
nor \U$25660 ( \33808 , \33803 , \33807 );
nand \U$25661 ( \33809 , \33801 , \33808 );
and \U$25662 ( \33810 , \33809 , \33569 );
or \U$25663 ( \33811 , \33799 , \33810 );
and \U$25665 ( \33812 , \33811 , 1'b1 );
or \U$25667 ( \33813 , \33812 , 1'b0 );
buf \U$25668 ( \33814 , \33813 );
_DC r23a72_GF_IsGateDCbyConstraint ( \33815_nR23a72 , \33814 , \21944 );
buf \U$25669 ( \33816 , \33815_nR23a72 );
not \U$25670 ( \33817 , \33257 );
and \U$25671 ( \33818 , RIdc30d68_5745, \33817 );
not \U$25672 ( \33819 , RIdc30d68_5745);
or \U$25673 ( \33820 , \33819 , \32779 );
buf \U$25674 ( \33821 , RIb886be8_12);
and \U$25675 ( \33822 , \32781 , \33821 );
buf \U$25676 ( \33823 , RIb838b28_180);
buf \U$25677 ( \33824 , \33823 );
not \U$25678 ( \33825 , \33053 );
and \U$25679 ( \33826 , \33824 , \33825 );
nor \U$25680 ( \33827 , \33822 , \33826 );
nand \U$25681 ( \33828 , \33820 , \33827 );
and \U$25682 ( \33829 , \33828 , \33257 );
or \U$25683 ( \33830 , \33818 , \33829 );
and \U$25685 ( \33831 , \33830 , 1'b1 );
or \U$25687 ( \33832 , \33831 , 1'b0 );
buf \U$25688 ( \33833 , \33832 );
_DC r23a74_GF_IsGateDCbyConstraint ( \33834_nR23a74 , \33833 , \21944 );
buf \U$25689 ( \33835 , \33834_nR23a74 );
not \U$25690 ( \33836 , \33297 );
and \U$25691 ( \33837 , RIdde3e10_5746, \33836 );
not \U$25692 ( \33838 , RIdde3e10_5746);
or \U$25693 ( \33839 , \33838 , \32949 );
buf \U$25694 ( \33840 , \23322 );
and \U$25695 ( \33841 , \32690 , \33840 );
buf \U$25696 ( \33842 , RIb838ba0_179);
buf \U$25697 ( \33843 , \33842 );
not \U$25698 ( \33844 , \32811 );
and \U$25699 ( \33845 , \33843 , \33844 );
nor \U$25700 ( \33846 , \33841 , \33845 );
nand \U$25701 ( \33847 , \33839 , \33846 );
and \U$25702 ( \33848 , \33847 , \33297 );
or \U$25703 ( \33849 , \33837 , \33848 );
and \U$25705 ( \33850 , \33849 , 1'b1 );
or \U$25707 ( \33851 , \33850 , 1'b0 );
buf \U$25708 ( \33852 , \33851 );
_DC r23a76_GF_IsGateDCbyConstraint ( \33853_nR23a76 , \33852 , \21944 );
buf \U$25709 ( \33854 , \33853_nR23a76 );
not \U$25710 ( \33855 , \33569 );
and \U$25711 ( \33856 , RIddce948_5747, \33855 );
not \U$25712 ( \33857 , RIddce948_5747);
or \U$25713 ( \33858 , \33857 , \32968 );
buf \U$25714 ( \33859 , \28547 );
and \U$25715 ( \33860 , \32739 , \33859 );
buf \U$25716 ( \33861 , RIb838c18_178);
buf \U$25717 ( \33862 , \33861 );
not \U$25718 ( \33863 , \32974 );
and \U$25719 ( \33864 , \33862 , \33863 );
nor \U$25720 ( \33865 , \33860 , \33864 );
nand \U$25721 ( \33866 , \33858 , \33865 );
and \U$25722 ( \33867 , \33866 , \33569 );
or \U$25723 ( \33868 , \33856 , \33867 );
and \U$25725 ( \33869 , \33868 , 1'b1 );
or \U$25727 ( \33870 , \33869 , 1'b0 );
buf \U$25728 ( \33871 , \33870 );
_DC r23a78_GF_IsGateDCbyConstraint ( \33872_nR23a78 , \33871 , \21944 );
buf \U$25729 ( \33873 , \33872_nR23a78 );
buf \U$25730 ( \33874 , \33296 );
not \U$25731 ( \33875 , \33874 );
and \U$25732 ( \33876 , RIdb96b50_5748, \33875 );
not \U$25733 ( \33877 , RIdb96b50_5748);
or \U$25734 ( \33878 , \33877 , \32688 );
buf \U$25735 ( \33879 , \28568 );
and \U$25736 ( \33880 , \32690 , \33879 );
buf \U$25737 ( \33881 , RIb838c90_177);
buf \U$25738 ( \33882 , \33881 );
not \U$25739 ( \33883 , \32852 );
and \U$25740 ( \33884 , \33882 , \33883 );
nor \U$25741 ( \33885 , \33880 , \33884 );
nand \U$25742 ( \33886 , \33878 , \33885 );
and \U$25743 ( \33887 , \33886 , \33874 );
or \U$25744 ( \33888 , \33876 , \33887 );
and \U$25746 ( \33889 , \33888 , 1'b1 );
or \U$25748 ( \33890 , \33889 , 1'b0 );
buf \U$25749 ( \33891 , \33890 );
_DC r23a7c_GF_IsGateDCbyConstraint ( \33892_nR23a7c , \33891 , \21944 );
buf \U$25750 ( \33893 , \33892_nR23a7c );
not \U$25751 ( \33894 , \33874 );
and \U$25752 ( \33895 , RIda0b300_5749, \33894 );
not \U$25753 ( \33896 , RIda0b300_5749);
or \U$25754 ( \33897 , \33896 , \32910 );
buf \U$25755 ( \33898 , RIb886dc8_8);
buf \U$25756 ( \33899 , \33898 );
and \U$25757 ( \33900 , \32781 , \33899 );
buf \U$25758 ( \33901 , RIb838d08_176);
buf \U$25759 ( \33902 , \33901 );
not \U$25760 ( \33903 , \32874 );
and \U$25761 ( \33904 , \33902 , \33903 );
nor \U$25762 ( \33905 , \33900 , \33904 );
nand \U$25763 ( \33906 , \33897 , \33905 );
and \U$25764 ( \33907 , \33906 , \33874 );
or \U$25765 ( \33908 , \33895 , \33907 );
and \U$25767 ( \33909 , \33908 , 1'b1 );
or \U$25769 ( \33910 , \33909 , 1'b0 );
buf \U$25770 ( \33911 , \33910 );
_DC r23a7e_GF_IsGateDCbyConstraint ( \33912_nR23a7e , \33911 , \21944 );
buf \U$25771 ( \33913 , \33912_nR23a7e );
not \U$25772 ( \33914 , \33569 );
and \U$25773 ( \33915 , RIdc00960_5750, \33914 );
not \U$25774 ( \33916 , RIdc00960_5750);
or \U$25775 ( \33917 , \33916 , \32779 );
buf \U$25776 ( \33918 , \23403 );
and \U$25777 ( \33919 , \32781 , \33918 );
buf \U$25778 ( \33920 , RIb838d80_175);
buf \U$25779 ( \33921 , \33920 );
not \U$25780 ( \33922 , \32974 );
and \U$25781 ( \33923 , \33921 , \33922 );
nor \U$25782 ( \33924 , \33919 , \33923 );
nand \U$25783 ( \33925 , \33917 , \33924 );
and \U$25784 ( \33926 , \33925 , \33569 );
or \U$25785 ( \33927 , \33915 , \33926 );
and \U$25787 ( \33928 , \33927 , 1'b1 );
or \U$25789 ( \33929 , \33928 , 1'b0 );
buf \U$25790 ( \33930 , \33929 );
_DC r23a80_GF_IsGateDCbyConstraint ( \33931_nR23a80 , \33930 , \21944 );
buf \U$25791 ( \33932 , \33931_nR23a80 );
not \U$25792 ( \33933 , \33257 );
and \U$25793 ( \33934 , RIdb708e8_5751, \33933 );
not \U$25794 ( \33935 , RIdb708e8_5751);
or \U$25795 ( \33936 , \33935 , \32949 );
buf \U$25796 ( \33937 , \23423 );
and \U$25797 ( \33938 , \32690 , \33937 );
buf \U$25798 ( \33939 , RIb838df8_174);
buf \U$25799 ( \33940 , \33939 );
not \U$25800 ( \33941 , \32895 );
and \U$25801 ( \33942 , \33940 , \33941 );
nor \U$25802 ( \33943 , \33938 , \33942 );
nand \U$25803 ( \33944 , \33936 , \33943 );
and \U$25804 ( \33945 , \33944 , \33257 );
or \U$25805 ( \33946 , \33934 , \33945 );
and \U$25807 ( \33947 , \33946 , 1'b1 );
or \U$25809 ( \33948 , \33947 , 1'b0 );
buf \U$25810 ( \33949 , \33948 );
_DC r23a82_GF_IsGateDCbyConstraint ( \33950_nR23a82 , \33949 , \21944 );
buf \U$25811 ( \33951 , \33950_nR23a82 );
not \U$25812 ( \33952 , \33257 );
and \U$25813 ( \33953 , RIdc692d0_5752, \33952 );
not \U$25814 ( \33954 , RIdc692d0_5752);
not \U$25815 ( \33955 , \32680 );
nor \U$25816 ( \33956 , \32678 , \33955 );
nand \U$25817 ( \33957 , \33956 , \32682 );
not \U$25818 ( \33958 , \33957 );
not \U$25819 ( \33959 , \32670 );
or \U$25820 ( \33960 , \32672 , \33959 );
not \U$25821 ( \33961 , \33960 );
nand \U$25822 ( \33962 , \32664 , \33961 );
not \U$25823 ( \33963 , \33962 );
or \U$25824 ( \33964 , \33958 , \33963 );
not \U$25825 ( \33965 , \33964 );
not \U$25826 ( \33966 , \33965 );
or \U$25827 ( \33967 , \33954 , \33966 );
not \U$25828 ( \33968 , \33957 );
not \U$25829 ( \33969 , \33968 );
not \U$25830 ( \33970 , \33969 );
and \U$25831 ( \33971 , \32694 , \33970 );
not \U$25832 ( \33972 , \33971 );
not \U$25833 ( \33973 , \32691 );
not \U$25834 ( \33974 , \33962 );
buf \U$25835 ( \33975 , \33974 );
not \U$25836 ( \33976 , \33975 );
or \U$25837 ( \33977 , \33973 , \33976 );
nand \U$25838 ( \33978 , \33967 , \33972 , \33977 );
and \U$25839 ( \33979 , \33978 , \33257 );
or \U$25840 ( \33980 , \33953 , \33979 );
and \U$25842 ( \33981 , \33980 , 1'b1 );
or \U$25844 ( \33982 , \33981 , 1'b0 );
buf \U$25845 ( \33983 , \33982 );
_DC r23a8c_GF_IsGateDCbyConstraint ( \33984_nR23a8c , \33983 , \21944 );
buf \U$25846 ( \33985 , \33984_nR23a8c );
not \U$25847 ( \33986 , \33569 );
and \U$25848 ( \33987 , RIdf7e930_5753, \33986 );
not \U$25849 ( \33988 , RIdf7e930_5753);
not \U$25850 ( \33989 , \33965 );
or \U$25851 ( \33990 , \33988 , \33989 );
not \U$25852 ( \33991 , \33968 );
not \U$25853 ( \33992 , \33991 );
and \U$25854 ( \33993 , \32722 , \33992 );
not \U$25855 ( \33994 , \33993 );
not \U$25856 ( \33995 , \32719 );
not \U$25857 ( \33996 , \33975 );
or \U$25858 ( \33997 , \33995 , \33996 );
nand \U$25859 ( \33998 , \33990 , \33994 , \33997 );
and \U$25860 ( \33999 , \33998 , \33569 );
or \U$25861 ( \34000 , \33987 , \33999 );
and \U$25863 ( \34001 , \34000 , 1'b1 );
or \U$25865 ( \34002 , \34001 , 1'b0 );
buf \U$25866 ( \34003 , \34002 );
_DC r23aa2_GF_IsGateDCbyConstraint ( \34004_nR23aa2 , \34003 , \21944 );
buf \U$25867 ( \34005 , \34004_nR23aa2 );
not \U$25868 ( \34006 , \33257 );
and \U$25869 ( \34007 , RIdf8d6d8_5754, \34006 );
not \U$25870 ( \34008 , RIdf8d6d8_5754);
or \U$25871 ( \34009 , \34008 , \33989 );
not \U$25872 ( \34010 , \33969 );
and \U$25873 ( \34011 , \32743 , \34010 );
not \U$25874 ( \34012 , \34011 );
not \U$25875 ( \34013 , \32740 );
not \U$25876 ( \34014 , \33975 );
or \U$25877 ( \34015 , \34013 , \34014 );
nand \U$25878 ( \34016 , \34009 , \34012 , \34015 );
and \U$25879 ( \34017 , \34016 , \33257 );
or \U$25880 ( \34018 , \34007 , \34017 );
and \U$25882 ( \34019 , \34018 , 1'b1 );
or \U$25884 ( \34020 , \34019 , 1'b0 );
buf \U$25885 ( \34021 , \34020 );
_DC r23ab8_GF_IsGateDCbyConstraint ( \34022_nR23ab8 , \34021 , \21944 );
buf \U$25886 ( \34023 , \34022_nR23ab8 );
not \U$25887 ( \34024 , \33874 );
and \U$25888 ( \34025 , RIdf9f978_5755, \34024 );
not \U$25889 ( \34026 , RIdf9f978_5755);
or \U$25890 ( \34027 , \34026 , \33989 );
not \U$25891 ( \34028 , \33968 );
not \U$25892 ( \34029 , \34028 );
and \U$25893 ( \34030 , \32764 , \34029 );
not \U$25894 ( \34031 , \34030 );
not \U$25895 ( \34032 , \32761 );
buf \U$25896 ( \34033 , \33974 );
not \U$25897 ( \34034 , \34033 );
or \U$25898 ( \34035 , \34032 , \34034 );
nand \U$25899 ( \34036 , \34027 , \34031 , \34035 );
and \U$25900 ( \34037 , \34036 , \33874 );
or \U$25901 ( \34038 , \34025 , \34037 );
and \U$25903 ( \34039 , \34038 , 1'b1 );
or \U$25905 ( \34040 , \34039 , 1'b0 );
buf \U$25906 ( \34041 , \34040 );
_DC r23ace_GF_IsGateDCbyConstraint ( \34042_nR23ace , \34041 , \21944 );
buf \U$25907 ( \34043 , \34042_nR23ace );
not \U$25908 ( \34044 , \33569 );
and \U$25909 ( \34045 , RIdfa6f20_5756, \34044 );
not \U$25910 ( \34046 , RIdfa6f20_5756);
not \U$25911 ( \34047 , \33965 );
or \U$25912 ( \34048 , \34046 , \34047 );
not \U$25913 ( \34049 , \33969 );
and \U$25914 ( \34050 , \32786 , \34049 );
not \U$25915 ( \34051 , \34050 );
not \U$25916 ( \34052 , \32783 );
not \U$25917 ( \34053 , \34033 );
or \U$25918 ( \34054 , \34052 , \34053 );
nand \U$25919 ( \34055 , \34048 , \34051 , \34054 );
and \U$25920 ( \34056 , \34055 , \33569 );
or \U$25921 ( \34057 , \34045 , \34056 );
and \U$25923 ( \34058 , \34057 , 1'b1 );
or \U$25925 ( \34059 , \34058 , 1'b0 );
buf \U$25926 ( \34060 , \34059 );
_DC r23ae4_GF_IsGateDCbyConstraint ( \34061_nR23ae4 , \34060 , \21944 );
buf \U$25927 ( \34062 , \34061_nR23ae4 );
not \U$25928 ( \34063 , \33336 );
and \U$25929 ( \34064 , RIdfaf968_5757, \34063 );
not \U$25930 ( \34065 , RIdfaf968_5757);
or \U$25931 ( \34066 , \34065 , \33964 );
not \U$25932 ( \34067 , \34028 );
and \U$25933 ( \34068 , \32806 , \34067 );
not \U$25934 ( \34069 , \34068 );
not \U$25935 ( \34070 , \32804 );
buf \U$25936 ( \34071 , \33974 );
not \U$25937 ( \34072 , \34071 );
or \U$25938 ( \34073 , \34070 , \34072 );
nand \U$25939 ( \34074 , \34066 , \34069 , \34073 );
and \U$25940 ( \34075 , \34074 , \33336 );
or \U$25941 ( \34076 , \34064 , \34075 );
and \U$25943 ( \34077 , \34076 , 1'b1 );
or \U$25945 ( \34078 , \34077 , 1'b0 );
buf \U$25946 ( \34079 , \34078 );
_DC r23afa_GF_IsGateDCbyConstraint ( \34080_nR23afa , \34079 , \21944 );
buf \U$25947 ( \34081 , \34080_nR23afa );
not \U$25948 ( \34082 , \33336 );
and \U$25949 ( \34083 , RIdfb74b0_5758, \34082 );
not \U$25950 ( \34084 , RIdfb74b0_5758);
or \U$25951 ( \34085 , \34084 , \33989 );
not \U$25952 ( \34086 , \33968 );
not \U$25953 ( \34087 , \34086 );
and \U$25954 ( \34088 , \32829 , \34087 );
not \U$25955 ( \34089 , \34088 );
not \U$25956 ( \34090 , \32827 );
not \U$25957 ( \34091 , \34033 );
or \U$25958 ( \34092 , \34090 , \34091 );
nand \U$25959 ( \34093 , \34085 , \34089 , \34092 );
and \U$25960 ( \34094 , \34093 , \33336 );
or \U$25961 ( \34095 , \34083 , \34094 );
and \U$25963 ( \34096 , \34095 , 1'b1 );
or \U$25965 ( \34097 , \34096 , 1'b0 );
buf \U$25966 ( \34098 , \34097 );
_DC r23b04_GF_IsGateDCbyConstraint ( \34099_nR23b04 , \34098 , \21944 );
buf \U$25967 ( \34100 , \34099_nR23b04 );
not \U$25968 ( \34101 , \33569 );
and \U$25969 ( \34102 , RIddf5a98_5759, \34101 );
not \U$25970 ( \34103 , RIddf5a98_5759);
or \U$25971 ( \34104 , \34103 , \33989 );
not \U$25972 ( \34105 , \34086 );
and \U$25973 ( \34106 , \32851 , \34105 );
not \U$25974 ( \34107 , \34106 );
not \U$25975 ( \34108 , \32848 );
not \U$25976 ( \34109 , \34071 );
or \U$25977 ( \34110 , \34108 , \34109 );
nand \U$25978 ( \34111 , \34104 , \34107 , \34110 );
and \U$25979 ( \34112 , \34111 , \33569 );
or \U$25980 ( \34113 , \34102 , \34112 );
and \U$25982 ( \34114 , \34113 , 1'b1 );
or \U$25984 ( \34115 , \34114 , 1'b0 );
buf \U$25985 ( \34116 , \34115 );
_DC r23b06_GF_IsGateDCbyConstraint ( \34117_nR23b06 , \34116 , \21944 );
buf \U$25986 ( \34118 , \34117_nR23b06 );
not \U$25987 ( \34119 , \33874 );
and \U$25988 ( \34120 , RIde028d8_5760, \34119 );
not \U$25989 ( \34121 , RIde028d8_5760);
or \U$25990 ( \34122 , \34121 , \33989 );
not \U$25991 ( \34123 , \33991 );
and \U$25992 ( \34124 , \32873 , \34123 );
not \U$25993 ( \34125 , \34124 );
not \U$25994 ( \34126 , \32870 );
not \U$25995 ( \34127 , \34033 );
or \U$25996 ( \34128 , \34126 , \34127 );
nand \U$25997 ( \34129 , \34122 , \34125 , \34128 );
and \U$25998 ( \34130 , \34129 , \33874 );
or \U$25999 ( \34131 , \34120 , \34130 );
and \U$26001 ( \34132 , \34131 , 1'b1 );
or \U$26003 ( \34133 , \34132 , 1'b0 );
buf \U$26004 ( \34134 , \34133 );
_DC r23b08_GF_IsGateDCbyConstraint ( \34135_nR23b08 , \34134 , \21944 );
buf \U$26005 ( \34136 , \34135_nR23b08 );
not \U$26006 ( \34137 , \33874 );
and \U$26007 ( \34138 , RIe036620_5761, \34137 );
not \U$26008 ( \34139 , RIe036620_5761);
or \U$26009 ( \34140 , \34139 , \33966 );
not \U$26010 ( \34141 , \33969 );
and \U$26011 ( \34142 , \32894 , \34141 );
not \U$26012 ( \34143 , \34142 );
not \U$26013 ( \34144 , \32891 );
not \U$26014 ( \34145 , \34033 );
or \U$26015 ( \34146 , \34144 , \34145 );
nand \U$26016 ( \34147 , \34140 , \34143 , \34146 );
and \U$26017 ( \34148 , \34147 , \33874 );
or \U$26018 ( \34149 , \34138 , \34148 );
and \U$26020 ( \34150 , \34149 , 1'b1 );
or \U$26022 ( \34151 , \34150 , 1'b0 );
buf \U$26023 ( \34152 , \34151 );
_DC r23b0a_GF_IsGateDCbyConstraint ( \34153_nR23b0a , \34152 , \21944 );
buf \U$26024 ( \34154 , \34153_nR23b0a );
not \U$26025 ( \34155 , \33569 );
and \U$26026 ( \34156 , RIe027530_5762, \34155 );
not \U$26027 ( \34157 , RIe027530_5762);
or \U$26028 ( \34158 , \34157 , \34047 );
not \U$26029 ( \34159 , \33991 );
and \U$26030 ( \34160 , \32914 , \34159 );
not \U$26031 ( \34161 , \34160 );
not \U$26032 ( \34162 , \32912 );
not \U$26033 ( \34163 , \34071 );
or \U$26034 ( \34164 , \34162 , \34163 );
nand \U$26035 ( \34165 , \34158 , \34161 , \34164 );
and \U$26036 ( \34166 , \34165 , \33569 );
or \U$26037 ( \34167 , \34156 , \34166 );
and \U$26039 ( \34168 , \34167 , 1'b1 );
or \U$26041 ( \34169 , \34168 , 1'b0 );
buf \U$26042 ( \34170 , \34169 );
_DC r23a8e_GF_IsGateDCbyConstraint ( \34171_nR23a8e , \34170 , \21944 );
buf \U$26043 ( \34172 , \34171_nR23a8e );
not \U$26044 ( \34173 , \33336 );
and \U$26045 ( \34174 , RIe01deb8_5763, \34173 );
not \U$26046 ( \34175 , RIe01deb8_5763);
or \U$26047 ( \34176 , \34175 , \33964 );
not \U$26048 ( \34177 , \34028 );
and \U$26049 ( \34178 , \32934 , \34177 );
not \U$26050 ( \34179 , \34178 );
not \U$26051 ( \34180 , \32931 );
not \U$26052 ( \34181 , \33975 );
or \U$26053 ( \34182 , \34180 , \34181 );
nand \U$26054 ( \34183 , \34176 , \34179 , \34182 );
and \U$26055 ( \34184 , \34183 , \33336 );
or \U$26056 ( \34185 , \34174 , \34184 );
and \U$26058 ( \34186 , \34185 , 1'b1 );
or \U$26060 ( \34187 , \34186 , 1'b0 );
buf \U$26061 ( \34188 , \34187 );
_DC r23a90_GF_IsGateDCbyConstraint ( \34189_nR23a90 , \34188 , \21944 );
buf \U$26062 ( \34190 , \34189_nR23a90 );
not \U$26063 ( \34191 , \33336 );
and \U$26064 ( \34192 , RIe00b3a8_5764, \34191 );
not \U$26065 ( \34193 , RIe00b3a8_5764);
or \U$26066 ( \34194 , \34193 , \33989 );
not \U$26067 ( \34195 , \34086 );
and \U$26068 ( \34196 , \32953 , \34195 );
not \U$26069 ( \34197 , \34196 );
not \U$26070 ( \34198 , \32951 );
not \U$26071 ( \34199 , \33975 );
or \U$26072 ( \34200 , \34198 , \34199 );
nand \U$26073 ( \34201 , \34194 , \34197 , \34200 );
and \U$26074 ( \34202 , \34201 , \33336 );
or \U$26075 ( \34203 , \34192 , \34202 );
and \U$26077 ( \34204 , \34203 , 1'b1 );
or \U$26079 ( \34205 , \34204 , 1'b0 );
buf \U$26080 ( \34206 , \34205 );
_DC r23a92_GF_IsGateDCbyConstraint ( \34207_nR23a92 , \34206 , \21944 );
buf \U$26081 ( \34208 , \34207_nR23a92 );
not \U$26082 ( \34209 , \33569 );
and \U$26083 ( \34210 , RIdffd938_5765, \34209 );
not \U$26084 ( \34211 , RIdffd938_5765);
or \U$26085 ( \34212 , \34211 , \33966 );
not \U$26086 ( \34213 , \33969 );
and \U$26087 ( \34214 , \32973 , \34213 );
not \U$26088 ( \34215 , \34214 );
not \U$26089 ( \34216 , \32970 );
not \U$26090 ( \34217 , \33975 );
or \U$26091 ( \34218 , \34216 , \34217 );
nand \U$26092 ( \34219 , \34212 , \34215 , \34218 );
and \U$26093 ( \34220 , \34219 , \33569 );
or \U$26094 ( \34221 , \34210 , \34220 );
and \U$26096 ( \34222 , \34221 , 1'b1 );
or \U$26098 ( \34223 , \34222 , 1'b0 );
buf \U$26099 ( \34224 , \34223 );
_DC r23a94_GF_IsGateDCbyConstraint ( \34225_nR23a94 , \34224 , \21944 );
buf \U$26100 ( \34226 , \34225_nR23a94 );
not \U$26101 ( \34227 , \33336 );
and \U$26102 ( \34228 , RIdfefb08_5766, \34227 );
not \U$26103 ( \34229 , RIdfefb08_5766);
or \U$26104 ( \34230 , \34229 , \33966 );
not \U$26105 ( \34231 , \33991 );
and \U$26106 ( \34232 , \32994 , \34231 );
not \U$26107 ( \34233 , \34232 );
not \U$26108 ( \34234 , \32991 );
not \U$26109 ( \34235 , \34071 );
or \U$26110 ( \34236 , \34234 , \34235 );
nand \U$26111 ( \34237 , \34230 , \34233 , \34236 );
and \U$26112 ( \34238 , \34237 , \33336 );
or \U$26113 ( \34239 , \34228 , \34238 );
and \U$26115 ( \34240 , \34239 , 1'b1 );
or \U$26117 ( \34241 , \34240 , 1'b0 );
buf \U$26118 ( \34242 , \34241 );
_DC r23a96_GF_IsGateDCbyConstraint ( \34243_nR23a96 , \34242 , \21944 );
buf \U$26119 ( \34244 , \34243_nR23a96 );
not \U$26120 ( \34245 , \33874 );
and \U$26121 ( \34246 , RIdfe0838_5767, \34245 );
not \U$26122 ( \34247 , RIdfe0838_5767);
or \U$26123 ( \34248 , \34247 , \33966 );
not \U$26124 ( \34249 , \34028 );
and \U$26125 ( \34250 , \33014 , \34249 );
not \U$26126 ( \34251 , \34250 );
not \U$26127 ( \34252 , \33011 );
not \U$26128 ( \34253 , \33974 );
or \U$26129 ( \34254 , \34252 , \34253 );
nand \U$26130 ( \34255 , \34248 , \34251 , \34254 );
and \U$26131 ( \34256 , \34255 , \33874 );
or \U$26132 ( \34257 , \34246 , \34256 );
and \U$26134 ( \34258 , \34257 , 1'b1 );
or \U$26136 ( \34259 , \34258 , 1'b0 );
buf \U$26137 ( \34260 , \34259 );
_DC r23a98_GF_IsGateDCbyConstraint ( \34261_nR23a98 , \34260 , \21944 );
buf \U$26138 ( \34262 , \34261_nR23a98 );
not \U$26139 ( \34263 , \33296 );
and \U$26140 ( \34264 , RIdfd6680_5768, \34263 );
not \U$26141 ( \34265 , RIdfd6680_5768);
or \U$26142 ( \34266 , \34265 , \33989 );
not \U$26143 ( \34267 , \34086 );
and \U$26144 ( \34268 , \33033 , \34267 );
not \U$26145 ( \34269 , \34268 );
not \U$26146 ( \34270 , \33030 );
not \U$26147 ( \34271 , \34071 );
or \U$26148 ( \34272 , \34270 , \34271 );
nand \U$26149 ( \34273 , \34266 , \34269 , \34272 );
and \U$26150 ( \34274 , \34273 , \33296 );
or \U$26151 ( \34275 , \34264 , \34274 );
and \U$26153 ( \34276 , \34275 , 1'b1 );
or \U$26155 ( \34277 , \34276 , 1'b0 );
buf \U$26156 ( \34278 , \34277 );
_DC r23a9a_GF_IsGateDCbyConstraint ( \34279_nR23a9a , \34278 , \21944 );
buf \U$26157 ( \34280 , \34279_nR23a9a );
not \U$26158 ( \34281 , \33336 );
and \U$26159 ( \34282 , RIe1084d0_5769, \34281 );
not \U$26160 ( \34283 , RIe1084d0_5769);
or \U$26161 ( \34284 , \34283 , \33989 );
not \U$26162 ( \34285 , \34086 );
and \U$26163 ( \34286 , \33052 , \34285 );
not \U$26164 ( \34287 , \34286 );
not \U$26165 ( \34288 , \33050 );
not \U$26166 ( \34289 , \33974 );
or \U$26167 ( \34290 , \34288 , \34289 );
nand \U$26168 ( \34291 , \34284 , \34287 , \34290 );
and \U$26169 ( \34292 , \34291 , \33336 );
or \U$26170 ( \34293 , \34282 , \34292 );
and \U$26172 ( \34294 , \34293 , 1'b1 );
or \U$26174 ( \34295 , \34294 , 1'b0 );
buf \U$26175 ( \34296 , \34295 );
_DC r23a9c_GF_IsGateDCbyConstraint ( \34297_nR23a9c , \34296 , \21944 );
buf \U$26176 ( \34298 , \34297_nR23a9c );
not \U$26177 ( \34299 , \33874 );
and \U$26178 ( \34300 , RIe10ad98_5770, \34299 );
not \U$26179 ( \34301 , RIe10ad98_5770);
or \U$26180 ( \34302 , \34301 , \33966 );
not \U$26181 ( \34303 , \33958 );
not \U$26182 ( \34304 , \34303 );
and \U$26183 ( \34305 , \33071 , \34304 );
not \U$26184 ( \34306 , \34305 );
not \U$26185 ( \34307 , \33069 );
not \U$26186 ( \34308 , \34033 );
or \U$26187 ( \34309 , \34307 , \34308 );
nand \U$26188 ( \34310 , \34302 , \34306 , \34309 );
and \U$26189 ( \34311 , \34310 , \33874 );
or \U$26190 ( \34312 , \34300 , \34311 );
and \U$26192 ( \34313 , \34312 , 1'b1 );
or \U$26194 ( \34314 , \34313 , 1'b0 );
buf \U$26195 ( \34315 , \34314 );
_DC r23a9e_GF_IsGateDCbyConstraint ( \34316_nR23a9e , \34315 , \21944 );
buf \U$26196 ( \34317 , \34316_nR23a9e );
buf \U$26197 ( \34318 , \32665 );
not \U$26198 ( \34319 , \34318 );
and \U$26199 ( \34320 , RIe10e470_5771, \34319 );
not \U$26200 ( \34321 , RIe10e470_5771);
or \U$26201 ( \34322 , \34321 , \33964 );
not \U$26202 ( \34323 , \33969 );
and \U$26203 ( \34324 , \33091 , \34323 );
not \U$26204 ( \34325 , \34324 );
not \U$26205 ( \34326 , \33088 );
not \U$26206 ( \34327 , \33975 );
or \U$26207 ( \34328 , \34326 , \34327 );
nand \U$26208 ( \34329 , \34322 , \34325 , \34328 );
and \U$26209 ( \34330 , \34329 , \34318 );
or \U$26210 ( \34331 , \34320 , \34330 );
and \U$26212 ( \34332 , \34331 , 1'b1 );
or \U$26214 ( \34333 , \34332 , 1'b0 );
buf \U$26215 ( \34334 , \34333 );
_DC r23aa0_GF_IsGateDCbyConstraint ( \34335_nR23aa0 , \34334 , \21944 );
buf \U$26216 ( \34336 , \34335_nR23aa0 );
not \U$26217 ( \34337 , \33874 );
and \U$26218 ( \34338 , RIe110d38_5772, \34337 );
not \U$26219 ( \34339 , RIe110d38_5772);
or \U$26220 ( \34340 , \34339 , \33966 );
not \U$26221 ( \34341 , \33969 );
and \U$26222 ( \34342 , \33110 , \34341 );
not \U$26223 ( \34343 , \34342 );
not \U$26224 ( \34344 , \33107 );
not \U$26225 ( \34345 , \33974 );
or \U$26226 ( \34346 , \34344 , \34345 );
nand \U$26227 ( \34347 , \34340 , \34343 , \34346 );
and \U$26228 ( \34348 , \34347 , \33874 );
or \U$26229 ( \34349 , \34338 , \34348 );
and \U$26231 ( \34350 , \34349 , 1'b1 );
or \U$26233 ( \34351 , \34350 , 1'b0 );
buf \U$26234 ( \34352 , \34351 );
_DC r23aa4_GF_IsGateDCbyConstraint ( \34353_nR23aa4 , \34352 , \21944 );
buf \U$26235 ( \34354 , \34353_nR23aa4 );
not \U$26236 ( \34355 , \33874 );
and \U$26237 ( \34356 , RIe113ab0_5773, \34355 );
not \U$26238 ( \34357 , RIe113ab0_5773);
or \U$26239 ( \34358 , \34357 , \33964 );
not \U$26240 ( \34359 , \33969 );
and \U$26241 ( \34360 , \33129 , \34359 );
not \U$26242 ( \34361 , \34360 );
not \U$26243 ( \34362 , \33126 );
not \U$26244 ( \34363 , \33974 );
or \U$26245 ( \34364 , \34362 , \34363 );
nand \U$26246 ( \34365 , \34358 , \34361 , \34364 );
and \U$26247 ( \34366 , \34365 , \33874 );
or \U$26248 ( \34367 , \34356 , \34366 );
and \U$26250 ( \34368 , \34367 , 1'b1 );
or \U$26252 ( \34369 , \34368 , 1'b0 );
buf \U$26253 ( \34370 , \34369 );
_DC r23aa6_GF_IsGateDCbyConstraint ( \34371_nR23aa6 , \34370 , \21944 );
buf \U$26254 ( \34372 , \34371_nR23aa6 );
not \U$26255 ( \34373 , \32755 );
and \U$26256 ( \34374 , RIe116cd8_5774, \34373 );
not \U$26257 ( \34375 , RIe116cd8_5774);
or \U$26258 ( \34376 , \34375 , \34047 );
not \U$26259 ( \34377 , \33969 );
and \U$26260 ( \34378 , \33149 , \34377 );
not \U$26261 ( \34379 , \34378 );
not \U$26262 ( \34380 , \33146 );
not \U$26263 ( \34381 , \33975 );
or \U$26264 ( \34382 , \34380 , \34381 );
nand \U$26265 ( \34383 , \34376 , \34379 , \34382 );
and \U$26266 ( \34384 , \34383 , \32755 );
or \U$26267 ( \34385 , \34374 , \34384 );
and \U$26269 ( \34386 , \34385 , 1'b1 );
or \U$26271 ( \34387 , \34386 , 1'b0 );
buf \U$26272 ( \34388 , \34387 );
_DC r23aa8_GF_IsGateDCbyConstraint ( \34389_nR23aa8 , \34388 , \21944 );
buf \U$26273 ( \34390 , \34389_nR23aa8 );
not \U$26274 ( \34391 , \33336 );
and \U$26275 ( \34392 , RIe119a50_5775, \34391 );
not \U$26276 ( \34393 , RIe119a50_5775);
or \U$26277 ( \34394 , \34393 , \34047 );
not \U$26278 ( \34395 , \33991 );
and \U$26279 ( \34396 , \33167 , \34395 );
not \U$26280 ( \34397 , \34396 );
not \U$26281 ( \34398 , \33165 );
not \U$26282 ( \34399 , \33974 );
or \U$26283 ( \34400 , \34398 , \34399 );
nand \U$26284 ( \34401 , \34394 , \34397 , \34400 );
and \U$26285 ( \34402 , \34401 , \33336 );
or \U$26286 ( \34403 , \34392 , \34402 );
and \U$26288 ( \34404 , \34403 , 1'b1 );
or \U$26290 ( \34405 , \34404 , 1'b0 );
buf \U$26291 ( \34406 , \34405 );
_DC r23aaa_GF_IsGateDCbyConstraint ( \34407_nR23aaa , \34406 , \21944 );
buf \U$26292 ( \34408 , \34407_nR23aaa );
not \U$26293 ( \34409 , \33336 );
and \U$26294 ( \34410 , RIe11cc78_5776, \34409 );
not \U$26295 ( \34411 , RIe11cc78_5776);
or \U$26296 ( \34412 , \34411 , \33989 );
not \U$26297 ( \34413 , \34086 );
and \U$26298 ( \34414 , \33187 , \34413 );
not \U$26299 ( \34415 , \34414 );
not \U$26300 ( \34416 , \33184 );
not \U$26301 ( \34417 , \34071 );
or \U$26302 ( \34418 , \34416 , \34417 );
nand \U$26303 ( \34419 , \34412 , \34415 , \34418 );
and \U$26304 ( \34420 , \34419 , \33336 );
or \U$26305 ( \34421 , \34410 , \34420 );
and \U$26307 ( \34422 , \34421 , 1'b1 );
or \U$26309 ( \34423 , \34422 , 1'b0 );
buf \U$26310 ( \34424 , \34423 );
_DC r23aac_GF_IsGateDCbyConstraint ( \34425_nR23aac , \34424 , \21944 );
buf \U$26311 ( \34426 , \34425_nR23aac );
not \U$26312 ( \34427 , \33217 );
and \U$26313 ( \34428 , RIe11f9f0_5777, \34427 );
not \U$26314 ( \34429 , RIe11f9f0_5777);
or \U$26315 ( \34430 , \34429 , \34047 );
not \U$26316 ( \34431 , \33969 );
and \U$26317 ( \34432 , \33205 , \34431 );
not \U$26318 ( \34433 , \34432 );
not \U$26319 ( \34434 , \33203 );
not \U$26320 ( \34435 , \33975 );
or \U$26321 ( \34436 , \34434 , \34435 );
nand \U$26322 ( \34437 , \34430 , \34433 , \34436 );
and \U$26323 ( \34438 , \34437 , \33217 );
or \U$26324 ( \34439 , \34428 , \34438 );
and \U$26326 ( \34440 , \34439 , 1'b1 );
or \U$26328 ( \34441 , \34440 , 1'b0 );
buf \U$26329 ( \34442 , \34441 );
_DC r23aae_GF_IsGateDCbyConstraint ( \34443_nR23aae , \34442 , \21944 );
buf \U$26330 ( \34444 , \34443_nR23aae );
not \U$26331 ( \34445 , \33336 );
and \U$26332 ( \34446 , RIe122c18_5778, \34445 );
not \U$26333 ( \34447 , RIe122c18_5778);
or \U$26334 ( \34448 , \34447 , \33989 );
not \U$26335 ( \34449 , \34303 );
and \U$26336 ( \34450 , \33226 , \34449 );
not \U$26337 ( \34451 , \34450 );
not \U$26338 ( \34452 , \33223 );
not \U$26339 ( \34453 , \33974 );
or \U$26340 ( \34454 , \34452 , \34453 );
nand \U$26341 ( \34455 , \34448 , \34451 , \34454 );
and \U$26342 ( \34456 , \34455 , \33336 );
or \U$26343 ( \34457 , \34446 , \34456 );
and \U$26345 ( \34458 , \34457 , 1'b1 );
or \U$26347 ( \34459 , \34458 , 1'b0 );
buf \U$26348 ( \34460 , \34459 );
_DC r23ab0_GF_IsGateDCbyConstraint ( \34461_nR23ab0 , \34460 , \21944 );
buf \U$26349 ( \34462 , \34461_nR23ab0 );
not \U$26350 ( \34463 , \33874 );
and \U$26351 ( \34464 , RIe125990_5779, \34463 );
not \U$26352 ( \34465 , RIe125990_5779);
or \U$26353 ( \34466 , \34465 , \33964 );
not \U$26354 ( \34467 , \34303 );
and \U$26355 ( \34468 , \33245 , \34467 );
not \U$26356 ( \34469 , \34468 );
not \U$26357 ( \34470 , \33242 );
not \U$26358 ( \34471 , \34033 );
or \U$26359 ( \34472 , \34470 , \34471 );
nand \U$26360 ( \34473 , \34466 , \34469 , \34472 );
and \U$26361 ( \34474 , \34473 , \33874 );
or \U$26362 ( \34475 , \34464 , \34474 );
and \U$26364 ( \34476 , \34475 , 1'b1 );
or \U$26366 ( \34477 , \34476 , 1'b0 );
buf \U$26367 ( \34478 , \34477 );
_DC r23ab2_GF_IsGateDCbyConstraint ( \34479_nR23ab2 , \34478 , \21944 );
buf \U$26368 ( \34480 , \34479_nR23ab2 );
not \U$26369 ( \34481 , \32666 );
and \U$26370 ( \34482 , RIe128258_5780, \34481 );
not \U$26371 ( \34483 , RIe128258_5780);
or \U$26372 ( \34484 , \34483 , \33966 );
not \U$26373 ( \34485 , \34303 );
and \U$26374 ( \34486 , \33265 , \34485 );
not \U$26375 ( \34487 , \34486 );
not \U$26376 ( \34488 , \33262 );
not \U$26377 ( \34489 , \33975 );
or \U$26378 ( \34490 , \34488 , \34489 );
nand \U$26379 ( \34491 , \34484 , \34487 , \34490 );
and \U$26380 ( \34492 , \34491 , \32666 );
or \U$26381 ( \34493 , \34482 , \34492 );
and \U$26383 ( \34494 , \34493 , 1'b1 );
or \U$26385 ( \34495 , \34494 , 1'b0 );
buf \U$26386 ( \34496 , \34495 );
_DC r23ab4_GF_IsGateDCbyConstraint ( \34497_nR23ab4 , \34496 , \21944 );
buf \U$26387 ( \34498 , \34497_nR23ab4 );
not \U$26388 ( \34499 , \33336 );
and \U$26389 ( \34500 , RIe12b930_5781, \34499 );
not \U$26390 ( \34501 , RIe12b930_5781);
or \U$26391 ( \34502 , \34501 , \33966 );
not \U$26392 ( \34503 , \34303 );
and \U$26393 ( \34504 , \33284 , \34503 );
not \U$26394 ( \34505 , \34504 );
not \U$26395 ( \34506 , \33281 );
not \U$26396 ( \34507 , \33975 );
or \U$26397 ( \34508 , \34506 , \34507 );
nand \U$26398 ( \34509 , \34502 , \34505 , \34508 );
and \U$26399 ( \34510 , \34509 , \33336 );
or \U$26400 ( \34511 , \34500 , \34510 );
and \U$26402 ( \34512 , \34511 , 1'b1 );
or \U$26404 ( \34513 , \34512 , 1'b0 );
buf \U$26405 ( \34514 , \34513 );
_DC r23ab6_GF_IsGateDCbyConstraint ( \34515_nR23ab6 , \34514 , \21944 );
buf \U$26406 ( \34516 , \34515_nR23ab6 );
not \U$26407 ( \34517 , \33336 );
and \U$26408 ( \34518 , RIe12e1f8_5782, \34517 );
not \U$26409 ( \34519 , RIe12e1f8_5782);
or \U$26410 ( \34520 , \34519 , \33966 );
not \U$26411 ( \34521 , \33991 );
and \U$26412 ( \34522 , \33305 , \34521 );
not \U$26413 ( \34523 , \34522 );
not \U$26414 ( \34524 , \33303 );
not \U$26415 ( \34525 , \33974 );
or \U$26416 ( \34526 , \34524 , \34525 );
nand \U$26417 ( \34527 , \34520 , \34523 , \34526 );
and \U$26418 ( \34528 , \34527 , \33336 );
or \U$26419 ( \34529 , \34518 , \34528 );
and \U$26421 ( \34530 , \34529 , 1'b1 );
or \U$26423 ( \34531 , \34530 , 1'b0 );
buf \U$26424 ( \34532 , \34531 );
_DC r23aba_GF_IsGateDCbyConstraint ( \34533_nR23aba , \34532 , \21944 );
buf \U$26425 ( \34534 , \34533_nR23aba );
not \U$26426 ( \34535 , \33568 );
and \U$26427 ( \34536 , RIe1308e0_5783, \34535 );
not \U$26428 ( \34537 , RIe1308e0_5783);
or \U$26429 ( \34538 , \34537 , \33966 );
not \U$26430 ( \34539 , \33969 );
and \U$26431 ( \34540 , \33324 , \34539 );
not \U$26432 ( \34541 , \34540 );
not \U$26433 ( \34542 , \33321 );
not \U$26434 ( \34543 , \33975 );
or \U$26435 ( \34544 , \34542 , \34543 );
nand \U$26436 ( \34545 , \34538 , \34541 , \34544 );
and \U$26437 ( \34546 , \34545 , \33568 );
or \U$26438 ( \34547 , \34536 , \34546 );
and \U$26440 ( \34548 , \34547 , 1'b1 );
or \U$26442 ( \34549 , \34548 , 1'b0 );
buf \U$26443 ( \34550 , \34549 );
_DC r23abc_GF_IsGateDCbyConstraint ( \34551_nR23abc , \34550 , \21944 );
buf \U$26444 ( \34552 , \34551_nR23abc );
not \U$26445 ( \34553 , \33874 );
and \U$26446 ( \34554 , RIe132398_5784, \34553 );
not \U$26447 ( \34555 , RIe132398_5784);
or \U$26448 ( \34556 , \34555 , \34047 );
not \U$26449 ( \34557 , \33991 );
and \U$26450 ( \34558 , \33344 , \34557 );
not \U$26451 ( \34559 , \34558 );
not \U$26452 ( \34560 , \33341 );
not \U$26453 ( \34561 , \33975 );
or \U$26454 ( \34562 , \34560 , \34561 );
nand \U$26455 ( \34563 , \34556 , \34559 , \34562 );
and \U$26456 ( \34564 , \34563 , \33874 );
or \U$26457 ( \34565 , \34554 , \34564 );
and \U$26459 ( \34566 , \34565 , 1'b1 );
or \U$26461 ( \34567 , \34566 , 1'b0 );
buf \U$26462 ( \34568 , \34567 );
_DC r23abe_GF_IsGateDCbyConstraint ( \34569_nR23abe , \34568 , \21944 );
buf \U$26463 ( \34570 , \34569_nR23abe );
not \U$26464 ( \34571 , \33874 );
and \U$26465 ( \34572 , RIe134300_5785, \34571 );
not \U$26466 ( \34573 , RIe134300_5785);
or \U$26467 ( \34574 , \34573 , \33964 );
not \U$26468 ( \34575 , \34028 );
and \U$26469 ( \34576 , \33363 , \34575 );
not \U$26470 ( \34577 , \34576 );
not \U$26471 ( \34578 , \33360 );
not \U$26472 ( \34579 , \33974 );
or \U$26473 ( \34580 , \34578 , \34579 );
nand \U$26474 ( \34581 , \34574 , \34577 , \34580 );
and \U$26475 ( \34582 , \34581 , \33874 );
or \U$26476 ( \34583 , \34572 , \34582 );
and \U$26478 ( \34584 , \34583 , 1'b1 );
or \U$26480 ( \34585 , \34584 , 1'b0 );
buf \U$26481 ( \34586 , \34585 );
_DC r23ac0_GF_IsGateDCbyConstraint ( \34587_nR23ac0 , \34586 , \21944 );
buf \U$26482 ( \34588 , \34587_nR23ac0 );
not \U$26483 ( \34589 , \33568 );
and \U$26484 ( \34590 , RIe135ae8_5786, \34589 );
not \U$26485 ( \34591 , RIe135ae8_5786);
or \U$26486 ( \34592 , \34591 , \33964 );
not \U$26487 ( \34593 , \34086 );
and \U$26488 ( \34594 , \33382 , \34593 );
not \U$26489 ( \34595 , \34594 );
not \U$26490 ( \34596 , \33379 );
not \U$26491 ( \34597 , \33975 );
or \U$26492 ( \34598 , \34596 , \34597 );
nand \U$26493 ( \34599 , \34592 , \34595 , \34598 );
and \U$26494 ( \34600 , \34599 , \33568 );
or \U$26495 ( \34601 , \34590 , \34600 );
and \U$26497 ( \34602 , \34601 , 1'b1 );
or \U$26499 ( \34603 , \34602 , 1'b0 );
buf \U$26500 ( \34604 , \34603 );
_DC r23ac2_GF_IsGateDCbyConstraint ( \34605_nR23ac2 , \34604 , \21944 );
buf \U$26501 ( \34606 , \34605_nR23ac2 );
not \U$26502 ( \34607 , \33336 );
and \U$26503 ( \34608 , RIe137258_5787, \34607 );
not \U$26504 ( \34609 , RIe137258_5787);
or \U$26505 ( \34610 , \34609 , \33989 );
not \U$26506 ( \34611 , \33969 );
and \U$26507 ( \34612 , \33402 , \34611 );
not \U$26508 ( \34613 , \34612 );
not \U$26509 ( \34614 , \33399 );
not \U$26510 ( \34615 , \33975 );
or \U$26511 ( \34616 , \34614 , \34615 );
nand \U$26512 ( \34617 , \34610 , \34613 , \34616 );
and \U$26513 ( \34618 , \34617 , \33336 );
or \U$26514 ( \34619 , \34608 , \34618 );
and \U$26516 ( \34620 , \34619 , 1'b1 );
or \U$26518 ( \34621 , \34620 , 1'b0 );
buf \U$26519 ( \34622 , \34621 );
_DC r23ac4_GF_IsGateDCbyConstraint ( \34623_nR23ac4 , \34622 , \21944 );
buf \U$26520 ( \34624 , \34623_nR23ac4 );
not \U$26521 ( \34625 , \32864 );
and \U$26522 ( \34626 , RIe138608_5788, \34625 );
not \U$26523 ( \34627 , RIe138608_5788);
or \U$26524 ( \34628 , \34627 , \33989 );
not \U$26525 ( \34629 , \33969 );
and \U$26526 ( \34630 , \33422 , \34629 );
not \U$26527 ( \34631 , \34630 );
not \U$26528 ( \34632 , \33419 );
not \U$26529 ( \34633 , \34033 );
or \U$26530 ( \34634 , \34632 , \34633 );
nand \U$26531 ( \34635 , \34628 , \34631 , \34634 );
and \U$26532 ( \34636 , \34635 , \32864 );
or \U$26533 ( \34637 , \34626 , \34636 );
and \U$26535 ( \34638 , \34637 , 1'b1 );
or \U$26537 ( \34639 , \34638 , 1'b0 );
buf \U$26538 ( \34640 , \34639 );
_DC r23ac6_GF_IsGateDCbyConstraint ( \34641_nR23ac6 , \34640 , \21944 );
buf \U$26539 ( \34642 , \34641_nR23ac6 );
not \U$26540 ( \34643 , \34318 );
and \U$26541 ( \34644 , RIe139850_5789, \34643 );
not \U$26542 ( \34645 , RIe139850_5789);
or \U$26543 ( \34646 , \34645 , \33964 );
not \U$26544 ( \34647 , \34028 );
and \U$26545 ( \34648 , \33440 , \34647 );
not \U$26546 ( \34649 , \34648 );
not \U$26547 ( \34650 , \33438 );
not \U$26548 ( \34651 , \33974 );
or \U$26549 ( \34652 , \34650 , \34651 );
nand \U$26550 ( \34653 , \34646 , \34649 , \34652 );
and \U$26551 ( \34654 , \34653 , \34318 );
or \U$26552 ( \34655 , \34644 , \34654 );
and \U$26554 ( \34656 , \34655 , 1'b1 );
or \U$26556 ( \34657 , \34656 , 1'b0 );
buf \U$26557 ( \34658 , \34657 );
_DC r23ac8_GF_IsGateDCbyConstraint ( \34659_nR23ac8 , \34658 , \21944 );
buf \U$26558 ( \34660 , \34659_nR23ac8 );
buf \U$26559 ( \34661 , \32841 );
not \U$26560 ( \34662 , \34661 );
and \U$26561 ( \34663 , RIe13ab88_5790, \34662 );
not \U$26562 ( \34664 , RIe13ab88_5790);
or \U$26563 ( \34665 , \34664 , \34047 );
not \U$26564 ( \34666 , \34086 );
and \U$26565 ( \34667 , \33459 , \34666 );
not \U$26566 ( \34668 , \34667 );
not \U$26567 ( \34669 , \33456 );
not \U$26568 ( \34670 , \33975 );
or \U$26569 ( \34671 , \34669 , \34670 );
nand \U$26570 ( \34672 , \34665 , \34668 , \34671 );
and \U$26571 ( \34673 , \34672 , \34661 );
or \U$26572 ( \34674 , \34663 , \34673 );
and \U$26574 ( \34675 , \34674 , 1'b1 );
or \U$26576 ( \34676 , \34675 , 1'b0 );
buf \U$26577 ( \34677 , \34676 );
_DC r23aca_GF_IsGateDCbyConstraint ( \34678_nR23aca , \34677 , \21944 );
buf \U$26578 ( \34679 , \34678_nR23aca );
not \U$26579 ( \34680 , \34661 );
and \U$26580 ( \34681 , RIe13c028_5791, \34680 );
not \U$26581 ( \34682 , RIe13c028_5791);
or \U$26582 ( \34683 , \34682 , \33966 );
not \U$26583 ( \34684 , \33969 );
and \U$26584 ( \34685 , \33478 , \34684 );
not \U$26585 ( \34686 , \34685 );
not \U$26586 ( \34687 , \33475 );
not \U$26587 ( \34688 , \33975 );
or \U$26588 ( \34689 , \34687 , \34688 );
nand \U$26589 ( \34690 , \34683 , \34686 , \34689 );
and \U$26590 ( \34691 , \34690 , \34661 );
or \U$26591 ( \34692 , \34681 , \34691 );
and \U$26593 ( \34693 , \34692 , 1'b1 );
or \U$26595 ( \34694 , \34693 , 1'b0 );
buf \U$26596 ( \34695 , \34694 );
_DC r23acc_GF_IsGateDCbyConstraint ( \34696_nR23acc , \34695 , \21944 );
buf \U$26597 ( \34697 , \34696_nR23acc );
buf \U$26598 ( \34698 , \32665 );
not \U$26599 ( \34699 , \34698 );
and \U$26600 ( \34700 , RIe13d5b8_5792, \34699 );
not \U$26601 ( \34701 , RIe13d5b8_5792);
or \U$26602 ( \34702 , \34701 , \33966 );
not \U$26603 ( \34703 , \34086 );
and \U$26604 ( \34704 , \33497 , \34703 );
not \U$26605 ( \34705 , \34704 );
not \U$26606 ( \34706 , \33494 );
not \U$26607 ( \34707 , \33974 );
or \U$26608 ( \34708 , \34706 , \34707 );
nand \U$26609 ( \34709 , \34702 , \34705 , \34708 );
and \U$26610 ( \34710 , \34709 , \34698 );
or \U$26611 ( \34711 , \34700 , \34710 );
and \U$26613 ( \34712 , \34711 , 1'b1 );
or \U$26615 ( \34713 , \34712 , 1'b0 );
buf \U$26616 ( \34714 , \34713 );
_DC r23ad0_GF_IsGateDCbyConstraint ( \34715_nR23ad0 , \34714 , \21944 );
buf \U$26617 ( \34716 , \34715_nR23ad0 );
not \U$26618 ( \34717 , \32864 );
and \U$26619 ( \34718 , RIe13ead0_5793, \34717 );
not \U$26620 ( \34719 , RIe13ead0_5793);
or \U$26621 ( \34720 , \34719 , \34047 );
not \U$26622 ( \34721 , \34028 );
and \U$26623 ( \34722 , \33517 , \34721 );
not \U$26624 ( \34723 , \34722 );
not \U$26625 ( \34724 , \33514 );
not \U$26626 ( \34725 , \34071 );
or \U$26627 ( \34726 , \34724 , \34725 );
nand \U$26628 ( \34727 , \34720 , \34723 , \34726 );
and \U$26629 ( \34728 , \34727 , \32864 );
or \U$26630 ( \34729 , \34718 , \34728 );
and \U$26632 ( \34730 , \34729 , 1'b1 );
or \U$26634 ( \34731 , \34730 , 1'b0 );
buf \U$26635 ( \34732 , \34731 );
_DC r23ad2_GF_IsGateDCbyConstraint ( \34733_nR23ad2 , \34732 , \21944 );
buf \U$26636 ( \34734 , \34733_nR23ad2 );
not \U$26637 ( \34735 , \34661 );
and \U$26638 ( \34736 , RIe13fef8_5794, \34735 );
not \U$26639 ( \34737 , RIe13fef8_5794);
or \U$26640 ( \34738 , \34737 , \33989 );
not \U$26641 ( \34739 , \33991 );
and \U$26642 ( \34740 , \33537 , \34739 );
not \U$26643 ( \34741 , \34740 );
not \U$26644 ( \34742 , \33534 );
not \U$26645 ( \34743 , \34033 );
or \U$26646 ( \34744 , \34742 , \34743 );
nand \U$26647 ( \34745 , \34738 , \34741 , \34744 );
and \U$26648 ( \34746 , \34745 , \34661 );
or \U$26649 ( \34747 , \34736 , \34746 );
and \U$26651 ( \34748 , \34747 , 1'b1 );
or \U$26653 ( \34749 , \34748 , 1'b0 );
buf \U$26654 ( \34750 , \34749 );
_DC r23ad4_GF_IsGateDCbyConstraint ( \34751_nR23ad4 , \34750 , \21944 );
buf \U$26655 ( \34752 , \34751_nR23ad4 );
not \U$26656 ( \34753 , \33568 );
and \U$26657 ( \34754 , RIe141230_5795, \34753 );
not \U$26658 ( \34755 , RIe141230_5795);
or \U$26659 ( \34756 , \34755 , \33966 );
not \U$26660 ( \34757 , \34303 );
and \U$26661 ( \34758 , \33556 , \34757 );
not \U$26662 ( \34759 , \34758 );
not \U$26663 ( \34760 , \33553 );
not \U$26664 ( \34761 , \34071 );
or \U$26665 ( \34762 , \34760 , \34761 );
nand \U$26666 ( \34763 , \34756 , \34759 , \34762 );
and \U$26667 ( \34764 , \34763 , \33568 );
or \U$26668 ( \34765 , \34754 , \34764 );
and \U$26670 ( \34766 , \34765 , 1'b1 );
or \U$26672 ( \34767 , \34766 , 1'b0 );
buf \U$26673 ( \34768 , \34767 );
_DC r23ad6_GF_IsGateDCbyConstraint ( \34769_nR23ad6 , \34768 , \21944 );
buf \U$26674 ( \34770 , \34769_nR23ad6 );
not \U$26675 ( \34771 , \34661 );
and \U$26676 ( \34772 , RIe142568_5796, \34771 );
not \U$26677 ( \34773 , RIe142568_5796);
or \U$26678 ( \34774 , \34773 , \34047 );
not \U$26679 ( \34775 , \34303 );
and \U$26680 ( \34776 , \33576 , \34775 );
not \U$26681 ( \34777 , \34776 );
not \U$26682 ( \34778 , \33574 );
not \U$26683 ( \34779 , \33974 );
or \U$26684 ( \34780 , \34778 , \34779 );
nand \U$26685 ( \34781 , \34774 , \34777 , \34780 );
and \U$26686 ( \34782 , \34781 , \34661 );
or \U$26687 ( \34783 , \34772 , \34782 );
and \U$26689 ( \34784 , \34783 , 1'b1 );
or \U$26691 ( \34785 , \34784 , 1'b0 );
buf \U$26692 ( \34786 , \34785 );
_DC r23ad8_GF_IsGateDCbyConstraint ( \34787_nR23ad8 , \34786 , \21944 );
buf \U$26693 ( \34788 , \34787_nR23ad8 );
not \U$26694 ( \34789 , \34661 );
and \U$26695 ( \34790 , RIe1434e0_5797, \34789 );
not \U$26696 ( \34791 , RIe1434e0_5797);
or \U$26697 ( \34792 , \34791 , \33989 );
not \U$26698 ( \34793 , \33991 );
and \U$26699 ( \34794 , \33594 , \34793 );
not \U$26700 ( \34795 , \34794 );
not \U$26701 ( \34796 , \33592 );
not \U$26702 ( \34797 , \34071 );
or \U$26703 ( \34798 , \34796 , \34797 );
nand \U$26704 ( \34799 , \34792 , \34795 , \34798 );
and \U$26705 ( \34800 , \34799 , \34661 );
or \U$26706 ( \34801 , \34790 , \34800 );
and \U$26708 ( \34802 , \34801 , 1'b1 );
or \U$26710 ( \34803 , \34802 , 1'b0 );
buf \U$26711 ( \34804 , \34803 );
_DC r23ada_GF_IsGateDCbyConstraint ( \34805_nR23ada , \34804 , \21944 );
buf \U$26712 ( \34806 , \34805_nR23ada );
not \U$26713 ( \34807 , \33296 );
and \U$26714 ( \34808 , RIe144638_5798, \34807 );
not \U$26715 ( \34809 , RIe144638_5798);
or \U$26716 ( \34810 , \34809 , \34047 );
not \U$26717 ( \34811 , \34086 );
and \U$26718 ( \34812 , \33612 , \34811 );
not \U$26719 ( \34813 , \34812 );
not \U$26720 ( \34814 , \33610 );
not \U$26721 ( \34815 , \33975 );
or \U$26722 ( \34816 , \34814 , \34815 );
nand \U$26723 ( \34817 , \34810 , \34813 , \34816 );
and \U$26724 ( \34818 , \34817 , \33296 );
or \U$26725 ( \34819 , \34808 , \34818 );
and \U$26727 ( \34820 , \34819 , 1'b1 );
or \U$26729 ( \34821 , \34820 , 1'b0 );
buf \U$26730 ( \34822 , \34821 );
_DC r23adc_GF_IsGateDCbyConstraint ( \34823_nR23adc , \34822 , \21944 );
buf \U$26731 ( \34824 , \34823_nR23adc );
not \U$26732 ( \34825 , \32864 );
and \U$26733 ( \34826 , RIe145880_5799, \34825 );
not \U$26734 ( \34827 , RIe145880_5799);
or \U$26735 ( \34828 , \34827 , \33964 );
not \U$26736 ( \34829 , \33969 );
and \U$26737 ( \34830 , \33632 , \34829 );
not \U$26738 ( \34831 , \34830 );
not \U$26739 ( \34832 , \33629 );
not \U$26740 ( \34833 , \34071 );
or \U$26741 ( \34834 , \34832 , \34833 );
nand \U$26742 ( \34835 , \34828 , \34831 , \34834 );
and \U$26743 ( \34836 , \34835 , \32864 );
or \U$26744 ( \34837 , \34826 , \34836 );
and \U$26746 ( \34838 , \34837 , 1'b1 );
or \U$26748 ( \34839 , \34838 , 1'b0 );
buf \U$26749 ( \34840 , \34839 );
_DC r23ade_GF_IsGateDCbyConstraint ( \34841_nR23ade , \34840 , \21944 );
buf \U$26750 ( \34842 , \34841_nR23ade );
not \U$26751 ( \34843 , \32864 );
and \U$26752 ( \34844 , RIe146ac8_5800, \34843 );
not \U$26753 ( \34845 , RIe146ac8_5800);
or \U$26754 ( \34846 , \34845 , \33989 );
not \U$26755 ( \34847 , \34303 );
and \U$26756 ( \34848 , \33651 , \34847 );
not \U$26757 ( \34849 , \34848 );
not \U$26758 ( \34850 , \33648 );
not \U$26759 ( \34851 , \34033 );
or \U$26760 ( \34852 , \34850 , \34851 );
nand \U$26761 ( \34853 , \34846 , \34849 , \34852 );
and \U$26762 ( \34854 , \34853 , \32864 );
or \U$26763 ( \34855 , \34844 , \34854 );
and \U$26765 ( \34856 , \34855 , 1'b1 );
or \U$26767 ( \34857 , \34856 , 1'b0 );
buf \U$26768 ( \34858 , \34857 );
_DC r23ae0_GF_IsGateDCbyConstraint ( \34859_nR23ae0 , \34858 , \21944 );
buf \U$26769 ( \34860 , \34859_nR23ae0 );
not \U$26770 ( \34861 , \32841 );
and \U$26771 ( \34862 , RIe1486e8_5801, \34861 );
not \U$26772 ( \34863 , RIe1486e8_5801);
or \U$26773 ( \34864 , \34863 , \33966 );
not \U$26774 ( \34865 , \34303 );
and \U$26775 ( \34866 , \33671 , \34865 );
not \U$26776 ( \34867 , \34866 );
not \U$26777 ( \34868 , \33668 );
not \U$26778 ( \34869 , \34071 );
or \U$26779 ( \34870 , \34868 , \34869 );
nand \U$26780 ( \34871 , \34864 , \34867 , \34870 );
and \U$26781 ( \34872 , \34871 , \32841 );
or \U$26782 ( \34873 , \34862 , \34872 );
and \U$26784 ( \34874 , \34873 , 1'b1 );
or \U$26786 ( \34875 , \34874 , 1'b0 );
buf \U$26787 ( \34876 , \34875 );
_DC r23ae2_GF_IsGateDCbyConstraint ( \34877_nR23ae2 , \34876 , \21944 );
buf \U$26788 ( \34878 , \34877_nR23ae2 );
not \U$26789 ( \34879 , \32864 );
and \U$26790 ( \34880 , RIe149f48_5802, \34879 );
not \U$26791 ( \34881 , RIe149f48_5802);
or \U$26792 ( \34882 , \34881 , \33964 );
not \U$26793 ( \34883 , \33991 );
and \U$26794 ( \34884 , \33691 , \34883 );
not \U$26795 ( \34885 , \34884 );
not \U$26796 ( \34886 , \33688 );
not \U$26797 ( \34887 , \34033 );
or \U$26798 ( \34888 , \34886 , \34887 );
nand \U$26799 ( \34889 , \34882 , \34885 , \34888 );
and \U$26800 ( \34890 , \34889 , \32864 );
or \U$26801 ( \34891 , \34880 , \34890 );
and \U$26803 ( \34892 , \34891 , 1'b1 );
or \U$26805 ( \34893 , \34892 , 1'b0 );
buf \U$26806 ( \34894 , \34893 );
_DC r23ae6_GF_IsGateDCbyConstraint ( \34895_nR23ae6 , \34894 , \21944 );
buf \U$26807 ( \34896 , \34895_nR23ae6 );
not \U$26808 ( \34897 , \34661 );
and \U$26809 ( \34898 , RIe14b550_5803, \34897 );
not \U$26810 ( \34899 , RIe14b550_5803);
or \U$26811 ( \34900 , \34899 , \34047 );
not \U$26812 ( \34901 , \34028 );
and \U$26813 ( \34902 , \33709 , \34901 );
not \U$26814 ( \34903 , \34902 );
not \U$26815 ( \34904 , \33707 );
not \U$26816 ( \34905 , \34071 );
or \U$26817 ( \34906 , \34904 , \34905 );
nand \U$26818 ( \34907 , \34900 , \34903 , \34906 );
and \U$26819 ( \34908 , \34907 , \34661 );
or \U$26820 ( \34909 , \34898 , \34908 );
and \U$26822 ( \34910 , \34909 , 1'b1 );
or \U$26824 ( \34911 , \34910 , 1'b0 );
buf \U$26825 ( \34912 , \34911 );
_DC r23ae8_GF_IsGateDCbyConstraint ( \34913_nR23ae8 , \34912 , \21944 );
buf \U$26826 ( \34914 , \34913_nR23ae8 );
buf \U$26827 ( \34915 , \32665 );
buf \U$26828 ( \34916 , \34915 );
not \U$26829 ( \34917 , \34916 );
and \U$26830 ( \34918 , RIe14c978_5804, \34917 );
not \U$26831 ( \34919 , RIe14c978_5804);
or \U$26832 ( \34920 , \34919 , \33964 );
not \U$26833 ( \34921 , \34086 );
and \U$26834 ( \34922 , \33728 , \34921 );
not \U$26835 ( \34923 , \34922 );
not \U$26836 ( \34924 , \33725 );
not \U$26837 ( \34925 , \34071 );
or \U$26838 ( \34926 , \34924 , \34925 );
nand \U$26839 ( \34927 , \34920 , \34923 , \34926 );
and \U$26840 ( \34928 , \34927 , \34916 );
or \U$26841 ( \34929 , \34918 , \34928 );
and \U$26843 ( \34930 , \34929 , 1'b1 );
or \U$26845 ( \34931 , \34930 , 1'b0 );
buf \U$26846 ( \34932 , \34931 );
_DC r23aea_GF_IsGateDCbyConstraint ( \34933_nR23aea , \34932 , \21944 );
buf \U$26847 ( \34934 , \34933_nR23aea );
not \U$26848 ( \34935 , \32864 );
and \U$26849 ( \34936 , RIe14e430_5805, \34935 );
not \U$26850 ( \34937 , RIe14e430_5805);
or \U$26851 ( \34938 , \34937 , \33966 );
not \U$26852 ( \34939 , \34086 );
and \U$26853 ( \34940 , \33746 , \34939 );
not \U$26854 ( \34941 , \34940 );
not \U$26855 ( \34942 , \33744 );
not \U$26856 ( \34943 , \34033 );
or \U$26857 ( \34944 , \34942 , \34943 );
nand \U$26858 ( \34945 , \34938 , \34941 , \34944 );
and \U$26859 ( \34946 , \34945 , \32864 );
or \U$26860 ( \34947 , \34936 , \34946 );
and \U$26862 ( \34948 , \34947 , 1'b1 );
or \U$26864 ( \34949 , \34948 , 1'b0 );
buf \U$26865 ( \34950 , \34949 );
_DC r23aec_GF_IsGateDCbyConstraint ( \34951_nR23aec , \34950 , \21944 );
buf \U$26866 ( \34952 , \34951_nR23aec );
not \U$26867 ( \34953 , \32864 );
and \U$26868 ( \34954 , RIe0865e8_5806, \34953 );
not \U$26869 ( \34955 , RIe0865e8_5806);
or \U$26870 ( \34956 , \34955 , \33989 );
not \U$26871 ( \34957 , \34028 );
and \U$26872 ( \34958 , \33766 , \34957 );
not \U$26873 ( \34959 , \34958 );
not \U$26874 ( \34960 , \33763 );
not \U$26875 ( \34961 , \34071 );
or \U$26876 ( \34962 , \34960 , \34961 );
nand \U$26877 ( \34963 , \34956 , \34959 , \34962 );
and \U$26878 ( \34964 , \34963 , \32864 );
or \U$26879 ( \34965 , \34954 , \34964 );
and \U$26881 ( \34966 , \34965 , 1'b1 );
or \U$26883 ( \34967 , \34966 , 1'b0 );
buf \U$26884 ( \34968 , \34967 );
_DC r23aee_GF_IsGateDCbyConstraint ( \34969_nR23aee , \34968 , \21944 );
buf \U$26885 ( \34970 , \34969_nR23aee );
not \U$26886 ( \34971 , \34916 );
and \U$26887 ( \34972 , RIe087f38_5807, \34971 );
not \U$26888 ( \34973 , RIe087f38_5807);
or \U$26889 ( \34974 , \34973 , \33964 );
not \U$26890 ( \34975 , \33969 );
and \U$26891 ( \34976 , \33786 , \34975 );
not \U$26892 ( \34977 , \34976 );
not \U$26893 ( \34978 , \33783 );
not \U$26894 ( \34979 , \34033 );
or \U$26895 ( \34980 , \34978 , \34979 );
nand \U$26896 ( \34981 , \34974 , \34977 , \34980 );
and \U$26897 ( \34982 , \34981 , \34916 );
or \U$26898 ( \34983 , \34972 , \34982 );
and \U$26900 ( \34984 , \34983 , 1'b1 );
or \U$26902 ( \34985 , \34984 , 1'b0 );
buf \U$26903 ( \34986 , \34985 );
_DC r23af0_GF_IsGateDCbyConstraint ( \34987_nR23af0 , \34986 , \21944 );
buf \U$26904 ( \34988 , \34987_nR23af0 );
not \U$26905 ( \34989 , \34661 );
and \U$26906 ( \34990 , RIe089db0_5808, \34989 );
not \U$26907 ( \34991 , RIe089db0_5808);
or \U$26908 ( \34992 , \34991 , \33966 );
not \U$26909 ( \34993 , \33991 );
and \U$26910 ( \34994 , \33805 , \34993 );
not \U$26911 ( \34995 , \34994 );
not \U$26912 ( \34996 , \33802 );
not \U$26913 ( \34997 , \34033 );
or \U$26914 ( \34998 , \34996 , \34997 );
nand \U$26915 ( \34999 , \34992 , \34995 , \34998 );
and \U$26916 ( \35000 , \34999 , \34661 );
or \U$26917 ( \35001 , \34990 , \35000 );
and \U$26919 ( \35002 , \35001 , 1'b1 );
or \U$26921 ( \35003 , \35002 , 1'b0 );
buf \U$26922 ( \35004 , \35003 );
_DC r23af2_GF_IsGateDCbyConstraint ( \35005_nR23af2 , \35004 , \21944 );
buf \U$26923 ( \35006 , \35005_nR23af2 );
not \U$26924 ( \35007 , \34661 );
and \U$26925 ( \35008 , RIe08b7f0_5809, \35007 );
not \U$26926 ( \35009 , RIe08b7f0_5809);
or \U$26927 ( \35010 , \35009 , \34047 );
not \U$26928 ( \35011 , \34028 );
and \U$26929 ( \35012 , \33824 , \35011 );
not \U$26930 ( \35013 , \35012 );
not \U$26931 ( \35014 , \33821 );
not \U$26932 ( \35015 , \34071 );
or \U$26933 ( \35016 , \35014 , \35015 );
nand \U$26934 ( \35017 , \35010 , \35013 , \35016 );
and \U$26935 ( \35018 , \35017 , \34661 );
or \U$26936 ( \35019 , \35008 , \35018 );
and \U$26938 ( \35020 , \35019 , 1'b1 );
or \U$26940 ( \35021 , \35020 , 1'b0 );
buf \U$26941 ( \35022 , \35021 );
_DC r23af4_GF_IsGateDCbyConstraint ( \35023_nR23af4 , \35022 , \21944 );
buf \U$26942 ( \35024 , \35023_nR23af4 );
not \U$26943 ( \35025 , \34916 );
and \U$26944 ( \35026 , RIe08d578_5810, \35025 );
not \U$26945 ( \35027 , RIe08d578_5810);
or \U$26946 ( \35028 , \35027 , \33989 );
not \U$26947 ( \35029 , \34086 );
and \U$26948 ( \35030 , \33843 , \35029 );
not \U$26949 ( \35031 , \35030 );
not \U$26950 ( \35032 , \33840 );
not \U$26951 ( \35033 , \34071 );
or \U$26952 ( \35034 , \35032 , \35033 );
nand \U$26953 ( \35035 , \35028 , \35031 , \35034 );
and \U$26954 ( \35036 , \35035 , \34916 );
or \U$26955 ( \35037 , \35026 , \35036 );
and \U$26957 ( \35038 , \35037 , 1'b1 );
or \U$26959 ( \35039 , \35038 , 1'b0 );
buf \U$26960 ( \35040 , \35039 );
_DC r23af6_GF_IsGateDCbyConstraint ( \35041_nR23af6 , \35040 , \21944 );
buf \U$26961 ( \35042 , \35041_nR23af6 );
not \U$26962 ( \35043 , \32864 );
and \U$26963 ( \35044 , RIe08f120_5811, \35043 );
not \U$26964 ( \35045 , RIe08f120_5811);
or \U$26965 ( \35046 , \35045 , \33964 );
not \U$26966 ( \35047 , \33991 );
and \U$26967 ( \35048 , \33862 , \35047 );
not \U$26968 ( \35049 , \35048 );
not \U$26969 ( \35050 , \33859 );
not \U$26970 ( \35051 , \34033 );
or \U$26971 ( \35052 , \35050 , \35051 );
nand \U$26972 ( \35053 , \35046 , \35049 , \35052 );
and \U$26973 ( \35054 , \35053 , \32864 );
or \U$26974 ( \35055 , \35044 , \35054 );
and \U$26976 ( \35056 , \35055 , 1'b1 );
or \U$26978 ( \35057 , \35056 , 1'b0 );
buf \U$26979 ( \35058 , \35057 );
_DC r23af8_GF_IsGateDCbyConstraint ( \35059_nR23af8 , \35058 , \21944 );
buf \U$26980 ( \35060 , \35059_nR23af8 );
not \U$26981 ( \35061 , \32864 );
and \U$26982 ( \35062 , RIe091100_5812, \35061 );
not \U$26983 ( \35063 , RIe091100_5812);
or \U$26984 ( \35064 , \35063 , \33966 );
not \U$26985 ( \35065 , \33969 );
and \U$26986 ( \35066 , \33882 , \35065 );
not \U$26987 ( \35067 , \35066 );
not \U$26988 ( \35068 , \33879 );
not \U$26989 ( \35069 , \34033 );
or \U$26990 ( \35070 , \35068 , \35069 );
nand \U$26991 ( \35071 , \35064 , \35067 , \35070 );
and \U$26992 ( \35072 , \35071 , \32864 );
or \U$26993 ( \35073 , \35062 , \35072 );
and \U$26995 ( \35074 , \35073 , 1'b1 );
or \U$26997 ( \35075 , \35074 , 1'b0 );
buf \U$26998 ( \35076 , \35075 );
_DC r23afc_GF_IsGateDCbyConstraint ( \35077_nR23afc , \35076 , \21944 );
buf \U$26999 ( \35078 , \35077_nR23afc );
not \U$27000 ( \35079 , \34916 );
and \U$27001 ( \35080 , RIe093248_5813, \35079 );
not \U$27002 ( \35081 , RIe093248_5813);
or \U$27003 ( \35082 , \35081 , \33966 );
not \U$27004 ( \35083 , \33969 );
and \U$27005 ( \35084 , \33902 , \35083 );
not \U$27006 ( \35085 , \35084 );
not \U$27007 ( \35086 , \33899 );
not \U$27008 ( \35087 , \34033 );
or \U$27009 ( \35088 , \35086 , \35087 );
nand \U$27010 ( \35089 , \35082 , \35085 , \35088 );
and \U$27011 ( \35090 , \35089 , \34916 );
or \U$27012 ( \35091 , \35080 , \35090 );
and \U$27014 ( \35092 , \35091 , 1'b1 );
or \U$27016 ( \35093 , \35092 , 1'b0 );
buf \U$27017 ( \35094 , \35093 );
_DC r23afe_GF_IsGateDCbyConstraint ( \35095_nR23afe , \35094 , \21944 );
buf \U$27018 ( \35096 , \35095_nR23afe );
not \U$27019 ( \35097 , \34661 );
and \U$27020 ( \35098 , RIe0950c0_5814, \35097 );
not \U$27021 ( \35099 , RIe0950c0_5814);
or \U$27022 ( \35100 , \35099 , \33989 );
not \U$27023 ( \35101 , \34303 );
and \U$27024 ( \35102 , \33921 , \35101 );
not \U$27025 ( \35103 , \35102 );
not \U$27026 ( \35104 , \33918 );
not \U$27027 ( \35105 , \34071 );
or \U$27028 ( \35106 , \35104 , \35105 );
nand \U$27029 ( \35107 , \35100 , \35103 , \35106 );
and \U$27030 ( \35108 , \35107 , \34661 );
or \U$27031 ( \35109 , \35098 , \35108 );
and \U$27033 ( \35110 , \35109 , 1'b1 );
or \U$27035 ( \35111 , \35110 , 1'b0 );
buf \U$27036 ( \35112 , \35111 );
_DC r23b00_GF_IsGateDCbyConstraint ( \35113_nR23b00 , \35112 , \21944 );
buf \U$27037 ( \35114 , \35113_nR23b00 );
not \U$27038 ( \35115 , \34916 );
and \U$27039 ( \35116 , RIe096998_5815, \35115 );
not \U$27040 ( \35117 , RIe096998_5815);
or \U$27041 ( \35118 , \35117 , \33966 );
not \U$27042 ( \35119 , \34086 );
and \U$27043 ( \35120 , \33940 , \35119 );
not \U$27044 ( \35121 , \35120 );
not \U$27045 ( \35122 , \33937 );
not \U$27046 ( \35123 , \34071 );
or \U$27047 ( \35124 , \35122 , \35123 );
nand \U$27048 ( \35125 , \35118 , \35121 , \35124 );
and \U$27049 ( \35126 , \35125 , \34916 );
or \U$27050 ( \35127 , \35116 , \35126 );
and \U$27052 ( \35128 , \35127 , 1'b1 );
or \U$27054 ( \35129 , \35128 , 1'b0 );
buf \U$27055 ( \35130 , \35129 );
_DC r23b02_GF_IsGateDCbyConstraint ( \35131_nR23b02 , \35130 , \21944 );
buf \U$27056 ( \35132 , \35131_nR23b02 );
not \U$27057 ( \35133 , \32864 );
and \U$27058 ( \35134 , RIe0986a8_5816, \35133 );
not \U$27059 ( \35135 , RIe0986a8_5816);
not \U$27060 ( \35136 , \32678 );
nor \U$27061 ( \35137 , \32680 , \35136 );
nand \U$27062 ( \35138 , \35137 , \32682 );
not \U$27063 ( \35139 , \35138 );
not \U$27064 ( \35140 , \32672 );
or \U$27065 ( \35141 , \32670 , \35140 );
not \U$27066 ( \35142 , \35141 );
nand \U$27067 ( \35143 , \32664 , \35142 );
not \U$27068 ( \35144 , \35143 );
or \U$27069 ( \35145 , \35139 , \35144 );
not \U$27070 ( \35146 , \35145 );
not \U$27071 ( \35147 , \35146 );
or \U$27072 ( \35148 , \35135 , \35147 );
not \U$27073 ( \35149 , \35138 );
not \U$27074 ( \35150 , \35149 );
not \U$27075 ( \35151 , \35150 );
and \U$27076 ( \35152 , \32694 , \35151 );
not \U$27077 ( \35153 , \35152 );
not \U$27078 ( \35154 , \35143 );
buf \U$27079 ( \35155 , \35154 );
not \U$27080 ( \35156 , \35155 );
or \U$27081 ( \35157 , \33973 , \35156 );
nand \U$27082 ( \35158 , \35148 , \35153 , \35157 );
and \U$27083 ( \35159 , \35158 , \32864 );
or \U$27084 ( \35160 , \35134 , \35159 );
and \U$27086 ( \35161 , \35160 , 1'b1 );
or \U$27088 ( \35162 , \35161 , 1'b0 );
buf \U$27089 ( \35163 , \35162 );
_DC r23b0c_GF_IsGateDCbyConstraint ( \35164_nR23b0c , \35163 , \21944 );
buf \U$27090 ( \35165 , \35164_nR23b0c );
not \U$27091 ( \35166 , \34916 );
and \U$27092 ( \35167 , RIe1cfd18_5817, \35166 );
not \U$27093 ( \35168 , RIe1cfd18_5817);
not \U$27094 ( \35169 , \35146 );
or \U$27095 ( \35170 , \35168 , \35169 );
not \U$27096 ( \35171 , \35150 );
and \U$27097 ( \35172 , \32722 , \35171 );
not \U$27098 ( \35173 , \35172 );
not \U$27099 ( \35174 , \35155 );
or \U$27100 ( \35175 , \33995 , \35174 );
nand \U$27101 ( \35176 , \35170 , \35173 , \35175 );
and \U$27102 ( \35177 , \35176 , \34916 );
or \U$27103 ( \35178 , \35167 , \35177 );
and \U$27105 ( \35179 , \35178 , 1'b1 );
or \U$27107 ( \35180 , \35179 , 1'b0 );
buf \U$27108 ( \35181 , \35180 );
_DC r23b22_GF_IsGateDCbyConstraint ( \35182_nR23b22 , \35181 , \21944 );
buf \U$27109 ( \35183 , \35182_nR23b22 );
not \U$27110 ( \35184 , \34661 );
and \U$27111 ( \35185 , RIe1ce080_5818, \35184 );
not \U$27112 ( \35186 , RIe1ce080_5818);
or \U$27113 ( \35187 , \35186 , \35169 );
not \U$27114 ( \35188 , \35139 );
not \U$27115 ( \35189 , \35188 );
and \U$27116 ( \35190 , \32743 , \35189 );
not \U$27117 ( \35191 , \35190 );
not \U$27118 ( \35192 , \35155 );
or \U$27119 ( \35193 , \34013 , \35192 );
nand \U$27120 ( \35194 , \35187 , \35191 , \35193 );
and \U$27121 ( \35195 , \35194 , \34661 );
or \U$27122 ( \35196 , \35185 , \35195 );
and \U$27124 ( \35197 , \35196 , 1'b1 );
or \U$27126 ( \35198 , \35197 , 1'b0 );
buf \U$27127 ( \35199 , \35198 );
_DC r23b38_GF_IsGateDCbyConstraint ( \35200_nR23b38 , \35199 , \21944 );
buf \U$27128 ( \35201 , \35200_nR23b38 );
not \U$27129 ( \35202 , \32864 );
and \U$27130 ( \35203 , RIe1cc550_5819, \35202 );
not \U$27131 ( \35204 , RIe1cc550_5819);
or \U$27132 ( \35205 , \35204 , \35169 );
not \U$27133 ( \35206 , \35150 );
and \U$27134 ( \35207 , \32764 , \35206 );
not \U$27135 ( \35208 , \35207 );
buf \U$27136 ( \35209 , \35154 );
not \U$27137 ( \35210 , \35209 );
or \U$27138 ( \35211 , \34032 , \35210 );
nand \U$27139 ( \35212 , \35205 , \35208 , \35211 );
and \U$27140 ( \35213 , \35212 , \32864 );
or \U$27141 ( \35214 , \35203 , \35213 );
and \U$27143 ( \35215 , \35214 , 1'b1 );
or \U$27145 ( \35216 , \35215 , 1'b0 );
buf \U$27146 ( \35217 , \35216 );
_DC r23b4e_GF_IsGateDCbyConstraint ( \35218_nR23b4e , \35217 , \21944 );
buf \U$27147 ( \35219 , \35218_nR23b4e );
not \U$27148 ( \35220 , \34916 );
and \U$27149 ( \35221 , RIe1ca048_5820, \35220 );
not \U$27150 ( \35222 , RIe1ca048_5820);
not \U$27151 ( \35223 , \35146 );
or \U$27152 ( \35224 , \35222 , \35223 );
not \U$27153 ( \35225 , \35188 );
and \U$27154 ( \35226 , \32786 , \35225 );
not \U$27155 ( \35227 , \35226 );
not \U$27156 ( \35228 , \35209 );
or \U$27157 ( \35229 , \34052 , \35228 );
nand \U$27158 ( \35230 , \35224 , \35227 , \35229 );
and \U$27159 ( \35231 , \35230 , \34916 );
or \U$27160 ( \35232 , \35221 , \35231 );
and \U$27162 ( \35233 , \35232 , 1'b1 );
or \U$27164 ( \35234 , \35233 , 1'b0 );
buf \U$27165 ( \35235 , \35234 );
_DC r23b64_GF_IsGateDCbyConstraint ( \35236_nR23b64 , \35235 , \21944 );
buf \U$27166 ( \35237 , \35236_nR23b64 );
not \U$27167 ( \35238 , \34661 );
and \U$27168 ( \35239 , RIe1c78e8_5821, \35238 );
not \U$27169 ( \35240 , RIe1c78e8_5821);
not \U$27170 ( \35241 , \35146 );
or \U$27171 ( \35242 , \35240 , \35241 );
not \U$27172 ( \35243 , \35149 );
not \U$27173 ( \35244 , \35243 );
and \U$27174 ( \35245 , \32806 , \35244 );
not \U$27175 ( \35246 , \35245 );
buf \U$27176 ( \35247 , \35154 );
not \U$27177 ( \35248 , \35247 );
or \U$27178 ( \35249 , \34070 , \35248 );
nand \U$27179 ( \35250 , \35242 , \35246 , \35249 );
and \U$27180 ( \35251 , \35250 , \34661 );
or \U$27181 ( \35252 , \35239 , \35251 );
and \U$27183 ( \35253 , \35252 , 1'b1 );
or \U$27185 ( \35254 , \35253 , 1'b0 );
buf \U$27186 ( \35255 , \35254 );
_DC r23b7a_GF_IsGateDCbyConstraint ( \35256_nR23b7a , \35255 , \21944 );
buf \U$27187 ( \35257 , \35256_nR23b7a );
not \U$27188 ( \35258 , \32864 );
and \U$27189 ( \35259 , RIe1c4f30_5822, \35258 );
not \U$27190 ( \35260 , RIe1c4f30_5822);
or \U$27191 ( \35261 , \35260 , \35169 );
not \U$27192 ( \35262 , \35188 );
and \U$27193 ( \35263 , \32829 , \35262 );
not \U$27194 ( \35264 , \35263 );
nand \U$27195 ( \35265 , \32827 , \35209 );
nand \U$27196 ( \35266 , \35261 , \35264 , \35265 );
and \U$27197 ( \35267 , \35266 , \32864 );
or \U$27198 ( \35268 , \35259 , \35267 );
and \U$27200 ( \35269 , \35268 , 1'b1 );
or \U$27202 ( \35270 , \35269 , 1'b0 );
buf \U$27203 ( \35271 , \35270 );
_DC r23b84_GF_IsGateDCbyConstraint ( \35272_nR23b84 , \35271 , \21944 );
buf \U$27204 ( \35273 , \35272_nR23b84 );
not \U$27205 ( \35274 , \34916 );
and \U$27206 ( \35275 , RIe1c26e0_5823, \35274 );
not \U$27207 ( \35276 , RIe1c26e0_5823);
or \U$27208 ( \35277 , \35276 , \35169 );
not \U$27209 ( \35278 , \35150 );
and \U$27210 ( \35279 , \32851 , \35278 );
not \U$27211 ( \35280 , \35279 );
not \U$27212 ( \35281 , \35247 );
or \U$27213 ( \35282 , \34108 , \35281 );
nand \U$27214 ( \35283 , \35277 , \35280 , \35282 );
and \U$27215 ( \35284 , \35283 , \34916 );
or \U$27216 ( \35285 , \35275 , \35284 );
and \U$27218 ( \35286 , \35285 , 1'b1 );
or \U$27220 ( \35287 , \35286 , 1'b0 );
buf \U$27221 ( \35288 , \35287 );
_DC r23b86_GF_IsGateDCbyConstraint ( \35289_nR23b86 , \35288 , \21944 );
buf \U$27222 ( \35290 , \35289_nR23b86 );
not \U$27223 ( \35291 , \34661 );
and \U$27224 ( \35292 , RIe1c0b38_5824, \35291 );
not \U$27225 ( \35293 , RIe1c0b38_5824);
or \U$27226 ( \35294 , \35293 , \35147 );
not \U$27227 ( \35295 , \35243 );
and \U$27228 ( \35296 , \32873 , \35295 );
not \U$27229 ( \35297 , \35296 );
not \U$27230 ( \35298 , \35209 );
or \U$27231 ( \35299 , \34126 , \35298 );
nand \U$27232 ( \35300 , \35294 , \35297 , \35299 );
and \U$27233 ( \35301 , \35300 , \34661 );
or \U$27234 ( \35302 , \35292 , \35301 );
and \U$27236 ( \35303 , \35302 , 1'b1 );
or \U$27238 ( \35304 , \35303 , 1'b0 );
buf \U$27239 ( \35305 , \35304 );
_DC r23b88_GF_IsGateDCbyConstraint ( \35306_nR23b88 , \35305 , \21944 );
buf \U$27240 ( \35307 , \35306_nR23b88 );
not \U$27241 ( \35308 , \32842 );
and \U$27242 ( \35309 , RIe1be9f0_5825, \35308 );
not \U$27243 ( \35310 , RIe1be9f0_5825);
not \U$27244 ( \35311 , \35146 );
or \U$27245 ( \35312 , \35310 , \35311 );
not \U$27246 ( \35313 , \35139 );
not \U$27247 ( \35314 , \35313 );
and \U$27248 ( \35315 , \32894 , \35314 );
not \U$27249 ( \35316 , \35315 );
not \U$27250 ( \35317 , \35209 );
or \U$27251 ( \35318 , \34144 , \35317 );
nand \U$27252 ( \35319 , \35312 , \35316 , \35318 );
and \U$27253 ( \35320 , \35319 , \32842 );
or \U$27254 ( \35321 , \35309 , \35320 );
and \U$27256 ( \35322 , \35321 , 1'b1 );
or \U$27258 ( \35323 , \35322 , 1'b0 );
buf \U$27259 ( \35324 , \35323 );
_DC r23b8a_GF_IsGateDCbyConstraint ( \35325_nR23b8a , \35324 , \21944 );
buf \U$27260 ( \35326 , \35325_nR23b8a );
not \U$27261 ( \35327 , \34916 );
and \U$27262 ( \35328 , RIe1bcce0_5826, \35327 );
not \U$27263 ( \35329 , RIe1bcce0_5826);
or \U$27264 ( \35330 , \35329 , \35223 );
not \U$27265 ( \35331 , \35313 );
and \U$27266 ( \35332 , \32914 , \35331 );
not \U$27267 ( \35333 , \35332 );
not \U$27268 ( \35334 , \35247 );
or \U$27269 ( \35335 , \34162 , \35334 );
nand \U$27270 ( \35336 , \35330 , \35333 , \35335 );
and \U$27271 ( \35337 , \35336 , \34916 );
or \U$27272 ( \35338 , \35328 , \35337 );
and \U$27274 ( \35339 , \35338 , 1'b1 );
or \U$27276 ( \35340 , \35339 , 1'b0 );
buf \U$27277 ( \35341 , \35340 );
_DC r23b0e_GF_IsGateDCbyConstraint ( \35342_nR23b0e , \35341 , \21944 );
buf \U$27278 ( \35343 , \35342_nR23b0e );
not \U$27279 ( \35344 , \32842 );
and \U$27280 ( \35345 , RIe1baf58_5827, \35344 );
not \U$27281 ( \35346 , RIe1baf58_5827);
or \U$27282 ( \35347 , \35346 , \35241 );
not \U$27283 ( \35348 , \35139 );
not \U$27284 ( \35349 , \35348 );
and \U$27285 ( \35350 , \32934 , \35349 );
not \U$27286 ( \35351 , \35350 );
nand \U$27287 ( \35352 , \32931 , \35155 );
nand \U$27288 ( \35353 , \35347 , \35351 , \35352 );
and \U$27289 ( \35354 , \35353 , \32842 );
or \U$27290 ( \35355 , \35345 , \35354 );
and \U$27292 ( \35356 , \35355 , 1'b1 );
or \U$27294 ( \35357 , \35356 , 1'b0 );
buf \U$27295 ( \35358 , \35357 );
_DC r23b10_GF_IsGateDCbyConstraint ( \35359_nR23b10 , \35358 , \21944 );
buf \U$27296 ( \35360 , \35359_nR23b10 );
not \U$27297 ( \35361 , \33296 );
and \U$27298 ( \35362 , RIe1b9158_5828, \35361 );
not \U$27299 ( \35363 , RIe1b9158_5828);
or \U$27300 ( \35364 , \35363 , \35169 );
not \U$27301 ( \35365 , \35139 );
not \U$27302 ( \35366 , \35365 );
and \U$27303 ( \35367 , \32953 , \35366 );
not \U$27304 ( \35368 , \35367 );
not \U$27305 ( \35369 , \35155 );
or \U$27306 ( \35370 , \34198 , \35369 );
nand \U$27307 ( \35371 , \35364 , \35368 , \35370 );
and \U$27308 ( \35372 , \35371 , \33296 );
or \U$27309 ( \35373 , \35362 , \35372 );
and \U$27311 ( \35374 , \35373 , 1'b1 );
or \U$27313 ( \35375 , \35374 , 1'b0 );
buf \U$27314 ( \35376 , \35375 );
_DC r23b12_GF_IsGateDCbyConstraint ( \35377_nR23b12 , \35376 , \21944 );
buf \U$27315 ( \35378 , \35377_nR23b12 );
not \U$27316 ( \35379 , \34916 );
and \U$27317 ( \35380 , RIe1b6908_5829, \35379 );
not \U$27318 ( \35381 , RIe1b6908_5829);
or \U$27319 ( \35382 , \35381 , \35311 );
not \U$27320 ( \35383 , \35150 );
and \U$27321 ( \35384 , \32973 , \35383 );
not \U$27322 ( \35385 , \35384 );
not \U$27323 ( \35386 , \35155 );
or \U$27324 ( \35387 , \34216 , \35386 );
nand \U$27325 ( \35388 , \35382 , \35385 , \35387 );
and \U$27326 ( \35389 , \35388 , \34916 );
or \U$27327 ( \35390 , \35380 , \35389 );
and \U$27329 ( \35391 , \35390 , 1'b1 );
or \U$27331 ( \35392 , \35391 , 1'b0 );
buf \U$27332 ( \35393 , \35392 );
_DC r23b14_GF_IsGateDCbyConstraint ( \35394_nR23b14 , \35393 , \21944 );
buf \U$27333 ( \35395 , \35394_nR23b14 );
not \U$27334 ( \35396 , \32842 );
and \U$27335 ( \35397 , RIe1b3b90_5830, \35396 );
not \U$27336 ( \35398 , RIe1b3b90_5830);
or \U$27337 ( \35399 , \35398 , \35311 );
not \U$27338 ( \35400 , \35313 );
and \U$27339 ( \35401 , \32994 , \35400 );
not \U$27340 ( \35402 , \35401 );
not \U$27341 ( \35403 , \35247 );
or \U$27342 ( \35404 , \34234 , \35403 );
nand \U$27343 ( \35405 , \35399 , \35402 , \35404 );
and \U$27344 ( \35406 , \35405 , \32842 );
or \U$27345 ( \35407 , \35397 , \35406 );
and \U$27347 ( \35408 , \35407 , 1'b1 );
or \U$27349 ( \35409 , \35408 , 1'b0 );
buf \U$27350 ( \35410 , \35409 );
_DC r23b16_GF_IsGateDCbyConstraint ( \35411_nR23b16 , \35410 , \21944 );
buf \U$27351 ( \35412 , \35411_nR23b16 );
not \U$27352 ( \35413 , \34661 );
and \U$27353 ( \35414 , RIe1b1d18_5831, \35413 );
not \U$27354 ( \35415 , RIe1b1d18_5831);
or \U$27355 ( \35416 , \35415 , \35311 );
not \U$27356 ( \35417 , \35348 );
and \U$27357 ( \35418 , \33014 , \35417 );
not \U$27358 ( \35419 , \35418 );
not \U$27359 ( \35420 , \35209 );
or \U$27360 ( \35421 , \34252 , \35420 );
nand \U$27361 ( \35422 , \35416 , \35419 , \35421 );
and \U$27362 ( \35423 , \35422 , \34661 );
or \U$27363 ( \35424 , \35414 , \35423 );
and \U$27365 ( \35425 , \35424 , 1'b1 );
or \U$27367 ( \35426 , \35425 , 1'b0 );
buf \U$27368 ( \35427 , \35426 );
_DC r23b18_GF_IsGateDCbyConstraint ( \35428_nR23b18 , \35427 , \21944 );
buf \U$27369 ( \35429 , \35428_nR23b18 );
not \U$27370 ( \35430 , \34916 );
and \U$27371 ( \35431 , RIe1aff90_5832, \35430 );
not \U$27372 ( \35432 , RIe1aff90_5832);
or \U$27373 ( \35433 , \35432 , \35147 );
not \U$27374 ( \35434 , \35365 );
and \U$27375 ( \35435 , \33033 , \35434 );
not \U$27376 ( \35436 , \35435 );
not \U$27377 ( \35437 , \35247 );
or \U$27378 ( \35438 , \34270 , \35437 );
nand \U$27379 ( \35439 , \35433 , \35436 , \35438 );
and \U$27380 ( \35440 , \35439 , \34916 );
or \U$27381 ( \35441 , \35431 , \35440 );
and \U$27383 ( \35442 , \35441 , 1'b1 );
or \U$27385 ( \35443 , \35442 , 1'b0 );
buf \U$27386 ( \35444 , \35443 );
_DC r23b1a_GF_IsGateDCbyConstraint ( \35445_nR23b1a , \35444 , \21944 );
buf \U$27387 ( \35446 , \35445_nR23b1a );
not \U$27388 ( \35447 , \32842 );
and \U$27389 ( \35448 , RIe1ae2f8_5833, \35447 );
not \U$27390 ( \35449 , RIe1ae2f8_5833);
or \U$27391 ( \35450 , \35449 , \35169 );
not \U$27392 ( \35451 , \35188 );
and \U$27393 ( \35452 , \33052 , \35451 );
not \U$27394 ( \35453 , \35452 );
not \U$27395 ( \35454 , \35154 );
or \U$27396 ( \35455 , \34288 , \35454 );
nand \U$27397 ( \35456 , \35450 , \35453 , \35455 );
and \U$27398 ( \35457 , \35456 , \32842 );
or \U$27399 ( \35458 , \35448 , \35457 );
and \U$27401 ( \35459 , \35458 , 1'b1 );
or \U$27403 ( \35460 , \35459 , 1'b0 );
buf \U$27404 ( \35461 , \35460 );
_DC r23b1c_GF_IsGateDCbyConstraint ( \35462_nR23b1c , \35461 , \21944 );
buf \U$27405 ( \35463 , \35462_nR23b1c );
not \U$27406 ( \35464 , \33217 );
and \U$27407 ( \35465 , RIe1ab940_5834, \35464 );
not \U$27408 ( \35466 , RIe1ab940_5834);
or \U$27409 ( \35467 , \35466 , \35147 );
not \U$27410 ( \35468 , \35188 );
and \U$27411 ( \35469 , \33071 , \35468 );
not \U$27412 ( \35470 , \35469 );
not \U$27413 ( \35471 , \35209 );
or \U$27414 ( \35472 , \34307 , \35471 );
nand \U$27415 ( \35473 , \35467 , \35470 , \35472 );
and \U$27416 ( \35474 , \35473 , \33217 );
or \U$27417 ( \35475 , \35465 , \35474 );
and \U$27419 ( \35476 , \35475 , 1'b1 );
or \U$27421 ( \35477 , \35476 , 1'b0 );
buf \U$27422 ( \35478 , \35477 );
_DC r23b1e_GF_IsGateDCbyConstraint ( \35479_nR23b1e , \35478 , \21944 );
buf \U$27423 ( \35480 , \35479_nR23b1e );
not \U$27424 ( \35481 , \34916 );
and \U$27425 ( \35482 , RIe1a8628_5835, \35481 );
not \U$27426 ( \35483 , RIe1a8628_5835);
or \U$27427 ( \35484 , \35483 , \35241 );
not \U$27428 ( \35485 , \35188 );
and \U$27429 ( \35486 , \33091 , \35485 );
not \U$27430 ( \35487 , \35486 );
not \U$27431 ( \35488 , \35155 );
or \U$27432 ( \35489 , \34326 , \35488 );
nand \U$27433 ( \35490 , \35484 , \35487 , \35489 );
and \U$27434 ( \35491 , \35490 , \34916 );
or \U$27435 ( \35492 , \35482 , \35491 );
and \U$27437 ( \35493 , \35492 , 1'b1 );
or \U$27439 ( \35494 , \35493 , 1'b0 );
buf \U$27440 ( \35495 , \35494 );
_DC r23b20_GF_IsGateDCbyConstraint ( \35496_nR23b20 , \35495 , \21944 );
buf \U$27441 ( \35497 , \35496_nR23b20 );
not \U$27442 ( \35498 , \32842 );
and \U$27443 ( \35499 , RIe1a6030_5836, \35498 );
not \U$27444 ( \35500 , RIe1a6030_5836);
or \U$27445 ( \35501 , \35500 , \35311 );
not \U$27446 ( \35502 , \35243 );
and \U$27447 ( \35503 , \33110 , \35502 );
not \U$27448 ( \35504 , \35503 );
not \U$27449 ( \35505 , \35154 );
or \U$27450 ( \35506 , \34344 , \35505 );
nand \U$27451 ( \35507 , \35501 , \35504 , \35506 );
and \U$27452 ( \35508 , \35507 , \32842 );
or \U$27453 ( \35509 , \35499 , \35508 );
and \U$27455 ( \35510 , \35509 , 1'b1 );
or \U$27457 ( \35511 , \35510 , 1'b0 );
buf \U$27458 ( \35512 , \35511 );
_DC r23b24_GF_IsGateDCbyConstraint ( \35513_nR23b24 , \35512 , \21944 );
buf \U$27459 ( \35514 , \35513_nR23b24 );
not \U$27460 ( \35515 , \34661 );
and \U$27461 ( \35516 , RIe1a2d90_5837, \35515 );
not \U$27462 ( \35517 , RIe1a2d90_5837);
or \U$27463 ( \35518 , \35517 , \35241 );
not \U$27464 ( \35519 , \35313 );
and \U$27465 ( \35520 , \33129 , \35519 );
not \U$27466 ( \35521 , \35520 );
not \U$27467 ( \35522 , \35154 );
or \U$27468 ( \35523 , \34362 , \35522 );
nand \U$27469 ( \35524 , \35518 , \35521 , \35523 );
and \U$27470 ( \35525 , \35524 , \34661 );
or \U$27471 ( \35526 , \35516 , \35525 );
and \U$27473 ( \35527 , \35526 , 1'b1 );
or \U$27475 ( \35528 , \35527 , 1'b0 );
buf \U$27476 ( \35529 , \35528 );
_DC r23b26_GF_IsGateDCbyConstraint ( \35530_nR23b26 , \35529 , \21944 );
buf \U$27477 ( \35531 , \35530_nR23b26 );
buf \U$27478 ( \35532 , \34915 );
not \U$27479 ( \35533 , \35532 );
and \U$27480 ( \35534 , RIe1a0540_5838, \35533 );
not \U$27481 ( \35535 , RIe1a0540_5838);
or \U$27482 ( \35536 , \35535 , \35223 );
not \U$27483 ( \35537 , \35150 );
and \U$27484 ( \35538 , \33149 , \35537 );
not \U$27485 ( \35539 , \35538 );
not \U$27486 ( \35540 , \35155 );
or \U$27487 ( \35541 , \34380 , \35540 );
nand \U$27488 ( \35542 , \35536 , \35539 , \35541 );
and \U$27489 ( \35543 , \35542 , \35532 );
or \U$27490 ( \35544 , \35534 , \35543 );
and \U$27492 ( \35545 , \35544 , 1'b1 );
or \U$27494 ( \35546 , \35545 , 1'b0 );
buf \U$27495 ( \35547 , \35546 );
_DC r23b28_GF_IsGateDCbyConstraint ( \35548_nR23b28 , \35547 , \21944 );
buf \U$27496 ( \35549 , \35548_nR23b28 );
not \U$27497 ( \35550 , \32842 );
and \U$27498 ( \35551 , RIe19da20_5839, \35550 );
not \U$27499 ( \35552 , RIe19da20_5839);
or \U$27500 ( \35553 , \35552 , \35223 );
not \U$27501 ( \35554 , \35243 );
and \U$27502 ( \35555 , \33167 , \35554 );
not \U$27503 ( \35556 , \35555 );
not \U$27504 ( \35557 , \35154 );
or \U$27505 ( \35558 , \34398 , \35557 );
nand \U$27506 ( \35559 , \35553 , \35556 , \35558 );
and \U$27507 ( \35560 , \35559 , \32842 );
or \U$27508 ( \35561 , \35551 , \35560 );
and \U$27510 ( \35562 , \35561 , 1'b1 );
or \U$27512 ( \35563 , \35562 , 1'b0 );
buf \U$27513 ( \35564 , \35563 );
_DC r23b2a_GF_IsGateDCbyConstraint ( \35565_nR23b2a , \35564 , \21944 );
buf \U$27514 ( \35566 , \35565_nR23b2a );
not \U$27515 ( \35567 , \33336 );
and \U$27516 ( \35568 , RIe19a870_5840, \35567 );
not \U$27517 ( \35569 , RIe19a870_5840);
or \U$27518 ( \35570 , \35569 , \35147 );
not \U$27519 ( \35571 , \35313 );
and \U$27520 ( \35572 , \33187 , \35571 );
not \U$27521 ( \35573 , \35572 );
not \U$27522 ( \35574 , \35154 );
or \U$27523 ( \35575 , \34416 , \35574 );
nand \U$27524 ( \35576 , \35570 , \35573 , \35575 );
and \U$27525 ( \35577 , \35576 , \33336 );
or \U$27526 ( \35578 , \35568 , \35577 );
and \U$27528 ( \35579 , \35578 , 1'b1 );
or \U$27530 ( \35580 , \35579 , 1'b0 );
buf \U$27531 ( \35581 , \35580 );
_DC r23b2c_GF_IsGateDCbyConstraint ( \35582_nR23b2c , \35581 , \21944 );
buf \U$27532 ( \35583 , \35582_nR23b2c );
not \U$27533 ( \35584 , \35532 );
and \U$27534 ( \35585 , RIe197cd8_5841, \35584 );
not \U$27535 ( \35586 , RIe197cd8_5841);
or \U$27536 ( \35587 , \35586 , \35223 );
not \U$27537 ( \35588 , \35365 );
and \U$27538 ( \35589 , \33205 , \35588 );
not \U$27539 ( \35590 , \35589 );
not \U$27540 ( \35591 , \35155 );
or \U$27541 ( \35592 , \34434 , \35591 );
nand \U$27542 ( \35593 , \35587 , \35590 , \35592 );
and \U$27543 ( \35594 , \35593 , \35532 );
or \U$27544 ( \35595 , \35585 , \35594 );
and \U$27546 ( \35596 , \35595 , 1'b1 );
or \U$27548 ( \35597 , \35596 , 1'b0 );
buf \U$27549 ( \35598 , \35597 );
_DC r23b2e_GF_IsGateDCbyConstraint ( \35599_nR23b2e , \35598 , \21944 );
buf \U$27550 ( \35600 , \35599_nR23b2e );
not \U$27551 ( \35601 , \32842 );
and \U$27552 ( \35602 , RIe195410_5842, \35601 );
not \U$27553 ( \35603 , RIe195410_5842);
or \U$27554 ( \35604 , \35603 , \35147 );
not \U$27555 ( \35605 , \35313 );
and \U$27556 ( \35606 , \33226 , \35605 );
not \U$27557 ( \35607 , \35606 );
not \U$27558 ( \35608 , \35154 );
or \U$27559 ( \35609 , \34452 , \35608 );
nand \U$27560 ( \35610 , \35604 , \35607 , \35609 );
and \U$27561 ( \35611 , \35610 , \32842 );
or \U$27562 ( \35612 , \35602 , \35611 );
and \U$27564 ( \35613 , \35612 , 1'b1 );
or \U$27566 ( \35614 , \35613 , 1'b0 );
buf \U$27567 ( \35615 , \35614 );
_DC r23b30_GF_IsGateDCbyConstraint ( \35616_nR23b30 , \35615 , \21944 );
buf \U$27568 ( \35617 , \35616_nR23b30 );
not \U$27569 ( \35618 , \33218 );
and \U$27570 ( \35619 , RIe192e90_5843, \35618 );
not \U$27571 ( \35620 , RIe192e90_5843);
or \U$27572 ( \35621 , \35620 , \35241 );
not \U$27573 ( \35622 , \35150 );
and \U$27574 ( \35623 , \33245 , \35622 );
not \U$27575 ( \35624 , \35623 );
not \U$27576 ( \35625 , \35209 );
or \U$27577 ( \35626 , \34470 , \35625 );
nand \U$27578 ( \35627 , \35621 , \35624 , \35626 );
and \U$27579 ( \35628 , \35627 , \33218 );
or \U$27580 ( \35629 , \35619 , \35628 );
and \U$27582 ( \35630 , \35629 , 1'b1 );
or \U$27584 ( \35631 , \35630 , 1'b0 );
buf \U$27585 ( \35632 , \35631 );
_DC r23b32_GF_IsGateDCbyConstraint ( \35633_nR23b32 , \35632 , \21944 );
buf \U$27586 ( \35634 , \35633_nR23b32 );
not \U$27587 ( \35635 , \35532 );
and \U$27588 ( \35636 , RIe190460_5844, \35635 );
not \U$27589 ( \35637 , RIe190460_5844);
or \U$27590 ( \35638 , \35637 , \35311 );
not \U$27591 ( \35639 , \35365 );
and \U$27592 ( \35640 , \33265 , \35639 );
not \U$27593 ( \35641 , \35640 );
not \U$27594 ( \35642 , \35155 );
or \U$27595 ( \35643 , \34488 , \35642 );
nand \U$27596 ( \35644 , \35638 , \35641 , \35643 );
and \U$27597 ( \35645 , \35644 , \35532 );
or \U$27598 ( \35646 , \35636 , \35645 );
and \U$27600 ( \35647 , \35646 , 1'b1 );
or \U$27602 ( \35648 , \35647 , 1'b0 );
buf \U$27603 ( \35649 , \35648 );
_DC r23b34_GF_IsGateDCbyConstraint ( \35650_nR23b34 , \35649 , \21944 );
buf \U$27604 ( \35651 , \35650_nR23b34 );
not \U$27605 ( \35652 , \32842 );
and \U$27606 ( \35653 , RIe18e0c0_5845, \35652 );
not \U$27607 ( \35654 , RIe18e0c0_5845);
or \U$27608 ( \35655 , \35654 , \35147 );
not \U$27609 ( \35656 , \35150 );
and \U$27610 ( \35657 , \33284 , \35656 );
not \U$27611 ( \35658 , \35657 );
not \U$27612 ( \35659 , \35155 );
or \U$27613 ( \35660 , \34506 , \35659 );
nand \U$27614 ( \35661 , \35655 , \35658 , \35660 );
and \U$27615 ( \35662 , \35661 , \32842 );
or \U$27616 ( \35663 , \35653 , \35662 );
and \U$27618 ( \35664 , \35663 , 1'b1 );
or \U$27620 ( \35665 , \35664 , 1'b0 );
buf \U$27621 ( \35666 , \35665 );
_DC r23b36_GF_IsGateDCbyConstraint ( \35667_nR23b36 , \35666 , \21944 );
buf \U$27622 ( \35668 , \35667_nR23b36 );
not \U$27623 ( \35669 , \32755 );
and \U$27624 ( \35670 , RIe18bc30_5846, \35669 );
not \U$27625 ( \35671 , RIe18bc30_5846);
or \U$27626 ( \35672 , \35671 , \35311 );
not \U$27627 ( \35673 , \35313 );
and \U$27628 ( \35674 , \33305 , \35673 );
not \U$27629 ( \35675 , \35674 );
not \U$27630 ( \35676 , \35247 );
or \U$27631 ( \35677 , \34524 , \35676 );
nand \U$27632 ( \35678 , \35672 , \35675 , \35677 );
and \U$27633 ( \35679 , \35678 , \32755 );
or \U$27634 ( \35680 , \35670 , \35679 );
and \U$27636 ( \35681 , \35680 , 1'b1 );
or \U$27638 ( \35682 , \35681 , 1'b0 );
buf \U$27639 ( \35683 , \35682 );
_DC r23b3a_GF_IsGateDCbyConstraint ( \35684_nR23b3a , \35683 , \21944 );
buf \U$27640 ( \35685 , \35684_nR23b3a );
not \U$27641 ( \35686 , \35532 );
and \U$27642 ( \35687 , RIe189098_5847, \35686 );
not \U$27643 ( \35688 , RIe189098_5847);
or \U$27644 ( \35689 , \35688 , \35147 );
not \U$27645 ( \35690 , \35150 );
and \U$27646 ( \35691 , \33324 , \35690 );
not \U$27647 ( \35692 , \35691 );
not \U$27648 ( \35693 , \35154 );
or \U$27649 ( \35694 , \34542 , \35693 );
nand \U$27650 ( \35695 , \35689 , \35692 , \35694 );
and \U$27651 ( \35696 , \35695 , \35532 );
or \U$27652 ( \35697 , \35687 , \35696 );
and \U$27654 ( \35698 , \35697 , 1'b1 );
or \U$27656 ( \35699 , \35698 , 1'b0 );
buf \U$27657 ( \35700 , \35699 );
_DC r23b3c_GF_IsGateDCbyConstraint ( \35701_nR23b3c , \35700 , \21944 );
buf \U$27658 ( \35702 , \35701_nR23b3c );
not \U$27659 ( \35703 , \32842 );
and \U$27660 ( \35704 , RIe186c08_5848, \35703 );
not \U$27661 ( \35705 , RIe186c08_5848);
or \U$27662 ( \35706 , \35705 , \35223 );
not \U$27663 ( \35707 , \35313 );
and \U$27664 ( \35708 , \33344 , \35707 );
not \U$27665 ( \35709 , \35708 );
not \U$27666 ( \35710 , \35155 );
or \U$27667 ( \35711 , \34560 , \35710 );
nand \U$27668 ( \35712 , \35706 , \35709 , \35711 );
and \U$27669 ( \35713 , \35712 , \32842 );
or \U$27670 ( \35714 , \35704 , \35713 );
and \U$27672 ( \35715 , \35714 , 1'b1 );
or \U$27674 ( \35716 , \35715 , 1'b0 );
buf \U$27675 ( \35717 , \35716 );
_DC r23b3e_GF_IsGateDCbyConstraint ( \35718_nR23b3e , \35717 , \21944 );
buf \U$27676 ( \35719 , \35718_nR23b3e );
not \U$27677 ( \35720 , \34661 );
and \U$27678 ( \35721 , RIe1839e0_5849, \35720 );
not \U$27679 ( \35722 , RIe1839e0_5849);
or \U$27680 ( \35723 , \35722 , \35241 );
not \U$27681 ( \35724 , \35348 );
and \U$27682 ( \35725 , \33363 , \35724 );
not \U$27683 ( \35726 , \35725 );
not \U$27684 ( \35727 , \35154 );
or \U$27685 ( \35728 , \34578 , \35727 );
nand \U$27686 ( \35729 , \35723 , \35726 , \35728 );
and \U$27687 ( \35730 , \35729 , \34661 );
or \U$27688 ( \35731 , \35721 , \35730 );
and \U$27690 ( \35732 , \35731 , 1'b1 );
or \U$27692 ( \35733 , \35732 , 1'b0 );
buf \U$27693 ( \35734 , \35733 );
_DC r23b40_GF_IsGateDCbyConstraint ( \35735_nR23b40 , \35734 , \21944 );
buf \U$27694 ( \35736 , \35735_nR23b40 );
not \U$27695 ( \35737 , \35532 );
and \U$27696 ( \35738 , RIe1817a8_5850, \35737 );
not \U$27697 ( \35739 , RIe1817a8_5850);
or \U$27698 ( \35740 , \35739 , \35241 );
not \U$27699 ( \35741 , \35365 );
and \U$27700 ( \35742 , \33382 , \35741 );
not \U$27701 ( \35743 , \35742 );
not \U$27702 ( \35744 , \35155 );
or \U$27703 ( \35745 , \34596 , \35744 );
nand \U$27704 ( \35746 , \35740 , \35743 , \35745 );
and \U$27705 ( \35747 , \35746 , \35532 );
or \U$27706 ( \35748 , \35738 , \35747 );
and \U$27708 ( \35749 , \35748 , 1'b1 );
or \U$27710 ( \35750 , \35749 , 1'b0 );
buf \U$27711 ( \35751 , \35750 );
_DC r23b42_GF_IsGateDCbyConstraint ( \35752_nR23b42 , \35751 , \21944 );
buf \U$27712 ( \35753 , \35752_nR23b42 );
not \U$27713 ( \35754 , \32842 );
and \U$27714 ( \35755 , RIe17fb88_5851, \35754 );
not \U$27715 ( \35756 , RIe17fb88_5851);
or \U$27716 ( \35757 , \35756 , \35169 );
not \U$27717 ( \35758 , \35188 );
and \U$27718 ( \35759 , \33402 , \35758 );
not \U$27719 ( \35760 , \35759 );
not \U$27720 ( \35761 , \35155 );
or \U$27721 ( \35762 , \34614 , \35761 );
nand \U$27722 ( \35763 , \35757 , \35760 , \35762 );
and \U$27723 ( \35764 , \35763 , \32842 );
or \U$27724 ( \35765 , \35755 , \35764 );
and \U$27726 ( \35766 , \35765 , 1'b1 );
or \U$27728 ( \35767 , \35766 , 1'b0 );
buf \U$27729 ( \35768 , \35767 );
_DC r23b44_GF_IsGateDCbyConstraint ( \35769_nR23b44 , \35768 , \21944 );
buf \U$27730 ( \35770 , \35769_nR23b44 );
not \U$27731 ( \35771 , \32864 );
and \U$27732 ( \35772 , RIe17def0_5852, \35771 );
not \U$27733 ( \35773 , RIe17def0_5852);
or \U$27734 ( \35774 , \35773 , \35169 );
not \U$27735 ( \35775 , \35150 );
and \U$27736 ( \35776 , \33422 , \35775 );
not \U$27737 ( \35777 , \35776 );
not \U$27738 ( \35778 , \35154 );
or \U$27739 ( \35779 , \34632 , \35778 );
nand \U$27740 ( \35780 , \35774 , \35777 , \35779 );
and \U$27741 ( \35781 , \35780 , \32864 );
or \U$27742 ( \35782 , \35772 , \35781 );
and \U$27744 ( \35783 , \35782 , 1'b1 );
or \U$27746 ( \35784 , \35783 , 1'b0 );
buf \U$27747 ( \35785 , \35784 );
_DC r23b46_GF_IsGateDCbyConstraint ( \35786_nR23b46 , \35785 , \21944 );
buf \U$27748 ( \35787 , \35786_nR23b46 );
not \U$27749 ( \35788 , \35532 );
and \U$27750 ( \35789 , RIe17c3c0_5853, \35788 );
not \U$27751 ( \35790 , RIe17c3c0_5853);
or \U$27752 ( \35791 , \35790 , \35241 );
not \U$27753 ( \35792 , \35348 );
and \U$27754 ( \35793 , \33440 , \35792 );
not \U$27755 ( \35794 , \35793 );
not \U$27756 ( \35795 , \35154 );
or \U$27757 ( \35796 , \34650 , \35795 );
nand \U$27758 ( \35797 , \35791 , \35794 , \35796 );
and \U$27759 ( \35798 , \35797 , \35532 );
or \U$27760 ( \35799 , \35789 , \35798 );
and \U$27762 ( \35800 , \35799 , 1'b1 );
or \U$27764 ( \35801 , \35800 , 1'b0 );
buf \U$27765 ( \35802 , \35801 );
_DC r23b48_GF_IsGateDCbyConstraint ( \35803_nR23b48 , \35802 , \21944 );
buf \U$27766 ( \35804 , \35803_nR23b48 );
not \U$27767 ( \35805 , \32842 );
and \U$27768 ( \35806 , RIe17a458_5854, \35805 );
not \U$27769 ( \35807 , RIe17a458_5854);
or \U$27770 ( \35808 , \35807 , \35223 );
not \U$27771 ( \35809 , \35365 );
and \U$27772 ( \35810 , \33459 , \35809 );
not \U$27773 ( \35811 , \35810 );
not \U$27774 ( \35812 , \35155 );
or \U$27775 ( \35813 , \34669 , \35812 );
nand \U$27776 ( \35814 , \35808 , \35811 , \35813 );
and \U$27777 ( \35815 , \35814 , \32842 );
or \U$27778 ( \35816 , \35806 , \35815 );
and \U$27780 ( \35817 , \35816 , 1'b1 );
or \U$27782 ( \35818 , \35817 , 1'b0 );
buf \U$27783 ( \35819 , \35818 );
_DC r23b4a_GF_IsGateDCbyConstraint ( \35820_nR23b4a , \35819 , \21944 );
buf \U$27784 ( \35821 , \35820_nR23b4a );
not \U$27785 ( \35822 , \33217 );
and \U$27786 ( \35823 , RIe1781a8_5855, \35822 );
not \U$27787 ( \35824 , RIe1781a8_5855);
or \U$27788 ( \35825 , \35824 , \35311 );
not \U$27789 ( \35826 , \35188 );
and \U$27790 ( \35827 , \33478 , \35826 );
not \U$27791 ( \35828 , \35827 );
not \U$27792 ( \35829 , \35155 );
or \U$27793 ( \35830 , \34687 , \35829 );
nand \U$27794 ( \35831 , \35825 , \35828 , \35830 );
and \U$27795 ( \35832 , \35831 , \33217 );
or \U$27796 ( \35833 , \35823 , \35832 );
and \U$27798 ( \35834 , \35833 , 1'b1 );
or \U$27800 ( \35835 , \35834 , 1'b0 );
buf \U$27801 ( \35836 , \35835 );
_DC r23b4c_GF_IsGateDCbyConstraint ( \35837_nR23b4c , \35836 , \21944 );
buf \U$27802 ( \35838 , \35837_nR23b4c );
not \U$27803 ( \35839 , \35532 );
and \U$27804 ( \35840 , RIe176240_5856, \35839 );
not \U$27805 ( \35841 , RIe176240_5856);
or \U$27806 ( \35842 , \35841 , \35311 );
not \U$27807 ( \35843 , \35150 );
and \U$27808 ( \35844 , \33497 , \35843 );
not \U$27809 ( \35845 , \35844 );
not \U$27810 ( \35846 , \35155 );
or \U$27811 ( \35847 , \34706 , \35846 );
nand \U$27812 ( \35848 , \35842 , \35845 , \35847 );
and \U$27813 ( \35849 , \35848 , \35532 );
or \U$27814 ( \35850 , \35840 , \35849 );
and \U$27816 ( \35851 , \35850 , 1'b1 );
or \U$27818 ( \35852 , \35851 , 1'b0 );
buf \U$27819 ( \35853 , \35852 );
_DC r23b50_GF_IsGateDCbyConstraint ( \35854_nR23b50 , \35853 , \21944 );
buf \U$27820 ( \35855 , \35854_nR23b50 );
not \U$27821 ( \35856 , \32842 );
and \U$27822 ( \35857 , RIe174530_5857, \35856 );
not \U$27823 ( \35858 , RIe174530_5857);
or \U$27824 ( \35859 , \35858 , \35223 );
not \U$27825 ( \35860 , \35243 );
and \U$27826 ( \35861 , \33517 , \35860 );
not \U$27827 ( \35862 , \35861 );
not \U$27828 ( \35863 , \35247 );
or \U$27829 ( \35864 , \34724 , \35863 );
nand \U$27830 ( \35865 , \35859 , \35862 , \35864 );
and \U$27831 ( \35866 , \35865 , \32842 );
or \U$27832 ( \35867 , \35857 , \35866 );
and \U$27834 ( \35868 , \35867 , 1'b1 );
or \U$27836 ( \35869 , \35868 , 1'b0 );
buf \U$27837 ( \35870 , \35869 );
_DC r23b52_GF_IsGateDCbyConstraint ( \35871_nR23b52 , \35870 , \21944 );
buf \U$27838 ( \35872 , \35871_nR23b52 );
not \U$27839 ( \35873 , \32864 );
and \U$27840 ( \35874 , RIe172988_5858, \35873 );
not \U$27841 ( \35875 , RIe172988_5858);
or \U$27842 ( \35876 , \35875 , \35169 );
not \U$27843 ( \35877 , \35313 );
and \U$27844 ( \35878 , \33537 , \35877 );
not \U$27845 ( \35879 , \35878 );
not \U$27846 ( \35880 , \35209 );
or \U$27847 ( \35881 , \34742 , \35880 );
nand \U$27848 ( \35882 , \35876 , \35879 , \35881 );
and \U$27849 ( \35883 , \35882 , \32864 );
or \U$27850 ( \35884 , \35874 , \35883 );
and \U$27852 ( \35885 , \35884 , 1'b1 );
or \U$27854 ( \35886 , \35885 , 1'b0 );
buf \U$27855 ( \35887 , \35886 );
_DC r23b54_GF_IsGateDCbyConstraint ( \35888_nR23b54 , \35887 , \21944 );
buf \U$27856 ( \35889 , \35888_nR23b54 );
not \U$27857 ( \35890 , \35532 );
and \U$27858 ( \35891 , RIe16fc70_5859, \35890 );
not \U$27859 ( \35892 , RIe16fc70_5859);
or \U$27860 ( \35893 , \35892 , \35311 );
not \U$27861 ( \35894 , \35348 );
and \U$27862 ( \35895 , \33556 , \35894 );
not \U$27863 ( \35896 , \35895 );
not \U$27864 ( \35897 , \35247 );
or \U$27865 ( \35898 , \34760 , \35897 );
nand \U$27866 ( \35899 , \35893 , \35896 , \35898 );
and \U$27867 ( \35900 , \35899 , \35532 );
or \U$27868 ( \35901 , \35891 , \35900 );
and \U$27870 ( \35902 , \35901 , 1'b1 );
or \U$27872 ( \35903 , \35902 , 1'b0 );
buf \U$27873 ( \35904 , \35903 );
_DC r23b56_GF_IsGateDCbyConstraint ( \35905_nR23b56 , \35904 , \21944 );
buf \U$27874 ( \35906 , \35905_nR23b56 );
not \U$27875 ( \35907 , \32842 );
and \U$27876 ( \35908 , RIe16e140_5860, \35907 );
not \U$27877 ( \35909 , RIe16e140_5860);
or \U$27878 ( \35910 , \35909 , \35223 );
not \U$27879 ( \35911 , \35243 );
and \U$27880 ( \35912 , \33576 , \35911 );
not \U$27881 ( \35913 , \35912 );
not \U$27882 ( \35914 , \35154 );
or \U$27883 ( \35915 , \34778 , \35914 );
nand \U$27884 ( \35916 , \35910 , \35913 , \35915 );
and \U$27885 ( \35917 , \35916 , \32842 );
or \U$27886 ( \35918 , \35908 , \35917 );
and \U$27888 ( \35919 , \35918 , 1'b1 );
or \U$27890 ( \35920 , \35919 , 1'b0 );
buf \U$27891 ( \35921 , \35920 );
_DC r23b58_GF_IsGateDCbyConstraint ( \35922_nR23b58 , \35921 , \21944 );
buf \U$27892 ( \35923 , \35922_nR23b58 );
not \U$27893 ( \35924 , \33218 );
and \U$27894 ( \35925 , RIe16c1d8_5861, \35924 );
not \U$27895 ( \35926 , RIe16c1d8_5861);
or \U$27896 ( \35927 , \35926 , \35147 );
not \U$27897 ( \35928 , \35313 );
and \U$27898 ( \35929 , \33594 , \35928 );
not \U$27899 ( \35930 , \35929 );
not \U$27900 ( \35931 , \35247 );
or \U$27901 ( \35932 , \34796 , \35931 );
nand \U$27902 ( \35933 , \35927 , \35930 , \35932 );
and \U$27903 ( \35934 , \35933 , \33218 );
or \U$27904 ( \35935 , \35925 , \35934 );
and \U$27906 ( \35936 , \35935 , 1'b1 );
or \U$27908 ( \35937 , \35936 , 1'b0 );
buf \U$27909 ( \35938 , \35937 );
_DC r23b5a_GF_IsGateDCbyConstraint ( \35939_nR23b5a , \35938 , \21944 );
buf \U$27910 ( \35940 , \35939_nR23b5a );
not \U$27911 ( \35941 , \35532 );
and \U$27912 ( \35942 , RIe16a5b8_5862, \35941 );
not \U$27913 ( \35943 , RIe16a5b8_5862);
or \U$27914 ( \35944 , \35943 , \35223 );
not \U$27915 ( \35945 , \35243 );
and \U$27916 ( \35946 , \33612 , \35945 );
not \U$27917 ( \35947 , \35946 );
not \U$27918 ( \35948 , \35155 );
or \U$27919 ( \35949 , \34814 , \35948 );
nand \U$27920 ( \35950 , \35944 , \35947 , \35949 );
and \U$27921 ( \35951 , \35950 , \35532 );
or \U$27922 ( \35952 , \35942 , \35951 );
and \U$27924 ( \35953 , \35952 , 1'b1 );
or \U$27926 ( \35954 , \35953 , 1'b0 );
buf \U$27927 ( \35955 , \35954 );
_DC r23b5c_GF_IsGateDCbyConstraint ( \35956_nR23b5c , \35955 , \21944 );
buf \U$27928 ( \35957 , \35956_nR23b5c );
not \U$27929 ( \35958 , \34915 );
and \U$27930 ( \35959 , RIe168a88_5863, \35958 );
not \U$27931 ( \35960 , RIe168a88_5863);
or \U$27932 ( \35961 , \35960 , \35241 );
not \U$27933 ( \35962 , \35313 );
and \U$27934 ( \35963 , \33632 , \35962 );
not \U$27935 ( \35964 , \35963 );
not \U$27936 ( \35965 , \35247 );
or \U$27937 ( \35966 , \34832 , \35965 );
nand \U$27938 ( \35967 , \35961 , \35964 , \35966 );
and \U$27939 ( \35968 , \35967 , \34915 );
or \U$27940 ( \35969 , \35959 , \35968 );
and \U$27942 ( \35970 , \35969 , 1'b1 );
or \U$27944 ( \35971 , \35970 , 1'b0 );
buf \U$27945 ( \35972 , \35971 );
_DC r23b5e_GF_IsGateDCbyConstraint ( \35973_nR23b5e , \35972 , \21944 );
buf \U$27946 ( \35974 , \35973_nR23b5e );
not \U$27947 ( \35975 , \33218 );
and \U$27948 ( \35976 , RIe167138_5864, \35975 );
not \U$27949 ( \35977 , RIe167138_5864);
or \U$27950 ( \35978 , \35977 , \35147 );
not \U$27951 ( \35979 , \35313 );
and \U$27952 ( \35980 , \33651 , \35979 );
not \U$27953 ( \35981 , \35980 );
not \U$27954 ( \35982 , \35209 );
or \U$27955 ( \35983 , \34850 , \35982 );
nand \U$27956 ( \35984 , \35978 , \35981 , \35983 );
and \U$27957 ( \35985 , \35984 , \33218 );
or \U$27958 ( \35986 , \35976 , \35985 );
and \U$27960 ( \35987 , \35986 , 1'b1 );
or \U$27962 ( \35988 , \35987 , 1'b0 );
buf \U$27963 ( \35989 , \35988 );
_DC r23b60_GF_IsGateDCbyConstraint ( \35990_nR23b60 , \35989 , \21944 );
buf \U$27964 ( \35991 , \35990_nR23b60 );
not \U$27965 ( \35992 , \35532 );
and \U$27966 ( \35993 , RIe39c680_5865, \35992 );
not \U$27967 ( \35994 , RIe39c680_5865);
or \U$27968 ( \35995 , \35994 , \35147 );
not \U$27969 ( \35996 , \35313 );
and \U$27970 ( \35997 , \33671 , \35996 );
not \U$27971 ( \35998 , \35997 );
not \U$27972 ( \35999 , \35247 );
or \U$27973 ( \36000 , \34868 , \35999 );
nand \U$27974 ( \36001 , \35995 , \35998 , \36000 );
and \U$27975 ( \36002 , \36001 , \35532 );
or \U$27976 ( \36003 , \35993 , \36002 );
and \U$27978 ( \36004 , \36003 , 1'b1 );
or \U$27980 ( \36005 , \36004 , 1'b0 );
buf \U$27981 ( \36006 , \36005 );
_DC r23b62_GF_IsGateDCbyConstraint ( \36007_nR23b62 , \36006 , \21944 );
buf \U$27982 ( \36008 , \36007_nR23b62 );
not \U$27983 ( \36009 , \34698 );
and \U$27984 ( \36010 , RIe39ce78_5866, \36009 );
not \U$27985 ( \36011 , RIe39ce78_5866);
or \U$27986 ( \36012 , \36011 , \35241 );
not \U$27987 ( \36013 , \35313 );
and \U$27988 ( \36014 , \33691 , \36013 );
not \U$27989 ( \36015 , \36014 );
not \U$27990 ( \36016 , \35209 );
or \U$27991 ( \36017 , \34886 , \36016 );
nand \U$27992 ( \36018 , \36012 , \36015 , \36017 );
and \U$27993 ( \36019 , \36018 , \34698 );
or \U$27994 ( \36020 , \36010 , \36019 );
and \U$27996 ( \36021 , \36020 , 1'b1 );
or \U$27998 ( \36022 , \36021 , 1'b0 );
buf \U$27999 ( \36023 , \36022 );
_DC r23b66_GF_IsGateDCbyConstraint ( \36024_nR23b66 , \36023 , \21944 );
buf \U$28000 ( \36025 , \36024_nR23b66 );
not \U$28001 ( \36026 , \33218 );
and \U$28002 ( \36027 , RIe39d670_5867, \36026 );
not \U$28003 ( \36028 , RIe39d670_5867);
or \U$28004 ( \36029 , \36028 , \35223 );
not \U$28005 ( \36030 , \35348 );
and \U$28006 ( \36031 , \33709 , \36030 );
not \U$28007 ( \36032 , \36031 );
not \U$28008 ( \36033 , \35247 );
or \U$28009 ( \36034 , \34904 , \36033 );
nand \U$28010 ( \36035 , \36029 , \36032 , \36034 );
and \U$28011 ( \36036 , \36035 , \33218 );
or \U$28012 ( \36037 , \36027 , \36036 );
and \U$28014 ( \36038 , \36037 , 1'b1 );
or \U$28016 ( \36039 , \36038 , 1'b0 );
buf \U$28017 ( \36040 , \36039 );
_DC r23b68_GF_IsGateDCbyConstraint ( \36041_nR23b68 , \36040 , \21944 );
buf \U$28018 ( \36042 , \36041_nR23b68 );
not \U$28019 ( \36043 , \35532 );
and \U$28020 ( \36044 , RIe39de68_5868, \36043 );
not \U$28021 ( \36045 , RIe39de68_5868);
or \U$28022 ( \36046 , \36045 , \35241 );
not \U$28023 ( \36047 , \35365 );
and \U$28024 ( \36048 , \33728 , \36047 );
not \U$28025 ( \36049 , \36048 );
not \U$28026 ( \36050 , \35247 );
or \U$28027 ( \36051 , \34924 , \36050 );
nand \U$28028 ( \36052 , \36046 , \36049 , \36051 );
and \U$28029 ( \36053 , \36052 , \35532 );
or \U$28030 ( \36054 , \36044 , \36053 );
and \U$28032 ( \36055 , \36054 , 1'b1 );
or \U$28034 ( \36056 , \36055 , 1'b0 );
buf \U$28035 ( \36057 , \36056 );
_DC r23b6a_GF_IsGateDCbyConstraint ( \36058_nR23b6a , \36057 , \21944 );
buf \U$28036 ( \36059 , \36058_nR23b6a );
not \U$28037 ( \36060 , \32755 );
and \U$28038 ( \36061 , RIe39e660_5869, \36060 );
not \U$28039 ( \36062 , RIe39e660_5869);
or \U$28040 ( \36063 , \36062 , \35147 );
not \U$28041 ( \36064 , \35188 );
and \U$28042 ( \36065 , \33746 , \36064 );
not \U$28043 ( \36066 , \36065 );
not \U$28044 ( \36067 , \35209 );
or \U$28045 ( \36068 , \34942 , \36067 );
nand \U$28046 ( \36069 , \36063 , \36066 , \36068 );
and \U$28047 ( \36070 , \36069 , \32755 );
or \U$28048 ( \36071 , \36061 , \36070 );
and \U$28050 ( \36072 , \36071 , 1'b1 );
or \U$28052 ( \36073 , \36072 , 1'b0 );
buf \U$28053 ( \36074 , \36073 );
_DC r23b6c_GF_IsGateDCbyConstraint ( \36075_nR23b6c , \36074 , \21944 );
buf \U$28054 ( \36076 , \36075_nR23b6c );
not \U$28055 ( \36077 , \33218 );
and \U$28056 ( \36078 , RIe39ee58_5870, \36077 );
not \U$28057 ( \36079 , RIe39ee58_5870);
or \U$28058 ( \36080 , \36079 , \35169 );
not \U$28059 ( \36081 , \35348 );
and \U$28060 ( \36082 , \33766 , \36081 );
not \U$28061 ( \36083 , \36082 );
not \U$28062 ( \36084 , \35247 );
or \U$28063 ( \36085 , \34960 , \36084 );
nand \U$28064 ( \36086 , \36080 , \36083 , \36085 );
and \U$28065 ( \36087 , \36086 , \33218 );
or \U$28066 ( \36088 , \36078 , \36087 );
and \U$28068 ( \36089 , \36088 , 1'b1 );
or \U$28070 ( \36090 , \36089 , 1'b0 );
buf \U$28071 ( \36091 , \36090 );
_DC r23b6e_GF_IsGateDCbyConstraint ( \36092_nR23b6e , \36091 , \21944 );
buf \U$28072 ( \36093 , \36092_nR23b6e );
not \U$28073 ( \36094 , \35532 );
and \U$28074 ( \36095 , RIe39f650_5871, \36094 );
not \U$28075 ( \36096 , RIe39f650_5871);
or \U$28076 ( \36097 , \36096 , \35241 );
not \U$28077 ( \36098 , \35188 );
and \U$28078 ( \36099 , \33786 , \36098 );
not \U$28079 ( \36100 , \36099 );
not \U$28080 ( \36101 , \35209 );
or \U$28081 ( \36102 , \34978 , \36101 );
nand \U$28082 ( \36103 , \36097 , \36100 , \36102 );
and \U$28083 ( \36104 , \36103 , \35532 );
or \U$28084 ( \36105 , \36095 , \36104 );
and \U$28086 ( \36106 , \36105 , 1'b1 );
or \U$28088 ( \36107 , \36106 , 1'b0 );
buf \U$28089 ( \36108 , \36107 );
_DC r23b70_GF_IsGateDCbyConstraint ( \36109_nR23b70 , \36108 , \21944 );
buf \U$28090 ( \36110 , \36109_nR23b70 );
not \U$28091 ( \36111 , \34698 );
and \U$28092 ( \36112 , RIe39fe48_5872, \36111 );
not \U$28093 ( \36113 , RIe39fe48_5872);
or \U$28094 ( \36114 , \36113 , \35311 );
not \U$28095 ( \36115 , \35313 );
and \U$28096 ( \36116 , \33805 , \36115 );
not \U$28097 ( \36117 , \36116 );
not \U$28098 ( \36118 , \35209 );
or \U$28099 ( \36119 , \34996 , \36118 );
nand \U$28100 ( \36120 , \36114 , \36117 , \36119 );
and \U$28101 ( \36121 , \36120 , \34698 );
or \U$28102 ( \36122 , \36112 , \36121 );
and \U$28104 ( \36123 , \36122 , 1'b1 );
or \U$28106 ( \36124 , \36123 , 1'b0 );
buf \U$28107 ( \36125 , \36124 );
_DC r23b72_GF_IsGateDCbyConstraint ( \36126_nR23b72 , \36125 , \21944 );
buf \U$28108 ( \36127 , \36126_nR23b72 );
not \U$28109 ( \36128 , \33218 );
and \U$28110 ( \36129 , RIe3a0640_5873, \36128 );
not \U$28111 ( \36130 , RIe3a0640_5873);
or \U$28112 ( \36131 , \36130 , \35223 );
not \U$28113 ( \36132 , \35348 );
and \U$28114 ( \36133 , \33824 , \36132 );
not \U$28115 ( \36134 , \36133 );
not \U$28116 ( \36135 , \35247 );
or \U$28117 ( \36136 , \35014 , \36135 );
nand \U$28118 ( \36137 , \36131 , \36134 , \36136 );
and \U$28119 ( \36138 , \36137 , \33218 );
or \U$28120 ( \36139 , \36129 , \36138 );
and \U$28122 ( \36140 , \36139 , 1'b1 );
or \U$28124 ( \36141 , \36140 , 1'b0 );
buf \U$28125 ( \36142 , \36141 );
_DC r23b74_GF_IsGateDCbyConstraint ( \36143_nR23b74 , \36142 , \21944 );
buf \U$28126 ( \36144 , \36143_nR23b74 );
buf \U$28127 ( \36145 , \34318 );
not \U$28128 ( \36146 , \36145 );
and \U$28129 ( \36147 , RIe3a0e38_5874, \36146 );
not \U$28130 ( \36148 , RIe3a0e38_5874);
or \U$28131 ( \36149 , \36148 , \35169 );
not \U$28132 ( \36150 , \35365 );
and \U$28133 ( \36151 , \33843 , \36150 );
not \U$28134 ( \36152 , \36151 );
not \U$28135 ( \36153 , \35247 );
or \U$28136 ( \36154 , \35032 , \36153 );
nand \U$28137 ( \36155 , \36149 , \36152 , \36154 );
and \U$28138 ( \36156 , \36155 , \36145 );
or \U$28139 ( \36157 , \36147 , \36156 );
and \U$28141 ( \36158 , \36157 , 1'b1 );
or \U$28143 ( \36159 , \36158 , 1'b0 );
buf \U$28144 ( \36160 , \36159 );
_DC r23b76_GF_IsGateDCbyConstraint ( \36161_nR23b76 , \36160 , \21944 );
buf \U$28145 ( \36162 , \36161_nR23b76 );
not \U$28146 ( \36163 , \34698 );
and \U$28147 ( \36164 , RIe3a1630_5875, \36163 );
not \U$28148 ( \36165 , RIe3a1630_5875);
or \U$28149 ( \36166 , \36165 , \35241 );
not \U$28150 ( \36167 , \35150 );
and \U$28151 ( \36168 , \33862 , \36167 );
not \U$28152 ( \36169 , \36168 );
not \U$28153 ( \36170 , \35209 );
or \U$28154 ( \36171 , \35050 , \36170 );
nand \U$28155 ( \36172 , \36166 , \36169 , \36171 );
and \U$28156 ( \36173 , \36172 , \34698 );
or \U$28157 ( \36174 , \36164 , \36173 );
and \U$28159 ( \36175 , \36174 , 1'b1 );
or \U$28161 ( \36176 , \36175 , 1'b0 );
buf \U$28162 ( \36177 , \36176 );
_DC r23b78_GF_IsGateDCbyConstraint ( \36178_nR23b78 , \36177 , \21944 );
buf \U$28163 ( \36179 , \36178_nR23b78 );
not \U$28164 ( \36180 , \33218 );
and \U$28165 ( \36181 , RIe3a1e28_5876, \36180 );
not \U$28166 ( \36182 , RIe3a1e28_5876);
or \U$28167 ( \36183 , \36182 , \35147 );
not \U$28168 ( \36184 , \35313 );
and \U$28169 ( \36185 , \33882 , \36184 );
not \U$28170 ( \36186 , \36185 );
not \U$28171 ( \36187 , \35209 );
or \U$28172 ( \36188 , \35068 , \36187 );
nand \U$28173 ( \36189 , \36183 , \36186 , \36188 );
and \U$28174 ( \36190 , \36189 , \33218 );
or \U$28175 ( \36191 , \36181 , \36190 );
and \U$28177 ( \36192 , \36191 , 1'b1 );
or \U$28179 ( \36193 , \36192 , 1'b0 );
buf \U$28180 ( \36194 , \36193 );
_DC r23b7c_GF_IsGateDCbyConstraint ( \36195_nR23b7c , \36194 , \21944 );
buf \U$28181 ( \36196 , \36195_nR23b7c );
not \U$28182 ( \36197 , \36145 );
and \U$28183 ( \36198 , RIe3a2620_5877, \36197 );
not \U$28184 ( \36199 , RIe3a2620_5877);
or \U$28185 ( \36200 , \36199 , \35311 );
not \U$28186 ( \36201 , \35348 );
and \U$28187 ( \36202 , \33902 , \36201 );
not \U$28188 ( \36203 , \36202 );
not \U$28189 ( \36204 , \35209 );
or \U$28190 ( \36205 , \35086 , \36204 );
nand \U$28191 ( \36206 , \36200 , \36203 , \36205 );
and \U$28192 ( \36207 , \36206 , \36145 );
or \U$28193 ( \36208 , \36198 , \36207 );
and \U$28195 ( \36209 , \36208 , 1'b1 );
or \U$28197 ( \36210 , \36209 , 1'b0 );
buf \U$28198 ( \36211 , \36210 );
_DC r23b7e_GF_IsGateDCbyConstraint ( \36212_nR23b7e , \36211 , \21944 );
buf \U$28199 ( \36213 , \36212_nR23b7e );
not \U$28200 ( \36214 , \34698 );
and \U$28201 ( \36215 , RIe3a2e18_5878, \36214 );
not \U$28202 ( \36216 , RIe3a2e18_5878);
or \U$28203 ( \36217 , \36216 , \35169 );
not \U$28204 ( \36218 , \35243 );
and \U$28205 ( \36219 , \33921 , \36218 );
not \U$28206 ( \36220 , \36219 );
not \U$28207 ( \36221 , \35247 );
or \U$28208 ( \36222 , \35104 , \36221 );
nand \U$28209 ( \36223 , \36217 , \36220 , \36222 );
and \U$28210 ( \36224 , \36223 , \34698 );
or \U$28211 ( \36225 , \36215 , \36224 );
and \U$28213 ( \36226 , \36225 , 1'b1 );
or \U$28215 ( \36227 , \36226 , 1'b0 );
buf \U$28216 ( \36228 , \36227 );
_DC r23b80_GF_IsGateDCbyConstraint ( \36229_nR23b80 , \36228 , \21944 );
buf \U$28217 ( \36230 , \36229_nR23b80 );
not \U$28218 ( \36231 , \33218 );
and \U$28219 ( \36232 , RIe3a3610_5879, \36231 );
not \U$28220 ( \36233 , RIe3a3610_5879);
or \U$28221 ( \36234 , \36233 , \35311 );
not \U$28222 ( \36235 , \35365 );
and \U$28223 ( \36236 , \33940 , \36235 );
not \U$28224 ( \36237 , \36236 );
not \U$28225 ( \36238 , \35247 );
or \U$28226 ( \36239 , \35122 , \36238 );
nand \U$28227 ( \36240 , \36234 , \36237 , \36239 );
and \U$28228 ( \36241 , \36240 , \33218 );
or \U$28229 ( \36242 , \36232 , \36241 );
and \U$28231 ( \36243 , \36242 , 1'b1 );
or \U$28233 ( \36244 , \36243 , 1'b0 );
buf \U$28234 ( \36245 , \36244 );
_DC r23b82_GF_IsGateDCbyConstraint ( \36246_nR23b82 , \36245 , \21944 );
buf \U$28235 ( \36247 , \36246_nR23b82 );
not \U$28236 ( \36248 , \36145 );
and \U$28237 ( \36249 , RIe3a3e08_5880, \36248 );
not \U$28238 ( \36250 , RIe3a3e08_5880);
nand \U$28239 ( \36251 , \32672 , \32670 );
not \U$28240 ( \36252 , \36251 );
nand \U$28241 ( \36253 , \32664 , \36252 );
not \U$28242 ( \36254 , \36253 );
nand \U$28243 ( \36255 , \32680 , \32678 );
not \U$28244 ( \36256 , \32682 );
or \U$28245 ( \36257 , \36255 , \36256 );
not \U$28246 ( \36258 , \36257 );
or \U$28247 ( \36259 , \36254 , \36258 );
buf \U$28248 ( \36260 , \36259 );
or \U$28249 ( \36261 , \36250 , \36260 );
not \U$28250 ( \36262 , \36253 );
buf \U$28251 ( \36263 , \36262 );
nand \U$28252 ( \36264 , \32691 , \36263 );
buf \U$28253 ( \36265 , \36258 );
nand \U$28254 ( \36266 , \32694 , \36265 );
nand \U$28255 ( \36267 , \36261 , \36264 , \36266 );
and \U$28256 ( \36268 , \36267 , \36145 );
or \U$28257 ( \36269 , \36249 , \36268 );
and \U$28259 ( \36270 , \36269 , 1'b1 );
or \U$28261 ( \36271 , \36270 , 1'b0 );
buf \U$28262 ( \36272 , \36271 );
_DC r23b8c_GF_IsGateDCbyConstraint ( \36273_nR23b8c , \36272 , \21944 );
buf \U$28263 ( \36274 , \36273_nR23b8c );
not \U$28264 ( \36275 , \34698 );
and \U$28265 ( \36276 , RIe3a4600_5881, \36275 );
not \U$28266 ( \36277 , RIe3a4600_5881);
buf \U$28267 ( \36278 , \36259 );
or \U$28268 ( \36279 , \36277 , \36278 );
buf \U$28269 ( \36280 , \36262 );
nand \U$28270 ( \36281 , \32719 , \36280 );
nand \U$28271 ( \36282 , \32722 , \36265 );
nand \U$28272 ( \36283 , \36279 , \36281 , \36282 );
and \U$28273 ( \36284 , \36283 , \34698 );
or \U$28274 ( \36285 , \36276 , \36284 );
and \U$28276 ( \36286 , \36285 , 1'b1 );
or \U$28278 ( \36287 , \36286 , 1'b0 );
buf \U$28279 ( \36288 , \36287 );
_DC r23ba2_GF_IsGateDCbyConstraint ( \36289_nR23ba2 , \36288 , \21944 );
buf \U$28280 ( \36290 , \36289_nR23ba2 );
not \U$28281 ( \36291 , \33218 );
and \U$28282 ( \36292 , RIe3a4df8_5882, \36291 );
not \U$28283 ( \36293 , RIe3a4df8_5882);
buf \U$28284 ( \36294 , \36259 );
or \U$28285 ( \36295 , \36293 , \36294 );
nand \U$28286 ( \36296 , \32740 , \36263 );
buf \U$28287 ( \36297 , \36258 );
nand \U$28288 ( \36298 , \32743 , \36297 );
nand \U$28289 ( \36299 , \36295 , \36296 , \36298 );
and \U$28290 ( \36300 , \36299 , \33218 );
or \U$28291 ( \36301 , \36292 , \36300 );
and \U$28293 ( \36302 , \36301 , 1'b1 );
or \U$28295 ( \36303 , \36302 , 1'b0 );
buf \U$28296 ( \36304 , \36303 );
_DC r23bb8_GF_IsGateDCbyConstraint ( \36305_nR23bb8 , \36304 , \21944 );
buf \U$28297 ( \36306 , \36305_nR23bb8 );
not \U$28298 ( \36307 , \36145 );
and \U$28299 ( \36308 , RIe3a55f0_5883, \36307 );
not \U$28300 ( \36309 , RIe3a55f0_5883);
buf \U$28301 ( \36310 , \36259 );
or \U$28302 ( \36311 , \36309 , \36310 );
nand \U$28303 ( \36312 , \32761 , \36280 );
nand \U$28304 ( \36313 , \32764 , \36265 );
nand \U$28305 ( \36314 , \36311 , \36312 , \36313 );
and \U$28306 ( \36315 , \36314 , \36145 );
or \U$28307 ( \36316 , \36308 , \36315 );
and \U$28309 ( \36317 , \36316 , 1'b1 );
or \U$28311 ( \36318 , \36317 , 1'b0 );
buf \U$28312 ( \36319 , \36318 );
_DC r23bce_GF_IsGateDCbyConstraint ( \36320_nR23bce , \36319 , \21944 );
buf \U$28313 ( \36321 , \36320_nR23bce );
not \U$28314 ( \36322 , \34915 );
and \U$28315 ( \36323 , RIe3a5de8_5884, \36322 );
not \U$28316 ( \36324 , RIe3a5de8_5884);
or \U$28317 ( \36325 , \36324 , \36260 );
buf \U$28318 ( \36326 , \36262 );
nand \U$28319 ( \36327 , \32783 , \36326 );
nand \U$28320 ( \36328 , \32786 , \36265 );
nand \U$28321 ( \36329 , \36325 , \36327 , \36328 );
and \U$28322 ( \36330 , \36329 , \34915 );
or \U$28323 ( \36331 , \36323 , \36330 );
and \U$28325 ( \36332 , \36331 , 1'b1 );
or \U$28327 ( \36333 , \36332 , 1'b0 );
buf \U$28328 ( \36334 , \36333 );
_DC r23be4_GF_IsGateDCbyConstraint ( \36335_nR23be4 , \36334 , \21944 );
buf \U$28329 ( \36336 , \36335_nR23be4 );
not \U$28330 ( \36337 , \33218 );
and \U$28331 ( \36338 , RIe3a65e0_5885, \36337 );
not \U$28332 ( \36339 , RIe3a65e0_5885);
or \U$28333 ( \36340 , \36339 , \36278 );
nand \U$28334 ( \36341 , \32804 , \36280 );
buf \U$28335 ( \36342 , \36258 );
nand \U$28336 ( \36343 , \32806 , \36342 );
nand \U$28337 ( \36344 , \36340 , \36341 , \36343 );
and \U$28338 ( \36345 , \36344 , \33218 );
or \U$28339 ( \36346 , \36338 , \36345 );
and \U$28341 ( \36347 , \36346 , 1'b1 );
or \U$28343 ( \36348 , \36347 , 1'b0 );
buf \U$28344 ( \36349 , \36348 );
_DC r23bfa_GF_IsGateDCbyConstraint ( \36350_nR23bfa , \36349 , \21944 );
buf \U$28345 ( \36351 , \36350_nR23bfa );
not \U$28346 ( \36352 , \36145 );
and \U$28347 ( \36353 , RIe3a6dd8_5886, \36352 );
not \U$28348 ( \36354 , RIe3a6dd8_5886);
or \U$28349 ( \36355 , \36354 , \36294 );
nand \U$28350 ( \36356 , \32827 , \36326 );
nand \U$28351 ( \36357 , \32829 , \36342 );
nand \U$28352 ( \36358 , \36355 , \36356 , \36357 );
and \U$28353 ( \36359 , \36358 , \36145 );
or \U$28354 ( \36360 , \36353 , \36359 );
and \U$28356 ( \36361 , \36360 , 1'b1 );
or \U$28358 ( \36362 , \36361 , 1'b0 );
buf \U$28359 ( \36363 , \36362 );
_DC r23c04_GF_IsGateDCbyConstraint ( \36364_nR23c04 , \36363 , \21944 );
buf \U$28360 ( \36365 , \36364_nR23c04 );
not \U$28361 ( \36366 , \34318 );
and \U$28362 ( \36367 , RIe3a75d0_5887, \36366 );
not \U$28363 ( \36368 , RIe3a75d0_5887);
or \U$28364 ( \36369 , \36368 , \36278 );
nand \U$28365 ( \36370 , \32848 , \36280 );
buf \U$28366 ( \36371 , \36258 );
nand \U$28367 ( \36372 , \32851 , \36371 );
nand \U$28368 ( \36373 , \36369 , \36370 , \36372 );
and \U$28369 ( \36374 , \36373 , \34318 );
or \U$28370 ( \36375 , \36367 , \36374 );
and \U$28372 ( \36376 , \36375 , 1'b1 );
or \U$28374 ( \36377 , \36376 , 1'b0 );
buf \U$28375 ( \36378 , \36377 );
_DC r23c06_GF_IsGateDCbyConstraint ( \36379_nR23c06 , \36378 , \21944 );
buf \U$28376 ( \36380 , \36379_nR23c06 );
not \U$28377 ( \36381 , \33218 );
and \U$28378 ( \36382 , RIe3a7dc8_5888, \36381 );
not \U$28379 ( \36383 , RIe3a7dc8_5888);
or \U$28380 ( \36384 , \36383 , \36260 );
nand \U$28381 ( \36385 , \32870 , \36326 );
nand \U$28382 ( \36386 , \32873 , \36297 );
nand \U$28383 ( \36387 , \36384 , \36385 , \36386 );
and \U$28384 ( \36388 , \36387 , \33218 );
or \U$28385 ( \36389 , \36382 , \36388 );
and \U$28387 ( \36390 , \36389 , 1'b1 );
or \U$28389 ( \36391 , \36390 , 1'b0 );
buf \U$28390 ( \36392 , \36391 );
_DC r23c08_GF_IsGateDCbyConstraint ( \36393_nR23c08 , \36392 , \21944 );
buf \U$28391 ( \36394 , \36393_nR23c08 );
not \U$28392 ( \36395 , \36145 );
and \U$28393 ( \36396 , RIe3a85c0_5889, \36395 );
not \U$28394 ( \36397 , RIe3a85c0_5889);
buf \U$28395 ( \36398 , \36259 );
or \U$28396 ( \36399 , \36397 , \36398 );
nand \U$28397 ( \36400 , \32891 , \36280 );
nand \U$28398 ( \36401 , \32894 , \36265 );
nand \U$28399 ( \36402 , \36399 , \36400 , \36401 );
and \U$28400 ( \36403 , \36402 , \36145 );
or \U$28401 ( \36404 , \36396 , \36403 );
and \U$28403 ( \36405 , \36404 , 1'b1 );
or \U$28405 ( \36406 , \36405 , 1'b0 );
buf \U$28406 ( \36407 , \36406 );
_DC r23c0a_GF_IsGateDCbyConstraint ( \36408_nR23c0a , \36407 , \21944 );
buf \U$28407 ( \36409 , \36408_nR23c0a );
not \U$28408 ( \36410 , \34698 );
and \U$28409 ( \36411 , RIe3a8db8_5890, \36410 );
not \U$28410 ( \36412 , RIe3a8db8_5890);
or \U$28411 ( \36413 , \36412 , \36398 );
nand \U$28412 ( \36414 , \32912 , \36263 );
nand \U$28413 ( \36415 , \32914 , \36297 );
nand \U$28414 ( \36416 , \36413 , \36414 , \36415 );
and \U$28415 ( \36417 , \36416 , \34698 );
or \U$28416 ( \36418 , \36411 , \36417 );
and \U$28418 ( \36419 , \36418 , 1'b1 );
or \U$28420 ( \36420 , \36419 , 1'b0 );
buf \U$28421 ( \36421 , \36420 );
_DC r23b8e_GF_IsGateDCbyConstraint ( \36422_nR23b8e , \36421 , \21944 );
buf \U$28422 ( \36423 , \36422_nR23b8e );
not \U$28423 ( \36424 , \33218 );
and \U$28424 ( \36425 , RIe3a95b0_5891, \36424 );
not \U$28425 ( \36426 , RIe3a95b0_5891);
or \U$28426 ( \36427 , \36426 , \36310 );
nand \U$28427 ( \36428 , \32931 , \36263 );
nand \U$28428 ( \36429 , \32934 , \36342 );
nand \U$28429 ( \36430 , \36427 , \36428 , \36429 );
and \U$28430 ( \36431 , \36430 , \33218 );
or \U$28431 ( \36432 , \36425 , \36431 );
and \U$28433 ( \36433 , \36432 , 1'b1 );
or \U$28435 ( \36434 , \36433 , 1'b0 );
buf \U$28436 ( \36435 , \36434 );
_DC r23b90_GF_IsGateDCbyConstraint ( \36436_nR23b90 , \36435 , \21944 );
buf \U$28437 ( \36437 , \36436_nR23b90 );
not \U$28438 ( \36438 , \36145 );
and \U$28439 ( \36439 , RIe3a9da8_5892, \36438 );
not \U$28440 ( \36440 , RIe3a9da8_5892);
or \U$28441 ( \36441 , \36440 , \36294 );
nand \U$28442 ( \36442 , \32951 , \36280 );
nand \U$28443 ( \36443 , \32953 , \36265 );
nand \U$28444 ( \36444 , \36441 , \36442 , \36443 );
and \U$28445 ( \36445 , \36444 , \36145 );
or \U$28446 ( \36446 , \36439 , \36445 );
and \U$28448 ( \36447 , \36446 , 1'b1 );
or \U$28450 ( \36448 , \36447 , 1'b0 );
buf \U$28451 ( \36449 , \36448 );
_DC r23b92_GF_IsGateDCbyConstraint ( \36450_nR23b92 , \36449 , \21944 );
buf \U$28452 ( \36451 , \36450_nR23b92 );
not \U$28453 ( \36452 , \34915 );
and \U$28454 ( \36453 , RIe3aa5a0_5893, \36452 );
not \U$28455 ( \36454 , RIe3aa5a0_5893);
or \U$28456 ( \36455 , \36454 , \36310 );
nand \U$28457 ( \36456 , \32970 , \36280 );
nand \U$28458 ( \36457 , \32973 , \36371 );
nand \U$28459 ( \36458 , \36455 , \36456 , \36457 );
and \U$28460 ( \36459 , \36458 , \34915 );
or \U$28461 ( \36460 , \36453 , \36459 );
and \U$28463 ( \36461 , \36460 , 1'b1 );
or \U$28465 ( \36462 , \36461 , 1'b0 );
buf \U$28466 ( \36463 , \36462 );
_DC r23b94_GF_IsGateDCbyConstraint ( \36464_nR23b94 , \36463 , \21944 );
buf \U$28467 ( \36465 , \36464_nR23b94 );
not \U$28468 ( \36466 , \33218 );
and \U$28469 ( \36467 , RIe3aad98_5894, \36466 );
not \U$28470 ( \36468 , RIe3aad98_5894);
or \U$28471 ( \36469 , \36468 , \36278 );
nand \U$28472 ( \36470 , \32991 , \36326 );
nand \U$28473 ( \36471 , \32994 , \36297 );
nand \U$28474 ( \36472 , \36469 , \36470 , \36471 );
and \U$28475 ( \36473 , \36472 , \33218 );
or \U$28476 ( \36474 , \36467 , \36473 );
and \U$28478 ( \36475 , \36474 , 1'b1 );
or \U$28480 ( \36476 , \36475 , 1'b0 );
buf \U$28481 ( \36477 , \36476 );
_DC r23b96_GF_IsGateDCbyConstraint ( \36478_nR23b96 , \36477 , \21944 );
buf \U$28482 ( \36479 , \36478_nR23b96 );
not \U$28483 ( \36480 , \36145 );
and \U$28484 ( \36481 , RIe3ab590_5895, \36480 );
not \U$28485 ( \36482 , RIe3ab590_5895);
or \U$28486 ( \36483 , \36482 , \36260 );
nand \U$28487 ( \36484 , \33011 , \36262 );
nand \U$28488 ( \36485 , \33014 , \36342 );
nand \U$28489 ( \36486 , \36483 , \36484 , \36485 );
and \U$28490 ( \36487 , \36486 , \36145 );
or \U$28491 ( \36488 , \36481 , \36487 );
and \U$28493 ( \36489 , \36488 , 1'b1 );
or \U$28495 ( \36490 , \36489 , 1'b0 );
buf \U$28496 ( \36491 , \36490 );
_DC r23b98_GF_IsGateDCbyConstraint ( \36492_nR23b98 , \36491 , \21944 );
buf \U$28497 ( \36493 , \36492_nR23b98 );
not \U$28498 ( \36494 , \34318 );
and \U$28499 ( \36495 , RIe3abd88_5896, \36494 );
not \U$28500 ( \36496 , RIe3abd88_5896);
or \U$28501 ( \36497 , \36496 , \36398 );
nand \U$28502 ( \36498 , \33030 , \36326 );
nand \U$28503 ( \36499 , \33033 , \36371 );
nand \U$28504 ( \36500 , \36497 , \36498 , \36499 );
and \U$28505 ( \36501 , \36500 , \34318 );
or \U$28506 ( \36502 , \36495 , \36501 );
and \U$28508 ( \36503 , \36502 , 1'b1 );
or \U$28510 ( \36504 , \36503 , 1'b0 );
buf \U$28511 ( \36505 , \36504 );
_DC r23b9a_GF_IsGateDCbyConstraint ( \36506_nR23b9a , \36505 , \21944 );
buf \U$28512 ( \36507 , \36506_nR23b9a );
not \U$28513 ( \36508 , \32755 );
and \U$28514 ( \36509 , RIe3ac580_5897, \36508 );
not \U$28515 ( \36510 , RIe3ac580_5897);
or \U$28516 ( \36511 , \36510 , \36310 );
nand \U$28517 ( \36512 , \33050 , \36263 );
nand \U$28518 ( \36513 , \33052 , \36342 );
nand \U$28519 ( \36514 , \36511 , \36512 , \36513 );
and \U$28520 ( \36515 , \36514 , \32755 );
or \U$28521 ( \36516 , \36509 , \36515 );
and \U$28523 ( \36517 , \36516 , 1'b1 );
or \U$28525 ( \36518 , \36517 , 1'b0 );
buf \U$28526 ( \36519 , \36518 );
_DC r23b9c_GF_IsGateDCbyConstraint ( \36520_nR23b9c , \36519 , \21944 );
buf \U$28527 ( \36521 , \36520_nR23b9c );
not \U$28528 ( \36522 , \36145 );
and \U$28529 ( \36523 , RIe3acd78_5898, \36522 );
not \U$28530 ( \36524 , RIe3acd78_5898);
or \U$28531 ( \36525 , \36524 , \36294 );
nand \U$28532 ( \36526 , \33069 , \36326 );
nand \U$28533 ( \36527 , \33071 , \36297 );
nand \U$28534 ( \36528 , \36525 , \36526 , \36527 );
and \U$28535 ( \36529 , \36528 , \36145 );
or \U$28536 ( \36530 , \36523 , \36529 );
and \U$28538 ( \36531 , \36530 , 1'b1 );
or \U$28540 ( \36532 , \36531 , 1'b0 );
buf \U$28541 ( \36533 , \36532 );
_DC r23b9e_GF_IsGateDCbyConstraint ( \36534_nR23b9e , \36533 , \21944 );
buf \U$28542 ( \36535 , \36534_nR23b9e );
buf \U$28543 ( \36536 , \34698 );
not \U$28544 ( \36537 , \36536 );
and \U$28545 ( \36538 , RIe3ad570_5899, \36537 );
not \U$28546 ( \36539 , RIe3ad570_5899);
or \U$28547 ( \36540 , \36539 , \36294 );
nand \U$28548 ( \36541 , \33088 , \36262 );
nand \U$28549 ( \36542 , \33091 , \36371 );
nand \U$28550 ( \36543 , \36540 , \36541 , \36542 );
and \U$28551 ( \36544 , \36543 , \36536 );
or \U$28552 ( \36545 , \36538 , \36544 );
and \U$28554 ( \36546 , \36545 , 1'b1 );
or \U$28556 ( \36547 , \36546 , 1'b0 );
buf \U$28557 ( \36548 , \36547 );
_DC r23ba0_GF_IsGateDCbyConstraint ( \36549_nR23ba0 , \36548 , \21944 );
buf \U$28558 ( \36550 , \36549_nR23ba0 );
not \U$28559 ( \36551 , \33296 );
and \U$28560 ( \36552 , RIe3add68_5900, \36551 );
not \U$28561 ( \36553 , RIe3add68_5900);
or \U$28562 ( \36554 , \36553 , \36260 );
nand \U$28563 ( \36555 , \33107 , \36263 );
nand \U$28564 ( \36556 , \33110 , \36342 );
nand \U$28565 ( \36557 , \36554 , \36555 , \36556 );
and \U$28566 ( \36558 , \36557 , \33296 );
or \U$28567 ( \36559 , \36552 , \36558 );
and \U$28569 ( \36560 , \36559 , 1'b1 );
or \U$28571 ( \36561 , \36560 , 1'b0 );
buf \U$28572 ( \36562 , \36561 );
_DC r23ba4_GF_IsGateDCbyConstraint ( \36563_nR23ba4 , \36562 , \21944 );
buf \U$28573 ( \36564 , \36563_nR23ba4 );
not \U$28574 ( \36565 , \36145 );
and \U$28575 ( \36566 , RIe3ae560_5901, \36565 );
not \U$28576 ( \36567 , RIe3ae560_5901);
or \U$28577 ( \36568 , \36567 , \36398 );
nand \U$28578 ( \36569 , \33126 , \36263 );
nand \U$28579 ( \36570 , \33129 , \36265 );
nand \U$28580 ( \36571 , \36568 , \36569 , \36570 );
and \U$28581 ( \36572 , \36571 , \36145 );
or \U$28582 ( \36573 , \36566 , \36572 );
and \U$28584 ( \36574 , \36573 , 1'b1 );
or \U$28586 ( \36575 , \36574 , 1'b0 );
buf \U$28587 ( \36576 , \36575 );
_DC r23ba6_GF_IsGateDCbyConstraint ( \36577_nR23ba6 , \36576 , \21944 );
buf \U$28588 ( \36578 , \36577_nR23ba6 );
not \U$28589 ( \36579 , \36536 );
and \U$28590 ( \36580 , RIe3aed58_5902, \36579 );
not \U$28591 ( \36581 , RIe3aed58_5902);
or \U$28592 ( \36582 , \36581 , \36278 );
nand \U$28593 ( \36583 , \33146 , \36326 );
nand \U$28594 ( \36584 , \33149 , \36265 );
nand \U$28595 ( \36585 , \36582 , \36583 , \36584 );
and \U$28596 ( \36586 , \36585 , \36536 );
or \U$28597 ( \36587 , \36580 , \36586 );
and \U$28599 ( \36588 , \36587 , 1'b1 );
or \U$28601 ( \36589 , \36588 , 1'b0 );
buf \U$28602 ( \36590 , \36589 );
_DC r23ba8_GF_IsGateDCbyConstraint ( \36591_nR23ba8 , \36590 , \21944 );
buf \U$28603 ( \36592 , \36591_nR23ba8 );
not \U$28604 ( \36593 , \33296 );
and \U$28605 ( \36594 , RIe3af550_5903, \36593 );
not \U$28606 ( \36595 , RIe3af550_5903);
or \U$28607 ( \36596 , \36595 , \36310 );
nand \U$28608 ( \36597 , \33165 , \36280 );
nand \U$28609 ( \36598 , \33167 , \36371 );
nand \U$28610 ( \36599 , \36596 , \36597 , \36598 );
and \U$28611 ( \36600 , \36599 , \33296 );
or \U$28612 ( \36601 , \36594 , \36600 );
and \U$28614 ( \36602 , \36601 , 1'b1 );
or \U$28616 ( \36603 , \36602 , 1'b0 );
buf \U$28617 ( \36604 , \36603 );
_DC r23baa_GF_IsGateDCbyConstraint ( \36605_nR23baa , \36604 , \21944 );
buf \U$28618 ( \36606 , \36605_nR23baa );
not \U$28619 ( \36607 , \36145 );
and \U$28620 ( \36608 , RIe3afd48_5904, \36607 );
not \U$28621 ( \36609 , RIe3afd48_5904);
or \U$28622 ( \36610 , \36609 , \36294 );
nand \U$28623 ( \36611 , \33184 , \36262 );
nand \U$28624 ( \36612 , \33187 , \36265 );
nand \U$28625 ( \36613 , \36610 , \36611 , \36612 );
and \U$28626 ( \36614 , \36613 , \36145 );
or \U$28627 ( \36615 , \36608 , \36614 );
and \U$28629 ( \36616 , \36615 , 1'b1 );
or \U$28631 ( \36617 , \36616 , 1'b0 );
buf \U$28632 ( \36618 , \36617 );
_DC r23bac_GF_IsGateDCbyConstraint ( \36619_nR23bac , \36618 , \21944 );
buf \U$28633 ( \36620 , \36619_nR23bac );
not \U$28634 ( \36621 , \36536 );
and \U$28635 ( \36622 , RIe3b0540_5905, \36621 );
not \U$28636 ( \36623 , RIe3b0540_5905);
or \U$28637 ( \36624 , \36623 , \36278 );
nand \U$28638 ( \36625 , \33203 , \36326 );
nand \U$28639 ( \36626 , \33205 , \36265 );
nand \U$28640 ( \36627 , \36624 , \36625 , \36626 );
and \U$28641 ( \36628 , \36627 , \36536 );
or \U$28642 ( \36629 , \36622 , \36628 );
and \U$28644 ( \36630 , \36629 , 1'b1 );
or \U$28646 ( \36631 , \36630 , 1'b0 );
buf \U$28647 ( \36632 , \36631 );
_DC r23bae_GF_IsGateDCbyConstraint ( \36633_nR23bae , \36632 , \21944 );
buf \U$28648 ( \36634 , \36633_nR23bae );
not \U$28649 ( \36635 , \33568 );
and \U$28650 ( \36636 , RIe3b0d38_5906, \36635 );
not \U$28651 ( \36637 , RIe3b0d38_5906);
or \U$28652 ( \36638 , \36637 , \36260 );
nand \U$28653 ( \36639 , \33223 , \36263 );
nand \U$28654 ( \36640 , \33226 , \36297 );
nand \U$28655 ( \36641 , \36638 , \36639 , \36640 );
and \U$28656 ( \36642 , \36641 , \33568 );
or \U$28657 ( \36643 , \36636 , \36642 );
and \U$28659 ( \36644 , \36643 , 1'b1 );
or \U$28661 ( \36645 , \36644 , 1'b0 );
buf \U$28662 ( \36646 , \36645 );
_DC r23bb0_GF_IsGateDCbyConstraint ( \36647_nR23bb0 , \36646 , \21944 );
buf \U$28663 ( \36648 , \36647_nR23bb0 );
not \U$28664 ( \36649 , \36145 );
and \U$28665 ( \36650 , RIe3b1530_5907, \36649 );
not \U$28666 ( \36651 , RIe3b1530_5907);
or \U$28667 ( \36652 , \36651 , \36260 );
nand \U$28668 ( \36653 , \33242 , \36262 );
nand \U$28669 ( \36654 , \33245 , \36265 );
nand \U$28670 ( \36655 , \36652 , \36653 , \36654 );
and \U$28671 ( \36656 , \36655 , \36145 );
or \U$28672 ( \36657 , \36650 , \36656 );
and \U$28674 ( \36658 , \36657 , 1'b1 );
or \U$28676 ( \36659 , \36658 , 1'b0 );
buf \U$28677 ( \36660 , \36659 );
_DC r23bb2_GF_IsGateDCbyConstraint ( \36661_nR23bb2 , \36660 , \21944 );
buf \U$28678 ( \36662 , \36661_nR23bb2 );
not \U$28679 ( \36663 , \36536 );
and \U$28680 ( \36664 , RIe3b1d28_5908, \36663 );
not \U$28681 ( \36665 , RIe3b1d28_5908);
or \U$28682 ( \36666 , \36665 , \36398 );
nand \U$28683 ( \36667 , \33262 , \36262 );
nand \U$28684 ( \36668 , \33265 , \36371 );
nand \U$28685 ( \36669 , \36666 , \36667 , \36668 );
and \U$28686 ( \36670 , \36669 , \36536 );
or \U$28687 ( \36671 , \36664 , \36670 );
and \U$28689 ( \36672 , \36671 , 1'b1 );
or \U$28691 ( \36673 , \36672 , 1'b0 );
buf \U$28692 ( \36674 , \36673 );
_DC r23bb4_GF_IsGateDCbyConstraint ( \36675_nR23bb4 , \36674 , \21944 );
buf \U$28693 ( \36676 , \36675_nR23bb4 );
not \U$28694 ( \36677 , \34915 );
and \U$28695 ( \36678 , RIe3b2520_5909, \36677 );
not \U$28696 ( \36679 , RIe3b2520_5909);
or \U$28697 ( \36680 , \36679 , \36310 );
nand \U$28698 ( \36681 , \33281 , \36263 );
nand \U$28699 ( \36682 , \33284 , \36371 );
nand \U$28700 ( \36683 , \36680 , \36681 , \36682 );
and \U$28701 ( \36684 , \36683 , \34915 );
or \U$28702 ( \36685 , \36678 , \36684 );
and \U$28704 ( \36686 , \36685 , 1'b1 );
or \U$28706 ( \36687 , \36686 , 1'b0 );
buf \U$28707 ( \36688 , \36687 );
_DC r23bb6_GF_IsGateDCbyConstraint ( \36689_nR23bb6 , \36688 , \21944 );
buf \U$28708 ( \36690 , \36689_nR23bb6 );
buf \U$28709 ( \36691 , \34915 );
not \U$28710 ( \36692 , \36691 );
and \U$28711 ( \36693 , RIe3b2d18_5910, \36692 );
not \U$28712 ( \36694 , RIe3b2d18_5910);
or \U$28713 ( \36695 , \36694 , \36278 );
nand \U$28714 ( \36696 , \33303 , \36263 );
nand \U$28715 ( \36697 , \33305 , \36342 );
nand \U$28716 ( \36698 , \36695 , \36696 , \36697 );
and \U$28717 ( \36699 , \36698 , \36691 );
or \U$28718 ( \36700 , \36693 , \36699 );
and \U$28720 ( \36701 , \36700 , 1'b1 );
or \U$28722 ( \36702 , \36701 , 1'b0 );
buf \U$28723 ( \36703 , \36702 );
_DC r23bba_GF_IsGateDCbyConstraint ( \36704_nR23bba , \36703 , \21944 );
buf \U$28724 ( \36705 , \36704_nR23bba );
not \U$28725 ( \36706 , \36536 );
and \U$28726 ( \36707 , RIe3b3510_5911, \36706 );
not \U$28727 ( \36708 , RIe3b3510_5911);
or \U$28728 ( \36709 , \36708 , \36398 );
nand \U$28729 ( \36710 , \33321 , \36262 );
nand \U$28730 ( \36711 , \33324 , \36297 );
nand \U$28731 ( \36712 , \36709 , \36710 , \36711 );
and \U$28732 ( \36713 , \36712 , \36536 );
or \U$28733 ( \36714 , \36707 , \36713 );
and \U$28735 ( \36715 , \36714 , 1'b1 );
or \U$28737 ( \36716 , \36715 , 1'b0 );
buf \U$28738 ( \36717 , \36716 );
_DC r23bbc_GF_IsGateDCbyConstraint ( \36718_nR23bbc , \36717 , \21944 );
buf \U$28739 ( \36719 , \36718_nR23bbc );
not \U$28740 ( \36720 , \33568 );
and \U$28741 ( \36721 , RIe3b3d08_5912, \36720 );
not \U$28742 ( \36722 , RIe3b3d08_5912);
or \U$28743 ( \36723 , \36722 , \36260 );
nand \U$28744 ( \36724 , \33341 , \36263 );
nand \U$28745 ( \36725 , \33344 , \36371 );
nand \U$28746 ( \36726 , \36723 , \36724 , \36725 );
and \U$28747 ( \36727 , \36726 , \33568 );
or \U$28748 ( \36728 , \36721 , \36727 );
and \U$28750 ( \36729 , \36728 , 1'b1 );
or \U$28752 ( \36730 , \36729 , 1'b0 );
buf \U$28753 ( \36731 , \36730 );
_DC r23bbe_GF_IsGateDCbyConstraint ( \36732_nR23bbe , \36731 , \21944 );
buf \U$28754 ( \36733 , \36732_nR23bbe );
not \U$28755 ( \36734 , \36691 );
and \U$28756 ( \36735 , RIe3b4500_5913, \36734 );
not \U$28757 ( \36736 , RIe3b4500_5913);
or \U$28758 ( \36737 , \36736 , \36398 );
nand \U$28759 ( \36738 , \33360 , \36326 );
nand \U$28760 ( \36739 , \33363 , \36371 );
nand \U$28761 ( \36740 , \36737 , \36738 , \36739 );
and \U$28762 ( \36741 , \36740 , \36691 );
or \U$28763 ( \36742 , \36735 , \36741 );
and \U$28765 ( \36743 , \36742 , 1'b1 );
or \U$28767 ( \36744 , \36743 , 1'b0 );
buf \U$28768 ( \36745 , \36744 );
_DC r23bc0_GF_IsGateDCbyConstraint ( \36746_nR23bc0 , \36745 , \21944 );
buf \U$28769 ( \36747 , \36746_nR23bc0 );
not \U$28770 ( \36748 , \36536 );
and \U$28771 ( \36749 , RIe3b4cf8_5914, \36748 );
not \U$28772 ( \36750 , RIe3b4cf8_5914);
or \U$28773 ( \36751 , \36750 , \36310 );
nand \U$28774 ( \36752 , \33379 , \36263 );
nand \U$28775 ( \36753 , \33382 , \36342 );
nand \U$28776 ( \36754 , \36751 , \36752 , \36753 );
and \U$28777 ( \36755 , \36754 , \36536 );
or \U$28778 ( \36756 , \36749 , \36755 );
and \U$28780 ( \36757 , \36756 , 1'b1 );
or \U$28782 ( \36758 , \36757 , 1'b0 );
buf \U$28783 ( \36759 , \36758 );
_DC r23bc2_GF_IsGateDCbyConstraint ( \36760_nR23bc2 , \36759 , \21944 );
buf \U$28784 ( \36761 , \36760_nR23bc2 );
not \U$28785 ( \36762 , \33568 );
and \U$28786 ( \36763 , RIe3b54f0_5915, \36762 );
not \U$28787 ( \36764 , RIe3b54f0_5915);
or \U$28788 ( \36765 , \36764 , \36294 );
nand \U$28789 ( \36766 , \33399 , \36263 );
nand \U$28790 ( \36767 , \33402 , \36297 );
nand \U$28791 ( \36768 , \36765 , \36766 , \36767 );
and \U$28792 ( \36769 , \36768 , \33568 );
or \U$28793 ( \36770 , \36763 , \36769 );
and \U$28795 ( \36771 , \36770 , 1'b1 );
or \U$28797 ( \36772 , \36771 , 1'b0 );
buf \U$28798 ( \36773 , \36772 );
_DC r23bc4_GF_IsGateDCbyConstraint ( \36774_nR23bc4 , \36773 , \21944 );
buf \U$28799 ( \36775 , \36774_nR23bc4 );
not \U$28800 ( \36776 , \36691 );
and \U$28801 ( \36777 , RIe3b5ce8_5916, \36776 );
not \U$28802 ( \36778 , RIe3b5ce8_5916);
or \U$28803 ( \36779 , \36778 , \36310 );
nand \U$28804 ( \36780 , \33419 , \36262 );
nand \U$28805 ( \36781 , \33422 , \36297 );
nand \U$28806 ( \36782 , \36779 , \36780 , \36781 );
and \U$28807 ( \36783 , \36782 , \36691 );
or \U$28808 ( \36784 , \36777 , \36783 );
and \U$28810 ( \36785 , \36784 , 1'b1 );
or \U$28812 ( \36786 , \36785 , 1'b0 );
buf \U$28813 ( \36787 , \36786 );
_DC r23bc6_GF_IsGateDCbyConstraint ( \36788_nR23bc6 , \36787 , \21944 );
buf \U$28814 ( \36789 , \36788_nR23bc6 );
not \U$28815 ( \36790 , \36536 );
and \U$28816 ( \36791 , RIe3b64e0_5917, \36790 );
not \U$28817 ( \36792 , RIe3b64e0_5917);
or \U$28818 ( \36793 , \36792 , \36278 );
nand \U$28819 ( \36794 , \33438 , \36263 );
nand \U$28820 ( \36795 , \33440 , \36342 );
nand \U$28821 ( \36796 , \36793 , \36794 , \36795 );
and \U$28822 ( \36797 , \36796 , \36536 );
or \U$28823 ( \36798 , \36791 , \36797 );
and \U$28825 ( \36799 , \36798 , 1'b1 );
or \U$28827 ( \36800 , \36799 , 1'b0 );
buf \U$28828 ( \36801 , \36800 );
_DC r23bc8_GF_IsGateDCbyConstraint ( \36802_nR23bc8 , \36801 , \21944 );
buf \U$28829 ( \36803 , \36802_nR23bc8 );
not \U$28830 ( \36804 , \32755 );
and \U$28831 ( \36805 , RIe3b6cd8_5918, \36804 );
not \U$28832 ( \36806 , RIe3b6cd8_5918);
or \U$28833 ( \36807 , \36806 , \36260 );
nand \U$28834 ( \36808 , \33456 , \36263 );
nand \U$28835 ( \36809 , \33459 , \36297 );
nand \U$28836 ( \36810 , \36807 , \36808 , \36809 );
and \U$28837 ( \36811 , \36810 , \32755 );
or \U$28838 ( \36812 , \36805 , \36811 );
and \U$28840 ( \36813 , \36812 , 1'b1 );
or \U$28842 ( \36814 , \36813 , 1'b0 );
buf \U$28843 ( \36815 , \36814 );
_DC r23bca_GF_IsGateDCbyConstraint ( \36816_nR23bca , \36815 , \21944 );
buf \U$28844 ( \36817 , \36816_nR23bca );
not \U$28845 ( \36818 , \36691 );
and \U$28846 ( \36819 , RIe3b74d0_5919, \36818 );
not \U$28847 ( \36820 , RIe3b74d0_5919);
or \U$28848 ( \36821 , \36820 , \36398 );
nand \U$28849 ( \36822 , \33475 , \36280 );
nand \U$28850 ( \36823 , \33478 , \36297 );
nand \U$28851 ( \36824 , \36821 , \36822 , \36823 );
and \U$28852 ( \36825 , \36824 , \36691 );
or \U$28853 ( \36826 , \36819 , \36825 );
and \U$28855 ( \36827 , \36826 , 1'b1 );
or \U$28857 ( \36828 , \36827 , 1'b0 );
buf \U$28858 ( \36829 , \36828 );
_DC r23bcc_GF_IsGateDCbyConstraint ( \36830_nR23bcc , \36829 , \21944 );
buf \U$28859 ( \36831 , \36830_nR23bcc );
not \U$28860 ( \36832 , \36536 );
and \U$28861 ( \36833 , RIe3b7cc8_5920, \36832 );
not \U$28862 ( \36834 , RIe3b7cc8_5920);
or \U$28863 ( \36835 , \36834 , \36294 );
nand \U$28864 ( \36836 , \33494 , \36280 );
nand \U$28865 ( \36837 , \33497 , \36371 );
nand \U$28866 ( \36838 , \36835 , \36836 , \36837 );
and \U$28867 ( \36839 , \36838 , \36536 );
or \U$28868 ( \36840 , \36833 , \36839 );
and \U$28870 ( \36841 , \36840 , 1'b1 );
or \U$28872 ( \36842 , \36841 , 1'b0 );
buf \U$28873 ( \36843 , \36842 );
_DC r23bd0_GF_IsGateDCbyConstraint ( \36844_nR23bd0 , \36843 , \21944 );
buf \U$28874 ( \36845 , \36844_nR23bd0 );
not \U$28875 ( \36846 , \33296 );
and \U$28876 ( \36847 , RIe3b84c0_5921, \36846 );
not \U$28877 ( \36848 , RIe3b84c0_5921);
or \U$28878 ( \36849 , \36848 , \36294 );
nand \U$28879 ( \36850 , \33514 , \36326 );
nand \U$28880 ( \36851 , \33517 , \36265 );
nand \U$28881 ( \36852 , \36849 , \36850 , \36851 );
and \U$28882 ( \36853 , \36852 , \33296 );
or \U$28883 ( \36854 , \36847 , \36853 );
and \U$28885 ( \36855 , \36854 , 1'b1 );
or \U$28887 ( \36856 , \36855 , 1'b0 );
buf \U$28888 ( \36857 , \36856 );
_DC r23bd2_GF_IsGateDCbyConstraint ( \36858_nR23bd2 , \36857 , \21944 );
buf \U$28889 ( \36859 , \36858_nR23bd2 );
not \U$28890 ( \36860 , \36691 );
and \U$28891 ( \36861 , RIe3b8cb8_5922, \36860 );
not \U$28892 ( \36862 , RIe3b8cb8_5922);
or \U$28893 ( \36863 , \36862 , \36278 );
nand \U$28894 ( \36864 , \33534 , \36263 );
nand \U$28895 ( \36865 , \33537 , \36297 );
nand \U$28896 ( \36866 , \36863 , \36864 , \36865 );
and \U$28897 ( \36867 , \36866 , \36691 );
or \U$28898 ( \36868 , \36861 , \36867 );
and \U$28900 ( \36869 , \36868 , 1'b1 );
or \U$28902 ( \36870 , \36869 , 1'b0 );
buf \U$28903 ( \36871 , \36870 );
_DC r23bd4_GF_IsGateDCbyConstraint ( \36872_nR23bd4 , \36871 , \21944 );
buf \U$28904 ( \36873 , \36872_nR23bd4 );
not \U$28905 ( \36874 , \36536 );
and \U$28906 ( \36875 , RIe3b94b0_5923, \36874 );
not \U$28907 ( \36876 , RIe3b94b0_5923);
or \U$28908 ( \36877 , \36876 , \36260 );
nand \U$28909 ( \36878 , \33553 , \36262 );
nand \U$28910 ( \36879 , \33556 , \36371 );
nand \U$28911 ( \36880 , \36877 , \36878 , \36879 );
and \U$28912 ( \36881 , \36880 , \36536 );
or \U$28913 ( \36882 , \36875 , \36881 );
and \U$28915 ( \36883 , \36882 , 1'b1 );
or \U$28917 ( \36884 , \36883 , 1'b0 );
buf \U$28918 ( \36885 , \36884 );
_DC r23bd6_GF_IsGateDCbyConstraint ( \36886_nR23bd6 , \36885 , \21944 );
buf \U$28919 ( \36887 , \36886_nR23bd6 );
not \U$28920 ( \36888 , \33568 );
and \U$28921 ( \36889 , RIe3b9ca8_5924, \36888 );
not \U$28922 ( \36890 , RIe3b9ca8_5924);
or \U$28923 ( \36891 , \36890 , \36398 );
nand \U$28924 ( \36892 , \33574 , \36280 );
nand \U$28925 ( \36893 , \33576 , \36371 );
nand \U$28926 ( \36894 , \36891 , \36892 , \36893 );
and \U$28927 ( \36895 , \36894 , \33568 );
or \U$28928 ( \36896 , \36889 , \36895 );
and \U$28930 ( \36897 , \36896 , 1'b1 );
or \U$28932 ( \36898 , \36897 , 1'b0 );
buf \U$28933 ( \36899 , \36898 );
_DC r23bd8_GF_IsGateDCbyConstraint ( \36900_nR23bd8 , \36899 , \21944 );
buf \U$28934 ( \36901 , \36900_nR23bd8 );
not \U$28935 ( \36902 , \36691 );
and \U$28936 ( \36903 , RIe3ba4a0_5925, \36902 );
not \U$28937 ( \36904 , RIe3ba4a0_5925);
or \U$28938 ( \36905 , \36904 , \36278 );
nand \U$28939 ( \36906 , \33592 , \36326 );
nand \U$28940 ( \36907 , \33594 , \36297 );
nand \U$28941 ( \36908 , \36905 , \36906 , \36907 );
and \U$28942 ( \36909 , \36908 , \36691 );
or \U$28943 ( \36910 , \36903 , \36909 );
and \U$28945 ( \36911 , \36910 , 1'b1 );
or \U$28947 ( \36912 , \36911 , 1'b0 );
buf \U$28948 ( \36913 , \36912 );
_DC r23bda_GF_IsGateDCbyConstraint ( \36914_nR23bda , \36913 , \21944 );
buf \U$28949 ( \36915 , \36914_nR23bda );
not \U$28950 ( \36916 , \36536 );
and \U$28951 ( \36917 , RIe3bac98_5926, \36916 );
not \U$28952 ( \36918 , RIe3bac98_5926);
or \U$28953 ( \36919 , \36918 , \36310 );
nand \U$28954 ( \36920 , \33610 , \36280 );
nand \U$28955 ( \36921 , \33612 , \36297 );
nand \U$28956 ( \36922 , \36919 , \36920 , \36921 );
and \U$28957 ( \36923 , \36922 , \36536 );
or \U$28958 ( \36924 , \36917 , \36923 );
and \U$28960 ( \36925 , \36924 , 1'b1 );
or \U$28962 ( \36926 , \36925 , 1'b0 );
buf \U$28963 ( \36927 , \36926 );
_DC r23bdc_GF_IsGateDCbyConstraint ( \36928_nR23bdc , \36927 , \21944 );
buf \U$28964 ( \36929 , \36928_nR23bdc );
not \U$28965 ( \36930 , \34915 );
and \U$28966 ( \36931 , RIe3bb490_5927, \36930 );
not \U$28967 ( \36932 , RIe3bb490_5927);
or \U$28968 ( \36933 , \36932 , \36294 );
nand \U$28969 ( \36934 , \33629 , \36280 );
nand \U$28970 ( \36935 , \33632 , \36265 );
nand \U$28971 ( \36936 , \36933 , \36934 , \36935 );
and \U$28972 ( \36937 , \36936 , \34915 );
or \U$28973 ( \36938 , \36931 , \36937 );
and \U$28975 ( \36939 , \36938 , 1'b1 );
or \U$28977 ( \36940 , \36939 , 1'b0 );
buf \U$28978 ( \36941 , \36940 );
_DC r23bde_GF_IsGateDCbyConstraint ( \36942_nR23bde , \36941 , \21944 );
buf \U$28979 ( \36943 , \36942_nR23bde );
not \U$28980 ( \36944 , \36691 );
and \U$28981 ( \36945 , RIe3bbc88_5928, \36944 );
not \U$28982 ( \36946 , RIe3bbc88_5928);
or \U$28983 ( \36947 , \36946 , \36278 );
nand \U$28984 ( \36948 , \33648 , \36263 );
nand \U$28985 ( \36949 , \33651 , \36371 );
nand \U$28986 ( \36950 , \36947 , \36948 , \36949 );
and \U$28987 ( \36951 , \36950 , \36691 );
or \U$28988 ( \36952 , \36945 , \36951 );
and \U$28990 ( \36953 , \36952 , 1'b1 );
or \U$28992 ( \36954 , \36953 , 1'b0 );
buf \U$28993 ( \36955 , \36954 );
_DC r23be0_GF_IsGateDCbyConstraint ( \36956_nR23be0 , \36955 , \21944 );
buf \U$28994 ( \36957 , \36956_nR23be0 );
not \U$28995 ( \36958 , \36536 );
and \U$28996 ( \36959 , RIe3bc480_5929, \36958 );
not \U$28997 ( \36960 , RIe3bc480_5929);
or \U$28998 ( \36961 , \36960 , \36260 );
nand \U$28999 ( \36962 , \33668 , \36326 );
nand \U$29000 ( \36963 , \33671 , \36265 );
nand \U$29001 ( \36964 , \36961 , \36962 , \36963 );
and \U$29002 ( \36965 , \36964 , \36536 );
or \U$29003 ( \36966 , \36959 , \36965 );
and \U$29005 ( \36967 , \36966 , 1'b1 );
or \U$29007 ( \36968 , \36967 , 1'b0 );
buf \U$29008 ( \36969 , \36968 );
_DC r23be2_GF_IsGateDCbyConstraint ( \36970_nR23be2 , \36969 , \21944 );
buf \U$29009 ( \36971 , \36970_nR23be2 );
not \U$29010 ( \36972 , \32755 );
and \U$29011 ( \36973 , RIe3bcc78_5930, \36972 );
not \U$29012 ( \36974 , RIe3bcc78_5930);
or \U$29013 ( \36975 , \36974 , \36398 );
nand \U$29014 ( \36976 , \33688 , \36280 );
nand \U$29015 ( \36977 , \33691 , \36265 );
nand \U$29016 ( \36978 , \36975 , \36976 , \36977 );
and \U$29017 ( \36979 , \36978 , \32755 );
or \U$29018 ( \36980 , \36973 , \36979 );
and \U$29020 ( \36981 , \36980 , 1'b1 );
or \U$29022 ( \36982 , \36981 , 1'b0 );
buf \U$29023 ( \36983 , \36982 );
_DC r23be6_GF_IsGateDCbyConstraint ( \36984_nR23be6 , \36983 , \21944 );
buf \U$29024 ( \36985 , \36984_nR23be6 );
not \U$29025 ( \36986 , \36691 );
and \U$29026 ( \36987 , RIe3bd470_5931, \36986 );
not \U$29027 ( \36988 , RIe3bd470_5931);
or \U$29028 ( \36989 , \36988 , \36310 );
nand \U$29029 ( \36990 , \33707 , \36263 );
nand \U$29030 ( \36991 , \33709 , \36342 );
nand \U$29031 ( \36992 , \36989 , \36990 , \36991 );
and \U$29032 ( \36993 , \36992 , \36691 );
or \U$29033 ( \36994 , \36987 , \36993 );
and \U$29035 ( \36995 , \36994 , 1'b1 );
or \U$29037 ( \36996 , \36995 , 1'b0 );
buf \U$29038 ( \36997 , \36996 );
_DC r23be8_GF_IsGateDCbyConstraint ( \36998_nR23be8 , \36997 , \21944 );
buf \U$29039 ( \36999 , \36998_nR23be8 );
not \U$29040 ( \37000 , \36536 );
and \U$29041 ( \37001 , RIe3bdc68_5932, \37000 );
not \U$29042 ( \37002 , RIe3bdc68_5932);
or \U$29043 ( \37003 , \37002 , \36294 );
nand \U$29044 ( \37004 , \33725 , \36280 );
nand \U$29045 ( \37005 , \33728 , \36371 );
nand \U$29046 ( \37006 , \37003 , \37004 , \37005 );
and \U$29047 ( \37007 , \37006 , \36536 );
or \U$29048 ( \37008 , \37001 , \37007 );
and \U$29050 ( \37009 , \37008 , 1'b1 );
or \U$29052 ( \37010 , \37009 , 1'b0 );
buf \U$29053 ( \37011 , \37010 );
_DC r23bea_GF_IsGateDCbyConstraint ( \37012_nR23bea , \37011 , \21944 );
buf \U$29054 ( \37013 , \37012_nR23bea );
not \U$29055 ( \37014 , \34318 );
and \U$29056 ( \37015 , RIe3be460_5933, \37014 );
not \U$29057 ( \37016 , RIe3be460_5933);
or \U$29058 ( \37017 , \37016 , \36278 );
nand \U$29059 ( \37018 , \33744 , \36326 );
nand \U$29060 ( \37019 , \33746 , \36342 );
nand \U$29061 ( \37020 , \37017 , \37018 , \37019 );
and \U$29062 ( \37021 , \37020 , \34318 );
or \U$29063 ( \37022 , \37015 , \37021 );
and \U$29065 ( \37023 , \37022 , 1'b1 );
or \U$29067 ( \37024 , \37023 , 1'b0 );
buf \U$29068 ( \37025 , \37024 );
_DC r23bec_GF_IsGateDCbyConstraint ( \37026_nR23bec , \37025 , \21944 );
buf \U$29069 ( \37027 , \37026_nR23bec );
not \U$29070 ( \37028 , \36691 );
and \U$29071 ( \37029 , RIe3bec58_5934, \37028 );
not \U$29072 ( \37030 , RIe3bec58_5934);
or \U$29073 ( \37031 , \37030 , \36398 );
nand \U$29074 ( \37032 , \33763 , \36280 );
nand \U$29075 ( \37033 , \33766 , \36342 );
nand \U$29076 ( \37034 , \37031 , \37032 , \37033 );
and \U$29077 ( \37035 , \37034 , \36691 );
or \U$29078 ( \37036 , \37029 , \37035 );
and \U$29080 ( \37037 , \37036 , 1'b1 );
or \U$29082 ( \37038 , \37037 , 1'b0 );
buf \U$29083 ( \37039 , \37038 );
_DC r23bee_GF_IsGateDCbyConstraint ( \37040_nR23bee , \37039 , \21944 );
buf \U$29084 ( \37041 , \37040_nR23bee );
not \U$29085 ( \37042 , \32756 );
and \U$29086 ( \37043 , RIe3bf450_5935, \37042 );
not \U$29087 ( \37044 , RIe3bf450_5935);
or \U$29088 ( \37045 , \37044 , \36260 );
nand \U$29089 ( \37046 , \33783 , \36326 );
nand \U$29090 ( \37047 , \33786 , \36371 );
nand \U$29091 ( \37048 , \37045 , \37046 , \37047 );
and \U$29092 ( \37049 , \37048 , \32756 );
or \U$29093 ( \37050 , \37043 , \37049 );
and \U$29095 ( \37051 , \37050 , 1'b1 );
or \U$29097 ( \37052 , \37051 , 1'b0 );
buf \U$29098 ( \37053 , \37052 );
_DC r23bf0_GF_IsGateDCbyConstraint ( \37054_nR23bf0 , \37053 , \21944 );
buf \U$29099 ( \37055 , \37054_nR23bf0 );
not \U$29100 ( \37056 , \34318 );
and \U$29101 ( \37057 , RIe3bfc48_5936, \37056 );
not \U$29102 ( \37058 , RIe3bfc48_5936);
or \U$29103 ( \37059 , \37058 , \36398 );
nand \U$29104 ( \37060 , \33802 , \36326 );
nand \U$29105 ( \37061 , \33805 , \36342 );
nand \U$29106 ( \37062 , \37059 , \37060 , \37061 );
and \U$29107 ( \37063 , \37062 , \34318 );
or \U$29108 ( \37064 , \37057 , \37063 );
and \U$29110 ( \37065 , \37064 , 1'b1 );
or \U$29112 ( \37066 , \37065 , 1'b0 );
buf \U$29113 ( \37067 , \37066 );
_DC r23bf2_GF_IsGateDCbyConstraint ( \37068_nR23bf2 , \37067 , \21944 );
buf \U$29114 ( \37069 , \37068_nR23bf2 );
not \U$29115 ( \37070 , \36691 );
and \U$29116 ( \37071 , RIe3c0440_5937, \37070 );
not \U$29117 ( \37072 , RIe3c0440_5937);
or \U$29118 ( \37073 , \37072 , \36310 );
nand \U$29119 ( \37074 , \33821 , \36280 );
nand \U$29120 ( \37075 , \33824 , \36265 );
nand \U$29121 ( \37076 , \37073 , \37074 , \37075 );
and \U$29122 ( \37077 , \37076 , \36691 );
or \U$29123 ( \37078 , \37071 , \37077 );
and \U$29125 ( \37079 , \37078 , 1'b1 );
or \U$29127 ( \37080 , \37079 , 1'b0 );
buf \U$29128 ( \37081 , \37080 );
_DC r23bf4_GF_IsGateDCbyConstraint ( \37082_nR23bf4 , \37081 , \21944 );
buf \U$29129 ( \37083 , \37082_nR23bf4 );
not \U$29130 ( \37084 , \32756 );
and \U$29131 ( \37085 , RIe3c0c38_5938, \37084 );
not \U$29132 ( \37086 , RIe3c0c38_5938);
or \U$29133 ( \37087 , \37086 , \36294 );
nand \U$29134 ( \37088 , \33840 , \36280 );
nand \U$29135 ( \37089 , \33843 , \36371 );
nand \U$29136 ( \37090 , \37087 , \37088 , \37089 );
and \U$29137 ( \37091 , \37090 , \32756 );
or \U$29138 ( \37092 , \37085 , \37091 );
and \U$29140 ( \37093 , \37092 , 1'b1 );
or \U$29142 ( \37094 , \37093 , 1'b0 );
buf \U$29143 ( \37095 , \37094 );
_DC r23bf6_GF_IsGateDCbyConstraint ( \37096_nR23bf6 , \37095 , \21944 );
buf \U$29144 ( \37097 , \37096_nR23bf6 );
not \U$29145 ( \37098 , \34318 );
and \U$29146 ( \37099 , RIe3c1430_5939, \37098 );
not \U$29147 ( \37100 , RIe3c1430_5939);
or \U$29148 ( \37101 , \37100 , \36310 );
nand \U$29149 ( \37102 , \33859 , \36326 );
nand \U$29150 ( \37103 , \33862 , \36297 );
nand \U$29151 ( \37104 , \37101 , \37102 , \37103 );
and \U$29152 ( \37105 , \37104 , \34318 );
or \U$29153 ( \37106 , \37099 , \37105 );
and \U$29155 ( \37107 , \37106 , 1'b1 );
or \U$29157 ( \37108 , \37107 , 1'b0 );
buf \U$29158 ( \37109 , \37108 );
_DC r23bf8_GF_IsGateDCbyConstraint ( \37110_nR23bf8 , \37109 , \21944 );
buf \U$29159 ( \37111 , \37110_nR23bf8 );
not \U$29160 ( \37112 , \36691 );
and \U$29161 ( \37113 , RIe3c1c28_5940, \37112 );
not \U$29162 ( \37114 , RIe3c1c28_5940);
or \U$29163 ( \37115 , \37114 , \36260 );
nand \U$29164 ( \37116 , \33879 , \36326 );
nand \U$29165 ( \37117 , \33882 , \36265 );
nand \U$29166 ( \37118 , \37115 , \37116 , \37117 );
and \U$29167 ( \37119 , \37118 , \36691 );
or \U$29168 ( \37120 , \37113 , \37119 );
and \U$29170 ( \37121 , \37120 , 1'b1 );
or \U$29172 ( \37122 , \37121 , 1'b0 );
buf \U$29173 ( \37123 , \37122 );
_DC r23bfc_GF_IsGateDCbyConstraint ( \37124_nR23bfc , \37123 , \21944 );
buf \U$29174 ( \37125 , \37124_nR23bfc );
not \U$29175 ( \37126 , \32756 );
and \U$29176 ( \37127 , RIe3c2420_5941, \37126 );
not \U$29177 ( \37128 , RIe3c2420_5941);
or \U$29178 ( \37129 , \37128 , \36398 );
nand \U$29179 ( \37130 , \33899 , \36326 );
nand \U$29180 ( \37131 , \33902 , \36297 );
nand \U$29181 ( \37132 , \37129 , \37130 , \37131 );
and \U$29182 ( \37133 , \37132 , \32756 );
or \U$29183 ( \37134 , \37127 , \37133 );
and \U$29185 ( \37135 , \37134 , 1'b1 );
or \U$29187 ( \37136 , \37135 , 1'b0 );
buf \U$29188 ( \37137 , \37136 );
_DC r23bfe_GF_IsGateDCbyConstraint ( \37138_nR23bfe , \37137 , \21944 );
buf \U$29189 ( \37139 , \37138_nR23bfe );
not \U$29190 ( \37140 , \34318 );
and \U$29191 ( \37141 , RIe3c2c18_5942, \37140 );
not \U$29192 ( \37142 , RIe3c2c18_5942);
or \U$29193 ( \37143 , \37142 , \36310 );
nand \U$29194 ( \37144 , \33918 , \36280 );
nand \U$29195 ( \37145 , \33921 , \36342 );
nand \U$29196 ( \37146 , \37143 , \37144 , \37145 );
and \U$29197 ( \37147 , \37146 , \34318 );
or \U$29198 ( \37148 , \37141 , \37147 );
and \U$29200 ( \37149 , \37148 , 1'b1 );
or \U$29202 ( \37150 , \37149 , 1'b0 );
buf \U$29203 ( \37151 , \37150 );
_DC r23c00_GF_IsGateDCbyConstraint ( \37152_nR23c00 , \37151 , \21944 );
buf \U$29204 ( \37153 , \37152_nR23c00 );
not \U$29205 ( \37154 , \36691 );
and \U$29206 ( \37155 , RIe3c3410_5943, \37154 );
not \U$29207 ( \37156 , RIe3c3410_5943);
or \U$29208 ( \37157 , \37156 , \36294 );
nand \U$29209 ( \37158 , \33937 , \36280 );
nand \U$29210 ( \37159 , \33940 , \36297 );
nand \U$29211 ( \37160 , \37157 , \37158 , \37159 );
and \U$29212 ( \37161 , \37160 , \36691 );
or \U$29213 ( \37162 , \37155 , \37161 );
and \U$29215 ( \37163 , \37162 , 1'b1 );
or \U$29217 ( \37164 , \37163 , 1'b0 );
buf \U$29218 ( \37165 , \37164 );
_DC r23c02_GF_IsGateDCbyConstraint ( \37166_nR23c02 , \37165 , \21944 );
buf \U$29219 ( \37167 , \37166_nR23c02 );
or \U$29220 ( \37168 , \32657 , \32682 );
not \U$29221 ( \37169 , \37168 );
not \U$29222 ( \37170 , \37169 );
and \U$29223 ( \37171 , RIe202f10_5656, \37170 );
not \U$29224 ( \37172 , RIe202f10_5656);
not \U$29225 ( \37173 , \37172 );
not \U$29226 ( \37174 , \32676 );
and \U$29227 ( \37175 , \37173 , \37174 );
buf \U$29228 ( \37176 , RIb86fc68_77);
buf \U$29229 ( \37177 , \37176 );
and \U$29230 ( \37178 , \37177 , \32676 );
or \U$29231 ( \37179 , \37175 , \37178 );
and \U$29232 ( \37180 , \37179 , \37169 );
or \U$29233 ( \37181 , \37171 , \37180 );
and \U$29235 ( \37182 , \37181 , 1'b1 );
or \U$29237 ( \37183 , \37182 , 1'b0 );
buf \U$29238 ( \37184 , \37183 );
_DC r239cc_GF_IsGateDCbyConstraint ( \37185_nR239cc , \37184 , \21944 );
buf \U$29239 ( \37186 , \37185_nR239cc );
not \U$29240 ( \37187 , \37168 );
not \U$29241 ( \37188 , \37187 );
and \U$29242 ( \37189 , RIe202448_5657, \37188 );
not \U$29243 ( \37190 , RIe202448_5657);
not \U$29244 ( \37191 , \37190 );
not \U$29245 ( \37192 , \32676 );
and \U$29246 ( \37193 , \37191 , \37192 );
buf \U$29247 ( \37194 , RIb86fce0_76);
buf \U$29248 ( \37195 , \37194 );
and \U$29249 ( \37196 , \37195 , \32676 );
or \U$29250 ( \37197 , \37193 , \37196 );
and \U$29251 ( \37198 , \37197 , \37187 );
or \U$29252 ( \37199 , \37189 , \37198 );
and \U$29254 ( \37200 , \37199 , 1'b1 );
or \U$29256 ( \37201 , \37200 , 1'b0 );
buf \U$29257 ( \37202 , \37201 );
_DC r239ce_GF_IsGateDCbyConstraint ( \37203_nR239ce , \37202 , \21944 );
buf \U$29258 ( \37204 , \37203_nR239ce );
not \U$29259 ( \37205 , \37169 );
and \U$29260 ( \37206 , RIe201980_5658, \37205 );
not \U$29261 ( \37207 , RIe201980_5658);
not \U$29262 ( \37208 , \37207 );
not \U$29263 ( \37209 , \32676 );
and \U$29264 ( \37210 , \37208 , \37209 );
buf \U$29265 ( \37211 , \26703 );
and \U$29266 ( \37212 , \37211 , \32676 );
or \U$29267 ( \37213 , \37210 , \37212 );
and \U$29268 ( \37214 , \37213 , \37169 );
or \U$29269 ( \37215 , \37206 , \37214 );
and \U$29271 ( \37216 , \37215 , 1'b1 );
or \U$29273 ( \37217 , \37216 , 1'b0 );
buf \U$29274 ( \37218 , \37217 );
_DC r239d0_GF_IsGateDCbyConstraint ( \37219_nR239d0 , \37218 , \21944 );
buf \U$29275 ( \37220 , \37219_nR239d0 );
not \U$29276 ( \37221 , \37169 );
and \U$29277 ( \37222 , RIe200e40_5659, \37221 );
not \U$29278 ( \37223 , RIe200e40_5659);
not \U$29279 ( \37224 , \37223 );
not \U$29280 ( \37225 , \32676 );
and \U$29281 ( \37226 , \37224 , \37225 );
buf \U$29282 ( \37227 , RIb87e8a8_74);
buf \U$29283 ( \37228 , \37227 );
and \U$29284 ( \37229 , \37228 , \32676 );
or \U$29285 ( \37230 , \37226 , \37229 );
and \U$29286 ( \37231 , \37230 , \37169 );
or \U$29287 ( \37232 , \37222 , \37231 );
and \U$29289 ( \37233 , \37232 , 1'b1 );
or \U$29291 ( \37234 , \37233 , 1'b0 );
buf \U$29292 ( \37235 , \37234 );
_DC r239d2_GF_IsGateDCbyConstraint ( \37236_nR239d2 , \37235 , \21944 );
buf \U$29293 ( \37237 , \37236_nR239d2 );
not \U$29294 ( \37238 , \37169 );
and \U$29295 ( \37239 , RIe2000a8_5660, \37238 );
not \U$29296 ( \37240 , RIe2000a8_5660);
not \U$29297 ( \37241 , \37240 );
not \U$29298 ( \37242 , \32676 );
and \U$29299 ( \37243 , \37241 , \37242 );
buf \U$29300 ( \37244 , RIb87e920_73);
buf \U$29301 ( \37245 , \37244 );
and \U$29302 ( \37246 , \37245 , \32676 );
or \U$29303 ( \37247 , \37243 , \37246 );
and \U$29304 ( \37248 , \37247 , \37169 );
or \U$29305 ( \37249 , \37239 , \37248 );
and \U$29307 ( \37250 , \37249 , 1'b1 );
or \U$29309 ( \37251 , \37250 , 1'b0 );
buf \U$29310 ( \37252 , \37251 );
_DC r239d4_GF_IsGateDCbyConstraint ( \37253_nR239d4 , \37252 , \21944 );
buf \U$29311 ( \37254 , \37253_nR239d4 );
not \U$29312 ( \37255 , \37187 );
and \U$29313 ( \37256 , RIe1ff310_5661, \37255 );
not \U$29314 ( \37257 , RIe1ff310_5661);
not \U$29315 ( \37258 , \37257 );
not \U$29316 ( \37259 , \32676 );
and \U$29317 ( \37260 , \37258 , \37259 );
buf \U$29318 ( \37261 , RIb87e998_72);
buf \U$29319 ( \37262 , \37261 );
and \U$29320 ( \37263 , \37262 , \32676 );
or \U$29321 ( \37264 , \37260 , \37263 );
and \U$29322 ( \37265 , \37264 , \37187 );
or \U$29323 ( \37266 , \37256 , \37265 );
and \U$29325 ( \37267 , \37266 , 1'b1 );
or \U$29327 ( \37268 , \37267 , 1'b0 );
buf \U$29328 ( \37269 , \37268 );
_DC r239d6_GF_IsGateDCbyConstraint ( \37270_nR239d6 , \37269 , \21944 );
buf \U$29329 ( \37271 , \37270_nR239d6 );
not \U$29330 ( \37272 , \37169 );
and \U$29331 ( \37273 , RIe1fe668_5662, \37272 );
not \U$29332 ( \37274 , RIe1fe668_5662);
not \U$29333 ( \37275 , \37274 );
not \U$29334 ( \37276 , \32676 );
and \U$29335 ( \37277 , \37275 , \37276 );
buf \U$29336 ( \37278 , RIb87ea10_71);
buf \U$29337 ( \37279 , \37278 );
and \U$29338 ( \37280 , \37279 , \32676 );
or \U$29339 ( \37281 , \37277 , \37280 );
and \U$29340 ( \37282 , \37281 , \37169 );
or \U$29341 ( \37283 , \37273 , \37282 );
and \U$29343 ( \37284 , \37283 , 1'b1 );
or \U$29345 ( \37285 , \37284 , 1'b0 );
buf \U$29346 ( \37286 , \37285 );
_DC r239d8_GF_IsGateDCbyConstraint ( \37287_nR239d8 , \37286 , \21944 );
buf \U$29347 ( \37288 , \37287_nR239d8 );
not \U$29348 ( \37289 , \37187 );
and \U$29349 ( \37290 , RIe1fd9c0_5663, \37289 );
not \U$29350 ( \37291 , RIe1fd9c0_5663);
not \U$29351 ( \37292 , \37291 );
not \U$29352 ( \37293 , \32676 );
and \U$29353 ( \37294 , \37292 , \37293 );
buf \U$29354 ( \37295 , RIb87ea88_70);
buf \U$29355 ( \37296 , \37295 );
and \U$29356 ( \37297 , \37296 , \32676 );
or \U$29357 ( \37298 , \37294 , \37297 );
and \U$29358 ( \37299 , \37298 , \37187 );
or \U$29359 ( \37300 , \37290 , \37299 );
and \U$29361 ( \37301 , \37300 , 1'b1 );
or \U$29363 ( \37302 , \37301 , 1'b0 );
buf \U$29364 ( \37303 , \37302 );
_DC r239da_GF_IsGateDCbyConstraint ( \37304_nR239da , \37303 , \21944 );
buf \U$29365 ( \37305 , \37304_nR239da );
not \U$29366 ( \37306 , \37169 );
and \U$29367 ( \37307 , RIe1fce80_5664, \37306 );
not \U$29368 ( \37308 , RIe1fce80_5664);
not \U$29369 ( \37309 , \37308 );
not \U$29370 ( \37310 , \33961 );
and \U$29371 ( \37311 , \37309 , \37310 );
and \U$29372 ( \37312 , \37177 , \33961 );
or \U$29373 ( \37313 , \37311 , \37312 );
and \U$29374 ( \37314 , \37313 , \37169 );
or \U$29375 ( \37315 , \37307 , \37314 );
and \U$29377 ( \37316 , \37315 , 1'b1 );
or \U$29379 ( \37317 , \37316 , 1'b0 );
buf \U$29380 ( \37318 , \37317 );
_DC r239dc_GF_IsGateDCbyConstraint ( \37319_nR239dc , \37318 , \21944 );
buf \U$29381 ( \37320 , \37319_nR239dc );
not \U$29382 ( \37321 , \37187 );
and \U$29383 ( \37322 , RIe1fc340_5665, \37321 );
not \U$29384 ( \37323 , RIe1fc340_5665);
not \U$29385 ( \37324 , \37323 );
not \U$29386 ( \37325 , \33961 );
and \U$29387 ( \37326 , \37324 , \37325 );
and \U$29388 ( \37327 , \37195 , \33961 );
or \U$29389 ( \37328 , \37326 , \37327 );
and \U$29390 ( \37329 , \37328 , \37187 );
or \U$29391 ( \37330 , \37322 , \37329 );
and \U$29393 ( \37331 , \37330 , 1'b1 );
or \U$29395 ( \37332 , \37331 , 1'b0 );
buf \U$29396 ( \37333 , \37332 );
_DC r239de_GF_IsGateDCbyConstraint ( \37334_nR239de , \37333 , \21944 );
buf \U$29397 ( \37335 , \37334_nR239de );
not \U$29398 ( \37336 , \37169 );
and \U$29399 ( \37337 , RIe1fb878_5666, \37336 );
not \U$29400 ( \37338 , RIe1fb878_5666);
not \U$29401 ( \37339 , \37338 );
not \U$29402 ( \37340 , \33961 );
and \U$29403 ( \37341 , \37339 , \37340 );
and \U$29404 ( \37342 , \37211 , \33961 );
or \U$29405 ( \37343 , \37341 , \37342 );
and \U$29406 ( \37344 , \37343 , \37169 );
or \U$29407 ( \37345 , \37337 , \37344 );
and \U$29409 ( \37346 , \37345 , 1'b1 );
or \U$29411 ( \37347 , \37346 , 1'b0 );
buf \U$29412 ( \37348 , \37347 );
_DC r239e0_GF_IsGateDCbyConstraint ( \37349_nR239e0 , \37348 , \21944 );
buf \U$29413 ( \37350 , \37349_nR239e0 );
not \U$29414 ( \37351 , \37187 );
and \U$29415 ( \37352 , RIe1facc0_5667, \37351 );
not \U$29416 ( \37353 , RIe1facc0_5667);
not \U$29417 ( \37354 , \37353 );
not \U$29418 ( \37355 , \33961 );
and \U$29419 ( \37356 , \37354 , \37355 );
and \U$29420 ( \37357 , \37228 , \33961 );
or \U$29421 ( \37358 , \37356 , \37357 );
and \U$29422 ( \37359 , \37358 , \37187 );
or \U$29423 ( \37360 , \37352 , \37359 );
and \U$29425 ( \37361 , \37360 , 1'b1 );
or \U$29427 ( \37362 , \37361 , 1'b0 );
buf \U$29428 ( \37363 , \37362 );
_DC r239e2_GF_IsGateDCbyConstraint ( \37364_nR239e2 , \37363 , \21944 );
buf \U$29429 ( \37365 , \37364_nR239e2 );
not \U$29430 ( \37366 , \37169 );
and \U$29431 ( \37367 , RIe1fa090_5668, \37366 );
not \U$29432 ( \37368 , RIe1fa090_5668);
not \U$29433 ( \37369 , \37368 );
not \U$29434 ( \37370 , \33961 );
and \U$29435 ( \37371 , \37369 , \37370 );
and \U$29436 ( \37372 , \37245 , \33961 );
or \U$29437 ( \37373 , \37371 , \37372 );
and \U$29438 ( \37374 , \37373 , \37169 );
or \U$29439 ( \37375 , \37367 , \37374 );
and \U$29441 ( \37376 , \37375 , 1'b1 );
or \U$29443 ( \37377 , \37376 , 1'b0 );
buf \U$29444 ( \37378 , \37377 );
_DC r239e4_GF_IsGateDCbyConstraint ( \37379_nR239e4 , \37378 , \21944 );
buf \U$29445 ( \37380 , \37379_nR239e4 );
not \U$29446 ( \37381 , \37187 );
and \U$29447 ( \37382 , RIe1f9118_5669, \37381 );
not \U$29448 ( \37383 , RIe1f9118_5669);
not \U$29449 ( \37384 , \37383 );
not \U$29450 ( \37385 , \33961 );
and \U$29451 ( \37386 , \37384 , \37385 );
and \U$29452 ( \37387 , \37262 , \33961 );
or \U$29453 ( \37388 , \37386 , \37387 );
and \U$29454 ( \37389 , \37388 , \37187 );
or \U$29455 ( \37390 , \37382 , \37389 );
and \U$29457 ( \37391 , \37390 , 1'b1 );
or \U$29459 ( \37392 , \37391 , 1'b0 );
buf \U$29460 ( \37393 , \37392 );
_DC r239e6_GF_IsGateDCbyConstraint ( \37394_nR239e6 , \37393 , \21944 );
buf \U$29461 ( \37395 , \37394_nR239e6 );
not \U$29462 ( \37396 , \37169 );
and \U$29463 ( \37397 , RIe1f7fc0_5670, \37396 );
not \U$29464 ( \37398 , RIe1f7fc0_5670);
not \U$29465 ( \37399 , \37398 );
not \U$29466 ( \37400 , \33961 );
and \U$29467 ( \37401 , \37399 , \37400 );
and \U$29468 ( \37402 , \37279 , \33961 );
or \U$29469 ( \37403 , \37401 , \37402 );
and \U$29470 ( \37404 , \37403 , \37169 );
or \U$29471 ( \37405 , \37397 , \37404 );
and \U$29473 ( \37406 , \37405 , 1'b1 );
or \U$29475 ( \37407 , \37406 , 1'b0 );
buf \U$29476 ( \37408 , \37407 );
_DC r239e8_GF_IsGateDCbyConstraint ( \37409_nR239e8 , \37408 , \21944 );
buf \U$29477 ( \37410 , \37409_nR239e8 );
not \U$29478 ( \37411 , \37187 );
and \U$29479 ( \37412 , RIe1f69b8_5671, \37411 );
not \U$29480 ( \37413 , RIe1f69b8_5671);
not \U$29481 ( \37414 , \37413 );
not \U$29482 ( \37415 , \33961 );
and \U$29483 ( \37416 , \37414 , \37415 );
and \U$29484 ( \37417 , \37296 , \33961 );
or \U$29485 ( \37418 , \37416 , \37417 );
and \U$29486 ( \37419 , \37418 , \37187 );
or \U$29487 ( \37420 , \37412 , \37419 );
and \U$29489 ( \37421 , \37420 , 1'b1 );
or \U$29491 ( \37422 , \37421 , 1'b0 );
buf \U$29492 ( \37423 , \37422 );
_DC r239ea_GF_IsGateDCbyConstraint ( \37424_nR239ea , \37423 , \21944 );
buf \U$29493 ( \37425 , \37424_nR239ea );
not \U$29494 ( \37426 , \37169 );
and \U$29495 ( \37427 , RIe1f5860_5672, \37426 );
not \U$29496 ( \37428 , RIe1f5860_5672);
not \U$29497 ( \37429 , \37428 );
not \U$29498 ( \37430 , \35142 );
and \U$29499 ( \37431 , \37429 , \37430 );
and \U$29500 ( \37432 , \37177 , \35142 );
or \U$29501 ( \37433 , \37431 , \37432 );
and \U$29502 ( \37434 , \37433 , \37169 );
or \U$29503 ( \37435 , \37427 , \37434 );
and \U$29505 ( \37436 , \37435 , 1'b1 );
or \U$29507 ( \37437 , \37436 , 1'b0 );
buf \U$29508 ( \37438 , \37437 );
_DC r239ec_GF_IsGateDCbyConstraint ( \37439_nR239ec , \37438 , \21944 );
buf \U$29509 ( \37440 , \37439_nR239ec );
not \U$29510 ( \37441 , \37169 );
and \U$29511 ( \37442 , RIe1f4258_5673, \37441 );
not \U$29512 ( \37443 , RIe1f4258_5673);
not \U$29513 ( \37444 , \37443 );
not \U$29514 ( \37445 , \35142 );
and \U$29515 ( \37446 , \37444 , \37445 );
and \U$29516 ( \37447 , \37195 , \35142 );
or \U$29517 ( \37448 , \37446 , \37447 );
and \U$29518 ( \37449 , \37448 , \37169 );
or \U$29519 ( \37450 , \37442 , \37449 );
and \U$29521 ( \37451 , \37450 , 1'b1 );
or \U$29523 ( \37452 , \37451 , 1'b0 );
buf \U$29524 ( \37453 , \37452 );
_DC r239ee_GF_IsGateDCbyConstraint ( \37454_nR239ee , \37453 , \21944 );
buf \U$29525 ( \37455 , \37454_nR239ee );
not \U$29526 ( \37456 , \37169 );
and \U$29527 ( \37457 , RIe1f3100_5674, \37456 );
not \U$29528 ( \37458 , RIe1f3100_5674);
not \U$29529 ( \37459 , \37458 );
not \U$29530 ( \37460 , \35142 );
and \U$29531 ( \37461 , \37459 , \37460 );
and \U$29532 ( \37462 , \37211 , \35142 );
or \U$29533 ( \37463 , \37461 , \37462 );
and \U$29534 ( \37464 , \37463 , \37169 );
or \U$29535 ( \37465 , \37457 , \37464 );
and \U$29537 ( \37466 , \37465 , 1'b1 );
or \U$29539 ( \37467 , \37466 , 1'b0 );
buf \U$29540 ( \37468 , \37467 );
_DC r239f0_GF_IsGateDCbyConstraint ( \37469_nR239f0 , \37468 , \21944 );
buf \U$29541 ( \37470 , \37469_nR239f0 );
not \U$29542 ( \37471 , \37169 );
and \U$29543 ( \37472 , RIe1f1fa8_5675, \37471 );
not \U$29544 ( \37473 , RIe1f1fa8_5675);
not \U$29545 ( \37474 , \37473 );
not \U$29546 ( \37475 , \35142 );
and \U$29547 ( \37476 , \37474 , \37475 );
and \U$29548 ( \37477 , \37228 , \35142 );
or \U$29549 ( \37478 , \37476 , \37477 );
and \U$29550 ( \37479 , \37478 , \37169 );
or \U$29551 ( \37480 , \37472 , \37479 );
and \U$29553 ( \37481 , \37480 , 1'b1 );
or \U$29555 ( \37482 , \37481 , 1'b0 );
buf \U$29556 ( \37483 , \37482 );
_DC r239f2_GF_IsGateDCbyConstraint ( \37484_nR239f2 , \37483 , \21944 );
buf \U$29557 ( \37485 , \37484_nR239f2 );
not \U$29558 ( \37486 , \37169 );
and \U$29559 ( \37487 , RIe1f09a0_5676, \37486 );
not \U$29560 ( \37488 , RIe1f09a0_5676);
not \U$29561 ( \37489 , \37488 );
not \U$29562 ( \37490 , \35142 );
and \U$29563 ( \37491 , \37489 , \37490 );
and \U$29564 ( \37492 , \37245 , \35142 );
or \U$29565 ( \37493 , \37491 , \37492 );
and \U$29566 ( \37494 , \37493 , \37169 );
or \U$29567 ( \37495 , \37487 , \37494 );
and \U$29569 ( \37496 , \37495 , 1'b1 );
or \U$29571 ( \37497 , \37496 , 1'b0 );
buf \U$29572 ( \37498 , \37497 );
_DC r239f4_GF_IsGateDCbyConstraint ( \37499_nR239f4 , \37498 , \21944 );
buf \U$29573 ( \37500 , \37499_nR239f4 );
not \U$29574 ( \37501 , \37169 );
and \U$29575 ( \37502 , RIe1ef848_5677, \37501 );
not \U$29576 ( \37503 , RIe1ef848_5677);
not \U$29577 ( \37504 , \37503 );
not \U$29578 ( \37505 , \35142 );
and \U$29579 ( \37506 , \37504 , \37505 );
and \U$29580 ( \37507 , \37262 , \35142 );
or \U$29581 ( \37508 , \37506 , \37507 );
and \U$29582 ( \37509 , \37508 , \37169 );
or \U$29583 ( \37510 , \37502 , \37509 );
and \U$29585 ( \37511 , \37510 , 1'b1 );
or \U$29587 ( \37512 , \37511 , 1'b0 );
buf \U$29588 ( \37513 , \37512 );
_DC r239f6_GF_IsGateDCbyConstraint ( \37514_nR239f6 , \37513 , \21944 );
buf \U$29589 ( \37515 , \37514_nR239f6 );
not \U$29590 ( \37516 , \37169 );
and \U$29591 ( \37517 , RIe1ee240_5678, \37516 );
not \U$29592 ( \37518 , RIe1ee240_5678);
not \U$29593 ( \37519 , \37518 );
not \U$29594 ( \37520 , \35142 );
and \U$29595 ( \37521 , \37519 , \37520 );
and \U$29596 ( \37522 , \37279 , \35142 );
or \U$29597 ( \37523 , \37521 , \37522 );
and \U$29598 ( \37524 , \37523 , \37169 );
or \U$29599 ( \37525 , \37517 , \37524 );
and \U$29601 ( \37526 , \37525 , 1'b1 );
or \U$29603 ( \37527 , \37526 , 1'b0 );
buf \U$29604 ( \37528 , \37527 );
_DC r239f8_GF_IsGateDCbyConstraint ( \37529_nR239f8 , \37528 , \21944 );
buf \U$29605 ( \37530 , \37529_nR239f8 );
not \U$29606 ( \37531 , \37169 );
and \U$29607 ( \37532 , RIe1ed0e8_5679, \37531 );
not \U$29608 ( \37533 , RIe1ed0e8_5679);
not \U$29609 ( \37534 , \37533 );
not \U$29610 ( \37535 , \35142 );
and \U$29611 ( \37536 , \37534 , \37535 );
and \U$29612 ( \37537 , \37296 , \35142 );
or \U$29613 ( \37538 , \37536 , \37537 );
and \U$29614 ( \37539 , \37538 , \37169 );
or \U$29615 ( \37540 , \37532 , \37539 );
and \U$29617 ( \37541 , \37540 , 1'b1 );
or \U$29619 ( \37542 , \37541 , 1'b0 );
buf \U$29620 ( \37543 , \37542 );
_DC r239fa_GF_IsGateDCbyConstraint ( \37544_nR239fa , \37543 , \21944 );
buf \U$29621 ( \37545 , \37544_nR239fa );
not \U$29622 ( \37546 , \37169 );
and \U$29623 ( \37547 , RIe1ebae0_5680, \37546 );
not \U$29624 ( \37548 , RIe1ebae0_5680);
not \U$29625 ( \37549 , \37548 );
not \U$29626 ( \37550 , \36252 );
and \U$29627 ( \37551 , \37549 , \37550 );
and \U$29628 ( \37552 , \37177 , \36252 );
or \U$29629 ( \37553 , \37551 , \37552 );
and \U$29630 ( \37554 , \37553 , \37169 );
or \U$29631 ( \37555 , \37547 , \37554 );
and \U$29633 ( \37556 , \37555 , 1'b1 );
or \U$29635 ( \37557 , \37556 , 1'b0 );
buf \U$29636 ( \37558 , \37557 );
_DC r239fc_GF_IsGateDCbyConstraint ( \37559_nR239fc , \37558 , \21944 );
buf \U$29637 ( \37560 , \37559_nR239fc );
not \U$29638 ( \37561 , \37187 );
and \U$29639 ( \37562 , RIe1ea988_5681, \37561 );
not \U$29640 ( \37563 , RIe1ea988_5681);
not \U$29641 ( \37564 , \37563 );
not \U$29642 ( \37565 , \36252 );
and \U$29643 ( \37566 , \37564 , \37565 );
and \U$29644 ( \37567 , \37195 , \36252 );
or \U$29645 ( \37568 , \37566 , \37567 );
and \U$29646 ( \37569 , \37568 , \37187 );
or \U$29647 ( \37570 , \37562 , \37569 );
and \U$29649 ( \37571 , \37570 , 1'b1 );
or \U$29651 ( \37572 , \37571 , 1'b0 );
buf \U$29652 ( \37573 , \37572 );
_DC r239fe_GF_IsGateDCbyConstraint ( \37574_nR239fe , \37573 , \21944 );
buf \U$29653 ( \37575 , \37574_nR239fe );
not \U$29654 ( \37576 , \37187 );
and \U$29655 ( \37577 , RIe1e9830_5682, \37576 );
not \U$29656 ( \37578 , RIe1e9830_5682);
not \U$29657 ( \37579 , \37578 );
not \U$29658 ( \37580 , \36252 );
and \U$29659 ( \37581 , \37579 , \37580 );
and \U$29660 ( \37582 , \37211 , \36252 );
or \U$29661 ( \37583 , \37581 , \37582 );
and \U$29662 ( \37584 , \37583 , \37187 );
or \U$29663 ( \37585 , \37577 , \37584 );
and \U$29665 ( \37586 , \37585 , 1'b1 );
or \U$29667 ( \37587 , \37586 , 1'b0 );
buf \U$29668 ( \37588 , \37587 );
_DC r23a00_GF_IsGateDCbyConstraint ( \37589_nR23a00 , \37588 , \21944 );
buf \U$29669 ( \37590 , \37589_nR23a00 );
not \U$29670 ( \37591 , \37187 );
and \U$29671 ( \37592 , RIe1e8228_5683, \37591 );
not \U$29672 ( \37593 , RIe1e8228_5683);
not \U$29673 ( \37594 , \37593 );
not \U$29674 ( \37595 , \36252 );
and \U$29675 ( \37596 , \37594 , \37595 );
and \U$29676 ( \37597 , \37228 , \36252 );
or \U$29677 ( \37598 , \37596 , \37597 );
and \U$29678 ( \37599 , \37598 , \37187 );
or \U$29679 ( \37600 , \37592 , \37599 );
and \U$29681 ( \37601 , \37600 , 1'b1 );
or \U$29683 ( \37602 , \37601 , 1'b0 );
buf \U$29684 ( \37603 , \37602 );
_DC r23a02_GF_IsGateDCbyConstraint ( \37604_nR23a02 , \37603 , \21944 );
buf \U$29685 ( \37605 , \37604_nR23a02 );
not \U$29686 ( \37606 , \37187 );
and \U$29687 ( \37607 , RIe1e70d0_5684, \37606 );
not \U$29688 ( \37608 , RIe1e70d0_5684);
not \U$29689 ( \37609 , \37608 );
not \U$29690 ( \37610 , \36252 );
and \U$29691 ( \37611 , \37609 , \37610 );
and \U$29692 ( \37612 , \37245 , \36252 );
or \U$29693 ( \37613 , \37611 , \37612 );
and \U$29694 ( \37614 , \37613 , \37187 );
or \U$29695 ( \37615 , \37607 , \37614 );
and \U$29697 ( \37616 , \37615 , 1'b1 );
or \U$29699 ( \37617 , \37616 , 1'b0 );
buf \U$29700 ( \37618 , \37617 );
_DC r23a04_GF_IsGateDCbyConstraint ( \37619_nR23a04 , \37618 , \21944 );
buf \U$29701 ( \37620 , \37619_nR23a04 );
not \U$29702 ( \37621 , \37187 );
and \U$29703 ( \37622 , RIe1e5ac8_5685, \37621 );
not \U$29704 ( \37623 , RIe1e5ac8_5685);
not \U$29705 ( \37624 , \37623 );
not \U$29706 ( \37625 , \36252 );
and \U$29707 ( \37626 , \37624 , \37625 );
and \U$29708 ( \37627 , \37262 , \36252 );
or \U$29709 ( \37628 , \37626 , \37627 );
and \U$29710 ( \37629 , \37628 , \37187 );
or \U$29711 ( \37630 , \37622 , \37629 );
and \U$29713 ( \37631 , \37630 , 1'b1 );
or \U$29715 ( \37632 , \37631 , 1'b0 );
buf \U$29716 ( \37633 , \37632 );
_DC r23a06_GF_IsGateDCbyConstraint ( \37634_nR23a06 , \37633 , \21944 );
buf \U$29717 ( \37635 , \37634_nR23a06 );
not \U$29718 ( \37636 , \37187 );
and \U$29719 ( \37637 , RIe1e4970_5686, \37636 );
not \U$29720 ( \37638 , RIe1e4970_5686);
not \U$29721 ( \37639 , \37638 );
not \U$29722 ( \37640 , \36252 );
and \U$29723 ( \37641 , \37639 , \37640 );
and \U$29724 ( \37642 , \37279 , \36252 );
or \U$29725 ( \37643 , \37641 , \37642 );
and \U$29726 ( \37644 , \37643 , \37187 );
or \U$29727 ( \37645 , \37637 , \37644 );
and \U$29729 ( \37646 , \37645 , 1'b1 );
or \U$29731 ( \37647 , \37646 , 1'b0 );
buf \U$29732 ( \37648 , \37647 );
_DC r23a08_GF_IsGateDCbyConstraint ( \37649_nR23a08 , \37648 , \21944 );
buf \U$29733 ( \37650 , \37649_nR23a08 );
not \U$29734 ( \37651 , \37169 );
and \U$29735 ( \37652 , RIe1e3368_5687, \37651 );
not \U$29736 ( \37653 , RIe1e3368_5687);
not \U$29737 ( \37654 , \37653 );
not \U$29738 ( \37655 , \36252 );
and \U$29739 ( \37656 , \37654 , \37655 );
and \U$29740 ( \37657 , \37296 , \36252 );
or \U$29741 ( \37658 , \37656 , \37657 );
and \U$29742 ( \37659 , \37658 , \37169 );
or \U$29743 ( \37660 , \37652 , \37659 );
and \U$29745 ( \37661 , \37660 , 1'b1 );
or \U$29747 ( \37662 , \37661 , 1'b0 );
buf \U$29748 ( \37663 , \37662 );
_DC r23a0a_GF_IsGateDCbyConstraint ( \37664_nR23a0a , \37663 , \21944 );
buf \U$29749 ( \37665 , \37664_nR23a0a );
buf \U$29750 ( \37666 , RIb7b9680_245);
buf \U$29751 ( \37667 , RIb79b3b0_273);
nand \U$29752 ( \37668 , \37667 , \32662 );
not \U$29753 ( \37669 , \37668 );
and \U$29754 ( \37670 , \37666 , \37669 );
and \U$29755 ( \37671 , RIe4520c0_5970, \37668 );
or \U$29756 ( \37672 , \37670 , \37671 );
and \U$29758 ( \37673 , \37672 , 1'b1 );
or \U$29760 ( \37674 , \37673 , 1'b0 );
buf \U$29761 ( \37675 , \37674 );
_DC r23c24_GF_IsGateDCbyConstraint ( \37676_nR23c24 , \37675 , \21944 );
buf \U$29762 ( \37677 , \37676_nR23c24 );
not \U$29763 ( \37678 , \37668 );
not \U$29764 ( \37679 , \37678 );
and \U$29765 ( \37680 , RIe438440_5990, \37679 );
buf \U$29766 ( \37681 , RIb7b96f8_244);
and \U$29767 ( \37682 , \37681 , \37678 );
or \U$29768 ( \37683 , \37680 , \37682 );
and \U$29770 ( \37684 , \37683 , 1'b1 );
or \U$29772 ( \37685 , \37684 , 1'b0 );
buf \U$29773 ( \37686 , \37685 );
_DC r23c26_GF_IsGateDCbyConstraint ( \37687_nR23c26 , \37686 , \21944 );
buf \U$29774 ( \37688 , \37687_nR23c26 );
not \U$29775 ( \37689 , \37678 );
and \U$29776 ( \37690 , RIe4390e8_5989, \37689 );
buf \U$29777 ( \37691 , RIb7c20c8_243);
and \U$29778 ( \37692 , \37691 , \37678 );
or \U$29779 ( \37693 , \37690 , \37692 );
and \U$29781 ( \37694 , \37693 , 1'b1 );
or \U$29783 ( \37695 , \37694 , 1'b0 );
buf \U$29784 ( \37696 , \37695 );
_DC r23c28_GF_IsGateDCbyConstraint ( \37697_nR23c28 , \37696 , \21944 );
buf \U$29785 ( \37698 , \37697_nR23c28 );
not \U$29786 ( \37699 , \37678 );
and \U$29787 ( \37700 , RIe439f70_5988, \37699 );
buf \U$29788 ( \37701 , RIb7c5728_242);
and \U$29789 ( \37702 , \37701 , \37678 );
or \U$29790 ( \37703 , \37700 , \37702 );
and \U$29792 ( \37704 , \37703 , 1'b1 );
or \U$29794 ( \37705 , \37704 , 1'b0 );
buf \U$29795 ( \37706 , \37705 );
_DC r23c2a_GF_IsGateDCbyConstraint ( \37707_nR23c2a , \37706 , \21944 );
buf \U$29796 ( \37708 , \37707_nR23c2a );
not \U$29797 ( \37709 , \37678 );
and \U$29798 ( \37710 , RIe43ad80_5987, \37709 );
buf \U$29799 ( \37711 , RIb7c57a0_241);
and \U$29800 ( \37712 , \37711 , \37678 );
or \U$29801 ( \37713 , \37710 , \37712 );
and \U$29803 ( \37714 , \37713 , 1'b1 );
or \U$29805 ( \37715 , \37714 , 1'b0 );
buf \U$29806 ( \37716 , \37715 );
_DC r23c2c_GF_IsGateDCbyConstraint ( \37717_nR23c2c , \37716 , \21944 );
buf \U$29807 ( \37718 , \37717_nR23c2c );
not \U$29808 ( \37719 , \37678 );
and \U$29809 ( \37720 , RIe43ba28_5986, \37719 );
buf \U$29810 ( \37721 , RIb7c5818_240);
and \U$29811 ( \37722 , \37721 , \37678 );
or \U$29812 ( \37723 , \37720 , \37722 );
and \U$29814 ( \37724 , \37723 , 1'b1 );
or \U$29816 ( \37725 , \37724 , 1'b0 );
buf \U$29817 ( \37726 , \37725 );
_DC r23c2e_GF_IsGateDCbyConstraint ( \37727_nR23c2e , \37726 , \21944 );
buf \U$29818 ( \37728 , \37727_nR23c2e );
not \U$29819 ( \37729 , \37678 );
and \U$29820 ( \37730 , RIe43c7c0_5985, \37729 );
buf \U$29821 ( \37731 , RIb7c5890_239);
and \U$29822 ( \37732 , \37731 , \37678 );
or \U$29823 ( \37733 , \37730 , \37732 );
and \U$29825 ( \37734 , \37733 , 1'b1 );
or \U$29827 ( \37735 , \37734 , 1'b0 );
buf \U$29828 ( \37736 , \37735 );
_DC r23c30_GF_IsGateDCbyConstraint ( \37737_nR23c30 , \37736 , \21944 );
buf \U$29829 ( \37738 , \37737_nR23c30 );
not \U$29830 ( \37739 , \37678 );
and \U$29831 ( \37740 , RIe43d5d0_5984, \37739 );
buf \U$29832 ( \37741 , RIb7c5908_238);
and \U$29833 ( \37742 , \37741 , \37678 );
or \U$29834 ( \37743 , \37740 , \37742 );
and \U$29836 ( \37744 , \37743 , 1'b1 );
or \U$29838 ( \37745 , \37744 , 1'b0 );
buf \U$29839 ( \37746 , \37745 );
_DC r23c32_GF_IsGateDCbyConstraint ( \37747_nR23c32 , \37746 , \21944 );
buf \U$29840 ( \37748 , \37747_nR23c32 );
not \U$29841 ( \37749 , \37678 );
and \U$29842 ( \37750 , RIe445e38_5974, \37749 );
buf \U$29843 ( \37751 , RIb7a09f0_266);
and \U$29844 ( \37752 , \37751 , \37678 );
or \U$29845 ( \37753 , \37750 , \37752 );
and \U$29847 ( \37754 , \37753 , 1'b1 );
or \U$29849 ( \37755 , \37754 , 1'b0 );
buf \U$29850 ( \37756 , \37755 );
_DC r23c22_GF_IsGateDCbyConstraint ( \37757_nR23c22 , \37756 , \21944 );
buf \U$29851 ( \37758 , \37757_nR23c22 );
not \U$29852 ( \37759 , \37678 );
and \U$29853 ( \37760 , RIe441c98_5979, \37759 );
buf \U$29854 ( \37761 , RIb7a0a68_265);
and \U$29855 ( \37762 , \37761 , \37678 );
or \U$29856 ( \37763 , \37760 , \37762 );
and \U$29858 ( \37764 , \37763 , 1'b1 );
or \U$29860 ( \37765 , \37764 , 1'b0 );
buf \U$29861 ( \37766 , \37765 );
_DC r23c34_GF_IsGateDCbyConstraint ( \37767_nR23c34 , \37766 , \21944 );
buf \U$29862 ( \37768 , \37767_nR23c34 );
not \U$29863 ( \37769 , \37678 );
and \U$29864 ( \37770 , RIe4429b8_5978, \37769 );
buf \U$29865 ( \37771 , RIb7a0ae0_264);
and \U$29866 ( \37772 , \37771 , \37678 );
or \U$29867 ( \37773 , \37770 , \37772 );
and \U$29869 ( \37774 , \37773 , 1'b1 );
or \U$29871 ( \37775 , \37774 , 1'b0 );
buf \U$29872 ( \37776 , \37775 );
_DC r23c36_GF_IsGateDCbyConstraint ( \37777_nR23c36 , \37776 , \21944 );
buf \U$29873 ( \37778 , \37777_nR23c36 );
not \U$29874 ( \37779 , \37678 );
and \U$29875 ( \37780 , RIe443750_5977, \37779 );
buf \U$29876 ( \37781 , RIb7a0b58_263);
and \U$29877 ( \37782 , \37781 , \37678 );
or \U$29878 ( \37783 , \37780 , \37782 );
and \U$29880 ( \37784 , \37783 , 1'b1 );
or \U$29882 ( \37785 , \37784 , 1'b0 );
buf \U$29883 ( \37786 , \37785 );
_DC r23c38_GF_IsGateDCbyConstraint ( \37787_nR23c38 , \37786 , \21944 );
buf \U$29884 ( \37788 , \37787_nR23c38 );
not \U$29885 ( \37789 , \37678 );
and \U$29886 ( \37790 , RIe437630_5991, \37789 );
buf \U$29887 ( \37791 , RIb7a0bd0_262);
and \U$29888 ( \37792 , \37791 , \37678 );
or \U$29889 ( \37793 , \37790 , \37792 );
and \U$29891 ( \37794 , \37793 , 1'b1 );
or \U$29893 ( \37795 , \37794 , 1'b0 );
buf \U$29894 ( \37796 , \37795 );
_DC r23c3a_GF_IsGateDCbyConstraint ( \37797_nR23c3a , \37796 , \21944 );
buf \U$29895 ( \37798 , \37797_nR23c3a );
buf \U$29896 ( \37799 , RIb839668_156);
buf \U$29897 ( \37800 , \37799 );
not \U$29898 ( \37801 , \37800 );
not \U$29899 ( \37802 , \37801 );
buf \U$29900 ( \37803 , RIb839848_152);
and \U$29901 ( \37804 , \37803 , \32652 );
buf \U$29902 ( \37805 , RIb8396e0_155);
nand \U$29903 ( \37806 , \37805 , \32652 );
not \U$29904 ( \37807 , \37806 );
buf \U$29905 ( \37808 , \37807 );
or \U$29906 ( \37809 , \37802 , \37804 , \37808 );
nand \U$29907 ( \37810 , \37809 , \32652 );
not \U$29908 ( \37811 , \37810 );
not \U$29909 ( \37812 , RIe455e28_5964);
or \U$29910 ( \37813 , \37811 , \37812 );
nand \U$29911 ( \37814 , \37806 , \37801 );
not \U$29912 ( \37815 , RIe4554c8_5965);
not \U$29913 ( \37816 , \37815 );
or \U$29914 ( \37817 , \37812 , \37816 );
not \U$29915 ( \37818 , \37817 );
nand \U$29916 ( \37819 , RIe454988_5966, \37818 );
or \U$29917 ( \37820 , \37814 , \37819 );
xor \U$29918 ( \37821 , \37812 , \37815 );
nor \U$29919 ( \37822 , \37821 , \37818 );
nand \U$29920 ( \37823 , \32652 , \37806 , \37800 );
or \U$29921 ( \37824 , \37822 , \37823 );
not \U$29922 ( \37825 , \37814 );
nand \U$29923 ( \37826 , \37804 , \37819 , \37825 );
not \U$29924 ( \37827 , RIe454988_5966);
nor \U$29925 ( \37828 , \37815 , \37827 );
xor \U$29926 ( \37829 , \37812 , \37828 );
or \U$29927 ( \37830 , \37826 , \37829 );
nand \U$29928 ( \37831 , \37813 , \37820 , \37824 , \37830 );
not \U$29929 ( \37832 , RIe45c278_5954);
not \U$29930 ( \37833 , RIe45cdb8_5953);
not \U$29931 ( \37834 , RIe45d880_5952);
not \U$29932 ( \37835 , \37834 );
nand \U$29933 ( \37836 , \37832 , \37833 , \37835 );
not \U$29934 ( \37837 , \37836 );
not \U$29935 ( \37838 , \37837 );
buf \U$29936 ( \37839 , RIb79b4a0_271);
and \U$29937 ( \37840 , \13923 , \8863 );
buf \U$29938 ( \37841 , \37840 );
nand \U$29939 ( \37842 , \37839 , \37841 );
not \U$29940 ( \37843 , \37842 );
not \U$29941 ( \37844 , \37843 );
and \U$29942 ( \37845 , \37835 , \37844 );
nor \U$29943 ( \37846 , \37833 , \37832 );
xnor \U$29944 ( \37847 , \37834 , \37846 );
and \U$29945 ( \37848 , \37847 , \37843 );
or \U$29946 ( \37849 , \37845 , \37848 );
not \U$29947 ( \37850 , \37849 );
and \U$29948 ( \37851 , \37838 , \37850 );
buf \U$29949 ( \37852 , RIb79b338_274);
buf \U$29950 ( \37853 , \37852 );
nand \U$29951 ( \37854 , \37841 , \37853 );
not \U$29952 ( \37855 , \37854 );
nor \U$29953 ( \37856 , \37851 , \37855 );
not \U$29954 ( \37857 , \37856 );
and \U$29955 ( \37858 , \37831 , \37857 );
not \U$29956 ( \37859 , RIe444fb0_5975);
nor \U$29957 ( \37860 , \37858 , \37859 );
nand \U$29958 ( \37861 , \37860 , \37672 );
not \U$29959 ( \37862 , \37861 );
not \U$29960 ( \37863 , \37831 );
and \U$29961 ( \37864 , \37863 , \37856 );
or \U$29962 ( \37865 , \37811 , \37827 );
or \U$29963 ( \37866 , \37814 , \37819 );
or \U$29964 ( \37867 , \37826 , RIe454988_5966);
nand \U$29965 ( \37868 , \37800 , \32652 );
not \U$29966 ( \37869 , \37868 );
nand \U$29967 ( \37870 , \37869 , \37805 );
not \U$29968 ( \37871 , \37870 );
nand \U$29969 ( \37872 , RIe454988_5966, \37817 );
and \U$29970 ( \37873 , \37819 , \37872 );
or \U$29971 ( \37874 , \37873 , \37868 );
and \U$29972 ( \37875 , \37874 , \37806 );
or \U$29973 ( \37876 , \37871 , \37875 );
nand \U$29974 ( \37877 , \37865 , \37866 , \37867 , \37876 );
not \U$29975 ( \37878 , \37877 );
xor \U$29976 ( \37879 , \37815 , \37827 );
not \U$29977 ( \37880 , \37826 );
and \U$29978 ( \37881 , \37879 , \37880 );
not \U$29979 ( \37882 , \37815 );
not \U$29980 ( \37883 , \37882 );
not \U$29981 ( \37884 , \37810 );
or \U$29982 ( \37885 , \37883 , \37884 );
not \U$29983 ( \37886 , \37823 );
nand \U$29984 ( \37887 , \37815 , \37817 , \37886 );
nand \U$29985 ( \37888 , \37885 , \37887 , \37870 );
or \U$29986 ( \37889 , \37881 , \37888 );
xor \U$29987 ( \37890 , \37833 , \37832 );
and \U$29988 ( \37891 , \37854 , \37843 );
and \U$29989 ( \37892 , \37890 , \37836 , \37891 );
not \U$29990 ( \37893 , \37833 );
and \U$29991 ( \37894 , \37842 , \37893 , \37854 );
or \U$29992 ( \37895 , \37892 , \37894 );
not \U$29993 ( \37896 , \37895 );
or \U$29994 ( \37897 , \37889 , \37896 );
and \U$29995 ( \37898 , \37832 , \37836 , \37891 );
not \U$29996 ( \37899 , \37832 );
and \U$29997 ( \37900 , \37842 , \37899 , \37854 );
nor \U$29998 ( \37901 , \37898 , \37900 );
nand \U$29999 ( \37902 , \37897 , \37901 );
or \U$30000 ( \37903 , \37878 , \37902 );
nand \U$30001 ( \37904 , \37889 , \37896 );
nand \U$30002 ( \37905 , \37903 , \37904 );
not \U$30003 ( \37906 , \37905 );
nor \U$30004 ( \37907 , \37864 , \37906 );
not \U$30005 ( \37908 , \37907 );
and \U$30006 ( \37909 , \37862 , \37908 );
not \U$30007 ( \37910 , RIe45a478_5957);
not \U$30008 ( \37911 , \37910 );
or \U$30009 ( \37912 , RIe45aec8_5956, \37911 );
not \U$30010 ( \37913 , \37912 );
and \U$30011 ( \37914 , \37913 , RIe45b8a0_5955);
nand \U$30012 ( \37915 , \32658 , \32662 );
not \U$30013 ( \37916 , \37915 );
or \U$30014 ( \37917 , \37666 , \37859 );
nand \U$30015 ( \37918 , \37917 , \32658 , \32662 );
nor \U$30016 ( \37919 , \37843 , \37855 );
nand \U$30017 ( \37920 , \37916 , \37918 , \37919 );
or \U$30018 ( \37921 , \37914 , \37920 );
nand \U$30019 ( \37922 , \32658 , \32662 );
not \U$30020 ( \37923 , \37922 );
not \U$30021 ( \37924 , \37923 );
not \U$30022 ( \37925 , \37912 );
not \U$30023 ( \37926 , \37925 );
or \U$30024 ( \37927 , RIe45b8a0_5955, \37926 );
nand \U$30025 ( \37928 , \37924 , \37891 , \37927 );
nand \U$30026 ( \37929 , \37921 , \37928 );
not \U$30027 ( \37930 , \37929 );
nand \U$30028 ( \37931 , \37925 , \37922 );
not \U$30029 ( \37932 , \37923 );
or \U$30030 ( \37933 , \37910 , \37932 );
not \U$30031 ( \37934 , \37933 );
not \U$30032 ( \37935 , RIe45aec8_5956);
and \U$30033 ( \37936 , \37934 , \37935 );
not \U$30034 ( \37937 , \37910 );
xnor \U$30035 ( \37938 , \37923 , \37937 );
not \U$30036 ( \37939 , \37938 );
and \U$30037 ( \37940 , \37939 , RIe45aec8_5956);
or \U$30038 ( \37941 , \37936 , \37940 );
not \U$30039 ( \37942 , \37941 );
and \U$30040 ( \37943 , \37931 , \37942 );
or \U$30041 ( \37944 , \37930 , \37943 );
not \U$30042 ( \37945 , \37855 );
not \U$30043 ( \37946 , \37918 );
not \U$30044 ( \37947 , \37946 );
xnor \U$30045 ( \37948 , \37843 , \37923 );
and \U$30046 ( \37949 , \37945 , \37947 , \37948 );
not \U$30047 ( \37950 , \37949 );
not \U$30048 ( \37951 , \37950 );
and \U$30049 ( \37952 , \37951 , RIe45aec8_5956);
nand \U$30050 ( \37953 , \37946 , \37854 );
not \U$30051 ( \37954 , \37953 );
and \U$30052 ( \37955 , RIe4534e8_5968, \37954 );
nor \U$30053 ( \37956 , \37952 , \37955 );
nand \U$30054 ( \37957 , \37944 , \37956 );
not \U$30055 ( \37958 , \37953 );
and \U$30056 ( \37959 , RIe452b88_5969, \37958 );
not \U$30057 ( \37960 , \37951 );
not \U$30058 ( \37961 , \37910 );
and \U$30059 ( \37962 , \37960 , \37961 );
not \U$30060 ( \37963 , \37929 );
and \U$30061 ( \37964 , \37963 , \37910 );
or \U$30062 ( \37965 , \37962 , \37964 );
not \U$30063 ( \37966 , \37965 );
or \U$30064 ( \37967 , \37959 , \37966 );
nor \U$30065 ( \37968 , \37957 , \37967 );
not \U$30066 ( \37969 , \37953 );
and \U$30067 ( \37970 , RIe453fb0_5967, \37969 );
or \U$30068 ( \37971 , \37923 , \37925 );
nand \U$30069 ( \37972 , RIe45aec8_5956, \37937 );
nand \U$30070 ( \37973 , \37971 , \37972 );
xnor \U$30071 ( \37974 , \37973 , \37922 );
nor \U$30072 ( \37975 , \37930 , \37974 );
not \U$30073 ( \37976 , \37975 );
not \U$30074 ( \37977 , RIe45b8a0_5955);
and \U$30075 ( \37978 , \37976 , \37977 );
not \U$30076 ( \37979 , \37951 );
not \U$30077 ( \37980 , \37974 );
and \U$30078 ( \37981 , \37979 , \37980 );
nand \U$30079 ( \37982 , \37920 , \37928 );
nor \U$30080 ( \37983 , \37951 , \37982 );
nor \U$30081 ( \37984 , \37981 , \37983 );
not \U$30082 ( \37985 , \37984 );
and \U$30083 ( \37986 , \37985 , RIe45b8a0_5955);
or \U$30084 ( \37987 , \37978 , \37986 );
not \U$30085 ( \37988 , \37987 );
or \U$30086 ( \37989 , \37970 , \37988 );
not \U$30087 ( \37990 , \37989 );
and \U$30088 ( \37991 , \37968 , \37990 );
or \U$30089 ( \37992 , \37909 , \37991 );
not \U$30090 ( \37993 , \37992 );
and \U$30092 ( \37994 , \37993 , 1'b1 );
or \U$30094 ( \37995 , \37994 , 1'b0 );
buf \U$30095 ( \37996 , \37995 );
_DC r23c20_GF_IsGateDCbyConstraint ( \37997_nR23c20 , \37996 , \21944 );
buf \U$30096 ( \37998 , \37997_nR23c20 );
and \U$30098 ( \37999 , \37967 , 1'b1 );
or \U$30100 ( \38000 , \37999 , 1'b0 );
buf \U$30101 ( \38001 , \38000 );
_DC r23c52_GF_IsGateDCbyConstraint ( \38002_nR23c52 , \38001 , \21944 );
buf \U$30102 ( \38003 , \38002_nR23c52 );
and \U$30104 ( \38004 , \37957 , 1'b1 );
or \U$30106 ( \38005 , \38004 , 1'b0 );
buf \U$30107 ( \38006 , \38005 );
_DC r23c54_GF_IsGateDCbyConstraint ( \38007_nR23c54 , \38006 , \21944 );
buf \U$30108 ( \38008 , \38007_nR23c54 );
and \U$30110 ( \38009 , \37989 , 1'b1 );
or \U$30112 ( \38010 , \38009 , 1'b0 );
buf \U$30113 ( \38011 , \38010 );
_DC r23c56_GF_IsGateDCbyConstraint ( \38012_nR23c56 , \38011 , \21944 );
buf \U$30114 ( \38013 , \38012_nR23c56 );
not \U$30115 ( \38014 , \21810 );
nand \U$30116 ( \38015 , \38014 , \21812 , RIe546098_6850);
nor \U$30117 ( \38016 , \21809 , \38015 );
buf \U$30118 ( \38017 , \38016 );
buf \U$30119 ( \38018 , \38017 );
not \U$30120 ( \38019 , \22095 );
buf \U$30121 ( \38020 , \38019 );
buf \U$30122 ( \38021 , \38020 );
nand \U$30123 ( \38022 , \38018 , \38021 );
not \U$30124 ( \38023 , \38022 );
buf \U$30125 ( \38024 , \8825 );
buf \U$30126 ( \38025 , \38024 );
not \U$30127 ( \38026 , \27242 );
and \U$30128 ( \38027 , \38026 , \21694 );
buf \U$30129 ( \38028 , \38027 );
buf \U$30130 ( \38029 , \38028 );
nand \U$30131 ( \38030 , \38025 , \38029 );
not \U$30132 ( \38031 , \38030 );
or \U$30133 ( \38032 , \38023 , \38031 );
buf \U$30134 ( \38033 , \38032 );
buf \U$30135 ( \38034 , \38033 );
not \U$30136 ( \38035 , \38034 );
and \U$30137 ( \38036 , RIe116b70_5293, \38035 );
not \U$30138 ( \38037 , RIe116b70_5293);
buf \U$30139 ( \38038 , \22109 );
buf \U$30140 ( \38039 , \27371 );
not \U$30141 ( \38040 , \38039 );
not \U$30142 ( \38041 , \38040 );
or \U$30143 ( \38042 , \38038 , \38041 );
not \U$30144 ( \38043 , \38042 );
nand \U$30145 ( \38044 , \38030 , \38043 );
not \U$30146 ( \38045 , \27378 );
buf \U$30147 ( \38046 , \38045 );
buf \U$30148 ( \38047 , RIeab7058_6894);
or \U$30149 ( \38048 , \38046 , \38047 , \38030 );
buf \U$30150 ( \38049 , \38048 );
and \U$30151 ( \38050 , \38044 , \38049 );
not \U$30152 ( \38051 , \38050 );
or \U$30153 ( \38052 , \38037 , \38051 );
not \U$30154 ( \38053 , \38044 );
buf \U$30155 ( \38054 , \38053 );
buf \U$30156 ( \38055 , \22131 );
and \U$30157 ( \38056 , \38054 , \38055 );
buf \U$30158 ( \38057 , RIb7c5980_237);
buf \U$30159 ( \38058 , \38057 );
not \U$30160 ( \38059 , \38049 );
and \U$30161 ( \38060 , \38058 , \38059 );
nor \U$30162 ( \38061 , \38056 , \38060 );
nand \U$30163 ( \38062 , \38052 , \38061 );
and \U$30164 ( \38063 , \38062 , \38034 );
or \U$30165 ( \38064 , \38036 , \38063 );
and \U$30167 ( \38065 , \38064 , 1'b1 );
or \U$30169 ( \38066 , \38065 , 1'b0 );
buf \U$30170 ( \38067 , \38066 );
_DC r23774_GF_IsGateDCbyConstraint ( \38068_nR23774 , \38067 , \21944 );
buf \U$30171 ( \38069 , \38068_nR23774 );
not \U$30172 ( \38070 , \38034 );
and \U$30173 ( \38071 , RIe115a18_5294, \38070 );
not \U$30174 ( \38072 , RIe115a18_5294);
not \U$30175 ( \38073 , \38046 );
not \U$30176 ( \38074 , \38047 );
and \U$30177 ( \38075 , \38073 , \38074 , \38031 );
not \U$30178 ( \38076 , \38075 );
buf \U$30179 ( \38077 , \38076 );
and \U$30180 ( \38078 , \38044 , \38077 );
not \U$30181 ( \38079 , \38078 );
or \U$30182 ( \38080 , \38072 , \38079 );
buf \U$30183 ( \38081 , \38053 );
buf \U$30184 ( \38082 , RIb87eb78_68);
buf \U$30185 ( \38083 , \38082 );
and \U$30186 ( \38084 , \38081 , \38083 );
buf \U$30187 ( \38085 , \22161 );
buf \U$30188 ( \38086 , \38048 );
not \U$30189 ( \38087 , \38086 );
and \U$30190 ( \38088 , \38085 , \38087 );
nor \U$30191 ( \38089 , \38084 , \38088 );
nand \U$30192 ( \38090 , \38080 , \38089 );
and \U$30193 ( \38091 , \38090 , \38034 );
or \U$30194 ( \38092 , \38071 , \38091 );
and \U$30196 ( \38093 , \38092 , 1'b1 );
or \U$30198 ( \38094 , \38093 , 1'b0 );
buf \U$30199 ( \38095 , \38094 );
_DC r2378a_GF_IsGateDCbyConstraint ( \38096_nR2378a , \38095 , \21944 );
buf \U$30200 ( \38097 , \38096_nR2378a );
not \U$30201 ( \38098 , \38034 );
and \U$30202 ( \38099 , RIe114410_5295, \38098 );
not \U$30203 ( \38100 , RIe114410_5295);
or \U$30204 ( \38101 , \38100 , \38051 );
buf \U$30205 ( \38102 , RIb87ebf0_67);
and \U$30206 ( \38103 , \38081 , \38102 );
buf \U$30207 ( \38104 , RIb7c5a70_235);
buf \U$30208 ( \38105 , \38104 );
not \U$30209 ( \38106 , \38049 );
and \U$30210 ( \38107 , \38105 , \38106 );
nor \U$30211 ( \38108 , \38103 , \38107 );
nand \U$30212 ( \38109 , \38101 , \38108 );
and \U$30213 ( \38110 , \38109 , \38034 );
or \U$30214 ( \38111 , \38099 , \38110 );
and \U$30216 ( \38112 , \38111 , 1'b1 );
or \U$30218 ( \38113 , \38112 , 1'b0 );
buf \U$30219 ( \38114 , \38113 );
_DC r237a0_GF_IsGateDCbyConstraint ( \38115_nR237a0 , \38114 , \21944 );
buf \U$30220 ( \38116 , \38115_nR237a0 );
buf \U$30221 ( \38117 , \38033 );
not \U$30222 ( \38118 , \38117 );
and \U$30223 ( \38119 , RIe1132b8_5296, \38118 );
not \U$30224 ( \38120 , RIe1132b8_5296);
not \U$30225 ( \38121 , \38078 );
or \U$30226 ( \38122 , \38120 , \38121 );
buf \U$30227 ( \38123 , \22202 );
and \U$30228 ( \38124 , \38081 , \38123 );
buf \U$30229 ( \38125 , RIb7cade0_234);
buf \U$30230 ( \38126 , \38125 );
not \U$30231 ( \38127 , \38077 );
and \U$30232 ( \38128 , \38126 , \38127 );
nor \U$30233 ( \38129 , \38124 , \38128 );
nand \U$30234 ( \38130 , \38122 , \38129 );
and \U$30235 ( \38131 , \38130 , \38117 );
or \U$30236 ( \38132 , \38119 , \38131 );
and \U$30238 ( \38133 , \38132 , 1'b1 );
or \U$30240 ( \38134 , \38133 , 1'b0 );
buf \U$30241 ( \38135 , \38134 );
_DC r237b6_GF_IsGateDCbyConstraint ( \38136_nR237b6 , \38135 , \21944 );
buf \U$30242 ( \38137 , \38136_nR237b6 );
not \U$30243 ( \38138 , \38117 );
and \U$30244 ( \38139 , RIe111cb0_5297, \38138 );
not \U$30245 ( \38140 , RIe111cb0_5297);
not \U$30246 ( \38141 , \38050 );
or \U$30247 ( \38142 , \38140 , \38141 );
buf \U$30248 ( \38143 , RIb885310_65);
and \U$30249 ( \38144 , \38054 , \38143 );
buf \U$30250 ( \38145 , \22226 );
not \U$30251 ( \38146 , \38086 );
and \U$30252 ( \38147 , \38145 , \38146 );
nor \U$30253 ( \38148 , \38144 , \38147 );
nand \U$30254 ( \38149 , \38142 , \38148 );
and \U$30255 ( \38150 , \38149 , \38117 );
or \U$30256 ( \38151 , \38139 , \38150 );
and \U$30258 ( \38152 , \38151 , 1'b1 );
or \U$30260 ( \38153 , \38152 , 1'b0 );
buf \U$30261 ( \38154 , \38153 );
_DC r237cc_GF_IsGateDCbyConstraint ( \38155_nR237cc , \38154 , \21944 );
buf \U$30262 ( \38156 , \38155_nR237cc );
not \U$30263 ( \38157 , \38034 );
and \U$30264 ( \38158 , RIe110b58_5298, \38157 );
not \U$30265 ( \38159 , RIe110b58_5298);
not \U$30266 ( \38160 , \38078 );
or \U$30267 ( \38161 , \38159 , \38160 );
buf \U$30268 ( \38162 , \38053 );
buf \U$30269 ( \38163 , \32803 );
and \U$30270 ( \38164 , \38162 , \38163 );
buf \U$30271 ( \38165 , RIb7caed0_232);
buf \U$30272 ( \38166 , \38165 );
not \U$30273 ( \38167 , \38046 );
not \U$30274 ( \38168 , \38047 );
and \U$30275 ( \38169 , \38167 , \38168 , \38031 );
not \U$30276 ( \38170 , \38169 );
buf \U$30277 ( \38171 , \38170 );
not \U$30278 ( \38172 , \38171 );
and \U$30279 ( \38173 , \38166 , \38172 );
nor \U$30280 ( \38174 , \38164 , \38173 );
nand \U$30281 ( \38175 , \38161 , \38174 );
and \U$30282 ( \38176 , \38175 , \38034 );
or \U$30283 ( \38177 , \38158 , \38176 );
and \U$30285 ( \38178 , \38177 , 1'b1 );
or \U$30287 ( \38179 , \38178 , 1'b0 );
buf \U$30288 ( \38180 , \38179 );
_DC r237e2_GF_IsGateDCbyConstraint ( \38181_nR237e2 , \38180 , \21944 );
buf \U$30289 ( \38182 , \38181_nR237e2 );
not \U$30290 ( \38183 , \38034 );
and \U$30291 ( \38184 , RIe10f550_5299, \38183 );
not \U$30292 ( \38185 , RIe10f550_5299);
not \U$30293 ( \38186 , \38050 );
or \U$30294 ( \38187 , \38185 , \38186 );
buf \U$30295 ( \38188 , RIb885400_63);
and \U$30296 ( \38189 , \38054 , \38188 );
buf \U$30297 ( \38190 , RIb7caf48_231);
buf \U$30298 ( \38191 , \38190 );
not \U$30299 ( \38192 , \38077 );
and \U$30300 ( \38193 , \38191 , \38192 );
nor \U$30301 ( \38194 , \38189 , \38193 );
nand \U$30302 ( \38195 , \38187 , \38194 );
and \U$30303 ( \38196 , \38195 , \38034 );
or \U$30304 ( \38197 , \38184 , \38196 );
and \U$30306 ( \38198 , \38197 , 1'b1 );
or \U$30308 ( \38199 , \38198 , 1'b0 );
buf \U$30309 ( \38200 , \38199 );
_DC r237ec_GF_IsGateDCbyConstraint ( \38201_nR237ec , \38200 , \21944 );
buf \U$30310 ( \38202 , \38201_nR237ec );
not \U$30311 ( \38203 , \38034 );
and \U$30312 ( \38204 , RIe10e3f8_5300, \38203 );
not \U$30313 ( \38205 , RIe10e3f8_5300);
or \U$30314 ( \38206 , \38205 , \38160 );
buf \U$30315 ( \38207 , \32847 );
and \U$30316 ( \38208 , \38162 , \38207 );
buf \U$30317 ( \38209 , RIb7cafc0_230);
buf \U$30318 ( \38210 , \38209 );
buf \U$30319 ( \38211 , \38170 );
not \U$30320 ( \38212 , \38211 );
and \U$30321 ( \38213 , \38210 , \38212 );
nor \U$30322 ( \38214 , \38208 , \38213 );
nand \U$30323 ( \38215 , \38206 , \38214 );
and \U$30324 ( \38216 , \38215 , \38034 );
or \U$30325 ( \38217 , \38204 , \38216 );
and \U$30327 ( \38218 , \38217 , 1'b1 );
or \U$30329 ( \38219 , \38218 , 1'b0 );
buf \U$30330 ( \38220 , \38219 );
_DC r237ee_GF_IsGateDCbyConstraint ( \38221_nR237ee , \38220 , \21944 );
buf \U$30331 ( \38222 , \38221_nR237ee );
buf \U$30332 ( \38223 , \38033 );
not \U$30333 ( \38224 , \38223 );
and \U$30334 ( \38225 , RIe10d2a0_5301, \38224 );
not \U$30335 ( \38226 , RIe10d2a0_5301);
or \U$30336 ( \38227 , \38226 , \38121 );
buf \U$30337 ( \38228 , \22313 );
and \U$30338 ( \38229 , \38162 , \38228 );
buf \U$30339 ( \38230 , \22316 );
buf \U$30340 ( \38231 , \38170 );
not \U$30341 ( \38232 , \38231 );
and \U$30342 ( \38233 , \38230 , \38232 );
nor \U$30343 ( \38234 , \38229 , \38233 );
nand \U$30344 ( \38235 , \38227 , \38234 );
and \U$30345 ( \38236 , \38235 , \38223 );
or \U$30346 ( \38237 , \38225 , \38236 );
and \U$30348 ( \38238 , \38237 , 1'b1 );
or \U$30350 ( \38239 , \38238 , 1'b0 );
buf \U$30351 ( \38240 , \38239 );
_DC r237f0_GF_IsGateDCbyConstraint ( \38241_nR237f0 , \38240 , \21944 );
buf \U$30352 ( \38242 , \38241_nR237f0 );
not \U$30353 ( \38243 , \38117 );
and \U$30354 ( \38244 , RIe10bc98_5302, \38243 );
not \U$30355 ( \38245 , RIe10bc98_5302);
or \U$30356 ( \38246 , \38245 , \38160 );
buf \U$30357 ( \38247 , \22334 );
and \U$30358 ( \38248 , \38054 , \38247 );
buf \U$30359 ( \38249 , RIb7cb0b0_228);
buf \U$30360 ( \38250 , \38249 );
buf \U$30361 ( \38251 , \38076 );
not \U$30362 ( \38252 , \38251 );
and \U$30363 ( \38253 , \38250 , \38252 );
nor \U$30364 ( \38254 , \38248 , \38253 );
nand \U$30365 ( \38255 , \38246 , \38254 );
and \U$30366 ( \38256 , \38255 , \38117 );
or \U$30367 ( \38257 , \38244 , \38256 );
and \U$30369 ( \38258 , \38257 , 1'b1 );
or \U$30371 ( \38259 , \38258 , 1'b0 );
buf \U$30372 ( \38260 , \38259 );
_DC r237f2_GF_IsGateDCbyConstraint ( \38261_nR237f2 , \38260 , \21944 );
buf \U$30373 ( \38262 , \38261_nR237f2 );
not \U$30374 ( \38263 , \38034 );
and \U$30375 ( \38264 , RIe10ab40_5303, \38263 );
not \U$30376 ( \38265 , RIe10ab40_5303);
not \U$30377 ( \38266 , \38050 );
or \U$30378 ( \38267 , \38265 , \38266 );
buf \U$30379 ( \38268 , \38053 );
buf \U$30380 ( \38269 , RIb8855e0_59);
and \U$30381 ( \38270 , \38268 , \38269 );
buf \U$30382 ( \38271 , \27608 );
not \U$30383 ( \38272 , \38171 );
and \U$30384 ( \38273 , \38271 , \38272 );
nor \U$30385 ( \38274 , \38270 , \38273 );
nand \U$30386 ( \38275 , \38267 , \38274 );
and \U$30387 ( \38276 , \38275 , \38034 );
or \U$30388 ( \38277 , \38264 , \38276 );
and \U$30390 ( \38278 , \38277 , 1'b1 );
or \U$30392 ( \38279 , \38278 , 1'b0 );
buf \U$30393 ( \38280 , \38279 );
_DC r23776_GF_IsGateDCbyConstraint ( \38281_nR23776 , \38280 , \21944 );
buf \U$30394 ( \38282 , \38281_nR23776 );
not \U$30395 ( \38283 , \38223 );
and \U$30396 ( \38284 , RIe109538_5304, \38283 );
not \U$30397 ( \38285 , RIe109538_5304);
or \U$30398 ( \38286 , \38285 , \38141 );
buf \U$30399 ( \38287 , \22376 );
and \U$30400 ( \38288 , \38081 , \38287 );
buf \U$30401 ( \38289 , RIb7d00d8_226);
buf \U$30402 ( \38290 , \38289 );
not \U$30403 ( \38291 , \38211 );
and \U$30404 ( \38292 , \38290 , \38291 );
nor \U$30405 ( \38293 , \38288 , \38292 );
nand \U$30406 ( \38294 , \38286 , \38293 );
and \U$30407 ( \38295 , \38294 , \38223 );
or \U$30408 ( \38296 , \38284 , \38295 );
and \U$30410 ( \38297 , \38296 , 1'b1 );
or \U$30412 ( \38298 , \38297 , 1'b0 );
buf \U$30413 ( \38299 , \38298 );
_DC r23778_GF_IsGateDCbyConstraint ( \38300_nR23778 , \38299 , \21944 );
buf \U$30414 ( \38301 , \38300_nR23778 );
not \U$30415 ( \38302 , \38034 );
and \U$30416 ( \38303 , RIe1083e0_5305, \38302 );
not \U$30417 ( \38304 , RIe1083e0_5305);
not \U$30418 ( \38305 , \38050 );
or \U$30419 ( \38306 , \38304 , \38305 );
buf \U$30420 ( \38307 , RIb8856d0_57);
and \U$30421 ( \38308 , \38162 , \38307 );
buf \U$30422 ( \38309 , \27647 );
not \U$30423 ( \38310 , \38231 );
and \U$30424 ( \38311 , \38309 , \38310 );
nor \U$30425 ( \38312 , \38308 , \38311 );
nand \U$30426 ( \38313 , \38306 , \38312 );
and \U$30427 ( \38314 , \38313 , \38034 );
or \U$30428 ( \38315 , \38303 , \38314 );
and \U$30430 ( \38316 , \38315 , 1'b1 );
or \U$30432 ( \38317 , \38316 , 1'b0 );
buf \U$30433 ( \38318 , \38317 );
_DC r2377a_GF_IsGateDCbyConstraint ( \38319_nR2377a , \38318 , \21944 );
buf \U$30434 ( \38320 , \38319_nR2377a );
not \U$30435 ( \38321 , \38034 );
and \U$30436 ( \38322 , RIe106dd8_5306, \38321 );
not \U$30437 ( \38323 , RIe106dd8_5306);
or \U$30438 ( \38324 , \38323 , \38079 );
buf \U$30439 ( \38325 , RIb885748_56);
and \U$30440 ( \38326 , \38081 , \38325 );
buf \U$30441 ( \38327 , RIb826e28_224);
buf \U$30442 ( \38328 , \38327 );
buf \U$30443 ( \38329 , \38076 );
not \U$30444 ( \38330 , \38329 );
and \U$30445 ( \38331 , \38328 , \38330 );
nor \U$30446 ( \38332 , \38326 , \38331 );
nand \U$30447 ( \38333 , \38324 , \38332 );
and \U$30448 ( \38334 , \38333 , \38034 );
or \U$30449 ( \38335 , \38322 , \38334 );
and \U$30451 ( \38336 , \38335 , 1'b1 );
or \U$30453 ( \38337 , \38336 , 1'b0 );
buf \U$30454 ( \38338 , \38337 );
_DC r2377c_GF_IsGateDCbyConstraint ( \38339_nR2377c , \38338 , \21944 );
buf \U$30455 ( \38340 , \38339_nR2377c );
not \U$30456 ( \38341 , \38223 );
and \U$30457 ( \38342 , RIdfd3728_5307, \38341 );
not \U$30458 ( \38343 , RIdfd3728_5307);
or \U$30459 ( \38344 , \38343 , \38121 );
buf \U$30460 ( \38345 , RIb8857c0_55);
buf \U$30461 ( \38346 , \38345 );
and \U$30462 ( \38347 , \38081 , \38346 );
buf \U$30463 ( \38348 , RIb826ea0_223);
buf \U$30464 ( \38349 , \38348 );
not \U$30465 ( \38350 , \38251 );
and \U$30466 ( \38351 , \38349 , \38350 );
nor \U$30467 ( \38352 , \38347 , \38351 );
nand \U$30468 ( \38353 , \38344 , \38352 );
and \U$30469 ( \38354 , \38353 , \38223 );
or \U$30470 ( \38355 , \38342 , \38354 );
and \U$30472 ( \38356 , \38355 , 1'b1 );
or \U$30474 ( \38357 , \38356 , 1'b0 );
buf \U$30475 ( \38358 , \38357 );
_DC r2377e_GF_IsGateDCbyConstraint ( \38359_nR2377e , \38358 , \21944 );
buf \U$30476 ( \38360 , \38359_nR2377e );
not \U$30477 ( \38361 , \38117 );
and \U$30478 ( \38362 , RIdfd71c0_5308, \38361 );
not \U$30479 ( \38363 , RIdfd71c0_5308);
or \U$30480 ( \38364 , \38363 , \38051 );
buf \U$30481 ( \38365 , RIb885838_54);
and \U$30482 ( \38366 , \38268 , \38365 );
buf \U$30483 ( \38367 , RIb826f18_222);
buf \U$30484 ( \38368 , \38367 );
not \U$30485 ( \38369 , \38077 );
and \U$30486 ( \38370 , \38368 , \38369 );
nor \U$30487 ( \38371 , \38366 , \38370 );
nand \U$30488 ( \38372 , \38364 , \38371 );
and \U$30489 ( \38373 , \38372 , \38117 );
or \U$30490 ( \38374 , \38362 , \38373 );
and \U$30492 ( \38375 , \38374 , 1'b1 );
or \U$30494 ( \38376 , \38375 , 1'b0 );
buf \U$30495 ( \38377 , \38376 );
_DC r23780_GF_IsGateDCbyConstraint ( \38378_nR23780 , \38377 , \21944 );
buf \U$30496 ( \38379 , \38378_nR23780 );
not \U$30497 ( \38380 , \38117 );
and \U$30498 ( \38381 , RIdfdc8f0_5309, \38380 );
not \U$30499 ( \38382 , RIdfdc8f0_5309);
or \U$30500 ( \38383 , \38382 , \38266 );
buf \U$30501 ( \38384 , \22477 );
and \U$30502 ( \38385 , \38268 , \38384 );
buf \U$30503 ( \38386 , RIb826f90_221);
buf \U$30504 ( \38387 , \38386 );
not \U$30505 ( \38388 , \38086 );
and \U$30506 ( \38389 , \38387 , \38388 );
nor \U$30507 ( \38390 , \38385 , \38389 );
nand \U$30508 ( \38391 , \38383 , \38390 );
and \U$30509 ( \38392 , \38391 , \38117 );
or \U$30510 ( \38393 , \38381 , \38392 );
and \U$30512 ( \38394 , \38393 , 1'b1 );
or \U$30514 ( \38395 , \38394 , 1'b0 );
buf \U$30515 ( \38396 , \38395 );
_DC r23782_GF_IsGateDCbyConstraint ( \38397_nR23782 , \38396 , \21944 );
buf \U$30516 ( \38398 , \38397_nR23782 );
not \U$30517 ( \38399 , \38223 );
and \U$30518 ( \38400 , RIdfe0b80_5310, \38399 );
not \U$30519 ( \38401 , RIdfe0b80_5310);
or \U$30520 ( \38402 , \38401 , \38141 );
buf \U$30521 ( \38403 , \22497 );
and \U$30522 ( \38404 , \38081 , \38403 );
buf \U$30523 ( \38405 , RIb8293a8_220);
buf \U$30524 ( \38406 , \38405 );
buf \U$30525 ( \38407 , \38048 );
not \U$30526 ( \38408 , \38407 );
and \U$30527 ( \38409 , \38406 , \38408 );
nor \U$30528 ( \38410 , \38404 , \38409 );
nand \U$30529 ( \38411 , \38402 , \38410 );
and \U$30530 ( \38412 , \38411 , \38223 );
or \U$30531 ( \38413 , \38400 , \38412 );
and \U$30533 ( \38414 , \38413 , 1'b1 );
or \U$30535 ( \38415 , \38414 , 1'b0 );
buf \U$30536 ( \38416 , \38415 );
_DC r23784_GF_IsGateDCbyConstraint ( \38417_nR23784 , \38416 , \21944 );
buf \U$30537 ( \38418 , \38417_nR23784 );
not \U$30538 ( \38419 , \38117 );
and \U$30539 ( \38420 , RIdfe6760_5311, \38419 );
not \U$30540 ( \38421 , RIdfe6760_5311);
or \U$30541 ( \38422 , \38421 , \38305 );
buf \U$30542 ( \38423 , RIb8859a0_51);
and \U$30543 ( \38424 , \38081 , \38423 );
buf \U$30544 ( \38425 , \27759 );
not \U$30545 ( \38426 , \38086 );
and \U$30546 ( \38427 , \38425 , \38426 );
nor \U$30547 ( \38428 , \38424 , \38427 );
nand \U$30548 ( \38429 , \38422 , \38428 );
and \U$30549 ( \38430 , \38429 , \38117 );
or \U$30550 ( \38431 , \38420 , \38430 );
and \U$30552 ( \38432 , \38431 , 1'b1 );
or \U$30554 ( \38433 , \38432 , 1'b0 );
buf \U$30555 ( \38434 , \38433 );
_DC r23786_GF_IsGateDCbyConstraint ( \38435_nR23786 , \38434 , \21944 );
buf \U$30556 ( \38436 , \38435_nR23786 );
not \U$30557 ( \38437 , \38034 );
and \U$30558 ( \38438 , RIdfeb788_5312, \38437 );
not \U$30559 ( \38439 , RIdfeb788_5312);
or \U$30560 ( \38440 , \38439 , \38186 );
buf \U$30561 ( \38441 , \33087 );
and \U$30562 ( \38442 , \38081 , \38441 );
buf \U$30563 ( \38443 , \22541 );
not \U$30564 ( \38444 , \38049 );
and \U$30565 ( \38445 , \38443 , \38444 );
nor \U$30566 ( \38446 , \38442 , \38445 );
nand \U$30567 ( \38447 , \38440 , \38446 );
and \U$30568 ( \38448 , \38447 , \38034 );
or \U$30569 ( \38449 , \38438 , \38448 );
and \U$30571 ( \38450 , \38449 , 1'b1 );
or \U$30573 ( \38451 , \38450 , 1'b0 );
buf \U$30574 ( \38452 , \38451 );
_DC r23788_GF_IsGateDCbyConstraint ( \38453_nR23788 , \38452 , \21944 );
buf \U$30575 ( \38454 , \38453_nR23788 );
not \U$30576 ( \38455 , \38223 );
and \U$30577 ( \38456 , RIdff1f98_5313, \38455 );
not \U$30578 ( \38457 , RIdff1f98_5313);
or \U$30579 ( \38458 , \38457 , \38121 );
buf \U$30580 ( \38459 , \22558 );
and \U$30581 ( \38460 , \38268 , \38459 );
buf \U$30582 ( \38461 , RIb829510_217);
buf \U$30583 ( \38462 , \38461 );
not \U$30584 ( \38463 , \38407 );
and \U$30585 ( \38464 , \38462 , \38463 );
nor \U$30586 ( \38465 , \38460 , \38464 );
nand \U$30587 ( \38466 , \38458 , \38465 );
and \U$30588 ( \38467 , \38466 , \38223 );
or \U$30589 ( \38468 , \38456 , \38467 );
and \U$30591 ( \38469 , \38468 , 1'b1 );
or \U$30593 ( \38470 , \38469 , 1'b0 );
buf \U$30594 ( \38471 , \38470 );
_DC r2378c_GF_IsGateDCbyConstraint ( \38472_nR2378c , \38471 , \21944 );
buf \U$30595 ( \38473 , \38472_nR2378c );
not \U$30596 ( \38474 , \38117 );
and \U$30597 ( \38475 , RIdff7f38_5314, \38474 );
not \U$30598 ( \38476 , RIdff7f38_5314);
or \U$30599 ( \38477 , \38476 , \38160 );
buf \U$30600 ( \38478 , \22578 );
and \U$30601 ( \38479 , \38054 , \38478 );
buf \U$30602 ( \38480 , RIb829588_216);
buf \U$30603 ( \38481 , \38480 );
not \U$30604 ( \38482 , \38171 );
and \U$30605 ( \38483 , \38481 , \38482 );
nor \U$30606 ( \38484 , \38479 , \38483 );
nand \U$30607 ( \38485 , \38477 , \38484 );
and \U$30608 ( \38486 , \38485 , \38117 );
or \U$30609 ( \38487 , \38475 , \38486 );
and \U$30611 ( \38488 , \38487 , 1'b1 );
or \U$30613 ( \38489 , \38488 , 1'b0 );
buf \U$30614 ( \38490 , \38489 );
_DC r2378e_GF_IsGateDCbyConstraint ( \38491_nR2378e , \38490 , \21944 );
buf \U$30615 ( \38492 , \38491_nR2378e );
not \U$30616 ( \38493 , \38117 );
and \U$30617 ( \38494 , RIdffe400_5315, \38493 );
not \U$30618 ( \38495 , RIdffe400_5315);
or \U$30619 ( \38496 , \38495 , \38186 );
buf \U$30620 ( \38497 , \33145 );
and \U$30621 ( \38498 , \38162 , \38497 );
buf \U$30622 ( \38499 , RIb829600_215);
buf \U$30623 ( \38500 , \38499 );
not \U$30624 ( \38501 , \38211 );
and \U$30625 ( \38502 , \38500 , \38501 );
nor \U$30626 ( \38503 , \38498 , \38502 );
nand \U$30627 ( \38504 , \38496 , \38503 );
and \U$30628 ( \38505 , \38504 , \38117 );
or \U$30629 ( \38506 , \38494 , \38505 );
and \U$30631 ( \38507 , \38506 , 1'b1 );
or \U$30633 ( \38508 , \38507 , 1'b0 );
buf \U$30634 ( \38509 , \38508 );
_DC r23790_GF_IsGateDCbyConstraint ( \38510_nR23790 , \38509 , \21944 );
buf \U$30635 ( \38511 , \38510_nR23790 );
not \U$30636 ( \38512 , \38223 );
and \U$30637 ( \38513 , RIe005750_5316, \38512 );
not \U$30638 ( \38514 , RIe005750_5316);
or \U$30639 ( \38515 , \38514 , \38160 );
buf \U$30640 ( \38516 , RIb885bf8_46);
and \U$30641 ( \38517 , \38054 , \38516 );
buf \U$30642 ( \38518 , \27853 );
not \U$30643 ( \38519 , \38231 );
and \U$30644 ( \38520 , \38518 , \38519 );
nor \U$30645 ( \38521 , \38517 , \38520 );
nand \U$30646 ( \38522 , \38515 , \38521 );
and \U$30647 ( \38523 , \38522 , \38223 );
or \U$30648 ( \38524 , \38513 , \38523 );
and \U$30650 ( \38525 , \38524 , 1'b1 );
or \U$30652 ( \38526 , \38525 , 1'b0 );
buf \U$30653 ( \38527 , \38526 );
_DC r23792_GF_IsGateDCbyConstraint ( \38528_nR23792 , \38527 , \21944 );
buf \U$30654 ( \38529 , \38528_nR23792 );
not \U$30655 ( \38530 , \38034 );
and \U$30656 ( \38531 , RIe00b420_5317, \38530 );
not \U$30657 ( \38532 , RIe00b420_5317);
or \U$30658 ( \38533 , \38532 , \38121 );
buf \U$30659 ( \38534 , \22639 );
and \U$30660 ( \38535 , \38268 , \38534 );
buf \U$30661 ( \38536 , RIb8296f0_213);
buf \U$30662 ( \38537 , \38536 );
not \U$30663 ( \38538 , \38171 );
and \U$30664 ( \38539 , \38537 , \38538 );
nor \U$30665 ( \38540 , \38535 , \38539 );
nand \U$30666 ( \38541 , \38533 , \38540 );
and \U$30667 ( \38542 , \38541 , \38034 );
or \U$30668 ( \38543 , \38531 , \38542 );
and \U$30670 ( \38544 , \38543 , 1'b1 );
or \U$30672 ( \38545 , \38544 , 1'b0 );
buf \U$30673 ( \38546 , \38545 );
_DC r23794_GF_IsGateDCbyConstraint ( \38547_nR23794 , \38546 , \21944 );
buf \U$30674 ( \38548 , \38547_nR23794 );
not \U$30675 ( \38549 , \38034 );
and \U$30676 ( \38550 , RIe0132b0_5318, \38549 );
not \U$30677 ( \38551 , RIe0132b0_5318);
or \U$30678 ( \38552 , \38551 , \38160 );
buf \U$30679 ( \38553 , RIb885ce8_44);
and \U$30680 ( \38554 , \38081 , \38553 );
buf \U$30681 ( \38555 , \27891 );
not \U$30682 ( \38556 , \38211 );
and \U$30683 ( \38557 , \38555 , \38556 );
nor \U$30684 ( \38558 , \38554 , \38557 );
nand \U$30685 ( \38559 , \38552 , \38558 );
and \U$30686 ( \38560 , \38559 , \38034 );
or \U$30687 ( \38561 , \38550 , \38560 );
and \U$30689 ( \38562 , \38561 , 1'b1 );
or \U$30691 ( \38563 , \38562 , 1'b0 );
buf \U$30692 ( \38564 , \38563 );
_DC r23796_GF_IsGateDCbyConstraint ( \38565_nR23796 , \38564 , \21944 );
buf \U$30693 ( \38566 , \38565_nR23796 );
not \U$30694 ( \38567 , \38223 );
and \U$30695 ( \38568 , RIe0193b8_5319, \38567 );
not \U$30696 ( \38569 , RIe0193b8_5319);
or \U$30697 ( \38570 , \38569 , \38079 );
buf \U$30698 ( \38571 , \22680 );
and \U$30699 ( \38572 , \38268 , \38571 );
buf \U$30700 ( \38573 , \22683 );
not \U$30701 ( \38574 , \38407 );
and \U$30702 ( \38575 , \38573 , \38574 );
nor \U$30703 ( \38576 , \38572 , \38575 );
nand \U$30704 ( \38577 , \38570 , \38576 );
and \U$30705 ( \38578 , \38577 , \38223 );
or \U$30706 ( \38579 , \38568 , \38578 );
and \U$30708 ( \38580 , \38579 , 1'b1 );
or \U$30710 ( \38581 , \38580 , 1'b0 );
buf \U$30711 ( \38582 , \38581 );
_DC r23798_GF_IsGateDCbyConstraint ( \38583_nR23798 , \38582 , \21944 );
buf \U$30712 ( \38584 , \38583_nR23798 );
not \U$30713 ( \38585 , \38117 );
and \U$30714 ( \38586 , RIe0202d0_5320, \38585 );
not \U$30715 ( \38587 , RIe0202d0_5320);
or \U$30716 ( \38588 , \38587 , \38121 );
buf \U$30717 ( \38589 , RIb885dd8_42);
and \U$30718 ( \38590 , \38268 , \38589 );
buf \U$30719 ( \38591 , \27929 );
not \U$30720 ( \38592 , \38329 );
and \U$30721 ( \38593 , \38591 , \38592 );
nor \U$30722 ( \38594 , \38590 , \38593 );
nand \U$30723 ( \38595 , \38588 , \38594 );
and \U$30724 ( \38596 , \38595 , \38117 );
or \U$30725 ( \38597 , \38586 , \38596 );
and \U$30727 ( \38598 , \38597 , 1'b1 );
or \U$30729 ( \38599 , \38598 , 1'b0 );
buf \U$30730 ( \38600 , \38599 );
_DC r2379a_GF_IsGateDCbyConstraint ( \38601_nR2379a , \38600 , \21944 );
buf \U$30731 ( \38602 , \38601_nR2379a );
buf \U$30732 ( \38603 , \38032 );
not \U$30733 ( \38604 , \38603 );
and \U$30734 ( \38605 , RIe023de0_5321, \38604 );
not \U$30735 ( \38606 , RIe023de0_5321);
or \U$30736 ( \38607 , \38606 , \38079 );
buf \U$30737 ( \38608 , RIb885e50_41);
buf \U$30738 ( \38609 , \38608 );
and \U$30739 ( \38610 , \38081 , \38609 );
buf \U$30740 ( \38611 , RIb82dc50_209);
buf \U$30741 ( \38612 , \38611 );
not \U$30742 ( \38613 , \38251 );
and \U$30743 ( \38614 , \38612 , \38613 );
nor \U$30744 ( \38615 , \38610 , \38614 );
nand \U$30745 ( \38616 , \38607 , \38615 );
and \U$30746 ( \38617 , \38616 , \38603 );
or \U$30747 ( \38618 , \38605 , \38617 );
and \U$30749 ( \38619 , \38618 , 1'b1 );
or \U$30751 ( \38620 , \38619 , 1'b0 );
buf \U$30752 ( \38621 , \38620 );
_DC r2379c_GF_IsGateDCbyConstraint ( \38622_nR2379c , \38621 , \21944 );
buf \U$30753 ( \38623 , \38622_nR2379c );
not \U$30754 ( \38624 , \38223 );
and \U$30755 ( \38625 , RIe027878_5322, \38624 );
not \U$30756 ( \38626 , RIe027878_5322);
or \U$30757 ( \38627 , \38626 , \38160 );
not \U$30758 ( \38628 , \38081 );
not \U$30759 ( \38629 , \38628 );
buf \U$30760 ( \38630 , RIb885ec8_40);
and \U$30761 ( \38631 , \38629 , \38630 );
buf \U$30762 ( \38632 , RIb82dcc8_208);
buf \U$30763 ( \38633 , \38632 );
not \U$30764 ( \38634 , \38077 );
and \U$30765 ( \38635 , \38633 , \38634 );
nor \U$30766 ( \38636 , \38631 , \38635 );
nand \U$30767 ( \38637 , \38627 , \38636 );
and \U$30768 ( \38638 , \38637 , \38223 );
or \U$30769 ( \38639 , \38625 , \38638 );
and \U$30771 ( \38640 , \38639 , 1'b1 );
or \U$30773 ( \38641 , \38640 , 1'b0 );
buf \U$30774 ( \38642 , \38641 );
_DC r2379e_GF_IsGateDCbyConstraint ( \38643_nR2379e , \38642 , \21944 );
buf \U$30775 ( \38644 , \38643_nR2379e );
buf \U$30776 ( \38645 , \38033 );
not \U$30777 ( \38646 , \38645 );
and \U$30778 ( \38647 , RIe02ccd8_5323, \38646 );
not \U$30779 ( \38648 , RIe02ccd8_5323);
or \U$30780 ( \38649 , \38648 , \38266 );
buf \U$30781 ( \38650 , \33302 );
and \U$30782 ( \38651 , \38268 , \38650 );
buf \U$30783 ( \38652 , RIb82dd40_207);
buf \U$30784 ( \38653 , \38652 );
not \U$30785 ( \38654 , \38086 );
and \U$30786 ( \38655 , \38653 , \38654 );
nor \U$30787 ( \38656 , \38651 , \38655 );
nand \U$30788 ( \38657 , \38649 , \38656 );
and \U$30789 ( \38658 , \38657 , \38645 );
or \U$30790 ( \38659 , \38647 , \38658 );
and \U$30792 ( \38660 , \38659 , 1'b1 );
or \U$30794 ( \38661 , \38660 , 1'b0 );
buf \U$30795 ( \38662 , \38661 );
_DC r237a2_GF_IsGateDCbyConstraint ( \38663_nR237a2 , \38662 , \21944 );
buf \U$30796 ( \38664 , \38663_nR237a2 );
not \U$30797 ( \38665 , \38645 );
and \U$30798 ( \38666 , RIe0322a0_5324, \38665 );
not \U$30799 ( \38667 , RIe0322a0_5324);
or \U$30800 ( \38668 , \38667 , \38051 );
buf \U$30801 ( \38669 , RIb885fb8_38);
buf \U$30802 ( \38670 , \38669 );
and \U$30803 ( \38671 , \38268 , \38670 );
buf \U$30804 ( \38672 , RIb82ddb8_206);
buf \U$30805 ( \38673 , \38672 );
not \U$30806 ( \38674 , \38407 );
and \U$30807 ( \38675 , \38673 , \38674 );
nor \U$30808 ( \38676 , \38671 , \38675 );
nand \U$30809 ( \38677 , \38668 , \38676 );
and \U$30810 ( \38678 , \38677 , \38645 );
or \U$30811 ( \38679 , \38666 , \38678 );
and \U$30813 ( \38680 , \38679 , 1'b1 );
or \U$30815 ( \38681 , \38680 , 1'b0 );
buf \U$30816 ( \38682 , \38681 );
_DC r237a4_GF_IsGateDCbyConstraint ( \38683_nR237a4 , \38682 , \21944 );
buf \U$30817 ( \38684 , \38683_nR237a4 );
not \U$30818 ( \38685 , \38223 );
and \U$30819 ( \38686 , RIe038768_5325, \38685 );
not \U$30820 ( \38687 , RIe038768_5325);
or \U$30821 ( \38688 , \38687 , \38266 );
buf \U$30822 ( \38689 , RIb886030_37);
buf \U$30823 ( \38690 , \38689 );
and \U$30824 ( \38691 , \38081 , \38690 );
buf \U$30825 ( \38692 , RIb82de30_205);
buf \U$30826 ( \38693 , \38692 );
not \U$30827 ( \38694 , \38231 );
and \U$30828 ( \38695 , \38693 , \38694 );
nor \U$30829 ( \38696 , \38691 , \38695 );
nand \U$30830 ( \38697 , \38688 , \38696 );
and \U$30831 ( \38698 , \38697 , \38223 );
or \U$30832 ( \38699 , \38686 , \38698 );
and \U$30834 ( \38700 , \38699 , 1'b1 );
or \U$30836 ( \38701 , \38700 , 1'b0 );
buf \U$30837 ( \38702 , \38701 );
_DC r237a6_GF_IsGateDCbyConstraint ( \38703_nR237a6 , \38702 , \21944 );
buf \U$30838 ( \38704 , \38703_nR237a6 );
buf \U$30839 ( \38705 , \38032 );
not \U$30840 ( \38706 , \38705 );
and \U$30841 ( \38707 , RIe03c728_5326, \38706 );
not \U$30842 ( \38708 , RIe03c728_5326);
or \U$30843 ( \38709 , \38708 , \38141 );
buf \U$30844 ( \38710 , \22822 );
and \U$30845 ( \38711 , \38268 , \38710 );
buf \U$30846 ( \38712 , RIb832228_204);
buf \U$30847 ( \38713 , \38712 );
not \U$30848 ( \38714 , \38329 );
and \U$30849 ( \38715 , \38713 , \38714 );
nor \U$30850 ( \38716 , \38711 , \38715 );
nand \U$30851 ( \38717 , \38709 , \38716 );
and \U$30852 ( \38718 , \38717 , \38705 );
or \U$30853 ( \38719 , \38707 , \38718 );
and \U$30855 ( \38720 , \38719 , 1'b1 );
or \U$30857 ( \38721 , \38720 , 1'b0 );
buf \U$30858 ( \38722 , \38721 );
_DC r237a8_GF_IsGateDCbyConstraint ( \38723_nR237a8 , \38722 , \21944 );
buf \U$30859 ( \38724 , \38723_nR237a8 );
not \U$30860 ( \38725 , \38645 );
and \U$30861 ( \38726 , RIde01258_5327, \38725 );
not \U$30862 ( \38727 , RIde01258_5327);
or \U$30863 ( \38728 , \38727 , \38305 );
not \U$30864 ( \38729 , \38081 );
not \U$30865 ( \38730 , \38729 );
buf \U$30866 ( \38731 , RIb886120_35);
and \U$30867 ( \38732 , \38730 , \38731 );
buf \U$30868 ( \38733 , RIb8322a0_203);
buf \U$30869 ( \38734 , \38733 );
not \U$30870 ( \38735 , \38171 );
and \U$30871 ( \38736 , \38734 , \38735 );
nor \U$30872 ( \38737 , \38732 , \38736 );
nand \U$30873 ( \38738 , \38728 , \38737 );
and \U$30874 ( \38739 , \38738 , \38645 );
or \U$30875 ( \38740 , \38726 , \38739 );
and \U$30877 ( \38741 , \38740 , 1'b1 );
or \U$30879 ( \38742 , \38741 , 1'b0 );
buf \U$30880 ( \38743 , \38742 );
_DC r237aa_GF_IsGateDCbyConstraint ( \38744_nR237aa , \38743 , \21944 );
buf \U$30881 ( \38745 , \38744_nR237aa );
not \U$30882 ( \38746 , \38223 );
and \U$30883 ( \38747 , RIddfd748_5328, \38746 );
not \U$30884 ( \38748 , RIddfd748_5328);
or \U$30885 ( \38749 , \38748 , \38186 );
not \U$30886 ( \38750 , \38268 );
not \U$30887 ( \38751 , \38750 );
buf \U$30888 ( \38752 , RIb886198_34);
and \U$30889 ( \38753 , \38751 , \38752 );
buf \U$30890 ( \38754 , \22865 );
not \U$30891 ( \38755 , \38171 );
and \U$30892 ( \38756 , \38754 , \38755 );
nor \U$30893 ( \38757 , \38753 , \38756 );
nand \U$30894 ( \38758 , \38749 , \38757 );
and \U$30895 ( \38759 , \38758 , \38223 );
or \U$30896 ( \38760 , \38747 , \38759 );
and \U$30898 ( \38761 , \38760 , 1'b1 );
or \U$30900 ( \38762 , \38761 , 1'b0 );
buf \U$30901 ( \38763 , \38762 );
_DC r237ac_GF_IsGateDCbyConstraint ( \38764_nR237ac , \38763 , \21944 );
buf \U$30902 ( \38765 , \38764_nR237ac );
not \U$30903 ( \38766 , \38645 );
and \U$30904 ( \38767 , RIddf9788_5329, \38766 );
not \U$30905 ( \38768 , RIddf9788_5329);
or \U$30906 ( \38769 , \38768 , \38079 );
not \U$30907 ( \38770 , \38750 );
buf \U$30908 ( \38771 , \22882 );
and \U$30909 ( \38772 , \38770 , \38771 );
buf \U$30910 ( \38773 , \22885 );
not \U$30911 ( \38774 , \38211 );
and \U$30912 ( \38775 , \38773 , \38774 );
nor \U$30913 ( \38776 , \38772 , \38775 );
nand \U$30914 ( \38777 , \38769 , \38776 );
and \U$30915 ( \38778 , \38777 , \38645 );
or \U$30916 ( \38779 , \38767 , \38778 );
and \U$30918 ( \38780 , \38779 , 1'b1 );
or \U$30920 ( \38781 , \38780 , 1'b0 );
buf \U$30921 ( \38782 , \38781 );
_DC r237ae_GF_IsGateDCbyConstraint ( \38783_nR237ae , \38782 , \21944 );
buf \U$30922 ( \38784 , \38783_nR237ae );
not \U$30923 ( \38785 , \38645 );
and \U$30924 ( \38786 , RIddf3d88_5330, \38785 );
not \U$30925 ( \38787 , RIddf3d88_5330);
or \U$30926 ( \38788 , \38787 , \38141 );
buf \U$30927 ( \38789 , \22904 );
and \U$30928 ( \38790 , \38268 , \38789 );
buf \U$30929 ( \38791 , RIb832408_200);
buf \U$30930 ( \38792 , \38791 );
not \U$30931 ( \38793 , \38231 );
and \U$30932 ( \38794 , \38792 , \38793 );
nor \U$30933 ( \38795 , \38790 , \38794 );
nand \U$30934 ( \38796 , \38788 , \38795 );
and \U$30935 ( \38797 , \38796 , \38645 );
or \U$30936 ( \38798 , \38786 , \38797 );
and \U$30938 ( \38799 , \38798 , 1'b1 );
or \U$30940 ( \38800 , \38799 , 1'b0 );
buf \U$30941 ( \38801 , \38800 );
_DC r237b0_GF_IsGateDCbyConstraint ( \38802_nR237b0 , \38801 , \21944 );
buf \U$30942 ( \38803 , \38802_nR237b0 );
not \U$30943 ( \38804 , \38223 );
and \U$30944 ( \38805 , RIdfba228_5331, \38804 );
not \U$30945 ( \38806 , RIdfba228_5331);
or \U$30946 ( \38807 , \38806 , \38305 );
buf \U$30947 ( \38808 , RIb886300_31);
and \U$30948 ( \38809 , \38268 , \38808 );
buf \U$30949 ( \38810 , \22927 );
not \U$30950 ( \38811 , \38329 );
and \U$30951 ( \38812 , \38810 , \38811 );
nor \U$30952 ( \38813 , \38809 , \38812 );
nand \U$30953 ( \38814 , \38807 , \38813 );
and \U$30954 ( \38815 , \38814 , \38223 );
or \U$30955 ( \38816 , \38805 , \38815 );
and \U$30957 ( \38817 , \38816 , 1'b1 );
or \U$30959 ( \38818 , \38817 , 1'b0 );
buf \U$30960 ( \38819 , \38818 );
_DC r237b2_GF_IsGateDCbyConstraint ( \38820_nR237b2 , \38819 , \21944 );
buf \U$30961 ( \38821 , \38820_nR237b2 );
buf \U$30962 ( \38822 , \38032 );
not \U$30963 ( \38823 , \38822 );
and \U$30964 ( \38824 , RIdfb5e30_5332, \38823 );
not \U$30965 ( \38825 , RIdfb5e30_5332);
or \U$30966 ( \38826 , \38825 , \38186 );
buf \U$30967 ( \38827 , RIb886378_30);
and \U$30968 ( \38828 , \38054 , \38827 );
buf \U$30969 ( \38829 , \22947 );
not \U$30970 ( \38830 , \38251 );
and \U$30971 ( \38831 , \38829 , \38830 );
nor \U$30972 ( \38832 , \38828 , \38831 );
nand \U$30973 ( \38833 , \38826 , \38832 );
and \U$30974 ( \38834 , \38833 , \38822 );
or \U$30975 ( \38835 , \38824 , \38834 );
and \U$30977 ( \38836 , \38835 , 1'b1 );
or \U$30979 ( \38837 , \38836 , 1'b0 );
buf \U$30980 ( \38838 , \38837 );
_DC r237b4_GF_IsGateDCbyConstraint ( \38839_nR237b4 , \38838 , \21944 );
buf \U$30981 ( \38840 , \38839_nR237b4 );
not \U$30982 ( \38841 , \38822 );
and \U$30983 ( \38842 , RIdfb2aa0_5333, \38841 );
not \U$30984 ( \38843 , RIdfb2aa0_5333);
or \U$30985 ( \38844 , \38843 , \38121 );
buf \U$30986 ( \38845 , \22964 );
and \U$30987 ( \38846 , \38162 , \38845 );
buf \U$30988 ( \38847 , \28179 );
not \U$30989 ( \38848 , \38251 );
and \U$30990 ( \38849 , \38847 , \38848 );
nor \U$30991 ( \38850 , \38846 , \38849 );
nand \U$30992 ( \38851 , \38844 , \38850 );
and \U$30993 ( \38852 , \38851 , \38822 );
or \U$30994 ( \38853 , \38842 , \38852 );
and \U$30996 ( \38854 , \38853 , 1'b1 );
or \U$30998 ( \38855 , \38854 , 1'b0 );
buf \U$30999 ( \38856 , \38855 );
_DC r237b8_GF_IsGateDCbyConstraint ( \38857_nR237b8 , \38856 , \21944 );
buf \U$31000 ( \38858 , \38857_nR237b8 );
not \U$31001 ( \38859 , \38223 );
and \U$31002 ( \38860 , RIdfaec48_5334, \38859 );
not \U$31003 ( \38861 , RIdfaec48_5334);
or \U$31004 ( \38862 , \38861 , \38160 );
buf \U$31005 ( \38863 , RIb886468_28);
and \U$31006 ( \38864 , \38162 , \38863 );
buf \U$31007 ( \38865 , \28198 );
not \U$31008 ( \38866 , \38077 );
and \U$31009 ( \38867 , \38865 , \38866 );
nor \U$31010 ( \38868 , \38864 , \38867 );
nand \U$31011 ( \38869 , \38862 , \38868 );
and \U$31012 ( \38870 , \38869 , \38223 );
or \U$31013 ( \38871 , \38860 , \38870 );
and \U$31015 ( \38872 , \38871 , 1'b1 );
or \U$31017 ( \38873 , \38872 , 1'b0 );
buf \U$31018 ( \38874 , \38873 );
_DC r237ba_GF_IsGateDCbyConstraint ( \38875_nR237ba , \38874 , \21944 );
buf \U$31019 ( \38876 , \38875_nR237ba );
not \U$31020 ( \38877 , \38705 );
and \U$31021 ( \38878 , RIdfabf48_5335, \38877 );
not \U$31022 ( \38879 , RIdfabf48_5335);
or \U$31023 ( \38880 , \38879 , \38079 );
buf \U$31024 ( \38881 , RIb8864e0_27);
and \U$31025 ( \38882 , \38054 , \38881 );
buf \U$31026 ( \38883 , \28217 );
not \U$31027 ( \38884 , \38211 );
and \U$31028 ( \38885 , \38883 , \38884 );
nor \U$31029 ( \38886 , \38882 , \38885 );
nand \U$31030 ( \38887 , \38880 , \38886 );
and \U$31031 ( \38888 , \38887 , \38705 );
or \U$31032 ( \38889 , \38878 , \38888 );
and \U$31034 ( \38890 , \38889 , 1'b1 );
or \U$31036 ( \38891 , \38890 , 1'b0 );
buf \U$31037 ( \38892 , \38891 );
_DC r237bc_GF_IsGateDCbyConstraint ( \38893_nR237bc , \38892 , \21944 );
buf \U$31038 ( \38894 , \38893_nR237bc );
not \U$31039 ( \38895 , \38645 );
and \U$31040 ( \38896 , RIdfa97e8_5336, \38895 );
not \U$31041 ( \38897 , RIdfa97e8_5336);
or \U$31042 ( \38898 , \38897 , \38121 );
buf \U$31043 ( \38899 , \23022 );
and \U$31044 ( \38900 , \38268 , \38899 );
buf \U$31045 ( \38901 , RIb838498_194);
buf \U$31046 ( \38902 , \38901 );
not \U$31047 ( \38903 , \38049 );
and \U$31048 ( \38904 , \38902 , \38903 );
nor \U$31049 ( \38905 , \38900 , \38904 );
nand \U$31050 ( \38906 , \38898 , \38905 );
and \U$31051 ( \38907 , \38906 , \38645 );
or \U$31052 ( \38908 , \38896 , \38907 );
and \U$31054 ( \38909 , \38908 , 1'b1 );
or \U$31056 ( \38910 , \38909 , 1'b0 );
buf \U$31057 ( \38911 , \38910 );
_DC r237be_GF_IsGateDCbyConstraint ( \38912_nR237be , \38911 , \21944 );
buf \U$31058 ( \38913 , \38912_nR237be );
buf \U$31059 ( \38914 , \38822 );
not \U$31060 ( \38915 , \38914 );
and \U$31061 ( \38916 , RIdfa5e40_5337, \38915 );
not \U$31062 ( \38917 , RIdfa5e40_5337);
or \U$31063 ( \38918 , \38917 , \38051 );
buf \U$31064 ( \38919 , RIb8865d0_25);
and \U$31065 ( \38920 , \38081 , \38919 );
buf \U$31066 ( \38921 , \28256 );
not \U$31067 ( \38922 , \38086 );
and \U$31068 ( \38923 , \38921 , \38922 );
nor \U$31069 ( \38924 , \38920 , \38923 );
nand \U$31070 ( \38925 , \38918 , \38924 );
and \U$31071 ( \38926 , \38925 , \38914 );
or \U$31072 ( \38927 , \38916 , \38926 );
and \U$31074 ( \38928 , \38927 , 1'b1 );
or \U$31076 ( \38929 , \38928 , 1'b0 );
buf \U$31077 ( \38930 , \38929 );
_DC r237c0_GF_IsGateDCbyConstraint ( \38931_nR237c0 , \38930 , \21944 );
buf \U$31078 ( \38932 , \38931_nR237c0 );
not \U$31079 ( \38933 , \38603 );
and \U$31080 ( \38934 , RIdfa2f60_5338, \38933 );
not \U$31081 ( \38935 , RIdfa2f60_5338);
or \U$31082 ( \38936 , \38935 , \38266 );
buf \U$31083 ( \38937 , RIb886648_24);
and \U$31084 ( \38938 , \38162 , \38937 );
buf \U$31085 ( \38939 , RIb838588_192);
buf \U$31086 ( \38940 , \38939 );
not \U$31087 ( \38941 , \38407 );
and \U$31088 ( \38942 , \38940 , \38941 );
nor \U$31089 ( \38943 , \38938 , \38942 );
nand \U$31090 ( \38944 , \38936 , \38943 );
and \U$31091 ( \38945 , \38944 , \38603 );
or \U$31092 ( \38946 , \38934 , \38945 );
and \U$31094 ( \38947 , \38946 , 1'b1 );
or \U$31096 ( \38948 , \38947 , 1'b0 );
buf \U$31097 ( \38949 , \38948 );
_DC r237c2_GF_IsGateDCbyConstraint ( \38950_nR237c2 , \38949 , \21944 );
buf \U$31098 ( \38951 , \38950_nR237c2 );
not \U$31099 ( \38952 , \38645 );
and \U$31100 ( \38953 , RIdf9e4d8_5339, \38952 );
not \U$31101 ( \38954 , RIdf9e4d8_5339);
or \U$31102 ( \38955 , \38954 , \38121 );
buf \U$31103 ( \38956 , RIb8866c0_23);
and \U$31104 ( \38957 , \38162 , \38956 );
buf \U$31105 ( \38958 , \28294 );
not \U$31106 ( \38959 , \38171 );
and \U$31107 ( \38960 , \38958 , \38959 );
nor \U$31108 ( \38961 , \38957 , \38960 );
nand \U$31109 ( \38962 , \38955 , \38961 );
and \U$31110 ( \38963 , \38962 , \38645 );
or \U$31111 ( \38964 , \38953 , \38963 );
and \U$31113 ( \38965 , \38964 , 1'b1 );
or \U$31115 ( \38966 , \38965 , 1'b0 );
buf \U$31116 ( \38967 , \38966 );
_DC r237c4_GF_IsGateDCbyConstraint ( \38968_nR237c4 , \38967 , \21944 );
buf \U$31117 ( \38969 , \38968_nR237c4 );
not \U$31118 ( \38970 , \38914 );
and \U$31119 ( \38971 , RIdf99618_5340, \38970 );
not \U$31120 ( \38972 , RIdf99618_5340);
or \U$31121 ( \38973 , \38972 , \38160 );
buf \U$31122 ( \38974 , \23104 );
and \U$31123 ( \38975 , \38162 , \38974 );
buf \U$31124 ( \38976 , RIb838678_190);
buf \U$31125 ( \38977 , \38976 );
not \U$31126 ( \38978 , \38211 );
and \U$31127 ( \38979 , \38977 , \38978 );
nor \U$31128 ( \38980 , \38975 , \38979 );
nand \U$31129 ( \38981 , \38973 , \38980 );
and \U$31130 ( \38982 , \38981 , \38914 );
or \U$31131 ( \38983 , \38971 , \38982 );
and \U$31133 ( \38984 , \38983 , 1'b1 );
or \U$31135 ( \38985 , \38984 , 1'b0 );
buf \U$31136 ( \38986 , \38985 );
_DC r237c6_GF_IsGateDCbyConstraint ( \38987_nR237c6 , \38986 , \21944 );
buf \U$31137 ( \38988 , \38987_nR237c6 );
not \U$31138 ( \38989 , \38645 );
and \U$31139 ( \38990 , RIdf90f90_5341, \38989 );
not \U$31140 ( \38991 , RIdf90f90_5341);
or \U$31141 ( \38992 , \38991 , \38079 );
buf \U$31142 ( \38993 , RIb8867b0_21);
and \U$31143 ( \38994 , \38054 , \38993 );
buf \U$31144 ( \38995 , \23127 );
not \U$31145 ( \38996 , \38231 );
and \U$31146 ( \38997 , \38995 , \38996 );
nor \U$31147 ( \38998 , \38994 , \38997 );
nand \U$31148 ( \38999 , \38992 , \38998 );
and \U$31149 ( \39000 , \38999 , \38645 );
or \U$31150 ( \39001 , \38990 , \39000 );
and \U$31152 ( \39002 , \39001 , 1'b1 );
or \U$31154 ( \39003 , \39002 , 1'b0 );
buf \U$31155 ( \39004 , \39003 );
_DC r237c8_GF_IsGateDCbyConstraint ( \39005_nR237c8 , \39004 , \21944 );
buf \U$31156 ( \39006 , \39005_nR237c8 );
not \U$31157 ( \39007 , \38645 );
and \U$31158 ( \39008 , RIdf8ae88_5342, \39007 );
not \U$31159 ( \39009 , RIdf8ae88_5342);
or \U$31160 ( \39010 , \39009 , \38079 );
buf \U$31161 ( \39011 , \33667 );
and \U$31162 ( \39012 , \38054 , \39011 );
buf \U$31163 ( \39013 , RIb838768_188);
buf \U$31164 ( \39014 , \39013 );
not \U$31165 ( \39015 , \38049 );
and \U$31166 ( \39016 , \39014 , \39015 );
nor \U$31167 ( \39017 , \39012 , \39016 );
nand \U$31168 ( \39018 , \39010 , \39017 );
and \U$31169 ( \39019 , \39018 , \38645 );
or \U$31170 ( \39020 , \39008 , \39019 );
and \U$31172 ( \39021 , \39020 , 1'b1 );
or \U$31174 ( \39022 , \39021 , 1'b0 );
buf \U$31175 ( \39023 , \39022 );
_DC r237ca_GF_IsGateDCbyConstraint ( \39024_nR237ca , \39023 , \21944 );
buf \U$31176 ( \39025 , \39024_nR237ca );
not \U$31177 ( \39026 , \38914 );
and \U$31178 ( \39027 , RIdf848d0_5343, \39026 );
not \U$31179 ( \39028 , RIdf848d0_5343);
or \U$31180 ( \39029 , \39028 , \38305 );
buf \U$31181 ( \39030 , \23164 );
and \U$31182 ( \39031 , \38162 , \39030 );
buf \U$31183 ( \39032 , RIb8387e0_187);
buf \U$31184 ( \39033 , \39032 );
not \U$31185 ( \39034 , \38231 );
and \U$31186 ( \39035 , \39033 , \39034 );
nor \U$31187 ( \39036 , \39031 , \39035 );
nand \U$31188 ( \39037 , \39029 , \39036 );
and \U$31189 ( \39038 , \39037 , \38914 );
or \U$31190 ( \39039 , \39027 , \39038 );
and \U$31192 ( \39040 , \39039 , 1'b1 );
or \U$31194 ( \39041 , \39040 , 1'b0 );
buf \U$31195 ( \39042 , \39041 );
_DC r237ce_GF_IsGateDCbyConstraint ( \39043_nR237ce , \39042 , \21944 );
buf \U$31196 ( \39044 , \39043_nR237ce );
buf \U$31197 ( \39045 , \38032 );
not \U$31198 ( \39046 , \39045 );
and \U$31199 ( \39047 , RIdf7c248_5344, \39046 );
not \U$31200 ( \39048 , RIdf7c248_5344);
or \U$31201 ( \39049 , \39048 , \38186 );
buf \U$31202 ( \39050 , RIb886918_18);
buf \U$31203 ( \39051 , \39050 );
and \U$31204 ( \39052 , \38162 , \39051 );
buf \U$31205 ( \39053 , RIb838858_186);
buf \U$31206 ( \39054 , \39053 );
not \U$31207 ( \39055 , \38329 );
and \U$31208 ( \39056 , \39054 , \39055 );
nor \U$31209 ( \39057 , \39052 , \39056 );
nand \U$31210 ( \39058 , \39049 , \39057 );
and \U$31211 ( \39059 , \39058 , \39045 );
or \U$31212 ( \39060 , \39047 , \39059 );
and \U$31214 ( \39061 , \39060 , 1'b1 );
or \U$31216 ( \39062 , \39061 , 1'b0 );
buf \U$31217 ( \39063 , \39062 );
_DC r237d0_GF_IsGateDCbyConstraint ( \39064_nR237d0 , \39063 , \21944 );
buf \U$31218 ( \39065 , \39064_nR237d0 );
buf \U$31219 ( \39066 , \38032 );
not \U$31220 ( \39067 , \39066 );
and \U$31221 ( \39068 , RIdf76140_5345, \39067 );
not \U$31222 ( \39069 , RIdf76140_5345);
or \U$31223 ( \39070 , \39069 , \38079 );
buf \U$31224 ( \39071 , \23203 );
and \U$31225 ( \39072 , \38054 , \39071 );
buf \U$31226 ( \39073 , RIb8388d0_185);
buf \U$31227 ( \39074 , \39073 );
not \U$31228 ( \39075 , \38251 );
and \U$31229 ( \39076 , \39074 , \39075 );
nor \U$31230 ( \39077 , \39072 , \39076 );
nand \U$31231 ( \39078 , \39070 , \39077 );
and \U$31232 ( \39079 , \39078 , \39066 );
or \U$31233 ( \39080 , \39068 , \39079 );
and \U$31235 ( \39081 , \39080 , 1'b1 );
or \U$31237 ( \39082 , \39081 , 1'b0 );
buf \U$31238 ( \39083 , \39082 );
_DC r237d2_GF_IsGateDCbyConstraint ( \39084_nR237d2 , \39083 , \21944 );
buf \U$31239 ( \39085 , \39084_nR237d2 );
not \U$31240 ( \39086 , \38914 );
and \U$31241 ( \39087 , RIdc56298_5346, \39086 );
not \U$31242 ( \39088 , RIdc56298_5346);
or \U$31243 ( \39089 , \39088 , \38121 );
buf \U$31244 ( \39090 , RIb886a08_16);
and \U$31245 ( \39091 , \38054 , \39090 );
buf \U$31246 ( \39092 , RIb838948_184);
buf \U$31247 ( \39093 , \39092 );
not \U$31248 ( \39094 , \38077 );
and \U$31249 ( \39095 , \39093 , \39094 );
nor \U$31250 ( \39096 , \39091 , \39095 );
nand \U$31251 ( \39097 , \39089 , \39096 );
and \U$31252 ( \39098 , \39097 , \38914 );
or \U$31253 ( \39099 , \39087 , \39098 );
and \U$31255 ( \39100 , \39099 , 1'b1 );
or \U$31257 ( \39101 , \39100 , 1'b0 );
buf \U$31258 ( \39102 , \39101 );
_DC r237d4_GF_IsGateDCbyConstraint ( \39103_nR237d4 , \39102 , \21944 );
buf \U$31259 ( \39104 , \39103_nR237d4 );
not \U$31260 ( \39105 , \38645 );
and \U$31261 ( \39106 , RIdd75f50_5347, \39105 );
not \U$31262 ( \39107 , RIdd75f50_5347);
or \U$31263 ( \39108 , \39107 , \38160 );
buf \U$31264 ( \39109 , \33762 );
and \U$31265 ( \39110 , \38162 , \39109 );
buf \U$31266 ( \39111 , RIb8389c0_183);
buf \U$31267 ( \39112 , \39111 );
not \U$31268 ( \39113 , \38049 );
and \U$31269 ( \39114 , \39112 , \39113 );
nor \U$31270 ( \39115 , \39110 , \39114 );
nand \U$31271 ( \39116 , \39108 , \39115 );
and \U$31272 ( \39117 , \39116 , \38645 );
or \U$31273 ( \39118 , \39106 , \39117 );
and \U$31275 ( \39119 , \39118 , 1'b1 );
or \U$31277 ( \39120 , \39119 , 1'b0 );
buf \U$31278 ( \39121 , \39120 );
_DC r237d6_GF_IsGateDCbyConstraint ( \39122_nR237d6 , \39121 , \21944 );
buf \U$31279 ( \39123 , \39122_nR237d6 );
not \U$31280 ( \39124 , \38645 );
and \U$31281 ( \39125 , RIdd9d6b8_5348, \39124 );
not \U$31282 ( \39126 , RIdd9d6b8_5348);
or \U$31283 ( \39127 , \39126 , \38051 );
buf \U$31284 ( \39128 , RIb886af8_14);
and \U$31285 ( \39129 , \38268 , \39128 );
buf \U$31286 ( \39130 , RIb838a38_182);
buf \U$31287 ( \39131 , \39130 );
not \U$31288 ( \39132 , \38086 );
and \U$31289 ( \39133 , \39131 , \39132 );
nor \U$31290 ( \39134 , \39129 , \39133 );
nand \U$31291 ( \39135 , \39127 , \39134 );
and \U$31292 ( \39136 , \39135 , \38645 );
or \U$31293 ( \39137 , \39125 , \39136 );
and \U$31295 ( \39138 , \39137 , 1'b1 );
or \U$31297 ( \39139 , \39138 , 1'b0 );
buf \U$31298 ( \39140 , \39139 );
_DC r237d8_GF_IsGateDCbyConstraint ( \39141_nR237d8 , \39140 , \21944 );
buf \U$31299 ( \39142 , \39141_nR237d8 );
not \U$31300 ( \39143 , \38914 );
and \U$31301 ( \39144 , RIdb67180_5349, \39143 );
not \U$31302 ( \39145 , RIdb67180_5349);
or \U$31303 ( \39146 , \39145 , \38266 );
not \U$31304 ( \39147 , \38044 );
buf \U$31305 ( \39148 , \23283 );
and \U$31306 ( \39149 , \39147 , \39148 );
buf \U$31307 ( \39150 , RIb838ab0_181);
buf \U$31308 ( \39151 , \39150 );
not \U$31309 ( \39152 , \38407 );
and \U$31310 ( \39153 , \39151 , \39152 );
nor \U$31311 ( \39154 , \39149 , \39153 );
nand \U$31312 ( \39155 , \39146 , \39154 );
and \U$31313 ( \39156 , \39155 , \38914 );
or \U$31314 ( \39157 , \39144 , \39156 );
and \U$31316 ( \39158 , \39157 , 1'b1 );
or \U$31318 ( \39159 , \39158 , 1'b0 );
buf \U$31319 ( \39160 , \39159 );
_DC r237da_GF_IsGateDCbyConstraint ( \39161_nR237da , \39160 , \21944 );
buf \U$31320 ( \39162 , \39161_nR237da );
buf \U$31321 ( \39163 , \38032 );
not \U$31322 ( \39164 , \39163 );
and \U$31323 ( \39165 , RIdc198c0_5350, \39164 );
not \U$31324 ( \39166 , RIdc198c0_5350);
or \U$31325 ( \39167 , \39166 , \38141 );
buf \U$31326 ( \39168 , RIb886be8_12);
buf \U$31327 ( \39169 , \39168 );
and \U$31328 ( \39170 , \38054 , \39169 );
buf \U$31329 ( \39171 , \23305 );
not \U$31330 ( \39172 , \38407 );
and \U$31331 ( \39173 , \39171 , \39172 );
nor \U$31332 ( \39174 , \39170 , \39173 );
nand \U$31333 ( \39175 , \39167 , \39174 );
and \U$31334 ( \39176 , \39175 , \39163 );
or \U$31335 ( \39177 , \39165 , \39176 );
and \U$31337 ( \39178 , \39177 , 1'b1 );
or \U$31339 ( \39179 , \39178 , 1'b0 );
buf \U$31340 ( \39180 , \39179 );
_DC r237dc_GF_IsGateDCbyConstraint ( \39181_nR237dc , \39180 , \21944 );
buf \U$31341 ( \39182 , \39181_nR237dc );
not \U$31342 ( \39183 , \38645 );
and \U$31343 ( \39184 , RIdc008e8_5351, \39183 );
not \U$31344 ( \39185 , RIdc008e8_5351);
or \U$31345 ( \39186 , \39185 , \38305 );
buf \U$31346 ( \39187 , RIb886c60_11);
buf \U$31347 ( \39188 , \39187 );
and \U$31348 ( \39189 , \38081 , \39188 );
buf \U$31349 ( \39190 , \23325 );
not \U$31350 ( \39191 , \38171 );
and \U$31351 ( \39192 , \39190 , \39191 );
nor \U$31352 ( \39193 , \39189 , \39192 );
nand \U$31353 ( \39194 , \39186 , \39193 );
and \U$31354 ( \39195 , \39194 , \38645 );
or \U$31355 ( \39196 , \39184 , \39195 );
and \U$31357 ( \39197 , \39196 , 1'b1 );
or \U$31359 ( \39198 , \39197 , 1'b0 );
buf \U$31360 ( \39199 , \39198 );
_DC r237de_GF_IsGateDCbyConstraint ( \39200_nR237de , \39199 , \21944 );
buf \U$31361 ( \39201 , \39200_nR237de );
not \U$31362 ( \39202 , \38914 );
and \U$31363 ( \39203 , RIdacdc88_5352, \39202 );
not \U$31364 ( \39204 , RIdacdc88_5352);
or \U$31365 ( \39205 , \39204 , \38079 );
not \U$31366 ( \39206 , \38162 );
not \U$31367 ( \39207 , \39206 );
buf \U$31368 ( \39208 , \28547 );
and \U$31369 ( \39209 , \39207 , \39208 );
buf \U$31370 ( \39210 , RIb838c18_178);
buf \U$31371 ( \39211 , \39210 );
not \U$31372 ( \39212 , \38329 );
and \U$31373 ( \39213 , \39211 , \39212 );
nor \U$31374 ( \39214 , \39209 , \39213 );
nand \U$31375 ( \39215 , \39205 , \39214 );
and \U$31376 ( \39216 , \39215 , \38914 );
or \U$31377 ( \39217 , \39203 , \39216 );
and \U$31379 ( \39218 , \39217 , 1'b1 );
or \U$31381 ( \39219 , \39218 , 1'b0 );
buf \U$31382 ( \39220 , \39219 );
_DC r237e0_GF_IsGateDCbyConstraint ( \39221_nR237e0 , \39220 , \21944 );
buf \U$31383 ( \39222 , \39221_nR237e0 );
not \U$31384 ( \39223 , \38645 );
and \U$31385 ( \39224 , RId8fd180_5353, \39223 );
not \U$31386 ( \39225 , RId8fd180_5353);
or \U$31387 ( \39226 , \39225 , \38051 );
buf \U$31388 ( \39227 , \23363 );
and \U$31389 ( \39228 , \38162 , \39227 );
buf \U$31390 ( \39229 , RIb838c90_177);
buf \U$31391 ( \39230 , \39229 );
not \U$31392 ( \39231 , \38211 );
and \U$31393 ( \39232 , \39230 , \39231 );
nor \U$31394 ( \39233 , \39228 , \39232 );
nand \U$31395 ( \39234 , \39226 , \39233 );
and \U$31396 ( \39235 , \39234 , \38645 );
or \U$31397 ( \39236 , \39224 , \39235 );
and \U$31399 ( \39237 , \39236 , 1'b1 );
or \U$31401 ( \39238 , \39237 , 1'b0 );
buf \U$31402 ( \39239 , \39238 );
_DC r237e4_GF_IsGateDCbyConstraint ( \39240_nR237e4 , \39239 , \21944 );
buf \U$31403 ( \39241 , \39240_nR237e4 );
not \U$31404 ( \39242 , \38645 );
and \U$31405 ( \39243 , RIdb353b0_5354, \39242 );
not \U$31406 ( \39244 , RIdb353b0_5354);
or \U$31407 ( \39245 , \39244 , \38266 );
not \U$31408 ( \39246 , \39206 );
buf \U$31409 ( \39247 , \23383 );
and \U$31410 ( \39248 , \39246 , \39247 );
buf \U$31411 ( \39249 , RIb838d08_176);
buf \U$31412 ( \39250 , \39249 );
not \U$31413 ( \39251 , \38231 );
and \U$31414 ( \39252 , \39250 , \39251 );
nor \U$31415 ( \39253 , \39248 , \39252 );
nand \U$31416 ( \39254 , \39245 , \39253 );
and \U$31417 ( \39255 , \39254 , \38645 );
or \U$31418 ( \39256 , \39243 , \39255 );
and \U$31420 ( \39257 , \39256 , 1'b1 );
or \U$31422 ( \39258 , \39257 , 1'b0 );
buf \U$31423 ( \39259 , \39258 );
_DC r237e6_GF_IsGateDCbyConstraint ( \39260_nR237e6 , \39259 , \21944 );
buf \U$31424 ( \39261 , \39260_nR237e6 );
not \U$31425 ( \39262 , \38914 );
and \U$31426 ( \39263 , RIdbdbca0_5355, \39262 );
not \U$31427 ( \39264 , RIdbdbca0_5355);
or \U$31428 ( \39265 , \39264 , \38141 );
buf \U$31429 ( \39266 , RIb886e40_7);
and \U$31430 ( \39267 , \38162 , \39266 );
buf \U$31431 ( \39268 , RIb838d80_175);
buf \U$31432 ( \39269 , \39268 );
not \U$31433 ( \39270 , \38329 );
and \U$31434 ( \39271 , \39269 , \39270 );
nor \U$31435 ( \39272 , \39267 , \39271 );
nand \U$31436 ( \39273 , \39265 , \39272 );
and \U$31437 ( \39274 , \39273 , \38914 );
or \U$31438 ( \39275 , \39263 , \39274 );
and \U$31440 ( \39276 , \39275 , 1'b1 );
or \U$31442 ( \39277 , \39276 , 1'b0 );
buf \U$31443 ( \39278 , \39277 );
_DC r237e8_GF_IsGateDCbyConstraint ( \39279_nR237e8 , \39278 , \21944 );
buf \U$31444 ( \39280 , \39279_nR237e8 );
not \U$31445 ( \39281 , \39045 );
and \U$31446 ( \39282 , RIdb8b8b8_5356, \39281 );
not \U$31447 ( \39283 , RIdb8b8b8_5356);
or \U$31448 ( \39284 , \39283 , \38305 );
buf \U$31449 ( \39285 , RIb886eb8_6);
and \U$31450 ( \39286 , \38054 , \39285 );
buf \U$31451 ( \39287 , RIb838df8_174);
buf \U$31452 ( \39288 , \39287 );
not \U$31453 ( \39289 , \38251 );
and \U$31454 ( \39290 , \39288 , \39289 );
nor \U$31455 ( \39291 , \39286 , \39290 );
nand \U$31456 ( \39292 , \39284 , \39291 );
and \U$31457 ( \39293 , \39292 , \39045 );
or \U$31458 ( \39294 , \39282 , \39293 );
and \U$31460 ( \39295 , \39294 , 1'b1 );
or \U$31462 ( \39296 , \39295 , 1'b0 );
buf \U$31463 ( \39297 , \39296 );
_DC r237ea_GF_IsGateDCbyConstraint ( \39298_nR237ea , \39297 , \21944 );
buf \U$31464 ( \39299 , \39298_nR237ea );
not \U$31465 ( \39300 , \39066 );
and \U$31466 ( \39301 , RIddb1a28_5357, \39300 );
not \U$31467 ( \39302 , RIddb1a28_5357);
not \U$31468 ( \39303 , \38047 );
nor \U$31469 ( \39304 , \38046 , \39303 );
and \U$31470 ( \39305 , \39304 , \38031 );
not \U$31471 ( \39306 , \38038 );
or \U$31472 ( \39307 , \38039 , \39306 );
not \U$31473 ( \39308 , \39307 );
nand \U$31474 ( \39309 , \38030 , \39308 );
not \U$31475 ( \39310 , \39309 );
or \U$31476 ( \39311 , \39305 , \39310 );
not \U$31477 ( \39312 , \39311 );
not \U$31478 ( \39313 , \39312 );
or \U$31479 ( \39314 , \39302 , \39313 );
not \U$31480 ( \39315 , \39305 );
not \U$31481 ( \39316 , \39315 );
and \U$31482 ( \39317 , \38058 , \39316 );
not \U$31483 ( \39318 , \39317 );
not \U$31484 ( \39319 , \38055 );
not \U$31485 ( \39320 , \39309 );
buf \U$31486 ( \39321 , \39320 );
not \U$31487 ( \39322 , \39321 );
or \U$31488 ( \39323 , \39319 , \39322 );
nand \U$31489 ( \39324 , \39314 , \39318 , \39323 );
and \U$31490 ( \39325 , \39324 , \39066 );
or \U$31491 ( \39326 , \39301 , \39325 );
and \U$31493 ( \39327 , \39326 , 1'b1 );
or \U$31495 ( \39328 , \39327 , 1'b0 );
buf \U$31496 ( \39329 , \39328 );
_DC r237f4_GF_IsGateDCbyConstraint ( \39330_nR237f4 , \39329 , \21944 );
buf \U$31497 ( \39331 , \39330_nR237f4 );
not \U$31498 ( \39332 , \38914 );
and \U$31499 ( \39333 , RIddc60e0_5358, \39332 );
not \U$31500 ( \39334 , RIddc60e0_5358);
not \U$31501 ( \39335 , \39312 );
or \U$31502 ( \39336 , \39334 , \39335 );
not \U$31503 ( \39337 , \39305 );
not \U$31504 ( \39338 , \39337 );
and \U$31505 ( \39339 , \38085 , \39338 );
not \U$31506 ( \39340 , \39339 );
not \U$31507 ( \39341 , \38083 );
buf \U$31508 ( \39342 , \39320 );
not \U$31509 ( \39343 , \39342 );
or \U$31510 ( \39344 , \39341 , \39343 );
nand \U$31511 ( \39345 , \39336 , \39340 , \39344 );
and \U$31512 ( \39346 , \39345 , \38914 );
or \U$31513 ( \39347 , \39333 , \39346 );
and \U$31515 ( \39348 , \39347 , 1'b1 );
or \U$31517 ( \39349 , \39348 , 1'b0 );
buf \U$31518 ( \39350 , \39349 );
_DC r2380a_GF_IsGateDCbyConstraint ( \39351_nR2380a , \39350 , \21944 );
buf \U$31519 ( \39352 , \39351_nR2380a );
not \U$31520 ( \39353 , \39163 );
and \U$31521 ( \39354 , RIddd3cb8_5359, \39353 );
not \U$31522 ( \39355 , RIddd3cb8_5359);
not \U$31523 ( \39356 , \39312 );
or \U$31524 ( \39357 , \39355 , \39356 );
not \U$31525 ( \39358 , \39315 );
and \U$31526 ( \39359 , \38105 , \39358 );
not \U$31527 ( \39360 , \39359 );
not \U$31528 ( \39361 , \38102 );
not \U$31529 ( \39362 , \39321 );
or \U$31530 ( \39363 , \39361 , \39362 );
nand \U$31531 ( \39364 , \39357 , \39360 , \39363 );
and \U$31532 ( \39365 , \39364 , \39163 );
or \U$31533 ( \39366 , \39354 , \39365 );
and \U$31535 ( \39367 , \39366 , 1'b1 );
or \U$31537 ( \39368 , \39367 , 1'b0 );
buf \U$31538 ( \39369 , \39368 );
_DC r23820_GF_IsGateDCbyConstraint ( \39370_nR23820 , \39369 , \21944 );
buf \U$31539 ( \39371 , \39370_nR23820 );
not \U$31540 ( \39372 , \39045 );
and \U$31541 ( \39373 , RIdddeaa0_5360, \39372 );
not \U$31542 ( \39374 , RIdddeaa0_5360);
not \U$31543 ( \39375 , \39312 );
or \U$31544 ( \39376 , \39374 , \39375 );
not \U$31545 ( \39377 , \39305 );
not \U$31546 ( \39378 , \39377 );
and \U$31547 ( \39379 , \38126 , \39378 );
not \U$31548 ( \39380 , \39379 );
not \U$31549 ( \39381 , \38123 );
not \U$31550 ( \39382 , \39342 );
or \U$31551 ( \39383 , \39381 , \39382 );
nand \U$31552 ( \39384 , \39376 , \39380 , \39383 );
and \U$31553 ( \39385 , \39384 , \39045 );
or \U$31554 ( \39386 , \39373 , \39385 );
and \U$31556 ( \39387 , \39386 , 1'b1 );
or \U$31558 ( \39388 , \39387 , 1'b0 );
buf \U$31559 ( \39389 , \39388 );
_DC r23836_GF_IsGateDCbyConstraint ( \39390_nR23836 , \39389 , \21944 );
buf \U$31560 ( \39391 , \39390_nR23836 );
not \U$31561 ( \39392 , \38914 );
and \U$31562 ( \39393 , RIdde50d0_5361, \39392 );
not \U$31563 ( \39394 , RIdde50d0_5361);
or \U$31564 ( \39395 , \39394 , \39375 );
not \U$31565 ( \39396 , \39315 );
and \U$31566 ( \39397 , \38145 , \39396 );
not \U$31567 ( \39398 , \39397 );
not \U$31568 ( \39399 , \38143 );
buf \U$31569 ( \39400 , \39320 );
not \U$31570 ( \39401 , \39400 );
or \U$31571 ( \39402 , \39399 , \39401 );
nand \U$31572 ( \39403 , \39395 , \39398 , \39402 );
and \U$31573 ( \39404 , \39403 , \38914 );
or \U$31574 ( \39405 , \39393 , \39404 );
and \U$31576 ( \39406 , \39405 , 1'b1 );
or \U$31578 ( \39407 , \39406 , 1'b0 );
buf \U$31579 ( \39408 , \39407 );
_DC r2384c_GF_IsGateDCbyConstraint ( \39409_nR2384c , \39408 , \21944 );
buf \U$31580 ( \39410 , \39409_nR2384c );
buf \U$31581 ( \39411 , \38032 );
not \U$31582 ( \39412 , \39411 );
and \U$31583 ( \39413 , RIddeee50_5362, \39412 );
not \U$31584 ( \39414 , RIddeee50_5362);
or \U$31585 ( \39415 , \39414 , \39375 );
not \U$31586 ( \39416 , \39315 );
and \U$31587 ( \39417 , \38166 , \39416 );
not \U$31588 ( \39418 , \39417 );
not \U$31589 ( \39419 , \38163 );
not \U$31590 ( \39420 , \39342 );
or \U$31591 ( \39421 , \39419 , \39420 );
nand \U$31592 ( \39422 , \39415 , \39418 , \39421 );
and \U$31593 ( \39423 , \39422 , \39411 );
or \U$31594 ( \39424 , \39413 , \39423 );
and \U$31596 ( \39425 , \39424 , 1'b1 );
or \U$31598 ( \39426 , \39425 , 1'b0 );
buf \U$31599 ( \39427 , \39426 );
_DC r23862_GF_IsGateDCbyConstraint ( \39428_nR23862 , \39427 , \21944 );
buf \U$31600 ( \39429 , \39428_nR23862 );
not \U$31601 ( \39430 , \39411 );
and \U$31602 ( \39431 , RIdc2bb60_5363, \39430 );
not \U$31603 ( \39432 , RIdc2bb60_5363);
or \U$31604 ( \39433 , \39432 , \39335 );
not \U$31605 ( \39434 , \39305 );
not \U$31606 ( \39435 , \39434 );
and \U$31607 ( \39436 , \38191 , \39435 );
not \U$31608 ( \39437 , \39436 );
not \U$31609 ( \39438 , \38188 );
not \U$31610 ( \39439 , \39400 );
or \U$31611 ( \39440 , \39438 , \39439 );
nand \U$31612 ( \39441 , \39433 , \39437 , \39440 );
and \U$31613 ( \39442 , \39441 , \39411 );
or \U$31614 ( \39443 , \39431 , \39442 );
and \U$31616 ( \39444 , \39443 , 1'b1 );
or \U$31618 ( \39445 , \39444 , 1'b0 );
buf \U$31619 ( \39446 , \39445 );
_DC r2386c_GF_IsGateDCbyConstraint ( \39447_nR2386c , \39446 , \21944 );
buf \U$31620 ( \39448 , \39447_nR2386c );
not \U$31621 ( \39449 , \38914 );
and \U$31622 ( \39450 , RIdc34788_5364, \39449 );
not \U$31623 ( \39451 , RIdc34788_5364);
or \U$31624 ( \39452 , \39451 , \39375 );
not \U$31625 ( \39453 , \39377 );
and \U$31626 ( \39454 , \38210 , \39453 );
not \U$31627 ( \39455 , \39454 );
not \U$31628 ( \39456 , \38207 );
not \U$31629 ( \39457 , \39342 );
or \U$31630 ( \39458 , \39456 , \39457 );
nand \U$31631 ( \39459 , \39452 , \39455 , \39458 );
and \U$31632 ( \39460 , \39459 , \38914 );
or \U$31633 ( \39461 , \39450 , \39460 );
and \U$31635 ( \39462 , \39461 , 1'b1 );
or \U$31637 ( \39463 , \39462 , 1'b0 );
buf \U$31638 ( \39464 , \39463 );
_DC r2386e_GF_IsGateDCbyConstraint ( \39465_nR2386e , \39464 , \21944 );
buf \U$31639 ( \39466 , \39465_nR2386e );
not \U$31640 ( \39467 , \38645 );
and \U$31641 ( \39468 , RIde6e7b8_5365, \39467 );
not \U$31642 ( \39469 , RIde6e7b8_5365);
or \U$31643 ( \39470 , \39469 , \39313 );
not \U$31644 ( \39471 , \39337 );
and \U$31645 ( \39472 , \38230 , \39471 );
not \U$31646 ( \39473 , \39472 );
not \U$31647 ( \39474 , \38228 );
not \U$31648 ( \39475 , \39400 );
or \U$31649 ( \39476 , \39474 , \39475 );
nand \U$31650 ( \39477 , \39470 , \39473 , \39476 );
and \U$31651 ( \39478 , \39477 , \38645 );
or \U$31652 ( \39479 , \39468 , \39478 );
and \U$31654 ( \39480 , \39479 , 1'b1 );
or \U$31656 ( \39481 , \39480 , 1'b0 );
buf \U$31657 ( \39482 , \39481 );
_DC r23870_GF_IsGateDCbyConstraint ( \39483_nR23870 , \39482 , \21944 );
buf \U$31658 ( \39484 , \39483_nR23870 );
not \U$31659 ( \39485 , \39066 );
and \U$31660 ( \39486 , RIde62ad0_5366, \39485 );
not \U$31661 ( \39487 , RIde62ad0_5366);
or \U$31662 ( \39488 , \39487 , \39313 );
not \U$31663 ( \39489 , \39337 );
and \U$31664 ( \39490 , \38250 , \39489 );
not \U$31665 ( \39491 , \39490 );
not \U$31666 ( \39492 , \38247 );
not \U$31667 ( \39493 , \39400 );
or \U$31668 ( \39494 , \39492 , \39493 );
nand \U$31669 ( \39495 , \39488 , \39491 , \39494 );
and \U$31670 ( \39496 , \39495 , \39066 );
or \U$31671 ( \39497 , \39486 , \39496 );
and \U$31673 ( \39498 , \39497 , 1'b1 );
or \U$31675 ( \39499 , \39498 , 1'b0 );
buf \U$31676 ( \39500 , \39499 );
_DC r23872_GF_IsGateDCbyConstraint ( \39501_nR23872 , \39500 , \21944 );
buf \U$31677 ( \39502 , \39501_nR23872 );
not \U$31678 ( \39503 , \38914 );
and \U$31679 ( \39504 , RIde55510_5367, \39503 );
not \U$31680 ( \39505 , RIde55510_5367);
not \U$31681 ( \39506 , \39312 );
or \U$31682 ( \39507 , \39505 , \39506 );
not \U$31683 ( \39508 , \39315 );
and \U$31684 ( \39509 , \38271 , \39508 );
not \U$31685 ( \39510 , \39509 );
not \U$31686 ( \39511 , \38269 );
not \U$31687 ( \39512 , \39321 );
or \U$31688 ( \39513 , \39511 , \39512 );
nand \U$31689 ( \39514 , \39507 , \39510 , \39513 );
and \U$31690 ( \39515 , \39514 , \38914 );
or \U$31691 ( \39516 , \39504 , \39515 );
and \U$31693 ( \39517 , \39516 , 1'b1 );
or \U$31695 ( \39518 , \39517 , 1'b0 );
buf \U$31696 ( \39519 , \39518 );
_DC r237f6_GF_IsGateDCbyConstraint ( \39520_nR237f6 , \39519 , \21944 );
buf \U$31697 ( \39521 , \39520_nR237f6 );
not \U$31698 ( \39522 , \38822 );
and \U$31699 ( \39523 , RIde4a188_5368, \39522 );
not \U$31700 ( \39524 , RIde4a188_5368);
or \U$31701 ( \39525 , \39524 , \39335 );
not \U$31702 ( \39526 , \39337 );
and \U$31703 ( \39527 , \38290 , \39526 );
not \U$31704 ( \39528 , \39527 );
not \U$31705 ( \39529 , \38287 );
not \U$31706 ( \39530 , \39321 );
or \U$31707 ( \39531 , \39529 , \39530 );
nand \U$31708 ( \39532 , \39525 , \39528 , \39531 );
and \U$31709 ( \39533 , \39532 , \38822 );
or \U$31710 ( \39534 , \39523 , \39533 );
and \U$31712 ( \39535 , \39534 , 1'b1 );
or \U$31714 ( \39536 , \39535 , 1'b0 );
buf \U$31715 ( \39537 , \39536 );
_DC r237f8_GF_IsGateDCbyConstraint ( \39538_nR237f8 , \39537 , \21944 );
buf \U$31716 ( \39539 , \39538_nR237f8 );
not \U$31717 ( \39540 , \38822 );
and \U$31718 ( \39541 , RIde36d90_5369, \39540 );
not \U$31719 ( \39542 , RIde36d90_5369);
or \U$31720 ( \39543 , \39542 , \39335 );
not \U$31721 ( \39544 , \39315 );
and \U$31722 ( \39545 , \38309 , \39544 );
not \U$31723 ( \39546 , \39545 );
not \U$31724 ( \39547 , \38307 );
not \U$31725 ( \39548 , \39321 );
or \U$31726 ( \39549 , \39547 , \39548 );
nand \U$31727 ( \39550 , \39543 , \39546 , \39549 );
and \U$31728 ( \39551 , \39550 , \38822 );
or \U$31729 ( \39552 , \39541 , \39551 );
and \U$31731 ( \39553 , \39552 , 1'b1 );
or \U$31733 ( \39554 , \39553 , 1'b0 );
buf \U$31734 ( \39555 , \39554 );
_DC r237fa_GF_IsGateDCbyConstraint ( \39556_nR237fa , \39555 , \21944 );
buf \U$31735 ( \39557 , \39556_nR237fa );
not \U$31736 ( \39558 , \38914 );
and \U$31737 ( \39559 , RIde29c80_5370, \39558 );
not \U$31738 ( \39560 , RIde29c80_5370);
or \U$31739 ( \39561 , \39560 , \39335 );
not \U$31740 ( \39562 , \39315 );
and \U$31741 ( \39563 , \38328 , \39562 );
not \U$31742 ( \39564 , \39563 );
not \U$31743 ( \39565 , \38325 );
not \U$31744 ( \39566 , \39321 );
or \U$31745 ( \39567 , \39565 , \39566 );
nand \U$31746 ( \39568 , \39561 , \39564 , \39567 );
and \U$31747 ( \39569 , \39568 , \38914 );
or \U$31748 ( \39570 , \39559 , \39569 );
and \U$31750 ( \39571 , \39570 , 1'b1 );
or \U$31752 ( \39572 , \39571 , 1'b0 );
buf \U$31753 ( \39573 , \39572 );
_DC r237fc_GF_IsGateDCbyConstraint ( \39574_nR237fc , \39573 , \21944 );
buf \U$31754 ( \39575 , \39574_nR237fc );
not \U$31755 ( \39576 , \39066 );
and \U$31756 ( \39577 , RIde1c210_5371, \39576 );
not \U$31757 ( \39578 , RIde1c210_5371);
or \U$31758 ( \39579 , \39578 , \39313 );
not \U$31759 ( \39580 , \39337 );
and \U$31760 ( \39581 , \38349 , \39580 );
not \U$31761 ( \39582 , \39581 );
not \U$31762 ( \39583 , \38346 );
not \U$31763 ( \39584 , \39321 );
or \U$31764 ( \39585 , \39583 , \39584 );
nand \U$31765 ( \39586 , \39579 , \39582 , \39585 );
and \U$31766 ( \39587 , \39586 , \39066 );
or \U$31767 ( \39588 , \39577 , \39587 );
and \U$31769 ( \39589 , \39588 , 1'b1 );
or \U$31771 ( \39590 , \39589 , 1'b0 );
buf \U$31772 ( \39591 , \39590 );
_DC r237fe_GF_IsGateDCbyConstraint ( \39592_nR237fe , \39591 , \21944 );
buf \U$31773 ( \39593 , \39592_nR237fe );
not \U$31774 ( \39594 , \38645 );
and \U$31775 ( \39595 , RIde0cb08_5372, \39594 );
not \U$31776 ( \39596 , RIde0cb08_5372);
or \U$31777 ( \39597 , \39596 , \39313 );
not \U$31778 ( \39598 , \39315 );
and \U$31779 ( \39599 , \38368 , \39598 );
not \U$31780 ( \39600 , \39599 );
not \U$31781 ( \39601 , \38365 );
not \U$31782 ( \39602 , \39400 );
or \U$31783 ( \39603 , \39601 , \39602 );
nand \U$31784 ( \39604 , \39597 , \39600 , \39603 );
and \U$31785 ( \39605 , \39604 , \38645 );
or \U$31786 ( \39606 , \39595 , \39605 );
and \U$31788 ( \39607 , \39606 , 1'b1 );
or \U$31790 ( \39608 , \39607 , 1'b0 );
buf \U$31791 ( \39609 , \39608 );
_DC r23800_GF_IsGateDCbyConstraint ( \39610_nR23800 , \39609 , \21944 );
buf \U$31792 ( \39611 , \39610_nR23800 );
not \U$31793 ( \39612 , \39411 );
and \U$31794 ( \39613 , RIe03d4c0_5373, \39612 );
not \U$31795 ( \39614 , RIe03d4c0_5373);
or \U$31796 ( \39615 , \39614 , \39506 );
not \U$31797 ( \39616 , \39315 );
and \U$31798 ( \39617 , \38387 , \39616 );
not \U$31799 ( \39618 , \39617 );
not \U$31800 ( \39619 , \38384 );
not \U$31801 ( \39620 , \39400 );
or \U$31802 ( \39621 , \39619 , \39620 );
nand \U$31803 ( \39622 , \39615 , \39618 , \39621 );
and \U$31804 ( \39623 , \39622 , \39411 );
or \U$31805 ( \39624 , \39613 , \39623 );
and \U$31807 ( \39625 , \39624 , 1'b1 );
or \U$31809 ( \39626 , \39625 , 1'b0 );
buf \U$31810 ( \39627 , \39626 );
_DC r23802_GF_IsGateDCbyConstraint ( \39628_nR23802 , \39627 , \21944 );
buf \U$31811 ( \39629 , \39628_nR23802 );
not \U$31812 ( \39630 , \38705 );
and \U$31813 ( \39631 , RIe040b98_5374, \39630 );
not \U$31814 ( \39632 , RIe040b98_5374);
or \U$31815 ( \39633 , \39632 , \39335 );
not \U$31816 ( \39634 , \39434 );
and \U$31817 ( \39635 , \38406 , \39634 );
not \U$31818 ( \39636 , \39635 );
not \U$31819 ( \39637 , \38403 );
not \U$31820 ( \39638 , \39320 );
or \U$31821 ( \39639 , \39637 , \39638 );
nand \U$31822 ( \39640 , \39633 , \39636 , \39639 );
and \U$31823 ( \39641 , \39640 , \38705 );
or \U$31824 ( \39642 , \39631 , \39641 );
and \U$31826 ( \39643 , \39642 , 1'b1 );
or \U$31828 ( \39644 , \39643 , 1'b0 );
buf \U$31829 ( \39645 , \39644 );
_DC r23804_GF_IsGateDCbyConstraint ( \39646_nR23804 , \39645 , \21944 );
buf \U$31830 ( \39647 , \39646_nR23804 );
not \U$31831 ( \39648 , \38117 );
and \U$31832 ( \39649 , RIe043460_5375, \39648 );
not \U$31833 ( \39650 , RIe043460_5375);
or \U$31834 ( \39651 , \39650 , \39356 );
not \U$31835 ( \39652 , \39337 );
and \U$31836 ( \39653 , \38425 , \39652 );
not \U$31837 ( \39654 , \39653 );
not \U$31838 ( \39655 , \38423 );
not \U$31839 ( \39656 , \39400 );
or \U$31840 ( \39657 , \39655 , \39656 );
nand \U$31841 ( \39658 , \39651 , \39654 , \39657 );
and \U$31842 ( \39659 , \39658 , \38117 );
or \U$31843 ( \39660 , \39649 , \39659 );
and \U$31845 ( \39661 , \39660 , 1'b1 );
or \U$31847 ( \39662 , \39661 , 1'b0 );
buf \U$31848 ( \39663 , \39662 );
_DC r23806_GF_IsGateDCbyConstraint ( \39664_nR23806 , \39663 , \21944 );
buf \U$31849 ( \39665 , \39664_nR23806 );
not \U$31850 ( \39666 , \39163 );
and \U$31851 ( \39667 , RIe046b38_5376, \39666 );
not \U$31852 ( \39668 , RIe046b38_5376);
or \U$31853 ( \39669 , \39668 , \39375 );
not \U$31854 ( \39670 , \39434 );
and \U$31855 ( \39671 , \38443 , \39670 );
not \U$31856 ( \39672 , \39671 );
not \U$31857 ( \39673 , \38441 );
not \U$31858 ( \39674 , \39321 );
or \U$31859 ( \39675 , \39673 , \39674 );
nand \U$31860 ( \39676 , \39669 , \39672 , \39675 );
and \U$31861 ( \39677 , \39676 , \39163 );
or \U$31862 ( \39678 , \39667 , \39677 );
and \U$31864 ( \39679 , \39678 , 1'b1 );
or \U$31866 ( \39680 , \39679 , 1'b0 );
buf \U$31867 ( \39681 , \39680 );
_DC r23808_GF_IsGateDCbyConstraint ( \39682_nR23808 , \39681 , \21944 );
buf \U$31868 ( \39683 , \39682_nR23808 );
not \U$31869 ( \39684 , \38117 );
and \U$31870 ( \39685 , RIe049400_5377, \39684 );
not \U$31871 ( \39686 , RIe049400_5377);
or \U$31872 ( \39687 , \39686 , \39313 );
not \U$31873 ( \39688 , \39337 );
and \U$31874 ( \39689 , \38462 , \39688 );
not \U$31875 ( \39690 , \39689 );
not \U$31876 ( \39691 , \38459 );
not \U$31877 ( \39692 , \39320 );
or \U$31878 ( \39693 , \39691 , \39692 );
nand \U$31879 ( \39694 , \39687 , \39690 , \39693 );
and \U$31880 ( \39695 , \39694 , \38117 );
or \U$31881 ( \39696 , \39685 , \39695 );
and \U$31883 ( \39697 , \39696 , 1'b1 );
or \U$31885 ( \39698 , \39697 , 1'b0 );
buf \U$31886 ( \39699 , \39698 );
_DC r2380c_GF_IsGateDCbyConstraint ( \39700_nR2380c , \39699 , \21944 );
buf \U$31887 ( \39701 , \39700_nR2380c );
not \U$31888 ( \39702 , \38117 );
and \U$31889 ( \39703 , RIe04c178_5378, \39702 );
not \U$31890 ( \39704 , RIe04c178_5378);
or \U$31891 ( \39705 , \39704 , \39356 );
not \U$31892 ( \39706 , \39434 );
and \U$31893 ( \39707 , \38481 , \39706 );
not \U$31894 ( \39708 , \39707 );
not \U$31895 ( \39709 , \38478 );
not \U$31896 ( \39710 , \39342 );
or \U$31897 ( \39711 , \39709 , \39710 );
nand \U$31898 ( \39712 , \39705 , \39708 , \39711 );
and \U$31899 ( \39713 , \39712 , \38117 );
or \U$31900 ( \39714 , \39703 , \39713 );
and \U$31902 ( \39715 , \39714 , 1'b1 );
or \U$31904 ( \39716 , \39715 , 1'b0 );
buf \U$31905 ( \39717 , \39716 );
_DC r2380e_GF_IsGateDCbyConstraint ( \39718_nR2380e , \39717 , \21944 );
buf \U$31906 ( \39719 , \39718_nR2380e );
not \U$31907 ( \39720 , \38603 );
and \U$31908 ( \39721 , RIe04f3a0_5379, \39720 );
not \U$31909 ( \39722 , RIe04f3a0_5379);
or \U$31910 ( \39723 , \39722 , \39506 );
not \U$31911 ( \39724 , \39337 );
and \U$31912 ( \39725 , \38500 , \39724 );
not \U$31913 ( \39726 , \39725 );
not \U$31914 ( \39727 , \38497 );
not \U$31915 ( \39728 , \39321 );
or \U$31916 ( \39729 , \39727 , \39728 );
nand \U$31917 ( \39730 , \39723 , \39726 , \39729 );
and \U$31918 ( \39731 , \39730 , \38603 );
or \U$31919 ( \39732 , \39721 , \39731 );
and \U$31921 ( \39733 , \39732 , 1'b1 );
or \U$31923 ( \39734 , \39733 , 1'b0 );
buf \U$31924 ( \39735 , \39734 );
_DC r23810_GF_IsGateDCbyConstraint ( \39736_nR23810 , \39735 , \21944 );
buf \U$31925 ( \39737 , \39736_nR23810 );
not \U$31926 ( \39738 , \39411 );
and \U$31927 ( \39739 , RIe052118_5380, \39738 );
not \U$31928 ( \39740 , RIe052118_5380);
or \U$31929 ( \39741 , \39740 , \39506 );
not \U$31930 ( \39742 , \39377 );
and \U$31931 ( \39743 , \38518 , \39742 );
not \U$31932 ( \39744 , \39743 );
not \U$31933 ( \39745 , \38516 );
not \U$31934 ( \39746 , \39342 );
or \U$31935 ( \39747 , \39745 , \39746 );
nand \U$31936 ( \39748 , \39741 , \39744 , \39747 );
and \U$31937 ( \39749 , \39748 , \39411 );
or \U$31938 ( \39750 , \39739 , \39749 );
and \U$31940 ( \39751 , \39750 , 1'b1 );
or \U$31942 ( \39752 , \39751 , 1'b0 );
buf \U$31943 ( \39753 , \39752 );
_DC r23812_GF_IsGateDCbyConstraint ( \39754_nR23812 , \39753 , \21944 );
buf \U$31944 ( \39755 , \39754_nR23812 );
not \U$31945 ( \39756 , \38603 );
and \U$31946 ( \39757 , RIe055340_5381, \39756 );
not \U$31947 ( \39758 , RIe055340_5381);
or \U$31948 ( \39759 , \39758 , \39375 );
not \U$31949 ( \39760 , \39337 );
and \U$31950 ( \39761 , \38537 , \39760 );
not \U$31951 ( \39762 , \39761 );
not \U$31952 ( \39763 , \38534 );
not \U$31953 ( \39764 , \39320 );
or \U$31954 ( \39765 , \39763 , \39764 );
nand \U$31955 ( \39766 , \39759 , \39762 , \39765 );
and \U$31956 ( \39767 , \39766 , \38603 );
or \U$31957 ( \39768 , \39757 , \39767 );
and \U$31959 ( \39769 , \39768 , 1'b1 );
or \U$31961 ( \39770 , \39769 , 1'b0 );
buf \U$31962 ( \39771 , \39770 );
_DC r23814_GF_IsGateDCbyConstraint ( \39772_nR23814 , \39771 , \21944 );
buf \U$31963 ( \39773 , \39772_nR23814 );
not \U$31964 ( \39774 , \38033 );
and \U$31965 ( \39775 , RIe0580b8_5382, \39774 );
not \U$31966 ( \39776 , RIe0580b8_5382);
or \U$31967 ( \39777 , \39776 , \39506 );
not \U$31968 ( \39778 , \39337 );
and \U$31969 ( \39779 , \38555 , \39778 );
not \U$31970 ( \39780 , \39779 );
not \U$31971 ( \39781 , \38553 );
not \U$31972 ( \39782 , \39342 );
or \U$31973 ( \39783 , \39781 , \39782 );
nand \U$31974 ( \39784 , \39777 , \39780 , \39783 );
and \U$31975 ( \39785 , \39784 , \38033 );
or \U$31976 ( \39786 , \39775 , \39785 );
and \U$31978 ( \39787 , \39786 , 1'b1 );
or \U$31980 ( \39788 , \39787 , 1'b0 );
buf \U$31981 ( \39789 , \39788 );
_DC r23816_GF_IsGateDCbyConstraint ( \39790_nR23816 , \39789 , \21944 );
buf \U$31982 ( \39791 , \39790_nR23816 );
not \U$31983 ( \39792 , \39411 );
and \U$31984 ( \39793 , RIe05b2e0_5383, \39792 );
not \U$31985 ( \39794 , RIe05b2e0_5383);
or \U$31986 ( \39795 , \39794 , \39356 );
not \U$31987 ( \39796 , \39377 );
and \U$31988 ( \39797 , \38573 , \39796 );
not \U$31989 ( \39798 , \39797 );
not \U$31990 ( \39799 , \38571 );
not \U$31991 ( \39800 , \39320 );
or \U$31992 ( \39801 , \39799 , \39800 );
nand \U$31993 ( \39802 , \39795 , \39798 , \39801 );
and \U$31994 ( \39803 , \39802 , \39411 );
or \U$31995 ( \39804 , \39793 , \39803 );
and \U$31997 ( \39805 , \39804 , 1'b1 );
or \U$31999 ( \39806 , \39805 , 1'b0 );
buf \U$32000 ( \39807 , \39806 );
_DC r23818_GF_IsGateDCbyConstraint ( \39808_nR23818 , \39807 , \21944 );
buf \U$32001 ( \39809 , \39808_nR23818 );
not \U$32002 ( \39810 , \38117 );
and \U$32003 ( \39811 , RIe05e058_5384, \39810 );
not \U$32004 ( \39812 , RIe05e058_5384);
or \U$32005 ( \39813 , \39812 , \39375 );
not \U$32006 ( \39814 , \39377 );
and \U$32007 ( \39815 , \38591 , \39814 );
not \U$32008 ( \39816 , \39815 );
not \U$32009 ( \39817 , \38589 );
not \U$32010 ( \39818 , \39342 );
or \U$32011 ( \39819 , \39817 , \39818 );
nand \U$32012 ( \39820 , \39813 , \39816 , \39819 );
and \U$32013 ( \39821 , \39820 , \38117 );
or \U$32014 ( \39822 , \39811 , \39821 );
and \U$32016 ( \39823 , \39822 , 1'b1 );
or \U$32018 ( \39824 , \39823 , 1'b0 );
buf \U$32019 ( \39825 , \39824 );
_DC r2381a_GF_IsGateDCbyConstraint ( \39826_nR2381a , \39825 , \21944 );
buf \U$32020 ( \39827 , \39826_nR2381a );
not \U$32021 ( \39828 , \38822 );
and \U$32022 ( \39829 , RIe060920_5385, \39828 );
not \U$32023 ( \39830 , RIe060920_5385);
or \U$32024 ( \39831 , \39830 , \39356 );
not \U$32025 ( \39832 , \39337 );
and \U$32026 ( \39833 , \38612 , \39832 );
not \U$32027 ( \39834 , \39833 );
not \U$32028 ( \39835 , \38609 );
not \U$32029 ( \39836 , \39321 );
or \U$32030 ( \39837 , \39835 , \39836 );
nand \U$32031 ( \39838 , \39831 , \39834 , \39837 );
and \U$32032 ( \39839 , \39838 , \38822 );
or \U$32033 ( \39840 , \39829 , \39839 );
and \U$32035 ( \39841 , \39840 , 1'b1 );
or \U$32037 ( \39842 , \39841 , 1'b0 );
buf \U$32038 ( \39843 , \39842 );
_DC r2381c_GF_IsGateDCbyConstraint ( \39844_nR2381c , \39843 , \21944 );
buf \U$32039 ( \39845 , \39844_nR2381c );
not \U$32040 ( \39846 , \38705 );
and \U$32041 ( \39847 , RIe063ff8_5386, \39846 );
not \U$32042 ( \39848 , RIe063ff8_5386);
or \U$32043 ( \39849 , \39848 , \39375 );
not \U$32044 ( \39850 , \39377 );
and \U$32045 ( \39851 , \38633 , \39850 );
not \U$32046 ( \39852 , \39851 );
not \U$32047 ( \39853 , \38630 );
not \U$32048 ( \39854 , \39321 );
or \U$32049 ( \39855 , \39853 , \39854 );
nand \U$32050 ( \39856 , \39849 , \39852 , \39855 );
and \U$32051 ( \39857 , \39856 , \38705 );
or \U$32052 ( \39858 , \39847 , \39857 );
and \U$32054 ( \39859 , \39858 , 1'b1 );
or \U$32056 ( \39860 , \39859 , 1'b0 );
buf \U$32057 ( \39861 , \39860 );
_DC r2381e_GF_IsGateDCbyConstraint ( \39862_nR2381e , \39861 , \21944 );
buf \U$32058 ( \39863 , \39862_nR2381e );
not \U$32059 ( \39864 , \39411 );
and \U$32060 ( \39865 , RIe0662a8_5387, \39864 );
not \U$32061 ( \39866 , RIe0662a8_5387);
or \U$32062 ( \39867 , \39866 , \39506 );
not \U$32063 ( \39868 , \39377 );
and \U$32064 ( \39869 , \38653 , \39868 );
not \U$32065 ( \39870 , \39869 );
not \U$32066 ( \39871 , \38650 );
not \U$32067 ( \39872 , \39320 );
or \U$32068 ( \39873 , \39871 , \39872 );
nand \U$32069 ( \39874 , \39867 , \39870 , \39873 );
and \U$32070 ( \39875 , \39874 , \39411 );
or \U$32071 ( \39876 , \39865 , \39875 );
and \U$32073 ( \39877 , \39876 , 1'b1 );
or \U$32075 ( \39878 , \39877 , 1'b0 );
buf \U$32076 ( \39879 , \39878 );
_DC r23822_GF_IsGateDCbyConstraint ( \39880_nR23822 , \39879 , \21944 );
buf \U$32077 ( \39881 , \39880_nR23822 );
not \U$32078 ( \39882 , \38822 );
and \U$32079 ( \39883 , RIe068288_5388, \39882 );
not \U$32080 ( \39884 , RIe068288_5388);
or \U$32081 ( \39885 , \39884 , \39335 );
not \U$32082 ( \39886 , \39315 );
and \U$32083 ( \39887 , \38673 , \39886 );
not \U$32084 ( \39888 , \39887 );
not \U$32085 ( \39889 , \38670 );
not \U$32086 ( \39890 , \39320 );
or \U$32087 ( \39891 , \39889 , \39890 );
nand \U$32088 ( \39892 , \39885 , \39888 , \39891 );
and \U$32089 ( \39893 , \39892 , \38822 );
or \U$32090 ( \39894 , \39883 , \39893 );
and \U$32092 ( \39895 , \39894 , 1'b1 );
or \U$32094 ( \39896 , \39895 , 1'b0 );
buf \U$32095 ( \39897 , \39896 );
_DC r23824_GF_IsGateDCbyConstraint ( \39898_nR23824 , \39897 , \21944 );
buf \U$32096 ( \39899 , \39898_nR23824 );
not \U$32097 ( \39900 , \38705 );
and \U$32098 ( \39901 , RIe069a70_5389, \39900 );
not \U$32099 ( \39902 , RIe069a70_5389);
or \U$32100 ( \39903 , \39902 , \39335 );
not \U$32101 ( \39904 , \39315 );
and \U$32102 ( \39905 , \38693 , \39904 );
not \U$32103 ( \39906 , \39905 );
not \U$32104 ( \39907 , \38690 );
not \U$32105 ( \39908 , \39321 );
or \U$32106 ( \39909 , \39907 , \39908 );
nand \U$32107 ( \39910 , \39903 , \39906 , \39909 );
and \U$32108 ( \39911 , \39910 , \38705 );
or \U$32109 ( \39912 , \39901 , \39911 );
and \U$32111 ( \39913 , \39912 , 1'b1 );
or \U$32113 ( \39914 , \39913 , 1'b0 );
buf \U$32114 ( \39915 , \39914 );
_DC r23826_GF_IsGateDCbyConstraint ( \39916_nR23826 , \39915 , \21944 );
buf \U$32115 ( \39917 , \39916_nR23826 );
not \U$32116 ( \39918 , \38603 );
and \U$32117 ( \39919 , RIe06b870_5390, \39918 );
not \U$32118 ( \39920 , RIe06b870_5390);
or \U$32119 ( \39921 , \39920 , \39356 );
not \U$32120 ( \39922 , \39337 );
and \U$32121 ( \39923 , \38713 , \39922 );
not \U$32122 ( \39924 , \39923 );
not \U$32123 ( \39925 , \38710 );
not \U$32124 ( \39926 , \39342 );
or \U$32125 ( \39927 , \39925 , \39926 );
nand \U$32126 ( \39928 , \39921 , \39924 , \39927 );
and \U$32127 ( \39929 , \39928 , \38603 );
or \U$32128 ( \39930 , \39919 , \39929 );
and \U$32130 ( \39931 , \39930 , 1'b1 );
or \U$32132 ( \39932 , \39931 , 1'b0 );
buf \U$32133 ( \39933 , \39932 );
_DC r23828_GF_IsGateDCbyConstraint ( \39934_nR23828 , \39933 , \21944 );
buf \U$32134 ( \39935 , \39934_nR23828 );
not \U$32135 ( \39936 , \38822 );
and \U$32136 ( \39937 , RIe06cf68_5391, \39936 );
not \U$32137 ( \39938 , RIe06cf68_5391);
or \U$32138 ( \39939 , \39938 , \39313 );
not \U$32139 ( \39940 , \39315 );
and \U$32140 ( \39941 , \38734 , \39940 );
not \U$32141 ( \39942 , \39941 );
not \U$32142 ( \39943 , \38731 );
not \U$32143 ( \39944 , \39321 );
or \U$32144 ( \39945 , \39943 , \39944 );
nand \U$32145 ( \39946 , \39939 , \39942 , \39945 );
and \U$32146 ( \39947 , \39946 , \38822 );
or \U$32147 ( \39948 , \39937 , \39947 );
and \U$32149 ( \39949 , \39948 , 1'b1 );
or \U$32151 ( \39950 , \39949 , 1'b0 );
buf \U$32152 ( \39951 , \39950 );
_DC r2382a_GF_IsGateDCbyConstraint ( \39952_nR2382a , \39951 , \21944 );
buf \U$32153 ( \39953 , \39952_nR2382a );
not \U$32154 ( \39954 , \39163 );
and \U$32155 ( \39955 , RIe06e6d8_5392, \39954 );
not \U$32156 ( \39956 , RIe06e6d8_5392);
or \U$32157 ( \39957 , \39956 , \39356 );
not \U$32158 ( \39958 , \39434 );
and \U$32159 ( \39959 , \38754 , \39958 );
not \U$32160 ( \39960 , \39959 );
not \U$32161 ( \39961 , \38752 );
not \U$32162 ( \39962 , \39321 );
or \U$32163 ( \39963 , \39961 , \39962 );
nand \U$32164 ( \39964 , \39957 , \39960 , \39963 );
and \U$32165 ( \39965 , \39964 , \39163 );
or \U$32166 ( \39966 , \39955 , \39965 );
and \U$32168 ( \39967 , \39966 , 1'b1 );
or \U$32170 ( \39968 , \39967 , 1'b0 );
buf \U$32171 ( \39969 , \39968 );
_DC r2382c_GF_IsGateDCbyConstraint ( \39970_nR2382c , \39969 , \21944 );
buf \U$32172 ( \39971 , \39970_nR2382c );
not \U$32173 ( \39972 , \38603 );
and \U$32174 ( \39973 , RIe06fa10_5393, \39972 );
not \U$32175 ( \39974 , RIe06fa10_5393);
or \U$32176 ( \39975 , \39974 , \39375 );
not \U$32177 ( \39976 , \39315 );
and \U$32178 ( \39977 , \38773 , \39976 );
not \U$32179 ( \39978 , \39977 );
not \U$32180 ( \39979 , \38771 );
not \U$32181 ( \39980 , \39320 );
or \U$32182 ( \39981 , \39979 , \39980 );
nand \U$32183 ( \39982 , \39975 , \39978 , \39981 );
and \U$32184 ( \39983 , \39982 , \38603 );
or \U$32185 ( \39984 , \39973 , \39983 );
and \U$32187 ( \39985 , \39984 , 1'b1 );
or \U$32189 ( \39986 , \39985 , 1'b0 );
buf \U$32190 ( \39987 , \39986 );
_DC r2382e_GF_IsGateDCbyConstraint ( \39988_nR2382e , \39987 , \21944 );
buf \U$32191 ( \39989 , \39988_nR2382e );
not \U$32192 ( \39990 , \39045 );
and \U$32193 ( \39991 , RIe070eb0_5394, \39990 );
not \U$32194 ( \39992 , RIe070eb0_5394);
or \U$32195 ( \39993 , \39992 , \39356 );
not \U$32196 ( \39994 , \39377 );
and \U$32197 ( \39995 , \38792 , \39994 );
not \U$32198 ( \39996 , \39995 );
not \U$32199 ( \39997 , \38789 );
not \U$32200 ( \39998 , \39320 );
or \U$32201 ( \39999 , \39997 , \39998 );
nand \U$32202 ( \40000 , \39993 , \39996 , \39999 );
and \U$32203 ( \40001 , \40000 , \39045 );
or \U$32204 ( \40002 , \39991 , \40001 );
and \U$32206 ( \40003 , \40002 , 1'b1 );
or \U$32208 ( \40004 , \40003 , 1'b0 );
buf \U$32209 ( \40005 , \40004 );
_DC r23830_GF_IsGateDCbyConstraint ( \40006_nR23830 , \40005 , \21944 );
buf \U$32210 ( \40007 , \40006_nR23830 );
buf \U$32211 ( \40008 , \39045 );
not \U$32212 ( \40009 , \40008 );
and \U$32213 ( \40010 , RIe0721e8_5395, \40009 );
not \U$32214 ( \40011 , RIe0721e8_5395);
or \U$32215 ( \40012 , \40011 , \39335 );
not \U$32216 ( \40013 , \39315 );
and \U$32217 ( \40014 , \38810 , \40013 );
not \U$32218 ( \40015 , \40014 );
not \U$32219 ( \40016 , \38808 );
not \U$32220 ( \40017 , \39321 );
or \U$32221 ( \40018 , \40016 , \40017 );
nand \U$32222 ( \40019 , \40012 , \40015 , \40018 );
and \U$32223 ( \40020 , \40019 , \40008 );
or \U$32224 ( \40021 , \40010 , \40020 );
and \U$32226 ( \40022 , \40021 , 1'b1 );
or \U$32228 ( \40023 , \40022 , 1'b0 );
buf \U$32229 ( \40024 , \40023 );
_DC r23832_GF_IsGateDCbyConstraint ( \40025_nR23832 , \40024 , \21944 );
buf \U$32230 ( \40026 , \40025_nR23832 );
not \U$32231 ( \40027 , \40008 );
and \U$32232 ( \40028 , RIe073808_5396, \40027 );
not \U$32233 ( \40029 , RIe073808_5396);
or \U$32234 ( \40030 , \40029 , \39506 );
not \U$32235 ( \40031 , \39434 );
and \U$32236 ( \40032 , \38829 , \40031 );
not \U$32237 ( \40033 , \40032 );
not \U$32238 ( \40034 , \38827 );
not \U$32239 ( \40035 , \39321 );
or \U$32240 ( \40036 , \40034 , \40035 );
nand \U$32241 ( \40037 , \40030 , \40033 , \40036 );
and \U$32242 ( \40038 , \40037 , \40008 );
or \U$32243 ( \40039 , \40028 , \40038 );
and \U$32245 ( \40040 , \40039 , 1'b1 );
or \U$32247 ( \40041 , \40040 , 1'b0 );
buf \U$32248 ( \40042 , \40041 );
_DC r23834_GF_IsGateDCbyConstraint ( \40043_nR23834 , \40042 , \21944 );
buf \U$32249 ( \40044 , \40043_nR23834 );
not \U$32250 ( \40045 , \38033 );
and \U$32251 ( \40046 , RIe074960_5397, \40045 );
not \U$32252 ( \40047 , RIe074960_5397);
or \U$32253 ( \40048 , \40047 , \39506 );
not \U$32254 ( \40049 , \39377 );
and \U$32255 ( \40050 , \38847 , \40049 );
not \U$32256 ( \40051 , \40050 );
not \U$32257 ( \40052 , \38845 );
not \U$32258 ( \40053 , \39342 );
or \U$32259 ( \40054 , \40052 , \40053 );
nand \U$32260 ( \40055 , \40048 , \40051 , \40054 );
and \U$32261 ( \40056 , \40055 , \38033 );
or \U$32262 ( \40057 , \40046 , \40056 );
and \U$32264 ( \40058 , \40057 , 1'b1 );
or \U$32266 ( \40059 , \40058 , 1'b0 );
buf \U$32267 ( \40060 , \40059 );
_DC r23838_GF_IsGateDCbyConstraint ( \40061_nR23838 , \40060 , \21944 );
buf \U$32268 ( \40062 , \40061_nR23838 );
not \U$32269 ( \40063 , \38603 );
and \U$32270 ( \40064 , RIe0762b0_5398, \40063 );
not \U$32271 ( \40065 , RIe0762b0_5398);
or \U$32272 ( \40066 , \40065 , \39313 );
not \U$32273 ( \40067 , \39315 );
and \U$32274 ( \40068 , \38865 , \40067 );
not \U$32275 ( \40069 , \40068 );
not \U$32276 ( \40070 , \38863 );
not \U$32277 ( \40071 , \39400 );
or \U$32278 ( \40072 , \40070 , \40071 );
nand \U$32279 ( \40073 , \40066 , \40069 , \40072 );
and \U$32280 ( \40074 , \40073 , \38603 );
or \U$32281 ( \40075 , \40064 , \40074 );
and \U$32283 ( \40076 , \40075 , 1'b1 );
or \U$32285 ( \40077 , \40076 , 1'b0 );
buf \U$32286 ( \40078 , \40077 );
_DC r2383a_GF_IsGateDCbyConstraint ( \40079_nR2383a , \40078 , \21944 );
buf \U$32287 ( \40080 , \40079_nR2383a );
not \U$32288 ( \40081 , \40008 );
and \U$32289 ( \40082 , RIe0779a8_5399, \40081 );
not \U$32290 ( \40083 , RIe0779a8_5399);
or \U$32291 ( \40084 , \40083 , \39335 );
not \U$32292 ( \40085 , \39337 );
and \U$32293 ( \40086 , \38883 , \40085 );
not \U$32294 ( \40087 , \40086 );
not \U$32295 ( \40088 , \38881 );
not \U$32296 ( \40089 , \39400 );
or \U$32297 ( \40090 , \40088 , \40089 );
nand \U$32298 ( \40091 , \40084 , \40087 , \40090 );
and \U$32299 ( \40092 , \40091 , \40008 );
or \U$32300 ( \40093 , \40082 , \40092 );
and \U$32302 ( \40094 , \40093 , 1'b1 );
or \U$32304 ( \40095 , \40094 , 1'b0 );
buf \U$32305 ( \40096 , \40095 );
_DC r2383c_GF_IsGateDCbyConstraint ( \40097_nR2383c , \40096 , \21944 );
buf \U$32306 ( \40098 , \40097_nR2383c );
not \U$32307 ( \40099 , \39066 );
and \U$32308 ( \40100 , RIe079118_5400, \40099 );
not \U$32309 ( \40101 , RIe079118_5400);
or \U$32310 ( \40102 , \40101 , \39335 );
not \U$32311 ( \40103 , \39337 );
and \U$32312 ( \40104 , \38902 , \40103 );
not \U$32313 ( \40105 , \40104 );
not \U$32314 ( \40106 , \38899 );
not \U$32315 ( \40107 , \39321 );
or \U$32316 ( \40108 , \40106 , \40107 );
nand \U$32317 ( \40109 , \40102 , \40105 , \40108 );
and \U$32318 ( \40110 , \40109 , \39066 );
or \U$32319 ( \40111 , \40100 , \40110 );
and \U$32321 ( \40112 , \40111 , 1'b1 );
or \U$32323 ( \40113 , \40112 , 1'b0 );
buf \U$32324 ( \40114 , \40113 );
_DC r2383e_GF_IsGateDCbyConstraint ( \40115_nR2383e , \40114 , \21944 );
buf \U$32325 ( \40116 , \40115_nR2383e );
not \U$32326 ( \40117 , \40008 );
and \U$32327 ( \40118 , RIe07a798_5401, \40117 );
not \U$32328 ( \40119 , RIe07a798_5401);
or \U$32329 ( \40120 , \40119 , \39375 );
not \U$32330 ( \40121 , \39377 );
and \U$32331 ( \40122 , \38921 , \40121 );
not \U$32332 ( \40123 , \40122 );
not \U$32333 ( \40124 , \38919 );
not \U$32334 ( \40125 , \39400 );
or \U$32335 ( \40126 , \40124 , \40125 );
nand \U$32336 ( \40127 , \40120 , \40123 , \40126 );
and \U$32337 ( \40128 , \40127 , \40008 );
or \U$32338 ( \40129 , \40118 , \40128 );
and \U$32340 ( \40130 , \40129 , 1'b1 );
or \U$32342 ( \40131 , \40130 , 1'b0 );
buf \U$32343 ( \40132 , \40131 );
_DC r23840_GF_IsGateDCbyConstraint ( \40133_nR23840 , \40132 , \21944 );
buf \U$32344 ( \40134 , \40133_nR23840 );
not \U$32345 ( \40135 , \40008 );
and \U$32346 ( \40136 , RIe07bcb0_5402, \40135 );
not \U$32347 ( \40137 , RIe07bcb0_5402);
or \U$32348 ( \40138 , \40137 , \39313 );
not \U$32349 ( \40139 , \39315 );
and \U$32350 ( \40140 , \38940 , \40139 );
not \U$32351 ( \40141 , \40140 );
not \U$32352 ( \40142 , \38937 );
not \U$32353 ( \40143 , \39342 );
or \U$32354 ( \40144 , \40142 , \40143 );
nand \U$32355 ( \40145 , \40138 , \40141 , \40144 );
and \U$32356 ( \40146 , \40145 , \40008 );
or \U$32357 ( \40147 , \40136 , \40146 );
and \U$32359 ( \40148 , \40147 , 1'b1 );
or \U$32361 ( \40149 , \40148 , 1'b0 );
buf \U$32362 ( \40150 , \40149 );
_DC r23842_GF_IsGateDCbyConstraint ( \40151_nR23842 , \40150 , \21944 );
buf \U$32363 ( \40152 , \40151_nR23842 );
not \U$32364 ( \40153 , \38822 );
and \U$32365 ( \40154 , RIe07d768_5403, \40153 );
not \U$32366 ( \40155 , RIe07d768_5403);
or \U$32367 ( \40156 , \40155 , \39506 );
not \U$32368 ( \40157 , \39377 );
and \U$32369 ( \40158 , \38958 , \40157 );
not \U$32370 ( \40159 , \40158 );
not \U$32371 ( \40160 , \38956 );
not \U$32372 ( \40161 , \39400 );
or \U$32373 ( \40162 , \40160 , \40161 );
nand \U$32374 ( \40163 , \40156 , \40159 , \40162 );
and \U$32375 ( \40164 , \40163 , \38822 );
or \U$32376 ( \40165 , \40154 , \40164 );
and \U$32378 ( \40166 , \40165 , 1'b1 );
or \U$32380 ( \40167 , \40166 , 1'b0 );
buf \U$32381 ( \40168 , \40167 );
_DC r23844_GF_IsGateDCbyConstraint ( \40169_nR23844 , \40168 , \21944 );
buf \U$32382 ( \40170 , \40169_nR23844 );
not \U$32383 ( \40171 , \39163 );
and \U$32384 ( \40172 , RIe07f220_5404, \40171 );
not \U$32385 ( \40173 , RIe07f220_5404);
or \U$32386 ( \40174 , \40173 , \39356 );
not \U$32387 ( \40175 , \39315 );
and \U$32388 ( \40176 , \38977 , \40175 );
not \U$32389 ( \40177 , \40176 );
not \U$32390 ( \40178 , \38974 );
not \U$32391 ( \40179 , \39321 );
or \U$32392 ( \40180 , \40178 , \40179 );
nand \U$32393 ( \40181 , \40174 , \40177 , \40180 );
and \U$32394 ( \40182 , \40181 , \39163 );
or \U$32395 ( \40183 , \40172 , \40182 );
and \U$32397 ( \40184 , \40183 , 1'b1 );
or \U$32399 ( \40185 , \40184 , 1'b0 );
buf \U$32400 ( \40186 , \40185 );
_DC r23846_GF_IsGateDCbyConstraint ( \40187_nR23846 , \40186 , \21944 );
buf \U$32401 ( \40188 , \40187_nR23846 );
not \U$32402 ( \40189 , \39045 );
and \U$32403 ( \40190 , RIe080cd8_5405, \40189 );
not \U$32404 ( \40191 , RIe080cd8_5405);
or \U$32405 ( \40192 , \40191 , \39313 );
not \U$32406 ( \40193 , \39337 );
and \U$32407 ( \40194 , \38995 , \40193 );
not \U$32408 ( \40195 , \40194 );
not \U$32409 ( \40196 , \38993 );
not \U$32410 ( \40197 , \39321 );
or \U$32411 ( \40198 , \40196 , \40197 );
nand \U$32412 ( \40199 , \40192 , \40195 , \40198 );
and \U$32413 ( \40200 , \40199 , \39045 );
or \U$32414 ( \40201 , \40190 , \40200 );
and \U$32416 ( \40202 , \40201 , 1'b1 );
or \U$32418 ( \40203 , \40202 , 1'b0 );
buf \U$32419 ( \40204 , \40203 );
_DC r23848_GF_IsGateDCbyConstraint ( \40205_nR23848 , \40204 , \21944 );
buf \U$32420 ( \40206 , \40205_nR23848 );
not \U$32421 ( \40207 , \39163 );
and \U$32422 ( \40208 , RIe082088_5406, \40207 );
not \U$32423 ( \40209 , RIe082088_5406);
or \U$32424 ( \40210 , \40209 , \39335 );
not \U$32425 ( \40211 , \39377 );
and \U$32426 ( \40212 , \39014 , \40211 );
not \U$32427 ( \40213 , \40212 );
not \U$32428 ( \40214 , \39011 );
not \U$32429 ( \40215 , \39342 );
or \U$32430 ( \40216 , \40214 , \40215 );
nand \U$32431 ( \40217 , \40210 , \40213 , \40216 );
and \U$32432 ( \40218 , \40217 , \39163 );
or \U$32433 ( \40219 , \40208 , \40218 );
and \U$32435 ( \40220 , \40219 , 1'b1 );
or \U$32437 ( \40221 , \40220 , 1'b0 );
buf \U$32438 ( \40222 , \40221 );
_DC r2384a_GF_IsGateDCbyConstraint ( \40223_nR2384a , \40222 , \21944 );
buf \U$32439 ( \40224 , \40223_nR2384a );
not \U$32440 ( \40225 , \38603 );
and \U$32441 ( \40226 , RIe083078_5407, \40225 );
not \U$32442 ( \40227 , RIe083078_5407);
or \U$32443 ( \40228 , \40227 , \39356 );
not \U$32444 ( \40229 , \39337 );
and \U$32445 ( \40230 , \39033 , \40229 );
not \U$32446 ( \40231 , \40230 );
not \U$32447 ( \40232 , \39030 );
not \U$32448 ( \40233 , \39400 );
or \U$32449 ( \40234 , \40232 , \40233 );
nand \U$32450 ( \40235 , \40228 , \40231 , \40234 );
and \U$32451 ( \40236 , \40235 , \38603 );
or \U$32452 ( \40237 , \40226 , \40236 );
and \U$32454 ( \40238 , \40237 , 1'b1 );
or \U$32456 ( \40239 , \40238 , 1'b0 );
buf \U$32457 ( \40240 , \40239 );
_DC r2384e_GF_IsGateDCbyConstraint ( \40241_nR2384e , \40240 , \21944 );
buf \U$32458 ( \40242 , \40241_nR2384e );
not \U$32459 ( \40243 , \40008 );
and \U$32460 ( \40244 , RIe0843b0_5408, \40243 );
not \U$32461 ( \40245 , RIe0843b0_5408);
or \U$32462 ( \40246 , \40245 , \39375 );
not \U$32463 ( \40247 , \39377 );
and \U$32464 ( \40248 , \39054 , \40247 );
not \U$32465 ( \40249 , \40248 );
not \U$32466 ( \40250 , \39051 );
not \U$32467 ( \40251 , \39342 );
or \U$32468 ( \40252 , \40250 , \40251 );
nand \U$32469 ( \40253 , \40246 , \40249 , \40252 );
and \U$32470 ( \40254 , \40253 , \40008 );
or \U$32471 ( \40255 , \40244 , \40254 );
and \U$32473 ( \40256 , \40255 , 1'b1 );
or \U$32475 ( \40257 , \40256 , 1'b0 );
buf \U$32476 ( \40258 , \40257 );
_DC r23850_GF_IsGateDCbyConstraint ( \40259_nR23850 , \40258 , \21944 );
buf \U$32477 ( \40260 , \40259_nR23850 );
buf \U$32478 ( \40261 , \38705 );
not \U$32479 ( \40262 , \40261 );
and \U$32480 ( \40263 , RIdfbbbf0_5409, \40262 );
not \U$32481 ( \40264 , RIdfbbbf0_5409);
or \U$32482 ( \40265 , \40264 , \39313 );
not \U$32483 ( \40266 , \39315 );
and \U$32484 ( \40267 , \39074 , \40266 );
not \U$32485 ( \40268 , \40267 );
not \U$32486 ( \40269 , \39071 );
not \U$32487 ( \40270 , \39342 );
or \U$32488 ( \40271 , \40269 , \40270 );
nand \U$32489 ( \40272 , \40265 , \40268 , \40271 );
and \U$32490 ( \40273 , \40272 , \40261 );
or \U$32491 ( \40274 , \40263 , \40273 );
and \U$32493 ( \40275 , \40274 , 1'b1 );
or \U$32495 ( \40276 , \40275 , 1'b0 );
buf \U$32496 ( \40277 , \40276 );
_DC r23852_GF_IsGateDCbyConstraint ( \40278_nR23852 , \40277 , \21944 );
buf \U$32497 ( \40279 , \40278_nR23852 );
not \U$32498 ( \40280 , \38033 );
and \U$32499 ( \40281 , RIdfbd5b8_5410, \40280 );
not \U$32500 ( \40282 , RIdfbd5b8_5410);
or \U$32501 ( \40283 , \40282 , \39313 );
not \U$32502 ( \40284 , \39434 );
and \U$32503 ( \40285 , \39093 , \40284 );
not \U$32504 ( \40286 , \40285 );
not \U$32505 ( \40287 , \39090 );
not \U$32506 ( \40288 , \39400 );
or \U$32507 ( \40289 , \40287 , \40288 );
nand \U$32508 ( \40290 , \40283 , \40286 , \40289 );
and \U$32509 ( \40291 , \40290 , \38033 );
or \U$32510 ( \40292 , \40281 , \40291 );
and \U$32512 ( \40293 , \40292 , 1'b1 );
or \U$32514 ( \40294 , \40293 , 1'b0 );
buf \U$32515 ( \40295 , \40294 );
_DC r23854_GF_IsGateDCbyConstraint ( \40296_nR23854 , \40295 , \21944 );
buf \U$32516 ( \40297 , \40296_nR23854 );
not \U$32517 ( \40298 , \39045 );
and \U$32518 ( \40299 , RIdfbf3b8_5411, \40298 );
not \U$32519 ( \40300 , RIdfbf3b8_5411);
or \U$32520 ( \40301 , \40300 , \39506 );
not \U$32521 ( \40302 , \39377 );
and \U$32522 ( \40303 , \39112 , \40302 );
not \U$32523 ( \40304 , \40303 );
not \U$32524 ( \40305 , \39109 );
not \U$32525 ( \40306 , \39342 );
or \U$32526 ( \40307 , \40305 , \40306 );
nand \U$32527 ( \40308 , \40301 , \40304 , \40307 );
and \U$32528 ( \40309 , \40308 , \39045 );
or \U$32529 ( \40310 , \40299 , \40309 );
and \U$32531 ( \40311 , \40310 , 1'b1 );
or \U$32533 ( \40312 , \40311 , 1'b0 );
buf \U$32534 ( \40313 , \40312 );
_DC r23856_GF_IsGateDCbyConstraint ( \40314_nR23856 , \40313 , \21944 );
buf \U$32535 ( \40315 , \40314_nR23856 );
not \U$32536 ( \40316 , \40261 );
and \U$32537 ( \40317 , RIdfc15f0_5412, \40316 );
not \U$32538 ( \40318 , RIdfc15f0_5412);
or \U$32539 ( \40319 , \40318 , \39506 );
not \U$32540 ( \40320 , \39315 );
and \U$32541 ( \40321 , \39131 , \40320 );
not \U$32542 ( \40322 , \40321 );
not \U$32543 ( \40323 , \39128 );
not \U$32544 ( \40324 , \39400 );
or \U$32545 ( \40325 , \40323 , \40324 );
nand \U$32546 ( \40326 , \40319 , \40322 , \40325 );
and \U$32547 ( \40327 , \40326 , \40261 );
or \U$32548 ( \40328 , \40317 , \40327 );
and \U$32550 ( \40329 , \40328 , 1'b1 );
or \U$32552 ( \40330 , \40329 , 1'b0 );
buf \U$32553 ( \40331 , \40330 );
_DC r23858_GF_IsGateDCbyConstraint ( \40332_nR23858 , \40331 , \21944 );
buf \U$32554 ( \40333 , \40332_nR23858 );
not \U$32555 ( \40334 , \40008 );
and \U$32556 ( \40335 , RIdfc30a8_5413, \40334 );
not \U$32557 ( \40336 , RIdfc30a8_5413);
or \U$32558 ( \40337 , \40336 , \39356 );
not \U$32559 ( \40338 , \39315 );
and \U$32560 ( \40339 , \39151 , \40338 );
not \U$32561 ( \40340 , \40339 );
not \U$32562 ( \40341 , \39148 );
not \U$32563 ( \40342 , \39400 );
or \U$32564 ( \40343 , \40341 , \40342 );
nand \U$32565 ( \40344 , \40337 , \40340 , \40343 );
and \U$32566 ( \40345 , \40344 , \40008 );
or \U$32567 ( \40346 , \40335 , \40345 );
and \U$32569 ( \40347 , \40346 , 1'b1 );
or \U$32571 ( \40348 , \40347 , 1'b0 );
buf \U$32572 ( \40349 , \40348 );
_DC r2385a_GF_IsGateDCbyConstraint ( \40350_nR2385a , \40349 , \21944 );
buf \U$32573 ( \40351 , \40350_nR2385a );
not \U$32574 ( \40352 , \40008 );
and \U$32575 ( \40353 , RIdfc4f20_5414, \40352 );
not \U$32576 ( \40354 , RIdfc4f20_5414);
or \U$32577 ( \40355 , \40354 , \39375 );
not \U$32578 ( \40356 , \39434 );
and \U$32579 ( \40357 , \39171 , \40356 );
not \U$32580 ( \40358 , \40357 );
not \U$32581 ( \40359 , \39169 );
not \U$32582 ( \40360 , \39342 );
or \U$32583 ( \40361 , \40359 , \40360 );
nand \U$32584 ( \40362 , \40355 , \40358 , \40361 );
and \U$32585 ( \40363 , \40362 , \40008 );
or \U$32586 ( \40364 , \40353 , \40363 );
and \U$32588 ( \40365 , \40364 , 1'b1 );
or \U$32590 ( \40366 , \40365 , 1'b0 );
buf \U$32591 ( \40367 , \40366 );
_DC r2385c_GF_IsGateDCbyConstraint ( \40368_nR2385c , \40367 , \21944 );
buf \U$32592 ( \40369 , \40368_nR2385c );
not \U$32593 ( \40370 , \40261 );
and \U$32594 ( \40371 , RIdfc6f00_5415, \40370 );
not \U$32595 ( \40372 , RIdfc6f00_5415);
or \U$32596 ( \40373 , \40372 , \39375 );
not \U$32597 ( \40374 , \39337 );
and \U$32598 ( \40375 , \39190 , \40374 );
not \U$32599 ( \40376 , \40375 );
not \U$32600 ( \40377 , \39188 );
not \U$32601 ( \40378 , \39342 );
or \U$32602 ( \40379 , \40377 , \40378 );
nand \U$32603 ( \40380 , \40373 , \40376 , \40379 );
and \U$32604 ( \40381 , \40380 , \40261 );
or \U$32605 ( \40382 , \40371 , \40381 );
and \U$32607 ( \40383 , \40382 , 1'b1 );
or \U$32609 ( \40384 , \40383 , 1'b0 );
buf \U$32610 ( \40385 , \40384 );
_DC r2385e_GF_IsGateDCbyConstraint ( \40386_nR2385e , \40385 , \21944 );
buf \U$32611 ( \40387 , \40386_nR2385e );
not \U$32612 ( \40388 , \38822 );
and \U$32613 ( \40389 , RIdfc85f8_5416, \40388 );
not \U$32614 ( \40390 , RIdfc85f8_5416);
or \U$32615 ( \40391 , \40390 , \39506 );
not \U$32616 ( \40392 , \39337 );
and \U$32617 ( \40393 , \39211 , \40392 );
not \U$32618 ( \40394 , \40393 );
not \U$32619 ( \40395 , \39208 );
not \U$32620 ( \40396 , \39400 );
or \U$32621 ( \40397 , \40395 , \40396 );
nand \U$32622 ( \40398 , \40391 , \40394 , \40397 );
and \U$32623 ( \40399 , \40398 , \38822 );
or \U$32624 ( \40400 , \40389 , \40399 );
and \U$32626 ( \40401 , \40400 , 1'b1 );
or \U$32628 ( \40402 , \40401 , 1'b0 );
buf \U$32629 ( \40403 , \40402 );
_DC r23860_GF_IsGateDCbyConstraint ( \40404_nR23860 , \40403 , \21944 );
buf \U$32630 ( \40405 , \40404_nR23860 );
not \U$32631 ( \40406 , \38603 );
and \U$32632 ( \40407 , RIdfca3f8_5417, \40406 );
not \U$32633 ( \40408 , RIdfca3f8_5417);
or \U$32634 ( \40409 , \40408 , \39356 );
not \U$32635 ( \40410 , \39337 );
and \U$32636 ( \40411 , \39230 , \40410 );
not \U$32637 ( \40412 , \40411 );
not \U$32638 ( \40413 , \39227 );
not \U$32639 ( \40414 , \39400 );
or \U$32640 ( \40415 , \40413 , \40414 );
nand \U$32641 ( \40416 , \40409 , \40412 , \40415 );
and \U$32642 ( \40417 , \40416 , \38603 );
or \U$32643 ( \40418 , \40407 , \40417 );
and \U$32645 ( \40419 , \40418 , 1'b1 );
or \U$32647 ( \40420 , \40419 , 1'b0 );
buf \U$32648 ( \40421 , \40420 );
_DC r23864_GF_IsGateDCbyConstraint ( \40422_nR23864 , \40421 , \21944 );
buf \U$32649 ( \40423 , \40422_nR23864 );
not \U$32650 ( \40424 , \40261 );
and \U$32651 ( \40425 , RIdfcc720_5418, \40424 );
not \U$32652 ( \40426 , RIdfcc720_5418);
or \U$32653 ( \40427 , \40426 , \39335 );
not \U$32654 ( \40428 , \39337 );
and \U$32655 ( \40429 , \39250 , \40428 );
not \U$32656 ( \40430 , \40429 );
not \U$32657 ( \40431 , \39247 );
not \U$32658 ( \40432 , \39400 );
or \U$32659 ( \40433 , \40431 , \40432 );
nand \U$32660 ( \40434 , \40427 , \40430 , \40433 );
and \U$32661 ( \40435 , \40434 , \40261 );
or \U$32662 ( \40436 , \40425 , \40435 );
and \U$32664 ( \40437 , \40436 , 1'b1 );
or \U$32666 ( \40438 , \40437 , 1'b0 );
buf \U$32667 ( \40439 , \40438 );
_DC r23866_GF_IsGateDCbyConstraint ( \40440_nR23866 , \40439 , \21944 );
buf \U$32668 ( \40441 , \40440_nR23866 );
not \U$32669 ( \40442 , \40008 );
and \U$32670 ( \40443 , RIdfce8e0_5419, \40442 );
not \U$32671 ( \40444 , RIdfce8e0_5419);
or \U$32672 ( \40445 , \40444 , \39506 );
not \U$32673 ( \40446 , \39377 );
and \U$32674 ( \40447 , \39269 , \40446 );
not \U$32675 ( \40448 , \40447 );
not \U$32676 ( \40449 , \39266 );
not \U$32677 ( \40450 , \39342 );
or \U$32678 ( \40451 , \40449 , \40450 );
nand \U$32679 ( \40452 , \40445 , \40448 , \40451 );
and \U$32680 ( \40453 , \40452 , \40008 );
or \U$32681 ( \40454 , \40443 , \40453 );
and \U$32683 ( \40455 , \40454 , 1'b1 );
or \U$32685 ( \40456 , \40455 , 1'b0 );
buf \U$32686 ( \40457 , \40456 );
_DC r23868_GF_IsGateDCbyConstraint ( \40458_nR23868 , \40457 , \21944 );
buf \U$32687 ( \40459 , \40458_nR23868 );
not \U$32688 ( \40460 , \40261 );
and \U$32689 ( \40461 , RIe106478_5420, \40460 );
not \U$32690 ( \40462 , RIe106478_5420);
or \U$32691 ( \40463 , \40462 , \39356 );
not \U$32692 ( \40464 , \39434 );
and \U$32693 ( \40465 , \39288 , \40464 );
not \U$32694 ( \40466 , \40465 );
not \U$32695 ( \40467 , \39285 );
not \U$32696 ( \40468 , \39342 );
or \U$32697 ( \40469 , \40467 , \40468 );
nand \U$32698 ( \40470 , \40463 , \40466 , \40469 );
and \U$32699 ( \40471 , \40470 , \40261 );
or \U$32700 ( \40472 , \40461 , \40471 );
and \U$32702 ( \40473 , \40472 , 1'b1 );
or \U$32704 ( \40474 , \40473 , 1'b0 );
buf \U$32705 ( \40475 , \40474 );
_DC r2386a_GF_IsGateDCbyConstraint ( \40476_nR2386a , \40475 , \21944 );
buf \U$32706 ( \40477 , \40476_nR2386a );
not \U$32707 ( \40478 , \39045 );
and \U$32708 ( \40479 , RIe104948_5421, \40478 );
not \U$32709 ( \40480 , RIe104948_5421);
not \U$32710 ( \40481 , \38046 );
nor \U$32711 ( \40482 , \38047 , \40481 );
and \U$32712 ( \40483 , \40482 , \38031 );
not \U$32713 ( \40484 , \38039 );
or \U$32714 ( \40485 , \38038 , \40484 );
not \U$32715 ( \40486 , \40485 );
nand \U$32716 ( \40487 , \38030 , \40486 );
not \U$32717 ( \40488 , \40487 );
or \U$32718 ( \40489 , \40483 , \40488 );
not \U$32719 ( \40490 , \40489 );
not \U$32720 ( \40491 , \40490 );
or \U$32721 ( \40492 , \40480 , \40491 );
not \U$32722 ( \40493 , \40483 );
not \U$32723 ( \40494 , \40493 );
and \U$32724 ( \40495 , \38058 , \40494 );
not \U$32725 ( \40496 , \40495 );
not \U$32726 ( \40497 , \40487 );
buf \U$32727 ( \40498 , \40497 );
not \U$32728 ( \40499 , \40498 );
or \U$32729 ( \40500 , \39319 , \40499 );
nand \U$32730 ( \40501 , \40492 , \40496 , \40500 );
and \U$32731 ( \40502 , \40501 , \39045 );
or \U$32732 ( \40503 , \40479 , \40502 );
and \U$32734 ( \40504 , \40503 , 1'b1 );
or \U$32736 ( \40505 , \40504 , 1'b0 );
buf \U$32737 ( \40506 , \40505 );
_DC r23874_GF_IsGateDCbyConstraint ( \40507_nR23874 , \40506 , \21944 );
buf \U$32738 ( \40508 , \40507_nR23874 );
not \U$32739 ( \40509 , \40261 );
and \U$32740 ( \40510 , RIe102b48_5422, \40509 );
not \U$32741 ( \40511 , RIe102b48_5422);
not \U$32742 ( \40512 , \40490 );
or \U$32743 ( \40513 , \40511 , \40512 );
not \U$32744 ( \40514 , \40483 );
not \U$32745 ( \40515 , \40514 );
and \U$32746 ( \40516 , \38085 , \40515 );
not \U$32747 ( \40517 , \40516 );
buf \U$32748 ( \40518 , \40497 );
not \U$32749 ( \40519 , \40518 );
or \U$32750 ( \40520 , \39341 , \40519 );
nand \U$32751 ( \40521 , \40513 , \40517 , \40520 );
and \U$32752 ( \40522 , \40521 , \40261 );
or \U$32753 ( \40523 , \40510 , \40522 );
and \U$32755 ( \40524 , \40523 , 1'b1 );
or \U$32757 ( \40525 , \40524 , 1'b0 );
buf \U$32758 ( \40526 , \40525 );
_DC r2388a_GF_IsGateDCbyConstraint ( \40527_nR2388a , \40526 , \21944 );
buf \U$32759 ( \40528 , \40527_nR2388a );
not \U$32760 ( \40529 , \40008 );
and \U$32761 ( \40530 , RIe100f28_5423, \40529 );
not \U$32762 ( \40531 , RIe100f28_5423);
not \U$32763 ( \40532 , \40490 );
or \U$32764 ( \40533 , \40531 , \40532 );
not \U$32765 ( \40534 , \40493 );
and \U$32766 ( \40535 , \38105 , \40534 );
not \U$32767 ( \40536 , \40535 );
not \U$32768 ( \40537 , \40498 );
or \U$32769 ( \40538 , \39361 , \40537 );
nand \U$32770 ( \40539 , \40533 , \40536 , \40538 );
and \U$32771 ( \40540 , \40539 , \40008 );
or \U$32772 ( \40541 , \40530 , \40540 );
and \U$32774 ( \40542 , \40541 , 1'b1 );
or \U$32776 ( \40543 , \40542 , 1'b0 );
buf \U$32777 ( \40544 , \40543 );
_DC r238a0_GF_IsGateDCbyConstraint ( \40545_nR238a0 , \40544 , \21944 );
buf \U$32778 ( \40546 , \40545_nR238a0 );
not \U$32779 ( \40547 , \38822 );
and \U$32780 ( \40548 , RIe0fea20_5424, \40547 );
not \U$32781 ( \40549 , RIe0fea20_5424);
not \U$32782 ( \40550 , \40490 );
or \U$32783 ( \40551 , \40549 , \40550 );
not \U$32784 ( \40552 , \40514 );
and \U$32785 ( \40553 , \38126 , \40552 );
not \U$32786 ( \40554 , \40553 );
not \U$32787 ( \40555 , \40518 );
or \U$32788 ( \40556 , \39381 , \40555 );
nand \U$32789 ( \40557 , \40551 , \40554 , \40556 );
and \U$32790 ( \40558 , \40557 , \38822 );
or \U$32791 ( \40559 , \40548 , \40558 );
and \U$32793 ( \40560 , \40559 , 1'b1 );
or \U$32795 ( \40561 , \40560 , 1'b0 );
buf \U$32796 ( \40562 , \40561 );
_DC r238b6_GF_IsGateDCbyConstraint ( \40563_nR238b6 , \40562 , \21944 );
buf \U$32797 ( \40564 , \40563_nR238b6 );
not \U$32798 ( \40565 , \40261 );
and \U$32799 ( \40566 , RIe0fcd10_5425, \40565 );
not \U$32800 ( \40567 , RIe0fcd10_5425);
or \U$32801 ( \40568 , \40567 , \40550 );
not \U$32802 ( \40569 , \40493 );
and \U$32803 ( \40570 , \38145 , \40569 );
not \U$32804 ( \40571 , \40570 );
buf \U$32805 ( \40572 , \40497 );
not \U$32806 ( \40573 , \40572 );
or \U$32807 ( \40574 , \39399 , \40573 );
nand \U$32808 ( \40575 , \40568 , \40571 , \40574 );
and \U$32809 ( \40576 , \40575 , \40261 );
or \U$32810 ( \40577 , \40566 , \40576 );
and \U$32812 ( \40578 , \40577 , 1'b1 );
or \U$32814 ( \40579 , \40578 , 1'b0 );
buf \U$32815 ( \40580 , \40579 );
_DC r238cc_GF_IsGateDCbyConstraint ( \40581_nR238cc , \40580 , \21944 );
buf \U$32816 ( \40582 , \40581_nR238cc );
not \U$32817 ( \40583 , \40008 );
and \U$32818 ( \40584 , RIe0fa3d0_5426, \40583 );
not \U$32819 ( \40585 , RIe0fa3d0_5426);
or \U$32820 ( \40586 , \40585 , \40550 );
not \U$32821 ( \40587 , \40483 );
not \U$32822 ( \40588 , \40587 );
and \U$32823 ( \40589 , \38166 , \40588 );
not \U$32824 ( \40590 , \40589 );
not \U$32825 ( \40591 , \40518 );
or \U$32826 ( \40592 , \39419 , \40591 );
nand \U$32827 ( \40593 , \40586 , \40590 , \40592 );
and \U$32828 ( \40594 , \40593 , \40008 );
or \U$32829 ( \40595 , \40584 , \40594 );
and \U$32831 ( \40596 , \40595 , 1'b1 );
or \U$32833 ( \40597 , \40596 , 1'b0 );
buf \U$32834 ( \40598 , \40597 );
_DC r238e2_GF_IsGateDCbyConstraint ( \40599_nR238e2 , \40598 , \21944 );
buf \U$32835 ( \40600 , \40599_nR238e2 );
not \U$32836 ( \40601 , \39045 );
and \U$32837 ( \40602 , RIe0f7838_5427, \40601 );
not \U$32838 ( \40603 , RIe0f7838_5427);
or \U$32839 ( \40604 , \40603 , \40512 );
not \U$32840 ( \40605 , \40493 );
and \U$32841 ( \40606 , \38191 , \40605 );
not \U$32842 ( \40607 , \40606 );
not \U$32843 ( \40608 , \40572 );
or \U$32844 ( \40609 , \39438 , \40608 );
nand \U$32845 ( \40610 , \40604 , \40607 , \40609 );
and \U$32846 ( \40611 , \40610 , \39045 );
or \U$32847 ( \40612 , \40602 , \40611 );
and \U$32849 ( \40613 , \40612 , 1'b1 );
or \U$32851 ( \40614 , \40613 , 1'b0 );
buf \U$32852 ( \40615 , \40614 );
_DC r238ec_GF_IsGateDCbyConstraint ( \40616_nR238ec , \40615 , \21944 );
buf \U$32853 ( \40617 , \40616_nR238ec );
not \U$32854 ( \40618 , \40261 );
and \U$32855 ( \40619 , RIe0f5a38_5428, \40618 );
not \U$32856 ( \40620 , RIe0f5a38_5428);
or \U$32857 ( \40621 , \40620 , \40550 );
not \U$32858 ( \40622 , \40514 );
and \U$32859 ( \40623 , \38210 , \40622 );
not \U$32860 ( \40624 , \40623 );
not \U$32861 ( \40625 , \40518 );
or \U$32862 ( \40626 , \39456 , \40625 );
nand \U$32863 ( \40627 , \40621 , \40624 , \40626 );
and \U$32864 ( \40628 , \40627 , \40261 );
or \U$32865 ( \40629 , \40619 , \40628 );
and \U$32867 ( \40630 , \40629 , 1'b1 );
or \U$32869 ( \40631 , \40630 , 1'b0 );
buf \U$32870 ( \40632 , \40631 );
_DC r238ee_GF_IsGateDCbyConstraint ( \40633_nR238ee , \40632 , \21944 );
buf \U$32871 ( \40634 , \40633_nR238ee );
not \U$32872 ( \40635 , \40008 );
and \U$32873 ( \40636 , RIe0f3968_5429, \40635 );
not \U$32874 ( \40637 , RIe0f3968_5429);
or \U$32875 ( \40638 , \40637 , \40491 );
not \U$32876 ( \40639 , \40483 );
not \U$32877 ( \40640 , \40639 );
and \U$32878 ( \40641 , \38230 , \40640 );
not \U$32879 ( \40642 , \40641 );
not \U$32880 ( \40643 , \40572 );
or \U$32881 ( \40644 , \39474 , \40643 );
nand \U$32882 ( \40645 , \40638 , \40642 , \40644 );
and \U$32883 ( \40646 , \40645 , \40008 );
or \U$32884 ( \40647 , \40636 , \40646 );
and \U$32886 ( \40648 , \40647 , 1'b1 );
or \U$32888 ( \40649 , \40648 , 1'b0 );
buf \U$32889 ( \40650 , \40649 );
_DC r238f0_GF_IsGateDCbyConstraint ( \40651_nR238f0 , \40650 , \21944 );
buf \U$32890 ( \40652 , \40651_nR238f0 );
buf \U$32891 ( \40653 , \38603 );
not \U$32892 ( \40654 , \40653 );
and \U$32893 ( \40655 , RIe0f1b68_5430, \40654 );
not \U$32894 ( \40656 , RIe0f1b68_5430);
or \U$32895 ( \40657 , \40656 , \40491 );
not \U$32896 ( \40658 , \40514 );
and \U$32897 ( \40659 , \38250 , \40658 );
not \U$32898 ( \40660 , \40659 );
not \U$32899 ( \40661 , \40572 );
or \U$32900 ( \40662 , \39492 , \40661 );
nand \U$32901 ( \40663 , \40657 , \40660 , \40662 );
and \U$32902 ( \40664 , \40663 , \40653 );
or \U$32903 ( \40665 , \40655 , \40664 );
and \U$32905 ( \40666 , \40665 , 1'b1 );
or \U$32907 ( \40667 , \40666 , 1'b0 );
buf \U$32908 ( \40668 , \40667 );
_DC r238f2_GF_IsGateDCbyConstraint ( \40669_nR238f2 , \40668 , \21944 );
buf \U$32909 ( \40670 , \40669_nR238f2 );
not \U$32910 ( \40671 , \40261 );
and \U$32911 ( \40672 , RIe0f0290_5431, \40671 );
not \U$32912 ( \40673 , RIe0f0290_5431);
not \U$32913 ( \40674 , \40490 );
or \U$32914 ( \40675 , \40673 , \40674 );
not \U$32915 ( \40676 , \40639 );
and \U$32916 ( \40677 , \38271 , \40676 );
not \U$32917 ( \40678 , \40677 );
buf \U$32918 ( \40679 , \40497 );
not \U$32919 ( \40680 , \40679 );
or \U$32920 ( \40681 , \39511 , \40680 );
nand \U$32921 ( \40682 , \40675 , \40678 , \40681 );
and \U$32922 ( \40683 , \40682 , \40261 );
or \U$32923 ( \40684 , \40672 , \40683 );
and \U$32925 ( \40685 , \40684 , 1'b1 );
or \U$32927 ( \40686 , \40685 , 1'b0 );
buf \U$32928 ( \40687 , \40686 );
_DC r23876_GF_IsGateDCbyConstraint ( \40688_nR23876 , \40687 , \21944 );
buf \U$32929 ( \40689 , \40688_nR23876 );
buf \U$32930 ( \40690 , \39045 );
not \U$32931 ( \40691 , \40690 );
and \U$32932 ( \40692 , RIe0ee508_5432, \40691 );
not \U$32933 ( \40693 , RIe0ee508_5432);
or \U$32934 ( \40694 , \40693 , \40512 );
not \U$32935 ( \40695 , \40587 );
and \U$32936 ( \40696 , \38290 , \40695 );
not \U$32937 ( \40697 , \40696 );
not \U$32938 ( \40698 , \40498 );
or \U$32939 ( \40699 , \39529 , \40698 );
nand \U$32940 ( \40700 , \40694 , \40697 , \40699 );
and \U$32941 ( \40701 , \40700 , \40690 );
or \U$32942 ( \40702 , \40692 , \40701 );
and \U$32944 ( \40703 , \40702 , 1'b1 );
or \U$32946 ( \40704 , \40703 , 1'b0 );
buf \U$32947 ( \40705 , \40704 );
_DC r23878_GF_IsGateDCbyConstraint ( \40706_nR23878 , \40705 , \21944 );
buf \U$32948 ( \40707 , \40706_nR23878 );
not \U$32949 ( \40708 , \40653 );
and \U$32950 ( \40709 , RIe0ec690_5433, \40708 );
not \U$32951 ( \40710 , RIe0ec690_5433);
or \U$32952 ( \40711 , \40710 , \40512 );
not \U$32953 ( \40712 , \40483 );
not \U$32954 ( \40713 , \40712 );
and \U$32955 ( \40714 , \38309 , \40713 );
not \U$32956 ( \40715 , \40714 );
not \U$32957 ( \40716 , \40498 );
or \U$32958 ( \40717 , \39547 , \40716 );
nand \U$32959 ( \40718 , \40711 , \40715 , \40717 );
and \U$32960 ( \40719 , \40718 , \40653 );
or \U$32961 ( \40720 , \40709 , \40719 );
and \U$32963 ( \40721 , \40720 , 1'b1 );
or \U$32965 ( \40722 , \40721 , 1'b0 );
buf \U$32966 ( \40723 , \40722 );
_DC r2387a_GF_IsGateDCbyConstraint ( \40724_nR2387a , \40723 , \21944 );
buf \U$32967 ( \40725 , \40724_nR2387a );
not \U$32968 ( \40726 , \40261 );
and \U$32969 ( \40727 , RIe0eaea8_5434, \40726 );
not \U$32970 ( \40728 , RIe0eaea8_5434);
or \U$32971 ( \40729 , \40728 , \40512 );
not \U$32972 ( \40730 , \40493 );
and \U$32973 ( \40731 , \38328 , \40730 );
not \U$32974 ( \40732 , \40731 );
not \U$32975 ( \40733 , \40498 );
or \U$32976 ( \40734 , \39565 , \40733 );
nand \U$32977 ( \40735 , \40729 , \40732 , \40734 );
and \U$32978 ( \40736 , \40735 , \40261 );
or \U$32979 ( \40737 , \40727 , \40736 );
and \U$32981 ( \40738 , \40737 , 1'b1 );
or \U$32983 ( \40739 , \40738 , 1'b0 );
buf \U$32984 ( \40740 , \40739 );
_DC r2387c_GF_IsGateDCbyConstraint ( \40741_nR2387c , \40740 , \21944 );
buf \U$32985 ( \40742 , \40741_nR2387c );
not \U$32986 ( \40743 , \40690 );
and \U$32987 ( \40744 , RIe0e8658_5435, \40743 );
not \U$32988 ( \40745 , RIe0e8658_5435);
or \U$32989 ( \40746 , \40745 , \40491 );
not \U$32990 ( \40747 , \40639 );
and \U$32991 ( \40748 , \38349 , \40747 );
not \U$32992 ( \40749 , \40748 );
not \U$32993 ( \40750 , \40498 );
or \U$32994 ( \40751 , \39583 , \40750 );
nand \U$32995 ( \40752 , \40746 , \40749 , \40751 );
and \U$32996 ( \40753 , \40752 , \40690 );
or \U$32997 ( \40754 , \40744 , \40753 );
and \U$32999 ( \40755 , \40754 , 1'b1 );
or \U$33001 ( \40756 , \40755 , 1'b0 );
buf \U$33002 ( \40757 , \40756 );
_DC r2387e_GF_IsGateDCbyConstraint ( \40758_nR2387e , \40757 , \21944 );
buf \U$33003 ( \40759 , \40758_nR2387e );
not \U$33004 ( \40760 , \40653 );
and \U$33005 ( \40761 , RIe0e54a8_5436, \40760 );
not \U$33006 ( \40762 , RIe0e54a8_5436);
or \U$33007 ( \40763 , \40762 , \40491 );
not \U$33008 ( \40764 , \40587 );
and \U$33009 ( \40765 , \38368 , \40764 );
not \U$33010 ( \40766 , \40765 );
not \U$33011 ( \40767 , \40679 );
or \U$33012 ( \40768 , \39601 , \40767 );
nand \U$33013 ( \40769 , \40763 , \40766 , \40768 );
and \U$33014 ( \40770 , \40769 , \40653 );
or \U$33015 ( \40771 , \40761 , \40770 );
and \U$33017 ( \40772 , \40771 , 1'b1 );
or \U$33019 ( \40773 , \40772 , 1'b0 );
buf \U$33020 ( \40774 , \40773 );
_DC r23880_GF_IsGateDCbyConstraint ( \40775_nR23880 , \40774 , \21944 );
buf \U$33021 ( \40776 , \40775_nR23880 );
not \U$33022 ( \40777 , \40261 );
and \U$33023 ( \40778 , RIe0e2988_5437, \40777 );
not \U$33024 ( \40779 , RIe0e2988_5437);
or \U$33025 ( \40780 , \40779 , \40674 );
not \U$33026 ( \40781 , \40712 );
and \U$33027 ( \40782 , \38387 , \40781 );
not \U$33028 ( \40783 , \40782 );
not \U$33029 ( \40784 , \40572 );
or \U$33030 ( \40785 , \39619 , \40784 );
nand \U$33031 ( \40786 , \40780 , \40783 , \40785 );
and \U$33032 ( \40787 , \40786 , \40261 );
or \U$33033 ( \40788 , \40778 , \40787 );
and \U$33035 ( \40789 , \40788 , 1'b1 );
or \U$33037 ( \40790 , \40789 , 1'b0 );
buf \U$33038 ( \40791 , \40790 );
_DC r23882_GF_IsGateDCbyConstraint ( \40792_nR23882 , \40791 , \21944 );
buf \U$33039 ( \40793 , \40792_nR23882 );
not \U$33040 ( \40794 , \40690 );
and \U$33041 ( \40795 , RIe0e0228_5438, \40794 );
not \U$33042 ( \40796 , RIe0e0228_5438);
or \U$33043 ( \40797 , \40796 , \40512 );
not \U$33044 ( \40798 , \40712 );
and \U$33045 ( \40799 , \38406 , \40798 );
not \U$33046 ( \40800 , \40799 );
not \U$33047 ( \40801 , \40679 );
or \U$33048 ( \40802 , \39637 , \40801 );
nand \U$33049 ( \40803 , \40797 , \40800 , \40802 );
and \U$33050 ( \40804 , \40803 , \40690 );
or \U$33051 ( \40805 , \40795 , \40804 );
and \U$33053 ( \40806 , \40805 , 1'b1 );
or \U$33055 ( \40807 , \40806 , 1'b0 );
buf \U$33056 ( \40808 , \40807 );
_DC r23884_GF_IsGateDCbyConstraint ( \40809_nR23884 , \40808 , \21944 );
buf \U$33057 ( \40810 , \40809_nR23884 );
not \U$33058 ( \40811 , \40653 );
and \U$33059 ( \40812 , RIe0dd7f8_5439, \40811 );
not \U$33060 ( \40813 , RIe0dd7f8_5439);
or \U$33061 ( \40814 , \40813 , \40532 );
not \U$33062 ( \40815 , \40514 );
and \U$33063 ( \40816 , \38425 , \40815 );
not \U$33064 ( \40817 , \40816 );
not \U$33065 ( \40818 , \40572 );
or \U$33066 ( \40819 , \39655 , \40818 );
nand \U$33067 ( \40820 , \40814 , \40817 , \40819 );
and \U$33068 ( \40821 , \40820 , \40653 );
or \U$33069 ( \40822 , \40812 , \40821 );
and \U$33071 ( \40823 , \40822 , 1'b1 );
or \U$33073 ( \40824 , \40823 , 1'b0 );
buf \U$33074 ( \40825 , \40824 );
_DC r23886_GF_IsGateDCbyConstraint ( \40826_nR23886 , \40825 , \21944 );
buf \U$33075 ( \40827 , \40826_nR23886 );
not \U$33076 ( \40828 , \40261 );
and \U$33077 ( \40829 , RIe0da828_5440, \40828 );
not \U$33078 ( \40830 , RIe0da828_5440);
or \U$33079 ( \40831 , \40830 , \40550 );
not \U$33080 ( \40832 , \40514 );
and \U$33081 ( \40833 , \38443 , \40832 );
not \U$33082 ( \40834 , \40833 );
not \U$33083 ( \40835 , \40498 );
or \U$33084 ( \40836 , \39673 , \40835 );
nand \U$33085 ( \40837 , \40831 , \40834 , \40836 );
and \U$33086 ( \40838 , \40837 , \40261 );
or \U$33087 ( \40839 , \40829 , \40838 );
and \U$33089 ( \40840 , \40839 , 1'b1 );
or \U$33091 ( \40841 , \40840 , 1'b0 );
buf \U$33092 ( \40842 , \40841 );
_DC r23888_GF_IsGateDCbyConstraint ( \40843_nR23888 , \40842 , \21944 );
buf \U$33093 ( \40844 , \40843_nR23888 );
not \U$33094 ( \40845 , \40690 );
and \U$33095 ( \40846 , RIe0d7f60_5441, \40845 );
not \U$33096 ( \40847 , RIe0d7f60_5441);
or \U$33097 ( \40848 , \40847 , \40491 );
not \U$33098 ( \40849 , \40493 );
and \U$33099 ( \40850 , \38462 , \40849 );
not \U$33100 ( \40851 , \40850 );
not \U$33101 ( \40852 , \40679 );
or \U$33102 ( \40853 , \39691 , \40852 );
nand \U$33103 ( \40854 , \40848 , \40851 , \40853 );
and \U$33104 ( \40855 , \40854 , \40690 );
or \U$33105 ( \40856 , \40846 , \40855 );
and \U$33107 ( \40857 , \40856 , 1'b1 );
or \U$33109 ( \40858 , \40857 , 1'b0 );
buf \U$33110 ( \40859 , \40858 );
_DC r2388c_GF_IsGateDCbyConstraint ( \40860_nR2388c , \40859 , \21944 );
buf \U$33111 ( \40861 , \40860_nR2388c );
not \U$33112 ( \40862 , \40653 );
and \U$33113 ( \40863 , RIe0d4f18_5442, \40862 );
not \U$33114 ( \40864 , RIe0d4f18_5442);
or \U$33115 ( \40865 , \40864 , \40532 );
not \U$33116 ( \40866 , \40514 );
and \U$33117 ( \40867 , \38481 , \40866 );
not \U$33118 ( \40868 , \40867 );
not \U$33119 ( \40869 , \40518 );
or \U$33120 ( \40870 , \39709 , \40869 );
nand \U$33121 ( \40871 , \40865 , \40868 , \40870 );
and \U$33122 ( \40872 , \40871 , \40653 );
or \U$33123 ( \40873 , \40863 , \40872 );
and \U$33125 ( \40874 , \40873 , 1'b1 );
or \U$33127 ( \40875 , \40874 , 1'b0 );
buf \U$33128 ( \40876 , \40875 );
_DC r2388e_GF_IsGateDCbyConstraint ( \40877_nR2388e , \40876 , \21944 );
buf \U$33129 ( \40878 , \40877_nR2388e );
buf \U$33130 ( \40879 , \38705 );
not \U$33131 ( \40880 , \40879 );
and \U$33132 ( \40881 , RIe0d3280_5443, \40880 );
not \U$33133 ( \40882 , RIe0d3280_5443);
or \U$33134 ( \40883 , \40882 , \40674 );
not \U$33135 ( \40884 , \40514 );
and \U$33136 ( \40885 , \38500 , \40884 );
not \U$33137 ( \40886 , \40885 );
not \U$33138 ( \40887 , \40498 );
or \U$33139 ( \40888 , \39727 , \40887 );
nand \U$33140 ( \40889 , \40883 , \40886 , \40888 );
and \U$33141 ( \40890 , \40889 , \40879 );
or \U$33142 ( \40891 , \40881 , \40890 );
and \U$33144 ( \40892 , \40891 , 1'b1 );
or \U$33146 ( \40893 , \40892 , 1'b0 );
buf \U$33147 ( \40894 , \40893 );
_DC r23890_GF_IsGateDCbyConstraint ( \40895_nR23890 , \40894 , \21944 );
buf \U$33148 ( \40896 , \40895_nR23890 );
not \U$33149 ( \40897 , \40690 );
and \U$33150 ( \40898 , RIe0d02b0_5444, \40897 );
not \U$33151 ( \40899 , RIe0d02b0_5444);
or \U$33152 ( \40900 , \40899 , \40674 );
not \U$33153 ( \40901 , \40639 );
and \U$33154 ( \40902 , \38518 , \40901 );
not \U$33155 ( \40903 , \40902 );
not \U$33156 ( \40904 , \40518 );
or \U$33157 ( \40905 , \39745 , \40904 );
nand \U$33158 ( \40906 , \40900 , \40903 , \40905 );
and \U$33159 ( \40907 , \40906 , \40690 );
or \U$33160 ( \40908 , \40898 , \40907 );
and \U$33162 ( \40909 , \40908 , 1'b1 );
or \U$33164 ( \40910 , \40909 , 1'b0 );
buf \U$33165 ( \40911 , \40910 );
_DC r23892_GF_IsGateDCbyConstraint ( \40912_nR23892 , \40911 , \21944 );
buf \U$33166 ( \40913 , \40912_nR23892 );
not \U$33167 ( \40914 , \40653 );
and \U$33168 ( \40915 , RIe0cdad8_5445, \40914 );
not \U$33169 ( \40916 , RIe0cdad8_5445);
or \U$33170 ( \40917 , \40916 , \40550 );
not \U$33171 ( \40918 , \40639 );
and \U$33172 ( \40919 , \38537 , \40918 );
not \U$33173 ( \40920 , \40919 );
not \U$33174 ( \40921 , \40679 );
or \U$33175 ( \40922 , \39763 , \40921 );
nand \U$33176 ( \40923 , \40917 , \40920 , \40922 );
and \U$33177 ( \40924 , \40923 , \40653 );
or \U$33178 ( \40925 , \40915 , \40924 );
and \U$33180 ( \40926 , \40925 , 1'b1 );
or \U$33182 ( \40927 , \40926 , 1'b0 );
buf \U$33183 ( \40928 , \40927 );
_DC r23894_GF_IsGateDCbyConstraint ( \40929_nR23894 , \40928 , \21944 );
buf \U$33184 ( \40930 , \40929_nR23894 );
not \U$33185 ( \40931 , \40879 );
and \U$33186 ( \40932 , RIe0cae50_5446, \40931 );
not \U$33187 ( \40933 , RIe0cae50_5446);
or \U$33188 ( \40934 , \40933 , \40674 );
not \U$33189 ( \40935 , \40712 );
and \U$33190 ( \40936 , \38555 , \40935 );
not \U$33191 ( \40937 , \40936 );
not \U$33192 ( \40938 , \40518 );
or \U$33193 ( \40939 , \39781 , \40938 );
nand \U$33194 ( \40940 , \40934 , \40937 , \40939 );
and \U$33195 ( \40941 , \40940 , \40879 );
or \U$33196 ( \40942 , \40932 , \40941 );
and \U$33198 ( \40943 , \40942 , 1'b1 );
or \U$33200 ( \40944 , \40943 , 1'b0 );
buf \U$33201 ( \40945 , \40944 );
_DC r23896_GF_IsGateDCbyConstraint ( \40946_nR23896 , \40945 , \21944 );
buf \U$33202 ( \40947 , \40946_nR23896 );
not \U$33203 ( \40948 , \40690 );
and \U$33204 ( \40949 , RIe0c8150_5447, \40948 );
not \U$33205 ( \40950 , RIe0c8150_5447);
or \U$33206 ( \40951 , \40950 , \40532 );
not \U$33207 ( \40952 , \40712 );
and \U$33208 ( \40953 , \38573 , \40952 );
not \U$33209 ( \40954 , \40953 );
not \U$33210 ( \40955 , \40679 );
or \U$33211 ( \40956 , \39799 , \40955 );
nand \U$33212 ( \40957 , \40951 , \40954 , \40956 );
and \U$33213 ( \40958 , \40957 , \40690 );
or \U$33214 ( \40959 , \40949 , \40958 );
and \U$33216 ( \40960 , \40959 , 1'b1 );
or \U$33218 ( \40961 , \40960 , 1'b0 );
buf \U$33219 ( \40962 , \40961 );
_DC r23898_GF_IsGateDCbyConstraint ( \40963_nR23898 , \40962 , \21944 );
buf \U$33220 ( \40964 , \40963_nR23898 );
not \U$33221 ( \40965 , \40653 );
and \U$33222 ( \40966 , RIe0c5d38_5448, \40965 );
not \U$33223 ( \40967 , RIe0c5d38_5448);
or \U$33224 ( \40968 , \40967 , \40550 );
not \U$33225 ( \40969 , \40493 );
and \U$33226 ( \40970 , \38591 , \40969 );
not \U$33227 ( \40971 , \40970 );
not \U$33228 ( \40972 , \40679 );
or \U$33229 ( \40973 , \39817 , \40972 );
nand \U$33230 ( \40974 , \40968 , \40971 , \40973 );
and \U$33231 ( \40975 , \40974 , \40653 );
or \U$33232 ( \40976 , \40966 , \40975 );
and \U$33234 ( \40977 , \40976 , 1'b1 );
or \U$33236 ( \40978 , \40977 , 1'b0 );
buf \U$33237 ( \40979 , \40978 );
_DC r2389a_GF_IsGateDCbyConstraint ( \40980_nR2389a , \40979 , \21944 );
buf \U$33238 ( \40981 , \40980_nR2389a );
not \U$33239 ( \40982 , \40879 );
and \U$33240 ( \40983 , RIe0c3290_5449, \40982 );
not \U$33241 ( \40984 , RIe0c3290_5449);
or \U$33242 ( \40985 , \40984 , \40532 );
not \U$33243 ( \40986 , \40639 );
and \U$33244 ( \40987 , \38612 , \40986 );
not \U$33245 ( \40988 , \40987 );
not \U$33246 ( \40989 , \40498 );
or \U$33247 ( \40990 , \39835 , \40989 );
nand \U$33248 ( \40991 , \40985 , \40988 , \40990 );
and \U$33249 ( \40992 , \40991 , \40879 );
or \U$33250 ( \40993 , \40983 , \40992 );
and \U$33252 ( \40994 , \40993 , 1'b1 );
or \U$33254 ( \40995 , \40994 , 1'b0 );
buf \U$33255 ( \40996 , \40995 );
_DC r2389c_GF_IsGateDCbyConstraint ( \40997_nR2389c , \40996 , \21944 );
buf \U$33256 ( \40998 , \40997_nR2389c );
not \U$33257 ( \40999 , \40690 );
and \U$33258 ( \41000 , RIe0c0d88_5450, \40999 );
not \U$33259 ( \41001 , RIe0c0d88_5450);
or \U$33260 ( \41002 , \41001 , \40550 );
not \U$33261 ( \41003 , \40514 );
and \U$33262 ( \41004 , \38633 , \41003 );
not \U$33263 ( \41005 , \41004 );
not \U$33264 ( \41006 , \40498 );
or \U$33265 ( \41007 , \39853 , \41006 );
nand \U$33266 ( \41008 , \41002 , \41005 , \41007 );
and \U$33267 ( \41009 , \41008 , \40690 );
or \U$33268 ( \41010 , \41000 , \41009 );
and \U$33270 ( \41011 , \41010 , 1'b1 );
or \U$33272 ( \41012 , \41011 , 1'b0 );
buf \U$33273 ( \41013 , \41012 );
_DC r2389e_GF_IsGateDCbyConstraint ( \41014_nR2389e , \41013 , \21944 );
buf \U$33274 ( \41015 , \41014_nR2389e );
not \U$33275 ( \41016 , \40653 );
and \U$33276 ( \41017 , RIe0be628_5451, \41016 );
not \U$33277 ( \41018 , RIe0be628_5451);
or \U$33278 ( \41019 , \41018 , \40674 );
not \U$33279 ( \41020 , \40639 );
and \U$33280 ( \41021 , \38653 , \41020 );
not \U$33281 ( \41022 , \41021 );
not \U$33282 ( \41023 , \40679 );
or \U$33283 ( \41024 , \39871 , \41023 );
nand \U$33284 ( \41025 , \41019 , \41022 , \41024 );
and \U$33285 ( \41026 , \41025 , \40653 );
or \U$33286 ( \41027 , \41017 , \41026 );
and \U$33288 ( \41028 , \41027 , 1'b1 );
or \U$33290 ( \41029 , \41028 , 1'b0 );
buf \U$33291 ( \41030 , \41029 );
_DC r238a2_GF_IsGateDCbyConstraint ( \41031_nR238a2 , \41030 , \21944 );
buf \U$33292 ( \41032 , \41031_nR238a2 );
not \U$33293 ( \41033 , \40879 );
and \U$33294 ( \41034 , RIe0bbdd8_5452, \41033 );
not \U$33295 ( \41035 , RIe0bbdd8_5452);
or \U$33296 ( \41036 , \41035 , \40512 );
not \U$33297 ( \41037 , \40493 );
and \U$33298 ( \41038 , \38673 , \41037 );
not \U$33299 ( \41039 , \41038 );
not \U$33300 ( \41040 , \40679 );
or \U$33301 ( \41041 , \39889 , \41040 );
nand \U$33302 ( \41042 , \41036 , \41039 , \41041 );
and \U$33303 ( \41043 , \41042 , \40879 );
or \U$33304 ( \41044 , \41034 , \41043 );
and \U$33306 ( \41045 , \41044 , 1'b1 );
or \U$33308 ( \41046 , \41045 , 1'b0 );
buf \U$33309 ( \41047 , \41046 );
_DC r238a4_GF_IsGateDCbyConstraint ( \41048_nR238a4 , \41047 , \21944 );
buf \U$33310 ( \41049 , \41048_nR238a4 );
not \U$33311 ( \41050 , \40690 );
and \U$33312 ( \41051 , RIe0b91c8_5453, \41050 );
not \U$33313 ( \41052 , RIe0b91c8_5453);
or \U$33314 ( \41053 , \41052 , \40512 );
not \U$33315 ( \41054 , \40639 );
and \U$33316 ( \41055 , \38693 , \41054 );
not \U$33317 ( \41056 , \41055 );
not \U$33318 ( \41057 , \40498 );
or \U$33319 ( \41058 , \39907 , \41057 );
nand \U$33320 ( \41059 , \41053 , \41056 , \41058 );
and \U$33321 ( \41060 , \41059 , \40690 );
or \U$33322 ( \41061 , \41051 , \41060 );
and \U$33324 ( \41062 , \41061 , 1'b1 );
or \U$33326 ( \41063 , \41062 , 1'b0 );
buf \U$33327 ( \41064 , \41063 );
_DC r238a6_GF_IsGateDCbyConstraint ( \41065_nR238a6 , \41064 , \21944 );
buf \U$33328 ( \41066 , \41065_nR238a6 );
not \U$33329 ( \41067 , \40653 );
and \U$33330 ( \41068 , RIe0b5f28_5454, \41067 );
not \U$33331 ( \41069 , RIe0b5f28_5454);
or \U$33332 ( \41070 , \41069 , \40532 );
not \U$33333 ( \41071 , \40587 );
and \U$33334 ( \41072 , \38713 , \41071 );
not \U$33335 ( \41073 , \41072 );
not \U$33336 ( \41074 , \40679 );
or \U$33337 ( \41075 , \39925 , \41074 );
nand \U$33338 ( \41076 , \41070 , \41073 , \41075 );
and \U$33339 ( \41077 , \41076 , \40653 );
or \U$33340 ( \41078 , \41068 , \41077 );
and \U$33342 ( \41079 , \41078 , 1'b1 );
or \U$33344 ( \41080 , \41079 , 1'b0 );
buf \U$33345 ( \41081 , \41080 );
_DC r238a8_GF_IsGateDCbyConstraint ( \41082_nR238a8 , \41081 , \21944 );
buf \U$33346 ( \41083 , \41082_nR238a8 );
not \U$33347 ( \41084 , \40879 );
and \U$33348 ( \41085 , RIe0b3318_5455, \41084 );
not \U$33349 ( \41086 , RIe0b3318_5455);
or \U$33350 ( \41087 , \41086 , \40491 );
not \U$33351 ( \41088 , \40712 );
and \U$33352 ( \41089 , \38734 , \41088 );
not \U$33353 ( \41090 , \41089 );
not \U$33354 ( \41091 , \40498 );
or \U$33355 ( \41092 , \39943 , \41091 );
nand \U$33356 ( \41093 , \41087 , \41090 , \41092 );
and \U$33357 ( \41094 , \41093 , \40879 );
or \U$33358 ( \41095 , \41085 , \41094 );
and \U$33360 ( \41096 , \41095 , 1'b1 );
or \U$33362 ( \41097 , \41096 , 1'b0 );
buf \U$33363 ( \41098 , \41097 );
_DC r238aa_GF_IsGateDCbyConstraint ( \41099_nR238aa , \41098 , \21944 );
buf \U$33364 ( \41100 , \41099_nR238aa );
not \U$33365 ( \41101 , \40690 );
and \U$33366 ( \41102 , RIe0b02d0_5456, \41101 );
not \U$33367 ( \41103 , RIe0b02d0_5456);
or \U$33368 ( \41104 , \41103 , \40532 );
not \U$33369 ( \41105 , \40493 );
and \U$33370 ( \41106 , \38754 , \41105 );
not \U$33371 ( \41107 , \41106 );
not \U$33372 ( \41108 , \40679 );
or \U$33373 ( \41109 , \39961 , \41108 );
nand \U$33374 ( \41110 , \41104 , \41107 , \41109 );
and \U$33375 ( \41111 , \41110 , \40690 );
or \U$33376 ( \41112 , \41102 , \41111 );
and \U$33378 ( \41113 , \41112 , 1'b1 );
or \U$33380 ( \41114 , \41113 , 1'b0 );
buf \U$33381 ( \41115 , \41114 );
_DC r238ac_GF_IsGateDCbyConstraint ( \41116_nR238ac , \41115 , \21944 );
buf \U$33382 ( \41117 , \41116_nR238ac );
not \U$33383 ( \41118 , \40653 );
and \U$33384 ( \41119 , RIe0adeb8_5457, \41118 );
not \U$33385 ( \41120 , RIe0adeb8_5457);
or \U$33386 ( \41121 , \41120 , \40550 );
not \U$33387 ( \41122 , \40493 );
and \U$33388 ( \41123 , \38773 , \41122 );
not \U$33389 ( \41124 , \41123 );
not \U$33390 ( \41125 , \40679 );
or \U$33391 ( \41126 , \39979 , \41125 );
nand \U$33392 ( \41127 , \41121 , \41124 , \41126 );
and \U$33393 ( \41128 , \41127 , \40653 );
or \U$33394 ( \41129 , \41119 , \41128 );
and \U$33396 ( \41130 , \41129 , 1'b1 );
or \U$33398 ( \41131 , \41130 , 1'b0 );
buf \U$33399 ( \41132 , \41131 );
_DC r238ae_GF_IsGateDCbyConstraint ( \41133_nR238ae , \41132 , \21944 );
buf \U$33400 ( \41134 , \41133_nR238ae );
not \U$33401 ( \41135 , \40879 );
and \U$33402 ( \41136 , RIe0ac0b8_5458, \41135 );
not \U$33403 ( \41137 , RIe0ac0b8_5458);
or \U$33404 ( \41138 , \41137 , \40532 );
not \U$33405 ( \41139 , \40587 );
and \U$33406 ( \41140 , \38792 , \41139 );
not \U$33407 ( \41141 , \41140 );
not \U$33408 ( \41142 , \40679 );
or \U$33409 ( \41143 , \39997 , \41142 );
nand \U$33410 ( \41144 , \41138 , \41141 , \41143 );
and \U$33411 ( \41145 , \41144 , \40879 );
or \U$33412 ( \41146 , \41136 , \41145 );
and \U$33414 ( \41147 , \41146 , 1'b1 );
or \U$33416 ( \41148 , \41147 , 1'b0 );
buf \U$33417 ( \41149 , \41148 );
_DC r238b0_GF_IsGateDCbyConstraint ( \41150_nR238b0 , \41149 , \21944 );
buf \U$33418 ( \41151 , \41150_nR238b0 );
not \U$33419 ( \41152 , \40690 );
and \U$33420 ( \41153 , RIe0aa330_5459, \41152 );
not \U$33421 ( \41154 , RIe0aa330_5459);
or \U$33422 ( \41155 , \41154 , \40512 );
not \U$33423 ( \41156 , \40712 );
and \U$33424 ( \41157 , \38810 , \41156 );
not \U$33425 ( \41158 , \41157 );
not \U$33426 ( \41159 , \40679 );
or \U$33427 ( \41160 , \40016 , \41159 );
nand \U$33428 ( \41161 , \41155 , \41158 , \41160 );
and \U$33429 ( \41162 , \41161 , \40690 );
or \U$33430 ( \41163 , \41153 , \41162 );
and \U$33432 ( \41164 , \41163 , 1'b1 );
or \U$33434 ( \41165 , \41164 , 1'b0 );
buf \U$33435 ( \41166 , \41165 );
_DC r238b2_GF_IsGateDCbyConstraint ( \41167_nR238b2 , \41166 , \21944 );
buf \U$33436 ( \41168 , \41167_nR238b2 );
not \U$33437 ( \41169 , \40653 );
and \U$33438 ( \41170 , RIe0a83c8_5460, \41169 );
not \U$33439 ( \41171 , RIe0a83c8_5460);
or \U$33440 ( \41172 , \41171 , \40674 );
not \U$33441 ( \41173 , \40493 );
and \U$33442 ( \41174 , \38829 , \41173 );
not \U$33443 ( \41175 , \41174 );
not \U$33444 ( \41176 , \40498 );
or \U$33445 ( \41177 , \40034 , \41176 );
nand \U$33446 ( \41178 , \41172 , \41175 , \41177 );
and \U$33447 ( \41179 , \41178 , \40653 );
or \U$33448 ( \41180 , \41170 , \41179 );
and \U$33450 ( \41181 , \41180 , 1'b1 );
or \U$33452 ( \41182 , \41181 , 1'b0 );
buf \U$33453 ( \41183 , \41182 );
_DC r238b4_GF_IsGateDCbyConstraint ( \41184_nR238b4 , \41183 , \21944 );
buf \U$33454 ( \41185 , \41184_nR238b4 );
not \U$33455 ( \41186 , \40879 );
and \U$33456 ( \41187 , RIe0a6a00_5461, \41186 );
not \U$33457 ( \41188 , RIe0a6a00_5461);
or \U$33458 ( \41189 , \41188 , \40674 );
not \U$33459 ( \41190 , \40514 );
and \U$33460 ( \41191 , \38847 , \41190 );
not \U$33461 ( \41192 , \41191 );
not \U$33462 ( \41193 , \40518 );
or \U$33463 ( \41194 , \40052 , \41193 );
nand \U$33464 ( \41195 , \41189 , \41192 , \41194 );
and \U$33465 ( \41196 , \41195 , \40879 );
or \U$33466 ( \41197 , \41187 , \41196 );
and \U$33468 ( \41198 , \41197 , 1'b1 );
or \U$33470 ( \41199 , \41198 , 1'b0 );
buf \U$33471 ( \41200 , \41199 );
_DC r238b8_GF_IsGateDCbyConstraint ( \41201_nR238b8 , \41200 , \21944 );
buf \U$33472 ( \41202 , \41201_nR238b8 );
not \U$33473 ( \41203 , \40690 );
and \U$33474 ( \41204 , RIe0a40c0_5462, \41203 );
not \U$33475 ( \41205 , RIe0a40c0_5462);
or \U$33476 ( \41206 , \41205 , \40491 );
not \U$33477 ( \41207 , \40493 );
and \U$33478 ( \41208 , \38865 , \41207 );
not \U$33479 ( \41209 , \41208 );
not \U$33480 ( \41210 , \40572 );
or \U$33481 ( \41211 , \40070 , \41210 );
nand \U$33482 ( \41212 , \41206 , \41209 , \41211 );
and \U$33483 ( \41213 , \41212 , \40690 );
or \U$33484 ( \41214 , \41204 , \41213 );
and \U$33486 ( \41215 , \41214 , 1'b1 );
or \U$33488 ( \41216 , \41215 , 1'b0 );
buf \U$33489 ( \41217 , \41216 );
_DC r238ba_GF_IsGateDCbyConstraint ( \41218_nR238ba , \41217 , \21944 );
buf \U$33490 ( \41219 , \41218_nR238ba );
not \U$33491 ( \41220 , \40653 );
and \U$33492 ( \41221 , RIe0a2158_5463, \41220 );
not \U$33493 ( \41222 , RIe0a2158_5463);
or \U$33494 ( \41223 , \41222 , \40512 );
not \U$33495 ( \41224 , \40493 );
and \U$33496 ( \41225 , \38883 , \41224 );
not \U$33497 ( \41226 , \41225 );
not \U$33498 ( \41227 , \40679 );
or \U$33499 ( \41228 , \40088 , \41227 );
nand \U$33500 ( \41229 , \41223 , \41226 , \41228 );
and \U$33501 ( \41230 , \41229 , \40653 );
or \U$33502 ( \41231 , \41221 , \41230 );
and \U$33504 ( \41232 , \41231 , 1'b1 );
or \U$33506 ( \41233 , \41232 , 1'b0 );
buf \U$33507 ( \41234 , \41233 );
_DC r238bc_GF_IsGateDCbyConstraint ( \41235_nR238bc , \41234 , \21944 );
buf \U$33508 ( \41236 , \41235_nR238bc );
not \U$33509 ( \41237 , \40879 );
and \U$33510 ( \41238 , RIe0a0010_5464, \41237 );
not \U$33511 ( \41239 , RIe0a0010_5464);
or \U$33512 ( \41240 , \41239 , \40512 );
not \U$33513 ( \41241 , \40514 );
and \U$33514 ( \41242 , \38902 , \41241 );
not \U$33515 ( \41243 , \41242 );
not \U$33516 ( \41244 , \40498 );
or \U$33517 ( \41245 , \40106 , \41244 );
nand \U$33518 ( \41246 , \41240 , \41243 , \41245 );
and \U$33519 ( \41247 , \41246 , \40879 );
or \U$33520 ( \41248 , \41238 , \41247 );
and \U$33522 ( \41249 , \41248 , 1'b1 );
or \U$33524 ( \41250 , \41249 , 1'b0 );
buf \U$33525 ( \41251 , \41250 );
_DC r238be_GF_IsGateDCbyConstraint ( \41252_nR238be , \41251 , \21944 );
buf \U$33526 ( \41253 , \41252_nR238be );
not \U$33527 ( \41254 , \40690 );
and \U$33528 ( \41255 , RIe09e378_5465, \41254 );
not \U$33529 ( \41256 , RIe09e378_5465);
or \U$33530 ( \41257 , \41256 , \40550 );
not \U$33531 ( \41258 , \40493 );
and \U$33532 ( \41259 , \38921 , \41258 );
not \U$33533 ( \41260 , \41259 );
not \U$33534 ( \41261 , \40572 );
or \U$33535 ( \41262 , \40124 , \41261 );
nand \U$33536 ( \41263 , \41257 , \41260 , \41262 );
and \U$33537 ( \41264 , \41263 , \40690 );
or \U$33538 ( \41265 , \41255 , \41264 );
and \U$33540 ( \41266 , \41265 , 1'b1 );
or \U$33542 ( \41267 , \41266 , 1'b0 );
buf \U$33543 ( \41268 , \41267 );
_DC r238c0_GF_IsGateDCbyConstraint ( \41269_nR238c0 , \41268 , \21944 );
buf \U$33544 ( \41270 , \41269_nR238c0 );
buf \U$33545 ( \41271 , \38603 );
not \U$33546 ( \41272 , \41271 );
and \U$33547 ( \41273 , RIe09c668_5466, \41272 );
not \U$33548 ( \41274 , RIe09c668_5466);
or \U$33549 ( \41275 , \41274 , \40491 );
not \U$33550 ( \41276 , \40639 );
and \U$33551 ( \41277 , \38940 , \41276 );
not \U$33552 ( \41278 , \41277 );
not \U$33553 ( \41279 , \40679 );
or \U$33554 ( \41280 , \40142 , \41279 );
nand \U$33555 ( \41281 , \41275 , \41278 , \41280 );
and \U$33556 ( \41282 , \41281 , \41271 );
or \U$33557 ( \41283 , \41273 , \41282 );
and \U$33559 ( \41284 , \41283 , 1'b1 );
or \U$33561 ( \41285 , \41284 , 1'b0 );
buf \U$33562 ( \41286 , \41285 );
_DC r238c2_GF_IsGateDCbyConstraint ( \41287_nR238c2 , \41286 , \21944 );
buf \U$33563 ( \41288 , \41287_nR238c2 );
not \U$33564 ( \41289 , \40879 );
and \U$33565 ( \41290 , RIe09a8e0_5467, \41289 );
not \U$33566 ( \41291 , RIe09a8e0_5467);
or \U$33567 ( \41292 , \41291 , \40674 );
not \U$33568 ( \41293 , \40587 );
and \U$33569 ( \41294 , \38958 , \41293 );
not \U$33570 ( \41295 , \41294 );
not \U$33571 ( \41296 , \40572 );
or \U$33572 ( \41297 , \40160 , \41296 );
nand \U$33573 ( \41298 , \41292 , \41295 , \41297 );
and \U$33574 ( \41299 , \41298 , \40879 );
or \U$33575 ( \41300 , \41290 , \41299 );
and \U$33577 ( \41301 , \41300 , 1'b1 );
or \U$33579 ( \41302 , \41301 , 1'b0 );
buf \U$33580 ( \41303 , \41302 );
_DC r238c4_GF_IsGateDCbyConstraint ( \41304_nR238c4 , \41303 , \21944 );
buf \U$33581 ( \41305 , \41304_nR238c4 );
buf \U$33582 ( \41306 , \39163 );
not \U$33583 ( \41307 , \41306 );
and \U$33584 ( \41308 , RIe099080_5468, \41307 );
not \U$33585 ( \41309 , RIe099080_5468);
or \U$33586 ( \41310 , \41309 , \40532 );
not \U$33587 ( \41311 , \40514 );
and \U$33588 ( \41312 , \38977 , \41311 );
not \U$33589 ( \41313 , \41312 );
not \U$33590 ( \41314 , \40498 );
or \U$33591 ( \41315 , \40178 , \41314 );
nand \U$33592 ( \41316 , \41310 , \41313 , \41315 );
and \U$33593 ( \41317 , \41316 , \41306 );
or \U$33594 ( \41318 , \41308 , \41317 );
and \U$33596 ( \41319 , \41318 , 1'b1 );
or \U$33598 ( \41320 , \41319 , 1'b0 );
buf \U$33599 ( \41321 , \41320 );
_DC r238c6_GF_IsGateDCbyConstraint ( \41322_nR238c6 , \41321 , \21944 );
buf \U$33600 ( \41323 , \41322_nR238c6 );
not \U$33601 ( \41324 , \41271 );
and \U$33602 ( \41325 , RIe1d1cf8_5469, \41324 );
not \U$33603 ( \41326 , RIe1d1cf8_5469);
or \U$33604 ( \41327 , \41326 , \40491 );
not \U$33605 ( \41328 , \40514 );
and \U$33606 ( \41329 , \38995 , \41328 );
not \U$33607 ( \41330 , \41329 );
not \U$33608 ( \41331 , \40498 );
or \U$33609 ( \41332 , \40196 , \41331 );
nand \U$33610 ( \41333 , \41327 , \41330 , \41332 );
and \U$33611 ( \41334 , \41333 , \41271 );
or \U$33612 ( \41335 , \41325 , \41334 );
and \U$33614 ( \41336 , \41335 , 1'b1 );
or \U$33616 ( \41337 , \41336 , 1'b0 );
buf \U$33617 ( \41338 , \41337 );
_DC r238c8_GF_IsGateDCbyConstraint ( \41339_nR238c8 , \41338 , \21944 );
buf \U$33618 ( \41340 , \41339_nR238c8 );
not \U$33619 ( \41341 , \40879 );
and \U$33620 ( \41342 , RIe1d24f0_5470, \41341 );
not \U$33621 ( \41343 , RIe1d24f0_5470);
or \U$33622 ( \41344 , \41343 , \40512 );
not \U$33623 ( \41345 , \40712 );
and \U$33624 ( \41346 , \39014 , \41345 );
not \U$33625 ( \41347 , \41346 );
not \U$33626 ( \41348 , \40518 );
or \U$33627 ( \41349 , \40214 , \41348 );
nand \U$33628 ( \41350 , \41344 , \41347 , \41349 );
and \U$33629 ( \41351 , \41350 , \40879 );
or \U$33630 ( \41352 , \41342 , \41351 );
and \U$33632 ( \41353 , \41352 , 1'b1 );
or \U$33634 ( \41354 , \41353 , 1'b0 );
buf \U$33635 ( \41355 , \41354 );
_DC r238ca_GF_IsGateDCbyConstraint ( \41356_nR238ca , \41355 , \21944 );
buf \U$33636 ( \41357 , \41356_nR238ca );
not \U$33637 ( \41358 , \41306 );
and \U$33638 ( \41359 , RIe1d2ce8_5471, \41358 );
not \U$33639 ( \41360 , RIe1d2ce8_5471);
or \U$33640 ( \41361 , \41360 , \40532 );
not \U$33641 ( \41362 , \40639 );
and \U$33642 ( \41363 , \39033 , \41362 );
not \U$33643 ( \41364 , \41363 );
not \U$33644 ( \41365 , \40572 );
or \U$33645 ( \41366 , \40232 , \41365 );
nand \U$33646 ( \41367 , \41361 , \41364 , \41366 );
and \U$33647 ( \41368 , \41367 , \41306 );
or \U$33648 ( \41369 , \41359 , \41368 );
and \U$33650 ( \41370 , \41369 , 1'b1 );
or \U$33652 ( \41371 , \41370 , 1'b0 );
buf \U$33653 ( \41372 , \41371 );
_DC r238ce_GF_IsGateDCbyConstraint ( \41373_nR238ce , \41372 , \21944 );
buf \U$33654 ( \41374 , \41373_nR238ce );
not \U$33655 ( \41375 , \41271 );
and \U$33656 ( \41376 , RIe1d34e0_5472, \41375 );
not \U$33657 ( \41377 , RIe1d34e0_5472);
or \U$33658 ( \41378 , \41377 , \40550 );
not \U$33659 ( \41379 , \40587 );
and \U$33660 ( \41380 , \39054 , \41379 );
not \U$33661 ( \41381 , \41380 );
not \U$33662 ( \41382 , \40518 );
or \U$33663 ( \41383 , \40250 , \41382 );
nand \U$33664 ( \41384 , \41378 , \41381 , \41383 );
and \U$33665 ( \41385 , \41384 , \41271 );
or \U$33666 ( \41386 , \41376 , \41385 );
and \U$33668 ( \41387 , \41386 , 1'b1 );
or \U$33670 ( \41388 , \41387 , 1'b0 );
buf \U$33671 ( \41389 , \41388 );
_DC r238d0_GF_IsGateDCbyConstraint ( \41390_nR238d0 , \41389 , \21944 );
buf \U$33672 ( \41391 , \41390_nR238d0 );
not \U$33673 ( \41392 , \40879 );
and \U$33674 ( \41393 , RIe1d3cd8_5473, \41392 );
not \U$33675 ( \41394 , RIe1d3cd8_5473);
or \U$33676 ( \41395 , \41394 , \40491 );
not \U$33677 ( \41396 , \40712 );
and \U$33678 ( \41397 , \39074 , \41396 );
not \U$33679 ( \41398 , \41397 );
not \U$33680 ( \41399 , \40518 );
or \U$33681 ( \41400 , \40269 , \41399 );
nand \U$33682 ( \41401 , \41395 , \41398 , \41400 );
and \U$33683 ( \41402 , \41401 , \40879 );
or \U$33684 ( \41403 , \41393 , \41402 );
and \U$33686 ( \41404 , \41403 , 1'b1 );
or \U$33688 ( \41405 , \41404 , 1'b0 );
buf \U$33689 ( \41406 , \41405 );
_DC r238d2_GF_IsGateDCbyConstraint ( \41407_nR238d2 , \41406 , \21944 );
buf \U$33690 ( \41408 , \41407_nR238d2 );
not \U$33691 ( \41409 , \41306 );
and \U$33692 ( \41410 , RIe1d44d0_5474, \41409 );
not \U$33693 ( \41411 , RIe1d44d0_5474);
or \U$33694 ( \41412 , \41411 , \40491 );
not \U$33695 ( \41413 , \40712 );
and \U$33696 ( \41414 , \39093 , \41413 );
not \U$33697 ( \41415 , \41414 );
not \U$33698 ( \41416 , \40572 );
or \U$33699 ( \41417 , \40287 , \41416 );
nand \U$33700 ( \41418 , \41412 , \41415 , \41417 );
and \U$33701 ( \41419 , \41418 , \41306 );
or \U$33702 ( \41420 , \41410 , \41419 );
and \U$33704 ( \41421 , \41420 , 1'b1 );
or \U$33706 ( \41422 , \41421 , 1'b0 );
buf \U$33707 ( \41423 , \41422 );
_DC r238d4_GF_IsGateDCbyConstraint ( \41424_nR238d4 , \41423 , \21944 );
buf \U$33708 ( \41425 , \41424_nR238d4 );
not \U$33709 ( \41426 , \41271 );
and \U$33710 ( \41427 , RIe1d4cc8_5475, \41426 );
not \U$33711 ( \41428 , RIe1d4cc8_5475);
or \U$33712 ( \41429 , \41428 , \40674 );
not \U$33713 ( \41430 , \40587 );
and \U$33714 ( \41431 , \39112 , \41430 );
not \U$33715 ( \41432 , \41431 );
not \U$33716 ( \41433 , \40518 );
or \U$33717 ( \41434 , \40305 , \41433 );
nand \U$33718 ( \41435 , \41429 , \41432 , \41434 );
and \U$33719 ( \41436 , \41435 , \41271 );
or \U$33720 ( \41437 , \41427 , \41436 );
and \U$33722 ( \41438 , \41437 , 1'b1 );
or \U$33724 ( \41439 , \41438 , 1'b0 );
buf \U$33725 ( \41440 , \41439 );
_DC r238d6_GF_IsGateDCbyConstraint ( \41441_nR238d6 , \41440 , \21944 );
buf \U$33726 ( \41442 , \41441_nR238d6 );
not \U$33727 ( \41443 , \40879 );
and \U$33728 ( \41444 , RIe1d54c0_5476, \41443 );
not \U$33729 ( \41445 , RIe1d54c0_5476);
or \U$33730 ( \41446 , \41445 , \40674 );
not \U$33731 ( \41447 , \40493 );
and \U$33732 ( \41448 , \39131 , \41447 );
not \U$33733 ( \41449 , \41448 );
not \U$33734 ( \41450 , \40572 );
or \U$33735 ( \41451 , \40323 , \41450 );
nand \U$33736 ( \41452 , \41446 , \41449 , \41451 );
and \U$33737 ( \41453 , \41452 , \40879 );
or \U$33738 ( \41454 , \41444 , \41453 );
and \U$33740 ( \41455 , \41454 , 1'b1 );
or \U$33742 ( \41456 , \41455 , 1'b0 );
buf \U$33743 ( \41457 , \41456 );
_DC r238d8_GF_IsGateDCbyConstraint ( \41458_nR238d8 , \41457 , \21944 );
buf \U$33744 ( \41459 , \41458_nR238d8 );
not \U$33745 ( \41460 , \41306 );
and \U$33746 ( \41461 , RIe1d5cb8_5477, \41460 );
not \U$33747 ( \41462 , RIe1d5cb8_5477);
or \U$33748 ( \41463 , \41462 , \40532 );
not \U$33749 ( \41464 , \40639 );
and \U$33750 ( \41465 , \39151 , \41464 );
not \U$33751 ( \41466 , \41465 );
not \U$33752 ( \41467 , \40572 );
or \U$33753 ( \41468 , \40341 , \41467 );
nand \U$33754 ( \41469 , \41463 , \41466 , \41468 );
and \U$33755 ( \41470 , \41469 , \41306 );
or \U$33756 ( \41471 , \41461 , \41470 );
and \U$33758 ( \41472 , \41471 , 1'b1 );
or \U$33760 ( \41473 , \41472 , 1'b0 );
buf \U$33761 ( \41474 , \41473 );
_DC r238da_GF_IsGateDCbyConstraint ( \41475_nR238da , \41474 , \21944 );
buf \U$33762 ( \41476 , \41475_nR238da );
not \U$33763 ( \41477 , \41271 );
and \U$33764 ( \41478 , RIe1d64b0_5478, \41477 );
not \U$33765 ( \41479 , RIe1d64b0_5478);
or \U$33766 ( \41480 , \41479 , \40550 );
not \U$33767 ( \41481 , \40587 );
and \U$33768 ( \41482 , \39171 , \41481 );
not \U$33769 ( \41483 , \41482 );
not \U$33770 ( \41484 , \40518 );
or \U$33771 ( \41485 , \40359 , \41484 );
nand \U$33772 ( \41486 , \41480 , \41483 , \41485 );
and \U$33773 ( \41487 , \41486 , \41271 );
or \U$33774 ( \41488 , \41478 , \41487 );
and \U$33776 ( \41489 , \41488 , 1'b1 );
or \U$33778 ( \41490 , \41489 , 1'b0 );
buf \U$33779 ( \41491 , \41490 );
_DC r238dc_GF_IsGateDCbyConstraint ( \41492_nR238dc , \41491 , \21944 );
buf \U$33780 ( \41493 , \41492_nR238dc );
buf \U$33781 ( \41494 , \39066 );
not \U$33782 ( \41495 , \41494 );
and \U$33783 ( \41496 , RIe1d6ca8_5479, \41495 );
not \U$33784 ( \41497 , RIe1d6ca8_5479);
or \U$33785 ( \41498 , \41497 , \40550 );
not \U$33786 ( \41499 , \40712 );
and \U$33787 ( \41500 , \39190 , \41499 );
not \U$33788 ( \41501 , \41500 );
not \U$33789 ( \41502 , \40518 );
or \U$33790 ( \41503 , \40377 , \41502 );
nand \U$33791 ( \41504 , \41498 , \41501 , \41503 );
and \U$33792 ( \41505 , \41504 , \41494 );
or \U$33793 ( \41506 , \41496 , \41505 );
and \U$33795 ( \41507 , \41506 , 1'b1 );
or \U$33797 ( \41508 , \41507 , 1'b0 );
buf \U$33798 ( \41509 , \41508 );
_DC r238de_GF_IsGateDCbyConstraint ( \41510_nR238de , \41509 , \21944 );
buf \U$33799 ( \41511 , \41510_nR238de );
not \U$33800 ( \41512 , \41306 );
and \U$33801 ( \41513 , RIe1d74a0_5480, \41512 );
not \U$33802 ( \41514 , RIe1d74a0_5480);
or \U$33803 ( \41515 , \41514 , \40674 );
not \U$33804 ( \41516 , \40514 );
and \U$33805 ( \41517 , \39211 , \41516 );
not \U$33806 ( \41518 , \41517 );
not \U$33807 ( \41519 , \40572 );
or \U$33808 ( \41520 , \40395 , \41519 );
nand \U$33809 ( \41521 , \41515 , \41518 , \41520 );
and \U$33810 ( \41522 , \41521 , \41306 );
or \U$33811 ( \41523 , \41513 , \41522 );
and \U$33813 ( \41524 , \41523 , 1'b1 );
or \U$33815 ( \41525 , \41524 , 1'b0 );
buf \U$33816 ( \41526 , \41525 );
_DC r238e0_GF_IsGateDCbyConstraint ( \41527_nR238e0 , \41526 , \21944 );
buf \U$33817 ( \41528 , \41527_nR238e0 );
not \U$33818 ( \41529 , \41271 );
and \U$33819 ( \41530 , RIe1d7c98_5481, \41529 );
not \U$33820 ( \41531 , RIe1d7c98_5481);
or \U$33821 ( \41532 , \41531 , \40532 );
not \U$33822 ( \41533 , \40587 );
and \U$33823 ( \41534 , \39230 , \41533 );
not \U$33824 ( \41535 , \41534 );
not \U$33825 ( \41536 , \40572 );
or \U$33826 ( \41537 , \40413 , \41536 );
nand \U$33827 ( \41538 , \41532 , \41535 , \41537 );
and \U$33828 ( \41539 , \41538 , \41271 );
or \U$33829 ( \41540 , \41530 , \41539 );
and \U$33831 ( \41541 , \41540 , 1'b1 );
or \U$33833 ( \41542 , \41541 , 1'b0 );
buf \U$33834 ( \41543 , \41542 );
_DC r238e4_GF_IsGateDCbyConstraint ( \41544_nR238e4 , \41543 , \21944 );
buf \U$33835 ( \41545 , \41544_nR238e4 );
not \U$33836 ( \41546 , \41494 );
and \U$33837 ( \41547 , RIe1d8490_5482, \41546 );
not \U$33838 ( \41548 , RIe1d8490_5482);
or \U$33839 ( \41549 , \41548 , \40512 );
not \U$33840 ( \41550 , \40587 );
and \U$33841 ( \41551 , \39250 , \41550 );
not \U$33842 ( \41552 , \41551 );
not \U$33843 ( \41553 , \40572 );
or \U$33844 ( \41554 , \40431 , \41553 );
nand \U$33845 ( \41555 , \41549 , \41552 , \41554 );
and \U$33846 ( \41556 , \41555 , \41494 );
or \U$33847 ( \41557 , \41547 , \41556 );
and \U$33849 ( \41558 , \41557 , 1'b1 );
or \U$33851 ( \41559 , \41558 , 1'b0 );
buf \U$33852 ( \41560 , \41559 );
_DC r238e6_GF_IsGateDCbyConstraint ( \41561_nR238e6 , \41560 , \21944 );
buf \U$33853 ( \41562 , \41561_nR238e6 );
not \U$33854 ( \41563 , \41306 );
and \U$33855 ( \41564 , RIe1d8c88_5483, \41563 );
not \U$33856 ( \41565 , RIe1d8c88_5483);
or \U$33857 ( \41566 , \41565 , \40674 );
not \U$33858 ( \41567 , \40639 );
and \U$33859 ( \41568 , \39269 , \41567 );
not \U$33860 ( \41569 , \41568 );
not \U$33861 ( \41570 , \40518 );
or \U$33862 ( \41571 , \40449 , \41570 );
nand \U$33863 ( \41572 , \41566 , \41569 , \41571 );
and \U$33864 ( \41573 , \41572 , \41306 );
or \U$33865 ( \41574 , \41564 , \41573 );
and \U$33867 ( \41575 , \41574 , 1'b1 );
or \U$33869 ( \41576 , \41575 , 1'b0 );
buf \U$33870 ( \41577 , \41576 );
_DC r238e8_GF_IsGateDCbyConstraint ( \41578_nR238e8 , \41577 , \21944 );
buf \U$33871 ( \41579 , \41578_nR238e8 );
not \U$33872 ( \41580 , \41271 );
and \U$33873 ( \41581 , RIe1d9480_5484, \41580 );
not \U$33874 ( \41582 , RIe1d9480_5484);
or \U$33875 ( \41583 , \41582 , \40532 );
not \U$33876 ( \41584 , \40712 );
and \U$33877 ( \41585 , \39288 , \41584 );
not \U$33878 ( \41586 , \41585 );
not \U$33879 ( \41587 , \40518 );
or \U$33880 ( \41588 , \40467 , \41587 );
nand \U$33881 ( \41589 , \41583 , \41586 , \41588 );
and \U$33882 ( \41590 , \41589 , \41271 );
or \U$33883 ( \41591 , \41581 , \41590 );
and \U$33885 ( \41592 , \41591 , 1'b1 );
or \U$33887 ( \41593 , \41592 , 1'b0 );
buf \U$33888 ( \41594 , \41593 );
_DC r238ea_GF_IsGateDCbyConstraint ( \41595_nR238ea , \41594 , \21944 );
buf \U$33889 ( \41596 , \41595_nR238ea );
not \U$33890 ( \41597 , \41494 );
and \U$33891 ( \41598 , RIe1d9c78_5485, \41597 );
not \U$33892 ( \41599 , RIe1d9c78_5485);
nand \U$33893 ( \41600 , \38047 , \38046 );
not \U$33894 ( \41601 , \38031 );
or \U$33895 ( \41602 , \41600 , \41601 );
nand \U$33896 ( \41603 , \38039 , \38038 );
not \U$33897 ( \41604 , \41603 );
nand \U$33898 ( \41605 , \38030 , \41604 );
nand \U$33899 ( \41606 , \41602 , \41605 );
or \U$33900 ( \41607 , \41599 , \41606 );
not \U$33901 ( \41608 , \41605 );
buf \U$33902 ( \41609 , \41608 );
nand \U$33903 ( \41610 , \38055 , \41609 );
not \U$33904 ( \41611 , \41602 );
buf \U$33905 ( \41612 , \41611 );
nand \U$33906 ( \41613 , \38058 , \41612 );
nand \U$33907 ( \41614 , \41607 , \41610 , \41613 );
and \U$33908 ( \41615 , \41614 , \41494 );
or \U$33909 ( \41616 , \41598 , \41615 );
and \U$33911 ( \41617 , \41616 , 1'b1 );
or \U$33913 ( \41618 , \41617 , 1'b0 );
buf \U$33914 ( \41619 , \41618 );
_DC r238f4_GF_IsGateDCbyConstraint ( \41620_nR238f4 , \41619 , \21944 );
buf \U$33915 ( \41621 , \41620_nR238f4 );
not \U$33916 ( \41622 , \41306 );
and \U$33917 ( \41623 , RIe1da470_5486, \41622 );
not \U$33918 ( \41624 , RIe1da470_5486);
buf \U$33919 ( \41625 , \41606 );
or \U$33920 ( \41626 , \41624 , \41625 );
buf \U$33921 ( \41627 , \41608 );
nand \U$33922 ( \41628 , \38083 , \41627 );
nand \U$33923 ( \41629 , \38085 , \41612 );
nand \U$33924 ( \41630 , \41626 , \41628 , \41629 );
and \U$33925 ( \41631 , \41630 , \41306 );
or \U$33926 ( \41632 , \41623 , \41631 );
and \U$33928 ( \41633 , \41632 , 1'b1 );
or \U$33930 ( \41634 , \41633 , 1'b0 );
buf \U$33931 ( \41635 , \41634 );
_DC r2390a_GF_IsGateDCbyConstraint ( \41636_nR2390a , \41635 , \21944 );
buf \U$33932 ( \41637 , \41636_nR2390a );
not \U$33933 ( \41638 , \41271 );
and \U$33934 ( \41639 , RIe1dac68_5487, \41638 );
not \U$33935 ( \41640 , RIe1dac68_5487);
buf \U$33936 ( \41641 , \41606 );
or \U$33937 ( \41642 , \41640 , \41641 );
buf \U$33938 ( \41643 , \41608 );
nand \U$33939 ( \41644 , \38102 , \41643 );
buf \U$33940 ( \41645 , \41611 );
nand \U$33941 ( \41646 , \38105 , \41645 );
nand \U$33942 ( \41647 , \41642 , \41644 , \41646 );
and \U$33943 ( \41648 , \41647 , \41271 );
or \U$33944 ( \41649 , \41639 , \41648 );
and \U$33946 ( \41650 , \41649 , 1'b1 );
or \U$33948 ( \41651 , \41650 , 1'b0 );
buf \U$33949 ( \41652 , \41651 );
_DC r23920_GF_IsGateDCbyConstraint ( \41653_nR23920 , \41652 , \21944 );
buf \U$33950 ( \41654 , \41653_nR23920 );
not \U$33951 ( \41655 , \41494 );
and \U$33952 ( \41656 , RIe1db460_5488, \41655 );
not \U$33953 ( \41657 , RIe1db460_5488);
buf \U$33954 ( \41658 , \41606 );
or \U$33955 ( \41659 , \41657 , \41658 );
nand \U$33956 ( \41660 , \38123 , \41609 );
buf \U$33957 ( \41661 , \41611 );
nand \U$33958 ( \41662 , \38126 , \41661 );
nand \U$33959 ( \41663 , \41659 , \41660 , \41662 );
and \U$33960 ( \41664 , \41663 , \41494 );
or \U$33961 ( \41665 , \41656 , \41664 );
and \U$33963 ( \41666 , \41665 , 1'b1 );
or \U$33965 ( \41667 , \41666 , 1'b0 );
buf \U$33966 ( \41668 , \41667 );
_DC r23936_GF_IsGateDCbyConstraint ( \41669_nR23936 , \41668 , \21944 );
buf \U$33967 ( \41670 , \41669_nR23936 );
not \U$33968 ( \41671 , \41306 );
and \U$33969 ( \41672 , RIe1dbc58_5489, \41671 );
not \U$33970 ( \41673 , RIe1dbc58_5489);
or \U$33971 ( \41674 , \41673 , \41625 );
nand \U$33972 ( \41675 , \38143 , \41643 );
nand \U$33973 ( \41676 , \38145 , \41645 );
nand \U$33974 ( \41677 , \41674 , \41675 , \41676 );
and \U$33975 ( \41678 , \41677 , \41306 );
or \U$33976 ( \41679 , \41672 , \41678 );
and \U$33978 ( \41680 , \41679 , 1'b1 );
or \U$33980 ( \41681 , \41680 , 1'b0 );
buf \U$33981 ( \41682 , \41681 );
_DC r2394c_GF_IsGateDCbyConstraint ( \41683_nR2394c , \41682 , \21944 );
buf \U$33982 ( \41684 , \41683_nR2394c );
not \U$33983 ( \41685 , \41271 );
and \U$33984 ( \41686 , RIe1dc450_5490, \41685 );
not \U$33985 ( \41687 , RIe1dc450_5490);
or \U$33986 ( \41688 , \41687 , \41625 );
nand \U$33987 ( \41689 , \38163 , \41627 );
buf \U$33988 ( \41690 , \41611 );
nand \U$33989 ( \41691 , \38166 , \41690 );
nand \U$33990 ( \41692 , \41688 , \41689 , \41691 );
and \U$33991 ( \41693 , \41692 , \41271 );
or \U$33992 ( \41694 , \41686 , \41693 );
and \U$33994 ( \41695 , \41694 , 1'b1 );
or \U$33996 ( \41696 , \41695 , 1'b0 );
buf \U$33997 ( \41697 , \41696 );
_DC r23962_GF_IsGateDCbyConstraint ( \41698_nR23962 , \41697 , \21944 );
buf \U$33998 ( \41699 , \41698_nR23962 );
not \U$33999 ( \41700 , \41494 );
and \U$34000 ( \41701 , RIe1dcc48_5491, \41700 );
not \U$34001 ( \41702 , RIe1dcc48_5491);
or \U$34002 ( \41703 , \41702 , \41641 );
nand \U$34003 ( \41704 , \38188 , \41643 );
nand \U$34004 ( \41705 , \38191 , \41612 );
nand \U$34005 ( \41706 , \41703 , \41704 , \41705 );
and \U$34006 ( \41707 , \41706 , \41494 );
or \U$34007 ( \41708 , \41701 , \41707 );
and \U$34009 ( \41709 , \41708 , 1'b1 );
or \U$34011 ( \41710 , \41709 , 1'b0 );
buf \U$34012 ( \41711 , \41710 );
_DC r2396c_GF_IsGateDCbyConstraint ( \41712_nR2396c , \41711 , \21944 );
buf \U$34013 ( \41713 , \41712_nR2396c );
not \U$34014 ( \41714 , \41306 );
and \U$34015 ( \41715 , RIe1dd440_5492, \41714 );
not \U$34016 ( \41716 , RIe1dd440_5492);
or \U$34017 ( \41717 , \41716 , \41625 );
nand \U$34018 ( \41718 , \38207 , \41643 );
nand \U$34019 ( \41719 , \38210 , \41612 );
nand \U$34020 ( \41720 , \41717 , \41718 , \41719 );
and \U$34021 ( \41721 , \41720 , \41306 );
or \U$34022 ( \41722 , \41715 , \41721 );
and \U$34024 ( \41723 , \41722 , 1'b1 );
or \U$34026 ( \41724 , \41723 , 1'b0 );
buf \U$34027 ( \41725 , \41724 );
_DC r2396e_GF_IsGateDCbyConstraint ( \41726_nR2396e , \41725 , \21944 );
buf \U$34028 ( \41727 , \41726_nR2396e );
not \U$34029 ( \41728 , \41271 );
and \U$34030 ( \41729 , RIe1ddc38_5493, \41728 );
not \U$34031 ( \41730 , RIe1ddc38_5493);
or \U$34032 ( \41731 , \41730 , \41625 );
nand \U$34033 ( \41732 , \38228 , \41609 );
nand \U$34034 ( \41733 , \38230 , \41661 );
nand \U$34035 ( \41734 , \41731 , \41732 , \41733 );
and \U$34036 ( \41735 , \41734 , \41271 );
or \U$34037 ( \41736 , \41729 , \41735 );
and \U$34039 ( \41737 , \41736 , 1'b1 );
or \U$34041 ( \41738 , \41737 , 1'b0 );
buf \U$34042 ( \41739 , \41738 );
_DC r23970_GF_IsGateDCbyConstraint ( \41740_nR23970 , \41739 , \21944 );
buf \U$34043 ( \41741 , \41740_nR23970 );
not \U$34044 ( \41742 , \41494 );
and \U$34045 ( \41743 , RIe1de430_5494, \41742 );
not \U$34046 ( \41744 , RIe1de430_5494);
buf \U$34047 ( \41745 , \41606 );
or \U$34048 ( \41746 , \41744 , \41745 );
nand \U$34049 ( \41747 , \38247 , \41643 );
nand \U$34050 ( \41748 , \38250 , \41645 );
nand \U$34051 ( \41749 , \41746 , \41747 , \41748 );
and \U$34052 ( \41750 , \41749 , \41494 );
or \U$34053 ( \41751 , \41743 , \41750 );
and \U$34055 ( \41752 , \41751 , 1'b1 );
or \U$34057 ( \41753 , \41752 , 1'b0 );
buf \U$34058 ( \41754 , \41753 );
_DC r23972_GF_IsGateDCbyConstraint ( \41755_nR23972 , \41754 , \21944 );
buf \U$34059 ( \41756 , \41755_nR23972 );
not \U$34060 ( \41757 , \41306 );
and \U$34061 ( \41758 , RIe1dec28_5495, \41757 );
not \U$34062 ( \41759 , RIe1dec28_5495);
or \U$34063 ( \41760 , \41759 , \41745 );
nand \U$34064 ( \41761 , \38269 , \41609 );
nand \U$34065 ( \41762 , \38271 , \41690 );
nand \U$34066 ( \41763 , \41760 , \41761 , \41762 );
and \U$34067 ( \41764 , \41763 , \41306 );
or \U$34068 ( \41765 , \41758 , \41764 );
and \U$34070 ( \41766 , \41765 , 1'b1 );
or \U$34072 ( \41767 , \41766 , 1'b0 );
buf \U$34073 ( \41768 , \41767 );
_DC r238f6_GF_IsGateDCbyConstraint ( \41769_nR238f6 , \41768 , \21944 );
buf \U$34074 ( \41770 , \41769_nR238f6 );
not \U$34075 ( \41771 , \41271 );
and \U$34076 ( \41772 , RIe1df420_5496, \41771 );
not \U$34077 ( \41773 , RIe1df420_5496);
or \U$34078 ( \41774 , \41773 , \41658 );
nand \U$34079 ( \41775 , \38287 , \41643 );
nand \U$34080 ( \41776 , \38290 , \41645 );
nand \U$34081 ( \41777 , \41774 , \41775 , \41776 );
and \U$34082 ( \41778 , \41777 , \41271 );
or \U$34083 ( \41779 , \41772 , \41778 );
and \U$34085 ( \41780 , \41779 , 1'b1 );
or \U$34087 ( \41781 , \41780 , 1'b0 );
buf \U$34088 ( \41782 , \41781 );
_DC r238f8_GF_IsGateDCbyConstraint ( \41783_nR238f8 , \41782 , \21944 );
buf \U$34089 ( \41784 , \41783_nR238f8 );
not \U$34090 ( \41785 , \41494 );
and \U$34091 ( \41786 , RIe1dfc18_5497, \41785 );
not \U$34092 ( \41787 , RIe1dfc18_5497);
or \U$34093 ( \41788 , \41787 , \41641 );
nand \U$34094 ( \41789 , \38307 , \41627 );
nand \U$34095 ( \41790 , \38309 , \41690 );
nand \U$34096 ( \41791 , \41788 , \41789 , \41790 );
and \U$34097 ( \41792 , \41791 , \41494 );
or \U$34098 ( \41793 , \41786 , \41792 );
and \U$34100 ( \41794 , \41793 , 1'b1 );
or \U$34102 ( \41795 , \41794 , 1'b0 );
buf \U$34103 ( \41796 , \41795 );
_DC r238fa_GF_IsGateDCbyConstraint ( \41797_nR238fa , \41796 , \21944 );
buf \U$34104 ( \41798 , \41797_nR238fa );
not \U$34105 ( \41799 , \41306 );
and \U$34106 ( \41800 , RIe1e0410_5498, \41799 );
not \U$34107 ( \41801 , RIe1e0410_5498);
or \U$34108 ( \41802 , \41801 , \41658 );
nand \U$34109 ( \41803 , \38325 , \41643 );
nand \U$34110 ( \41804 , \38328 , \41661 );
nand \U$34111 ( \41805 , \41802 , \41803 , \41804 );
and \U$34112 ( \41806 , \41805 , \41306 );
or \U$34113 ( \41807 , \41800 , \41806 );
and \U$34115 ( \41808 , \41807 , 1'b1 );
or \U$34117 ( \41809 , \41808 , 1'b0 );
buf \U$34118 ( \41810 , \41809 );
_DC r238fc_GF_IsGateDCbyConstraint ( \41811_nR238fc , \41810 , \21944 );
buf \U$34119 ( \41812 , \41811_nR238fc );
not \U$34120 ( \41813 , \41271 );
and \U$34121 ( \41814 , RIe1e0c08_5499, \41813 );
not \U$34122 ( \41815 , RIe1e0c08_5499);
or \U$34123 ( \41816 , \41815 , \41625 );
buf \U$34124 ( \41817 , \41608 );
nand \U$34125 ( \41818 , \38346 , \41817 );
nand \U$34126 ( \41819 , \38349 , \41645 );
nand \U$34127 ( \41820 , \41816 , \41818 , \41819 );
and \U$34128 ( \41821 , \41820 , \41271 );
or \U$34129 ( \41822 , \41814 , \41821 );
and \U$34131 ( \41823 , \41822 , 1'b1 );
or \U$34133 ( \41824 , \41823 , 1'b0 );
buf \U$34134 ( \41825 , \41824 );
_DC r238fe_GF_IsGateDCbyConstraint ( \41826_nR238fe , \41825 , \21944 );
buf \U$34135 ( \41827 , \41826_nR238fe );
not \U$34136 ( \41828 , \41494 );
and \U$34137 ( \41829 , RIe1e1400_5500, \41828 );
not \U$34138 ( \41830 , RIe1e1400_5500);
or \U$34139 ( \41831 , \41830 , \41625 );
nand \U$34140 ( \41832 , \38365 , \41627 );
nand \U$34141 ( \41833 , \38368 , \41690 );
nand \U$34142 ( \41834 , \41831 , \41832 , \41833 );
and \U$34143 ( \41835 , \41834 , \41494 );
or \U$34144 ( \41836 , \41829 , \41835 );
and \U$34146 ( \41837 , \41836 , 1'b1 );
or \U$34148 ( \41838 , \41837 , 1'b0 );
buf \U$34149 ( \41839 , \41838 );
_DC r23900_GF_IsGateDCbyConstraint ( \41840_nR23900 , \41839 , \21944 );
buf \U$34150 ( \41841 , \41840_nR23900 );
not \U$34151 ( \41842 , \41306 );
and \U$34152 ( \41843 , RIe1e1bf8_5501, \41842 );
not \U$34153 ( \41844 , RIe1e1bf8_5501);
or \U$34154 ( \41845 , \41844 , \41745 );
nand \U$34155 ( \41846 , \38384 , \41609 );
nand \U$34156 ( \41847 , \38387 , \41612 );
nand \U$34157 ( \41848 , \41845 , \41846 , \41847 );
and \U$34158 ( \41849 , \41848 , \41306 );
or \U$34159 ( \41850 , \41843 , \41849 );
and \U$34161 ( \41851 , \41850 , 1'b1 );
or \U$34163 ( \41852 , \41851 , 1'b0 );
buf \U$34164 ( \41853 , \41852 );
_DC r23902_GF_IsGateDCbyConstraint ( \41854_nR23902 , \41853 , \21944 );
buf \U$34165 ( \41855 , \41854_nR23902 );
not \U$34166 ( \41856 , \39411 );
and \U$34167 ( \41857 , RIe1e23f0_5502, \41856 );
not \U$34168 ( \41858 , RIe1e23f0_5502);
or \U$34169 ( \41859 , \41858 , \41658 );
nand \U$34170 ( \41860 , \38403 , \41627 );
nand \U$34171 ( \41861 , \38406 , \41661 );
nand \U$34172 ( \41862 , \41859 , \41860 , \41861 );
and \U$34173 ( \41863 , \41862 , \39411 );
or \U$34174 ( \41864 , \41857 , \41863 );
and \U$34176 ( \41865 , \41864 , 1'b1 );
or \U$34178 ( \41866 , \41865 , 1'b0 );
buf \U$34179 ( \41867 , \41866 );
_DC r23904_GF_IsGateDCbyConstraint ( \41868_nR23904 , \41867 , \21944 );
buf \U$34180 ( \41869 , \41868_nR23904 );
not \U$34181 ( \41870 , \41494 );
and \U$34182 ( \41871 , RIe1e2be8_5503, \41870 );
not \U$34183 ( \41872 , RIe1e2be8_5503);
or \U$34184 ( \41873 , \41872 , \41641 );
nand \U$34185 ( \41874 , \38423 , \41609 );
nand \U$34186 ( \41875 , \38425 , \41661 );
nand \U$34187 ( \41876 , \41873 , \41874 , \41875 );
and \U$34188 ( \41877 , \41876 , \41494 );
or \U$34189 ( \41878 , \41871 , \41877 );
and \U$34191 ( \41879 , \41878 , 1'b1 );
or \U$34193 ( \41880 , \41879 , 1'b0 );
buf \U$34194 ( \41881 , \41880 );
_DC r23906_GF_IsGateDCbyConstraint ( \41882_nR23906 , \41881 , \21944 );
buf \U$34195 ( \41883 , \41882_nR23906 );
not \U$34196 ( \41884 , \39066 );
and \U$34197 ( \41885 , RIe1e33e0_5504, \41884 );
not \U$34198 ( \41886 , RIe1e33e0_5504);
or \U$34199 ( \41887 , \41886 , \41641 );
nand \U$34200 ( \41888 , \38441 , \41643 );
nand \U$34201 ( \41889 , \38443 , \41645 );
nand \U$34202 ( \41890 , \41887 , \41888 , \41889 );
and \U$34203 ( \41891 , \41890 , \39066 );
or \U$34204 ( \41892 , \41885 , \41891 );
and \U$34206 ( \41893 , \41892 , 1'b1 );
or \U$34208 ( \41894 , \41893 , 1'b0 );
buf \U$34209 ( \41895 , \41894 );
_DC r23908_GF_IsGateDCbyConstraint ( \41896_nR23908 , \41895 , \21944 );
buf \U$34210 ( \41897 , \41896_nR23908 );
not \U$34211 ( \41898 , \39411 );
and \U$34212 ( \41899 , RIe1e3bd8_5505, \41898 );
not \U$34213 ( \41900 , RIe1e3bd8_5505);
or \U$34214 ( \41901 , \41900 , \41745 );
nand \U$34215 ( \41902 , \38459 , \41609 );
nand \U$34216 ( \41903 , \38462 , \41645 );
nand \U$34217 ( \41904 , \41901 , \41902 , \41903 );
and \U$34218 ( \41905 , \41904 , \39411 );
or \U$34219 ( \41906 , \41899 , \41905 );
and \U$34221 ( \41907 , \41906 , 1'b1 );
or \U$34223 ( \41908 , \41907 , 1'b0 );
buf \U$34224 ( \41909 , \41908 );
_DC r2390c_GF_IsGateDCbyConstraint ( \41910_nR2390c , \41909 , \21944 );
buf \U$34225 ( \41911 , \41910_nR2390c );
not \U$34226 ( \41912 , \41494 );
and \U$34227 ( \41913 , RIe1e43d0_5506, \41912 );
not \U$34228 ( \41914 , RIe1e43d0_5506);
or \U$34229 ( \41915 , \41914 , \41745 );
nand \U$34230 ( \41916 , \38478 , \41817 );
nand \U$34231 ( \41917 , \38481 , \41690 );
nand \U$34232 ( \41918 , \41915 , \41916 , \41917 );
and \U$34233 ( \41919 , \41918 , \41494 );
or \U$34234 ( \41920 , \41913 , \41919 );
and \U$34236 ( \41921 , \41920 , 1'b1 );
or \U$34238 ( \41922 , \41921 , 1'b0 );
buf \U$34239 ( \41923 , \41922 );
_DC r2390e_GF_IsGateDCbyConstraint ( \41924_nR2390e , \41923 , \21944 );
buf \U$34240 ( \41925 , \41924_nR2390e );
not \U$34241 ( \41926 , \38705 );
and \U$34242 ( \41927 , RIe1e4bc8_5507, \41926 );
not \U$34243 ( \41928 , RIe1e4bc8_5507);
or \U$34244 ( \41929 , \41928 , \41625 );
nand \U$34245 ( \41930 , \38497 , \41817 );
nand \U$34246 ( \41931 , \38500 , \41612 );
nand \U$34247 ( \41932 , \41929 , \41930 , \41931 );
and \U$34248 ( \41933 , \41932 , \38705 );
or \U$34249 ( \41934 , \41927 , \41933 );
and \U$34251 ( \41935 , \41934 , 1'b1 );
or \U$34253 ( \41936 , \41935 , 1'b0 );
buf \U$34254 ( \41937 , \41936 );
_DC r23910_GF_IsGateDCbyConstraint ( \41938_nR23910 , \41937 , \21944 );
buf \U$34255 ( \41939 , \41938_nR23910 );
not \U$34256 ( \41940 , \39411 );
and \U$34257 ( \41941 , RIe1e53c0_5508, \41940 );
not \U$34258 ( \41942 , RIe1e53c0_5508);
or \U$34259 ( \41943 , \41942 , \41658 );
nand \U$34260 ( \41944 , \38516 , \41817 );
nand \U$34261 ( \41945 , \38518 , \41645 );
nand \U$34262 ( \41946 , \41943 , \41944 , \41945 );
and \U$34263 ( \41947 , \41946 , \39411 );
or \U$34264 ( \41948 , \41941 , \41947 );
and \U$34266 ( \41949 , \41948 , 1'b1 );
or \U$34268 ( \41950 , \41949 , 1'b0 );
buf \U$34269 ( \41951 , \41950 );
_DC r23912_GF_IsGateDCbyConstraint ( \41952_nR23912 , \41951 , \21944 );
buf \U$34270 ( \41953 , \41952_nR23912 );
not \U$34271 ( \41954 , \41494 );
and \U$34272 ( \41955 , RIe1e5bb8_5509, \41954 );
not \U$34273 ( \41956 , RIe1e5bb8_5509);
or \U$34274 ( \41957 , \41956 , \41641 );
nand \U$34275 ( \41958 , \38534 , \41609 );
nand \U$34276 ( \41959 , \38537 , \41661 );
nand \U$34277 ( \41960 , \41957 , \41958 , \41959 );
and \U$34278 ( \41961 , \41960 , \41494 );
or \U$34279 ( \41962 , \41955 , \41961 );
and \U$34281 ( \41963 , \41962 , 1'b1 );
or \U$34283 ( \41964 , \41963 , 1'b0 );
buf \U$34284 ( \41965 , \41964 );
_DC r23914_GF_IsGateDCbyConstraint ( \41966_nR23914 , \41965 , \21944 );
buf \U$34285 ( \41967 , \41966_nR23914 );
not \U$34286 ( \41968 , \38705 );
and \U$34287 ( \41969 , RIe1e63b0_5510, \41968 );
not \U$34288 ( \41970 , RIe1e63b0_5510);
or \U$34289 ( \41971 , \41970 , \41625 );
nand \U$34290 ( \41972 , \38553 , \41817 );
nand \U$34291 ( \41973 , \38555 , \41690 );
nand \U$34292 ( \41974 , \41971 , \41972 , \41973 );
and \U$34293 ( \41975 , \41974 , \38705 );
or \U$34294 ( \41976 , \41969 , \41975 );
and \U$34296 ( \41977 , \41976 , 1'b1 );
or \U$34298 ( \41978 , \41977 , 1'b0 );
buf \U$34299 ( \41979 , \41978 );
_DC r23916_GF_IsGateDCbyConstraint ( \41980_nR23916 , \41979 , \21944 );
buf \U$34300 ( \41981 , \41980_nR23916 );
not \U$34301 ( \41982 , \39411 );
and \U$34302 ( \41983 , RIe1e6ba8_5511, \41982 );
not \U$34303 ( \41984 , RIe1e6ba8_5511);
or \U$34304 ( \41985 , \41984 , \41625 );
nand \U$34305 ( \41986 , \38571 , \41643 );
nand \U$34306 ( \41987 , \38573 , \41690 );
nand \U$34307 ( \41988 , \41985 , \41986 , \41987 );
and \U$34308 ( \41989 , \41988 , \39411 );
or \U$34309 ( \41990 , \41983 , \41989 );
and \U$34311 ( \41991 , \41990 , 1'b1 );
or \U$34313 ( \41992 , \41991 , 1'b0 );
buf \U$34314 ( \41993 , \41992 );
_DC r23918_GF_IsGateDCbyConstraint ( \41994_nR23918 , \41993 , \21944 );
buf \U$34315 ( \41995 , \41994_nR23918 );
not \U$34316 ( \41996 , \41494 );
and \U$34317 ( \41997 , RIe1e73a0_5512, \41996 );
not \U$34318 ( \41998 , RIe1e73a0_5512);
or \U$34319 ( \41999 , \41998 , \41745 );
nand \U$34320 ( \42000 , \38589 , \41609 );
nand \U$34321 ( \42001 , \38591 , \41612 );
nand \U$34322 ( \42002 , \41999 , \42000 , \42001 );
and \U$34323 ( \42003 , \42002 , \41494 );
or \U$34324 ( \42004 , \41997 , \42003 );
and \U$34326 ( \42005 , \42004 , 1'b1 );
or \U$34328 ( \42006 , \42005 , 1'b0 );
buf \U$34329 ( \42007 , \42006 );
_DC r2391a_GF_IsGateDCbyConstraint ( \42008_nR2391a , \42007 , \21944 );
buf \U$34330 ( \42009 , \42008_nR2391a );
not \U$34331 ( \42010 , \39163 );
and \U$34332 ( \42011 , RIe1e7b98_5513, \42010 );
not \U$34333 ( \42012 , RIe1e7b98_5513);
or \U$34334 ( \42013 , \42012 , \41745 );
nand \U$34335 ( \42014 , \38609 , \41643 );
nand \U$34336 ( \42015 , \38612 , \41661 );
nand \U$34337 ( \42016 , \42013 , \42014 , \42015 );
and \U$34338 ( \42017 , \42016 , \39163 );
or \U$34339 ( \42018 , \42011 , \42017 );
and \U$34341 ( \42019 , \42018 , 1'b1 );
or \U$34343 ( \42020 , \42019 , 1'b0 );
buf \U$34344 ( \42021 , \42020 );
_DC r2391c_GF_IsGateDCbyConstraint ( \42022_nR2391c , \42021 , \21944 );
buf \U$34345 ( \42023 , \42022_nR2391c );
not \U$34346 ( \42024 , \39411 );
and \U$34347 ( \42025 , RIe1e8390_5514, \42024 );
not \U$34348 ( \42026 , RIe1e8390_5514);
or \U$34349 ( \42027 , \42026 , \41658 );
nand \U$34350 ( \42028 , \38630 , \41817 );
nand \U$34351 ( \42029 , \38633 , \41612 );
nand \U$34352 ( \42030 , \42027 , \42028 , \42029 );
and \U$34353 ( \42031 , \42030 , \39411 );
or \U$34354 ( \42032 , \42025 , \42031 );
and \U$34356 ( \42033 , \42032 , 1'b1 );
or \U$34358 ( \42034 , \42033 , 1'b0 );
buf \U$34359 ( \42035 , \42034 );
_DC r2391e_GF_IsGateDCbyConstraint ( \42036_nR2391e , \42035 , \21944 );
buf \U$34360 ( \42037 , \42036_nR2391e );
buf \U$34361 ( \42038 , \39066 );
not \U$34362 ( \42039 , \42038 );
and \U$34363 ( \42040 , RIe1e8b88_5515, \42039 );
not \U$34364 ( \42041 , RIe1e8b88_5515);
or \U$34365 ( \42042 , \42041 , \41625 );
nand \U$34366 ( \42043 , \38650 , \41817 );
nand \U$34367 ( \42044 , \38653 , \41661 );
nand \U$34368 ( \42045 , \42042 , \42043 , \42044 );
and \U$34369 ( \42046 , \42045 , \42038 );
or \U$34370 ( \42047 , \42040 , \42046 );
and \U$34372 ( \42048 , \42047 , 1'b1 );
or \U$34374 ( \42049 , \42048 , 1'b0 );
buf \U$34375 ( \42050 , \42049 );
_DC r23922_GF_IsGateDCbyConstraint ( \42051_nR23922 , \42050 , \21944 );
buf \U$34376 ( \42052 , \42051_nR23922 );
not \U$34377 ( \42053 , \39411 );
and \U$34378 ( \42054 , RIe1e9380_5516, \42053 );
not \U$34379 ( \42055 , RIe1e9380_5516);
or \U$34380 ( \42056 , \42055 , \41745 );
nand \U$34381 ( \42057 , \38670 , \41817 );
nand \U$34382 ( \42058 , \38673 , \41612 );
nand \U$34383 ( \42059 , \42056 , \42057 , \42058 );
and \U$34384 ( \42060 , \42059 , \39411 );
or \U$34385 ( \42061 , \42054 , \42060 );
and \U$34387 ( \42062 , \42061 , 1'b1 );
or \U$34389 ( \42063 , \42062 , 1'b0 );
buf \U$34390 ( \42064 , \42063 );
_DC r23924_GF_IsGateDCbyConstraint ( \42065_nR23924 , \42064 , \21944 );
buf \U$34391 ( \42066 , \42065_nR23924 );
not \U$34392 ( \42067 , \39411 );
and \U$34393 ( \42068 , RIe1e9b78_5517, \42067 );
not \U$34394 ( \42069 , RIe1e9b78_5517);
or \U$34395 ( \42070 , \42069 , \41625 );
nand \U$34396 ( \42071 , \38690 , \41609 );
nand \U$34397 ( \42072 , \38693 , \41690 );
nand \U$34398 ( \42073 , \42070 , \42071 , \42072 );
and \U$34399 ( \42074 , \42073 , \39411 );
or \U$34400 ( \42075 , \42068 , \42074 );
and \U$34402 ( \42076 , \42075 , 1'b1 );
or \U$34404 ( \42077 , \42076 , 1'b0 );
buf \U$34405 ( \42078 , \42077 );
_DC r23926_GF_IsGateDCbyConstraint ( \42079_nR23926 , \42078 , \21944 );
buf \U$34406 ( \42080 , \42079_nR23926 );
not \U$34407 ( \42081 , \42038 );
and \U$34408 ( \42082 , RIe1ea370_5518, \42081 );
not \U$34409 ( \42083 , RIe1ea370_5518);
or \U$34410 ( \42084 , \42083 , \41745 );
nand \U$34411 ( \42085 , \38710 , \41643 );
nand \U$34412 ( \42086 , \38713 , \41645 );
nand \U$34413 ( \42087 , \42084 , \42085 , \42086 );
and \U$34414 ( \42088 , \42087 , \42038 );
or \U$34415 ( \42089 , \42082 , \42088 );
and \U$34417 ( \42090 , \42089 , 1'b1 );
or \U$34419 ( \42091 , \42090 , 1'b0 );
buf \U$34420 ( \42092 , \42091 );
_DC r23928_GF_IsGateDCbyConstraint ( \42093_nR23928 , \42092 , \21944 );
buf \U$34421 ( \42094 , \42093_nR23928 );
not \U$34422 ( \42095 , \39163 );
and \U$34423 ( \42096 , RIe1eab68_5519, \42095 );
not \U$34424 ( \42097 , RIe1eab68_5519);
or \U$34425 ( \42098 , \42097 , \41658 );
nand \U$34426 ( \42099 , \38731 , \41643 );
nand \U$34427 ( \42100 , \38734 , \41690 );
nand \U$34428 ( \42101 , \42098 , \42099 , \42100 );
and \U$34429 ( \42102 , \42101 , \39163 );
or \U$34430 ( \42103 , \42096 , \42102 );
and \U$34432 ( \42104 , \42103 , 1'b1 );
or \U$34434 ( \42105 , \42104 , 1'b0 );
buf \U$34435 ( \42106 , \42105 );
_DC r2392a_GF_IsGateDCbyConstraint ( \42107_nR2392a , \42106 , \21944 );
buf \U$34436 ( \42108 , \42107_nR2392a );
not \U$34437 ( \42109 , \39411 );
and \U$34438 ( \42110 , RIe1eb360_5520, \42109 );
not \U$34439 ( \42111 , RIe1eb360_5520);
or \U$34440 ( \42112 , \42111 , \41641 );
nand \U$34441 ( \42113 , \38752 , \41627 );
nand \U$34442 ( \42114 , \38754 , \41661 );
nand \U$34443 ( \42115 , \42112 , \42113 , \42114 );
and \U$34444 ( \42116 , \42115 , \39411 );
or \U$34445 ( \42117 , \42110 , \42116 );
and \U$34447 ( \42118 , \42117 , 1'b1 );
or \U$34449 ( \42119 , \42118 , 1'b0 );
buf \U$34450 ( \42120 , \42119 );
_DC r2392c_GF_IsGateDCbyConstraint ( \42121_nR2392c , \42120 , \21944 );
buf \U$34451 ( \42122 , \42121_nR2392c );
not \U$34452 ( \42123 , \42038 );
and \U$34453 ( \42124 , RIe1ebb58_5521, \42123 );
not \U$34454 ( \42125 , RIe1ebb58_5521);
or \U$34455 ( \42126 , \42125 , \41658 );
nand \U$34456 ( \42127 , \38771 , \41627 );
nand \U$34457 ( \42128 , \38773 , \41645 );
nand \U$34458 ( \42129 , \42126 , \42127 , \42128 );
and \U$34459 ( \42130 , \42129 , \42038 );
or \U$34460 ( \42131 , \42124 , \42130 );
and \U$34462 ( \42132 , \42131 , 1'b1 );
or \U$34464 ( \42133 , \42132 , 1'b0 );
buf \U$34465 ( \42134 , \42133 );
_DC r2392e_GF_IsGateDCbyConstraint ( \42135_nR2392e , \42134 , \21944 );
buf \U$34466 ( \42136 , \42135_nR2392e );
not \U$34467 ( \42137 , \39163 );
and \U$34468 ( \42138 , RIe1ec350_5522, \42137 );
not \U$34469 ( \42139 , RIe1ec350_5522);
or \U$34470 ( \42140 , \42139 , \41625 );
nand \U$34471 ( \42141 , \38789 , \41609 );
nand \U$34472 ( \42142 , \38792 , \41690 );
nand \U$34473 ( \42143 , \42140 , \42141 , \42142 );
and \U$34474 ( \42144 , \42143 , \39163 );
or \U$34475 ( \42145 , \42138 , \42144 );
and \U$34477 ( \42146 , \42145 , 1'b1 );
or \U$34479 ( \42147 , \42146 , 1'b0 );
buf \U$34480 ( \42148 , \42147 );
_DC r23930_GF_IsGateDCbyConstraint ( \42149_nR23930 , \42148 , \21944 );
buf \U$34481 ( \42150 , \42149_nR23930 );
not \U$34482 ( \42151 , \39411 );
and \U$34483 ( \42152 , RIe1ecb48_5523, \42151 );
not \U$34484 ( \42153 , RIe1ecb48_5523);
or \U$34485 ( \42154 , \42153 , \41745 );
nand \U$34486 ( \42155 , \38808 , \41609 );
nand \U$34487 ( \42156 , \38810 , \41612 );
nand \U$34488 ( \42157 , \42154 , \42155 , \42156 );
and \U$34489 ( \42158 , \42157 , \39411 );
or \U$34490 ( \42159 , \42152 , \42158 );
and \U$34492 ( \42160 , \42159 , 1'b1 );
or \U$34494 ( \42161 , \42160 , 1'b0 );
buf \U$34495 ( \42162 , \42161 );
_DC r23932_GF_IsGateDCbyConstraint ( \42163_nR23932 , \42162 , \21944 );
buf \U$34496 ( \42164 , \42163_nR23932 );
not \U$34497 ( \42165 , \42038 );
and \U$34498 ( \42166 , RIe1ed340_5524, \42165 );
not \U$34499 ( \42167 , RIe1ed340_5524);
or \U$34500 ( \42168 , \42167 , \41745 );
nand \U$34501 ( \42169 , \38827 , \41817 );
nand \U$34502 ( \42170 , \38829 , \41645 );
nand \U$34503 ( \42171 , \42168 , \42169 , \42170 );
and \U$34504 ( \42172 , \42171 , \42038 );
or \U$34505 ( \42173 , \42166 , \42172 );
and \U$34507 ( \42174 , \42173 , 1'b1 );
or \U$34509 ( \42175 , \42174 , 1'b0 );
buf \U$34510 ( \42176 , \42175 );
_DC r23934_GF_IsGateDCbyConstraint ( \42177_nR23934 , \42176 , \21944 );
buf \U$34511 ( \42178 , \42177_nR23934 );
not \U$34512 ( \42179 , \39066 );
and \U$34513 ( \42180 , RIe1edb38_5525, \42179 );
not \U$34514 ( \42181 , RIe1edb38_5525);
or \U$34515 ( \42182 , \42181 , \41641 );
nand \U$34516 ( \42183 , \38845 , \41627 );
nand \U$34517 ( \42184 , \38847 , \41661 );
nand \U$34518 ( \42185 , \42182 , \42183 , \42184 );
and \U$34519 ( \42186 , \42185 , \39066 );
or \U$34520 ( \42187 , \42180 , \42186 );
and \U$34522 ( \42188 , \42187 , 1'b1 );
or \U$34524 ( \42189 , \42188 , 1'b0 );
buf \U$34525 ( \42190 , \42189 );
_DC r23938_GF_IsGateDCbyConstraint ( \42191_nR23938 , \42190 , \21944 );
buf \U$34526 ( \42192 , \42191_nR23938 );
not \U$34527 ( \42193 , \39411 );
and \U$34528 ( \42194 , RIe1ee330_5526, \42193 );
not \U$34529 ( \42195 , RIe1ee330_5526);
or \U$34530 ( \42196 , \42195 , \41641 );
nand \U$34531 ( \42197 , \38863 , \41627 );
nand \U$34532 ( \42198 , \38865 , \41690 );
nand \U$34533 ( \42199 , \42196 , \42197 , \42198 );
and \U$34534 ( \42200 , \42199 , \39411 );
or \U$34535 ( \42201 , \42194 , \42200 );
and \U$34537 ( \42202 , \42201 , 1'b1 );
or \U$34539 ( \42203 , \42202 , 1'b0 );
buf \U$34540 ( \42204 , \42203 );
_DC r2393a_GF_IsGateDCbyConstraint ( \42205_nR2393a , \42204 , \21944 );
buf \U$34541 ( \42206 , \42205_nR2393a );
not \U$34542 ( \42207 , \42038 );
and \U$34543 ( \42208 , RIe1eeb28_5527, \42207 );
not \U$34544 ( \42209 , RIe1eeb28_5527);
or \U$34545 ( \42210 , \42209 , \41625 );
nand \U$34546 ( \42211 , \38881 , \41609 );
nand \U$34547 ( \42212 , \38883 , \41612 );
nand \U$34548 ( \42213 , \42210 , \42211 , \42212 );
and \U$34549 ( \42214 , \42213 , \42038 );
or \U$34550 ( \42215 , \42208 , \42214 );
and \U$34552 ( \42216 , \42215 , 1'b1 );
or \U$34554 ( \42217 , \42216 , 1'b0 );
buf \U$34555 ( \42218 , \42217 );
_DC r2393c_GF_IsGateDCbyConstraint ( \42219_nR2393c , \42218 , \21944 );
buf \U$34556 ( \42220 , \42219_nR2393c );
not \U$34557 ( \42221 , \38705 );
and \U$34558 ( \42222 , RIe1ef320_5528, \42221 );
not \U$34559 ( \42223 , RIe1ef320_5528);
or \U$34560 ( \42224 , \42223 , \41641 );
nand \U$34561 ( \42225 , \38899 , \41627 );
nand \U$34562 ( \42226 , \38902 , \41612 );
nand \U$34563 ( \42227 , \42224 , \42225 , \42226 );
and \U$34564 ( \42228 , \42227 , \38705 );
or \U$34565 ( \42229 , \42222 , \42228 );
and \U$34567 ( \42230 , \42229 , 1'b1 );
or \U$34569 ( \42231 , \42230 , 1'b0 );
buf \U$34570 ( \42232 , \42231 );
_DC r2393e_GF_IsGateDCbyConstraint ( \42233_nR2393e , \42232 , \21944 );
buf \U$34571 ( \42234 , \42233_nR2393e );
not \U$34572 ( \42235 , \39411 );
and \U$34573 ( \42236 , RIe1efb18_5529, \42235 );
not \U$34574 ( \42237 , RIe1efb18_5529);
or \U$34575 ( \42238 , \42237 , \41745 );
nand \U$34576 ( \42239 , \38919 , \41627 );
nand \U$34577 ( \42240 , \38921 , \41661 );
nand \U$34578 ( \42241 , \42238 , \42239 , \42240 );
and \U$34579 ( \42242 , \42241 , \39411 );
or \U$34580 ( \42243 , \42236 , \42242 );
and \U$34582 ( \42244 , \42243 , 1'b1 );
or \U$34584 ( \42245 , \42244 , 1'b0 );
buf \U$34585 ( \42246 , \42245 );
_DC r23940_GF_IsGateDCbyConstraint ( \42247_nR23940 , \42246 , \21944 );
buf \U$34586 ( \42248 , \42247_nR23940 );
not \U$34587 ( \42249 , \42038 );
and \U$34588 ( \42250 , RIe1f0310_5530, \42249 );
not \U$34589 ( \42251 , RIe1f0310_5530);
or \U$34590 ( \42252 , \42251 , \41625 );
nand \U$34591 ( \42253 , \38937 , \41627 );
nand \U$34592 ( \42254 , \38940 , \41645 );
nand \U$34593 ( \42255 , \42252 , \42253 , \42254 );
and \U$34594 ( \42256 , \42255 , \42038 );
or \U$34595 ( \42257 , \42250 , \42256 );
and \U$34597 ( \42258 , \42257 , 1'b1 );
or \U$34599 ( \42259 , \42258 , 1'b0 );
buf \U$34600 ( \42260 , \42259 );
_DC r23942_GF_IsGateDCbyConstraint ( \42261_nR23942 , \42260 , \21944 );
buf \U$34601 ( \42262 , \42261_nR23942 );
not \U$34602 ( \42263 , \39163 );
and \U$34603 ( \42264 , RIe1f0b08_5531, \42263 );
not \U$34604 ( \42265 , RIe1f0b08_5531);
or \U$34605 ( \42266 , \42265 , \41658 );
nand \U$34606 ( \42267 , \38956 , \41627 );
nand \U$34607 ( \42268 , \38958 , \41645 );
nand \U$34608 ( \42269 , \42266 , \42267 , \42268 );
and \U$34609 ( \42270 , \42269 , \39163 );
or \U$34610 ( \42271 , \42264 , \42270 );
and \U$34612 ( \42272 , \42271 , 1'b1 );
or \U$34614 ( \42273 , \42272 , 1'b0 );
buf \U$34615 ( \42274 , \42273 );
_DC r23944_GF_IsGateDCbyConstraint ( \42275_nR23944 , \42274 , \21944 );
buf \U$34616 ( \42276 , \42275_nR23944 );
not \U$34617 ( \42277 , \39411 );
and \U$34618 ( \42278 , RIe1f1300_5532, \42277 );
not \U$34619 ( \42279 , RIe1f1300_5532);
or \U$34620 ( \42280 , \42279 , \41641 );
nand \U$34621 ( \42281 , \38974 , \41817 );
nand \U$34622 ( \42282 , \38977 , \41612 );
nand \U$34623 ( \42283 , \42280 , \42281 , \42282 );
and \U$34624 ( \42284 , \42283 , \39411 );
or \U$34625 ( \42285 , \42278 , \42284 );
and \U$34627 ( \42286 , \42285 , 1'b1 );
or \U$34629 ( \42287 , \42286 , 1'b0 );
buf \U$34630 ( \42288 , \42287 );
_DC r23946_GF_IsGateDCbyConstraint ( \42289_nR23946 , \42288 , \21944 );
buf \U$34631 ( \42290 , \42289_nR23946 );
not \U$34632 ( \42291 , \42038 );
and \U$34633 ( \42292 , RIe1f1af8_5533, \42291 );
not \U$34634 ( \42293 , RIe1f1af8_5533);
or \U$34635 ( \42294 , \42293 , \41625 );
nand \U$34636 ( \42295 , \38993 , \41817 );
nand \U$34637 ( \42296 , \38995 , \41690 );
nand \U$34638 ( \42297 , \42294 , \42295 , \42296 );
and \U$34639 ( \42298 , \42297 , \42038 );
or \U$34640 ( \42299 , \42292 , \42298 );
and \U$34642 ( \42300 , \42299 , 1'b1 );
or \U$34644 ( \42301 , \42300 , 1'b0 );
buf \U$34645 ( \42302 , \42301 );
_DC r23948_GF_IsGateDCbyConstraint ( \42303_nR23948 , \42302 , \21944 );
buf \U$34646 ( \42304 , \42303_nR23948 );
not \U$34647 ( \42305 , \38033 );
and \U$34648 ( \42306 , RIe1f22f0_5534, \42305 );
not \U$34649 ( \42307 , RIe1f22f0_5534);
or \U$34650 ( \42308 , \42307 , \41658 );
nand \U$34651 ( \42309 , \39011 , \41643 );
nand \U$34652 ( \42310 , \39014 , \41690 );
nand \U$34653 ( \42311 , \42308 , \42309 , \42310 );
and \U$34654 ( \42312 , \42311 , \38033 );
or \U$34655 ( \42313 , \42306 , \42312 );
and \U$34657 ( \42314 , \42313 , 1'b1 );
or \U$34659 ( \42315 , \42314 , 1'b0 );
buf \U$34660 ( \42316 , \42315 );
_DC r2394a_GF_IsGateDCbyConstraint ( \42317_nR2394a , \42316 , \21944 );
buf \U$34661 ( \42318 , \42317_nR2394a );
not \U$34662 ( \42319 , \39411 );
and \U$34663 ( \42320 , RIe1f2ae8_5535, \42319 );
not \U$34664 ( \42321 , RIe1f2ae8_5535);
or \U$34665 ( \42322 , \42321 , \41745 );
nand \U$34666 ( \42323 , \39030 , \41609 );
nand \U$34667 ( \42324 , \39033 , \41661 );
nand \U$34668 ( \42325 , \42322 , \42323 , \42324 );
and \U$34669 ( \42326 , \42325 , \39411 );
or \U$34670 ( \42327 , \42320 , \42326 );
and \U$34672 ( \42328 , \42327 , 1'b1 );
or \U$34674 ( \42329 , \42328 , 1'b0 );
buf \U$34675 ( \42330 , \42329 );
_DC r2394e_GF_IsGateDCbyConstraint ( \42331_nR2394e , \42330 , \21944 );
buf \U$34676 ( \42332 , \42331_nR2394e );
not \U$34677 ( \42333 , \42038 );
and \U$34678 ( \42334 , RIe1f32e0_5536, \42333 );
not \U$34679 ( \42335 , RIe1f32e0_5536);
or \U$34680 ( \42336 , \42335 , \41658 );
nand \U$34681 ( \42337 , \39051 , \41817 );
nand \U$34682 ( \42338 , \39054 , \41661 );
nand \U$34683 ( \42339 , \42336 , \42337 , \42338 );
and \U$34684 ( \42340 , \42339 , \42038 );
or \U$34685 ( \42341 , \42334 , \42340 );
and \U$34687 ( \42342 , \42341 , 1'b1 );
or \U$34689 ( \42343 , \42342 , 1'b0 );
buf \U$34690 ( \42344 , \42343 );
_DC r23950_GF_IsGateDCbyConstraint ( \42345_nR23950 , \42344 , \21944 );
buf \U$34691 ( \42346 , \42345_nR23950 );
not \U$34692 ( \42347 , \39066 );
and \U$34693 ( \42348 , RIe1f3ad8_5537, \42347 );
not \U$34694 ( \42349 , RIe1f3ad8_5537);
or \U$34695 ( \42350 , \42349 , \41641 );
nand \U$34696 ( \42351 , \39071 , \41627 );
nand \U$34697 ( \42352 , \39074 , \41690 );
nand \U$34698 ( \42353 , \42350 , \42351 , \42352 );
and \U$34699 ( \42354 , \42353 , \39066 );
or \U$34700 ( \42355 , \42348 , \42354 );
and \U$34702 ( \42356 , \42355 , 1'b1 );
or \U$34704 ( \42357 , \42356 , 1'b0 );
buf \U$34705 ( \42358 , \42357 );
_DC r23952_GF_IsGateDCbyConstraint ( \42359_nR23952 , \42358 , \21944 );
buf \U$34706 ( \42360 , \42359_nR23952 );
not \U$34707 ( \42361 , \39045 );
and \U$34708 ( \42362 , RIe1f42d0_5538, \42361 );
not \U$34709 ( \42363 , RIe1f42d0_5538);
or \U$34710 ( \42364 , \42363 , \41625 );
nand \U$34711 ( \42365 , \39090 , \41817 );
nand \U$34712 ( \42366 , \39093 , \41612 );
nand \U$34713 ( \42367 , \42364 , \42365 , \42366 );
and \U$34714 ( \42368 , \42367 , \39045 );
or \U$34715 ( \42369 , \42362 , \42368 );
and \U$34717 ( \42370 , \42369 , 1'b1 );
or \U$34719 ( \42371 , \42370 , 1'b0 );
buf \U$34720 ( \42372 , \42371 );
_DC r23954_GF_IsGateDCbyConstraint ( \42373_nR23954 , \42372 , \21944 );
buf \U$34721 ( \42374 , \42373_nR23954 );
not \U$34722 ( \42375 , \42038 );
and \U$34723 ( \42376 , RIe1f4ac8_5539, \42375 );
not \U$34724 ( \42377 , RIe1f4ac8_5539);
or \U$34725 ( \42378 , \42377 , \41745 );
nand \U$34726 ( \42379 , \39109 , \41609 );
nand \U$34727 ( \42380 , \39112 , \41612 );
nand \U$34728 ( \42381 , \42378 , \42379 , \42380 );
and \U$34729 ( \42382 , \42381 , \42038 );
or \U$34730 ( \42383 , \42376 , \42382 );
and \U$34732 ( \42384 , \42383 , 1'b1 );
or \U$34734 ( \42385 , \42384 , 1'b0 );
buf \U$34735 ( \42386 , \42385 );
_DC r23956_GF_IsGateDCbyConstraint ( \42387_nR23956 , \42386 , \21944 );
buf \U$34736 ( \42388 , \42387_nR23956 );
not \U$34737 ( \42389 , \38117 );
and \U$34738 ( \42390 , RIe1f52c0_5540, \42389 );
not \U$34739 ( \42391 , RIe1f52c0_5540);
or \U$34740 ( \42392 , \42391 , \41745 );
nand \U$34741 ( \42393 , \39128 , \41817 );
nand \U$34742 ( \42394 , \39131 , \41661 );
nand \U$34743 ( \42395 , \42392 , \42393 , \42394 );
and \U$34744 ( \42396 , \42395 , \38117 );
or \U$34745 ( \42397 , \42390 , \42396 );
and \U$34747 ( \42398 , \42397 , 1'b1 );
or \U$34749 ( \42399 , \42398 , 1'b0 );
buf \U$34750 ( \42400 , \42399 );
_DC r23958_GF_IsGateDCbyConstraint ( \42401_nR23958 , \42400 , \21944 );
buf \U$34751 ( \42402 , \42401_nR23958 );
not \U$34752 ( \42403 , \39163 );
and \U$34753 ( \42404 , RIe1f5ab8_5541, \42403 );
not \U$34754 ( \42405 , RIe1f5ab8_5541);
or \U$34755 ( \42406 , \42405 , \41745 );
nand \U$34756 ( \42407 , \39148 , \41627 );
nand \U$34757 ( \42408 , \39151 , \41645 );
nand \U$34758 ( \42409 , \42406 , \42407 , \42408 );
and \U$34759 ( \42410 , \42409 , \39163 );
or \U$34760 ( \42411 , \42404 , \42410 );
and \U$34762 ( \42412 , \42411 , 1'b1 );
or \U$34764 ( \42413 , \42412 , 1'b0 );
buf \U$34765 ( \42414 , \42413 );
_DC r2395a_GF_IsGateDCbyConstraint ( \42415_nR2395a , \42414 , \21944 );
buf \U$34766 ( \42416 , \42415_nR2395a );
not \U$34767 ( \42417 , \42038 );
and \U$34768 ( \42418 , RIe1f62b0_5542, \42417 );
not \U$34769 ( \42419 , RIe1f62b0_5542);
or \U$34770 ( \42420 , \42419 , \41658 );
nand \U$34771 ( \42421 , \39169 , \41817 );
nand \U$34772 ( \42422 , \39171 , \41645 );
nand \U$34773 ( \42423 , \42420 , \42421 , \42422 );
and \U$34774 ( \42424 , \42423 , \42038 );
or \U$34775 ( \42425 , \42418 , \42424 );
and \U$34777 ( \42426 , \42425 , 1'b1 );
or \U$34779 ( \42427 , \42426 , 1'b0 );
buf \U$34780 ( \42428 , \42427 );
_DC r2395c_GF_IsGateDCbyConstraint ( \42429_nR2395c , \42428 , \21944 );
buf \U$34781 ( \42430 , \42429_nR2395c );
not \U$34782 ( \42431 , \38117 );
and \U$34783 ( \42432 , RIe1f6aa8_5543, \42431 );
not \U$34784 ( \42433 , RIe1f6aa8_5543);
or \U$34785 ( \42434 , \42433 , \41641 );
nand \U$34786 ( \42435 , \39188 , \41609 );
nand \U$34787 ( \42436 , \39190 , \41612 );
nand \U$34788 ( \42437 , \42434 , \42435 , \42436 );
and \U$34789 ( \42438 , \42437 , \38117 );
or \U$34790 ( \42439 , \42432 , \42438 );
and \U$34792 ( \42440 , \42439 , 1'b1 );
or \U$34794 ( \42441 , \42440 , 1'b0 );
buf \U$34795 ( \42442 , \42441 );
_DC r2395e_GF_IsGateDCbyConstraint ( \42443_nR2395e , \42442 , \21944 );
buf \U$34796 ( \42444 , \42443_nR2395e );
not \U$34797 ( \42445 , \38033 );
and \U$34798 ( \42446 , RIe1f72a0_5544, \42445 );
not \U$34799 ( \42447 , RIe1f72a0_5544);
or \U$34800 ( \42448 , \42447 , \41658 );
nand \U$34801 ( \42449 , \39208 , \41609 );
nand \U$34802 ( \42450 , \39211 , \41690 );
nand \U$34803 ( \42451 , \42448 , \42449 , \42450 );
and \U$34804 ( \42452 , \42451 , \38033 );
or \U$34805 ( \42453 , \42446 , \42452 );
and \U$34807 ( \42454 , \42453 , 1'b1 );
or \U$34809 ( \42455 , \42454 , 1'b0 );
buf \U$34810 ( \42456 , \42455 );
_DC r23960_GF_IsGateDCbyConstraint ( \42457_nR23960 , \42456 , \21944 );
buf \U$34811 ( \42458 , \42457_nR23960 );
not \U$34812 ( \42459 , \42038 );
and \U$34813 ( \42460 , RIe1f7a98_5545, \42459 );
not \U$34814 ( \42461 , RIe1f7a98_5545);
or \U$34815 ( \42462 , \42461 , \41606 );
nand \U$34816 ( \42463 , \39227 , \41627 );
nand \U$34817 ( \42464 , \39230 , \41645 );
nand \U$34818 ( \42465 , \42462 , \42463 , \42464 );
and \U$34819 ( \42466 , \42465 , \42038 );
or \U$34820 ( \42467 , \42460 , \42466 );
and \U$34822 ( \42468 , \42467 , 1'b1 );
or \U$34824 ( \42469 , \42468 , 1'b0 );
buf \U$34825 ( \42470 , \42469 );
_DC r23964_GF_IsGateDCbyConstraint ( \42471_nR23964 , \42470 , \21944 );
buf \U$34826 ( \42472 , \42471_nR23964 );
not \U$34827 ( \42473 , \38117 );
and \U$34828 ( \42474 , RIe1f8290_5546, \42473 );
not \U$34829 ( \42475 , RIe1f8290_5546);
or \U$34830 ( \42476 , \42475 , \41745 );
nand \U$34831 ( \42477 , \39247 , \41627 );
nand \U$34832 ( \42478 , \39250 , \41661 );
nand \U$34833 ( \42479 , \42476 , \42477 , \42478 );
and \U$34834 ( \42480 , \42479 , \38117 );
or \U$34835 ( \42481 , \42474 , \42480 );
and \U$34837 ( \42482 , \42481 , 1'b1 );
or \U$34839 ( \42483 , \42482 , 1'b0 );
buf \U$34840 ( \42484 , \42483 );
_DC r23966_GF_IsGateDCbyConstraint ( \42485_nR23966 , \42484 , \21944 );
buf \U$34841 ( \42486 , \42485_nR23966 );
not \U$34842 ( \42487 , \38822 );
and \U$34843 ( \42488 , RIe1f8a88_5547, \42487 );
not \U$34844 ( \42489 , RIe1f8a88_5547);
or \U$34845 ( \42490 , \42489 , \41658 );
nand \U$34846 ( \42491 , \39266 , \41817 );
nand \U$34847 ( \42492 , \39269 , \41661 );
nand \U$34848 ( \42493 , \42490 , \42491 , \42492 );
and \U$34849 ( \42494 , \42493 , \38822 );
or \U$34850 ( \42495 , \42488 , \42494 );
and \U$34852 ( \42496 , \42495 , 1'b1 );
or \U$34854 ( \42497 , \42496 , 1'b0 );
buf \U$34855 ( \42498 , \42497 );
_DC r23968_GF_IsGateDCbyConstraint ( \42499_nR23968 , \42498 , \21944 );
buf \U$34856 ( \42500 , \42499_nR23968 );
not \U$34857 ( \42501 , \42038 );
and \U$34858 ( \42502 , RIe1f9280_5548, \42501 );
not \U$34859 ( \42503 , RIe1f9280_5548);
or \U$34860 ( \42504 , \42503 , \41641 );
nand \U$34861 ( \42505 , \39285 , \41817 );
nand \U$34862 ( \42506 , \39288 , \41690 );
nand \U$34863 ( \42507 , \42504 , \42505 , \42506 );
and \U$34864 ( \42508 , \42507 , \42038 );
or \U$34865 ( \42509 , \42502 , \42508 );
and \U$34867 ( \42510 , \42509 , 1'b1 );
or \U$34869 ( \42511 , \42510 , 1'b0 );
buf \U$34870 ( \42512 , \42511 );
_DC r2396a_GF_IsGateDCbyConstraint ( \42513_nR2396a , \42512 , \21944 );
buf \U$34871 ( \42514 , \42513_nR2396a );
nor \U$34872 ( \42515 , \38022 , \38031 );
not \U$34873 ( \42516 , \42515 );
not \U$34874 ( \42517 , \42516 );
not \U$34875 ( \42518 , \42517 );
and \U$34876 ( \42519 , RIe137870_5261, \42518 );
not \U$34877 ( \42520 , RIe137870_5261);
not \U$34878 ( \42521 , \42520 );
not \U$34879 ( \42522 , \38043 );
and \U$34880 ( \42523 , \42521 , \42522 );
buf \U$34881 ( \42524 , RIb86fc68_77);
buf \U$34882 ( \42525 , \42524 );
and \U$34883 ( \42526 , \42525 , \38043 );
or \U$34884 ( \42527 , \42523 , \42526 );
and \U$34885 ( \42528 , \42527 , \42517 );
or \U$34886 ( \42529 , \42519 , \42528 );
and \U$34888 ( \42530 , \42529 , 1'b1 );
or \U$34890 ( \42531 , \42530 , 1'b0 );
buf \U$34891 ( \42532 , \42531 );
_DC r23734_GF_IsGateDCbyConstraint ( \42533_nR23734 , \42532 , \21944 );
buf \U$34892 ( \42534 , \42533_nR23734 );
not \U$34893 ( \42535 , \42515 );
and \U$34894 ( \42536 , RIe136da8_5262, \42535 );
not \U$34895 ( \42537 , RIe136da8_5262);
not \U$34896 ( \42538 , \42537 );
not \U$34897 ( \42539 , \38043 );
and \U$34898 ( \42540 , \42538 , \42539 );
buf \U$34899 ( \42541 , RIb86fce0_76);
buf \U$34900 ( \42542 , \42541 );
and \U$34901 ( \42543 , \42542 , \38043 );
or \U$34902 ( \42544 , \42540 , \42543 );
and \U$34903 ( \42545 , \42544 , \42515 );
or \U$34904 ( \42546 , \42536 , \42545 );
and \U$34906 ( \42547 , \42546 , 1'b1 );
or \U$34908 ( \42548 , \42547 , 1'b0 );
buf \U$34909 ( \42549 , \42548 );
_DC r23736_GF_IsGateDCbyConstraint ( \42550_nR23736 , \42549 , \21944 );
buf \U$34910 ( \42551 , \42550_nR23736 );
not \U$34911 ( \42552 , \42517 );
and \U$34912 ( \42553 , RIe136358_5263, \42552 );
not \U$34913 ( \42554 , RIe136358_5263);
not \U$34914 ( \42555 , \42554 );
not \U$34915 ( \42556 , \38043 );
and \U$34916 ( \42557 , \42555 , \42556 );
buf \U$34917 ( \42558 , RIb86fd58_75);
buf \U$34918 ( \42559 , \42558 );
and \U$34919 ( \42560 , \42559 , \38043 );
or \U$34920 ( \42561 , \42557 , \42560 );
and \U$34921 ( \42562 , \42561 , \42517 );
or \U$34922 ( \42563 , \42553 , \42562 );
and \U$34924 ( \42564 , \42563 , 1'b1 );
or \U$34926 ( \42565 , \42564 , 1'b0 );
buf \U$34927 ( \42566 , \42565 );
_DC r23738_GF_IsGateDCbyConstraint ( \42567_nR23738 , \42566 , \21944 );
buf \U$34928 ( \42568 , \42567_nR23738 );
not \U$34929 ( \42569 , \42517 );
and \U$34930 ( \42570 , RIe135890_5264, \42569 );
not \U$34931 ( \42571 , RIe135890_5264);
not \U$34932 ( \42572 , \42571 );
not \U$34933 ( \42573 , \38043 );
and \U$34934 ( \42574 , \42572 , \42573 );
buf \U$34935 ( \42575 , RIb87e8a8_74);
buf \U$34936 ( \42576 , \42575 );
and \U$34937 ( \42577 , \42576 , \38043 );
or \U$34938 ( \42578 , \42574 , \42577 );
and \U$34939 ( \42579 , \42578 , \42517 );
or \U$34940 ( \42580 , \42570 , \42579 );
and \U$34942 ( \42581 , \42580 , 1'b1 );
or \U$34944 ( \42582 , \42581 , 1'b0 );
buf \U$34945 ( \42583 , \42582 );
_DC r2373a_GF_IsGateDCbyConstraint ( \42584_nR2373a , \42583 , \21944 );
buf \U$34946 ( \42585 , \42584_nR2373a );
not \U$34947 ( \42586 , \42517 );
and \U$34948 ( \42587 , RIe134d50_5265, \42586 );
not \U$34949 ( \42588 , RIe134d50_5265);
not \U$34950 ( \42589 , \42588 );
not \U$34951 ( \42590 , \38043 );
and \U$34952 ( \42591 , \42589 , \42590 );
buf \U$34953 ( \42592 , RIb87e920_73);
buf \U$34954 ( \42593 , \42592 );
and \U$34955 ( \42594 , \42593 , \38043 );
or \U$34956 ( \42595 , \42591 , \42594 );
and \U$34957 ( \42596 , \42595 , \42517 );
or \U$34958 ( \42597 , \42587 , \42596 );
and \U$34960 ( \42598 , \42597 , 1'b1 );
or \U$34962 ( \42599 , \42598 , 1'b0 );
buf \U$34963 ( \42600 , \42599 );
_DC r2373c_GF_IsGateDCbyConstraint ( \42601_nR2373c , \42600 , \21944 );
buf \U$34964 ( \42602 , \42601_nR2373c );
not \U$34965 ( \42603 , \42515 );
and \U$34966 ( \42604 , RIe134288_5266, \42603 );
not \U$34967 ( \42605 , RIe134288_5266);
not \U$34968 ( \42606 , \42605 );
not \U$34969 ( \42607 , \38043 );
and \U$34970 ( \42608 , \42606 , \42607 );
buf \U$34971 ( \42609 , RIb87e998_72);
buf \U$34972 ( \42610 , \42609 );
and \U$34973 ( \42611 , \42610 , \38043 );
or \U$34974 ( \42612 , \42608 , \42611 );
and \U$34975 ( \42613 , \42612 , \42515 );
or \U$34976 ( \42614 , \42604 , \42613 );
and \U$34978 ( \42615 , \42614 , 1'b1 );
or \U$34980 ( \42616 , \42615 , 1'b0 );
buf \U$34981 ( \42617 , \42616 );
_DC r2373e_GF_IsGateDCbyConstraint ( \42618_nR2373e , \42617 , \21944 );
buf \U$34982 ( \42619 , \42618_nR2373e );
not \U$34983 ( \42620 , \42517 );
and \U$34984 ( \42621 , RIe1337c0_5267, \42620 );
not \U$34985 ( \42622 , RIe1337c0_5267);
not \U$34986 ( \42623 , \42622 );
not \U$34987 ( \42624 , \38043 );
and \U$34988 ( \42625 , \42623 , \42624 );
buf \U$34989 ( \42626 , RIb87ea10_71);
buf \U$34990 ( \42627 , \42626 );
and \U$34991 ( \42628 , \42627 , \38043 );
or \U$34992 ( \42629 , \42625 , \42628 );
and \U$34993 ( \42630 , \42629 , \42517 );
or \U$34994 ( \42631 , \42621 , \42630 );
and \U$34996 ( \42632 , \42631 , 1'b1 );
or \U$34998 ( \42633 , \42632 , 1'b0 );
buf \U$34999 ( \42634 , \42633 );
_DC r23740_GF_IsGateDCbyConstraint ( \42635_nR23740 , \42634 , \21944 );
buf \U$35000 ( \42636 , \42635_nR23740 );
not \U$35001 ( \42637 , \42515 );
and \U$35002 ( \42638 , RIe132c08_5268, \42637 );
not \U$35003 ( \42639 , RIe132c08_5268);
not \U$35004 ( \42640 , \42639 );
not \U$35005 ( \42641 , \38043 );
and \U$35006 ( \42642 , \42640 , \42641 );
buf \U$35007 ( \42643 , RIb87ea88_70);
buf \U$35008 ( \42644 , \42643 );
and \U$35009 ( \42645 , \42644 , \38043 );
or \U$35010 ( \42646 , \42642 , \42645 );
and \U$35011 ( \42647 , \42646 , \42515 );
or \U$35012 ( \42648 , \42638 , \42647 );
and \U$35014 ( \42649 , \42648 , 1'b1 );
or \U$35016 ( \42650 , \42649 , 1'b0 );
buf \U$35017 ( \42651 , \42650 );
_DC r23742_GF_IsGateDCbyConstraint ( \42652_nR23742 , \42651 , \21944 );
buf \U$35018 ( \42653 , \42652_nR23742 );
not \U$35019 ( \42654 , \42517 );
and \U$35020 ( \42655 , RIe131fd8_5269, \42654 );
not \U$35021 ( \42656 , RIe131fd8_5269);
not \U$35022 ( \42657 , \42656 );
not \U$35023 ( \42658 , \39308 );
and \U$35024 ( \42659 , \42657 , \42658 );
and \U$35025 ( \42660 , \42525 , \39308 );
or \U$35026 ( \42661 , \42659 , \42660 );
and \U$35027 ( \42662 , \42661 , \42517 );
or \U$35028 ( \42663 , \42655 , \42662 );
and \U$35030 ( \42664 , \42663 , 1'b1 );
or \U$35032 ( \42665 , \42664 , 1'b0 );
buf \U$35033 ( \42666 , \42665 );
_DC r23744_GF_IsGateDCbyConstraint ( \42667_nR23744 , \42666 , \21944 );
buf \U$35034 ( \42668 , \42667_nR23744 );
not \U$35035 ( \42669 , \42515 );
and \U$35036 ( \42670 , RIe1313a8_5270, \42669 );
not \U$35037 ( \42671 , RIe1313a8_5270);
not \U$35038 ( \42672 , \42671 );
not \U$35039 ( \42673 , \39308 );
and \U$35040 ( \42674 , \42672 , \42673 );
and \U$35041 ( \42675 , \42542 , \39308 );
or \U$35042 ( \42676 , \42674 , \42675 );
and \U$35043 ( \42677 , \42676 , \42515 );
or \U$35044 ( \42678 , \42670 , \42677 );
and \U$35046 ( \42679 , \42678 , 1'b1 );
or \U$35048 ( \42680 , \42679 , 1'b0 );
buf \U$35049 ( \42681 , \42680 );
_DC r23746_GF_IsGateDCbyConstraint ( \42682_nR23746 , \42681 , \21944 );
buf \U$35050 ( \42683 , \42682_nR23746 );
not \U$35051 ( \42684 , \42517 );
and \U$35052 ( \42685 , RIe1307f0_5271, \42684 );
not \U$35053 ( \42686 , RIe1307f0_5271);
not \U$35054 ( \42687 , \42686 );
not \U$35055 ( \42688 , \39308 );
and \U$35056 ( \42689 , \42687 , \42688 );
and \U$35057 ( \42690 , \42559 , \39308 );
or \U$35058 ( \42691 , \42689 , \42690 );
and \U$35059 ( \42692 , \42691 , \42517 );
or \U$35060 ( \42693 , \42685 , \42692 );
and \U$35062 ( \42694 , \42693 , 1'b1 );
or \U$35064 ( \42695 , \42694 , 1'b0 );
buf \U$35065 ( \42696 , \42695 );
_DC r23748_GF_IsGateDCbyConstraint ( \42697_nR23748 , \42696 , \21944 );
buf \U$35066 ( \42698 , \42697_nR23748 );
not \U$35067 ( \42699 , \42515 );
and \U$35068 ( \42700 , RIe12fbc0_5272, \42699 );
not \U$35069 ( \42701 , RIe12fbc0_5272);
not \U$35070 ( \42702 , \42701 );
not \U$35071 ( \42703 , \39308 );
and \U$35072 ( \42704 , \42702 , \42703 );
and \U$35073 ( \42705 , \42576 , \39308 );
or \U$35074 ( \42706 , \42704 , \42705 );
and \U$35075 ( \42707 , \42706 , \42515 );
or \U$35076 ( \42708 , \42700 , \42707 );
and \U$35078 ( \42709 , \42708 , 1'b1 );
or \U$35080 ( \42710 , \42709 , 1'b0 );
buf \U$35081 ( \42711 , \42710 );
_DC r2374a_GF_IsGateDCbyConstraint ( \42712_nR2374a , \42711 , \21944 );
buf \U$35082 ( \42713 , \42712_nR2374a );
not \U$35083 ( \42714 , \42517 );
and \U$35084 ( \42715 , RIe12f080_5273, \42714 );
not \U$35085 ( \42716 , RIe12f080_5273);
not \U$35086 ( \42717 , \42716 );
not \U$35087 ( \42718 , \39308 );
and \U$35088 ( \42719 , \42717 , \42718 );
and \U$35089 ( \42720 , \42593 , \39308 );
or \U$35090 ( \42721 , \42719 , \42720 );
and \U$35091 ( \42722 , \42721 , \42517 );
or \U$35092 ( \42723 , \42715 , \42722 );
and \U$35094 ( \42724 , \42723 , 1'b1 );
or \U$35096 ( \42725 , \42724 , 1'b0 );
buf \U$35097 ( \42726 , \42725 );
_DC r2374c_GF_IsGateDCbyConstraint ( \42727_nR2374c , \42726 , \21944 );
buf \U$35098 ( \42728 , \42727_nR2374c );
not \U$35099 ( \42729 , \42515 );
and \U$35100 ( \42730 , RIe12da78_5274, \42729 );
not \U$35101 ( \42731 , RIe12da78_5274);
not \U$35102 ( \42732 , \42731 );
not \U$35103 ( \42733 , \39308 );
and \U$35104 ( \42734 , \42732 , \42733 );
and \U$35105 ( \42735 , \42610 , \39308 );
or \U$35106 ( \42736 , \42734 , \42735 );
and \U$35107 ( \42737 , \42736 , \42515 );
or \U$35108 ( \42738 , \42730 , \42737 );
and \U$35110 ( \42739 , \42738 , 1'b1 );
or \U$35112 ( \42740 , \42739 , 1'b0 );
buf \U$35113 ( \42741 , \42740 );
_DC r2374e_GF_IsGateDCbyConstraint ( \42742_nR2374e , \42741 , \21944 );
buf \U$35114 ( \42743 , \42742_nR2374e );
not \U$35115 ( \42744 , \42517 );
and \U$35116 ( \42745 , RIe12c920_5275, \42744 );
not \U$35117 ( \42746 , RIe12c920_5275);
not \U$35118 ( \42747 , \42746 );
not \U$35119 ( \42748 , \39308 );
and \U$35120 ( \42749 , \42747 , \42748 );
and \U$35121 ( \42750 , \42627 , \39308 );
or \U$35122 ( \42751 , \42749 , \42750 );
and \U$35123 ( \42752 , \42751 , \42517 );
or \U$35124 ( \42753 , \42745 , \42752 );
and \U$35126 ( \42754 , \42753 , 1'b1 );
or \U$35128 ( \42755 , \42754 , 1'b0 );
buf \U$35129 ( \42756 , \42755 );
_DC r23750_GF_IsGateDCbyConstraint ( \42757_nR23750 , \42756 , \21944 );
buf \U$35130 ( \42758 , \42757_nR23750 );
not \U$35131 ( \42759 , \42515 );
and \U$35132 ( \42760 , RIe12b318_5276, \42759 );
not \U$35133 ( \42761 , RIe12b318_5276);
not \U$35134 ( \42762 , \42761 );
not \U$35135 ( \42763 , \39308 );
and \U$35136 ( \42764 , \42762 , \42763 );
and \U$35137 ( \42765 , \42644 , \39308 );
or \U$35138 ( \42766 , \42764 , \42765 );
and \U$35139 ( \42767 , \42766 , \42515 );
or \U$35140 ( \42768 , \42760 , \42767 );
and \U$35142 ( \42769 , \42768 , 1'b1 );
or \U$35144 ( \42770 , \42769 , 1'b0 );
buf \U$35145 ( \42771 , \42770 );
_DC r23752_GF_IsGateDCbyConstraint ( \42772_nR23752 , \42771 , \21944 );
buf \U$35146 ( \42773 , \42772_nR23752 );
not \U$35147 ( \42774 , \42517 );
and \U$35148 ( \42775 , RIe12a1c0_5277, \42774 );
not \U$35149 ( \42776 , RIe12a1c0_5277);
not \U$35150 ( \42777 , \42776 );
not \U$35151 ( \42778 , \40486 );
and \U$35152 ( \42779 , \42777 , \42778 );
and \U$35153 ( \42780 , \42525 , \40486 );
or \U$35154 ( \42781 , \42779 , \42780 );
and \U$35155 ( \42782 , \42781 , \42517 );
or \U$35156 ( \42783 , \42775 , \42782 );
and \U$35158 ( \42784 , \42783 , 1'b1 );
or \U$35160 ( \42785 , \42784 , 1'b0 );
buf \U$35161 ( \42786 , \42785 );
_DC r23754_GF_IsGateDCbyConstraint ( \42787_nR23754 , \42786 , \21944 );
buf \U$35162 ( \42788 , \42787_nR23754 );
not \U$35163 ( \42789 , \42517 );
and \U$35164 ( \42790 , RIe128bb8_5278, \42789 );
not \U$35165 ( \42791 , RIe128bb8_5278);
not \U$35166 ( \42792 , \42791 );
not \U$35167 ( \42793 , \40486 );
and \U$35168 ( \42794 , \42792 , \42793 );
and \U$35169 ( \42795 , \42542 , \40486 );
or \U$35170 ( \42796 , \42794 , \42795 );
and \U$35171 ( \42797 , \42796 , \42517 );
or \U$35172 ( \42798 , \42790 , \42797 );
and \U$35174 ( \42799 , \42798 , 1'b1 );
or \U$35176 ( \42800 , \42799 , 1'b0 );
buf \U$35177 ( \42801 , \42800 );
_DC r23756_GF_IsGateDCbyConstraint ( \42802_nR23756 , \42801 , \21944 );
buf \U$35178 ( \42803 , \42802_nR23756 );
not \U$35179 ( \42804 , \42517 );
and \U$35180 ( \42805 , RIe127a60_5279, \42804 );
not \U$35181 ( \42806 , RIe127a60_5279);
not \U$35182 ( \42807 , \42806 );
not \U$35183 ( \42808 , \40486 );
and \U$35184 ( \42809 , \42807 , \42808 );
and \U$35185 ( \42810 , \42559 , \40486 );
or \U$35186 ( \42811 , \42809 , \42810 );
and \U$35187 ( \42812 , \42811 , \42517 );
or \U$35188 ( \42813 , \42805 , \42812 );
and \U$35190 ( \42814 , \42813 , 1'b1 );
or \U$35192 ( \42815 , \42814 , 1'b0 );
buf \U$35193 ( \42816 , \42815 );
_DC r23758_GF_IsGateDCbyConstraint ( \42817_nR23758 , \42816 , \21944 );
buf \U$35194 ( \42818 , \42817_nR23758 );
not \U$35195 ( \42819 , \42517 );
and \U$35196 ( \42820 , RIe126908_5280, \42819 );
not \U$35197 ( \42821 , RIe126908_5280);
not \U$35198 ( \42822 , \42821 );
not \U$35199 ( \42823 , \40486 );
and \U$35200 ( \42824 , \42822 , \42823 );
and \U$35201 ( \42825 , \42576 , \40486 );
or \U$35202 ( \42826 , \42824 , \42825 );
and \U$35203 ( \42827 , \42826 , \42517 );
or \U$35204 ( \42828 , \42820 , \42827 );
and \U$35206 ( \42829 , \42828 , 1'b1 );
or \U$35208 ( \42830 , \42829 , 1'b0 );
buf \U$35209 ( \42831 , \42830 );
_DC r2375a_GF_IsGateDCbyConstraint ( \42832_nR2375a , \42831 , \21944 );
buf \U$35210 ( \42833 , \42832_nR2375a );
not \U$35211 ( \42834 , \42517 );
and \U$35212 ( \42835 , RIe125300_5281, \42834 );
not \U$35213 ( \42836 , RIe125300_5281);
not \U$35214 ( \42837 , \42836 );
not \U$35215 ( \42838 , \40486 );
and \U$35216 ( \42839 , \42837 , \42838 );
and \U$35217 ( \42840 , \42593 , \40486 );
or \U$35218 ( \42841 , \42839 , \42840 );
and \U$35219 ( \42842 , \42841 , \42517 );
or \U$35220 ( \42843 , \42835 , \42842 );
and \U$35222 ( \42844 , \42843 , 1'b1 );
or \U$35224 ( \42845 , \42844 , 1'b0 );
buf \U$35225 ( \42846 , \42845 );
_DC r2375c_GF_IsGateDCbyConstraint ( \42847_nR2375c , \42846 , \21944 );
buf \U$35226 ( \42848 , \42847_nR2375c );
not \U$35227 ( \42849 , \42517 );
and \U$35228 ( \42850 , RIe1241a8_5282, \42849 );
not \U$35229 ( \42851 , RIe1241a8_5282);
not \U$35230 ( \42852 , \42851 );
not \U$35231 ( \42853 , \40486 );
and \U$35232 ( \42854 , \42852 , \42853 );
and \U$35233 ( \42855 , \42610 , \40486 );
or \U$35234 ( \42856 , \42854 , \42855 );
and \U$35235 ( \42857 , \42856 , \42517 );
or \U$35236 ( \42858 , \42850 , \42857 );
and \U$35238 ( \42859 , \42858 , 1'b1 );
or \U$35240 ( \42860 , \42859 , 1'b0 );
buf \U$35241 ( \42861 , \42860 );
_DC r2375e_GF_IsGateDCbyConstraint ( \42862_nR2375e , \42861 , \21944 );
buf \U$35242 ( \42863 , \42862_nR2375e );
not \U$35243 ( \42864 , \42517 );
and \U$35244 ( \42865 , RIe122ba0_5283, \42864 );
not \U$35245 ( \42866 , RIe122ba0_5283);
not \U$35246 ( \42867 , \42866 );
not \U$35247 ( \42868 , \40486 );
and \U$35248 ( \42869 , \42867 , \42868 );
and \U$35249 ( \42870 , \42627 , \40486 );
or \U$35250 ( \42871 , \42869 , \42870 );
and \U$35251 ( \42872 , \42871 , \42517 );
or \U$35252 ( \42873 , \42865 , \42872 );
and \U$35254 ( \42874 , \42873 , 1'b1 );
or \U$35256 ( \42875 , \42874 , 1'b0 );
buf \U$35257 ( \42876 , \42875 );
_DC r23760_GF_IsGateDCbyConstraint ( \42877_nR23760 , \42876 , \21944 );
buf \U$35258 ( \42878 , \42877_nR23760 );
not \U$35259 ( \42879 , \42517 );
and \U$35260 ( \42880 , RIe121a48_5284, \42879 );
not \U$35261 ( \42881 , RIe121a48_5284);
not \U$35262 ( \42882 , \42881 );
not \U$35263 ( \42883 , \40486 );
and \U$35264 ( \42884 , \42882 , \42883 );
and \U$35265 ( \42885 , \42644 , \40486 );
or \U$35266 ( \42886 , \42884 , \42885 );
and \U$35267 ( \42887 , \42886 , \42517 );
or \U$35268 ( \42888 , \42880 , \42887 );
and \U$35270 ( \42889 , \42888 , 1'b1 );
or \U$35272 ( \42890 , \42889 , 1'b0 );
buf \U$35273 ( \42891 , \42890 );
_DC r23762_GF_IsGateDCbyConstraint ( \42892_nR23762 , \42891 , \21944 );
buf \U$35274 ( \42893 , \42892_nR23762 );
not \U$35275 ( \42894 , \42517 );
and \U$35276 ( \42895 , RIe120440_5285, \42894 );
not \U$35277 ( \42896 , RIe120440_5285);
not \U$35278 ( \42897 , \42896 );
not \U$35279 ( \42898 , \41604 );
and \U$35280 ( \42899 , \42897 , \42898 );
and \U$35281 ( \42900 , \42525 , \41604 );
or \U$35282 ( \42901 , \42899 , \42900 );
and \U$35283 ( \42902 , \42901 , \42517 );
or \U$35284 ( \42903 , \42895 , \42902 );
and \U$35286 ( \42904 , \42903 , 1'b1 );
or \U$35288 ( \42905 , \42904 , 1'b0 );
buf \U$35289 ( \42906 , \42905 );
_DC r23764_GF_IsGateDCbyConstraint ( \42907_nR23764 , \42906 , \21944 );
buf \U$35290 ( \42908 , \42907_nR23764 );
not \U$35291 ( \42909 , \42515 );
and \U$35292 ( \42910 , RIe11f2e8_5286, \42909 );
not \U$35293 ( \42911 , RIe11f2e8_5286);
not \U$35294 ( \42912 , \42911 );
not \U$35295 ( \42913 , \41604 );
and \U$35296 ( \42914 , \42912 , \42913 );
and \U$35297 ( \42915 , \42542 , \41604 );
or \U$35298 ( \42916 , \42914 , \42915 );
and \U$35299 ( \42917 , \42916 , \42515 );
or \U$35300 ( \42918 , \42910 , \42917 );
and \U$35302 ( \42919 , \42918 , 1'b1 );
or \U$35304 ( \42920 , \42919 , 1'b0 );
buf \U$35305 ( \42921 , \42920 );
_DC r23766_GF_IsGateDCbyConstraint ( \42922_nR23766 , \42921 , \21944 );
buf \U$35306 ( \42923 , \42922_nR23766 );
not \U$35307 ( \42924 , \42515 );
and \U$35308 ( \42925 , RIe11e190_5287, \42924 );
not \U$35309 ( \42926 , RIe11e190_5287);
not \U$35310 ( \42927 , \42926 );
not \U$35311 ( \42928 , \41604 );
and \U$35312 ( \42929 , \42927 , \42928 );
and \U$35313 ( \42930 , \42559 , \41604 );
or \U$35314 ( \42931 , \42929 , \42930 );
and \U$35315 ( \42932 , \42931 , \42515 );
or \U$35316 ( \42933 , \42925 , \42932 );
and \U$35318 ( \42934 , \42933 , 1'b1 );
or \U$35320 ( \42935 , \42934 , 1'b0 );
buf \U$35321 ( \42936 , \42935 );
_DC r23768_GF_IsGateDCbyConstraint ( \42937_nR23768 , \42936 , \21944 );
buf \U$35322 ( \42938 , \42937_nR23768 );
not \U$35323 ( \42939 , \42515 );
and \U$35324 ( \42940 , RIe11cb88_5288, \42939 );
not \U$35325 ( \42941 , RIe11cb88_5288);
not \U$35326 ( \42942 , \42941 );
not \U$35327 ( \42943 , \41604 );
and \U$35328 ( \42944 , \42942 , \42943 );
and \U$35329 ( \42945 , \42576 , \41604 );
or \U$35330 ( \42946 , \42944 , \42945 );
and \U$35331 ( \42947 , \42946 , \42515 );
or \U$35332 ( \42948 , \42940 , \42947 );
and \U$35334 ( \42949 , \42948 , 1'b1 );
or \U$35336 ( \42950 , \42949 , 1'b0 );
buf \U$35337 ( \42951 , \42950 );
_DC r2376a_GF_IsGateDCbyConstraint ( \42952_nR2376a , \42951 , \21944 );
buf \U$35338 ( \42953 , \42952_nR2376a );
not \U$35339 ( \42954 , \42515 );
and \U$35340 ( \42955 , RIe11ba30_5289, \42954 );
not \U$35341 ( \42956 , RIe11ba30_5289);
not \U$35342 ( \42957 , \42956 );
not \U$35343 ( \42958 , \41604 );
and \U$35344 ( \42959 , \42957 , \42958 );
and \U$35345 ( \42960 , \42593 , \41604 );
or \U$35346 ( \42961 , \42959 , \42960 );
and \U$35347 ( \42962 , \42961 , \42515 );
or \U$35348 ( \42963 , \42955 , \42962 );
and \U$35350 ( \42964 , \42963 , 1'b1 );
or \U$35352 ( \42965 , \42964 , 1'b0 );
buf \U$35353 ( \42966 , \42965 );
_DC r2376c_GF_IsGateDCbyConstraint ( \42967_nR2376c , \42966 , \21944 );
buf \U$35354 ( \42968 , \42967_nR2376c );
not \U$35355 ( \42969 , \42515 );
and \U$35356 ( \42970 , RIe11a428_5290, \42969 );
not \U$35357 ( \42971 , RIe11a428_5290);
not \U$35358 ( \42972 , \42971 );
not \U$35359 ( \42973 , \41604 );
and \U$35360 ( \42974 , \42972 , \42973 );
and \U$35361 ( \42975 , \42610 , \41604 );
or \U$35362 ( \42976 , \42974 , \42975 );
and \U$35363 ( \42977 , \42976 , \42515 );
or \U$35364 ( \42978 , \42970 , \42977 );
and \U$35366 ( \42979 , \42978 , 1'b1 );
or \U$35368 ( \42980 , \42979 , 1'b0 );
buf \U$35369 ( \42981 , \42980 );
_DC r2376e_GF_IsGateDCbyConstraint ( \42982_nR2376e , \42981 , \21944 );
buf \U$35370 ( \42983 , \42982_nR2376e );
not \U$35371 ( \42984 , \42515 );
and \U$35372 ( \42985 , RIe1192d0_5291, \42984 );
not \U$35373 ( \42986 , RIe1192d0_5291);
not \U$35374 ( \42987 , \42986 );
not \U$35375 ( \42988 , \41604 );
and \U$35376 ( \42989 , \42987 , \42988 );
and \U$35377 ( \42990 , \42627 , \41604 );
or \U$35378 ( \42991 , \42989 , \42990 );
and \U$35379 ( \42992 , \42991 , \42515 );
or \U$35380 ( \42993 , \42985 , \42992 );
and \U$35382 ( \42994 , \42993 , 1'b1 );
or \U$35384 ( \42995 , \42994 , 1'b0 );
buf \U$35385 ( \42996 , \42995 );
_DC r23770_GF_IsGateDCbyConstraint ( \42997_nR23770 , \42996 , \21944 );
buf \U$35386 ( \42998 , \42997_nR23770 );
not \U$35387 ( \42999 , \42517 );
and \U$35388 ( \43000 , RIe117cc8_5292, \42999 );
not \U$35389 ( \43001 , RIe117cc8_5292);
not \U$35390 ( \43002 , \43001 );
not \U$35391 ( \43003 , \41604 );
and \U$35392 ( \43004 , \43002 , \43003 );
and \U$35393 ( \43005 , \42644 , \41604 );
or \U$35394 ( \43006 , \43004 , \43005 );
and \U$35395 ( \43007 , \43006 , \42517 );
or \U$35396 ( \43008 , \43000 , \43007 );
and \U$35398 ( \43009 , \43008 , 1'b1 );
or \U$35400 ( \43010 , \43009 , 1'b0 );
buf \U$35401 ( \43011 , \43010 );
_DC r23772_GF_IsGateDCbyConstraint ( \43012_nR23772 , \43011 , \21944 );
buf \U$35402 ( \43013 , \43012_nR23772 );
buf \U$35403 ( \43014 , \21699 );
not \U$35404 ( \43015 , \43014 );
buf \U$35405 ( \43016 , RIb79b3b0_273);
nand \U$35406 ( \43017 , \43016 , \38028 );
not \U$35407 ( \43018 , \43017 );
and \U$35408 ( \43019 , \43015 , \43018 );
not \U$35409 ( \43020 , RIe38a110_5575);
and \U$35410 ( \43021 , \43020 , \43017 );
or \U$35411 ( \43022 , \43019 , \43021 );
not \U$35412 ( \43023 , \43022 );
and \U$35414 ( \43024 , \43023 , 1'b1 );
or \U$35416 ( \43025 , \43024 , 1'b0 );
buf \U$35417 ( \43026 , \43025 );
_DC r2398c_GF_IsGateDCbyConstraint ( \43027_nR2398c , \43026 , \21944 );
buf \U$35418 ( \43028 , \43027_nR2398c );
not \U$35419 ( \43029 , \43017 );
not \U$35420 ( \43030 , \43029 );
and \U$35421 ( \43031 , RIe378410_5590, \43030 );
buf \U$35422 ( \43032 , RIb7b96f8_244);
and \U$35423 ( \43033 , \43032 , \43029 );
or \U$35424 ( \43034 , \43031 , \43033 );
and \U$35426 ( \43035 , \43034 , 1'b1 );
or \U$35428 ( \43036 , \43035 , 1'b0 );
buf \U$35429 ( \43037 , \43036 );
_DC r2398e_GF_IsGateDCbyConstraint ( \43038_nR2398e , \43037 , \21944 );
buf \U$35430 ( \43039 , \43038_nR2398e );
not \U$35431 ( \43040 , \43029 );
and \U$35432 ( \43041 , RIe379220_5589, \43040 );
buf \U$35433 ( \43042 , RIb7c20c8_243);
and \U$35434 ( \43043 , \43042 , \43029 );
or \U$35435 ( \43044 , \43041 , \43043 );
and \U$35437 ( \43045 , \43044 , 1'b1 );
or \U$35439 ( \43046 , \43045 , 1'b0 );
buf \U$35440 ( \43047 , \43046 );
_DC r23990_GF_IsGateDCbyConstraint ( \43048_nR23990 , \43047 , \21944 );
buf \U$35441 ( \43049 , \43048_nR23990 );
not \U$35442 ( \43050 , \43029 );
and \U$35443 ( \43051 , RIe379e50_5588, \43050 );
buf \U$35444 ( \43052 , RIb7c5728_242);
and \U$35445 ( \43053 , \43052 , \43029 );
or \U$35446 ( \43054 , \43051 , \43053 );
and \U$35448 ( \43055 , \43054 , 1'b1 );
or \U$35450 ( \43056 , \43055 , 1'b0 );
buf \U$35451 ( \43057 , \43056 );
_DC r23992_GF_IsGateDCbyConstraint ( \43058_nR23992 , \43057 , \21944 );
buf \U$35452 ( \43059 , \43058_nR23992 );
not \U$35453 ( \43060 , \43029 );
and \U$35454 ( \43061 , RIe26f4f8_5601, \43060 );
buf \U$35455 ( \43062 , RIb7c57a0_241);
and \U$35456 ( \43063 , \43062 , \43029 );
or \U$35457 ( \43064 , \43061 , \43063 );
and \U$35459 ( \43065 , \43064 , 1'b1 );
or \U$35461 ( \43066 , \43065 , 1'b0 );
buf \U$35462 ( \43067 , \43066 );
_DC r23994_GF_IsGateDCbyConstraint ( \43068_nR23994 , \43067 , \21944 );
buf \U$35463 ( \43069 , \43068_nR23994 );
not \U$35464 ( \43070 , \43029 );
and \U$35465 ( \43071 , RIe270290_5600, \43070 );
buf \U$35466 ( \43072 , RIb7c5818_240);
and \U$35467 ( \43073 , \43072 , \43029 );
or \U$35468 ( \43074 , \43071 , \43073 );
and \U$35470 ( \43075 , \43074 , 1'b1 );
or \U$35472 ( \43076 , \43075 , 1'b0 );
buf \U$35473 ( \43077 , \43076 );
_DC r23996_GF_IsGateDCbyConstraint ( \43078_nR23996 , \43077 , \21944 );
buf \U$35474 ( \43079 , \43078_nR23996 );
not \U$35475 ( \43080 , \43029 );
and \U$35476 ( \43081 , RIe270ec0_5599, \43080 );
buf \U$35477 ( \43082 , RIb7c5890_239);
and \U$35478 ( \43083 , \43082 , \43029 );
or \U$35479 ( \43084 , \43081 , \43083 );
and \U$35481 ( \43085 , \43084 , 1'b1 );
or \U$35483 ( \43086 , \43085 , 1'b0 );
buf \U$35484 ( \43087 , \43086 );
_DC r23998_GF_IsGateDCbyConstraint ( \43088_nR23998 , \43087 , \21944 );
buf \U$35485 ( \43089 , \43088_nR23998 );
not \U$35486 ( \43090 , \43029 );
and \U$35487 ( \43091 , RIe271be0_5598, \43090 );
buf \U$35488 ( \43092 , RIb7c5908_238);
and \U$35489 ( \43093 , \43092 , \43029 );
or \U$35490 ( \43094 , \43091 , \43093 );
and \U$35492 ( \43095 , \43094 , 1'b1 );
or \U$35494 ( \43096 , \43095 , 1'b0 );
buf \U$35495 ( \43097 , \43096 );
_DC r2399a_GF_IsGateDCbyConstraint ( \43098_nR2399a , \43097 , \21944 );
buf \U$35496 ( \43099 , \43098_nR2399a );
not \U$35497 ( \43100 , \43029 );
and \U$35498 ( \43101 , RIe37b908_5586, \43100 );
buf \U$35499 ( \43102 , RIb7a09f0_266);
and \U$35500 ( \43103 , \43102 , \43029 );
or \U$35501 ( \43104 , \43101 , \43103 );
and \U$35503 ( \43105 , \43104 , 1'b1 );
or \U$35505 ( \43106 , \43105 , 1'b0 );
buf \U$35506 ( \43107 , \43106 );
_DC r2398a_GF_IsGateDCbyConstraint ( \43108_nR2398a , \43107 , \21944 );
buf \U$35507 ( \43109 , \43108_nR2398a );
not \U$35508 ( \43110 , \43029 );
and \U$35509 ( \43111 , RIe375008_5594, \43110 );
buf \U$35510 ( \43112 , RIb7a0a68_265);
and \U$35511 ( \43113 , \43112 , \43029 );
or \U$35512 ( \43114 , \43111 , \43113 );
and \U$35514 ( \43115 , \43114 , 1'b1 );
or \U$35516 ( \43116 , \43115 , 1'b0 );
buf \U$35517 ( \43117 , \43116 );
_DC r2399c_GF_IsGateDCbyConstraint ( \43118_nR2399c , \43117 , \21944 );
buf \U$35518 ( \43119 , \43118_nR2399c );
not \U$35519 ( \43120 , \43029 );
and \U$35520 ( \43121 , RIe375da0_5593, \43120 );
buf \U$35521 ( \43122 , RIb7a0ae0_264);
and \U$35522 ( \43123 , \43122 , \43029 );
or \U$35523 ( \43124 , \43121 , \43123 );
and \U$35525 ( \43125 , \43124 , 1'b1 );
or \U$35527 ( \43126 , \43125 , 1'b0 );
buf \U$35528 ( \43127 , \43126 );
_DC r2399e_GF_IsGateDCbyConstraint ( \43128_nR2399e , \43127 , \21944 );
buf \U$35529 ( \43129 , \43128_nR2399e );
not \U$35530 ( \43130 , \43029 );
and \U$35531 ( \43131 , RIe376a48_5592, \43130 );
buf \U$35532 ( \43132 , RIb7a0b58_263);
and \U$35533 ( \43133 , \43132 , \43029 );
or \U$35534 ( \43134 , \43131 , \43133 );
and \U$35536 ( \43135 , \43134 , 1'b1 );
or \U$35538 ( \43136 , \43135 , 1'b0 );
buf \U$35539 ( \43137 , \43136 );
_DC r239a0_GF_IsGateDCbyConstraint ( \43138_nR239a0 , \43137 , \21944 );
buf \U$35540 ( \43139 , \43138_nR239a0 );
not \U$35541 ( \43140 , \43029 );
and \U$35542 ( \43141 , RIe377768_5591, \43140 );
buf \U$35543 ( \43142 , RIb7a0bd0_262);
and \U$35544 ( \43143 , \43142 , \43029 );
or \U$35545 ( \43144 , \43141 , \43143 );
and \U$35547 ( \43145 , \43144 , 1'b1 );
or \U$35549 ( \43146 , \43145 , 1'b0 );
buf \U$35550 ( \43147 , \43146 );
_DC r239a2_GF_IsGateDCbyConstraint ( \43148_nR239a2 , \43147 , \21944 );
buf \U$35551 ( \43149 , \43148_nR239a2 );
not \U$35552 ( \43150 , RIe3921f8_5562);
not \U$35553 ( \43151 , \43150 );
or \U$35554 ( \43152 , RIe392b58_5561, \43151 );
not \U$35555 ( \43153 , \43152 );
and \U$35556 ( \43154 , \43153 , RIe3934b8_5560);
nand \U$35557 ( \43155 , \38024 , \38028 );
not \U$35558 ( \43156 , \43155 );
not \U$35559 ( \43157 , RIe37f9b8_5584);
or \U$35560 ( \43158 , \43014 , \43157 );
nand \U$35561 ( \43159 , \43158 , \38024 , \38028 );
buf \U$35562 ( \43160 , RIb79b4a0_271);
not \U$35563 ( \43161 , \9810 );
and \U$35564 ( \43162 , \43161 , \13923 );
buf \U$35565 ( \43163 , \43162 );
nand \U$35566 ( \43164 , \43160 , \43163 );
not \U$35567 ( \43165 , \43164 );
buf \U$35568 ( \43166 , RIb79b338_274);
buf \U$35569 ( \43167 , \43166 );
nand \U$35570 ( \43168 , \43163 , \43167 );
not \U$35571 ( \43169 , \43168 );
nor \U$35572 ( \43170 , \43165 , \43169 );
nand \U$35573 ( \43171 , \43156 , \43159 , \43170 );
or \U$35574 ( \43172 , \43154 , \43171 );
nand \U$35575 ( \43173 , \38024 , \38028 );
not \U$35576 ( \43174 , \43173 );
not \U$35577 ( \43175 , \43174 );
and \U$35578 ( \43176 , \43168 , \43165 );
not \U$35579 ( \43177 , \43152 );
not \U$35580 ( \43178 , \43177 );
or \U$35581 ( \43179 , RIe3934b8_5560, \43178 );
nand \U$35582 ( \43180 , \43175 , \43176 , \43179 );
nand \U$35583 ( \43181 , \43172 , \43180 );
not \U$35584 ( \43182 , \43181 );
or \U$35585 ( \43183 , \43174 , \43177 );
not \U$35586 ( \43184 , \43150 );
nand \U$35587 ( \43185 , RIe392b58_5561, \43184 );
nand \U$35588 ( \43186 , \43183 , \43185 );
xnor \U$35589 ( \43187 , \43186 , \43173 );
nor \U$35590 ( \43188 , \43182 , \43187 );
not \U$35591 ( \43189 , \43188 );
not \U$35592 ( \43190 , RIe3934b8_5560);
and \U$35593 ( \43191 , \43189 , \43190 );
not \U$35594 ( \43192 , \43169 );
not \U$35595 ( \43193 , \43159 );
not \U$35596 ( \43194 , \43193 );
xnor \U$35597 ( \43195 , \43165 , \43174 );
and \U$35598 ( \43196 , \43192 , \43194 , \43195 );
not \U$35599 ( \43197 , \43196 );
not \U$35600 ( \43198 , \43197 );
not \U$35601 ( \43199 , \43198 );
not \U$35602 ( \43200 , \43187 );
and \U$35603 ( \43201 , \43199 , \43200 );
nand \U$35604 ( \43202 , \43171 , \43180 );
nor \U$35605 ( \43203 , \43198 , \43202 );
nor \U$35606 ( \43204 , \43201 , \43203 );
not \U$35607 ( \43205 , \43204 );
and \U$35608 ( \43206 , \43205 , RIe3934b8_5560);
or \U$35609 ( \43207 , \43191 , \43206 );
not \U$35610 ( \43208 , RIe38b9e8_5572);
nand \U$35611 ( \43209 , \43193 , \43168 );
not \U$35612 ( \43210 , \43209 );
not \U$35613 ( \43211 , \43210 );
or \U$35614 ( \43212 , \43208 , \43211 );
not \U$35615 ( \43213 , \43209 );
and \U$35616 ( \43214 , RIe38a908_5574, \43213 );
not \U$35617 ( \43215 , \43198 );
not \U$35618 ( \43216 , \43150 );
and \U$35619 ( \43217 , \43215 , \43216 );
not \U$35620 ( \43218 , \43181 );
and \U$35621 ( \43219 , \43218 , \43150 );
or \U$35622 ( \43220 , \43217 , \43219 );
not \U$35623 ( \43221 , \43220 );
or \U$35624 ( \43222 , \43214 , \43221 );
nand \U$35625 ( \43223 , \43177 , \43173 );
not \U$35626 ( \43224 , \43174 );
or \U$35627 ( \43225 , \43150 , \43224 );
not \U$35628 ( \43226 , \43225 );
not \U$35629 ( \43227 , RIe392b58_5561);
and \U$35630 ( \43228 , \43226 , \43227 );
xnor \U$35631 ( \43229 , \43174 , \43184 );
not \U$35632 ( \43230 , \43229 );
and \U$35633 ( \43231 , \43230 , RIe392b58_5561);
or \U$35634 ( \43232 , \43228 , \43231 );
not \U$35635 ( \43233 , \43232 );
and \U$35636 ( \43234 , \43223 , \43233 );
or \U$35637 ( \43235 , \43182 , \43234 );
and \U$35638 ( \43236 , \43198 , RIe392b58_5561);
not \U$35639 ( \43237 , \43209 );
and \U$35640 ( \43238 , RIe38b1f0_5573, \43237 );
nor \U$35641 ( \43239 , \43236 , \43238 );
nand \U$35642 ( \43240 , \43235 , \43239 );
nor \U$35643 ( \43241 , \43222 , \43240 );
and \U$35644 ( \43242 , \43207 , \43212 , \43241 );
buf \U$35645 ( \43243 , RIb839668_156);
buf \U$35646 ( \43244 , \43243 );
not \U$35647 ( \43245 , \43244 );
not \U$35648 ( \43246 , \43245 );
buf \U$35649 ( \43247 , RIb839848_152);
and \U$35650 ( \43248 , \43247 , \38017 );
buf \U$35651 ( \43249 , RIb8396e0_155);
nand \U$35652 ( \43250 , \43249 , \38017 );
not \U$35653 ( \43251 , \43250 );
or \U$35654 ( \43252 , \43246 , \43248 , \43251 );
nand \U$35655 ( \43253 , \43252 , \38017 );
not \U$35656 ( \43254 , \43253 );
not \U$35657 ( \43255 , RIe38da40_5569);
or \U$35658 ( \43256 , \43254 , \43255 );
nand \U$35659 ( \43257 , \43250 , \43245 );
not \U$35660 ( \43258 , RIe38cf78_5570);
not \U$35661 ( \43259 , \43258 );
or \U$35662 ( \43260 , \43255 , \43259 );
not \U$35663 ( \43261 , \43260 );
nand \U$35664 ( \43262 , RIe38c4b0_5571, \43261 );
or \U$35665 ( \43263 , \43257 , \43262 );
xor \U$35666 ( \43264 , \43255 , \43258 );
nor \U$35667 ( \43265 , \43264 , \43261 );
nand \U$35668 ( \43266 , \38017 , \43250 , \43244 );
or \U$35669 ( \43267 , \43265 , \43266 );
not \U$35670 ( \43268 , \43257 );
nand \U$35671 ( \43269 , \43248 , \43262 , \43268 );
not \U$35672 ( \43270 , RIe38c4b0_5571);
nor \U$35673 ( \43271 , \43258 , \43270 );
xor \U$35674 ( \43272 , \43255 , \43271 );
or \U$35675 ( \43273 , \43269 , \43272 );
nand \U$35676 ( \43274 , \43256 , \43263 , \43267 , \43273 );
not \U$35677 ( \43275 , RIe393e90_5559);
not \U$35678 ( \43276 , RIe394868_5558);
not \U$35679 ( \43277 , RIe3951c8_5557);
not \U$35680 ( \43278 , \43277 );
nand \U$35681 ( \43279 , \43275 , \43276 , \43278 );
not \U$35682 ( \43280 , \43279 );
not \U$35683 ( \43281 , \43280 );
not \U$35684 ( \43282 , \43165 );
and \U$35685 ( \43283 , \43278 , \43282 );
nor \U$35686 ( \43284 , \43276 , \43275 );
xnor \U$35687 ( \43285 , \43277 , \43284 );
and \U$35688 ( \43286 , \43285 , \43165 );
or \U$35689 ( \43287 , \43283 , \43286 );
not \U$35690 ( \43288 , \43287 );
and \U$35691 ( \43289 , \43281 , \43288 );
nor \U$35692 ( \43290 , \43289 , \43169 );
not \U$35693 ( \43291 , \43290 );
or \U$35694 ( \43292 , \43274 , \43291 );
or \U$35695 ( \43293 , \43254 , \43270 );
or \U$35696 ( \43294 , \43257 , \43262 );
or \U$35697 ( \43295 , \43269 , RIe38c4b0_5571);
nand \U$35698 ( \43296 , \43244 , \38017 );
not \U$35699 ( \43297 , \43296 );
nand \U$35700 ( \43298 , \43297 , \43249 );
not \U$35701 ( \43299 , \43298 );
nand \U$35702 ( \43300 , RIe38c4b0_5571, \43260 );
and \U$35703 ( \43301 , \43262 , \43300 );
or \U$35704 ( \43302 , \43301 , \43296 );
and \U$35705 ( \43303 , \43302 , \43250 );
or \U$35706 ( \43304 , \43299 , \43303 );
nand \U$35707 ( \43305 , \43293 , \43294 , \43295 , \43304 );
not \U$35708 ( \43306 , \43305 );
xor \U$35709 ( \43307 , \43258 , \43270 );
not \U$35710 ( \43308 , \43269 );
and \U$35711 ( \43309 , \43307 , \43308 );
not \U$35712 ( \43310 , \43258 );
not \U$35713 ( \43311 , \43310 );
not \U$35714 ( \43312 , \43253 );
or \U$35715 ( \43313 , \43311 , \43312 );
not \U$35716 ( \43314 , \43266 );
nand \U$35717 ( \43315 , \43258 , \43260 , \43314 );
nand \U$35718 ( \43316 , \43313 , \43315 , \43298 );
or \U$35719 ( \43317 , \43309 , \43316 );
xor \U$35720 ( \43318 , \43276 , \43275 );
and \U$35721 ( \43319 , \43318 , \43279 , \43176 );
not \U$35722 ( \43320 , \43276 );
and \U$35723 ( \43321 , \43164 , \43320 , \43168 );
or \U$35724 ( \43322 , \43319 , \43321 );
not \U$35725 ( \43323 , \43322 );
or \U$35726 ( \43324 , \43317 , \43323 );
and \U$35727 ( \43325 , \43275 , \43279 , \43176 );
not \U$35728 ( \43326 , \43275 );
and \U$35729 ( \43327 , \43164 , \43326 , \43168 );
or \U$35730 ( \43328 , \43325 , \43327 );
not \U$35731 ( \43329 , \43328 );
nand \U$35732 ( \43330 , \43324 , \43329 );
or \U$35733 ( \43331 , \43306 , \43330 );
nand \U$35734 ( \43332 , \43317 , \43323 );
nand \U$35735 ( \43333 , \43331 , \43332 );
nand \U$35736 ( \43334 , \43292 , \43333 );
and \U$35737 ( \43335 , \43274 , \43291 );
not \U$35738 ( \43336 , RIe37f9b8_5584);
nor \U$35739 ( \43337 , \43335 , \43336 , \43022 );
and \U$35740 ( \43338 , \43334 , \43337 );
nor \U$35741 ( \43339 , \43242 , \43338 );
and \U$35743 ( \43340 , \43339 , 1'b1 );
or \U$35745 ( \43341 , \43340 , 1'b0 );
buf \U$35746 ( \43342 , \43341 );
_DC r23988_GF_IsGateDCbyConstraint ( \43343_nR23988 , \43342 , \21944 );
buf \U$35747 ( \43344 , \43343_nR23988 );
and \U$35749 ( \43345 , \43222 , 1'b1 );
or \U$35751 ( \43346 , \43345 , 1'b0 );
buf \U$35752 ( \43347 , \43346 );
_DC r239ba_GF_IsGateDCbyConstraint ( \43348_nR239ba , \43347 , \21944 );
buf \U$35753 ( \43349 , \43348_nR239ba );
and \U$35755 ( \43350 , \43240 , 1'b1 );
or \U$35757 ( \43351 , \43350 , 1'b0 );
buf \U$35758 ( \43352 , \43351 );
_DC r239bc_GF_IsGateDCbyConstraint ( \43353_nR239bc , \43352 , \21944 );
buf \U$35759 ( \43354 , \43353_nR239bc );
nand \U$35760 ( \43355 , \43212 , \43207 );
and \U$35762 ( \43356 , \43355 , 1'b1 );
or \U$35764 ( \43357 , \43356 , 1'b0 );
buf \U$35765 ( \43358 , \43357 );
_DC r239be_GF_IsGateDCbyConstraint ( \43359_nR239be , \43358 , \21944 );
buf \U$35766 ( \43360 , \43359_nR239be );
nand \U$35767 ( \43361 , \21810 , \21812 , RIe546098_6850);
nor \U$35768 ( \43362 , \21809 , \43361 );
buf \U$35769 ( \43363 , \43362 );
buf \U$35770 ( \43364 , \43363 );
buf \U$35771 ( \43365 , \27351 );
buf \U$35772 ( \43366 , \43365 );
nand \U$35773 ( \43367 , \43364 , \43366 );
buf \U$35774 ( \43368 , RIb79b518_270);
buf \U$35776 ( \43369 , \43368 );
not \U$35777 ( \43370 , \27247 );
and \U$35778 ( \43371 , \21694 , \43370 );
buf \U$35779 ( \43372 , \43371 );
buf \U$35780 ( \43373 , \43372 );
nand \U$35781 ( \43374 , \43369 , \43373 );
and \U$35782 ( \43375 , \43367 , \43374 );
not \U$35783 ( \43376 , \43375 );
buf \U$35784 ( \43377 , \43376 );
buf \U$35785 ( \43378 , \43377 );
not \U$35786 ( \43379 , \43378 );
and \U$35787 ( \43380 , RIe04cad8_4898, \43379 );
not \U$35788 ( \43381 , RIe04cad8_4898);
buf \U$35789 ( \43382 , RIe667bb0_6885);
buf \U$35790 ( \43383 , \43382 );
buf \U$35791 ( \43384 , RIe667f70_6886);
buf \U$35792 ( \43385 , \43384 );
not \U$35793 ( \43386 , \43385 );
not \U$35794 ( \43387 , \43386 );
or \U$35795 ( \43388 , \43383 , \43387 );
not \U$35796 ( \43389 , \43388 );
nand \U$35797 ( \43390 , \43374 , \43389 );
not \U$35798 ( \43391 , \27378 );
buf \U$35799 ( \43392 , \43391 );
not \U$35800 ( \43393 , \43392 );
not \U$35801 ( \43394 , \22119 );
buf \U$35802 ( \43395 , \43394 );
not \U$35803 ( \43396 , \43395 );
not \U$35804 ( \43397 , \43374 );
and \U$35805 ( \43398 , \43393 , \43396 , \43397 );
not \U$35806 ( \43399 , \43398 );
buf \U$35807 ( \43400 , \43399 );
and \U$35808 ( \43401 , \43390 , \43400 );
not \U$35809 ( \43402 , \43401 );
or \U$35810 ( \43403 , \43381 , \43402 );
not \U$35811 ( \43404 , \43390 );
buf \U$35812 ( \43405 , \43404 );
buf \U$35813 ( \43406 , RIb87eb00_69);
buf \U$35814 ( \43407 , \43406 );
and \U$35815 ( \43408 , \43405 , \43407 );
buf \U$35816 ( \43409 , \22134 );
not \U$35817 ( \43410 , \43400 );
and \U$35818 ( \43411 , \43409 , \43410 );
nor \U$35819 ( \43412 , \43408 , \43411 );
nand \U$35820 ( \43413 , \43403 , \43412 );
and \U$35821 ( \43414 , \43413 , \43378 );
or \U$35822 ( \43415 , \43380 , \43414 );
and \U$35824 ( \43416 , \43415 , 1'b1 );
or \U$35826 ( \43417 , \43416 , 1'b0 );
buf \U$35827 ( \43418 , \43417 );
_DC r234dc_GF_IsGateDCbyConstraint ( \43419_nR234dc , \43418 , \21944 );
buf \U$35828 ( \43420 , \43419_nR234dc );
not \U$35829 ( \43421 , \43378 );
and \U$35830 ( \43422 , RIe04b980_4899, \43421 );
not \U$35831 ( \43423 , RIe04b980_4899);
and \U$35832 ( \43424 , \43390 , \43400 );
not \U$35833 ( \43425 , \43424 );
or \U$35834 ( \43426 , \43423 , \43425 );
buf \U$35835 ( \43427 , \43404 );
buf \U$35836 ( \43428 , \32718 );
and \U$35837 ( \43429 , \43427 , \43428 );
buf \U$35838 ( \43430 , \32721 );
buf \U$35839 ( \43431 , \43399 );
not \U$35840 ( \43432 , \43431 );
and \U$35841 ( \43433 , \43430 , \43432 );
nor \U$35842 ( \43434 , \43429 , \43433 );
nand \U$35843 ( \43435 , \43426 , \43434 );
and \U$35844 ( \43436 , \43435 , \43378 );
or \U$35845 ( \43437 , \43422 , \43436 );
and \U$35847 ( \43438 , \43437 , 1'b1 );
or \U$35849 ( \43439 , \43438 , 1'b0 );
buf \U$35850 ( \43440 , \43439 );
_DC r234f2_GF_IsGateDCbyConstraint ( \43441_nR234f2 , \43440 , \21944 );
buf \U$35851 ( \43442 , \43441_nR234f2 );
not \U$35852 ( \43443 , \43378 );
and \U$35853 ( \43444 , RIe04a378_4900, \43443 );
not \U$35854 ( \43445 , RIe04a378_4900);
or \U$35855 ( \43446 , \43445 , \43402 );
buf \U$35856 ( \43447 , RIb87ebf0_67);
buf \U$35857 ( \43448 , \43447 );
and \U$35858 ( \43449 , \43405 , \43448 );
buf \U$35859 ( \43450 , \32742 );
not \U$35860 ( \43451 , \43400 );
and \U$35861 ( \43452 , \43450 , \43451 );
nor \U$35862 ( \43453 , \43449 , \43452 );
nand \U$35863 ( \43454 , \43446 , \43453 );
and \U$35864 ( \43455 , \43454 , \43378 );
or \U$35865 ( \43456 , \43444 , \43455 );
and \U$35867 ( \43457 , \43456 , 1'b1 );
or \U$35869 ( \43458 , \43457 , 1'b0 );
buf \U$35870 ( \43459 , \43458 );
_DC r23508_GF_IsGateDCbyConstraint ( \43460_nR23508 , \43459 , \21944 );
buf \U$35871 ( \43461 , \43460_nR23508 );
not \U$35872 ( \43462 , \43377 );
and \U$35873 ( \43463 , RIe049220_4901, \43462 );
not \U$35874 ( \43464 , RIe049220_4901);
not \U$35875 ( \43465 , \43424 );
or \U$35876 ( \43466 , \43464 , \43465 );
buf \U$35877 ( \43467 , RIb882ca0_66);
buf \U$35878 ( \43468 , \43467 );
and \U$35879 ( \43469 , \43427 , \43468 );
buf \U$35880 ( \43470 , \32763 );
not \U$35881 ( \43471 , \43400 );
and \U$35882 ( \43472 , \43470 , \43471 );
nor \U$35883 ( \43473 , \43469 , \43472 );
nand \U$35884 ( \43474 , \43466 , \43473 );
and \U$35885 ( \43475 , \43474 , \43377 );
or \U$35886 ( \43476 , \43463 , \43475 );
and \U$35888 ( \43477 , \43476 , 1'b1 );
or \U$35890 ( \43478 , \43477 , 1'b0 );
buf \U$35891 ( \43479 , \43478 );
_DC r2351e_GF_IsGateDCbyConstraint ( \43480_nR2351e , \43479 , \21944 );
buf \U$35892 ( \43481 , \43480_nR2351e );
buf \U$35893 ( \43482 , \43376 );
not \U$35894 ( \43483 , \43482 );
and \U$35895 ( \43484 , RIe047c18_4902, \43483 );
not \U$35896 ( \43485 , RIe047c18_4902);
not \U$35897 ( \43486 , \43401 );
or \U$35898 ( \43487 , \43485 , \43486 );
buf \U$35899 ( \43488 , \22223 );
and \U$35900 ( \43489 , \43405 , \43488 );
buf \U$35901 ( \43490 , RIb7cae58_233);
buf \U$35902 ( \43491 , \43490 );
not \U$35903 ( \43492 , \43431 );
and \U$35904 ( \43493 , \43491 , \43492 );
nor \U$35905 ( \43494 , \43489 , \43493 );
nand \U$35906 ( \43495 , \43487 , \43494 );
and \U$35907 ( \43496 , \43495 , \43482 );
or \U$35908 ( \43497 , \43484 , \43496 );
and \U$35910 ( \43498 , \43497 , 1'b1 );
or \U$35912 ( \43499 , \43498 , 1'b0 );
buf \U$35913 ( \43500 , \43499 );
_DC r23534_GF_IsGateDCbyConstraint ( \43501_nR23534 , \43500 , \21944 );
buf \U$35914 ( \43502 , \43501_nR23534 );
not \U$35915 ( \43503 , \43378 );
and \U$35916 ( \43504 , RIe046ac0_4903, \43503 );
not \U$35917 ( \43505 , RIe046ac0_4903);
not \U$35918 ( \43506 , \43424 );
or \U$35919 ( \43507 , \43505 , \43506 );
buf \U$35920 ( \43508 , RIb885388_64);
and \U$35921 ( \43509 , \43405 , \43508 );
buf \U$35922 ( \43510 , \27506 );
not \U$35923 ( \43511 , \43392 );
not \U$35924 ( \43512 , \43395 );
and \U$35925 ( \43513 , \43511 , \43512 , \43397 );
not \U$35926 ( \43514 , \43513 );
not \U$35927 ( \43515 , \43514 );
and \U$35928 ( \43516 , \43510 , \43515 );
nor \U$35929 ( \43517 , \43509 , \43516 );
nand \U$35930 ( \43518 , \43507 , \43517 );
and \U$35931 ( \43519 , \43518 , \43378 );
or \U$35932 ( \43520 , \43504 , \43519 );
and \U$35934 ( \43521 , \43520 , 1'b1 );
or \U$35936 ( \43522 , \43521 , 1'b0 );
buf \U$35937 ( \43523 , \43522 );
_DC r2354a_GF_IsGateDCbyConstraint ( \43524_nR2354a , \43523 , \21944 );
buf \U$35938 ( \43525 , \43524_nR2354a );
not \U$35939 ( \43526 , \43378 );
and \U$35940 ( \43527 , RIe045968_4904, \43526 );
not \U$35941 ( \43528 , RIe045968_4904);
not \U$35942 ( \43529 , \43401 );
or \U$35943 ( \43530 , \43528 , \43529 );
buf \U$35944 ( \43531 , RIb885400_63);
buf \U$35945 ( \43532 , \43531 );
and \U$35946 ( \43533 , \43405 , \43532 );
buf \U$35947 ( \43534 , RIb7caf48_231);
buf \U$35948 ( \43535 , \43534 );
not \U$35949 ( \43536 , \43400 );
and \U$35950 ( \43537 , \43535 , \43536 );
nor \U$35951 ( \43538 , \43533 , \43537 );
nand \U$35952 ( \43539 , \43530 , \43538 );
and \U$35953 ( \43540 , \43539 , \43378 );
or \U$35954 ( \43541 , \43527 , \43540 );
and \U$35956 ( \43542 , \43541 , 1'b1 );
or \U$35958 ( \43543 , \43542 , 1'b0 );
buf \U$35959 ( \43544 , \43543 );
_DC r23554_GF_IsGateDCbyConstraint ( \43545_nR23554 , \43544 , \21944 );
buf \U$35960 ( \43546 , \43545_nR23554 );
not \U$35961 ( \43547 , \43378 );
and \U$35962 ( \43548 , RIe044360_4905, \43547 );
not \U$35963 ( \43549 , RIe044360_4905);
or \U$35964 ( \43550 , \43549 , \43506 );
buf \U$35965 ( \43551 , \43404 );
buf \U$35966 ( \43552 , RIb885478_62);
buf \U$35967 ( \43553 , \43552 );
and \U$35968 ( \43554 , \43551 , \43553 );
buf \U$35969 ( \43555 , \27545 );
buf \U$35970 ( \43556 , \43514 );
not \U$35971 ( \43557 , \43556 );
and \U$35972 ( \43558 , \43555 , \43557 );
nor \U$35973 ( \43559 , \43554 , \43558 );
nand \U$35974 ( \43560 , \43550 , \43559 );
and \U$35975 ( \43561 , \43560 , \43378 );
or \U$35976 ( \43562 , \43548 , \43561 );
and \U$35978 ( \43563 , \43562 , 1'b1 );
or \U$35980 ( \43564 , \43563 , 1'b0 );
buf \U$35981 ( \43565 , \43564 );
_DC r23556_GF_IsGateDCbyConstraint ( \43566_nR23556 , \43565 , \21944 );
buf \U$35982 ( \43567 , \43566_nR23556 );
buf \U$35983 ( \43568 , \43377 );
not \U$35984 ( \43569 , \43568 );
and \U$35985 ( \43570 , RIe043208_4906, \43569 );
not \U$35986 ( \43571 , RIe043208_4906);
or \U$35987 ( \43572 , \43571 , \43465 );
buf \U$35988 ( \43573 , \27564 );
and \U$35989 ( \43574 , \43427 , \43573 );
buf \U$35990 ( \43575 , RIb7cb038_229);
buf \U$35991 ( \43576 , \43575 );
buf \U$35992 ( \43577 , \43399 );
not \U$35993 ( \43578 , \43577 );
and \U$35994 ( \43579 , \43576 , \43578 );
nor \U$35995 ( \43580 , \43574 , \43579 );
nand \U$35996 ( \43581 , \43572 , \43580 );
and \U$35997 ( \43582 , \43581 , \43568 );
or \U$35998 ( \43583 , \43570 , \43582 );
and \U$36000 ( \43584 , \43583 , 1'b1 );
or \U$36002 ( \43585 , \43584 , 1'b0 );
buf \U$36003 ( \43586 , \43585 );
_DC r23558_GF_IsGateDCbyConstraint ( \43587_nR23558 , \43586 , \21944 );
buf \U$36004 ( \43588 , \43587_nR23558 );
buf \U$36005 ( \43589 , \43376 );
not \U$36006 ( \43590 , \43589 );
and \U$36007 ( \43591 , RIe041c00_4907, \43590 );
not \U$36008 ( \43592 , RIe041c00_4907);
or \U$36009 ( \43593 , \43592 , \43506 );
buf \U$36010 ( \43594 , RIb885568_60);
buf \U$36011 ( \43595 , \43594 );
and \U$36012 ( \43596 , \43551 , \43595 );
buf \U$36013 ( \43597 , \32893 );
not \U$36014 ( \43598 , \43392 );
not \U$36015 ( \43599 , \43395 );
and \U$36016 ( \43600 , \43598 , \43599 , \43397 );
not \U$36017 ( \43601 , \43600 );
not \U$36018 ( \43602 , \43601 );
and \U$36019 ( \43603 , \43597 , \43602 );
nor \U$36020 ( \43604 , \43596 , \43603 );
nand \U$36021 ( \43605 , \43593 , \43604 );
and \U$36022 ( \43606 , \43605 , \43589 );
or \U$36023 ( \43607 , \43591 , \43606 );
and \U$36025 ( \43608 , \43607 , 1'b1 );
or \U$36027 ( \43609 , \43608 , 1'b0 );
buf \U$36028 ( \43610 , \43609 );
_DC r2355a_GF_IsGateDCbyConstraint ( \43611_nR2355a , \43610 , \21944 );
buf \U$36029 ( \43612 , \43611_nR2355a );
not \U$36030 ( \43613 , \43378 );
and \U$36031 ( \43614 , RIe040aa8_4908, \43613 );
not \U$36032 ( \43615 , RIe040aa8_4908);
not \U$36033 ( \43616 , \43401 );
or \U$36034 ( \43617 , \43615 , \43616 );
buf \U$36035 ( \43618 , RIb8855e0_59);
buf \U$36036 ( \43619 , \43618 );
and \U$36037 ( \43620 , \43427 , \43619 );
buf \U$36038 ( \43621 , RIb7cb128_227);
buf \U$36039 ( \43622 , \43621 );
not \U$36040 ( \43623 , \43431 );
and \U$36041 ( \43624 , \43622 , \43623 );
nor \U$36042 ( \43625 , \43620 , \43624 );
nand \U$36043 ( \43626 , \43617 , \43625 );
and \U$36044 ( \43627 , \43626 , \43378 );
or \U$36045 ( \43628 , \43614 , \43627 );
and \U$36047 ( \43629 , \43628 , 1'b1 );
or \U$36049 ( \43630 , \43629 , 1'b0 );
buf \U$36050 ( \43631 , \43630 );
_DC r234de_GF_IsGateDCbyConstraint ( \43632_nR234de , \43631 , \21944 );
buf \U$36051 ( \43633 , \43632_nR234de );
not \U$36052 ( \43634 , \43568 );
and \U$36053 ( \43635 , RIe03f4a0_4909, \43634 );
not \U$36054 ( \43636 , RIe03f4a0_4909);
or \U$36055 ( \43637 , \43636 , \43486 );
buf \U$36056 ( \43638 , RIb885658_58);
and \U$36057 ( \43639 , \43551 , \43638 );
buf \U$36058 ( \43640 , \27627 );
not \U$36059 ( \43641 , \43556 );
and \U$36060 ( \43642 , \43640 , \43641 );
nor \U$36061 ( \43643 , \43639 , \43642 );
nand \U$36062 ( \43644 , \43637 , \43643 );
and \U$36063 ( \43645 , \43644 , \43568 );
or \U$36064 ( \43646 , \43635 , \43645 );
and \U$36066 ( \43647 , \43646 , 1'b1 );
or \U$36068 ( \43648 , \43647 , 1'b0 );
buf \U$36069 ( \43649 , \43648 );
_DC r234e0_GF_IsGateDCbyConstraint ( \43650_nR234e0 , \43649 , \21944 );
buf \U$36070 ( \43651 , \43650_nR234e0 );
not \U$36071 ( \43652 , \43378 );
and \U$36072 ( \43653 , RIe03e348_4910, \43652 );
not \U$36073 ( \43654 , RIe03e348_4910);
not \U$36074 ( \43655 , \43401 );
or \U$36075 ( \43656 , \43654 , \43655 );
buf \U$36076 ( \43657 , RIb8856d0_57);
buf \U$36077 ( \43658 , \43657 );
and \U$36078 ( \43659 , \43427 , \43658 );
buf \U$36079 ( \43660 , RIb8263d8_225);
buf \U$36080 ( \43661 , \43660 );
not \U$36081 ( \43662 , \43577 );
and \U$36082 ( \43663 , \43661 , \43662 );
nor \U$36083 ( \43664 , \43659 , \43663 );
nand \U$36084 ( \43665 , \43656 , \43664 );
and \U$36085 ( \43666 , \43665 , \43378 );
or \U$36086 ( \43667 , \43653 , \43666 );
and \U$36088 ( \43668 , \43667 , 1'b1 );
or \U$36090 ( \43669 , \43668 , 1'b0 );
buf \U$36091 ( \43670 , \43669 );
_DC r234e2_GF_IsGateDCbyConstraint ( \43671_nR234e2 , \43670 , \21944 );
buf \U$36092 ( \43672 , \43671_nR234e2 );
not \U$36093 ( \43673 , \43378 );
and \U$36094 ( \43674 , RIe03d1f0_4911, \43673 );
not \U$36095 ( \43675 , RIe03d1f0_4911);
or \U$36096 ( \43676 , \43675 , \43425 );
buf \U$36097 ( \43677 , RIb885748_56);
buf \U$36098 ( \43678 , \43677 );
and \U$36099 ( \43679 , \43551 , \43678 );
buf \U$36100 ( \43680 , \27667 );
not \U$36101 ( \43681 , \43601 );
and \U$36102 ( \43682 , \43680 , \43681 );
nor \U$36103 ( \43683 , \43679 , \43682 );
nand \U$36104 ( \43684 , \43676 , \43683 );
and \U$36105 ( \43685 , \43684 , \43378 );
or \U$36106 ( \43686 , \43674 , \43685 );
and \U$36108 ( \43687 , \43686 , 1'b1 );
or \U$36110 ( \43688 , \43687 , 1'b0 );
buf \U$36111 ( \43689 , \43688 );
_DC r234e4_GF_IsGateDCbyConstraint ( \43690_nR234e4 , \43689 , \21944 );
buf \U$36112 ( \43691 , \43690_nR234e4 );
not \U$36113 ( \43692 , \43568 );
and \U$36114 ( \43693 , RIde08bc0_4912, \43692 );
not \U$36115 ( \43694 , RIde08bc0_4912);
or \U$36116 ( \43695 , \43694 , \43465 );
buf \U$36117 ( \43696 , \32990 );
and \U$36118 ( \43697 , \43427 , \43696 );
buf \U$36119 ( \43698 , \32993 );
not \U$36120 ( \43699 , \43601 );
and \U$36121 ( \43700 , \43698 , \43699 );
nor \U$36122 ( \43701 , \43697 , \43700 );
nand \U$36123 ( \43702 , \43695 , \43701 );
and \U$36124 ( \43703 , \43702 , \43568 );
or \U$36125 ( \43704 , \43693 , \43703 );
and \U$36127 ( \43705 , \43704 , 1'b1 );
or \U$36129 ( \43706 , \43705 , 1'b0 );
buf \U$36130 ( \43707 , \43706 );
_DC r234e6_GF_IsGateDCbyConstraint ( \43708_nR234e6 , \43707 , \21944 );
buf \U$36131 ( \43709 , \43708_nR234e6 );
buf \U$36132 ( \43710 , \43376 );
not \U$36133 ( \43711 , \43710 );
and \U$36134 ( \43712 , RIde0d030_4913, \43711 );
not \U$36135 ( \43713 , RIde0d030_4913);
or \U$36136 ( \43714 , \43713 , \43402 );
buf \U$36137 ( \43715 , \33010 );
and \U$36138 ( \43716 , \43427 , \43715 );
buf \U$36139 ( \43717 , RIb826f18_222);
buf \U$36140 ( \43718 , \43717 );
not \U$36141 ( \43719 , \43577 );
and \U$36142 ( \43720 , \43718 , \43719 );
nor \U$36143 ( \43721 , \43716 , \43720 );
nand \U$36144 ( \43722 , \43714 , \43721 );
and \U$36145 ( \43723 , \43722 , \43710 );
or \U$36146 ( \43724 , \43712 , \43723 );
and \U$36148 ( \43725 , \43724 , 1'b1 );
or \U$36150 ( \43726 , \43725 , 1'b0 );
buf \U$36151 ( \43727 , \43726 );
_DC r234e8_GF_IsGateDCbyConstraint ( \43728_nR234e8 , \43727 , \21944 );
buf \U$36152 ( \43729 , \43728_nR234e8 );
buf \U$36153 ( \43730 , \43376 );
not \U$36154 ( \43731 , \43730 );
and \U$36155 ( \43732 , RIde131b0_4914, \43731 );
not \U$36156 ( \43733 , RIde131b0_4914);
or \U$36157 ( \43734 , \43733 , \43616 );
buf \U$36158 ( \43735 , RIb8858b0_53);
buf \U$36159 ( \43736 , \43735 );
and \U$36160 ( \43737 , \43404 , \43736 );
buf \U$36161 ( \43738 , \33032 );
not \U$36162 ( \43739 , \43431 );
and \U$36163 ( \43740 , \43738 , \43739 );
nor \U$36164 ( \43741 , \43737 , \43740 );
nand \U$36165 ( \43742 , \43734 , \43741 );
and \U$36166 ( \43743 , \43742 , \43730 );
or \U$36167 ( \43744 , \43732 , \43743 );
and \U$36169 ( \43745 , \43744 , 1'b1 );
or \U$36171 ( \43746 , \43745 , 1'b0 );
buf \U$36172 ( \43747 , \43746 );
_DC r234ea_GF_IsGateDCbyConstraint ( \43748_nR234ea , \43747 , \21944 );
buf \U$36173 ( \43749 , \43748_nR234ea );
not \U$36174 ( \43750 , \43568 );
and \U$36175 ( \43751 , RIde17968_4915, \43750 );
not \U$36176 ( \43752 , RIde17968_4915);
or \U$36177 ( \43753 , \43752 , \43486 );
buf \U$36178 ( \43754 , \33049 );
and \U$36179 ( \43755 , \43551 , \43754 );
buf \U$36180 ( \43756 , \27740 );
not \U$36181 ( \43757 , \43577 );
and \U$36182 ( \43758 , \43756 , \43757 );
nor \U$36183 ( \43759 , \43755 , \43758 );
nand \U$36184 ( \43760 , \43753 , \43759 );
and \U$36185 ( \43761 , \43760 , \43568 );
or \U$36186 ( \43762 , \43751 , \43761 );
and \U$36188 ( \43763 , \43762 , 1'b1 );
or \U$36190 ( \43764 , \43763 , 1'b0 );
buf \U$36191 ( \43765 , \43764 );
_DC r234ec_GF_IsGateDCbyConstraint ( \43766_nR234ec , \43765 , \21944 );
buf \U$36192 ( \43767 , \43766_nR234ec );
not \U$36193 ( \43768 , \43482 );
and \U$36194 ( \43769 , RIde1f528_4916, \43768 );
not \U$36195 ( \43770 , RIde1f528_4916);
or \U$36196 ( \43771 , \43770 , \43655 );
buf \U$36197 ( \43772 , RIb8859a0_51);
buf \U$36198 ( \43773 , \43772 );
and \U$36199 ( \43774 , \43405 , \43773 );
buf \U$36200 ( \43775 , RIb829420_219);
buf \U$36201 ( \43776 , \43775 );
not \U$36202 ( \43777 , \43431 );
and \U$36203 ( \43778 , \43776 , \43777 );
nor \U$36204 ( \43779 , \43774 , \43778 );
nand \U$36205 ( \43780 , \43771 , \43779 );
and \U$36206 ( \43781 , \43780 , \43482 );
or \U$36207 ( \43782 , \43769 , \43781 );
and \U$36209 ( \43783 , \43782 , 1'b1 );
or \U$36211 ( \43784 , \43783 , 1'b0 );
buf \U$36212 ( \43785 , \43784 );
_DC r234ee_GF_IsGateDCbyConstraint ( \43786_nR234ee , \43785 , \21944 );
buf \U$36213 ( \43787 , \43786_nR234ee );
not \U$36214 ( \43788 , \43378 );
and \U$36215 ( \43789 , RIde24e38_4917, \43788 );
not \U$36216 ( \43790 , RIde24e38_4917);
or \U$36217 ( \43791 , \43790 , \43529 );
buf \U$36218 ( \43792 , \22538 );
and \U$36219 ( \43793 , \43551 , \43792 );
buf \U$36220 ( \43794 , RIb829498_218);
buf \U$36221 ( \43795 , \43794 );
not \U$36222 ( \43796 , \43400 );
and \U$36223 ( \43797 , \43795 , \43796 );
nor \U$36224 ( \43798 , \43793 , \43797 );
nand \U$36225 ( \43799 , \43791 , \43798 );
and \U$36226 ( \43800 , \43799 , \43378 );
or \U$36227 ( \43801 , \43789 , \43800 );
and \U$36229 ( \43802 , \43801 , 1'b1 );
or \U$36231 ( \43803 , \43802 , 1'b0 );
buf \U$36232 ( \43804 , \43803 );
_DC r234f0_GF_IsGateDCbyConstraint ( \43805_nR234f0 , \43804 , \21944 );
buf \U$36233 ( \43806 , \43805_nR234f0 );
not \U$36234 ( \43807 , \43568 );
and \U$36235 ( \43808 , RIde29ed8_4918, \43807 );
not \U$36236 ( \43809 , RIde29ed8_4918);
or \U$36237 ( \43810 , \43809 , \43465 );
buf \U$36238 ( \43811 , \27795 );
and \U$36239 ( \43812 , \43551 , \43811 );
buf \U$36240 ( \43813 , \27798 );
not \U$36241 ( \43814 , \43577 );
and \U$36242 ( \43815 , \43813 , \43814 );
nor \U$36243 ( \43816 , \43812 , \43815 );
nand \U$36244 ( \43817 , \43810 , \43816 );
and \U$36245 ( \43818 , \43817 , \43568 );
or \U$36246 ( \43819 , \43808 , \43818 );
and \U$36248 ( \43820 , \43819 , 1'b1 );
or \U$36250 ( \43821 , \43820 , 1'b0 );
buf \U$36251 ( \43822 , \43821 );
_DC r234f4_GF_IsGateDCbyConstraint ( \43823_nR234f4 , \43822 , \21944 );
buf \U$36252 ( \43824 , \43823_nR234f4 );
not \U$36253 ( \43825 , \43589 );
and \U$36254 ( \43826 , RIde31390_4919, \43825 );
not \U$36255 ( \43827 , RIde31390_4919);
or \U$36256 ( \43828 , \43827 , \43506 );
buf \U$36257 ( \43829 , RIb885b08_48);
buf \U$36258 ( \43830 , \43829 );
and \U$36259 ( \43831 , \43404 , \43830 );
buf \U$36260 ( \43832 , \33128 );
not \U$36261 ( \43833 , \43431 );
and \U$36262 ( \43834 , \43832 , \43833 );
nor \U$36263 ( \43835 , \43831 , \43834 );
nand \U$36264 ( \43836 , \43828 , \43835 );
and \U$36265 ( \43837 , \43836 , \43589 );
or \U$36266 ( \43838 , \43826 , \43837 );
and \U$36268 ( \43839 , \43838 , 1'b1 );
or \U$36270 ( \43840 , \43839 , 1'b0 );
buf \U$36271 ( \43841 , \43840 );
_DC r234f6_GF_IsGateDCbyConstraint ( \43842_nR234f6 , \43841 , \21944 );
buf \U$36272 ( \43843 , \43842_nR234f6 );
not \U$36273 ( \43844 , \43589 );
and \U$36274 ( \43845 , RIde36e08_4920, \43844 );
not \U$36275 ( \43846 , RIde36e08_4920);
or \U$36276 ( \43847 , \43846 , \43529 );
not \U$36277 ( \43848 , \43390 );
buf \U$36278 ( \43849 , \33145 );
and \U$36279 ( \43850 , \43848 , \43849 );
buf \U$36280 ( \43851 , RIb829600_215);
buf \U$36281 ( \43852 , \43851 );
not \U$36282 ( \43853 , \43556 );
and \U$36283 ( \43854 , \43852 , \43853 );
nor \U$36284 ( \43855 , \43850 , \43854 );
nand \U$36285 ( \43856 , \43847 , \43855 );
and \U$36286 ( \43857 , \43856 , \43589 );
or \U$36287 ( \43858 , \43845 , \43857 );
and \U$36289 ( \43859 , \43858 , 1'b1 );
or \U$36291 ( \43860 , \43859 , 1'b0 );
buf \U$36292 ( \43861 , \43860 );
_DC r234f8_GF_IsGateDCbyConstraint ( \43862_nR234f8 , \43861 , \21944 );
buf \U$36293 ( \43863 , \43862_nR234f8 );
not \U$36294 ( \43864 , \43568 );
and \U$36295 ( \43865 , RIde3efe0_4921, \43864 );
not \U$36296 ( \43866 , RIde3efe0_4921);
or \U$36297 ( \43867 , \43866 , \43506 );
buf \U$36298 ( \43868 , RIb885bf8_46);
buf \U$36299 ( \43869 , \43868 );
and \U$36300 ( \43870 , \43404 , \43869 );
buf \U$36301 ( \43871 , RIb829678_214);
buf \U$36302 ( \43872 , \43871 );
not \U$36303 ( \43873 , \43556 );
and \U$36304 ( \43874 , \43872 , \43873 );
nor \U$36305 ( \43875 , \43870 , \43874 );
nand \U$36306 ( \43876 , \43867 , \43875 );
and \U$36307 ( \43877 , \43876 , \43568 );
or \U$36308 ( \43878 , \43865 , \43877 );
and \U$36310 ( \43879 , \43878 , 1'b1 );
or \U$36312 ( \43880 , \43879 , 1'b0 );
buf \U$36313 ( \43881 , \43880 );
_DC r234fa_GF_IsGateDCbyConstraint ( \43882_nR234fa , \43881 , \21944 );
buf \U$36314 ( \43883 , \43882_nR234fa );
not \U$36315 ( \43884 , \43378 );
and \U$36316 ( \43885 , RIde45070_4922, \43884 );
not \U$36317 ( \43886 , RIde45070_4922);
or \U$36318 ( \43887 , \43886 , \43465 );
buf \U$36319 ( \43888 , \22639 );
and \U$36320 ( \43889 , \43551 , \43888 );
buf \U$36321 ( \43890 , \27872 );
not \U$36322 ( \43891 , \43400 );
and \U$36323 ( \43892 , \43890 , \43891 );
nor \U$36324 ( \43893 , \43889 , \43892 );
nand \U$36325 ( \43894 , \43887 , \43893 );
and \U$36326 ( \43895 , \43894 , \43378 );
or \U$36327 ( \43896 , \43885 , \43895 );
and \U$36329 ( \43897 , \43896 , 1'b1 );
or \U$36331 ( \43898 , \43897 , 1'b0 );
buf \U$36332 ( \43899 , \43898 );
_DC r234fc_GF_IsGateDCbyConstraint ( \43900_nR234fc , \43899 , \21944 );
buf \U$36333 ( \43901 , \43900_nR234fc );
not \U$36334 ( \43902 , \43378 );
and \U$36335 ( \43903 , RIde4c9d8_4923, \43902 );
not \U$36336 ( \43904 , RIde4c9d8_4923);
or \U$36337 ( \43905 , \43904 , \43506 );
buf \U$36338 ( \43906 , RIb885ce8_44);
buf \U$36339 ( \43907 , \43906 );
and \U$36340 ( \43908 , \43404 , \43907 );
buf \U$36341 ( \43909 , RIb82dae8_212);
buf \U$36342 ( \43910 , \43909 );
not \U$36343 ( \43911 , \43556 );
and \U$36344 ( \43912 , \43910 , \43911 );
nor \U$36345 ( \43913 , \43908 , \43912 );
nand \U$36346 ( \43914 , \43905 , \43913 );
and \U$36347 ( \43915 , \43914 , \43378 );
or \U$36348 ( \43916 , \43903 , \43915 );
and \U$36350 ( \43917 , \43916 , 1'b1 );
or \U$36352 ( \43918 , \43917 , 1'b0 );
buf \U$36353 ( \43919 , \43918 );
_DC r234fe_GF_IsGateDCbyConstraint ( \43920_nR234fe , \43919 , \21944 );
buf \U$36354 ( \43921 , \43920_nR234fe );
not \U$36355 ( \43922 , \43568 );
and \U$36356 ( \43923 , RIde51b68_4924, \43922 );
not \U$36357 ( \43924 , RIde51b68_4924);
or \U$36358 ( \43925 , \43924 , \43425 );
buf \U$36359 ( \43926 , RIb885d60_43);
buf \U$36360 ( \43927 , \43926 );
and \U$36361 ( \43928 , \43427 , \43927 );
buf \U$36362 ( \43929 , \33225 );
not \U$36363 ( \43930 , \43577 );
and \U$36364 ( \43931 , \43929 , \43930 );
nor \U$36365 ( \43932 , \43928 , \43931 );
nand \U$36366 ( \43933 , \43925 , \43932 );
and \U$36367 ( \43934 , \43933 , \43568 );
or \U$36368 ( \43935 , \43923 , \43934 );
and \U$36370 ( \43936 , \43935 , 1'b1 );
or \U$36372 ( \43937 , \43936 , 1'b0 );
buf \U$36373 ( \43938 , \43937 );
_DC r23500_GF_IsGateDCbyConstraint ( \43939_nR23500 , \43938 , \21944 );
buf \U$36374 ( \43940 , \43939_nR23500 );
not \U$36375 ( \43941 , \43589 );
and \U$36376 ( \43942 , RIde553a8_4925, \43941 );
not \U$36377 ( \43943 , RIde553a8_4925);
or \U$36378 ( \43944 , \43943 , \43465 );
buf \U$36379 ( \43945 , RIb885dd8_42);
buf \U$36380 ( \43946 , \43945 );
and \U$36381 ( \43947 , \43404 , \43946 );
buf \U$36382 ( \43948 , RIb82dbd8_210);
buf \U$36383 ( \43949 , \43948 );
not \U$36384 ( \43950 , \43601 );
and \U$36385 ( \43951 , \43949 , \43950 );
nor \U$36386 ( \43952 , \43947 , \43951 );
nand \U$36387 ( \43953 , \43944 , \43952 );
and \U$36388 ( \43954 , \43953 , \43589 );
or \U$36389 ( \43955 , \43942 , \43954 );
and \U$36391 ( \43956 , \43955 , 1'b1 );
or \U$36393 ( \43957 , \43956 , 1'b0 );
buf \U$36394 ( \43958 , \43957 );
_DC r23502_GF_IsGateDCbyConstraint ( \43959_nR23502 , \43958 , \21944 );
buf \U$36395 ( \43960 , \43959_nR23502 );
buf \U$36396 ( \43961 , \43376 );
not \U$36397 ( \43962 , \43961 );
and \U$36398 ( \43963 , RIde59c50_4926, \43962 );
not \U$36399 ( \43964 , RIde59c50_4926);
or \U$36400 ( \43965 , \43964 , \43425 );
buf \U$36401 ( \43966 , \38608 );
and \U$36402 ( \43967 , \43427 , \43966 );
buf \U$36403 ( \43968 , RIb82dc50_209);
buf \U$36404 ( \43969 , \43968 );
not \U$36405 ( \43970 , \43577 );
and \U$36406 ( \43971 , \43969 , \43970 );
nor \U$36407 ( \43972 , \43967 , \43971 );
nand \U$36408 ( \43973 , \43965 , \43972 );
and \U$36409 ( \43974 , \43973 , \43961 );
or \U$36410 ( \43975 , \43963 , \43974 );
and \U$36412 ( \43976 , \43975 , 1'b1 );
or \U$36414 ( \43977 , \43976 , 1'b0 );
buf \U$36415 ( \43978 , \43977 );
_DC r23504_GF_IsGateDCbyConstraint ( \43979_nR23504 , \43978 , \21944 );
buf \U$36416 ( \43980 , \43979_nR23504 );
not \U$36417 ( \43981 , \43568 );
and \U$36418 ( \43982 , RIde5e390_4927, \43981 );
not \U$36419 ( \43983 , RIde5e390_4927);
or \U$36420 ( \43984 , \43983 , \43506 );
buf \U$36421 ( \43985 , \22740 );
and \U$36422 ( \43986 , \43405 , \43985 );
buf \U$36423 ( \43987 , \33283 );
not \U$36424 ( \43988 , \43577 );
and \U$36425 ( \43989 , \43987 , \43988 );
nor \U$36426 ( \43990 , \43986 , \43989 );
nand \U$36427 ( \43991 , \43984 , \43990 );
and \U$36428 ( \43992 , \43991 , \43568 );
or \U$36429 ( \43993 , \43982 , \43992 );
and \U$36431 ( \43994 , \43993 , 1'b1 );
or \U$36433 ( \43995 , \43994 , 1'b0 );
buf \U$36434 ( \43996 , \43995 );
_DC r23506_GF_IsGateDCbyConstraint ( \43997_nR23506 , \43996 , \21944 );
buf \U$36435 ( \43998 , \43997_nR23506 );
not \U$36436 ( \43999 , \43377 );
and \U$36437 ( \44000 , RIde65668_4928, \43999 );
not \U$36438 ( \44001 , RIde65668_4928);
or \U$36439 ( \44002 , \44001 , \43616 );
buf \U$36440 ( \44003 , RIb885f40_39);
and \U$36441 ( \44004 , \43427 , \44003 );
buf \U$36442 ( \44005 , RIb82dd40_207);
buf \U$36443 ( \44006 , \44005 );
not \U$36444 ( \44007 , \43431 );
and \U$36445 ( \44008 , \44006 , \44007 );
nor \U$36446 ( \44009 , \44004 , \44008 );
nand \U$36447 ( \44010 , \44002 , \44009 );
and \U$36448 ( \44011 , \44010 , \43377 );
or \U$36449 ( \44012 , \44000 , \44011 );
and \U$36451 ( \44013 , \44012 , 1'b1 );
or \U$36453 ( \44014 , \44013 , 1'b0 );
buf \U$36454 ( \44015 , \44014 );
_DC r2350a_GF_IsGateDCbyConstraint ( \44016_nR2350a , \44015 , \21944 );
buf \U$36455 ( \44017 , \44016_nR2350a );
buf \U$36456 ( \44018 , \43376 );
not \U$36457 ( \44019 , \44018 );
and \U$36458 ( \44020 , RIde6a4b0_4929, \44019 );
not \U$36459 ( \44021 , RIde6a4b0_4929);
or \U$36460 ( \44022 , \44021 , \43402 );
buf \U$36461 ( \44023 , \38669 );
and \U$36462 ( \44024 , \43551 , \44023 );
buf \U$36463 ( \44025 , \28008 );
not \U$36464 ( \44026 , \43577 );
and \U$36465 ( \44027 , \44025 , \44026 );
nor \U$36466 ( \44028 , \44024 , \44027 );
nand \U$36467 ( \44029 , \44022 , \44028 );
and \U$36468 ( \44030 , \44029 , \44018 );
or \U$36469 ( \44031 , \44020 , \44030 );
and \U$36471 ( \44032 , \44031 , 1'b1 );
or \U$36473 ( \44033 , \44032 , 1'b0 );
buf \U$36474 ( \44034 , \44033 );
_DC r2350c_GF_IsGateDCbyConstraint ( \44035_nR2350c , \44034 , \21944 );
buf \U$36475 ( \44036 , \44035_nR2350c );
not \U$36476 ( \44037 , \43568 );
and \U$36477 ( \44038 , RIde6f820_4930, \44037 );
not \U$36478 ( \44039 , RIde6f820_4930);
or \U$36479 ( \44040 , \44039 , \43616 );
buf \U$36480 ( \44041 , \38689 );
and \U$36481 ( \44042 , \43427 , \44041 );
buf \U$36482 ( \44043 , \28028 );
not \U$36483 ( \44044 , \43431 );
and \U$36484 ( \44045 , \44043 , \44044 );
nor \U$36485 ( \44046 , \44042 , \44045 );
nand \U$36486 ( \44047 , \44040 , \44046 );
and \U$36487 ( \44048 , \44047 , \43568 );
or \U$36488 ( \44049 , \44038 , \44048 );
and \U$36490 ( \44050 , \44049 , 1'b1 );
or \U$36492 ( \44051 , \44050 , 1'b0 );
buf \U$36493 ( \44052 , \44051 );
_DC r2350e_GF_IsGateDCbyConstraint ( \44053_nR2350e , \44052 , \21944 );
buf \U$36494 ( \44054 , \44053_nR2350e );
not \U$36495 ( \44055 , \43961 );
and \U$36496 ( \44056 , RIdf73710_4931, \44055 );
not \U$36497 ( \44057 , RIdf73710_4931);
or \U$36498 ( \44058 , \44057 , \43486 );
buf \U$36499 ( \44059 , RIb8860a8_36);
buf \U$36500 ( \44060 , \44059 );
and \U$36501 ( \44061 , \43405 , \44060 );
buf \U$36502 ( \44062 , \28047 );
not \U$36503 ( \44063 , \43601 );
and \U$36504 ( \44064 , \44062 , \44063 );
nor \U$36505 ( \44065 , \44061 , \44064 );
nand \U$36506 ( \44066 , \44058 , \44065 );
and \U$36507 ( \44067 , \44066 , \43961 );
or \U$36508 ( \44068 , \44056 , \44067 );
and \U$36510 ( \44069 , \44068 , 1'b1 );
or \U$36512 ( \44070 , \44069 , 1'b0 );
buf \U$36513 ( \44071 , \44070 );
_DC r23510_GF_IsGateDCbyConstraint ( \44072_nR23510 , \44071 , \21944 );
buf \U$36514 ( \44073 , \44072_nR23510 );
buf \U$36515 ( \44074 , \43376 );
not \U$36516 ( \44075 , \44074 );
and \U$36517 ( \44076 , RIdc38040_4932, \44075 );
not \U$36518 ( \44077 , RIdc38040_4932);
or \U$36519 ( \44078 , \44077 , \43655 );
buf \U$36520 ( \44079 , \22842 );
and \U$36521 ( \44080 , \43405 , \44079 );
buf \U$36522 ( \44081 , RIb8322a0_203);
buf \U$36523 ( \44082 , \44081 );
not \U$36524 ( \44083 , \43514 );
and \U$36525 ( \44084 , \44082 , \44083 );
nor \U$36526 ( \44085 , \44080 , \44084 );
nand \U$36527 ( \44086 , \44078 , \44085 );
and \U$36528 ( \44087 , \44086 , \44074 );
or \U$36529 ( \44088 , \44076 , \44087 );
and \U$36531 ( \44089 , \44088 , 1'b1 );
or \U$36533 ( \44090 , \44089 , 1'b0 );
buf \U$36534 ( \44091 , \44090 );
_DC r23512_GF_IsGateDCbyConstraint ( \44092_nR23512 , \44091 , \21944 );
buf \U$36535 ( \44093 , \44092_nR23512 );
not \U$36536 ( \44094 , \43568 );
and \U$36537 ( \44095 , RIdc32b68_4933, \44094 );
not \U$36538 ( \44096 , RIdc32b68_4933);
or \U$36539 ( \44097 , \44096 , \43529 );
buf \U$36540 ( \44098 , \22862 );
and \U$36541 ( \44099 , \43405 , \44098 );
buf \U$36542 ( \44100 , RIb832318_202);
buf \U$36543 ( \44101 , \44100 );
not \U$36544 ( \44102 , \43431 );
and \U$36545 ( \44103 , \44101 , \44102 );
nor \U$36546 ( \44104 , \44099 , \44103 );
nand \U$36547 ( \44105 , \44097 , \44104 );
and \U$36548 ( \44106 , \44105 , \43568 );
or \U$36549 ( \44107 , \44095 , \44106 );
and \U$36551 ( \44108 , \44107 , 1'b1 );
or \U$36553 ( \44109 , \44108 , 1'b0 );
buf \U$36554 ( \44110 , \44109 );
_DC r23514_GF_IsGateDCbyConstraint ( \44111_nR23514 , \44110 , \21944 );
buf \U$36555 ( \44112 , \44111_nR23514 );
not \U$36556 ( \44113 , \44018 );
and \U$36557 ( \44114 , RIdc2ee78_4934, \44113 );
not \U$36558 ( \44115 , RIdc2ee78_4934);
or \U$36559 ( \44116 , \44115 , \43425 );
buf \U$36560 ( \44117 , RIb886210_33);
and \U$36561 ( \44118 , \43427 , \44117 );
buf \U$36562 ( \44119 , \33421 );
not \U$36563 ( \44120 , \43556 );
and \U$36564 ( \44121 , \44119 , \44120 );
nor \U$36565 ( \44122 , \44118 , \44121 );
nand \U$36566 ( \44123 , \44116 , \44122 );
and \U$36567 ( \44124 , \44123 , \44018 );
or \U$36568 ( \44125 , \44114 , \44124 );
and \U$36570 ( \44126 , \44125 , 1'b1 );
or \U$36572 ( \44127 , \44126 , 1'b0 );
buf \U$36573 ( \44128 , \44127 );
_DC r23516_GF_IsGateDCbyConstraint ( \44129_nR23516 , \44128 , \21944 );
buf \U$36574 ( \44130 , \44129_nR23516 );
not \U$36575 ( \44131 , \44018 );
and \U$36576 ( \44132 , RIdc29bf8_4935, \44131 );
not \U$36577 ( \44133 , RIdc29bf8_4935);
or \U$36578 ( \44134 , \44133 , \43486 );
buf \U$36579 ( \44135 , RIb886288_32);
buf \U$36580 ( \44136 , \44135 );
and \U$36581 ( \44137 , \43427 , \44136 );
buf \U$36582 ( \44138 , RIb832408_200);
buf \U$36583 ( \44139 , \44138 );
not \U$36584 ( \44140 , \43431 );
and \U$36585 ( \44141 , \44139 , \44140 );
nor \U$36586 ( \44142 , \44137 , \44141 );
nand \U$36587 ( \44143 , \44134 , \44142 );
and \U$36588 ( \44144 , \44143 , \44018 );
or \U$36589 ( \44145 , \44132 , \44144 );
and \U$36591 ( \44146 , \44145 , 1'b1 );
or \U$36593 ( \44147 , \44146 , 1'b0 );
buf \U$36594 ( \44148 , \44147 );
_DC r23518_GF_IsGateDCbyConstraint ( \44149_nR23518 , \44148 , \21944 );
buf \U$36595 ( \44150 , \44149_nR23518 );
not \U$36596 ( \44151 , \43568 );
and \U$36597 ( \44152 , RIddf1628_4936, \44151 );
not \U$36598 ( \44153 , RIddf1628_4936);
or \U$36599 ( \44154 , \44153 , \43655 );
buf \U$36600 ( \44155 , RIb886300_31);
buf \U$36601 ( \44156 , \44155 );
and \U$36602 ( \44157 , \43404 , \44156 );
buf \U$36603 ( \44158 , RIb832480_199);
buf \U$36604 ( \44159 , \44158 );
not \U$36605 ( \44160 , \43601 );
and \U$36606 ( \44161 , \44159 , \44160 );
nor \U$36607 ( \44162 , \44157 , \44161 );
nand \U$36608 ( \44163 , \44154 , \44162 );
and \U$36609 ( \44164 , \44163 , \43568 );
or \U$36610 ( \44165 , \44152 , \44164 );
and \U$36612 ( \44166 , \44165 , 1'b1 );
or \U$36614 ( \44167 , \44166 , 1'b0 );
buf \U$36615 ( \44168 , \44167 );
_DC r2351a_GF_IsGateDCbyConstraint ( \44169_nR2351a , \44168 , \21944 );
buf \U$36616 ( \44170 , \44169_nR2351a );
not \U$36617 ( \44171 , \43961 );
and \U$36618 ( \44172 , RIddee388_4937, \44171 );
not \U$36619 ( \44173 , RIddee388_4937);
or \U$36620 ( \44174 , \44173 , \43529 );
buf \U$36621 ( \44175 , RIb886378_30);
buf \U$36622 ( \44176 , \44175 );
and \U$36623 ( \44177 , \43405 , \44176 );
buf \U$36624 ( \44178 , RIb8324f8_198);
buf \U$36625 ( \44179 , \44178 );
not \U$36626 ( \44180 , \43601 );
and \U$36627 ( \44181 , \44179 , \44180 );
nor \U$36628 ( \44182 , \44177 , \44181 );
nand \U$36629 ( \44183 , \44174 , \44182 );
and \U$36630 ( \44184 , \44183 , \43961 );
or \U$36631 ( \44185 , \44172 , \44184 );
and \U$36633 ( \44186 , \44185 , 1'b1 );
or \U$36635 ( \44187 , \44186 , 1'b0 );
buf \U$36636 ( \44188 , \44187 );
_DC r2351c_GF_IsGateDCbyConstraint ( \44189_nR2351c , \44188 , \21944 );
buf \U$36637 ( \44190 , \44189_nR2351c );
not \U$36638 ( \44191 , \43961 );
and \U$36639 ( \44192 , RIddeaa58_4938, \44191 );
not \U$36640 ( \44193 , RIddeaa58_4938);
or \U$36641 ( \44194 , \44193 , \43465 );
buf \U$36642 ( \44195 , RIb8863f0_29);
buf \U$36643 ( \44196 , \44195 );
and \U$36644 ( \44197 , \43404 , \44196 );
buf \U$36645 ( \44198 , \33496 );
not \U$36646 ( \44199 , \43601 );
and \U$36647 ( \44200 , \44198 , \44199 );
nor \U$36648 ( \44201 , \44197 , \44200 );
nand \U$36649 ( \44202 , \44194 , \44201 );
and \U$36650 ( \44203 , \44202 , \43961 );
or \U$36651 ( \44204 , \44192 , \44203 );
and \U$36653 ( \44205 , \44204 , 1'b1 );
or \U$36655 ( \44206 , \44205 , 1'b0 );
buf \U$36656 ( \44207 , \44206 );
_DC r23520_GF_IsGateDCbyConstraint ( \44208_nR23520 , \44207 , \21944 );
buf \U$36657 ( \44209 , \44208_nR23520 );
not \U$36658 ( \44210 , \43568 );
and \U$36659 ( \44211 , RIdde7a88_4939, \44210 );
not \U$36660 ( \44212 , RIdde7a88_4939);
or \U$36661 ( \44213 , \44212 , \43506 );
buf \U$36662 ( \44214 , \33513 );
and \U$36663 ( \44215 , \43404 , \44214 );
buf \U$36664 ( \44216 , \33516 );
not \U$36665 ( \44217 , \43577 );
and \U$36666 ( \44218 , \44216 , \44217 );
nor \U$36667 ( \44219 , \44215 , \44218 );
nand \U$36668 ( \44220 , \44213 , \44219 );
and \U$36669 ( \44221 , \44220 , \43568 );
or \U$36670 ( \44222 , \44211 , \44221 );
and \U$36672 ( \44223 , \44222 , 1'b1 );
or \U$36674 ( \44224 , \44223 , 1'b0 );
buf \U$36675 ( \44225 , \44224 );
_DC r23522_GF_IsGateDCbyConstraint ( \44226_nR23522 , \44225 , \21944 );
buf \U$36676 ( \44227 , \44226_nR23522 );
not \U$36677 ( \44228 , \43961 );
and \U$36678 ( \44229 , RIdde35a0_4940, \44228 );
not \U$36679 ( \44230 , RIdde35a0_4940);
or \U$36680 ( \44231 , \44230 , \43425 );
buf \U$36681 ( \44232 , \33533 );
and \U$36682 ( \44233 , \43427 , \44232 );
buf \U$36683 ( \44234 , \33536 );
not \U$36684 ( \44235 , \43556 );
and \U$36685 ( \44236 , \44234 , \44235 );
nor \U$36686 ( \44237 , \44233 , \44236 );
nand \U$36687 ( \44238 , \44231 , \44237 );
and \U$36688 ( \44239 , \44238 , \43961 );
or \U$36689 ( \44240 , \44229 , \44239 );
and \U$36691 ( \44241 , \44240 , 1'b1 );
or \U$36693 ( \44242 , \44241 , 1'b0 );
buf \U$36694 ( \44243 , \44242 );
_DC r23524_GF_IsGateDCbyConstraint ( \44244_nR23524 , \44243 , \21944 );
buf \U$36695 ( \44245 , \44244_nR23524 );
not \U$36696 ( \44246 , \44018 );
and \U$36697 ( \44247 , RIdde0cd8_4941, \44246 );
not \U$36698 ( \44248 , RIdde0cd8_4941);
or \U$36699 ( \44249 , \44248 , \43465 );
buf \U$36700 ( \44250 , RIb886558_26);
buf \U$36701 ( \44251 , \44250 );
and \U$36702 ( \44252 , \43405 , \44251 );
buf \U$36703 ( \44253 , \33555 );
not \U$36704 ( \44254 , \43400 );
and \U$36705 ( \44255 , \44253 , \44254 );
nor \U$36706 ( \44256 , \44252 , \44255 );
nand \U$36707 ( \44257 , \44249 , \44256 );
and \U$36708 ( \44258 , \44257 , \44018 );
or \U$36709 ( \44259 , \44247 , \44258 );
and \U$36711 ( \44260 , \44259 , 1'b1 );
or \U$36713 ( \44261 , \44260 , 1'b0 );
buf \U$36714 ( \44262 , \44261 );
_DC r23526_GF_IsGateDCbyConstraint ( \44263_nR23526 , \44262 , \21944 );
buf \U$36715 ( \44264 , \44263_nR23526 );
buf \U$36716 ( \44265 , \43589 );
not \U$36717 ( \44266 , \44265 );
and \U$36718 ( \44267 , RIddddf60_4942, \44266 );
not \U$36719 ( \44268 , RIddddf60_4942);
or \U$36720 ( \44269 , \44268 , \43402 );
buf \U$36721 ( \44270 , RIb8865d0_25);
buf \U$36722 ( \44271 , \44270 );
and \U$36723 ( \44272 , \43405 , \44271 );
buf \U$36724 ( \44273 , RIb838510_193);
buf \U$36725 ( \44274 , \44273 );
not \U$36726 ( \44275 , \43431 );
and \U$36727 ( \44276 , \44274 , \44275 );
nor \U$36728 ( \44277 , \44272 , \44276 );
nand \U$36729 ( \44278 , \44269 , \44277 );
and \U$36730 ( \44279 , \44278 , \44265 );
or \U$36731 ( \44280 , \44267 , \44279 );
and \U$36733 ( \44281 , \44280 , 1'b1 );
or \U$36735 ( \44282 , \44281 , 1'b0 );
buf \U$36736 ( \44283 , \44282 );
_DC r23528_GF_IsGateDCbyConstraint ( \44284_nR23528 , \44283 , \21944 );
buf \U$36737 ( \44285 , \44284_nR23528 );
not \U$36738 ( \44286 , \43961 );
and \U$36739 ( \44287 , RIdddb710_4943, \44286 );
not \U$36740 ( \44288 , RIdddb710_4943);
or \U$36741 ( \44289 , \44288 , \43616 );
buf \U$36742 ( \44290 , RIb886648_24);
buf \U$36743 ( \44291 , \44290 );
and \U$36744 ( \44292 , \43404 , \44291 );
buf \U$36745 ( \44293 , RIb838588_192);
buf \U$36746 ( \44294 , \44293 );
not \U$36747 ( \44295 , \43577 );
and \U$36748 ( \44296 , \44294 , \44295 );
nor \U$36749 ( \44297 , \44292 , \44296 );
nand \U$36750 ( \44298 , \44289 , \44297 );
and \U$36751 ( \44299 , \44298 , \43961 );
or \U$36752 ( \44300 , \44287 , \44299 );
and \U$36754 ( \44301 , \44300 , 1'b1 );
or \U$36756 ( \44302 , \44301 , 1'b0 );
buf \U$36757 ( \44303 , \44302 );
_DC r2352a_GF_IsGateDCbyConstraint ( \44304_nR2352a , \44303 , \21944 );
buf \U$36758 ( \44305 , \44304_nR2352a );
not \U$36759 ( \44306 , \44018 );
and \U$36760 ( \44307 , RIddd5e78_4944, \44306 );
not \U$36761 ( \44308 , RIddd5e78_4944);
or \U$36762 ( \44309 , \44308 , \43465 );
buf \U$36763 ( \44310 , RIb8866c0_23);
buf \U$36764 ( \44311 , \44310 );
and \U$36765 ( \44312 , \43405 , \44311 );
buf \U$36766 ( \44313 , RIb838600_191);
buf \U$36767 ( \44314 , \44313 );
not \U$36768 ( \44315 , \43514 );
and \U$36769 ( \44316 , \44314 , \44315 );
nor \U$36770 ( \44317 , \44312 , \44316 );
nand \U$36771 ( \44318 , \44309 , \44317 );
and \U$36772 ( \44319 , \44318 , \44018 );
or \U$36773 ( \44320 , \44307 , \44319 );
and \U$36775 ( \44321 , \44320 , 1'b1 );
or \U$36777 ( \44322 , \44321 , 1'b0 );
buf \U$36778 ( \44323 , \44322 );
_DC r2352c_GF_IsGateDCbyConstraint ( \44324_nR2352c , \44323 , \21944 );
buf \U$36779 ( \44325 , \44324_nR2352c );
not \U$36780 ( \44326 , \44265 );
and \U$36781 ( \44327 , RIddd2278_4945, \44326 );
not \U$36782 ( \44328 , RIddd2278_4945);
or \U$36783 ( \44329 , \44328 , \43506 );
buf \U$36784 ( \44330 , \33628 );
and \U$36785 ( \44331 , \43405 , \44330 );
buf \U$36786 ( \44332 , \33631 );
not \U$36787 ( \44333 , \43556 );
and \U$36788 ( \44334 , \44332 , \44333 );
nor \U$36789 ( \44335 , \44331 , \44334 );
nand \U$36790 ( \44336 , \44329 , \44335 );
and \U$36791 ( \44337 , \44336 , \44265 );
or \U$36792 ( \44338 , \44327 , \44337 );
and \U$36794 ( \44339 , \44338 , 1'b1 );
or \U$36796 ( \44340 , \44339 , 1'b0 );
buf \U$36797 ( \44341 , \44340 );
_DC r2352e_GF_IsGateDCbyConstraint ( \44342_nR2352e , \44341 , \21944 );
buf \U$36798 ( \44343 , \44342_nR2352e );
not \U$36799 ( \44344 , \44018 );
and \U$36800 ( \44345 , RIddcc080_4946, \44344 );
not \U$36801 ( \44346 , RIddcc080_4946);
or \U$36802 ( \44347 , \44346 , \43425 );
buf \U$36803 ( \44348 , RIb8867b0_21);
buf \U$36804 ( \44349 , \44348 );
and \U$36805 ( \44350 , \43404 , \44349 );
buf \U$36806 ( \44351 , RIb8386f0_189);
buf \U$36807 ( \44352 , \44351 );
not \U$36808 ( \44353 , \43556 );
and \U$36809 ( \44354 , \44352 , \44353 );
nor \U$36810 ( \44355 , \44350 , \44354 );
nand \U$36811 ( \44356 , \44347 , \44355 );
and \U$36812 ( \44357 , \44356 , \44018 );
or \U$36813 ( \44358 , \44345 , \44357 );
and \U$36815 ( \44359 , \44358 , 1'b1 );
or \U$36817 ( \44360 , \44359 , 1'b0 );
buf \U$36818 ( \44361 , \44360 );
_DC r23530_GF_IsGateDCbyConstraint ( \44362_nR23530 , \44361 , \21944 );
buf \U$36819 ( \44363 , \44362_nR23530 );
not \U$36820 ( \44364 , \44074 );
and \U$36821 ( \44365 , RIddc39f8_4947, \44364 );
not \U$36822 ( \44366 , RIddc39f8_4947);
or \U$36823 ( \44367 , \44366 , \43425 );
buf \U$36824 ( \44368 , RIb886828_20);
and \U$36825 ( \44369 , \43427 , \44368 );
buf \U$36826 ( \44370 , \33670 );
not \U$36827 ( \44371 , \43400 );
and \U$36828 ( \44372 , \44370 , \44371 );
nor \U$36829 ( \44373 , \44369 , \44372 );
nand \U$36830 ( \44374 , \44367 , \44373 );
and \U$36831 ( \44375 , \44374 , \44074 );
or \U$36832 ( \44376 , \44365 , \44375 );
and \U$36834 ( \44377 , \44376 , 1'b1 );
or \U$36836 ( \44378 , \44377 , 1'b0 );
buf \U$36837 ( \44379 , \44378 );
_DC r23532_GF_IsGateDCbyConstraint ( \44380_nR23532 , \44379 , \21944 );
buf \U$36838 ( \44381 , \44380_nR23532 );
not \U$36839 ( \44382 , \44265 );
and \U$36840 ( \44383 , RIddbd8f0_4948, \44382 );
not \U$36841 ( \44384 , RIddbd8f0_4948);
or \U$36842 ( \44385 , \44384 , \43655 );
buf \U$36843 ( \44386 , \33687 );
and \U$36844 ( \44387 , \43427 , \44386 );
buf \U$36845 ( \44388 , \33690 );
not \U$36846 ( \44389 , \43577 );
and \U$36847 ( \44390 , \44388 , \44389 );
nor \U$36848 ( \44391 , \44387 , \44390 );
nand \U$36849 ( \44392 , \44385 , \44391 );
and \U$36850 ( \44393 , \44392 , \44265 );
or \U$36851 ( \44394 , \44383 , \44393 );
and \U$36853 ( \44395 , \44394 , 1'b1 );
or \U$36855 ( \44396 , \44395 , 1'b0 );
buf \U$36856 ( \44397 , \44396 );
_DC r23536_GF_IsGateDCbyConstraint ( \44398_nR23536 , \44397 , \21944 );
buf \U$36857 ( \44399 , \44398_nR23536 );
not \U$36858 ( \44400 , \43961 );
and \U$36859 ( \44401 , RIddb5268_4949, \44400 );
not \U$36860 ( \44402 , RIddb5268_4949);
or \U$36861 ( \44403 , \44402 , \43529 );
buf \U$36862 ( \44404 , RIb886918_18);
buf \U$36863 ( \44405 , \44404 );
and \U$36864 ( \44406 , \43405 , \44405 );
buf \U$36865 ( \44407 , \28391 );
not \U$36866 ( \44408 , \43601 );
and \U$36867 ( \44409 , \44407 , \44408 );
nor \U$36868 ( \44410 , \44406 , \44409 );
nand \U$36869 ( \44411 , \44403 , \44410 );
and \U$36870 ( \44412 , \44411 , \43961 );
or \U$36871 ( \44413 , \44401 , \44412 );
and \U$36873 ( \44414 , \44413 , 1'b1 );
or \U$36875 ( \44415 , \44414 , 1'b0 );
buf \U$36876 ( \44416 , \44415 );
_DC r23538_GF_IsGateDCbyConstraint ( \44417_nR23538 , \44416 , \21944 );
buf \U$36877 ( \44418 , \44417_nR23538 );
not \U$36878 ( \44419 , \43961 );
and \U$36879 ( \44420 , RIddaf160_4950, \44419 );
not \U$36880 ( \44421 , RIddaf160_4950);
or \U$36881 ( \44422 , \44421 , \43425 );
buf \U$36882 ( \44423 , RIb886990_17);
and \U$36883 ( \44424 , \43551 , \44423 );
buf \U$36884 ( \44425 , \28411 );
not \U$36885 ( \44426 , \43577 );
and \U$36886 ( \44427 , \44425 , \44426 );
nor \U$36887 ( \44428 , \44424 , \44427 );
nand \U$36888 ( \44429 , \44422 , \44428 );
and \U$36889 ( \44430 , \44429 , \43961 );
or \U$36890 ( \44431 , \44420 , \44430 );
and \U$36892 ( \44432 , \44431 , 1'b1 );
or \U$36894 ( \44433 , \44432 , 1'b0 );
buf \U$36895 ( \44434 , \44433 );
_DC r2353a_GF_IsGateDCbyConstraint ( \44435_nR2353a , \44434 , \21944 );
buf \U$36896 ( \44436 , \44435_nR2353a );
not \U$36897 ( \44437 , \44265 );
and \U$36898 ( \44438 , RIdb7c228_4951, \44437 );
not \U$36899 ( \44439 , RIdb7c228_4951);
or \U$36900 ( \44440 , \44439 , \43465 );
buf \U$36901 ( \44441 , RIb886a08_16);
buf \U$36902 ( \44442 , \44441 );
and \U$36903 ( \44443 , \43405 , \44442 );
buf \U$36904 ( \44444 , RIb838948_184);
buf \U$36905 ( \44445 , \44444 );
not \U$36906 ( \44446 , \43577 );
and \U$36907 ( \44447 , \44445 , \44446 );
nor \U$36908 ( \44448 , \44443 , \44447 );
nand \U$36909 ( \44449 , \44440 , \44448 );
and \U$36910 ( \44450 , \44449 , \44265 );
or \U$36911 ( \44451 , \44438 , \44450 );
and \U$36913 ( \44452 , \44451 , 1'b1 );
or \U$36915 ( \44453 , \44452 , 1'b0 );
buf \U$36916 ( \44454 , \44453 );
_DC r2353c_GF_IsGateDCbyConstraint ( \44455_nR2353c , \44454 , \21944 );
buf \U$36917 ( \44456 , \44455_nR2353c );
not \U$36918 ( \44457 , \44018 );
and \U$36919 ( \44458 , RIdb96c40_4952, \44457 );
not \U$36920 ( \44459 , RIdb96c40_4952);
or \U$36921 ( \44460 , \44459 , \43506 );
buf \U$36922 ( \44461 , \33762 );
and \U$36923 ( \44462 , \43427 , \44461 );
buf \U$36924 ( \44463 , \28451 );
not \U$36925 ( \44464 , \43400 );
and \U$36926 ( \44465 , \44463 , \44464 );
nor \U$36927 ( \44466 , \44462 , \44465 );
nand \U$36928 ( \44467 , \44460 , \44466 );
and \U$36929 ( \44468 , \44467 , \44018 );
or \U$36930 ( \44469 , \44458 , \44468 );
and \U$36932 ( \44470 , \44469 , 1'b1 );
or \U$36934 ( \44471 , \44470 , 1'b0 );
buf \U$36935 ( \44472 , \44471 );
_DC r2353e_GF_IsGateDCbyConstraint ( \44473_nR2353e , \44472 , \21944 );
buf \U$36936 ( \44474 , \44473_nR2353e );
not \U$36937 ( \44475 , \43482 );
and \U$36938 ( \44476 , RIdbbbd38_4953, \44475 );
not \U$36939 ( \44477 , RIdbbbd38_4953);
or \U$36940 ( \44478 , \44477 , \43402 );
buf \U$36941 ( \44479 , \33782 );
and \U$36942 ( \44480 , \43405 , \44479 );
buf \U$36943 ( \44481 , \28470 );
not \U$36944 ( \44482 , \43431 );
and \U$36945 ( \44483 , \44481 , \44482 );
nor \U$36946 ( \44484 , \44480 , \44483 );
nand \U$36947 ( \44485 , \44478 , \44484 );
and \U$36948 ( \44486 , \44485 , \43482 );
or \U$36949 ( \44487 , \44476 , \44486 );
and \U$36951 ( \44488 , \44487 , 1'b1 );
or \U$36953 ( \44489 , \44488 , 1'b0 );
buf \U$36954 ( \44490 , \44489 );
_DC r23540_GF_IsGateDCbyConstraint ( \44491_nR23540 , \44490 , \21944 );
buf \U$36955 ( \44492 , \44491_nR23540 );
not \U$36956 ( \44493 , \44265 );
and \U$36957 ( \44494 , RIdbdcdf8_4954, \44493 );
not \U$36958 ( \44495 , RIdbdcdf8_4954);
or \U$36959 ( \44496 , \44495 , \43616 );
not \U$36960 ( \44497 , \43551 );
not \U$36961 ( \44498 , \44497 );
buf \U$36962 ( \44499 , RIb886b70_13);
buf \U$36963 ( \44500 , \44499 );
and \U$36964 ( \44501 , \44498 , \44500 );
buf \U$36965 ( \44502 , RIb838ab0_181);
buf \U$36966 ( \44503 , \44502 );
not \U$36967 ( \44504 , \43577 );
and \U$36968 ( \44505 , \44503 , \44504 );
nor \U$36969 ( \44506 , \44501 , \44505 );
nand \U$36970 ( \44507 , \44496 , \44506 );
and \U$36971 ( \44508 , \44507 , \44265 );
or \U$36972 ( \44509 , \44494 , \44508 );
and \U$36974 ( \44510 , \44509 , 1'b1 );
or \U$36976 ( \44511 , \44510 , 1'b0 );
buf \U$36977 ( \44512 , \44511 );
_DC r23542_GF_IsGateDCbyConstraint ( \44513_nR23542 , \44512 , \21944 );
buf \U$36978 ( \44514 , \44513_nR23542 );
not \U$36979 ( \44515 , \43961 );
and \U$36980 ( \44516 , RIdb5db80_4955, \44515 );
not \U$36981 ( \44517 , RIdb5db80_4955);
or \U$36982 ( \44518 , \44517 , \43486 );
not \U$36983 ( \44519 , \43551 );
not \U$36984 ( \44520 , \44519 );
buf \U$36985 ( \44521 , \28506 );
and \U$36986 ( \44522 , \44520 , \44521 );
buf \U$36987 ( \44523 , RIb838b28_180);
buf \U$36988 ( \44524 , \44523 );
not \U$36989 ( \44525 , \43577 );
and \U$36990 ( \44526 , \44524 , \44525 );
nor \U$36991 ( \44527 , \44522 , \44526 );
nand \U$36992 ( \44528 , \44518 , \44527 );
and \U$36993 ( \44529 , \44528 , \43961 );
or \U$36994 ( \44530 , \44516 , \44529 );
and \U$36996 ( \44531 , \44530 , 1'b1 );
or \U$36998 ( \44532 , \44531 , 1'b0 );
buf \U$36999 ( \44533 , \44532 );
_DC r23544_GF_IsGateDCbyConstraint ( \44534_nR23544 , \44533 , \21944 );
buf \U$37000 ( \44535 , \44534_nR23544 );
not \U$37001 ( \44536 , \43482 );
and \U$37002 ( \44537 , RIdb48190_4956, \44536 );
not \U$37003 ( \44538 , RIdb48190_4956);
or \U$37004 ( \44539 , \44538 , \43655 );
buf \U$37005 ( \44540 , \39187 );
and \U$37006 ( \44541 , \43427 , \44540 );
buf \U$37007 ( \44542 , RIb838ba0_179);
buf \U$37008 ( \44543 , \44542 );
not \U$37009 ( \44544 , \43514 );
and \U$37010 ( \44545 , \44543 , \44544 );
nor \U$37011 ( \44546 , \44541 , \44545 );
nand \U$37012 ( \44547 , \44539 , \44546 );
and \U$37013 ( \44548 , \44547 , \43482 );
or \U$37014 ( \44549 , \44537 , \44548 );
and \U$37016 ( \44550 , \44549 , 1'b1 );
or \U$37018 ( \44551 , \44550 , 1'b0 );
buf \U$37019 ( \44552 , \44551 );
_DC r23546_GF_IsGateDCbyConstraint ( \44553_nR23546 , \44552 , \21944 );
buf \U$37020 ( \44554 , \44553_nR23546 );
not \U$37021 ( \44555 , \44265 );
and \U$37022 ( \44556 , RIdb26ba8_4957, \44555 );
not \U$37023 ( \44557 , RIdb26ba8_4957);
or \U$37024 ( \44558 , \44557 , \43425 );
buf \U$37025 ( \44559 , \23342 );
and \U$37026 ( \44560 , \43551 , \44559 );
buf \U$37027 ( \44561 , \28550 );
not \U$37028 ( \44562 , \43601 );
and \U$37029 ( \44563 , \44561 , \44562 );
nor \U$37030 ( \44564 , \44560 , \44563 );
nand \U$37031 ( \44565 , \44558 , \44564 );
and \U$37032 ( \44566 , \44565 , \44265 );
or \U$37033 ( \44567 , \44556 , \44566 );
and \U$37035 ( \44568 , \44567 , 1'b1 );
or \U$37037 ( \44569 , \44568 , 1'b0 );
buf \U$37038 ( \44570 , \44569 );
_DC r23548_GF_IsGateDCbyConstraint ( \44571_nR23548 , \44570 , \21944 );
buf \U$37039 ( \44572 , \44571_nR23548 );
not \U$37040 ( \44573 , \43710 );
and \U$37041 ( \44574 , RId917aa8_4958, \44573 );
not \U$37042 ( \44575 , RId917aa8_4958);
or \U$37043 ( \44576 , \44575 , \43402 );
buf \U$37044 ( \44577 , \28568 );
and \U$37045 ( \44578 , \43551 , \44577 );
buf \U$37046 ( \44579 , \23366 );
not \U$37047 ( \44580 , \43556 );
and \U$37048 ( \44581 , \44579 , \44580 );
nor \U$37049 ( \44582 , \44578 , \44581 );
nand \U$37050 ( \44583 , \44576 , \44582 );
and \U$37051 ( \44584 , \44583 , \43710 );
or \U$37052 ( \44585 , \44574 , \44584 );
and \U$37054 ( \44586 , \44585 , 1'b1 );
or \U$37056 ( \44587 , \44586 , 1'b0 );
buf \U$37057 ( \44588 , \44587 );
_DC r2354c_GF_IsGateDCbyConstraint ( \44589_nR2354c , \44588 , \21944 );
buf \U$37058 ( \44590 , \44589_nR2354c );
buf \U$37059 ( \44591 , \43376 );
not \U$37060 ( \44592 , \44591 );
and \U$37061 ( \44593 , RId986da8_4959, \44592 );
not \U$37062 ( \44594 , RId986da8_4959);
or \U$37063 ( \44595 , \44594 , \43616 );
buf \U$37064 ( \44596 , RIb886dc8_8);
and \U$37065 ( \44597 , \43427 , \44596 );
buf \U$37066 ( \44598 , RIb838d08_176);
buf \U$37067 ( \44599 , \44598 );
not \U$37068 ( \44600 , \43431 );
and \U$37069 ( \44601 , \44599 , \44600 );
nor \U$37070 ( \44602 , \44597 , \44601 );
nand \U$37071 ( \44603 , \44595 , \44602 );
and \U$37072 ( \44604 , \44603 , \44591 );
or \U$37073 ( \44605 , \44593 , \44604 );
and \U$37075 ( \44606 , \44605 , 1'b1 );
or \U$37077 ( \44607 , \44606 , 1'b0 );
buf \U$37078 ( \44608 , \44607 );
_DC r2354e_GF_IsGateDCbyConstraint ( \44609_nR2354e , \44608 , \21944 );
buf \U$37079 ( \44610 , \44609_nR2354e );
not \U$37080 ( \44611 , \44265 );
and \U$37081 ( \44612 , RIda7eb60_4960, \44611 );
not \U$37082 ( \44613 , RIda7eb60_4960);
or \U$37083 ( \44614 , \44613 , \43486 );
buf \U$37084 ( \44615 , \28605 );
and \U$37085 ( \44616 , \43427 , \44615 );
buf \U$37086 ( \44617 , RIb838d80_175);
buf \U$37087 ( \44618 , \44617 );
not \U$37088 ( \44619 , \43601 );
and \U$37089 ( \44620 , \44618 , \44619 );
nor \U$37090 ( \44621 , \44616 , \44620 );
nand \U$37091 ( \44622 , \44614 , \44621 );
and \U$37092 ( \44623 , \44622 , \44265 );
or \U$37093 ( \44624 , \44612 , \44623 );
and \U$37095 ( \44625 , \44624 , 1'b1 );
or \U$37097 ( \44626 , \44625 , 1'b0 );
buf \U$37098 ( \44627 , \44626 );
_DC r23550_GF_IsGateDCbyConstraint ( \44628_nR23550 , \44627 , \21944 );
buf \U$37099 ( \44629 , \44628_nR23550 );
not \U$37100 ( \44630 , \43961 );
and \U$37101 ( \44631 , RIdaf90e0_4961, \44630 );
not \U$37102 ( \44632 , RIdaf90e0_4961);
or \U$37103 ( \44633 , \44632 , \43655 );
buf \U$37104 ( \44634 , \23423 );
and \U$37105 ( \44635 , \43405 , \44634 );
buf \U$37106 ( \44636 , \23426 );
not \U$37107 ( \44637 , \43601 );
and \U$37108 ( \44638 , \44636 , \44637 );
nor \U$37109 ( \44639 , \44635 , \44638 );
nand \U$37110 ( \44640 , \44633 , \44639 );
and \U$37111 ( \44641 , \44640 , \43961 );
or \U$37112 ( \44642 , \44631 , \44641 );
and \U$37114 ( \44643 , \44642 , 1'b1 );
or \U$37116 ( \44644 , \44643 , 1'b0 );
buf \U$37117 ( \44645 , \44644 );
_DC r23552_GF_IsGateDCbyConstraint ( \44646_nR23552 , \44645 , \21944 );
buf \U$37118 ( \44647 , \44646_nR23552 );
not \U$37119 ( \44648 , \43961 );
and \U$37120 ( \44649 , RIdab27a8_4962, \44648 );
not \U$37121 ( \44650 , RIdab27a8_4962);
not \U$37122 ( \44651 , \43395 );
nor \U$37123 ( \44652 , \43392 , \44651 );
nand \U$37124 ( \44653 , \44652 , \43397 );
not \U$37125 ( \44654 , \44653 );
not \U$37126 ( \44655 , \43383 );
or \U$37127 ( \44656 , \43385 , \44655 );
not \U$37128 ( \44657 , \44656 );
nand \U$37129 ( \44658 , \43374 , \44657 );
not \U$37130 ( \44659 , \44658 );
or \U$37131 ( \44660 , \44654 , \44659 );
not \U$37132 ( \44661 , \44660 );
not \U$37133 ( \44662 , \44661 );
or \U$37134 ( \44663 , \44650 , \44662 );
not \U$37135 ( \44664 , \44653 );
not \U$37136 ( \44665 , \44664 );
not \U$37137 ( \44666 , \44665 );
and \U$37138 ( \44667 , \43409 , \44666 );
not \U$37139 ( \44668 , \44667 );
not \U$37140 ( \44669 , \43407 );
not \U$37141 ( \44670 , \44658 );
buf \U$37142 ( \44671 , \44670 );
not \U$37143 ( \44672 , \44671 );
or \U$37144 ( \44673 , \44669 , \44672 );
nand \U$37145 ( \44674 , \44663 , \44668 , \44673 );
and \U$37146 ( \44675 , \44674 , \43961 );
or \U$37147 ( \44676 , \44649 , \44675 );
and \U$37149 ( \44677 , \44676 , 1'b1 );
or \U$37151 ( \44678 , \44677 , 1'b0 );
buf \U$37152 ( \44679 , \44678 );
_DC r2355c_GF_IsGateDCbyConstraint ( \44680_nR2355c , \44679 , \21944 );
buf \U$37153 ( \44681 , \44680_nR2355c );
not \U$37154 ( \44682 , \44265 );
and \U$37155 ( \44683 , RIdbf1ca8_4963, \44682 );
not \U$37156 ( \44684 , RIdbf1ca8_4963);
or \U$37157 ( \44685 , \44684 , \44662 );
not \U$37158 ( \44686 , \44654 );
not \U$37159 ( \44687 , \44686 );
and \U$37160 ( \44688 , \43430 , \44687 );
not \U$37161 ( \44689 , \44688 );
not \U$37162 ( \44690 , \43428 );
buf \U$37163 ( \44691 , \44670 );
not \U$37164 ( \44692 , \44691 );
or \U$37165 ( \44693 , \44690 , \44692 );
nand \U$37166 ( \44694 , \44685 , \44689 , \44693 );
and \U$37167 ( \44695 , \44694 , \44265 );
or \U$37168 ( \44696 , \44683 , \44695 );
and \U$37170 ( \44697 , \44696 , 1'b1 );
or \U$37172 ( \44698 , \44697 , 1'b0 );
buf \U$37173 ( \44699 , \44698 );
_DC r23572_GF_IsGateDCbyConstraint ( \44700_nR23572 , \44699 , \21944 );
buf \U$37174 ( \44701 , \44700_nR23572 );
not \U$37175 ( \44702 , \43961 );
and \U$37176 ( \44703 , RIdc00a50_4964, \44702 );
not \U$37177 ( \44704 , RIdc00a50_4964);
not \U$37178 ( \44705 , \44661 );
or \U$37179 ( \44706 , \44704 , \44705 );
not \U$37180 ( \44707 , \44665 );
and \U$37181 ( \44708 , \43450 , \44707 );
not \U$37182 ( \44709 , \44708 );
not \U$37183 ( \44710 , \43448 );
not \U$37184 ( \44711 , \44671 );
or \U$37185 ( \44712 , \44710 , \44711 );
nand \U$37186 ( \44713 , \44706 , \44709 , \44712 );
and \U$37187 ( \44714 , \44713 , \43961 );
or \U$37188 ( \44715 , \44703 , \44714 );
and \U$37190 ( \44716 , \44715 , 1'b1 );
or \U$37192 ( \44717 , \44716 , 1'b0 );
buf \U$37193 ( \44718 , \44717 );
_DC r23588_GF_IsGateDCbyConstraint ( \44719_nR23588 , \44718 , \21944 );
buf \U$37194 ( \44720 , \44719_nR23588 );
not \U$37195 ( \44721 , \44018 );
and \U$37196 ( \44722 , RIdc0fe88_4965, \44721 );
not \U$37197 ( \44723 , RIdc0fe88_4965);
not \U$37198 ( \44724 , \44661 );
or \U$37199 ( \44725 , \44723 , \44724 );
not \U$37200 ( \44726 , \44686 );
and \U$37201 ( \44727 , \43470 , \44726 );
not \U$37202 ( \44728 , \44727 );
not \U$37203 ( \44729 , \43468 );
not \U$37204 ( \44730 , \44671 );
or \U$37205 ( \44731 , \44729 , \44730 );
nand \U$37206 ( \44732 , \44725 , \44728 , \44731 );
and \U$37207 ( \44733 , \44732 , \44018 );
or \U$37208 ( \44734 , \44722 , \44733 );
and \U$37210 ( \44735 , \44734 , 1'b1 );
or \U$37212 ( \44736 , \44735 , 1'b0 );
buf \U$37213 ( \44737 , \44736 );
_DC r2359e_GF_IsGateDCbyConstraint ( \44738_nR2359e , \44737 , \21944 );
buf \U$37214 ( \44739 , \44738_nR2359e );
not \U$37215 ( \44740 , \44265 );
and \U$37216 ( \44741 , RIdc16080_4966, \44740 );
not \U$37217 ( \44742 , RIdc16080_4966);
or \U$37218 ( \44743 , \44742 , \44705 );
not \U$37219 ( \44744 , \44665 );
and \U$37220 ( \44745 , \43491 , \44744 );
not \U$37221 ( \44746 , \44745 );
not \U$37222 ( \44747 , \43488 );
not \U$37223 ( \44748 , \44691 );
or \U$37224 ( \44749 , \44747 , \44748 );
nand \U$37225 ( \44750 , \44743 , \44746 , \44749 );
and \U$37226 ( \44751 , \44750 , \44265 );
or \U$37227 ( \44752 , \44741 , \44751 );
and \U$37229 ( \44753 , \44752 , 1'b1 );
or \U$37231 ( \44754 , \44753 , 1'b0 );
buf \U$37232 ( \44755 , \44754 );
_DC r235b4_GF_IsGateDCbyConstraint ( \44756_nR235b4 , \44755 , \21944 );
buf \U$37233 ( \44757 , \44756_nR235b4 );
buf \U$37234 ( \44758 , \43482 );
not \U$37235 ( \44759 , \44758 );
and \U$37236 ( \44760 , RIdc1c098_4967, \44759 );
not \U$37237 ( \44761 , RIdc1c098_4967);
or \U$37238 ( \44762 , \44761 , \44705 );
not \U$37239 ( \44763 , \44654 );
not \U$37240 ( \44764 , \44763 );
and \U$37241 ( \44765 , \43510 , \44764 );
not \U$37242 ( \44766 , \44765 );
not \U$37243 ( \44767 , \43508 );
buf \U$37244 ( \44768 , \44670 );
not \U$37245 ( \44769 , \44768 );
or \U$37246 ( \44770 , \44767 , \44769 );
nand \U$37247 ( \44771 , \44762 , \44766 , \44770 );
and \U$37248 ( \44772 , \44771 , \44758 );
or \U$37249 ( \44773 , \44760 , \44772 );
and \U$37251 ( \44774 , \44773 , 1'b1 );
or \U$37253 ( \44775 , \44774 , 1'b0 );
buf \U$37254 ( \44776 , \44775 );
_DC r235ca_GF_IsGateDCbyConstraint ( \44777_nR235ca , \44776 , \21944 );
buf \U$37255 ( \44778 , \44777_nR235ca );
not \U$37256 ( \44779 , \44758 );
and \U$37257 ( \44780 , RIdc25080_4968, \44779 );
not \U$37258 ( \44781 , RIdc25080_4968);
or \U$37259 ( \44782 , \44781 , \44662 );
not \U$37260 ( \44783 , \44664 );
not \U$37261 ( \44784 , \44783 );
and \U$37262 ( \44785 , \43535 , \44784 );
not \U$37263 ( \44786 , \44785 );
not \U$37264 ( \44787 , \43532 );
not \U$37265 ( \44788 , \44691 );
or \U$37266 ( \44789 , \44787 , \44788 );
nand \U$37267 ( \44790 , \44782 , \44786 , \44789 );
and \U$37268 ( \44791 , \44790 , \44758 );
or \U$37269 ( \44792 , \44780 , \44791 );
and \U$37271 ( \44793 , \44792 , 1'b1 );
or \U$37273 ( \44794 , \44793 , 1'b0 );
buf \U$37274 ( \44795 , \44794 );
_DC r235d4_GF_IsGateDCbyConstraint ( \44796_nR235d4 , \44795 , \21944 );
buf \U$37275 ( \44797 , \44796_nR235d4 );
not \U$37276 ( \44798 , \44265 );
and \U$37277 ( \44799 , RIdb67810_4969, \44798 );
not \U$37278 ( \44800 , RIdb67810_4969);
not \U$37279 ( \44801 , \44661 );
or \U$37280 ( \44802 , \44800 , \44801 );
not \U$37281 ( \44803 , \44686 );
and \U$37282 ( \44804 , \43555 , \44803 );
not \U$37283 ( \44805 , \44804 );
not \U$37284 ( \44806 , \43553 );
not \U$37285 ( \44807 , \44768 );
or \U$37286 ( \44808 , \44806 , \44807 );
nand \U$37287 ( \44809 , \44802 , \44805 , \44808 );
and \U$37288 ( \44810 , \44809 , \44265 );
or \U$37289 ( \44811 , \44799 , \44810 );
and \U$37291 ( \44812 , \44811 , 1'b1 );
or \U$37293 ( \44813 , \44812 , 1'b0 );
buf \U$37294 ( \44814 , \44813 );
_DC r235d6_GF_IsGateDCbyConstraint ( \44815_nR235d6 , \44814 , \21944 );
buf \U$37295 ( \44816 , \44815_nR235d6 );
not \U$37296 ( \44817 , \43377 );
and \U$37297 ( \44818 , RIdda8518_4970, \44817 );
not \U$37298 ( \44819 , RIdda8518_4970);
or \U$37299 ( \44820 , \44819 , \44662 );
not \U$37300 ( \44821 , \44763 );
and \U$37301 ( \44822 , \43576 , \44821 );
not \U$37302 ( \44823 , \44822 );
not \U$37303 ( \44824 , \43573 );
not \U$37304 ( \44825 , \44768 );
or \U$37305 ( \44826 , \44824 , \44825 );
nand \U$37306 ( \44827 , \44820 , \44823 , \44826 );
and \U$37307 ( \44828 , \44827 , \43377 );
or \U$37308 ( \44829 , \44818 , \44828 );
and \U$37310 ( \44830 , \44829 , 1'b1 );
or \U$37312 ( \44831 , \44830 , 1'b0 );
buf \U$37313 ( \44832 , \44831 );
_DC r235d8_GF_IsGateDCbyConstraint ( \44833_nR235d8 , \44832 , \21944 );
buf \U$37314 ( \44834 , \44833_nR235d8 );
not \U$37315 ( \44835 , \43589 );
and \U$37316 ( \44836 , RIdd9d5c8_4971, \44835 );
not \U$37317 ( \44837 , RIdd9d5c8_4971);
or \U$37318 ( \44838 , \44837 , \44705 );
not \U$37319 ( \44839 , \44664 );
not \U$37320 ( \44840 , \44839 );
and \U$37321 ( \44841 , \43597 , \44840 );
not \U$37322 ( \44842 , \44841 );
not \U$37323 ( \44843 , \43595 );
not \U$37324 ( \44844 , \44671 );
or \U$37325 ( \44845 , \44843 , \44844 );
nand \U$37326 ( \44846 , \44838 , \44842 , \44845 );
and \U$37327 ( \44847 , \44846 , \43589 );
or \U$37328 ( \44848 , \44836 , \44847 );
and \U$37330 ( \44849 , \44848 , 1'b1 );
or \U$37332 ( \44850 , \44849 , 1'b0 );
buf \U$37333 ( \44851 , \44850 );
_DC r235da_GF_IsGateDCbyConstraint ( \44852_nR235da , \44851 , \21944 );
buf \U$37334 ( \44853 , \44852_nR235da );
not \U$37335 ( \44854 , \44265 );
and \U$37336 ( \44855 , RIdd8f270_4972, \44854 );
not \U$37337 ( \44856 , RIdd8f270_4972);
or \U$37338 ( \44857 , \44856 , \44801 );
not \U$37339 ( \44858 , \44839 );
and \U$37340 ( \44859 , \43622 , \44858 );
not \U$37341 ( \44860 , \44859 );
not \U$37342 ( \44861 , \43619 );
not \U$37343 ( \44862 , \44768 );
or \U$37344 ( \44863 , \44861 , \44862 );
nand \U$37345 ( \44864 , \44857 , \44860 , \44863 );
and \U$37346 ( \44865 , \44864 , \44265 );
or \U$37347 ( \44866 , \44855 , \44865 );
and \U$37349 ( \44867 , \44866 , 1'b1 );
or \U$37351 ( \44868 , \44867 , 1'b0 );
buf \U$37352 ( \44869 , \44868 );
_DC r2355e_GF_IsGateDCbyConstraint ( \44870_nR2355e , \44869 , \21944 );
buf \U$37353 ( \44871 , \44870_nR2355e );
not \U$37354 ( \44872 , \44758 );
and \U$37355 ( \44873 , RIdd82fe8_4973, \44872 );
not \U$37356 ( \44874 , RIdd82fe8_4973);
or \U$37357 ( \44875 , \44874 , \44662 );
not \U$37358 ( \44876 , \44664 );
not \U$37359 ( \44877 , \44876 );
and \U$37360 ( \44878 , \43640 , \44877 );
not \U$37361 ( \44879 , \44878 );
not \U$37362 ( \44880 , \43638 );
not \U$37363 ( \44881 , \44671 );
or \U$37364 ( \44882 , \44880 , \44881 );
nand \U$37365 ( \44883 , \44875 , \44879 , \44882 );
and \U$37366 ( \44884 , \44883 , \44758 );
or \U$37367 ( \44885 , \44873 , \44884 );
and \U$37369 ( \44886 , \44885 , 1'b1 );
or \U$37371 ( \44887 , \44886 , 1'b0 );
buf \U$37372 ( \44888 , \44887 );
_DC r23560_GF_IsGateDCbyConstraint ( \44889_nR23560 , \44888 , \21944 );
buf \U$37373 ( \44890 , \44889_nR23560 );
not \U$37374 ( \44891 , \44758 );
and \U$37375 ( \44892 , RIdd74150_4974, \44891 );
not \U$37376 ( \44893 , RIdd74150_4974);
or \U$37377 ( \44894 , \44893 , \44801 );
not \U$37378 ( \44895 , \44664 );
not \U$37379 ( \44896 , \44895 );
and \U$37380 ( \44897 , \43661 , \44896 );
not \U$37381 ( \44898 , \44897 );
not \U$37382 ( \44899 , \43658 );
not \U$37383 ( \44900 , \44768 );
or \U$37384 ( \44901 , \44899 , \44900 );
nand \U$37385 ( \44902 , \44894 , \44898 , \44901 );
and \U$37386 ( \44903 , \44902 , \44758 );
or \U$37387 ( \44904 , \44892 , \44903 );
and \U$37389 ( \44905 , \44904 , 1'b1 );
or \U$37391 ( \44906 , \44905 , 1'b0 );
buf \U$37392 ( \44907 , \44906 );
_DC r23562_GF_IsGateDCbyConstraint ( \44908_nR23562 , \44907 , \21944 );
buf \U$37393 ( \44909 , \44908_nR23562 );
not \U$37394 ( \44910 , \44265 );
and \U$37395 ( \44911 , RIdc641b8_4975, \44910 );
not \U$37396 ( \44912 , RIdc641b8_4975);
or \U$37397 ( \44913 , \44912 , \44662 );
not \U$37398 ( \44914 , \44665 );
and \U$37399 ( \44915 , \43680 , \44914 );
not \U$37400 ( \44916 , \44915 );
not \U$37401 ( \44917 , \43678 );
not \U$37402 ( \44918 , \44670 );
or \U$37403 ( \44919 , \44917 , \44918 );
nand \U$37404 ( \44920 , \44913 , \44916 , \44919 );
and \U$37405 ( \44921 , \44920 , \44265 );
or \U$37406 ( \44922 , \44911 , \44921 );
and \U$37408 ( \44923 , \44922 , 1'b1 );
or \U$37410 ( \44924 , \44923 , 1'b0 );
buf \U$37411 ( \44925 , \44924 );
_DC r23564_GF_IsGateDCbyConstraint ( \44926_nR23564 , \44925 , \21944 );
buf \U$37412 ( \44927 , \44926_nR23564 );
not \U$37413 ( \44928 , \44758 );
and \U$37414 ( \44929 , RIdc54600_4976, \44928 );
not \U$37415 ( \44930 , RIdc54600_4976);
or \U$37416 ( \44931 , \44930 , \44705 );
not \U$37417 ( \44932 , \44839 );
and \U$37418 ( \44933 , \43698 , \44932 );
not \U$37419 ( \44934 , \44933 );
not \U$37420 ( \44935 , \43696 );
not \U$37421 ( \44936 , \44768 );
or \U$37422 ( \44937 , \44935 , \44936 );
nand \U$37423 ( \44938 , \44931 , \44934 , \44937 );
and \U$37424 ( \44939 , \44938 , \44758 );
or \U$37425 ( \44940 , \44929 , \44939 );
and \U$37427 ( \44941 , \44940 , 1'b1 );
or \U$37429 ( \44942 , \44941 , 1'b0 );
buf \U$37430 ( \44943 , \44942 );
_DC r23566_GF_IsGateDCbyConstraint ( \44944_nR23566 , \44943 , \21944 );
buf \U$37431 ( \44945 , \44944_nR23566 );
not \U$37432 ( \44946 , \43710 );
and \U$37433 ( \44947 , RIdc46848_4977, \44946 );
not \U$37434 ( \44948 , RIdc46848_4977);
or \U$37435 ( \44949 , \44948 , \44724 );
not \U$37436 ( \44950 , \44876 );
and \U$37437 ( \44951 , \43718 , \44950 );
not \U$37438 ( \44952 , \44951 );
not \U$37439 ( \44953 , \43715 );
not \U$37440 ( \44954 , \44691 );
or \U$37441 ( \44955 , \44953 , \44954 );
nand \U$37442 ( \44956 , \44949 , \44952 , \44955 );
and \U$37443 ( \44957 , \44956 , \43710 );
or \U$37444 ( \44958 , \44947 , \44957 );
and \U$37446 ( \44959 , \44958 , 1'b1 );
or \U$37448 ( \44960 , \44959 , 1'b0 );
buf \U$37449 ( \44961 , \44960 );
_DC r23568_GF_IsGateDCbyConstraint ( \44962_nR23568 , \44961 , \21944 );
buf \U$37450 ( \44963 , \44962_nR23568 );
not \U$37451 ( \44964 , \43961 );
and \U$37452 ( \44965 , RIdc3b970_4978, \44964 );
not \U$37453 ( \44966 , RIdc3b970_4978);
or \U$37454 ( \44967 , \44966 , \44705 );
not \U$37455 ( \44968 , \44895 );
and \U$37456 ( \44969 , \43738 , \44968 );
not \U$37457 ( \44970 , \44969 );
not \U$37458 ( \44971 , \43736 );
not \U$37459 ( \44972 , \44768 );
or \U$37460 ( \44973 , \44971 , \44972 );
nand \U$37461 ( \44974 , \44967 , \44970 , \44973 );
and \U$37462 ( \44975 , \44974 , \43961 );
or \U$37463 ( \44976 , \44965 , \44975 );
and \U$37465 ( \44977 , \44976 , 1'b1 );
or \U$37467 ( \44978 , \44977 , 1'b0 );
buf \U$37468 ( \44979 , \44978 );
_DC r2356a_GF_IsGateDCbyConstraint ( \44980_nR2356a , \44979 , \21944 );
buf \U$37469 ( \44981 , \44980_nR2356a );
not \U$37470 ( \44982 , \44758 );
and \U$37471 ( \44983 , RIdf77220_4979, \44982 );
not \U$37472 ( \44984 , RIdf77220_4979);
or \U$37473 ( \44985 , \44984 , \44705 );
not \U$37474 ( \44986 , \44783 );
and \U$37475 ( \44987 , \43756 , \44986 );
not \U$37476 ( \44988 , \44987 );
not \U$37477 ( \44989 , \43754 );
not \U$37478 ( \44990 , \44691 );
or \U$37479 ( \44991 , \44989 , \44990 );
nand \U$37480 ( \44992 , \44985 , \44988 , \44991 );
and \U$37481 ( \44993 , \44992 , \44758 );
or \U$37482 ( \44994 , \44983 , \44993 );
and \U$37484 ( \44995 , \44994 , 1'b1 );
or \U$37486 ( \44996 , \44995 , 1'b0 );
buf \U$37487 ( \44997 , \44996 );
_DC r2356c_GF_IsGateDCbyConstraint ( \44998_nR2356c , \44997 , \21944 );
buf \U$37488 ( \44999 , \44998_nR2356c );
not \U$37489 ( \45000 , \44591 );
and \U$37490 ( \45001 , RIdf79f98_4980, \45000 );
not \U$37491 ( \45002 , RIdf79f98_4980);
or \U$37492 ( \45003 , \45002 , \44724 );
not \U$37493 ( \45004 , \44876 );
and \U$37494 ( \45005 , \43776 , \45004 );
not \U$37495 ( \45006 , \45005 );
not \U$37496 ( \45007 , \43773 );
not \U$37497 ( \45008 , \44691 );
or \U$37498 ( \45009 , \45007 , \45008 );
nand \U$37499 ( \45010 , \45003 , \45006 , \45009 );
and \U$37500 ( \45011 , \45010 , \44591 );
or \U$37501 ( \45012 , \45001 , \45011 );
and \U$37503 ( \45013 , \45012 , 1'b1 );
or \U$37505 ( \45014 , \45013 , 1'b0 );
buf \U$37506 ( \45015 , \45014 );
_DC r2356e_GF_IsGateDCbyConstraint ( \45016_nR2356e , \45015 , \21944 );
buf \U$37507 ( \45017 , \45016_nR2356e );
not \U$37508 ( \45018 , \43710 );
and \U$37509 ( \45019 , RIdf7c860_4981, \45018 );
not \U$37510 ( \45020 , RIdf7c860_4981);
or \U$37511 ( \45021 , \45020 , \44662 );
not \U$37512 ( \45022 , \44783 );
and \U$37513 ( \45023 , \43795 , \45022 );
not \U$37514 ( \45024 , \45023 );
not \U$37515 ( \45025 , \43792 );
not \U$37516 ( \45026 , \44671 );
or \U$37517 ( \45027 , \45025 , \45026 );
nand \U$37518 ( \45028 , \45021 , \45024 , \45027 );
and \U$37519 ( \45029 , \45028 , \43710 );
or \U$37520 ( \45030 , \45019 , \45029 );
and \U$37522 ( \45031 , \45030 , 1'b1 );
or \U$37524 ( \45032 , \45031 , 1'b0 );
buf \U$37525 ( \45033 , \45032 );
_DC r23570_GF_IsGateDCbyConstraint ( \45034_nR23570 , \45033 , \21944 );
buf \U$37526 ( \45035 , \45034_nR23570 );
not \U$37527 ( \45036 , \44074 );
and \U$37528 ( \45037 , RIdf7ff38_4982, \45036 );
not \U$37529 ( \45038 , RIdf7ff38_4982);
or \U$37530 ( \45039 , \45038 , \44724 );
not \U$37531 ( \45040 , \44763 );
and \U$37532 ( \45041 , \43813 , \45040 );
not \U$37533 ( \45042 , \45041 );
not \U$37534 ( \45043 , \43811 );
not \U$37535 ( \45044 , \44768 );
or \U$37536 ( \45045 , \45043 , \45044 );
nand \U$37537 ( \45046 , \45039 , \45042 , \45045 );
and \U$37538 ( \45047 , \45046 , \44074 );
or \U$37539 ( \45048 , \45037 , \45047 );
and \U$37541 ( \45049 , \45048 , 1'b1 );
or \U$37543 ( \45050 , \45049 , 1'b0 );
buf \U$37544 ( \45051 , \45050 );
_DC r23574_GF_IsGateDCbyConstraint ( \45052_nR23574 , \45051 , \21944 );
buf \U$37545 ( \45053 , \45052_nR23574 );
not \U$37546 ( \45054 , \43730 );
and \U$37547 ( \45055 , RIdf82800_4983, \45054 );
not \U$37548 ( \45056 , RIdf82800_4983);
or \U$37549 ( \45057 , \45056 , \44724 );
not \U$37550 ( \45058 , \44839 );
and \U$37551 ( \45059 , \43832 , \45058 );
not \U$37552 ( \45060 , \45059 );
not \U$37553 ( \45061 , \43830 );
not \U$37554 ( \45062 , \44671 );
or \U$37555 ( \45063 , \45061 , \45062 );
nand \U$37556 ( \45064 , \45057 , \45060 , \45063 );
and \U$37557 ( \45065 , \45064 , \43730 );
or \U$37558 ( \45066 , \45055 , \45065 );
and \U$37560 ( \45067 , \45066 , 1'b1 );
or \U$37562 ( \45068 , \45067 , 1'b0 );
buf \U$37563 ( \45069 , \45068 );
_DC r23576_GF_IsGateDCbyConstraint ( \45070_nR23576 , \45069 , \21944 );
buf \U$37564 ( \45071 , \45070_nR23576 );
not \U$37565 ( \45072 , \44074 );
and \U$37566 ( \45073 , RIdf85ed8_4984, \45072 );
not \U$37567 ( \45074 , RIdf85ed8_4984);
or \U$37568 ( \45075 , \45074 , \44705 );
not \U$37569 ( \45076 , \44686 );
and \U$37570 ( \45077 , \43852 , \45076 );
not \U$37571 ( \45078 , \45077 );
not \U$37572 ( \45079 , \43849 );
not \U$37573 ( \45080 , \44670 );
or \U$37574 ( \45081 , \45079 , \45080 );
nand \U$37575 ( \45082 , \45075 , \45078 , \45081 );
and \U$37576 ( \45083 , \45082 , \44074 );
or \U$37577 ( \45084 , \45073 , \45083 );
and \U$37579 ( \45085 , \45084 , 1'b1 );
or \U$37581 ( \45086 , \45085 , 1'b0 );
buf \U$37582 ( \45087 , \45086 );
_DC r23578_GF_IsGateDCbyConstraint ( \45088_nR23578 , \45087 , \21944 );
buf \U$37583 ( \45089 , \45088_nR23578 );
not \U$37584 ( \45090 , \44758 );
and \U$37585 ( \45091 , RIdf887a0_4985, \45090 );
not \U$37586 ( \45092 , RIdf887a0_4985);
or \U$37587 ( \45093 , \45092 , \44662 );
not \U$37588 ( \45094 , \44763 );
and \U$37589 ( \45095 , \43872 , \45094 );
not \U$37590 ( \45096 , \45095 );
not \U$37591 ( \45097 , \43869 );
not \U$37592 ( \45098 , \44768 );
or \U$37593 ( \45099 , \45097 , \45098 );
nand \U$37594 ( \45100 , \45093 , \45096 , \45099 );
and \U$37595 ( \45101 , \45100 , \44758 );
or \U$37596 ( \45102 , \45091 , \45101 );
and \U$37598 ( \45103 , \45102 , 1'b1 );
or \U$37600 ( \45104 , \45103 , 1'b0 );
buf \U$37601 ( \45105 , \45104 );
_DC r2357a_GF_IsGateDCbyConstraint ( \45106_nR2357a , \45105 , \21944 );
buf \U$37602 ( \45107 , \45106_nR2357a );
not \U$37603 ( \45108 , \44758 );
and \U$37604 ( \45109 , RIdf8be78_4986, \45108 );
not \U$37605 ( \45110 , RIdf8be78_4986);
or \U$37606 ( \45111 , \45110 , \44662 );
not \U$37607 ( \45112 , \44839 );
and \U$37608 ( \45113 , \43890 , \45112 );
not \U$37609 ( \45114 , \45113 );
not \U$37610 ( \45115 , \43888 );
not \U$37611 ( \45116 , \44670 );
or \U$37612 ( \45117 , \45115 , \45116 );
nand \U$37613 ( \45118 , \45111 , \45114 , \45117 );
and \U$37614 ( \45119 , \45118 , \44758 );
or \U$37615 ( \45120 , \45109 , \45119 );
and \U$37617 ( \45121 , \45120 , 1'b1 );
or \U$37619 ( \45122 , \45121 , 1'b0 );
buf \U$37620 ( \45123 , \45122 );
_DC r2357c_GF_IsGateDCbyConstraint ( \45124_nR2357c , \45123 , \21944 );
buf \U$37621 ( \45125 , \45124_nR2357c );
not \U$37622 ( \45126 , \43377 );
and \U$37623 ( \45127 , RIdf8e740_4987, \45126 );
not \U$37624 ( \45128 , RIdf8e740_4987);
or \U$37625 ( \45129 , \45128 , \44801 );
not \U$37626 ( \45130 , \44665 );
and \U$37627 ( \45131 , \43910 , \45130 );
not \U$37628 ( \45132 , \45131 );
not \U$37629 ( \45133 , \43907 );
not \U$37630 ( \45134 , \44691 );
or \U$37631 ( \45135 , \45133 , \45134 );
nand \U$37632 ( \45136 , \45129 , \45132 , \45135 );
and \U$37633 ( \45137 , \45136 , \43377 );
or \U$37634 ( \45138 , \45127 , \45137 );
and \U$37636 ( \45139 , \45138 , 1'b1 );
or \U$37638 ( \45140 , \45139 , 1'b0 );
buf \U$37639 ( \45141 , \45140 );
_DC r2357e_GF_IsGateDCbyConstraint ( \45142_nR2357e , \45141 , \21944 );
buf \U$37640 ( \45143 , \45142_nR2357e );
not \U$37641 ( \45144 , \44758 );
and \U$37642 ( \45145 , RIdf91008_4988, \45144 );
not \U$37643 ( \45146 , RIdf91008_4988);
or \U$37644 ( \45147 , \45146 , \44662 );
not \U$37645 ( \45148 , \44763 );
and \U$37646 ( \45149 , \43929 , \45148 );
not \U$37647 ( \45150 , \45149 );
not \U$37648 ( \45151 , \43927 );
not \U$37649 ( \45152 , \44671 );
or \U$37650 ( \45153 , \45151 , \45152 );
nand \U$37651 ( \45154 , \45147 , \45150 , \45153 );
and \U$37652 ( \45155 , \45154 , \44758 );
or \U$37653 ( \45156 , \45145 , \45155 );
and \U$37655 ( \45157 , \45156 , 1'b1 );
or \U$37657 ( \45158 , \45157 , 1'b0 );
buf \U$37658 ( \45159 , \45158 );
_DC r23580_GF_IsGateDCbyConstraint ( \45160_nR23580 , \45159 , \21944 );
buf \U$37659 ( \45161 , \45160_nR23580 );
not \U$37660 ( \45162 , \43482 );
and \U$37661 ( \45163 , RIdf946e0_4989, \45162 );
not \U$37662 ( \45164 , RIdf946e0_4989);
or \U$37663 ( \45165 , \45164 , \44705 );
not \U$37664 ( \45166 , \44686 );
and \U$37665 ( \45167 , \43949 , \45166 );
not \U$37666 ( \45168 , \45167 );
not \U$37667 ( \45169 , \43946 );
not \U$37668 ( \45170 , \44671 );
or \U$37669 ( \45171 , \45169 , \45170 );
nand \U$37670 ( \45172 , \45165 , \45168 , \45171 );
and \U$37671 ( \45173 , \45172 , \43482 );
or \U$37672 ( \45174 , \45163 , \45173 );
and \U$37674 ( \45175 , \45174 , 1'b1 );
or \U$37676 ( \45176 , \45175 , 1'b0 );
buf \U$37677 ( \45177 , \45176 );
_DC r23582_GF_IsGateDCbyConstraint ( \45178_nR23582 , \45177 , \21944 );
buf \U$37678 ( \45179 , \45178_nR23582 );
not \U$37679 ( \45180 , \43589 );
and \U$37680 ( \45181 , RIdf96fa8_4990, \45180 );
not \U$37681 ( \45182 , RIdf96fa8_4990);
or \U$37682 ( \45183 , \45182 , \44724 );
not \U$37683 ( \45184 , \44895 );
and \U$37684 ( \45185 , \43969 , \45184 );
not \U$37685 ( \45186 , \45185 );
not \U$37686 ( \45187 , \43966 );
not \U$37687 ( \45188 , \44671 );
or \U$37688 ( \45189 , \45187 , \45188 );
nand \U$37689 ( \45190 , \45183 , \45186 , \45189 );
and \U$37690 ( \45191 , \45190 , \43589 );
or \U$37691 ( \45192 , \45181 , \45191 );
and \U$37693 ( \45193 , \45192 , 1'b1 );
or \U$37695 ( \45194 , \45193 , 1'b0 );
buf \U$37696 ( \45195 , \45194 );
_DC r23584_GF_IsGateDCbyConstraint ( \45196_nR23584 , \45195 , \21944 );
buf \U$37697 ( \45197 , \45196_nR23584 );
not \U$37698 ( \45198 , \44758 );
and \U$37699 ( \45199 , RIdf9a680_4991, \45198 );
not \U$37700 ( \45200 , RIdf9a680_4991);
or \U$37701 ( \45201 , \45200 , \44724 );
not \U$37702 ( \45202 , \44839 );
and \U$37703 ( \45203 , \43987 , \45202 );
not \U$37704 ( \45204 , \45203 );
not \U$37705 ( \45205 , \43985 );
not \U$37706 ( \45206 , \44670 );
or \U$37707 ( \45207 , \45205 , \45206 );
nand \U$37708 ( \45208 , \45201 , \45204 , \45207 );
and \U$37709 ( \45209 , \45208 , \44758 );
or \U$37710 ( \45210 , \45199 , \45209 );
and \U$37712 ( \45211 , \45210 , 1'b1 );
or \U$37714 ( \45212 , \45211 , 1'b0 );
buf \U$37715 ( \45213 , \45212 );
_DC r23586_GF_IsGateDCbyConstraint ( \45214_nR23586 , \45213 , \21944 );
buf \U$37716 ( \45215 , \45214_nR23586 );
not \U$37717 ( \45216 , \44758 );
and \U$37718 ( \45217 , RIdf9ccf0_4992, \45216 );
not \U$37719 ( \45218 , RIdf9ccf0_4992);
or \U$37720 ( \45219 , \45218 , \44662 );
not \U$37721 ( \45220 , \44839 );
and \U$37722 ( \45221 , \44006 , \45220 );
not \U$37723 ( \45222 , \45221 );
not \U$37724 ( \45223 , \44003 );
not \U$37725 ( \45224 , \44768 );
or \U$37726 ( \45225 , \45223 , \45224 );
nand \U$37727 ( \45226 , \45219 , \45222 , \45225 );
and \U$37728 ( \45227 , \45226 , \44758 );
or \U$37729 ( \45228 , \45217 , \45227 );
and \U$37731 ( \45229 , \45228 , 1'b1 );
or \U$37733 ( \45230 , \45229 , 1'b0 );
buf \U$37734 ( \45231 , \45230 );
_DC r2358a_GF_IsGateDCbyConstraint ( \45232_nR2358a , \45231 , \21944 );
buf \U$37735 ( \45233 , \45232_nR2358a );
not \U$37736 ( \45234 , \43589 );
and \U$37737 ( \45235 , RIdf9ec58_4993, \45234 );
not \U$37738 ( \45236 , RIdf9ec58_4993);
or \U$37739 ( \45237 , \45236 , \44724 );
not \U$37740 ( \45238 , \44665 );
and \U$37741 ( \45239 , \44025 , \45238 );
not \U$37742 ( \45240 , \45239 );
not \U$37743 ( \45241 , \44023 );
not \U$37744 ( \45242 , \44670 );
or \U$37745 ( \45243 , \45241 , \45242 );
nand \U$37746 ( \45244 , \45237 , \45240 , \45243 );
and \U$37747 ( \45245 , \45244 , \43589 );
or \U$37748 ( \45246 , \45235 , \45245 );
and \U$37750 ( \45247 , \45246 , 1'b1 );
or \U$37752 ( \45248 , \45247 , 1'b0 );
buf \U$37753 ( \45249 , \45248 );
_DC r2358c_GF_IsGateDCbyConstraint ( \45250_nR2358c , \45249 , \21944 );
buf \U$37754 ( \45251 , \45250_nR2358c );
not \U$37755 ( \45252 , \44018 );
and \U$37756 ( \45253 , RIdfa04b8_4994, \45252 );
not \U$37757 ( \45254 , RIdfa04b8_4994);
or \U$37758 ( \45255 , \45254 , \44705 );
not \U$37759 ( \45256 , \44839 );
and \U$37760 ( \45257 , \44043 , \45256 );
not \U$37761 ( \45258 , \45257 );
not \U$37762 ( \45259 , \44041 );
not \U$37763 ( \45260 , \44768 );
or \U$37764 ( \45261 , \45259 , \45260 );
nand \U$37765 ( \45262 , \45255 , \45258 , \45261 );
and \U$37766 ( \45263 , \45262 , \44018 );
or \U$37767 ( \45264 , \45253 , \45263 );
and \U$37769 ( \45265 , \45264 , 1'b1 );
or \U$37771 ( \45266 , \45265 , 1'b0 );
buf \U$37772 ( \45267 , \45266 );
_DC r2358e_GF_IsGateDCbyConstraint ( \45268_nR2358e , \45267 , \21944 );
buf \U$37773 ( \45269 , \45268_nR2358e );
not \U$37774 ( \45270 , \43377 );
and \U$37775 ( \45271 , RIdfa1bb0_4995, \45270 );
not \U$37776 ( \45272 , RIdfa1bb0_4995);
or \U$37777 ( \45273 , \45272 , \44662 );
not \U$37778 ( \45274 , \44876 );
and \U$37779 ( \45275 , \44062 , \45274 );
not \U$37780 ( \45276 , \45275 );
not \U$37781 ( \45277 , \44060 );
not \U$37782 ( \45278 , \44671 );
or \U$37783 ( \45279 , \45277 , \45278 );
nand \U$37784 ( \45280 , \45273 , \45276 , \45279 );
and \U$37785 ( \45281 , \45280 , \43377 );
or \U$37786 ( \45282 , \45271 , \45281 );
and \U$37788 ( \45283 , \45282 , 1'b1 );
or \U$37790 ( \45284 , \45283 , 1'b0 );
buf \U$37791 ( \45285 , \45284 );
_DC r23590_GF_IsGateDCbyConstraint ( \45286_nR23590 , \45285 , \21944 );
buf \U$37792 ( \45287 , \45286_nR23590 );
not \U$37793 ( \45288 , \43589 );
and \U$37794 ( \45289 , RIdfa3b18_4996, \45288 );
not \U$37795 ( \45290 , RIdfa3b18_4996);
or \U$37796 ( \45291 , \45290 , \44662 );
not \U$37797 ( \45292 , \44895 );
and \U$37798 ( \45293 , \44082 , \45292 );
not \U$37799 ( \45294 , \45293 );
not \U$37800 ( \45295 , \44079 );
not \U$37801 ( \45296 , \44691 );
or \U$37802 ( \45297 , \45295 , \45296 );
nand \U$37803 ( \45298 , \45291 , \45294 , \45297 );
and \U$37804 ( \45299 , \45298 , \43589 );
or \U$37805 ( \45300 , \45289 , \45299 );
and \U$37807 ( \45301 , \45300 , 1'b1 );
or \U$37809 ( \45302 , \45301 , 1'b0 );
buf \U$37810 ( \45303 , \45302 );
_DC r23592_GF_IsGateDCbyConstraint ( \45304_nR23592 , \45303 , \21944 );
buf \U$37811 ( \45305 , \45304_nR23592 );
not \U$37812 ( \45306 , \44758 );
and \U$37813 ( \45307 , RIdfa4dd8_4997, \45306 );
not \U$37814 ( \45308 , RIdfa4dd8_4997);
or \U$37815 ( \45309 , \45308 , \44724 );
not \U$37816 ( \45310 , \44783 );
and \U$37817 ( \45311 , \44101 , \45310 );
not \U$37818 ( \45312 , \45311 );
not \U$37819 ( \45313 , \44098 );
not \U$37820 ( \45314 , \44671 );
or \U$37821 ( \45315 , \45313 , \45314 );
nand \U$37822 ( \45316 , \45309 , \45312 , \45315 );
and \U$37823 ( \45317 , \45316 , \44758 );
or \U$37824 ( \45318 , \45307 , \45317 );
and \U$37826 ( \45319 , \45318 , 1'b1 );
or \U$37828 ( \45320 , \45319 , 1'b0 );
buf \U$37829 ( \45321 , \45320 );
_DC r23594_GF_IsGateDCbyConstraint ( \45322_nR23594 , \45321 , \21944 );
buf \U$37830 ( \45323 , \45322_nR23594 );
buf \U$37831 ( \45324 , \43482 );
not \U$37832 ( \45325 , \45324 );
and \U$37833 ( \45326 , RIdfa6110_4998, \45325 );
not \U$37834 ( \45327 , RIdfa6110_4998);
or \U$37835 ( \45328 , \45327 , \44724 );
not \U$37836 ( \45329 , \44665 );
and \U$37837 ( \45330 , \44119 , \45329 );
not \U$37838 ( \45331 , \45330 );
not \U$37839 ( \45332 , \44117 );
not \U$37840 ( \45333 , \44670 );
or \U$37841 ( \45334 , \45332 , \45333 );
nand \U$37842 ( \45335 , \45328 , \45331 , \45334 );
and \U$37843 ( \45336 , \45335 , \45324 );
or \U$37844 ( \45337 , \45326 , \45336 );
and \U$37846 ( \45338 , \45337 , 1'b1 );
or \U$37848 ( \45339 , \45338 , 1'b0 );
buf \U$37849 ( \45340 , \45339 );
_DC r23596_GF_IsGateDCbyConstraint ( \45341_nR23596 , \45340 , \21944 );
buf \U$37850 ( \45342 , \45341_nR23596 );
not \U$37851 ( \45343 , \44074 );
and \U$37852 ( \45344 , RIdfa75b0_4999, \45343 );
not \U$37853 ( \45345 , RIdfa75b0_4999);
or \U$37854 ( \45346 , \45345 , \44801 );
not \U$37855 ( \45347 , \44876 );
and \U$37856 ( \45348 , \44139 , \45347 );
not \U$37857 ( \45349 , \45348 );
not \U$37858 ( \45350 , \44136 );
not \U$37859 ( \45351 , \44670 );
or \U$37860 ( \45352 , \45350 , \45351 );
nand \U$37861 ( \45353 , \45346 , \45349 , \45352 );
and \U$37862 ( \45354 , \45353 , \44074 );
or \U$37863 ( \45355 , \45344 , \45354 );
and \U$37865 ( \45356 , \45355 , 1'b1 );
or \U$37867 ( \45357 , \45356 , 1'b0 );
buf \U$37868 ( \45358 , \45357 );
_DC r23598_GF_IsGateDCbyConstraint ( \45359_nR23598 , \45358 , \21944 );
buf \U$37869 ( \45360 , \45359_nR23598 );
buf \U$37870 ( \45361 , \44074 );
not \U$37871 ( \45362 , \45361 );
and \U$37872 ( \45363 , RIdfa88e8_5000, \45362 );
not \U$37873 ( \45364 , RIdfa88e8_5000);
or \U$37874 ( \45365 , \45364 , \44724 );
not \U$37875 ( \45366 , \44895 );
and \U$37876 ( \45367 , \44159 , \45366 );
not \U$37877 ( \45368 , \45367 );
not \U$37878 ( \45369 , \44156 );
not \U$37879 ( \45370 , \44691 );
or \U$37880 ( \45371 , \45369 , \45370 );
nand \U$37881 ( \45372 , \45365 , \45368 , \45371 );
and \U$37882 ( \45373 , \45372 , \45361 );
or \U$37883 ( \45374 , \45363 , \45373 );
and \U$37885 ( \45375 , \45374 , 1'b1 );
or \U$37887 ( \45376 , \45375 , 1'b0 );
buf \U$37888 ( \45377 , \45376 );
_DC r2359a_GF_IsGateDCbyConstraint ( \45378_nR2359a , \45377 , \21944 );
buf \U$37889 ( \45379 , \45378_nR2359a );
not \U$37890 ( \45380 , \45361 );
and \U$37891 ( \45381 , RIdfa9d10_5001, \45380 );
not \U$37892 ( \45382 , RIdfa9d10_5001);
or \U$37893 ( \45383 , \45382 , \44801 );
not \U$37894 ( \45384 , \44783 );
and \U$37895 ( \45385 , \44179 , \45384 );
not \U$37896 ( \45386 , \45385 );
not \U$37897 ( \45387 , \44176 );
not \U$37898 ( \45388 , \44671 );
or \U$37899 ( \45389 , \45387 , \45388 );
nand \U$37900 ( \45390 , \45383 , \45386 , \45389 );
and \U$37901 ( \45391 , \45390 , \45361 );
or \U$37902 ( \45392 , \45381 , \45391 );
and \U$37904 ( \45393 , \45392 , 1'b1 );
or \U$37906 ( \45394 , \45393 , 1'b0 );
buf \U$37907 ( \45395 , \45394 );
_DC r2359c_GF_IsGateDCbyConstraint ( \45396_nR2359c , \45395 , \21944 );
buf \U$37908 ( \45397 , \45396_nR2359c );
not \U$37909 ( \45398 , \44018 );
and \U$37910 ( \45399 , RIdfab048_5002, \45398 );
not \U$37911 ( \45400 , RIdfab048_5002);
or \U$37912 ( \45401 , \45400 , \44801 );
not \U$37913 ( \45402 , \44686 );
and \U$37914 ( \45403 , \44198 , \45402 );
not \U$37915 ( \45404 , \45403 );
not \U$37916 ( \45405 , \44196 );
not \U$37917 ( \45406 , \44671 );
or \U$37918 ( \45407 , \45405 , \45406 );
nand \U$37919 ( \45408 , \45401 , \45404 , \45407 );
and \U$37920 ( \45409 , \45408 , \44018 );
or \U$37921 ( \45410 , \45399 , \45409 );
and \U$37923 ( \45411 , \45410 , 1'b1 );
or \U$37925 ( \45412 , \45411 , 1'b0 );
buf \U$37926 ( \45413 , \45412 );
_DC r235a0_GF_IsGateDCbyConstraint ( \45414_nR235a0 , \45413 , \21944 );
buf \U$37927 ( \45415 , \45414_nR235a0 );
not \U$37928 ( \45416 , \45324 );
and \U$37929 ( \45417 , RIdfac218_5003, \45416 );
not \U$37930 ( \45418 , RIdfac218_5003);
or \U$37931 ( \45419 , \45418 , \44705 );
not \U$37932 ( \45420 , \44763 );
and \U$37933 ( \45421 , \44216 , \45420 );
not \U$37934 ( \45422 , \45421 );
not \U$37935 ( \45423 , \44214 );
not \U$37936 ( \45424 , \44768 );
or \U$37937 ( \45425 , \45423 , \45424 );
nand \U$37938 ( \45426 , \45419 , \45422 , \45425 );
and \U$37939 ( \45427 , \45426 , \45324 );
or \U$37940 ( \45428 , \45417 , \45427 );
and \U$37942 ( \45429 , \45428 , 1'b1 );
or \U$37944 ( \45430 , \45429 , 1'b0 );
buf \U$37945 ( \45431 , \45430 );
_DC r235a2_GF_IsGateDCbyConstraint ( \45432_nR235a2 , \45431 , \21944 );
buf \U$37946 ( \45433 , \45432_nR235a2 );
not \U$37947 ( \45434 , \45361 );
and \U$37948 ( \45435 , RIdfad460_5004, \45434 );
not \U$37949 ( \45436 , RIdfad460_5004);
or \U$37950 ( \45437 , \45436 , \44705 );
not \U$37951 ( \45438 , \44839 );
and \U$37952 ( \45439 , \44234 , \45438 );
not \U$37953 ( \45440 , \45439 );
not \U$37954 ( \45441 , \44232 );
not \U$37955 ( \45442 , \44691 );
or \U$37956 ( \45443 , \45441 , \45442 );
nand \U$37957 ( \45444 , \45437 , \45440 , \45443 );
and \U$37958 ( \45445 , \45444 , \45361 );
or \U$37959 ( \45446 , \45435 , \45445 );
and \U$37961 ( \45447 , \45446 , 1'b1 );
or \U$37963 ( \45448 , \45447 , 1'b0 );
buf \U$37964 ( \45449 , \45448 );
_DC r235a4_GF_IsGateDCbyConstraint ( \45450_nR235a4 , \45449 , \21944 );
buf \U$37965 ( \45451 , \45450_nR235a4 );
not \U$37966 ( \45452 , \43482 );
and \U$37967 ( \45453 , RIdfaecc0_5005, \45452 );
not \U$37968 ( \45454 , RIdfaecc0_5005);
or \U$37969 ( \45455 , \45454 , \44801 );
not \U$37970 ( \45456 , \44665 );
and \U$37971 ( \45457 , \44253 , \45456 );
not \U$37972 ( \45458 , \45457 );
not \U$37973 ( \45459 , \44251 );
not \U$37974 ( \45460 , \44671 );
or \U$37975 ( \45461 , \45459 , \45460 );
nand \U$37976 ( \45462 , \45455 , \45458 , \45461 );
and \U$37977 ( \45463 , \45462 , \43482 );
or \U$37978 ( \45464 , \45453 , \45463 );
and \U$37980 ( \45465 , \45464 , 1'b1 );
or \U$37982 ( \45466 , \45465 , 1'b0 );
buf \U$37983 ( \45467 , \45466 );
_DC r235a6_GF_IsGateDCbyConstraint ( \45468_nR235a6 , \45467 , \21944 );
buf \U$37984 ( \45469 , \45468_nR235a6 );
not \U$37985 ( \45470 , \45361 );
and \U$37986 ( \45471 , RIdfb0610_5006, \45470 );
not \U$37987 ( \45472 , RIdfb0610_5006);
or \U$37988 ( \45473 , \45472 , \44705 );
not \U$37989 ( \45474 , \44686 );
and \U$37990 ( \45475 , \44274 , \45474 );
not \U$37991 ( \45476 , \45475 );
not \U$37992 ( \45477 , \44271 );
not \U$37993 ( \45478 , \44691 );
or \U$37994 ( \45479 , \45477 , \45478 );
nand \U$37995 ( \45480 , \45473 , \45476 , \45479 );
and \U$37996 ( \45481 , \45480 , \45361 );
or \U$37997 ( \45482 , \45471 , \45481 );
and \U$37999 ( \45483 , \45482 , 1'b1 );
or \U$38001 ( \45484 , \45483 , 1'b0 );
buf \U$38002 ( \45485 , \45484 );
_DC r235a8_GF_IsGateDCbyConstraint ( \45486_nR235a8 , \45485 , \21944 );
buf \U$38003 ( \45487 , \45486_nR235a8 );
not \U$38004 ( \45488 , \45361 );
and \U$38005 ( \45489 , RIdfb1c90_5007, \45488 );
not \U$38006 ( \45490 , RIdfb1c90_5007);
or \U$38007 ( \45491 , \45490 , \44705 );
not \U$38008 ( \45492 , \44839 );
and \U$38009 ( \45493 , \44294 , \45492 );
not \U$38010 ( \45494 , \45493 );
not \U$38011 ( \45495 , \44291 );
not \U$38012 ( \45496 , \44768 );
or \U$38013 ( \45497 , \45495 , \45496 );
nand \U$38014 ( \45498 , \45491 , \45494 , \45497 );
and \U$38015 ( \45499 , \45498 , \45361 );
or \U$38016 ( \45500 , \45489 , \45499 );
and \U$38018 ( \45501 , \45500 , 1'b1 );
or \U$38020 ( \45502 , \45501 , 1'b0 );
buf \U$38021 ( \45503 , \45502 );
_DC r235aa_GF_IsGateDCbyConstraint ( \45504_nR235aa , \45503 , \21944 );
buf \U$38022 ( \45505 , \45504_nR235aa );
not \U$38023 ( \45506 , \43589 );
and \U$38024 ( \45507 , RIdfb3310_5008, \45506 );
not \U$38025 ( \45508 , RIdfb3310_5008);
or \U$38026 ( \45509 , \45508 , \44662 );
not \U$38027 ( \45510 , \44763 );
and \U$38028 ( \45511 , \44314 , \45510 );
not \U$38029 ( \45512 , \45511 );
not \U$38030 ( \45513 , \44311 );
not \U$38031 ( \45514 , \44671 );
or \U$38032 ( \45515 , \45513 , \45514 );
nand \U$38033 ( \45516 , \45509 , \45512 , \45515 );
and \U$38034 ( \45517 , \45516 , \43589 );
or \U$38035 ( \45518 , \45507 , \45517 );
and \U$38037 ( \45519 , \45518 , 1'b1 );
or \U$38039 ( \45520 , \45519 , 1'b0 );
buf \U$38040 ( \45521 , \45520 );
_DC r235ac_GF_IsGateDCbyConstraint ( \45522_nR235ac , \45521 , \21944 );
buf \U$38041 ( \45523 , \45522_nR235ac );
not \U$38042 ( \45524 , \45324 );
and \U$38043 ( \45525 , RIdfb4828_5009, \45524 );
not \U$38044 ( \45526 , RIdfb4828_5009);
or \U$38045 ( \45527 , \45526 , \44724 );
not \U$38046 ( \45528 , \44839 );
and \U$38047 ( \45529 , \44332 , \45528 );
not \U$38048 ( \45530 , \45529 );
not \U$38049 ( \45531 , \44330 );
not \U$38050 ( \45532 , \44768 );
or \U$38051 ( \45533 , \45531 , \45532 );
nand \U$38052 ( \45534 , \45527 , \45530 , \45533 );
and \U$38053 ( \45535 , \45534 , \45324 );
or \U$38054 ( \45536 , \45525 , \45535 );
and \U$38056 ( \45537 , \45536 , 1'b1 );
or \U$38058 ( \45538 , \45537 , 1'b0 );
buf \U$38059 ( \45539 , \45538 );
_DC r235ae_GF_IsGateDCbyConstraint ( \45540_nR235ae , \45539 , \21944 );
buf \U$38060 ( \45541 , \45540_nR235ae );
not \U$38061 ( \45542 , \45324 );
and \U$38062 ( \45543 , RIdfb5d40_5010, \45542 );
not \U$38063 ( \45544 , RIdfb5d40_5010);
or \U$38064 ( \45545 , \45544 , \44705 );
not \U$38065 ( \45546 , \44895 );
and \U$38066 ( \45547 , \44352 , \45546 );
not \U$38067 ( \45548 , \45547 );
not \U$38068 ( \45549 , \44349 );
not \U$38069 ( \45550 , \44671 );
or \U$38070 ( \45551 , \45549 , \45550 );
nand \U$38071 ( \45552 , \45545 , \45548 , \45551 );
and \U$38072 ( \45553 , \45552 , \45324 );
or \U$38073 ( \45554 , \45543 , \45553 );
and \U$38075 ( \45555 , \45554 , 1'b1 );
or \U$38077 ( \45556 , \45555 , 1'b0 );
buf \U$38078 ( \45557 , \45556 );
_DC r235b0_GF_IsGateDCbyConstraint ( \45558_nR235b0 , \45557 , \21944 );
buf \U$38079 ( \45559 , \45558_nR235b0 );
not \U$38080 ( \45560 , \43710 );
and \U$38081 ( \45561 , RIdfb77f8_5011, \45560 );
not \U$38082 ( \45562 , RIdfb77f8_5011);
or \U$38083 ( \45563 , \45562 , \44801 );
not \U$38084 ( \45564 , \44839 );
and \U$38085 ( \45565 , \44370 , \45564 );
not \U$38086 ( \45566 , \45565 );
not \U$38087 ( \45567 , \44368 );
not \U$38088 ( \45568 , \44768 );
or \U$38089 ( \45569 , \45567 , \45568 );
nand \U$38090 ( \45570 , \45563 , \45566 , \45569 );
and \U$38091 ( \45571 , \45570 , \43710 );
or \U$38092 ( \45572 , \45561 , \45571 );
and \U$38094 ( \45573 , \45572 , 1'b1 );
or \U$38096 ( \45574 , \45573 , 1'b0 );
buf \U$38097 ( \45575 , \45574 );
_DC r235b2_GF_IsGateDCbyConstraint ( \45576_nR235b2 , \45575 , \21944 );
buf \U$38098 ( \45577 , \45576_nR235b2 );
not \U$38099 ( \45578 , \45324 );
and \U$38100 ( \45579 , RIdfb92b0_5012, \45578 );
not \U$38101 ( \45580 , RIdfb92b0_5012);
or \U$38102 ( \45581 , \45580 , \44705 );
not \U$38103 ( \45582 , \44839 );
and \U$38104 ( \45583 , \44388 , \45582 );
not \U$38105 ( \45584 , \45583 );
not \U$38106 ( \45585 , \44386 );
not \U$38107 ( \45586 , \44768 );
or \U$38108 ( \45587 , \45585 , \45586 );
nand \U$38109 ( \45588 , \45581 , \45584 , \45587 );
and \U$38110 ( \45589 , \45588 , \45324 );
or \U$38111 ( \45590 , \45579 , \45589 );
and \U$38113 ( \45591 , \45590 , 1'b1 );
or \U$38115 ( \45592 , \45591 , 1'b0 );
buf \U$38116 ( \45593 , \45592 );
_DC r235b6_GF_IsGateDCbyConstraint ( \45594_nR235b6 , \45593 , \21944 );
buf \U$38117 ( \45595 , \45594_nR235b6 );
not \U$38118 ( \45596 , \45361 );
and \U$38119 ( \45597 , RIdfba9a8_5013, \45596 );
not \U$38120 ( \45598 , RIdfba9a8_5013);
or \U$38121 ( \45599 , \45598 , \44801 );
not \U$38122 ( \45600 , \44876 );
and \U$38123 ( \45601 , \44407 , \45600 );
not \U$38124 ( \45602 , \45601 );
not \U$38125 ( \45603 , \44405 );
not \U$38126 ( \45604 , \44691 );
or \U$38127 ( \45605 , \45603 , \45604 );
nand \U$38128 ( \45606 , \45599 , \45602 , \45605 );
and \U$38129 ( \45607 , \45606 , \45361 );
or \U$38130 ( \45608 , \45597 , \45607 );
and \U$38132 ( \45609 , \45608 , 1'b1 );
or \U$38134 ( \45610 , \45609 , 1'b0 );
buf \U$38135 ( \45611 , \45610 );
_DC r235b8_GF_IsGateDCbyConstraint ( \45612_nR235b8 , \45611 , \21944 );
buf \U$38136 ( \45613 , \45612_nR235b8 );
buf \U$38137 ( \45614 , \44591 );
not \U$38138 ( \45615 , \45614 );
and \U$38139 ( \45616 , RIddf2ca8_5014, \45615 );
not \U$38140 ( \45617 , RIddf2ca8_5014);
or \U$38141 ( \45618 , \45617 , \44801 );
not \U$38142 ( \45619 , \44895 );
and \U$38143 ( \45620 , \44425 , \45619 );
not \U$38144 ( \45621 , \45620 );
not \U$38145 ( \45622 , \44423 );
not \U$38146 ( \45623 , \44768 );
or \U$38147 ( \45624 , \45622 , \45623 );
nand \U$38148 ( \45625 , \45618 , \45621 , \45624 );
and \U$38149 ( \45626 , \45625 , \45614 );
or \U$38150 ( \45627 , \45616 , \45626 );
and \U$38152 ( \45628 , \45627 , 1'b1 );
or \U$38154 ( \45629 , \45628 , 1'b0 );
buf \U$38155 ( \45630 , \45629 );
_DC r235ba_GF_IsGateDCbyConstraint ( \45631_nR235ba , \45630 , \21944 );
buf \U$38156 ( \45632 , \45631_nR235ba );
not \U$38157 ( \45633 , \45324 );
and \U$38158 ( \45634 , RIddf4580_5015, \45633 );
not \U$38159 ( \45635 , RIddf4580_5015);
or \U$38160 ( \45636 , \45635 , \44724 );
not \U$38161 ( \45637 , \44783 );
and \U$38162 ( \45638 , \44445 , \45637 );
not \U$38163 ( \45639 , \45638 );
not \U$38164 ( \45640 , \44442 );
not \U$38165 ( \45641 , \44768 );
or \U$38166 ( \45642 , \45640 , \45641 );
nand \U$38167 ( \45643 , \45636 , \45639 , \45642 );
and \U$38168 ( \45644 , \45643 , \45324 );
or \U$38169 ( \45645 , \45634 , \45644 );
and \U$38171 ( \45646 , \45645 , 1'b1 );
or \U$38173 ( \45647 , \45646 , 1'b0 );
buf \U$38174 ( \45648 , \45647 );
_DC r235bc_GF_IsGateDCbyConstraint ( \45649_nR235bc , \45648 , \21944 );
buf \U$38175 ( \45650 , \45649_nR235bc );
not \U$38176 ( \45651 , \45324 );
and \U$38177 ( \45652 , RIddf6308_5016, \45651 );
not \U$38178 ( \45653 , RIddf6308_5016);
or \U$38179 ( \45654 , \45653 , \44662 );
not \U$38180 ( \45655 , \44876 );
and \U$38181 ( \45656 , \44463 , \45655 );
not \U$38182 ( \45657 , \45656 );
not \U$38183 ( \45658 , \44461 );
not \U$38184 ( \45659 , \44671 );
or \U$38185 ( \45660 , \45658 , \45659 );
nand \U$38186 ( \45661 , \45654 , \45657 , \45660 );
and \U$38187 ( \45662 , \45661 , \45324 );
or \U$38188 ( \45663 , \45652 , \45662 );
and \U$38190 ( \45664 , \45663 , 1'b1 );
or \U$38192 ( \45665 , \45664 , 1'b0 );
buf \U$38193 ( \45666 , \45665 );
_DC r235be_GF_IsGateDCbyConstraint ( \45667_nR235be , \45666 , \21944 );
buf \U$38194 ( \45668 , \45667_nR235be );
not \U$38195 ( \45669 , \45614 );
and \U$38196 ( \45670 , RIddf8270_5017, \45669 );
not \U$38197 ( \45671 , RIddf8270_5017);
or \U$38198 ( \45672 , \45671 , \44662 );
not \U$38199 ( \45673 , \44665 );
and \U$38200 ( \45674 , \44481 , \45673 );
not \U$38201 ( \45675 , \45674 );
not \U$38202 ( \45676 , \44479 );
not \U$38203 ( \45677 , \44691 );
or \U$38204 ( \45678 , \45676 , \45677 );
nand \U$38205 ( \45679 , \45672 , \45675 , \45678 );
and \U$38206 ( \45680 , \45679 , \45614 );
or \U$38207 ( \45681 , \45670 , \45680 );
and \U$38209 ( \45682 , \45681 , 1'b1 );
or \U$38211 ( \45683 , \45682 , 1'b0 );
buf \U$38212 ( \45684 , \45683 );
_DC r235c0_GF_IsGateDCbyConstraint ( \45685_nR235c0 , \45684 , \21944 );
buf \U$38213 ( \45686 , \45685_nR235c0 );
not \U$38214 ( \45687 , \45361 );
and \U$38215 ( \45688 , RIddf9e90_5018, \45687 );
not \U$38216 ( \45689 , RIddf9e90_5018);
or \U$38217 ( \45690 , \45689 , \44724 );
not \U$38218 ( \45691 , \44839 );
and \U$38219 ( \45692 , \44503 , \45691 );
not \U$38220 ( \45693 , \45692 );
not \U$38221 ( \45694 , \44500 );
not \U$38222 ( \45695 , \44671 );
or \U$38223 ( \45696 , \45694 , \45695 );
nand \U$38224 ( \45697 , \45690 , \45693 , \45696 );
and \U$38225 ( \45698 , \45697 , \45361 );
or \U$38226 ( \45699 , \45688 , \45698 );
and \U$38228 ( \45700 , \45699 , 1'b1 );
or \U$38230 ( \45701 , \45700 , 1'b0 );
buf \U$38231 ( \45702 , \45701 );
_DC r235c2_GF_IsGateDCbyConstraint ( \45703_nR235c2 , \45702 , \21944 );
buf \U$38232 ( \45704 , \45703_nR235c2 );
not \U$38233 ( \45705 , \45361 );
and \U$38234 ( \45706 , RIddfbdf8_5019, \45705 );
not \U$38235 ( \45707 , RIddfbdf8_5019);
or \U$38236 ( \45708 , \45707 , \44724 );
not \U$38237 ( \45709 , \44876 );
and \U$38238 ( \45710 , \44524 , \45709 );
not \U$38239 ( \45711 , \45710 );
not \U$38240 ( \45712 , \44521 );
not \U$38241 ( \45713 , \44691 );
or \U$38242 ( \45714 , \45712 , \45713 );
nand \U$38243 ( \45715 , \45708 , \45711 , \45714 );
and \U$38244 ( \45716 , \45715 , \45361 );
or \U$38245 ( \45717 , \45706 , \45716 );
and \U$38247 ( \45718 , \45717 , 1'b1 );
or \U$38249 ( \45719 , \45718 , 1'b0 );
buf \U$38250 ( \45720 , \45719 );
_DC r235c4_GF_IsGateDCbyConstraint ( \45721_nR235c4 , \45720 , \21944 );
buf \U$38251 ( \45722 , \45721_nR235c4 );
not \U$38252 ( \45723 , \45614 );
and \U$38253 ( \45724 , RIddfdb08_5020, \45723 );
not \U$38254 ( \45725 , RIddfdb08_5020);
or \U$38255 ( \45726 , \45725 , \44801 );
not \U$38256 ( \45727 , \44895 );
and \U$38257 ( \45728 , \44543 , \45727 );
not \U$38258 ( \45729 , \45728 );
not \U$38259 ( \45730 , \44540 );
not \U$38260 ( \45731 , \44691 );
or \U$38261 ( \45732 , \45730 , \45731 );
nand \U$38262 ( \45733 , \45726 , \45729 , \45732 );
and \U$38263 ( \45734 , \45733 , \45614 );
or \U$38264 ( \45735 , \45724 , \45734 );
and \U$38266 ( \45736 , \45735 , 1'b1 );
or \U$38268 ( \45737 , \45736 , 1'b0 );
buf \U$38269 ( \45738 , \45737 );
_DC r235c6_GF_IsGateDCbyConstraint ( \45739_nR235c6 , \45738 , \21944 );
buf \U$38270 ( \45740 , \45739_nR235c6 );
not \U$38271 ( \45741 , \45324 );
and \U$38272 ( \45742 , RIddff548_5021, \45741 );
not \U$38273 ( \45743 , RIddff548_5021);
or \U$38274 ( \45744 , \45743 , \44705 );
not \U$38275 ( \45745 , \44686 );
and \U$38276 ( \45746 , \44561 , \45745 );
not \U$38277 ( \45747 , \45746 );
not \U$38278 ( \45748 , \44559 );
not \U$38279 ( \45749 , \44670 );
or \U$38280 ( \45750 , \45748 , \45749 );
nand \U$38281 ( \45751 , \45744 , \45747 , \45750 );
and \U$38282 ( \45752 , \45751 , \45324 );
or \U$38283 ( \45753 , \45742 , \45752 );
and \U$38285 ( \45754 , \45753 , 1'b1 );
or \U$38287 ( \45755 , \45754 , 1'b0 );
buf \U$38288 ( \45756 , \45755 );
_DC r235c8_GF_IsGateDCbyConstraint ( \45757_nR235c8 , \45756 , \21944 );
buf \U$38289 ( \45758 , \45757_nR235c8 );
not \U$38290 ( \45759 , \45324 );
and \U$38291 ( \45760 , RIde015a0_5022, \45759 );
not \U$38292 ( \45761 , RIde015a0_5022);
or \U$38293 ( \45762 , \45761 , \44705 );
not \U$38294 ( \45763 , \44839 );
and \U$38295 ( \45764 , \44579 , \45763 );
not \U$38296 ( \45765 , \45764 );
not \U$38297 ( \45766 , \44577 );
not \U$38298 ( \45767 , \44768 );
or \U$38299 ( \45768 , \45766 , \45767 );
nand \U$38300 ( \45769 , \45762 , \45765 , \45768 );
and \U$38301 ( \45770 , \45769 , \45324 );
or \U$38302 ( \45771 , \45760 , \45770 );
and \U$38304 ( \45772 , \45771 , 1'b1 );
or \U$38306 ( \45773 , \45772 , 1'b0 );
buf \U$38307 ( \45774 , \45773 );
_DC r235cc_GF_IsGateDCbyConstraint ( \45775_nR235cc , \45774 , \21944 );
buf \U$38308 ( \45776 , \45775_nR235cc );
not \U$38309 ( \45777 , \45614 );
and \U$38310 ( \45778 , RIde03508_5023, \45777 );
not \U$38311 ( \45779 , RIde03508_5023);
or \U$38312 ( \45780 , \45779 , \44662 );
not \U$38313 ( \45781 , \44876 );
and \U$38314 ( \45782 , \44599 , \45781 );
not \U$38315 ( \45783 , \45782 );
not \U$38316 ( \45784 , \44596 );
not \U$38317 ( \45785 , \44691 );
or \U$38318 ( \45786 , \45784 , \45785 );
nand \U$38319 ( \45787 , \45780 , \45783 , \45786 );
and \U$38320 ( \45788 , \45787 , \45614 );
or \U$38321 ( \45789 , \45778 , \45788 );
and \U$38323 ( \45790 , \45789 , 1'b1 );
or \U$38325 ( \45791 , \45790 , 1'b0 );
buf \U$38326 ( \45792 , \45791 );
_DC r235ce_GF_IsGateDCbyConstraint ( \45793_nR235ce , \45792 , \21944 );
buf \U$38327 ( \45794 , \45793_nR235ce );
not \U$38328 ( \45795 , \45361 );
and \U$38329 ( \45796 , RIde04fc0_5024, \45795 );
not \U$38330 ( \45797 , RIde04fc0_5024);
or \U$38331 ( \45798 , \45797 , \44705 );
not \U$38332 ( \45799 , \44763 );
and \U$38333 ( \45800 , \44618 , \45799 );
not \U$38334 ( \45801 , \45800 );
not \U$38335 ( \45802 , \44615 );
not \U$38336 ( \45803 , \44691 );
or \U$38337 ( \45804 , \45802 , \45803 );
nand \U$38338 ( \45805 , \45798 , \45801 , \45804 );
and \U$38339 ( \45806 , \45805 , \45361 );
or \U$38340 ( \45807 , \45796 , \45806 );
and \U$38342 ( \45808 , \45807 , 1'b1 );
or \U$38344 ( \45809 , \45808 , 1'b0 );
buf \U$38345 ( \45810 , \45809 );
_DC r235d0_GF_IsGateDCbyConstraint ( \45811_nR235d0 , \45810 , \21944 );
buf \U$38346 ( \45812 , \45811_nR235d0 );
not \U$38347 ( \45813 , \45614 );
and \U$38348 ( \45814 , RIe03bbe8_5025, \45813 );
not \U$38349 ( \45815 , RIe03bbe8_5025);
or \U$38350 ( \45816 , \45815 , \44724 );
not \U$38351 ( \45817 , \44895 );
and \U$38352 ( \45818 , \44636 , \45817 );
not \U$38353 ( \45819 , \45818 );
not \U$38354 ( \45820 , \44634 );
not \U$38355 ( \45821 , \44691 );
or \U$38356 ( \45822 , \45820 , \45821 );
nand \U$38357 ( \45823 , \45816 , \45819 , \45822 );
and \U$38358 ( \45824 , \45823 , \45614 );
or \U$38359 ( \45825 , \45814 , \45824 );
and \U$38361 ( \45826 , \45825 , 1'b1 );
or \U$38363 ( \45827 , \45826 , 1'b0 );
buf \U$38364 ( \45828 , \45827 );
_DC r235d2_GF_IsGateDCbyConstraint ( \45829_nR235d2 , \45828 , \21944 );
buf \U$38365 ( \45830 , \45829_nR235d2 );
not \U$38366 ( \45831 , \45324 );
and \U$38367 ( \45832 , RIe039cf8_5026, \45831 );
not \U$38368 ( \45833 , RIe039cf8_5026);
not \U$38369 ( \45834 , \43392 );
nor \U$38370 ( \45835 , \43395 , \45834 );
nand \U$38371 ( \45836 , \45835 , \43397 );
not \U$38372 ( \45837 , \45836 );
not \U$38373 ( \45838 , \43385 );
or \U$38374 ( \45839 , \43383 , \45838 );
not \U$38375 ( \45840 , \45839 );
nand \U$38376 ( \45841 , \43374 , \45840 );
not \U$38377 ( \45842 , \45841 );
or \U$38378 ( \45843 , \45837 , \45842 );
not \U$38379 ( \45844 , \45843 );
not \U$38380 ( \45845 , \45844 );
or \U$38381 ( \45846 , \45833 , \45845 );
not \U$38382 ( \45847 , \45836 );
not \U$38383 ( \45848 , \45847 );
not \U$38384 ( \45849 , \45848 );
and \U$38385 ( \45850 , \43409 , \45849 );
not \U$38386 ( \45851 , \45850 );
not \U$38387 ( \45852 , \45841 );
buf \U$38388 ( \45853 , \45852 );
not \U$38389 ( \45854 , \45853 );
or \U$38390 ( \45855 , \44669 , \45854 );
nand \U$38391 ( \45856 , \45846 , \45851 , \45855 );
and \U$38392 ( \45857 , \45856 , \45324 );
or \U$38393 ( \45858 , \45832 , \45857 );
and \U$38395 ( \45859 , \45858 , 1'b1 );
or \U$38397 ( \45860 , \45859 , 1'b0 );
buf \U$38398 ( \45861 , \45860 );
_DC r235dc_GF_IsGateDCbyConstraint ( \45862_nR235dc , \45861 , \21944 );
buf \U$38399 ( \45863 , \45862_nR235dc );
not \U$38400 ( \45864 , \45614 );
and \U$38401 ( \45865 , RIe038600_5027, \45864 );
not \U$38402 ( \45866 , RIe038600_5027);
or \U$38403 ( \45867 , \45866 , \45845 );
not \U$38404 ( \45868 , \45837 );
not \U$38405 ( \45869 , \45868 );
and \U$38406 ( \45870 , \43430 , \45869 );
not \U$38407 ( \45871 , \45870 );
buf \U$38408 ( \45872 , \45852 );
not \U$38409 ( \45873 , \45872 );
or \U$38410 ( \45874 , \44690 , \45873 );
nand \U$38411 ( \45875 , \45867 , \45871 , \45874 );
and \U$38412 ( \45876 , \45875 , \45614 );
or \U$38413 ( \45877 , \45865 , \45876 );
and \U$38415 ( \45878 , \45877 , 1'b1 );
or \U$38417 ( \45879 , \45878 , 1'b0 );
buf \U$38418 ( \45880 , \45879 );
_DC r235f2_GF_IsGateDCbyConstraint ( \45881_nR235f2 , \45880 , \21944 );
buf \U$38419 ( \45882 , \45881_nR235f2 );
not \U$38420 ( \45883 , \45361 );
and \U$38421 ( \45884 , RIe0363c8_5028, \45883 );
not \U$38422 ( \45885 , RIe0363c8_5028);
or \U$38423 ( \45886 , \45885 , \45845 );
not \U$38424 ( \45887 , \45848 );
and \U$38425 ( \45888 , \43450 , \45887 );
not \U$38426 ( \45889 , \45888 );
not \U$38427 ( \45890 , \45853 );
or \U$38428 ( \45891 , \44710 , \45890 );
nand \U$38429 ( \45892 , \45886 , \45889 , \45891 );
and \U$38430 ( \45893 , \45892 , \45361 );
or \U$38431 ( \45894 , \45884 , \45893 );
and \U$38433 ( \45895 , \45894 , 1'b1 );
or \U$38435 ( \45896 , \45895 , 1'b0 );
buf \U$38436 ( \45897 , \45896 );
_DC r23608_GF_IsGateDCbyConstraint ( \45898_nR23608 , \45897 , \21944 );
buf \U$38437 ( \45899 , \45898_nR23608 );
not \U$38438 ( \45900 , \45324 );
and \U$38439 ( \45901 , RIe033b78_5029, \45900 );
not \U$38440 ( \45902 , RIe033b78_5029);
not \U$38441 ( \45903 , \45844 );
or \U$38442 ( \45904 , \45902 , \45903 );
not \U$38443 ( \45905 , \45868 );
and \U$38444 ( \45906 , \43470 , \45905 );
not \U$38445 ( \45907 , \45906 );
not \U$38446 ( \45908 , \45853 );
or \U$38447 ( \45909 , \44729 , \45908 );
nand \U$38448 ( \45910 , \45904 , \45907 , \45909 );
and \U$38449 ( \45911 , \45910 , \45324 );
or \U$38450 ( \45912 , \45901 , \45911 );
and \U$38452 ( \45913 , \45912 , 1'b1 );
or \U$38454 ( \45914 , \45913 , 1'b0 );
buf \U$38455 ( \45915 , \45914 );
_DC r2361e_GF_IsGateDCbyConstraint ( \45916_nR2361e , \45915 , \21944 );
buf \U$38456 ( \45917 , \45916_nR2361e );
not \U$38457 ( \45918 , \45614 );
and \U$38458 ( \45919 , RIe031580_5030, \45918 );
not \U$38459 ( \45920 , RIe031580_5030);
not \U$38460 ( \45921 , \45844 );
or \U$38461 ( \45922 , \45920 , \45921 );
not \U$38462 ( \45923 , \45848 );
and \U$38463 ( \45924 , \43491 , \45923 );
not \U$38464 ( \45925 , \45924 );
not \U$38465 ( \45926 , \45872 );
or \U$38466 ( \45927 , \44747 , \45926 );
nand \U$38467 ( \45928 , \45922 , \45925 , \45927 );
and \U$38468 ( \45929 , \45928 , \45614 );
or \U$38469 ( \45930 , \45919 , \45929 );
and \U$38471 ( \45931 , \45930 , 1'b1 );
or \U$38473 ( \45932 , \45931 , 1'b0 );
buf \U$38474 ( \45933 , \45932 );
_DC r23634_GF_IsGateDCbyConstraint ( \45934_nR23634 , \45933 , \21944 );
buf \U$38475 ( \45935 , \45934_nR23634 );
not \U$38476 ( \45936 , \45361 );
and \U$38477 ( \45937 , RIe02ee98_5031, \45936 );
not \U$38478 ( \45938 , RIe02ee98_5031);
or \U$38479 ( \45939 , \45938 , \45921 );
not \U$38480 ( \45940 , \45837 );
not \U$38481 ( \45941 , \45940 );
and \U$38482 ( \45942 , \43510 , \45941 );
not \U$38483 ( \45943 , \45942 );
buf \U$38484 ( \45944 , \45852 );
not \U$38485 ( \45945 , \45944 );
or \U$38486 ( \45946 , \44767 , \45945 );
nand \U$38487 ( \45947 , \45939 , \45943 , \45946 );
and \U$38488 ( \45948 , \45947 , \45361 );
or \U$38489 ( \45949 , \45937 , \45948 );
and \U$38491 ( \45950 , \45949 , 1'b1 );
or \U$38493 ( \45951 , \45950 , 1'b0 );
buf \U$38494 ( \45952 , \45951 );
_DC r2364a_GF_IsGateDCbyConstraint ( \45953_nR2364a , \45952 , \21944 );
buf \U$38495 ( \45954 , \45953_nR2364a );
not \U$38496 ( \45955 , \45324 );
and \U$38497 ( \45956 , RIe02c4e0_5032, \45955 );
not \U$38498 ( \45957 , RIe02c4e0_5032);
or \U$38499 ( \45958 , \45957 , \45845 );
not \U$38500 ( \45959 , \45847 );
not \U$38501 ( \45960 , \45959 );
and \U$38502 ( \45961 , \43535 , \45960 );
not \U$38503 ( \45962 , \45961 );
not \U$38504 ( \45963 , \45872 );
or \U$38505 ( \45964 , \44787 , \45963 );
nand \U$38506 ( \45965 , \45958 , \45962 , \45964 );
and \U$38507 ( \45966 , \45965 , \45324 );
or \U$38508 ( \45967 , \45956 , \45966 );
and \U$38510 ( \45968 , \45967 , 1'b1 );
or \U$38512 ( \45969 , \45968 , 1'b0 );
buf \U$38513 ( \45970 , \45969 );
_DC r23654_GF_IsGateDCbyConstraint ( \45971_nR23654 , \45970 , \21944 );
buf \U$38514 ( \45972 , \45971_nR23654 );
not \U$38515 ( \45973 , \45614 );
and \U$38516 ( \45974 , RIe02a488_5033, \45973 );
not \U$38517 ( \45975 , RIe02a488_5033);
not \U$38518 ( \45976 , \45844 );
or \U$38519 ( \45977 , \45975 , \45976 );
not \U$38520 ( \45978 , \45868 );
and \U$38521 ( \45979 , \43555 , \45978 );
not \U$38522 ( \45980 , \45979 );
not \U$38523 ( \45981 , \45944 );
or \U$38524 ( \45982 , \44806 , \45981 );
nand \U$38525 ( \45983 , \45977 , \45980 , \45982 );
and \U$38526 ( \45984 , \45983 , \45614 );
or \U$38527 ( \45985 , \45974 , \45984 );
and \U$38529 ( \45986 , \45985 , 1'b1 );
or \U$38531 ( \45987 , \45986 , 1'b0 );
buf \U$38532 ( \45988 , \45987 );
_DC r23656_GF_IsGateDCbyConstraint ( \45989_nR23656 , \45988 , \21944 );
buf \U$38533 ( \45990 , \45989_nR23656 );
not \U$38534 ( \45991 , \45361 );
and \U$38535 ( \45992 , RIe028958_5034, \45991 );
not \U$38536 ( \45993 , RIe028958_5034);
or \U$38537 ( \45994 , \45993 , \45845 );
not \U$38538 ( \45995 , \45940 );
and \U$38539 ( \45996 , \43576 , \45995 );
not \U$38540 ( \45997 , \45996 );
not \U$38541 ( \45998 , \45944 );
or \U$38542 ( \45999 , \44824 , \45998 );
nand \U$38543 ( \46000 , \45994 , \45997 , \45999 );
and \U$38544 ( \46001 , \46000 , \45361 );
or \U$38545 ( \46002 , \45992 , \46001 );
and \U$38547 ( \46003 , \46002 , 1'b1 );
or \U$38549 ( \46004 , \46003 , 1'b0 );
buf \U$38550 ( \46005 , \46004 );
_DC r23658_GF_IsGateDCbyConstraint ( \46006_nR23658 , \46005 , \21944 );
buf \U$38551 ( \46007 , \46006_nR23658 );
buf \U$38552 ( \46008 , \44591 );
not \U$38553 ( \46009 , \46008 );
and \U$38554 ( \46010 , RIe026b58_5035, \46009 );
not \U$38555 ( \46011 , RIe026b58_5035);
or \U$38556 ( \46012 , \46011 , \45921 );
not \U$38557 ( \46013 , \45847 );
not \U$38558 ( \46014 , \46013 );
and \U$38559 ( \46015 , \43597 , \46014 );
not \U$38560 ( \46016 , \46015 );
not \U$38561 ( \46017 , \45853 );
or \U$38562 ( \46018 , \44843 , \46017 );
nand \U$38563 ( \46019 , \46012 , \46016 , \46018 );
and \U$38564 ( \46020 , \46019 , \46008 );
or \U$38565 ( \46021 , \46010 , \46020 );
and \U$38567 ( \46022 , \46021 , 1'b1 );
or \U$38569 ( \46023 , \46022 , 1'b0 );
buf \U$38570 ( \46024 , \46023 );
_DC r2365a_GF_IsGateDCbyConstraint ( \46025_nR2365a , \46024 , \21944 );
buf \U$38571 ( \46026 , \46025_nR2365a );
not \U$38572 ( \46027 , \45614 );
and \U$38573 ( \46028 , RIe025460_5036, \46027 );
not \U$38574 ( \46029 , RIe025460_5036);
or \U$38575 ( \46030 , \46029 , \45976 );
not \U$38576 ( \46031 , \46013 );
and \U$38577 ( \46032 , \43622 , \46031 );
not \U$38578 ( \46033 , \46032 );
not \U$38579 ( \46034 , \45944 );
or \U$38580 ( \46035 , \44861 , \46034 );
nand \U$38581 ( \46036 , \46030 , \46033 , \46035 );
and \U$38582 ( \46037 , \46036 , \45614 );
or \U$38583 ( \46038 , \46028 , \46037 );
and \U$38585 ( \46039 , \46038 , 1'b1 );
or \U$38587 ( \46040 , \46039 , 1'b0 );
buf \U$38588 ( \46041 , \46040 );
_DC r235de_GF_IsGateDCbyConstraint ( \46042_nR235de , \46041 , \21944 );
buf \U$38589 ( \46043 , \46042_nR235de );
buf \U$38590 ( \46044 , \44074 );
not \U$38591 ( \46045 , \46044 );
and \U$38592 ( \46046 , RIe023b88_5037, \46045 );
not \U$38593 ( \46047 , RIe023b88_5037);
or \U$38594 ( \46048 , \46047 , \45921 );
not \U$38595 ( \46049 , \45847 );
not \U$38596 ( \46050 , \46049 );
and \U$38597 ( \46051 , \43640 , \46050 );
not \U$38598 ( \46052 , \46051 );
not \U$38599 ( \46053 , \45853 );
or \U$38600 ( \46054 , \44880 , \46053 );
nand \U$38601 ( \46055 , \46048 , \46052 , \46054 );
and \U$38602 ( \46056 , \46055 , \46044 );
or \U$38603 ( \46057 , \46046 , \46056 );
and \U$38605 ( \46058 , \46057 , 1'b1 );
or \U$38607 ( \46059 , \46058 , 1'b0 );
buf \U$38608 ( \46060 , \46059 );
_DC r235e0_GF_IsGateDCbyConstraint ( \46061_nR235e0 , \46060 , \21944 );
buf \U$38609 ( \46062 , \46061_nR235e0 );
not \U$38610 ( \46063 , \46008 );
and \U$38611 ( \46064 , RIe021fe0_5038, \46063 );
not \U$38612 ( \46065 , RIe021fe0_5038);
or \U$38613 ( \46066 , \46065 , \45976 );
not \U$38614 ( \46067 , \45847 );
not \U$38615 ( \46068 , \46067 );
and \U$38616 ( \46069 , \43661 , \46068 );
not \U$38617 ( \46070 , \46069 );
not \U$38618 ( \46071 , \45944 );
or \U$38619 ( \46072 , \44899 , \46071 );
nand \U$38620 ( \46073 , \46066 , \46070 , \46072 );
and \U$38621 ( \46074 , \46073 , \46008 );
or \U$38622 ( \46075 , \46064 , \46074 );
and \U$38624 ( \46076 , \46075 , 1'b1 );
or \U$38626 ( \46077 , \46076 , 1'b0 );
buf \U$38627 ( \46078 , \46077 );
_DC r235e2_GF_IsGateDCbyConstraint ( \46079_nR235e2 , \46078 , \21944 );
buf \U$38628 ( \46080 , \46079_nR235e2 );
not \U$38629 ( \46081 , \45614 );
and \U$38630 ( \46082 , RIe020168_5039, \46081 );
not \U$38631 ( \46083 , RIe020168_5039);
or \U$38632 ( \46084 , \46083 , \45845 );
not \U$38633 ( \46085 , \45848 );
and \U$38634 ( \46086 , \43680 , \46085 );
not \U$38635 ( \46087 , \46086 );
buf \U$38636 ( \46088 , \45852 );
not \U$38637 ( \46089 , \46088 );
or \U$38638 ( \46090 , \44917 , \46089 );
nand \U$38639 ( \46091 , \46084 , \46087 , \46090 );
and \U$38640 ( \46092 , \46091 , \45614 );
or \U$38641 ( \46093 , \46082 , \46092 );
and \U$38643 ( \46094 , \46093 , 1'b1 );
or \U$38645 ( \46095 , \46094 , 1'b0 );
buf \U$38646 ( \46096 , \46095 );
_DC r235e4_GF_IsGateDCbyConstraint ( \46097_nR235e4 , \46096 , \21944 );
buf \U$38647 ( \46098 , \46097_nR235e4 );
not \U$38648 ( \46099 , \46044 );
and \U$38649 ( \46100 , RIe01dcd8_5040, \46099 );
not \U$38650 ( \46101 , RIe01dcd8_5040);
or \U$38651 ( \46102 , \46101 , \45845 );
not \U$38652 ( \46103 , \46013 );
and \U$38653 ( \46104 , \43698 , \46103 );
not \U$38654 ( \46105 , \46104 );
not \U$38655 ( \46106 , \46088 );
or \U$38656 ( \46107 , \44935 , \46106 );
nand \U$38657 ( \46108 , \46102 , \46105 , \46107 );
and \U$38658 ( \46109 , \46108 , \46044 );
or \U$38659 ( \46110 , \46100 , \46109 );
and \U$38661 ( \46111 , \46110 , 1'b1 );
or \U$38663 ( \46112 , \46111 , 1'b0 );
buf \U$38664 ( \46113 , \46112 );
_DC r235e6_GF_IsGateDCbyConstraint ( \46114_nR235e6 , \46113 , \21944 );
buf \U$38665 ( \46115 , \46114_nR235e6 );
not \U$38666 ( \46116 , \46008 );
and \U$38667 ( \46117 , RIe01b758_5041, \46116 );
not \U$38668 ( \46118 , RIe01b758_5041);
or \U$38669 ( \46119 , \46118 , \45903 );
not \U$38670 ( \46120 , \46049 );
and \U$38671 ( \46121 , \43718 , \46120 );
not \U$38672 ( \46122 , \46121 );
not \U$38673 ( \46123 , \46088 );
or \U$38674 ( \46124 , \44953 , \46123 );
nand \U$38675 ( \46125 , \46119 , \46122 , \46124 );
and \U$38676 ( \46126 , \46125 , \46008 );
or \U$38677 ( \46127 , \46117 , \46126 );
and \U$38679 ( \46128 , \46127 , 1'b1 );
or \U$38681 ( \46129 , \46128 , 1'b0 );
buf \U$38682 ( \46130 , \46129 );
_DC r235e8_GF_IsGateDCbyConstraint ( \46131_nR235e8 , \46130 , \21944 );
buf \U$38683 ( \46132 , \46131_nR235e8 );
not \U$38684 ( \46133 , \45614 );
and \U$38685 ( \46134 , RIe018440_5042, \46133 );
not \U$38686 ( \46135 , RIe018440_5042);
or \U$38687 ( \46136 , \46135 , \45921 );
not \U$38688 ( \46137 , \46067 );
and \U$38689 ( \46138 , \43738 , \46137 );
not \U$38690 ( \46139 , \46138 );
not \U$38691 ( \46140 , \45944 );
or \U$38692 ( \46141 , \44971 , \46140 );
nand \U$38693 ( \46142 , \46136 , \46139 , \46141 );
and \U$38694 ( \46143 , \46142 , \45614 );
or \U$38695 ( \46144 , \46134 , \46143 );
and \U$38697 ( \46145 , \46144 , 1'b1 );
or \U$38699 ( \46146 , \46145 , 1'b0 );
buf \U$38700 ( \46147 , \46146 );
_DC r235ea_GF_IsGateDCbyConstraint ( \46148_nR235ea , \46147 , \21944 );
buf \U$38701 ( \46149 , \46148_nR235ea );
not \U$38702 ( \46150 , \46044 );
and \U$38703 ( \46151 , RIe0157b8_5043, \46150 );
not \U$38704 ( \46152 , RIe0157b8_5043);
or \U$38705 ( \46153 , \46152 , \45921 );
not \U$38706 ( \46154 , \45959 );
and \U$38707 ( \46155 , \43756 , \46154 );
not \U$38708 ( \46156 , \46155 );
not \U$38709 ( \46157 , \45872 );
or \U$38710 ( \46158 , \44989 , \46157 );
nand \U$38711 ( \46159 , \46153 , \46156 , \46158 );
and \U$38712 ( \46160 , \46159 , \46044 );
or \U$38713 ( \46161 , \46151 , \46160 );
and \U$38715 ( \46162 , \46161 , 1'b1 );
or \U$38717 ( \46163 , \46162 , 1'b0 );
buf \U$38718 ( \46164 , \46163 );
_DC r235ec_GF_IsGateDCbyConstraint ( \46165_nR235ec , \46164 , \21944 );
buf \U$38719 ( \46166 , \46165_nR235ec );
not \U$38720 ( \46167 , \46008 );
and \U$38721 ( \46168 , RIe012590_5044, \46167 );
not \U$38722 ( \46169 , RIe012590_5044);
or \U$38723 ( \46170 , \46169 , \45903 );
not \U$38724 ( \46171 , \46049 );
and \U$38725 ( \46172 , \43776 , \46171 );
not \U$38726 ( \46173 , \46172 );
not \U$38727 ( \46174 , \46088 );
or \U$38728 ( \46175 , \45007 , \46174 );
nand \U$38729 ( \46176 , \46170 , \46173 , \46175 );
and \U$38730 ( \46177 , \46176 , \46008 );
or \U$38731 ( \46178 , \46168 , \46177 );
and \U$38733 ( \46179 , \46178 , 1'b1 );
or \U$38735 ( \46180 , \46179 , 1'b0 );
buf \U$38736 ( \46181 , \46180 );
_DC r235ee_GF_IsGateDCbyConstraint ( \46182_nR235ee , \46181 , \21944 );
buf \U$38737 ( \46183 , \46182_nR235ee );
not \U$38738 ( \46184 , \45614 );
and \U$38739 ( \46185 , RIe010628_5045, \46184 );
not \U$38740 ( \46186 , RIe010628_5045);
or \U$38741 ( \46187 , \46186 , \45845 );
not \U$38742 ( \46188 , \45959 );
and \U$38743 ( \46189 , \43795 , \46188 );
not \U$38744 ( \46190 , \46189 );
not \U$38745 ( \46191 , \45853 );
or \U$38746 ( \46192 , \45025 , \46191 );
nand \U$38747 ( \46193 , \46187 , \46190 , \46192 );
and \U$38748 ( \46194 , \46193 , \45614 );
or \U$38749 ( \46195 , \46185 , \46194 );
and \U$38751 ( \46196 , \46195 , 1'b1 );
or \U$38753 ( \46197 , \46196 , 1'b0 );
buf \U$38754 ( \46198 , \46197 );
_DC r235f0_GF_IsGateDCbyConstraint ( \46199_nR235f0 , \46198 , \21944 );
buf \U$38755 ( \46200 , \46199_nR235f0 );
not \U$38756 ( \46201 , \46044 );
and \U$38757 ( \46202 , RIe00d298_5046, \46201 );
not \U$38758 ( \46203 , RIe00d298_5046);
or \U$38759 ( \46204 , \46203 , \45903 );
not \U$38760 ( \46205 , \45940 );
and \U$38761 ( \46206 , \43813 , \46205 );
not \U$38762 ( \46207 , \46206 );
not \U$38763 ( \46208 , \45944 );
or \U$38764 ( \46209 , \45043 , \46208 );
nand \U$38765 ( \46210 , \46204 , \46207 , \46209 );
and \U$38766 ( \46211 , \46210 , \46044 );
or \U$38767 ( \46212 , \46202 , \46211 );
and \U$38769 ( \46213 , \46212 , 1'b1 );
or \U$38771 ( \46214 , \46213 , 1'b0 );
buf \U$38772 ( \46215 , \46214 );
_DC r235f4_GF_IsGateDCbyConstraint ( \46216_nR235f4 , \46215 , \21944 );
buf \U$38773 ( \46217 , \46216_nR235f4 );
not \U$38774 ( \46218 , \46008 );
and \U$38775 ( \46219 , RIe00a778_5047, \46218 );
not \U$38776 ( \46220 , RIe00a778_5047);
or \U$38777 ( \46221 , \46220 , \45903 );
not \U$38778 ( \46222 , \46013 );
and \U$38779 ( \46223 , \43832 , \46222 );
not \U$38780 ( \46224 , \46223 );
not \U$38781 ( \46225 , \46088 );
or \U$38782 ( \46226 , \45061 , \46225 );
nand \U$38783 ( \46227 , \46221 , \46224 , \46226 );
and \U$38784 ( \46228 , \46227 , \46008 );
or \U$38785 ( \46229 , \46219 , \46228 );
and \U$38787 ( \46230 , \46229 , 1'b1 );
or \U$38789 ( \46231 , \46230 , 1'b0 );
buf \U$38790 ( \46232 , \46231 );
_DC r235f6_GF_IsGateDCbyConstraint ( \46233_nR235f6 , \46232 , \21944 );
buf \U$38791 ( \46234 , \46233_nR235f6 );
buf \U$38792 ( \46235 , \43482 );
not \U$38793 ( \46236 , \46235 );
and \U$38794 ( \46237 , RIe007e38_5048, \46236 );
not \U$38795 ( \46238 , RIe007e38_5048);
or \U$38796 ( \46239 , \46238 , \45921 );
not \U$38797 ( \46240 , \45868 );
and \U$38798 ( \46241 , \43852 , \46240 );
not \U$38799 ( \46242 , \46241 );
not \U$38800 ( \46243 , \46088 );
or \U$38801 ( \46244 , \45079 , \46243 );
nand \U$38802 ( \46245 , \46239 , \46242 , \46244 );
and \U$38803 ( \46246 , \46245 , \46235 );
or \U$38804 ( \46247 , \46237 , \46246 );
and \U$38806 ( \46248 , \46247 , 1'b1 );
or \U$38808 ( \46249 , \46248 , 1'b0 );
buf \U$38809 ( \46250 , \46249 );
_DC r235f8_GF_IsGateDCbyConstraint ( \46251_nR235f8 , \46250 , \21944 );
buf \U$38810 ( \46252 , \46251_nR235f8 );
not \U$38811 ( \46253 , \46044 );
and \U$38812 ( \46254 , RIe004df0_5049, \46253 );
not \U$38813 ( \46255 , RIe004df0_5049);
or \U$38814 ( \46256 , \46255 , \45845 );
not \U$38815 ( \46257 , \45940 );
and \U$38816 ( \46258 , \43872 , \46257 );
not \U$38817 ( \46259 , \46258 );
not \U$38818 ( \46260 , \45944 );
or \U$38819 ( \46261 , \45097 , \46260 );
nand \U$38820 ( \46262 , \46256 , \46259 , \46261 );
and \U$38821 ( \46263 , \46262 , \46044 );
or \U$38822 ( \46264 , \46254 , \46263 );
and \U$38824 ( \46265 , \46264 , 1'b1 );
or \U$38826 ( \46266 , \46265 , 1'b0 );
buf \U$38827 ( \46267 , \46266 );
_DC r235fa_GF_IsGateDCbyConstraint ( \46268_nR235fa , \46267 , \21944 );
buf \U$38828 ( \46269 , \46268_nR235fa );
not \U$38829 ( \46270 , \46008 );
and \U$38830 ( \46271 , RIe0024b0_5050, \46270 );
not \U$38831 ( \46272 , RIe0024b0_5050);
or \U$38832 ( \46273 , \46272 , \45845 );
not \U$38833 ( \46274 , \46013 );
and \U$38834 ( \46275 , \43890 , \46274 );
not \U$38835 ( \46276 , \46275 );
not \U$38836 ( \46277 , \46088 );
or \U$38837 ( \46278 , \45115 , \46277 );
nand \U$38838 ( \46279 , \46273 , \46276 , \46278 );
and \U$38839 ( \46280 , \46279 , \46008 );
or \U$38840 ( \46281 , \46271 , \46280 );
and \U$38842 ( \46282 , \46281 , 1'b1 );
or \U$38844 ( \46283 , \46282 , 1'b0 );
buf \U$38845 ( \46284 , \46283 );
_DC r235fc_GF_IsGateDCbyConstraint ( \46285_nR235fc , \46284 , \21944 );
buf \U$38846 ( \46286 , \46285_nR235fc );
not \U$38847 ( \46287 , \46235 );
and \U$38848 ( \46288 , RIdfff558_5051, \46287 );
not \U$38849 ( \46289 , RIdfff558_5051);
or \U$38850 ( \46290 , \46289 , \45976 );
not \U$38851 ( \46291 , \45848 );
and \U$38852 ( \46292 , \43910 , \46291 );
not \U$38853 ( \46293 , \46292 );
not \U$38854 ( \46294 , \45872 );
or \U$38855 ( \46295 , \45133 , \46294 );
nand \U$38856 ( \46296 , \46290 , \46293 , \46295 );
and \U$38857 ( \46297 , \46296 , \46235 );
or \U$38858 ( \46298 , \46288 , \46297 );
and \U$38860 ( \46299 , \46298 , 1'b1 );
or \U$38862 ( \46300 , \46299 , 1'b0 );
buf \U$38863 ( \46301 , \46300 );
_DC r235fe_GF_IsGateDCbyConstraint ( \46302_nR235fe , \46301 , \21944 );
buf \U$38864 ( \46303 , \46302_nR235fe );
not \U$38865 ( \46304 , \46044 );
and \U$38866 ( \46305 , RIdffcd08_5052, \46304 );
not \U$38867 ( \46306 , RIdffcd08_5052);
or \U$38868 ( \46307 , \46306 , \45903 );
not \U$38869 ( \46308 , \45940 );
and \U$38870 ( \46309 , \43929 , \46308 );
not \U$38871 ( \46310 , \46309 );
not \U$38872 ( \46311 , \45853 );
or \U$38873 ( \46312 , \45151 , \46311 );
nand \U$38874 ( \46313 , \46307 , \46310 , \46312 );
and \U$38875 ( \46314 , \46313 , \46044 );
or \U$38876 ( \46315 , \46305 , \46314 );
and \U$38878 ( \46316 , \46315 , 1'b1 );
or \U$38880 ( \46317 , \46316 , 1'b0 );
buf \U$38881 ( \46318 , \46317 );
_DC r23600_GF_IsGateDCbyConstraint ( \46319_nR23600 , \46318 , \21944 );
buf \U$38882 ( \46320 , \46319_nR23600 );
not \U$38883 ( \46321 , \46008 );
and \U$38884 ( \46322 , RIdffa260_5053, \46321 );
not \U$38885 ( \46323 , RIdffa260_5053);
or \U$38886 ( \46324 , \46323 , \45921 );
not \U$38887 ( \46325 , \45868 );
and \U$38888 ( \46326 , \43949 , \46325 );
not \U$38889 ( \46327 , \46326 );
not \U$38890 ( \46328 , \45853 );
or \U$38891 ( \46329 , \45169 , \46328 );
nand \U$38892 ( \46330 , \46324 , \46327 , \46329 );
and \U$38893 ( \46331 , \46330 , \46008 );
or \U$38894 ( \46332 , \46322 , \46331 );
and \U$38896 ( \46333 , \46332 , 1'b1 );
or \U$38898 ( \46334 , \46333 , 1'b0 );
buf \U$38899 ( \46335 , \46334 );
_DC r23602_GF_IsGateDCbyConstraint ( \46336_nR23602 , \46335 , \21944 );
buf \U$38900 ( \46337 , \46336_nR23602 );
not \U$38901 ( \46338 , \46235 );
and \U$38902 ( \46339 , RIdff7b78_5054, \46338 );
not \U$38903 ( \46340 , RIdff7b78_5054);
or \U$38904 ( \46341 , \46340 , \45903 );
not \U$38905 ( \46342 , \46067 );
and \U$38906 ( \46343 , \43969 , \46342 );
not \U$38907 ( \46344 , \46343 );
not \U$38908 ( \46345 , \45853 );
or \U$38909 ( \46346 , \45187 , \46345 );
nand \U$38910 ( \46347 , \46341 , \46344 , \46346 );
and \U$38911 ( \46348 , \46347 , \46235 );
or \U$38912 ( \46349 , \46339 , \46348 );
and \U$38914 ( \46350 , \46349 , 1'b1 );
or \U$38916 ( \46351 , \46350 , 1'b0 );
buf \U$38917 ( \46352 , \46351 );
_DC r23604_GF_IsGateDCbyConstraint ( \46353_nR23604 , \46352 , \21944 );
buf \U$38918 ( \46354 , \46353_nR23604 );
not \U$38919 ( \46355 , \46044 );
and \U$38920 ( \46356 , RIdff4f68_5055, \46355 );
not \U$38921 ( \46357 , RIdff4f68_5055);
or \U$38922 ( \46358 , \46357 , \45976 );
not \U$38923 ( \46359 , \46013 );
and \U$38924 ( \46360 , \43987 , \46359 );
not \U$38925 ( \46361 , \46360 );
not \U$38926 ( \46362 , \46088 );
or \U$38927 ( \46363 , \45205 , \46362 );
nand \U$38928 ( \46364 , \46358 , \46361 , \46363 );
and \U$38929 ( \46365 , \46364 , \46044 );
or \U$38930 ( \46366 , \46356 , \46365 );
and \U$38932 ( \46367 , \46366 , 1'b1 );
or \U$38934 ( \46368 , \46367 , 1'b0 );
buf \U$38935 ( \46369 , \46368 );
_DC r23606_GF_IsGateDCbyConstraint ( \46370_nR23606 , \46369 , \21944 );
buf \U$38936 ( \46371 , \46370_nR23606 );
not \U$38937 ( \46372 , \46008 );
and \U$38938 ( \46373 , RIdff1ea8_5056, \46372 );
not \U$38939 ( \46374 , RIdff1ea8_5056);
or \U$38940 ( \46375 , \46374 , \45845 );
not \U$38941 ( \46376 , \46013 );
and \U$38942 ( \46377 , \44006 , \46376 );
not \U$38943 ( \46378 , \46377 );
not \U$38944 ( \46379 , \46088 );
or \U$38945 ( \46380 , \45223 , \46379 );
nand \U$38946 ( \46381 , \46375 , \46378 , \46380 );
and \U$38947 ( \46382 , \46381 , \46008 );
or \U$38948 ( \46383 , \46373 , \46382 );
and \U$38950 ( \46384 , \46383 , 1'b1 );
or \U$38952 ( \46385 , \46384 , 1'b0 );
buf \U$38953 ( \46386 , \46385 );
_DC r2360a_GF_IsGateDCbyConstraint ( \46387_nR2360a , \46386 , \21944 );
buf \U$38954 ( \46388 , \46387_nR2360a );
endmodule

