//
// Conformal-LEC Version 20.10-d132 (30-Jun-2020)
//
module top(RI2af433cd5b80_17,RI2af433cd5b08_16,RI2af433cd5a90_15,RI2af433cd5a18_14,RI2af433cd59a0_13,RI2af433cd5928_12,RI2af433cd58b0_11,RI2af433cd5838_10,RI2af433cd57c0_9,
        RI2af433cd5748_8,RI2af433cd56d0_7,RI2af433cd5658_6,RI2af433cd5bf8_18,RI2af433cd5c70_19,RI2af433cd5ce8_20,RI2af433cd5d60_21,RI2af433cd5dd8_22,RI2af433cd5e50_23,RI2af433cd5ec8_24,
        RI2af433cd5f40_25,RI2af433cd5fb8_26,RI2af433cd6030_27,RI2af433cd60a8_28,RI2af433cd6120_29,RI2af433cd6198_30,RI2af433cd6210_31,RI2af433cd6288_32,RI2af433cd6300_33,RI2af433cd6378_34,
        RI2af433cd63f0_35,RI2af433cd6468_36,RI2af433cd64e0_37,RI2af433cd6558_38,RI2af433cd65d0_39,RI2af433cd6648_40,RI2af433cd66c0_41,RI2af433cd6738_42,RI2af433cd67b0_43,RI2af433cd6828_44,
        RI2af433cd68a0_45,RI2af433cd6918_46,RI2af433cd6990_47,RI2af433cd6a08_48,RI2af433cd6a80_49,RI2af433cd6af8_50,RI2af433cd6b70_51,RI2af433cd6be8_52,RI2af433cd6c60_53,RI2af433cd6cd8_54,
        RI2af433cd6d50_55,RI2af433cd6dc8_56,RI2af433cd6e40_57,RI2af433cd6eb8_58,RI2af433cd6f30_59,RI2af433cd6fa8_60,RI2af433cd7020_61,RI2af433cd7098_62,RI2af433cd7110_63,RI2af433cd7188_64,
        RI2af433cd7200_65,RI2af433cd7278_66,RI2af433cd72f0_67,RI2af433cd7368_68,RI2af433cd73e0_69,RI2af433cd7458_70,RI2af433cd74d0_71,RI2af433cd7548_72,RI2af433cd75c0_73,RI2af433cd7638_74,
        RI2af433cd76b0_75,RI2af433cd7728_76,RI2af433cd77a0_77,RI2af433cd7818_78,RI2af433cd7890_79,RI2af433cd7908_80,RI2af433cd7980_81,RI2af433cd79f8_82,RI2af433cd7a70_83,RI2af433cd7ae8_84,
        RI2af433cd7b60_85,RI2af433cd7bd8_86,RI2af433cd7c50_87,RI2af433cd7cc8_88,RI2af433cd7d40_89,RI2af433cd7db8_90,RI2af433cd7e30_91,RI2af433cd7ea8_92,RI2af433cd7f20_93,RI2af433cd7f98_94,
        RI2af433cd8010_95,RI2af433cd8088_96,RI2af433cd8100_97,RI2af433cd8178_98,RI2af433cd81f0_99,RI2af433cd8268_100,RI2af433cd82e0_101,RI2af433cd8358_102,RI2af433cd83d0_103,RI2af433cd8448_104,
        RI2af433cd84c0_105,RI2af433cd8538_106,RI2af433cd85b0_107,RI2af433cd8628_108,RI2af433cd86a0_109,RI2af433cd8718_110,RI2af433cd8790_111,RI2af433cd8808_112,RI2af433cd8880_113,RI2af433cd88f8_114,
        RI2af433cd8970_115,RI2af433cd89e8_116,RI2af433cd8a60_117,RI2af433cd8ad8_118,RI2af433cd8b50_119,RI2af433cd8bc8_120,RI2af433cd8c40_121,RI2af433cd8cb8_122,RI2af433cd8d30_123,RI2af433cd8da8_124,
        RI2af433cd8e20_125,RI2af433cd8e98_126,RI2af433cd8f10_127,RI2af433cd8f88_128,RI2af433cd9000_129,RI2af433cd9078_130,RI2af433cd90f0_131,RI2af433cd9168_132,RI2af433cd91e0_133,RI2af433cd9258_134,
        RI2af433cd92d0_135,RI2af433cd9348_136,RI2af433cd93c0_137,RI2af433cd9438_138,RI2af433cd94b0_139,RI2af433cd9528_140,RI2af433cd95a0_141,RI2af433cd9618_142,RI2af433cd9690_143,RI2af433cd9708_144,
        RI2af433cd9780_145,RI2af433cd97f8_146,RI2af433cd9870_147,RI2af433cd98e8_148,RI2af433cd9960_149,RI2af433cd99d8_150,RI2af433cd9a50_151,RI2af433cd9ac8_152,RI2af433cd9b40_153,RI2af433cd9bb8_154,
        RI2af433cd9c30_155,RI2af433cd9ca8_156,RI2af433cd9d20_157,RI2af433cd9d98_158,RI2af433cd9e10_159,RI2af433cd9e88_160,RI2af433cd9f00_161,RI2af433cd9f78_162,RI2af433cd9ff0_163,RI2af433cda068_164,
        RI2af433cda0e0_165,RI2af433cda158_166,RI2af433cda1d0_167,RI2af433cda248_168,RI2af433cda2c0_169,RI2af433cda338_170,RI2af433cda3b0_171,RI2af433cda428_172,RI2af433cda4a0_173,RI2af433cda518_174,
        RI2af433cda590_175,RI2af433cda608_176,RI2af433cda680_177,RI2af433cda6f8_178,RI2af433cda770_179,RI2af433cda7e8_180,RI2af433cda860_181,RI2af433cda8d8_182,RI2af433cda950_183,RI2af433cda9c8_184,
        RI2af433cdaa40_185,RI2af433cdaab8_186,RI2af433cdab30_187,RI2af433cdaba8_188,RI2af433cdac20_189,RI2af433cdac98_190,RI2af433cdad10_191,RI2af433cdad88_192,RI2af433cdae00_193,RI2af433cdae78_194,
        RI2af433cdaef0_195,RI2af433cdaf68_196,RI2af433cdafe0_197,RI2af433cdb058_198,RI2af433cdb0d0_199,RI2af433cdb148_200,RI2af433cdb1c0_201,RI2af433cdb238_202,RI2af433cdb2b0_203,RI2af433cdb328_204,
        RI2af433cdb3a0_205,RI2af433cdb418_206,RI2af433cdb490_207,RI2af433cdb508_208,RI2af433cdb580_209,RI2af433cdb5f8_210,RI2af433cdb670_211,RI2af433cdb6e8_212,RI2af433cdb760_213,RI2af433cdb7d8_214,
        RI2af433cdb850_215,RI2af433cdb8c8_216,RI2af433cdb940_217,RI2af433cc8a70_1,RI2af433cd5478_2,RI2af433cd54f0_3,RI2af433cd5568_4,RI2af433cd55e0_5,R_da_9022e98,R_db_9022f40);
input RI2af433cd5b80_17,RI2af433cd5b08_16,RI2af433cd5a90_15,RI2af433cd5a18_14,RI2af433cd59a0_13,RI2af433cd5928_12,RI2af433cd58b0_11,RI2af433cd5838_10,RI2af433cd57c0_9,
        RI2af433cd5748_8,RI2af433cd56d0_7,RI2af433cd5658_6,RI2af433cd5bf8_18,RI2af433cd5c70_19,RI2af433cd5ce8_20,RI2af433cd5d60_21,RI2af433cd5dd8_22,RI2af433cd5e50_23,RI2af433cd5ec8_24,
        RI2af433cd5f40_25,RI2af433cd5fb8_26,RI2af433cd6030_27,RI2af433cd60a8_28,RI2af433cd6120_29,RI2af433cd6198_30,RI2af433cd6210_31,RI2af433cd6288_32,RI2af433cd6300_33,RI2af433cd6378_34,
        RI2af433cd63f0_35,RI2af433cd6468_36,RI2af433cd64e0_37,RI2af433cd6558_38,RI2af433cd65d0_39,RI2af433cd6648_40,RI2af433cd66c0_41,RI2af433cd6738_42,RI2af433cd67b0_43,RI2af433cd6828_44,
        RI2af433cd68a0_45,RI2af433cd6918_46,RI2af433cd6990_47,RI2af433cd6a08_48,RI2af433cd6a80_49,RI2af433cd6af8_50,RI2af433cd6b70_51,RI2af433cd6be8_52,RI2af433cd6c60_53,RI2af433cd6cd8_54,
        RI2af433cd6d50_55,RI2af433cd6dc8_56,RI2af433cd6e40_57,RI2af433cd6eb8_58,RI2af433cd6f30_59,RI2af433cd6fa8_60,RI2af433cd7020_61,RI2af433cd7098_62,RI2af433cd7110_63,RI2af433cd7188_64,
        RI2af433cd7200_65,RI2af433cd7278_66,RI2af433cd72f0_67,RI2af433cd7368_68,RI2af433cd73e0_69,RI2af433cd7458_70,RI2af433cd74d0_71,RI2af433cd7548_72,RI2af433cd75c0_73,RI2af433cd7638_74,
        RI2af433cd76b0_75,RI2af433cd7728_76,RI2af433cd77a0_77,RI2af433cd7818_78,RI2af433cd7890_79,RI2af433cd7908_80,RI2af433cd7980_81,RI2af433cd79f8_82,RI2af433cd7a70_83,RI2af433cd7ae8_84,
        RI2af433cd7b60_85,RI2af433cd7bd8_86,RI2af433cd7c50_87,RI2af433cd7cc8_88,RI2af433cd7d40_89,RI2af433cd7db8_90,RI2af433cd7e30_91,RI2af433cd7ea8_92,RI2af433cd7f20_93,RI2af433cd7f98_94,
        RI2af433cd8010_95,RI2af433cd8088_96,RI2af433cd8100_97,RI2af433cd8178_98,RI2af433cd81f0_99,RI2af433cd8268_100,RI2af433cd82e0_101,RI2af433cd8358_102,RI2af433cd83d0_103,RI2af433cd8448_104,
        RI2af433cd84c0_105,RI2af433cd8538_106,RI2af433cd85b0_107,RI2af433cd8628_108,RI2af433cd86a0_109,RI2af433cd8718_110,RI2af433cd8790_111,RI2af433cd8808_112,RI2af433cd8880_113,RI2af433cd88f8_114,
        RI2af433cd8970_115,RI2af433cd89e8_116,RI2af433cd8a60_117,RI2af433cd8ad8_118,RI2af433cd8b50_119,RI2af433cd8bc8_120,RI2af433cd8c40_121,RI2af433cd8cb8_122,RI2af433cd8d30_123,RI2af433cd8da8_124,
        RI2af433cd8e20_125,RI2af433cd8e98_126,RI2af433cd8f10_127,RI2af433cd8f88_128,RI2af433cd9000_129,RI2af433cd9078_130,RI2af433cd90f0_131,RI2af433cd9168_132,RI2af433cd91e0_133,RI2af433cd9258_134,
        RI2af433cd92d0_135,RI2af433cd9348_136,RI2af433cd93c0_137,RI2af433cd9438_138,RI2af433cd94b0_139,RI2af433cd9528_140,RI2af433cd95a0_141,RI2af433cd9618_142,RI2af433cd9690_143,RI2af433cd9708_144,
        RI2af433cd9780_145,RI2af433cd97f8_146,RI2af433cd9870_147,RI2af433cd98e8_148,RI2af433cd9960_149,RI2af433cd99d8_150,RI2af433cd9a50_151,RI2af433cd9ac8_152,RI2af433cd9b40_153,RI2af433cd9bb8_154,
        RI2af433cd9c30_155,RI2af433cd9ca8_156,RI2af433cd9d20_157,RI2af433cd9d98_158,RI2af433cd9e10_159,RI2af433cd9e88_160,RI2af433cd9f00_161,RI2af433cd9f78_162,RI2af433cd9ff0_163,RI2af433cda068_164,
        RI2af433cda0e0_165,RI2af433cda158_166,RI2af433cda1d0_167,RI2af433cda248_168,RI2af433cda2c0_169,RI2af433cda338_170,RI2af433cda3b0_171,RI2af433cda428_172,RI2af433cda4a0_173,RI2af433cda518_174,
        RI2af433cda590_175,RI2af433cda608_176,RI2af433cda680_177,RI2af433cda6f8_178,RI2af433cda770_179,RI2af433cda7e8_180,RI2af433cda860_181,RI2af433cda8d8_182,RI2af433cda950_183,RI2af433cda9c8_184,
        RI2af433cdaa40_185,RI2af433cdaab8_186,RI2af433cdab30_187,RI2af433cdaba8_188,RI2af433cdac20_189,RI2af433cdac98_190,RI2af433cdad10_191,RI2af433cdad88_192,RI2af433cdae00_193,RI2af433cdae78_194,
        RI2af433cdaef0_195,RI2af433cdaf68_196,RI2af433cdafe0_197,RI2af433cdb058_198,RI2af433cdb0d0_199,RI2af433cdb148_200,RI2af433cdb1c0_201,RI2af433cdb238_202,RI2af433cdb2b0_203,RI2af433cdb328_204,
        RI2af433cdb3a0_205,RI2af433cdb418_206,RI2af433cdb490_207,RI2af433cdb508_208,RI2af433cdb580_209,RI2af433cdb5f8_210,RI2af433cdb670_211,RI2af433cdb6e8_212,RI2af433cdb760_213,RI2af433cdb7d8_214,
        RI2af433cdb850_215,RI2af433cdb8c8_216,RI2af433cdb940_217,RI2af433cc8a70_1,RI2af433cd5478_2,RI2af433cd54f0_3,RI2af433cd5568_4,RI2af433cd55e0_5;
output R_da_9022e98,R_db_9022f40;

wire \220 , \221_N$2 , \222_ZERO , \223 , \224_N$1 , \225_ONE , \226 , \227 , \228 ,
         \229 , \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 , \238 ,
         \239 , \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 , \248 ,
         \249 , \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 , \258 ,
         \259 , \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 , \268 ,
         \269 , \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 , \278 ,
         \279 , \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 , \288 ,
         \289 , \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 , \298 ,
         \299 , \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 , \308 ,
         \309 , \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 , \318 ,
         \319 , \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 , \328 ,
         \329 , \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 , \338 ,
         \339 , \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 , \348 ,
         \349 , \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 ,
         \359 , \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 ,
         \369 , \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 ,
         \379 , \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 ,
         \389 , \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 ,
         \399 , \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 ,
         \409 , \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 ,
         \419 , \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 ,
         \429 , \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 ,
         \439 , \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 ,
         \449 , \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 ,
         \459 , \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 ,
         \469 , \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 ,
         \479 , \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 ,
         \489 , \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 ,
         \499 , \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 ,
         \509 , \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 ,
         \519 , \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 ,
         \529 , \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 ,
         \539 , \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 ,
         \549 , \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 ,
         \559 , \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 ,
         \569 , \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 ,
         \579 , \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 ,
         \589 , \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 ,
         \599 , \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 ,
         \609 , \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 ,
         \619 , \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 ,
         \629 , \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 ,
         \639 , \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 ,
         \649 , \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658_nR372 ,
         \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 ,
         \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 ,
         \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 ,
         \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 ,
         \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 ,
         \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 ,
         \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 ,
         \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 ,
         \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 ,
         \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 ,
         \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 ,
         \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 ,
         \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 ,
         \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 ,
         \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 ,
         \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 ,
         \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 ,
         \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 ,
         \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 ,
         \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 ,
         \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 ,
         \869 , \870 , \871 , \872 , \873 , \874 , \875_nR1bf , \876 , \877 , \878 ;
buf \U$labaj116 ( R_da_9022e98, \659 );
buf \U$labaj117 ( R_db_9022f40, \878 );
not \U$1 ( \226 , RI2af433cd59a0_13);
not \U$2 ( \227 , RI2af433cd5838_10);
not \U$3 ( \228 , RI2af433cd57c0_9);
nor \U$4 ( \229 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$5 ( \230 , RI2af433cd5b80_17, \229 );
not \U$6 ( \231 , RI2af433cd5b08_16);
not \U$7 ( \232 , RI2af433cd5a90_15);
not \U$8 ( \233 , RI2af433cd5a18_14);
nor \U$9 ( \234 , \231 , \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$10 ( \235 , RI2af433cd5bf8_18, \234 );
nor \U$11 ( \236 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$12 ( \237 , RI2af433cd5c70_19, \236 );
nor \U$13 ( \238 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$14 ( \239 , RI2af433cd5ce8_20, \238 );
nor \U$15 ( \240 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$16 ( \241 , RI2af433cd5d60_21, \240 );
nor \U$17 ( \242 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$18 ( \243 , RI2af433cd5dd8_22, \242 );
nor \U$19 ( \244 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$20 ( \245 , RI2af433cd5e50_23, \244 );
nor \U$21 ( \246 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$22 ( \247 , RI2af433cd5ec8_24, \246 );
nor \U$23 ( \248 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$24 ( \249 , RI2af433cd5f40_25, \248 );
not \U$25 ( \250 , RI2af433cd5928_12);
not \U$26 ( \251 , RI2af433cd58b0_11);
nor \U$27 ( \252 , \231 , \232 , \233 , \226 , \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$28 ( \253 , RI2af433cd5fb8_26, \252 );
nor \U$29 ( \254 , RI2af433cd5b08_16, \232 , \233 , \226 , \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$30 ( \255 , RI2af433cd6030_27, \254 );
nor \U$31 ( \256 , \231 , RI2af433cd5a90_15, \233 , \226 , \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$32 ( \257 , RI2af433cd60a8_28, \256 );
nor \U$33 ( \258 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$34 ( \259 , RI2af433cd6120_29, \258 );
nor \U$35 ( \260 , \231 , \232 , RI2af433cd5a18_14, \226 , \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$36 ( \261 , RI2af433cd6198_30, \260 );
nor \U$37 ( \262 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$38 ( \263 , RI2af433cd6210_31, \262 );
nor \U$39 ( \264 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$40 ( \265 , RI2af433cd6288_32, \264 );
nor \U$41 ( \266 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$42 ( \267 , RI2af433cd6300_33, \266 );
nor \U$43 ( \268 , \231 , \232 , \233 , RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$44 ( \269 , RI2af433cd6378_34, \268 );
nor \U$45 ( \270 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$46 ( \271 , RI2af433cd63f0_35, \270 );
nor \U$47 ( \272 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$48 ( \273 , RI2af433cd6468_36, \272 );
nor \U$49 ( \274 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$50 ( \275 , RI2af433cd64e0_37, \274 );
nor \U$51 ( \276 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$52 ( \277 , RI2af433cd6558_38, \276 );
nor \U$53 ( \278 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$54 ( \279 , RI2af433cd65d0_39, \278 );
nor \U$55 ( \280 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$56 ( \281 , RI2af433cd6648_40, \280 );
nor \U$57 ( \282 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$58 ( \283 , RI2af433cd66c0_41, \282 );
nor \U$59 ( \284 , \231 , \232 , \233 , \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$60 ( \285 , RI2af433cd6738_42, \284 );
nor \U$61 ( \286 , RI2af433cd5b08_16, \232 , \233 , \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$62 ( \287 , RI2af433cd67b0_43, \286 );
nor \U$63 ( \288 , \231 , RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$64 ( \289 , RI2af433cd6828_44, \288 );
nor \U$65 ( \290 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$66 ( \291 , RI2af433cd68a0_45, \290 );
nor \U$67 ( \292 , \231 , \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$68 ( \293 , RI2af433cd6918_46, \292 );
nor \U$69 ( \294 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$70 ( \295 , RI2af433cd6990_47, \294 );
nor \U$71 ( \296 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$72 ( \297 , RI2af433cd6a08_48, \296 );
nor \U$73 ( \298 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$74 ( \299 , RI2af433cd6a80_49, \298 );
nor \U$75 ( \300 , \231 , \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$76 ( \301 , RI2af433cd6af8_50, \300 );
nor \U$77 ( \302 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$78 ( \303 , RI2af433cd6b70_51, \302 );
nor \U$79 ( \304 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$80 ( \305 , RI2af433cd6be8_52, \304 );
nor \U$81 ( \306 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$82 ( \307 , RI2af433cd6c60_53, \306 );
nor \U$83 ( \308 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$84 ( \309 , RI2af433cd6cd8_54, \308 );
nor \U$85 ( \310 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$86 ( \311 , RI2af433cd6d50_55, \310 );
nor \U$87 ( \312 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$88 ( \313 , RI2af433cd6dc8_56, \312 );
nor \U$89 ( \314 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$90 ( \315 , RI2af433cd6e40_57, \314 );
nor \U$91 ( \316 , \231 , \232 , \233 , \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$92 ( \317 , RI2af433cd6eb8_58, \316 );
nor \U$93 ( \318 , RI2af433cd5b08_16, \232 , \233 , \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$94 ( \319 , RI2af433cd6f30_59, \318 );
nor \U$95 ( \320 , \231 , RI2af433cd5a90_15, \233 , \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$96 ( \321 , RI2af433cd6fa8_60, \320 );
nor \U$97 ( \322 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$98 ( \323 , RI2af433cd7020_61, \322 );
nor \U$99 ( \324 , \231 , \232 , RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$100 ( \325 , RI2af433cd7098_62, \324 );
nor \U$101 ( \326 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$102 ( \327 , RI2af433cd7110_63, \326 );
nor \U$103 ( \328 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$104 ( \329 , RI2af433cd7188_64, \328 );
nor \U$105 ( \330 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$106 ( \331 , RI2af433cd7200_65, \330 );
nor \U$107 ( \332 , \231 , \232 , \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$108 ( \333 , RI2af433cd7278_66, \332 );
nor \U$109 ( \334 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$110 ( \335 , RI2af433cd72f0_67, \334 );
nor \U$111 ( \336 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$112 ( \337 , RI2af433cd7368_68, \336 );
nor \U$113 ( \338 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$114 ( \339 , RI2af433cd73e0_69, \338 );
nor \U$115 ( \340 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$116 ( \341 , RI2af433cd7458_70, \340 );
nor \U$117 ( \342 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$118 ( \343 , RI2af433cd74d0_71, \342 );
nor \U$119 ( \344 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$120 ( \345 , RI2af433cd7548_72, \344 );
nor \U$121 ( \346 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$122 ( \347 , RI2af433cd75c0_73, \346 );
nor \U$123 ( \348 , \231 , \232 , \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$124 ( \349 , RI2af433cd7638_74, \348 );
nor \U$125 ( \350 , RI2af433cd5b08_16, \232 , \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$126 ( \351 , RI2af433cd76b0_75, \350 );
nor \U$127 ( \352 , \231 , RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$128 ( \353 , RI2af433cd7728_76, \352 );
nor \U$129 ( \354 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$130 ( \355 , RI2af433cd77a0_77, \354 );
nor \U$131 ( \356 , \231 , \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$132 ( \357 , RI2af433cd7818_78, \356 );
nor \U$133 ( \358 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$134 ( \359 , RI2af433cd7890_79, \358 );
nor \U$135 ( \360 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$136 ( \361 , RI2af433cd7908_80, \360 );
or \U$137 ( \362 , \230 , \235 , \237 , \239 , \241 , \243 , \245 , \247 , \249 , \253 , \255 , \257 , \259 , \261 , \263 , \265 , \267 , \269 , \271 , \273 , \275 , \277 , \279 , \281 , \283 , \285 , \287 , \289 , \291 , \293 , \295 , \297 , \299 , \301 , \303 , \305 , \307 , \309 , \311 , \313 , \315 , \317 , \319 , \321 , \323 , \325 , \327 , \329 , \331 , \333 , \335 , \337 , \339 , \341 , \343 , \345 , \347 , \349 , \351 , \353 , \355 , \357 , \359 , \361 );
nor \U$138 ( \363 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$139 ( \364 , RI2af433cd7980_81, \363 );
nor \U$140 ( \365 , \231 , \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$141 ( \366 , RI2af433cd79f8_82, \365 );
nor \U$142 ( \367 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$143 ( \368 , RI2af433cd7a70_83, \367 );
nor \U$144 ( \369 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$145 ( \370 , RI2af433cd7ae8_84, \369 );
nor \U$146 ( \371 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$147 ( \372 , RI2af433cd7b60_85, \371 );
nor \U$148 ( \373 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$149 ( \374 , RI2af433cd7bd8_86, \373 );
nor \U$150 ( \375 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$151 ( \376 , RI2af433cd7c50_87, \375 );
nor \U$152 ( \377 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$153 ( \378 , RI2af433cd7cc8_88, \377 );
nor \U$154 ( \379 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, \228 , RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$155 ( \380 , RI2af433cd7d40_89, \379 );
nor \U$156 ( \381 , \231 , \232 , \233 , \226 , \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$157 ( \382 , RI2af433cd7db8_90, \381 );
nor \U$158 ( \383 , RI2af433cd5b08_16, \232 , \233 , \226 , \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$159 ( \384 , RI2af433cd7e30_91, \383 );
nor \U$160 ( \385 , \231 , RI2af433cd5a90_15, \233 , \226 , \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$161 ( \386 , RI2af433cd7ea8_92, \385 );
nor \U$162 ( \387 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$163 ( \388 , RI2af433cd7f20_93, \387 );
nor \U$164 ( \389 , \231 , \232 , RI2af433cd5a18_14, \226 , \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$165 ( \390 , RI2af433cd7f98_94, \389 );
nor \U$166 ( \391 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$167 ( \392 , RI2af433cd8010_95, \391 );
nor \U$168 ( \393 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$169 ( \394 , RI2af433cd8088_96, \393 );
nor \U$170 ( \395 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$171 ( \396 , RI2af433cd8100_97, \395 );
nor \U$172 ( \397 , \231 , \232 , \233 , RI2af433cd59a0_13, \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$173 ( \398 , RI2af433cd8178_98, \397 );
nor \U$174 ( \399 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$175 ( \400 , RI2af433cd81f0_99, \399 );
nor \U$176 ( \401 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$177 ( \402 , RI2af433cd8268_100, \401 );
nor \U$178 ( \403 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$179 ( \404 , RI2af433cd82e0_101, \403 );
nor \U$180 ( \405 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$181 ( \406 , RI2af433cd8358_102, \405 );
nor \U$182 ( \407 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$183 ( \408 , RI2af433cd83d0_103, \407 );
nor \U$184 ( \409 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$185 ( \410 , RI2af433cd8448_104, \409 );
nor \U$186 ( \411 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$187 ( \412 , RI2af433cd84c0_105, \411 );
nor \U$188 ( \413 , \231 , \232 , \233 , \226 , RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$189 ( \414 , RI2af433cd8538_106, \413 );
nor \U$190 ( \415 , RI2af433cd5b08_16, \232 , \233 , \226 , RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$191 ( \416 , RI2af433cd85b0_107, \415 );
nor \U$192 ( \417 , \231 , RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$193 ( \418 , RI2af433cd8628_108, \417 );
nor \U$194 ( \419 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$195 ( \420 , RI2af433cd86a0_109, \419 );
nor \U$196 ( \421 , \231 , \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$197 ( \422 , RI2af433cd8718_110, \421 );
nor \U$198 ( \423 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$199 ( \424 , RI2af433cd8790_111, \423 );
nor \U$200 ( \425 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$201 ( \426 , RI2af433cd8808_112, \425 );
nor \U$202 ( \427 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$203 ( \428 , RI2af433cd8880_113, \427 );
nor \U$204 ( \429 , \231 , \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$205 ( \430 , RI2af433cd88f8_114, \429 );
nor \U$206 ( \431 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$207 ( \432 , RI2af433cd8970_115, \431 );
nor \U$208 ( \433 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$209 ( \434 , RI2af433cd89e8_116, \433 );
nor \U$210 ( \435 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$211 ( \436 , RI2af433cd8a60_117, \435 );
nor \U$212 ( \437 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$213 ( \438 , RI2af433cd8ad8_118, \437 );
nor \U$214 ( \439 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$215 ( \440 , RI2af433cd8b50_119, \439 );
nor \U$216 ( \441 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$217 ( \442 , RI2af433cd8bc8_120, \441 );
nor \U$218 ( \443 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$219 ( \444 , RI2af433cd8c40_121, \443 );
nor \U$220 ( \445 , \231 , \232 , \233 , \226 , \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$221 ( \446 , RI2af433cd8cb8_122, \445 );
nor \U$222 ( \447 , RI2af433cd5b08_16, \232 , \233 , \226 , \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$223 ( \448 , RI2af433cd8d30_123, \447 );
nor \U$224 ( \449 , \231 , RI2af433cd5a90_15, \233 , \226 , \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$225 ( \450 , RI2af433cd8da8_124, \449 );
nor \U$226 ( \451 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$227 ( \452 , RI2af433cd8e20_125, \451 );
nor \U$228 ( \453 , \231 , \232 , RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$229 ( \454 , RI2af433cd8e98_126, \453 );
nor \U$230 ( \455 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$231 ( \456 , RI2af433cd8f10_127, \455 );
nor \U$232 ( \457 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$233 ( \458 , RI2af433cd8f88_128, \457 );
nor \U$234 ( \459 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$235 ( \460 , RI2af433cd9000_129, \459 );
nor \U$236 ( \461 , \231 , \232 , \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$237 ( \462 , RI2af433cd9078_130, \461 );
nor \U$238 ( \463 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$239 ( \464 , RI2af433cd90f0_131, \463 );
nor \U$240 ( \465 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$241 ( \466 , RI2af433cd9168_132, \465 );
nor \U$242 ( \467 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$243 ( \468 , RI2af433cd91e0_133, \467 );
nor \U$244 ( \469 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$245 ( \470 , RI2af433cd9258_134, \469 );
nor \U$246 ( \471 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$247 ( \472 , RI2af433cd92d0_135, \471 );
nor \U$248 ( \473 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$249 ( \474 , RI2af433cd9348_136, \473 );
nor \U$250 ( \475 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$251 ( \476 , RI2af433cd93c0_137, \475 );
nor \U$252 ( \477 , \231 , \232 , \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$253 ( \478 , RI2af433cd9438_138, \477 );
nor \U$254 ( \479 , RI2af433cd5b08_16, \232 , \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$255 ( \480 , RI2af433cd94b0_139, \479 );
nor \U$256 ( \481 , \231 , RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$257 ( \482 , RI2af433cd9528_140, \481 );
nor \U$258 ( \483 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$259 ( \484 , RI2af433cd95a0_141, \483 );
nor \U$260 ( \485 , \231 , \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$261 ( \486 , RI2af433cd9618_142, \485 );
nor \U$262 ( \487 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$263 ( \488 , RI2af433cd9690_143, \487 );
nor \U$264 ( \489 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$265 ( \490 , RI2af433cd9708_144, \489 );
or \U$266 ( \491 , \364 , \366 , \368 , \370 , \372 , \374 , \376 , \378 , \380 , \382 , \384 , \386 , \388 , \390 , \392 , \394 , \396 , \398 , \400 , \402 , \404 , \406 , \408 , \410 , \412 , \414 , \416 , \418 , \420 , \422 , \424 , \426 , \428 , \430 , \432 , \434 , \436 , \438 , \440 , \442 , \444 , \446 , \448 , \450 , \452 , \454 , \456 , \458 , \460 , \462 , \464 , \466 , \468 , \470 , \472 , \474 , \476 , \478 , \480 , \482 , \484 , \486 , \488 , \490 );
nor \U$267 ( \492 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$268 ( \493 , RI2af433cd9780_145, \492 );
nor \U$269 ( \494 , \231 , \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$270 ( \495 , RI2af433cd97f8_146, \494 );
nor \U$271 ( \496 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$272 ( \497 , RI2af433cd9870_147, \496 );
nor \U$273 ( \498 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$274 ( \499 , RI2af433cd98e8_148, \498 );
nor \U$275 ( \500 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$276 ( \501 , RI2af433cd9960_149, \500 );
nor \U$277 ( \502 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$278 ( \503 , RI2af433cd99d8_150, \502 );
nor \U$279 ( \504 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$280 ( \505 , RI2af433cd9a50_151, \504 );
nor \U$281 ( \506 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$282 ( \507 , RI2af433cd9ac8_152, \506 );
nor \U$283 ( \508 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, \227 , RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$284 ( \509 , RI2af433cd9b40_153, \508 );
nor \U$285 ( \510 , \231 , \232 , \233 , \226 , \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$286 ( \511 , RI2af433cd9bb8_154, \510 );
nor \U$287 ( \512 , RI2af433cd5b08_16, \232 , \233 , \226 , \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$288 ( \513 , RI2af433cd9c30_155, \512 );
nor \U$289 ( \514 , \231 , RI2af433cd5a90_15, \233 , \226 , \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$290 ( \515 , RI2af433cd9ca8_156, \514 );
nor \U$291 ( \516 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$292 ( \517 , RI2af433cd9d20_157, \516 );
nor \U$293 ( \518 , \231 , \232 , RI2af433cd5a18_14, \226 , \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$294 ( \519 , RI2af433cd9d98_158, \518 );
nor \U$295 ( \520 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$296 ( \521 , RI2af433cd9e10_159, \520 );
nor \U$297 ( \522 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$298 ( \523 , RI2af433cd9e88_160, \522 );
nor \U$299 ( \524 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$300 ( \525 , RI2af433cd9f00_161, \524 );
nor \U$301 ( \526 , \231 , \232 , \233 , RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$302 ( \527 , RI2af433cd9f78_162, \526 );
nor \U$303 ( \528 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$304 ( \529 , RI2af433cd9ff0_163, \528 );
nor \U$305 ( \530 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$306 ( \531 , RI2af433cda068_164, \530 );
nor \U$307 ( \532 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$308 ( \533 , RI2af433cda0e0_165, \532 );
nor \U$309 ( \534 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$310 ( \535 , RI2af433cda158_166, \534 );
nor \U$311 ( \536 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$312 ( \537 , RI2af433cda1d0_167, \536 );
nor \U$313 ( \538 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$314 ( \539 , RI2af433cda248_168, \538 );
nor \U$315 ( \540 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$316 ( \541 , RI2af433cda2c0_169, \540 );
nor \U$317 ( \542 , \231 , \232 , \233 , \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$318 ( \543 , RI2af433cda338_170, \542 );
nor \U$319 ( \544 , RI2af433cd5b08_16, \232 , \233 , \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$320 ( \545 , RI2af433cda3b0_171, \544 );
nor \U$321 ( \546 , \231 , RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$322 ( \547 , RI2af433cda428_172, \546 );
nor \U$323 ( \548 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$324 ( \549 , RI2af433cda4a0_173, \548 );
nor \U$325 ( \550 , \231 , \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$326 ( \551 , RI2af433cda518_174, \550 );
nor \U$327 ( \552 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$328 ( \553 , RI2af433cda590_175, \552 );
nor \U$329 ( \554 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$330 ( \555 , RI2af433cda608_176, \554 );
nor \U$331 ( \556 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$332 ( \557 , RI2af433cda680_177, \556 );
nor \U$333 ( \558 , \231 , \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$334 ( \559 , RI2af433cda6f8_178, \558 );
nor \U$335 ( \560 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$336 ( \561 , RI2af433cda770_179, \560 );
nor \U$337 ( \562 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$338 ( \563 , RI2af433cda7e8_180, \562 );
nor \U$339 ( \564 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$340 ( \565 , RI2af433cda860_181, \564 );
nor \U$341 ( \566 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$342 ( \567 , RI2af433cda8d8_182, \566 );
nor \U$343 ( \568 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$344 ( \569 , RI2af433cda950_183, \568 );
nor \U$345 ( \570 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$346 ( \571 , RI2af433cda9c8_184, \570 );
nor \U$347 ( \572 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, \251 , RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$348 ( \573 , RI2af433cdaa40_185, \572 );
nor \U$349 ( \574 , \231 , \232 , \233 , \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$350 ( \575 , RI2af433cdaab8_186, \574 );
nor \U$351 ( \576 , RI2af433cd5b08_16, \232 , \233 , \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$352 ( \577 , RI2af433cdab30_187, \576 );
nor \U$353 ( \578 , \231 , RI2af433cd5a90_15, \233 , \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$354 ( \579 , RI2af433cdaba8_188, \578 );
nor \U$355 ( \580 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$356 ( \581 , RI2af433cdac20_189, \580 );
nor \U$357 ( \582 , \231 , \232 , RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$358 ( \583 , RI2af433cdac98_190, \582 );
nor \U$359 ( \584 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$360 ( \585 , RI2af433cdad10_191, \584 );
nor \U$361 ( \586 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$362 ( \587 , RI2af433cdad88_192, \586 );
nor \U$363 ( \588 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$364 ( \589 , RI2af433cdae00_193, \588 );
nor \U$365 ( \590 , \231 , \232 , \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$366 ( \591 , RI2af433cdae78_194, \590 );
nor \U$367 ( \592 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$368 ( \593 , RI2af433cdaef0_195, \592 );
nor \U$369 ( \594 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$370 ( \595 , RI2af433cdaf68_196, \594 );
nor \U$371 ( \596 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$372 ( \597 , RI2af433cdafe0_197, \596 );
nor \U$373 ( \598 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$374 ( \599 , RI2af433cdb058_198, \598 );
nor \U$375 ( \600 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$376 ( \601 , RI2af433cdb0d0_199, \600 );
nor \U$377 ( \602 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$378 ( \603 , RI2af433cdb148_200, \602 );
nor \U$379 ( \604 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, \250 , RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$380 ( \605 , RI2af433cdb1c0_201, \604 );
nor \U$381 ( \606 , \231 , \232 , \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$382 ( \607 , RI2af433cdb238_202, \606 );
nor \U$383 ( \608 , RI2af433cd5b08_16, \232 , \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$384 ( \609 , RI2af433cdb2b0_203, \608 );
nor \U$385 ( \610 , \231 , RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$386 ( \611 , RI2af433cdb328_204, \610 );
nor \U$387 ( \612 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$388 ( \613 , RI2af433cdb3a0_205, \612 );
nor \U$389 ( \614 , \231 , \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$390 ( \615 , RI2af433cdb418_206, \614 );
nor \U$391 ( \616 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$392 ( \617 , RI2af433cdb490_207, \616 );
nor \U$393 ( \618 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$394 ( \619 , RI2af433cdb508_208, \618 );
or \U$395 ( \620 , \493 , \495 , \497 , \499 , \501 , \503 , \505 , \507 , \509 , \511 , \513 , \515 , \517 , \519 , \521 , \523 , \525 , \527 , \529 , \531 , \533 , \535 , \537 , \539 , \541 , \543 , \545 , \547 , \549 , \551 , \553 , \555 , \557 , \559 , \561 , \563 , \565 , \567 , \569 , \571 , \573 , \575 , \577 , \579 , \581 , \583 , \585 , \587 , \589 , \591 , \593 , \595 , \597 , \599 , \601 , \603 , \605 , \607 , \609 , \611 , \613 , \615 , \617 , \619 );
nor \U$396 ( \621 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, \226 , RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$397 ( \622 , RI2af433cdb580_209, \621 );
nor \U$398 ( \623 , \231 , \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$399 ( \624 , RI2af433cdb5f8_210, \623 );
nor \U$400 ( \625 , RI2af433cd5b08_16, \232 , \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$401 ( \626 , RI2af433cdb670_211, \625 );
nor \U$402 ( \627 , \231 , RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$403 ( \628 , RI2af433cdb6e8_212, \627 );
nor \U$404 ( \629 , RI2af433cd5b08_16, RI2af433cd5a90_15, \233 , RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$405 ( \630 , RI2af433cdb760_213, \629 );
nor \U$406 ( \631 , \231 , \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$407 ( \632 , RI2af433cdb7d8_214, \631 );
nor \U$408 ( \633 , RI2af433cd5b08_16, \232 , RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$409 ( \634 , RI2af433cdb850_215, \633 );
nor \U$410 ( \635 , \231 , RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$411 ( \636 , RI2af433cdb8c8_216, \635 );
nor \U$412 ( \637 , RI2af433cd5b08_16, RI2af433cd5a90_15, RI2af433cd5a18_14, RI2af433cd59a0_13, RI2af433cd5928_12, RI2af433cd58b0_11, RI2af433cd5838_10, RI2af433cd57c0_9, RI2af433cd5748_8, RI2af433cd56d0_7, RI2af433cd5658_6);
and \U$413 ( \638 , RI2af433cdb940_217, \637 );
or \U$414 ( \639 , \622 , \624 , \626 , \628 , \630 , \632 , \634 , \636 , \638 );
or \U$415 ( \640 , \362 , \491 , \620 , \639 );
buf \U$416 ( \641 , RI2af433cd5748_8);
buf \U$417 ( \642 , RI2af433cd56d0_7);
buf \U$418 ( \643 , RI2af433cd5658_6);
buf \U$419 ( \644 , RI2af433cd5838_10);
buf \U$420 ( \645 , RI2af433cd57c0_9);
buf \U$421 ( \646 , RI2af433cd5928_12);
buf \U$422 ( \647 , RI2af433cd58b0_11);
buf \U$423 ( \648 , RI2af433cd59a0_13);
buf \U$424 ( \649 , RI2af433cd5b08_16);
buf \U$425 ( \650 , RI2af433cd5a90_15);
buf \U$426 ( \651 , RI2af433cd5a18_14);
or \U$427 ( \652 , \649 , \650 , \651 );
and \U$428 ( \653 , \648 , \652 );
or \U$429 ( \654 , \646 , \647 , \653 );
and \U$430 ( \655 , \644 , \645 , \654 );
or \U$431 ( \656 , \641 , \642 , \643 , \655 );
buf \U$432 ( \657 , \656 );
_DC r372 ( \658_nR372 , \640 , \657 );
buf \U$433 ( \659 , \658_nR372 );
xor \U$434 ( \660 , RI2af433cc8a70_1, RI2af433cd5478_2);
xor \U$435 ( \661 , RI2af433cd54f0_3, RI2af433cd5568_4);
xor \U$436 ( \662 , \660 , \661 );
xor \U$437 ( \663 , RI2af433cd55e0_5, RI2af433cd5658_6);
xor \U$438 ( \664 , RI2af433cd56d0_7, RI2af433cd5748_8);
xor \U$439 ( \665 , \663 , \664 );
xor \U$440 ( \666 , \662 , \665 );
xor \U$441 ( \667 , RI2af433cd57c0_9, RI2af433cd5838_10);
xor \U$442 ( \668 , RI2af433cd58b0_11, RI2af433cd5928_12);
xor \U$443 ( \669 , \667 , \668 );
xor \U$444 ( \670 , RI2af433cd59a0_13, RI2af433cd5a18_14);
xor \U$445 ( \671 , RI2af433cd5a90_15, RI2af433cd5b08_16);
xor \U$446 ( \672 , \670 , \671 );
xor \U$447 ( \673 , \669 , \672 );
xor \U$448 ( \674 , \666 , \673 );
xor \U$449 ( \675 , RI2af433cd5b80_17, RI2af433cd5bf8_18);
xor \U$450 ( \676 , RI2af433cd5c70_19, RI2af433cd5ce8_20);
xor \U$451 ( \677 , \675 , \676 );
xor \U$452 ( \678 , RI2af433cd5d60_21, RI2af433cd5dd8_22);
xor \U$453 ( \679 , RI2af433cd5e50_23, RI2af433cd5ec8_24);
xor \U$454 ( \680 , \678 , \679 );
xor \U$455 ( \681 , \677 , \680 );
xor \U$456 ( \682 , RI2af433cd5f40_25, RI2af433cd5fb8_26);
xor \U$457 ( \683 , RI2af433cd6030_27, RI2af433cd60a8_28);
xor \U$458 ( \684 , \682 , \683 );
xor \U$459 ( \685 , RI2af433cd6120_29, RI2af433cd6198_30);
xor \U$460 ( \686 , RI2af433cd6210_31, RI2af433cd6288_32);
xor \U$461 ( \687 , \685 , \686 );
xor \U$462 ( \688 , \684 , \687 );
xor \U$463 ( \689 , \681 , \688 );
xor \U$464 ( \690 , RI2af433cd6300_33, RI2af433cd6378_34);
xor \U$465 ( \691 , RI2af433cd63f0_35, RI2af433cd6468_36);
xor \U$466 ( \692 , \690 , \691 );
xor \U$467 ( \693 , RI2af433cd64e0_37, RI2af433cd6558_38);
xor \U$468 ( \694 , RI2af433cd65d0_39, RI2af433cd6648_40);
xor \U$469 ( \695 , \693 , \694 );
xor \U$470 ( \696 , \692 , \695 );
xor \U$471 ( \697 , RI2af433cd66c0_41, RI2af433cd6738_42);
xor \U$472 ( \698 , RI2af433cd67b0_43, RI2af433cd6828_44);
xor \U$473 ( \699 , \697 , \698 );
xor \U$474 ( \700 , RI2af433cd68a0_45, RI2af433cd6918_46);
xor \U$475 ( \701 , RI2af433cd6990_47, RI2af433cd6a08_48);
xor \U$476 ( \702 , \700 , \701 );
xor \U$477 ( \703 , \699 , \702 );
xor \U$478 ( \704 , \696 , \703 );
xor \U$479 ( \705 , \689 , \704 );
xor \U$480 ( \706 , RI2af433cd6a80_49, RI2af433cd6af8_50);
xor \U$481 ( \707 , RI2af433cd6b70_51, RI2af433cd6be8_52);
xor \U$482 ( \708 , \706 , \707 );
xor \U$483 ( \709 , RI2af433cd6c60_53, RI2af433cd6cd8_54);
xor \U$484 ( \710 , RI2af433cd6d50_55, RI2af433cd6dc8_56);
xor \U$485 ( \711 , \709 , \710 );
xor \U$486 ( \712 , \708 , \711 );
xor \U$487 ( \713 , RI2af433cd6e40_57, RI2af433cd6eb8_58);
xor \U$488 ( \714 , RI2af433cd6f30_59, RI2af433cd6fa8_60);
xor \U$489 ( \715 , \713 , \714 );
xor \U$490 ( \716 , RI2af433cd7020_61, RI2af433cd7098_62);
xor \U$491 ( \717 , RI2af433cd7110_63, RI2af433cd7188_64);
xor \U$492 ( \718 , \716 , \717 );
xor \U$493 ( \719 , \715 , \718 );
xor \U$494 ( \720 , \712 , \719 );
xor \U$495 ( \721 , RI2af433cd7200_65, RI2af433cd7278_66);
xor \U$496 ( \722 , RI2af433cd72f0_67, RI2af433cd7368_68);
xor \U$497 ( \723 , \721 , \722 );
xor \U$498 ( \724 , RI2af433cd73e0_69, RI2af433cd7458_70);
xor \U$499 ( \725 , RI2af433cd74d0_71, RI2af433cd7548_72);
xor \U$500 ( \726 , \724 , \725 );
xor \U$501 ( \727 , \723 , \726 );
xor \U$502 ( \728 , RI2af433cd75c0_73, RI2af433cd7638_74);
xor \U$503 ( \729 , RI2af433cd76b0_75, RI2af433cd7728_76);
xor \U$504 ( \730 , \728 , \729 );
xor \U$505 ( \731 , RI2af433cd77a0_77, RI2af433cd7818_78);
xor \U$506 ( \732 , RI2af433cd7890_79, RI2af433cd7908_80);
xor \U$507 ( \733 , \731 , \732 );
xor \U$508 ( \734 , \730 , \733 );
xor \U$509 ( \735 , \727 , \734 );
xor \U$510 ( \736 , \720 , \735 );
xor \U$511 ( \737 , \705 , \736 );
xor \U$512 ( \738 , RI2af433cd7980_81, RI2af433cd79f8_82);
xor \U$513 ( \739 , RI2af433cd7a70_83, RI2af433cd7ae8_84);
xor \U$514 ( \740 , \738 , \739 );
xor \U$515 ( \741 , RI2af433cd7b60_85, RI2af433cd7bd8_86);
xor \U$516 ( \742 , RI2af433cd7c50_87, RI2af433cd7cc8_88);
xor \U$517 ( \743 , \741 , \742 );
xor \U$518 ( \744 , \740 , \743 );
xor \U$519 ( \745 , RI2af433cd7d40_89, RI2af433cd7db8_90);
xor \U$520 ( \746 , RI2af433cd7e30_91, RI2af433cd7ea8_92);
xor \U$521 ( \747 , \745 , \746 );
xor \U$522 ( \748 , RI2af433cd7f20_93, RI2af433cd7f98_94);
xor \U$523 ( \749 , RI2af433cd8010_95, RI2af433cd8088_96);
xor \U$524 ( \750 , \748 , \749 );
xor \U$525 ( \751 , \747 , \750 );
xor \U$526 ( \752 , \744 , \751 );
xor \U$527 ( \753 , RI2af433cd8100_97, RI2af433cd8178_98);
xor \U$528 ( \754 , RI2af433cd81f0_99, RI2af433cd8268_100);
xor \U$529 ( \755 , \753 , \754 );
xor \U$530 ( \756 , RI2af433cd82e0_101, RI2af433cd8358_102);
xor \U$531 ( \757 , RI2af433cd83d0_103, RI2af433cd8448_104);
xor \U$532 ( \758 , \756 , \757 );
xor \U$533 ( \759 , \755 , \758 );
xor \U$534 ( \760 , RI2af433cd84c0_105, RI2af433cd8538_106);
xor \U$535 ( \761 , RI2af433cd85b0_107, RI2af433cd8628_108);
xor \U$536 ( \762 , \760 , \761 );
xor \U$537 ( \763 , RI2af433cd86a0_109, RI2af433cd8718_110);
xor \U$538 ( \764 , RI2af433cd8790_111, RI2af433cd8808_112);
xor \U$539 ( \765 , \763 , \764 );
xor \U$540 ( \766 , \762 , \765 );
xor \U$541 ( \767 , \759 , \766 );
xor \U$542 ( \768 , \752 , \767 );
xor \U$543 ( \769 , RI2af433cd8880_113, RI2af433cd88f8_114);
xor \U$544 ( \770 , RI2af433cd8970_115, RI2af433cd89e8_116);
xor \U$545 ( \771 , \769 , \770 );
xor \U$546 ( \772 , RI2af433cd8a60_117, RI2af433cd8ad8_118);
xor \U$547 ( \773 , RI2af433cd8b50_119, RI2af433cd8bc8_120);
xor \U$548 ( \774 , \772 , \773 );
xor \U$549 ( \775 , \771 , \774 );
xor \U$550 ( \776 , RI2af433cd8c40_121, RI2af433cd8cb8_122);
xor \U$551 ( \777 , RI2af433cd8d30_123, RI2af433cd8da8_124);
xor \U$552 ( \778 , \776 , \777 );
xor \U$553 ( \779 , RI2af433cd8e20_125, RI2af433cd8e98_126);
xor \U$554 ( \780 , RI2af433cd8f10_127, RI2af433cd8f88_128);
xor \U$555 ( \781 , \779 , \780 );
xor \U$556 ( \782 , \778 , \781 );
xor \U$557 ( \783 , \775 , \782 );
xor \U$558 ( \784 , RI2af433cd9000_129, RI2af433cd9078_130);
xor \U$559 ( \785 , RI2af433cd90f0_131, RI2af433cd9168_132);
xor \U$560 ( \786 , \784 , \785 );
xor \U$561 ( \787 , RI2af433cd91e0_133, RI2af433cd9258_134);
xor \U$562 ( \788 , RI2af433cd92d0_135, RI2af433cd9348_136);
xor \U$563 ( \789 , \787 , \788 );
xor \U$564 ( \790 , \786 , \789 );
xor \U$565 ( \791 , RI2af433cd93c0_137, RI2af433cd9438_138);
xor \U$566 ( \792 , RI2af433cd94b0_139, RI2af433cd9528_140);
xor \U$567 ( \793 , \791 , \792 );
xor \U$568 ( \794 , RI2af433cd95a0_141, RI2af433cd9618_142);
xor \U$569 ( \795 , RI2af433cd9690_143, RI2af433cd9708_144);
xor \U$570 ( \796 , \794 , \795 );
xor \U$571 ( \797 , \793 , \796 );
xor \U$572 ( \798 , \790 , \797 );
xor \U$573 ( \799 , \783 , \798 );
xor \U$574 ( \800 , \768 , \799 );
xor \U$575 ( \801 , \737 , \800 );
xor \U$576 ( \802 , RI2af433cd9780_145, RI2af433cd97f8_146);
xor \U$577 ( \803 , RI2af433cd9870_147, RI2af433cd98e8_148);
xor \U$578 ( \804 , \802 , \803 );
xor \U$579 ( \805 , RI2af433cd9960_149, RI2af433cd99d8_150);
xor \U$580 ( \806 , RI2af433cd9a50_151, RI2af433cd9ac8_152);
xor \U$581 ( \807 , \805 , \806 );
xor \U$582 ( \808 , \804 , \807 );
xor \U$583 ( \809 , RI2af433cd9b40_153, RI2af433cd9bb8_154);
xor \U$584 ( \810 , RI2af433cd9c30_155, RI2af433cd9ca8_156);
xor \U$585 ( \811 , \809 , \810 );
xor \U$586 ( \812 , RI2af433cd9d20_157, RI2af433cd9d98_158);
xor \U$587 ( \813 , RI2af433cd9e10_159, RI2af433cd9e88_160);
xor \U$588 ( \814 , \812 , \813 );
xor \U$589 ( \815 , \811 , \814 );
xor \U$590 ( \816 , \808 , \815 );
xor \U$591 ( \817 , RI2af433cd9f00_161, RI2af433cd9f78_162);
xor \U$592 ( \818 , RI2af433cd9ff0_163, RI2af433cda068_164);
xor \U$593 ( \819 , \817 , \818 );
xor \U$594 ( \820 , RI2af433cda0e0_165, RI2af433cda158_166);
xor \U$595 ( \821 , RI2af433cda1d0_167, RI2af433cda248_168);
xor \U$596 ( \822 , \820 , \821 );
xor \U$597 ( \823 , \819 , \822 );
xor \U$598 ( \824 , RI2af433cda2c0_169, RI2af433cda338_170);
xor \U$599 ( \825 , RI2af433cda3b0_171, RI2af433cda428_172);
xor \U$600 ( \826 , \824 , \825 );
xor \U$601 ( \827 , RI2af433cda4a0_173, RI2af433cda518_174);
xor \U$602 ( \828 , RI2af433cda590_175, RI2af433cda608_176);
xor \U$603 ( \829 , \827 , \828 );
xor \U$604 ( \830 , \826 , \829 );
xor \U$605 ( \831 , \823 , \830 );
xor \U$606 ( \832 , \816 , \831 );
xor \U$607 ( \833 , RI2af433cda680_177, RI2af433cda6f8_178);
xor \U$608 ( \834 , RI2af433cda770_179, RI2af433cda7e8_180);
xor \U$609 ( \835 , \833 , \834 );
xor \U$610 ( \836 , RI2af433cda860_181, RI2af433cda8d8_182);
xor \U$611 ( \837 , RI2af433cda950_183, RI2af433cda9c8_184);
xor \U$612 ( \838 , \836 , \837 );
xor \U$613 ( \839 , \835 , \838 );
xor \U$614 ( \840 , RI2af433cdaa40_185, RI2af433cdaab8_186);
xor \U$615 ( \841 , RI2af433cdab30_187, RI2af433cdaba8_188);
xor \U$616 ( \842 , \840 , \841 );
xor \U$617 ( \843 , RI2af433cdac20_189, RI2af433cdac98_190);
xor \U$618 ( \844 , RI2af433cdad10_191, RI2af433cdad88_192);
xor \U$619 ( \845 , \843 , \844 );
xor \U$620 ( \846 , \842 , \845 );
xor \U$621 ( \847 , \839 , \846 );
xor \U$622 ( \848 , RI2af433cdae00_193, RI2af433cdae78_194);
xor \U$623 ( \849 , RI2af433cdaef0_195, RI2af433cdaf68_196);
xor \U$624 ( \850 , \848 , \849 );
xor \U$625 ( \851 , RI2af433cdafe0_197, RI2af433cdb058_198);
xor \U$626 ( \852 , RI2af433cdb0d0_199, RI2af433cdb148_200);
xor \U$627 ( \853 , \851 , \852 );
xor \U$628 ( \854 , \850 , \853 );
xor \U$629 ( \855 , RI2af433cdb1c0_201, RI2af433cdb238_202);
xor \U$630 ( \856 , RI2af433cdb2b0_203, RI2af433cdb328_204);
xor \U$631 ( \857 , \855 , \856 );
xor \U$632 ( \858 , RI2af433cdb3a0_205, RI2af433cdb418_206);
xor \U$633 ( \859 , RI2af433cdb490_207, RI2af433cdb508_208);
xor \U$634 ( \860 , \858 , \859 );
xor \U$635 ( \861 , \857 , \860 );
xor \U$636 ( \862 , \854 , \861 );
xor \U$637 ( \863 , \847 , \862 );
xor \U$638 ( \864 , \832 , \863 );
xor \U$639 ( \865 , RI2af433cdb580_209, RI2af433cdb5f8_210);
xor \U$640 ( \866 , RI2af433cdb670_211, RI2af433cdb6e8_212);
xor \U$641 ( \867 , \865 , \866 );
xor \U$642 ( \868 , RI2af433cdb760_213, RI2af433cdb7d8_214);
xor \U$643 ( \869 , RI2af433cdb850_215, RI2af433cdb8c8_216);
xor \U$644 ( \870 , \868 , \869 );
xor \U$645 ( \871 , \867 , \870 );
xor \U$646 ( \872 , \871 , RI2af433cdb940_217);
xor \U$647 ( \873 , \864 , \872 );
xor \U$648 ( \874 , \801 , \873 );
_DC r1bf ( \875_nR1bf , 1'b0 , 1'b1 );
and \U$651 ( \876 , \874 , \875_nR1bf );
and \U$652 ( \877 , \674 , \876 );
buf \U$653 ( \878 , \877 );
endmodule

